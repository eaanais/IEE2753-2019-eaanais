* NGSPICE file created from FIR.ext - technology: scmos

* Black-box entry subcircuit for FILL abstract view
.subckt FILL gnd vdd
.ends

* Black-box entry subcircuit for OAI21X1 abstract view
.subckt OAI21X1 A B C gnd Y vdd
.ends

* Black-box entry subcircuit for NOR2X1 abstract view
.subckt NOR2X1 A B gnd Y vdd
.ends

* Black-box entry subcircuit for CLKBUF1 abstract view
.subckt CLKBUF1 A gnd Y vdd
.ends

* Black-box entry subcircuit for NAND2X1 abstract view
.subckt NAND2X1 A B gnd Y vdd
.ends

* Black-box entry subcircuit for NAND3X1 abstract view
.subckt NAND3X1 A B C gnd Y vdd
.ends

* Black-box entry subcircuit for INVX1 abstract view
.subckt INVX1 A gnd Y vdd
.ends

* Black-box entry subcircuit for DFFPOSX1 abstract view
.subckt DFFPOSX1 Q CLK D gnd vdd
.ends

* Black-box entry subcircuit for AOI21X1 abstract view
.subckt AOI21X1 A B C gnd Y vdd
.ends

* Black-box entry subcircuit for BUFX2 abstract view
.subckt BUFX2 A gnd Y vdd
.ends

* Black-box entry subcircuit for OAI22X1 abstract view
.subckt OAI22X1 A B C D gnd Y vdd
.ends

* Black-box entry subcircuit for DFFSR abstract view
.subckt DFFSR Q CLK R S D gnd vdd
.ends

* Black-box entry subcircuit for XOR2X1 abstract view
.subckt XOR2X1 A B gnd Y vdd
.ends

* Black-box entry subcircuit for OR2X2 abstract view
.subckt OR2X2 A B gnd Y vdd
.ends

* Black-box entry subcircuit for NOR3X1 abstract view
.subckt NOR3X1 A B C gnd Y vdd
.ends

* Black-box entry subcircuit for AND2X2 abstract view
.subckt AND2X2 A B gnd Y vdd
.ends

* Black-box entry subcircuit for AOI22X1 abstract view
.subckt AOI22X1 A B C D gnd Y vdd
.ends

* Black-box entry subcircuit for XNOR2X1 abstract view
.subckt XNOR2X1 A B gnd Y vdd
.ends

.subckt FIR clk rst din[0] din[1] din[2] din[3] din[4] din[5] din[6] din[7] dout[0]
+ dout[1] dout[2] dout[3] dout[4] dout[5] dout[6] dout[7]
XFILL_8_CLKBUF1_8 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_2_DFFSR_25 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_22_DFFSR_143 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_19_DFFSR_18 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_12_DFFSR_146 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_2_INVX1_297 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_1_NOR2X1_6 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_19_CLKBUF1_11 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_8_DFFSR_140 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_43_DFFSR_75 INVX1_4/gnd DFFSR_51/S FILL
XFILL_18_CLKBUF1_14 BUFX2_43/A DFFSR_23/S FILL
XFILL_49_DFFSR_171 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_5_OAI21X1_256 INVX1_2/gnd DFFSR_51/S FILL
XFILL_40_2_0 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_39_DFFSR_174 BUFX2_43/A DFFSR_97/S FILL
XFILL_17_CLKBUF1_17 INVX1_94/gnd DFFSR_25/S FILL
XFILL_1_INVX1_117 INVX1_4/gnd DFFSR_51/S FILL
XFILL_7_NAND3X1_106 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_27_DFFSR_25 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_29_DFFSR_177 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_16_CLKBUF1_20 INVX1_4/gnd DFFSR_51/S FILL
XFILL_16_DFFSR_65 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_38_4_1 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_15_CLKBUF1_23 INVX1_89/gnd DFFSR_2/S FILL
XFILL_11_DFFPOSX1_10 INVX1_8/gnd DFFSR_5/S FILL
XFILL_19_DFFSR_180 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_6_OAI21X1_190 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_3_XOR2X1_2 BUFX2_8/gnd DFFSR_10/S FILL
XOAI21X1_226 OR2X2_2/A AOI22X1_13/Y OAI21X1_223/C BUFX2_6/gnd NAND3X1_71/C DFFSR_91/S
+ OAI21X1
XFILL_6_OAI21X1_7 INVX1_8/gnd DFFSR_5/S FILL
XFILL_23_DFFSR_4 INVX1_4/gnd DFFSR_4/S FILL
XFILL_7_OAI21X1_124 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_42_DFFSR_101 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_7_DFFSR_79 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_5_DFFSR_177 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_24_DFFSR_72 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_35_DFFSR_32 INVX1_2/gnd DFFSR_1/S FILL
XFILL_32_DFFSR_104 INVX1_4/gnd DFFSR_4/S FILL
XFILL_22_DFFSR_107 BUFX2_36/A DFFSR_8/S FILL
XFILL_1_DFFPOSX1_21 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_12_DFFSR_110 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_6_BUFX2_17 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_2_INVX1_261 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_5_OAI21X1_220 BUFX2_43/A DFFSR_97/S FILL
XFILL_43_DFFSR_39 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_32_DFFSR_79 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_8_DFFSR_104 INVX1_4/gnd DFFSR_4/S FILL
XFILL_49_DFFSR_135 BUFX2_43/A DFFSR_97/S FILL
XFILL_16_DFFSR_29 INVX1_4/gnd DFFSR_4/S FILL
XFILL_39_DFFSR_138 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_29_DFFSR_141 INVX1_94/gnd DFFSR_25/S FILL
XFILL_46_1_2 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_6_OAI21X1_154 BUFX2_37/A DFFSR_8/S FILL
XFILL_19_DFFSR_144 INVX1_8/gnd DFFSR_5/S FILL
XFILL_5_CLKBUF1_9 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_20_DFFPOSX1_29 DFFSR_1/gnd DFFSR_9/S FILL
XNOR2X1_26 NOR2X1_26/A NOR2X1_26/B DFFSR_73/gnd NOR2X1_26/Y DFFSR_11/S NOR2X1
XFILL_4_NOR2X1_23 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_40_DFFSR_86 DFFSR_1/gnd DFFSR_9/S FILL
XOAI21X1_190 INVX1_214/Y INVX1_231/Y NAND2X1_190/Y BUFX2_5/gnd OAI21X1_190/Y DFFSR_6/S
+ OAI21X1
XFILL_6_NAND2X1_268 BUFX2_37/A DFFSR_8/S FILL
XFILL_3_INVX1_405 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_13_DFFSR_76 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_7_DFFSR_43 INVX1_94/gnd DFFSR_25/S FILL
XFILL_5_DFFSR_141 INVX1_94/gnd DFFSR_25/S FILL
XFILL_24_DFFSR_36 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_46_DFFSR_172 BUFX2_37/A DFFSR_8/S FILL
XFILL_14_0_0 BUFX2_37/A DFFSR_8/S FILL
XFILL_36_DFFSR_175 INVX1_23/gnd DFFSR_91/S FILL
XFILL_4_OAI21X1_250 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_26_DFFSR_178 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_16_DFFSR_181 INVX1_23/gnd DFFSR_186/S FILL
XFILL_12_2_1 BUFX2_36/A DFFSR_6/S FILL
XFILL_2_INVX1_225 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_48_DFFSR_93 INVX1_2/gnd DFFSR_51/S FILL
XFILL_6_NAND3X1_100 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_10_4_2 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_9_AND2X2_2 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_7_CLKBUF1_11 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_21_DFFSR_83 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_4_INVX1_37 INVX1_94/gnd DFFSR_52/S FILL
XFILL_32_DFFSR_43 INVX1_94/gnd DFFSR_25/S FILL
XFILL_4_DFFSR_90 INVX1_2/gnd DFFSR_1/S FILL
XFILL_6_CLKBUF1_14 BUFX2_43/A DFFSR_23/S FILL
XFILL_3_OAI21X1_8 BUFX2_36/A DFFSR_6/S FILL
XFILL_5_OAI21X1_184 BUFX2_19/gnd DFFSR_52/S FILL
XCLKBUF1_14 clk BUFX2_43/A CLKBUF1_14/Y DFFSR_23/S CLKBUF1
XFILL_5_CLKBUF1_17 INVX1_94/gnd DFFSR_25/S FILL
XFILL_39_DFFSR_102 INVX1_8/gnd DFFSR_7/S FILL
XFILL_3_BUFX2_28 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_29_DFFSR_105 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_5_4 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_2_DFFSR_178 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_4_CLKBUF1_20 INVX1_4/gnd DFFSR_51/S FILL
XFILL_3_CLKBUF1_23 INVX1_89/gnd DFFSR_2/S FILL
XFILL_19_DFFSR_108 INVX1_89/gnd DFFSR_2/S FILL
XFILL_6_OAI21X1_118 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_1_INVX1_84 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_40_DFFSR_50 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_0_DFFPOSX1_15 BUFX2_35/A DFFSR_14/S FILL
XOAI21X1_154 DFFSR_8/S INVX1_182/Y OAI21X1_154/C BUFX2_37/A DFFSR_154/D DFFSR_8/S
+ OAI21X1
XFILL_29_DFFSR_90 INVX1_2/gnd DFFSR_1/S FILL
XFILL_6_NAND2X1_232 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_3_INVX1_369 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_5_DFFSR_105 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_13_DFFSR_40 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_5_NAND3X1_130 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_46_DFFSR_136 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_4_OAI21X1_214 BUFX2_35/A DFFSR_97/S FILL
XNAND2X1_268 DFFSR_8/S DFFSR_165/Q BUFX2_37/A NAND2X1_268/Y DFFSR_8/S NAND2X1
XFILL_36_DFFSR_139 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_2_INVX1_189 BUFX2_35/A DFFSR_14/S FILL
XFILL_26_DFFSR_142 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_35_DFFSR_7 INVX1_8/gnd DFFSR_7/S FILL
XFILL_16_DFFSR_145 INVX1_23/gnd DFFSR_186/S FILL
XFILL_37_DFFSR_97 BUFX2_35/A DFFSR_97/S FILL
XFILL_48_DFFSR_57 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_5_OAI21X1_148 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_19_DFFPOSX1_23 INVX1_23/gnd DFFSR_91/S FILL
XFILL_4_DFFSR_54 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_1_NOR2X1_24 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_21_DFFSR_47 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_10_DFFSR_87 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_0_0_2 DFFSR_89/gnd DFFSR_92/S FILL
XNAND3X1_100 NAND3X1_98/B NAND3X1_98/C OR2X2_2/Y BUFX2_6/gnd AOI21X1_31/A DFFSR_14/S
+ NAND3X1
XFILL_2_DFFSR_142 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_0_INVX1_406 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_43_DFFSR_173 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_5_NAND2X1_262 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_33_DFFSR_176 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_23_DFFSR_179 INVX1_2/gnd DFFSR_1/S FILL
XFILL_40_DFFSR_14 BUFX2_35/A DFFSR_14/S FILL
XFILL_29_DFFSR_54 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_18_DFFSR_94 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_1_INVX1_48 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_13_DFFSR_182 INVX1_89/gnd DFFSR_36/S FILL
XFILL_47_2_0 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_3_OAI21X1_244 DFFSR_3/gnd DFFSR_4/S FILL
XOAI21X1_118 BUFX2_17/Y INVX1_133/Y OAI21X1_118/C DFFSR_73/gnd DFFSR_118/D DFFSR_11/S
+ OAI21X1
XFILL_6_NAND2X1_196 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_3_INVX1_333 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_46_DFFSR_100 INVX1_23/gnd DFFSR_186/S FILL
XFILL_0_BUFX2_39 BUFX2_43/A DFFSR_97/S FILL
XFILL_0_OAI21X1_9 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_45_4_1 INVX1_2/gnd DFFSR_1/S FILL
XNAND2X1_232 AND2X2_13/B AND2X2_13/A BUFX2_7/gnd NAND3X1_110/B DFFSR_54/S NAND2X1
XFILL_36_DFFSR_103 INVX1_8/gnd DFFSR_7/S FILL
XFILL_9_DFFSR_176 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_4_OAI21X1_178 INVX1_94/gnd DFFSR_25/S FILL
XFILL_26_DFFSR_106 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_16_DFFSR_109 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_37_DFFSR_61 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_2_INVX1_153 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_48_DFFSR_21 INVX1_2/gnd DFFSR_1/S FILL
XFILL_4_DFFSR_18 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_21_DFFSR_11 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_10_DFFSR_51 INVX1_2/gnd DFFSR_51/S FILL
XFILL_5_OAI21X1_112 INVX1_4/gnd DFFSR_4/S FILL
XFILL_0_INVX1_370 BUFX2_36/A DFFSR_8/S FILL
XFILL_2_DFFSR_106 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_45_DFFSR_68 BUFX2_35/A DFFSR_14/S FILL
XFILL_11_5_0 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_5_NAND2X1_226 BUFX2_36/A DFFSR_6/S FILL
XFILL_43_DFFSR_137 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_22_DFFSR_1 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_33_DFFSR_140 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_9_CLKBUF1_8 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_23_DFFSR_143 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_1_INVX1_12 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_4_NAND3X1_124 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_1_DFFSR_65 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_13_DFFSR_146 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_6_BUFX2_2 BUFX2_43/A DFFSR_23/S FILL
XFILL_29_DFFSR_18 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_18_DFFSR_58 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_3_OAI21X1_208 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_6_NAND2X1_160 INVX1_8/gnd DFFSR_5/S FILL
XFILL_3_INVX1_297 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_9_DFFSR_140 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_18_DFFPOSX1_17 BUFX2_37/A DFFSR_8/S FILL
XNAND2X1_196 NAND2X1_195/B AND2X2_7/Y BUFX2_7/gnd NAND3X1_22/C DFFSR_54/S NAND2X1
XFILL_50_DFFSR_171 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_4_OAI21X1_142 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_40_DFFSR_174 BUFX2_43/A DFFSR_97/S FILL
XFILL_2_INVX1_117 INVX1_4/gnd DFFSR_51/S FILL
XFILL_37_DFFSR_25 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_18_DFFPOSX1_2 INVX1_89/gnd DFFSR_36/S FILL
XFILL_30_DFFSR_177 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_9_DFFSR_72 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_26_DFFSR_65 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_17_DFFPOSX1_5 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_16_DFFPOSX1_8 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_4_NAND2X1_256 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_10_DFFSR_15 INVX1_8/gnd DFFSR_7/S FILL
XFILL_20_DFFSR_180 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_10_DFFSR_183 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_0_INVX1_334 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_21_0_0 INVX1_94/gnd DFFSR_25/S FILL
XFILL_7_OAI21X1_7 INVX1_8/gnd DFFSR_5/S FILL
XFILL_2_OAI21X1_238 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_8_DFFPOSX1_28 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_43_DFFSR_101 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_5_NAND2X1_190 BUFX2_35/A DFFSR_97/S FILL
XFILL_19_2_1 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_6_DFFSR_177 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_34_DFFSR_72 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_45_DFFSR_32 INVX1_2/gnd DFFSR_1/S FILL
XFILL_33_DFFSR_104 INVX1_4/gnd DFFSR_4/S FILL
XFILL_1_1_0 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_23_DFFSR_107 BUFX2_36/A DFFSR_8/S FILL
XFILL_17_4_2 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_18_DFFSR_22 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_1_DFFSR_29 INVX1_4/gnd DFFSR_4/S FILL
XFILL_3_OAI21X1_172 BUFX2_36/A DFFSR_6/S FILL
XFILL_10_OAI22X1_3 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_6_NAND2X1_124 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_13_DFFSR_110 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_3_INVX1_261 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_42_DFFSR_79 DFFSR_79/gnd DFFSR_36/S FILL
XNAND2X1_160 NAND3X1_1/C BUFX2_3/Y INVX1_8/gnd NAND2X1_160/Y DFFSR_5/S NAND2X1
XFILL_9_DFFSR_104 INVX1_4/gnd DFFSR_4/S FILL
XFILL_50_DFFSR_135 BUFX2_43/A DFFSR_97/S FILL
XFILL_3_NAND2X1_286 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_4_OAI21X1_106 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_15_DFFSR_69 BUFX2_43/A DFFSR_23/S FILL
XFILL_9_DFFSR_36 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_26_DFFSR_29 INVX1_4/gnd DFFSR_4/S FILL
XFILL_40_DFFSR_138 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_30_DFFSR_141 INVX1_94/gnd DFFSR_25/S FILL
XFILL_4_NAND2X1_220 BUFX2_35/A DFFSR_14/S FILL
XFILL_20_DFFSR_144 INVX1_8/gnd DFFSR_5/S FILL
XFILL_6_CLKBUF1_9 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_2_XOR2X1_6 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_10_DFFSR_147 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_13_DFFSR_8 BUFX2_36/A DFFSR_8/S FILL
XFILL_3_NAND3X1_118 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_5_NOR2X1_23 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_50_DFFSR_86 DFFSR_1/gnd DFFSR_9/S FILL
XINVX1_408 NAND2X1_3/B DFFSR_9/gnd INVX1_408/Y DFFSR_9/S INVX1
XFILL_0_INVX1_298 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_2_OAI21X1_202 BUFX2_35/A DFFSR_14/S FILL
XFILL_5_NAND2X1_154 BUFX2_37/A DFFSR_8/S FILL
XFILL_23_DFFSR_76 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_6_DFFSR_83 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_6_DFFSR_141 INVX1_94/gnd DFFSR_25/S FILL
XFILL_34_DFFSR_36 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_47_DFFSR_172 BUFX2_37/A DFFSR_8/S FILL
XFILL_37_DFFSR_175 INVX1_23/gnd DFFSR_91/S FILL
XFILL_5_BUFX2_21 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_27_DFFSR_178 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_17_DFFPOSX1_11 INVX1_4/gnd DFFSR_4/S FILL
XFILL_9_OAI21X1_97 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_3_INVX1_225 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_3_OAI21X1_136 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_17_DFFSR_181 INVX1_23/gnd DFFSR_186/S FILL
XFILL_7_0_2 BUFX2_35/A DFFSR_97/S FILL
XFILL_34_DFFSR_4 INVX1_4/gnd DFFSR_4/S FILL
XFILL_3_INVX1_77 BUFX2_37/A DFFSR_81/S FILL
XFILL_31_DFFSR_83 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_42_DFFSR_43 INVX1_94/gnd DFFSR_25/S FILL
XFILL_9_AOI21X1_13 INVX1_8/gnd DFFSR_7/S FILL
XFILL_4_OAI21X1_8 BUFX2_36/A DFFSR_6/S FILL
XNAND2X1_124 BUFX2_23/Y INVX1_131/A DFFSR_79/gnd NAND2X1_124/Y DFFSR_36/S NAND2X1
XFILL_3_NAND2X1_250 INVX1_8/gnd DFFSR_5/S FILL
XFILL_8_AOI21X1_16 BUFX2_43/A DFFSR_23/S FILL
XFILL_40_DFFSR_102 INVX1_8/gnd DFFSR_7/S FILL
XFILL_30_DFFSR_105 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_9_1 BUFX2_43/A DFFSR_97/S FILL
XFILL_7_AOI21X1_19 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_15_DFFSR_33 INVX1_94/gnd DFFSR_52/S FILL
XFILL_6_DFFPOSX1_2 INVX1_89/gnd DFFSR_36/S FILL
XFILL_3_DFFSR_178 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_1_OAI21X1_232 BUFX2_35/A DFFSR_97/S FILL
XFILL_6_AOI21X1_22 BUFX2_43/A DFFSR_97/S FILL
XDFFPOSX1_2 NAND3X1_1/C CLKBUF1_10/Y XOR2X1_1/Y INVX1_89/gnd DFFSR_36/S DFFPOSX1
XFILL_20_DFFSR_108 INVX1_89/gnd DFFSR_2/S FILL
XFILL_5_DFFPOSX1_5 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_5_AOI21X1_25 BUFX2_43/A DFFSR_97/S FILL
XAOI21X1_22 NAND3X1_37/Y NAND3X1_47/B OAI22X1_2/Y BUFX2_43/A AOI21X1_22/Y DFFSR_97/S
+ AOI21X1
XFILL_4_NAND2X1_184 BUFX2_37/A DFFSR_8/S FILL
XFILL_4_DFFPOSX1_8 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_7_DFFPOSX1_22 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_4_AOI21X1_28 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_10_DFFSR_111 INVX1_8/gnd DFFSR_5/S FILL
XFILL_3_AOI21X1_31 INVX1_23/gnd DFFSR_186/S FILL
XFILL_39_DFFSR_90 INVX1_2/gnd DFFSR_1/S FILL
XFILL_0_INVX1_262 INVX1_2/gnd DFFSR_1/S FILL
XFILL_50_DFFSR_50 DFFSR_73/gnd DFFSR_11/S FILL
XINVX1_372 INVX1_97/A DFFSR_73/gnd INVX1_372/Y DFFSR_57/S INVX1
XFILL_2_AOI21X1_34 INVX1_94/gnd DFFSR_25/S FILL
XFILL_2_OAI21X1_166 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_6_DFFSR_105 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_1_AOI21X1_37 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_6_DFFSR_47 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_23_DFFSR_40 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_12_DFFSR_80 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_5_NAND2X1_118 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_47_DFFSR_136 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_0_AOI21X1_40 DFFSR_3/gnd DFFSR_4/S FILL
XBUFX2_25 INVX1_1/Y BUFX2_5/gnd BUFX2_25/Y DFFSR_6/S BUFX2
XFILL_37_DFFSR_139 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_3_OAI21X1_100 INVX1_23/gnd DFFSR_91/S FILL
XFILL_26_DFFPOSX1_30 BUFX2_43/A DFFSR_97/S FILL
XFILL_14_7 BUFX2_36/A DFFSR_8/S FILL
XFILL_9_OAI21X1_61 BUFX2_36/A DFFSR_8/S FILL
XFILL_27_DFFSR_142 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_2_NAND2X1_280 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_17_DFFSR_145 INVX1_23/gnd DFFSR_186/S FILL
XFILL_3_INVX1_189 BUFX2_35/A DFFSR_14/S FILL
XFILL_47_DFFSR_97 BUFX2_35/A DFFSR_97/S FILL
XFILL_8_OAI21X1_64 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_8_AND2X2_6 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_6_NAND2X1_85 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_7_OAI21X1_67 INVX1_2/gnd DFFSR_1/S FILL
XFILL_18_5_0 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_2_NOR2X1_24 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_3_INVX1_41 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_0_OAI21X1_262 INVX1_89/gnd DFFSR_36/S FILL
XFILL_31_DFFSR_47 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_20_DFFSR_87 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_5_NAND2X1_88 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_3_DFFSR_94 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_3_NAND2X1_214 BUFX2_35/A DFFSR_97/S FILL
XNAND2X1_85 BUFX2_23/Y INVX1_87/A DFFSR_79/gnd OAI21X1_85/C DFFSR_45/S NAND2X1
XFILL_6_OAI21X1_70 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_4_NAND2X1_91 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_2_NAND3X1_112 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_1_INVX1_406 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_5_OAI21X1_73 DFFSR_73/gnd DFFSR_11/S FILL
XOAI21X1_70 BUFX2_17/Y INVX1_79/Y NAND2X1_70/Y DFFSR_73/gnd DFFSR_70/D DFFSR_57/S
+ OAI21X1
XFILL_44_DFFSR_173 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_3_DFFSR_142 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_4_OAI21X1_76 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_2_BUFX2_32 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_3_NAND2X1_94 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_4_NAND2X1_148 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_2_NAND2X1_97 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_1_OAI21X1_196 INVX1_94/gnd DFFSR_25/S FILL
XFILL_3_OAI21X1_79 INVX1_89/gnd DFFSR_36/S FILL
XFILL_1_DFFSR_7 INVX1_8/gnd DFFSR_7/S FILL
XFILL_34_DFFSR_176 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_2_OAI21X1_82 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_0_INVX1_226 BUFX2_35/A DFFSR_14/S FILL
XFILL_50_DFFSR_14 BUFX2_35/A DFFSR_14/S FILL
XINVX1_336 DFFSR_97/Q BUFX2_5/gnd INVX1_336/Y DFFSR_6/S INVX1
XFILL_39_DFFSR_54 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_1_OAI21X1_85 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_0_INVX1_88 INVX1_2/gnd DFFSR_1/S FILL
XFILL_24_DFFSR_179 INVX1_2/gnd DFFSR_1/S FILL
XFILL_28_DFFSR_94 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_14_DFFSR_182 INVX1_89/gnd DFFSR_36/S FILL
XFILL_0_OAI21X1_88 INVX1_4/gnd DFFSR_4/S FILL
XFILL_12_DFFSR_44 BUFX2_8/gnd DFFSR_10/S FILL
XBUFX2_3 BUFX2_2/A DFFSR_5/gnd BUFX2_3/Y DFFSR_2/S BUFX2
XFILL_4_INVX1_333 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_2_OAI21X1_130 INVX1_4/gnd DFFSR_4/S FILL
XFILL_6_DFFSR_11 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_47_DFFSR_100 INVX1_23/gnd DFFSR_186/S FILL
XFILL_1_OAI21X1_9 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_37_DFFSR_103 INVX1_8/gnd DFFSR_7/S FILL
XFILL_2_NAND2X1_244 INVX1_94/gnd DFFSR_52/S FILL
XFILL_27_DFFSR_106 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_0_DFFSR_179 INVX1_2/gnd DFFSR_1/S FILL
XFILL_47_DFFSR_61 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_3_INVX1_153 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_17_DFFSR_109 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_8_OAI21X1_28 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_28_0_0 INVX1_89/gnd DFFSR_36/S FILL
XFILL_7_OAI21X1_31 BUFX2_35/A DFFSR_97/S FILL
XFILL_3_DFFSR_58 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_31_DFFSR_11 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_6_NAND2X1_49 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_0_OAI21X1_226 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_6_DFFPOSX1_16 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_3_NAND2X1_178 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_5_NAND2X1_52 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_26_2_1 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_6_OAI21X1_34 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_20_DFFSR_51 INVX1_2/gnd DFFSR_51/S FILL
XFILL_8_1_0 BUFX2_43/A DFFSR_97/S FILL
XFILL_1_INVX1_370 BUFX2_36/A DFFSR_8/S FILL
XFILL_5_OAI21X1_37 INVX1_89/gnd DFFSR_2/S FILL
XFILL_4_NAND2X1_55 INVX1_89/gnd DFFSR_2/S FILL
XNAND2X1_49 INVX1_47/A DFFSR_11/S DFFSR_73/gnd NAND2X1_49/Y DFFSR_11/S NAND2X1
XFILL_24_4_2 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_4_OAI21X1_40 INVX1_8/gnd DFFSR_7/S FILL
XOAI21X1_34 DFFSR_1/S INVX1_39/Y NAND2X1_34/Y DFFSR_1/gnd DFFSR_34/D DFFSR_1/S OAI21X1
XFILL_3_DFFSR_106 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_3_NAND2X1_58 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_2_NAND2X1_61 BUFX2_37/A DFFSR_81/S FILL
XFILL_44_DFFSR_137 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_3_OAI21X1_43 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_46_DFFSR_7 INVX1_8/gnd DFFSR_7/S FILL
XFILL_1_OAI21X1_160 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_6_3_1 BUFX2_35/A DFFSR_14/S FILL
XFILL_2_OAI21X1_46 BUFX2_37/A DFFSR_81/S FILL
XFILL_34_DFFSR_140 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_4_NAND2X1_112 INVX1_4/gnd DFFSR_4/S FILL
XFILL_1_NAND2X1_64 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_11_AOI22X1_12 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_24_DFFSR_143 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_0_NAND2X1_67 INVX1_2/gnd DFFSR_1/S FILL
XFILL_1_OAI21X1_49 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_14_DFFSR_146 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_4_5_2 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_0_INVX1_190 BUFX2_43/A DFFSR_97/S FILL
XFILL_0_INVX1_52 BUFX2_37/A DFFSR_81/S FILL
XFILL_0_OAI21X1_52 INVX1_94/gnd DFFSR_25/S FILL
XFILL_17_DFFSR_98 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_39_DFFSR_18 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_28_DFFSR_58 DFFSR_3/gnd DFFSR_4/S FILL
XINVX1_300 INVX1_24/A BUFX2_16/gnd INVX1_300/Y DFFSR_11/S INVX1
XFILL_1_NAND2X1_274 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_4_INVX1_297 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_25_DFFPOSX1_24 BUFX2_43/A DFFSR_23/S FILL
XFILL_1_INVX1_9 BUFX2_36/A DFFSR_6/S FILL
XFILL_51_DFFSR_171 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_41_DFFSR_174 BUFX2_43/A DFFSR_97/S FILL
XFILL_0_DFFSR_143 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_2_NAND2X1_208 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_47_DFFSR_25 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_31_DFFSR_177 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_3_INVX1_117 INVX1_4/gnd DFFSR_51/S FILL
XFILL_36_DFFSR_65 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_1_NAND3X1_106 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_6_NAND2X1_13 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_0_OAI21X1_190 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_3_DFFSR_22 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_5_NAND2X1_16 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_20_DFFSR_15 INVX1_8/gnd DFFSR_7/S FILL
XFILL_21_DFFSR_180 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_11_DFFSR_183 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_3_NAND2X1_142 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_9_OAI21X1_245 DFFSR_5/gnd DFFSR_2/S FILL
XNAND2X1_13 DFFSR_11/S DFFSR_5/Q DFFSR_73/gnd NAND2X1_13/Y DFFSR_11/S NAND2X1
XFILL_1_INVX1_334 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_8_OAI21X1_7 INVX1_8/gnd DFFSR_5/S FILL
XFILL_11_OAI22X1_60 INVX1_8/gnd DFFSR_5/S FILL
XFILL_4_NAND2X1_19 DFFSR_1/gnd DFFSR_1/S FILL
XDFFPOSX1_16 INVX1_402/A CLKBUF1_14/Y AOI21X1_42/Y BUFX2_6/gnd DFFSR_91/S DFFPOSX1
XFILL_3_NAND2X1_22 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_2_NOR2X1_3 INVX1_94/gnd DFFSR_25/S FILL
XFILL_10_OAI22X1_63 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_12_DFFSR_5 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_44_DFFSR_101 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_2_NAND2X1_25 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_1_OAI21X1_124 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_7_DFFSR_177 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_44_DFFSR_72 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_34_DFFSR_104 INVX1_4/gnd DFFSR_4/S FILL
XFILL_24_DFFSR_107 BUFX2_36/A DFFSR_8/S FILL
XFILL_1_NAND2X1_28 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_2_OAI21X1_10 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_0_NAND2X1_31 BUFX2_43/A DFFSR_97/S FILL
XFILL_0_INVX1_16 BUFX2_43/A DFFSR_23/S FILL
XFILL_0_DFFSR_69 BUFX2_43/A DFFSR_23/S FILL
XFILL_17_DFFSR_62 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_8_NAND3X1_84 INVX1_94/gnd DFFSR_25/S FILL
XFILL_28_DFFSR_22 BUFX2_8/gnd DFFSR_10/S FILL
XINVX1_264 NOR2X1_1/A DFFSR_71/gnd INVX1_264/Y DFFSR_10/S INVX1
XFILL_0_INVX1_154 INVX1_8/gnd DFFSR_7/S FILL
XFILL_9_OAI22X1_66 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_1_OAI21X1_13 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_7_NAND3X1_87 INVX1_94/gnd DFFSR_52/S FILL
XFILL_1_NAND2X1_238 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_0_OAI21X1_16 INVX1_89/gnd DFFSR_36/S FILL
XFILL_14_DFFSR_110 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_6_NAND3X1_90 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_4_INVX1_261 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_5_NAND3X1_93 BUFX2_5/gnd DFFSR_23/S FILL
XNAND3X1_90 INVX1_258/A NAND3X1_90/B NAND3X1_90/C BUFX2_5/gnd NAND3X1_97/C DFFSR_23/S
+ NAND3X1
XFILL_4_NAND3X1_96 BUFX2_43/A DFFSR_97/S FILL
XFILL_33_DFFSR_1 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_3_NAND3X1_99 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_51_DFFSR_135 BUFX2_43/A DFFSR_97/S FILL
XFILL_2_NAND2X1_172 BUFX2_36/A DFFSR_6/S FILL
XFILL_0_DFFSR_107 BUFX2_36/A DFFSR_8/S FILL
XFILL_5_DFFPOSX1_10 INVX1_8/gnd DFFSR_5/S FILL
XFILL_25_DFFSR_69 BUFX2_43/A DFFSR_23/S FILL
XFILL_8_DFFSR_76 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_36_DFFSR_29 INVX1_4/gnd DFFSR_4/S FILL
XFILL_41_DFFSR_138 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_31_DFFSR_141 INVX1_94/gnd DFFSR_25/S FILL
XFILL_21_DFFSR_144 INVX1_8/gnd DFFSR_5/S FILL
XFILL_7_CLKBUF1_9 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_14_DFFPOSX1_29 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_11_DFFSR_147 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_0_OAI21X1_154 BUFX2_37/A DFFSR_8/S FILL
XFILL_9_OAI21X1_209 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_3_NAND2X1_106 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_6_NOR2X1_23 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_1_INVX1_298 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_0_NAND2X1_268 BUFX2_37/A DFFSR_8/S FILL
XFILL_33_DFFSR_76 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_44_DFFSR_36 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_10_OAI22X1_27 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_9_NAND3X1_45 BUFX2_35/A DFFSR_97/S FILL
XFILL_48_DFFSR_172 BUFX2_37/A DFFSR_8/S FILL
XFILL_24_DFFPOSX1_18 BUFX2_37/A DFFSR_8/S FILL
XFILL_7_DFFSR_141 INVX1_94/gnd DFFSR_25/S FILL
XFILL_38_DFFSR_175 INVX1_23/gnd DFFSR_91/S FILL
XFILL_8_NAND3X1_48 BUFX2_43/A DFFSR_23/S FILL
XFILL_9_OAI22X1_30 INVX1_94/gnd DFFSR_25/S FILL
XFILL_0_INVX1_118 BUFX2_37/A DFFSR_8/S FILL
XFILL_7_NAND3X1_51 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_0_DFFSR_33 INVX1_94/gnd DFFSR_52/S FILL
XFILL_25_5_0 DFFSR_71/gnd DFFSR_45/S FILL
XINVX1_228 AOI21X1_3/Y DFFSR_5/gnd INVX1_228/Y DFFSR_2/S INVX1
XFILL_8_OAI22X1_33 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_17_DFFSR_26 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_1_NAND2X1_202 BUFX2_35/A DFFSR_97/S FILL
XFILL_6_NAND3X1_54 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_4_INVX1_225 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_7_OAI22X1_36 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_28_DFFSR_178 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_18_DFFSR_181 INVX1_23/gnd DFFSR_186/S FILL
XFILL_6_OAI22X1_39 BUFX2_37/A DFFSR_8/S FILL
XFILL_5_NAND3X1_57 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_0_NAND3X1_100 BUFX2_6/gnd DFFSR_14/S FILL
XNAND3X1_54 NAND3X1_56/A NAND3X1_52/Y NAND3X1_53/Y BUFX2_7/gnd NAND3X1_54/Y DFFSR_54/S
+ NAND3X1
XFILL_4_NAND3X1_60 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_5_OAI22X1_42 INVX1_8/gnd DFFSR_7/S FILL
XFILL_3_NAND3X1_63 BUFX2_43/A DFFSR_23/S FILL
XFILL_5_OAI21X1_8 BUFX2_36/A DFFSR_6/S FILL
XOAI22X1_39 INVX1_337/Y OAI22X1_39/B INVX1_336/Y OAI22X1_39/D BUFX2_37/A NOR2X1_29/B
+ DFFSR_8/S OAI22X1
XFILL_41_DFFSR_83 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_4_OAI22X1_45 INVX1_89/gnd DFFSR_2/S FILL
XDFFSR_181 INVX1_411/A INVX1_1/A DFFSR_183/R DFFSR_186/S DFFSR_181/D INVX1_23/gnd
+ DFFSR_186/S DFFSR
XFILL_2_NAND3X1_66 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_3_OAI22X1_48 BUFX2_37/A DFFSR_81/S FILL
XFILL_2_NAND2X1_136 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_41_DFFSR_102 INVX1_8/gnd DFFSR_7/S FILL
XFILL_8_OAI21X1_239 INVX1_4/gnd DFFSR_4/S FILL
XFILL_31_DFFSR_105 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_25_DFFSR_33 INVX1_94/gnd DFFSR_52/S FILL
XFILL_8_DFFSR_40 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_4_DFFSR_178 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_14_DFFSR_73 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_1_NAND3X1_69 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_2_OAI22X1_51 BUFX2_7/gnd DFFSR_81/S FILL
XNAND2X1_2 DFFSR_5/S INVX1_407/A INVX1_8/gnd OAI21X1_2/C DFFSR_5/S NAND2X1
XFILL_0_NAND3X1_72 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_1_OAI22X1_54 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_21_DFFSR_108 INVX1_89/gnd DFFSR_2/S FILL
XFILL_0_OAI21X1_118 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_9_OAI21X1_173 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_11_DFFSR_111 INVX1_8/gnd DFFSR_5/S FILL
XFILL_0_OAI22X1_57 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_0_DFFSR_4 INVX1_4/gnd DFFSR_4/S FILL
XFILL_49_DFFSR_90 INVX1_2/gnd DFFSR_1/S FILL
XFILL_1_INVX1_262 INVX1_2/gnd DFFSR_1/S FILL
XOAI22X1_1 INVX1_213/Y NOR2X1_7/A INVX1_214/Y INVX1_216/Y BUFX2_36/A OAI22X1_1/Y DFFSR_8/S
+ OAI22X1
XFILL_7_DFFSR_105 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_0_NAND2X1_232 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_33_DFFSR_40 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_5_DFFSR_87 DFFSR_3/gnd DFFSR_4/S FILL
XINVX1_74 DFFSR_65/Q DFFSR_3/gnd INVX1_74/Y DFFSR_4/S INVX1
XFILL_22_DFFSR_80 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_48_DFFSR_136 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_35_0_0 BUFX2_17/gnd DFFSR_57/S FILL
XINVX1_192 BUFX2_2/Y BUFX2_35/A INVX1_192/Y DFFSR_14/S INVX1
XFILL_8_NAND3X1_12 INVX1_94/gnd DFFSR_52/S FILL
XFILL_38_DFFSR_139 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_4_BUFX2_25 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_28_DFFSR_142 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_7_NAND3X1_15 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_33_2_1 INVX1_8/gnd DFFSR_7/S FILL
XFILL_1_NAND2X1_166 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_18_DFFSR_145 INVX1_23/gnd DFFSR_186/S FILL
XFILL_4_INVX1_189 BUFX2_35/A DFFSR_14/S FILL
XFILL_6_NAND3X1_18 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_24_DFFSR_8 BUFX2_36/A DFFSR_8/S FILL
XFILL_5_NAND3X1_21 BUFX2_7/gnd DFFSR_81/S FILL
XNAND3X1_18 INVX1_229/A NOR3X1_1/A INVX1_228/Y DFFSR_5/gnd INVX1_236/A DFFSR_5/S NAND3X1
XFILL_4_NAND3X1_24 BUFX2_37/A DFFSR_8/S FILL
XFILL_3_NOR2X1_24 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_41_DFFSR_47 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_2_INVX1_81 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_31_4_2 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_30_DFFSR_87 DFFSR_3/gnd DFFSR_4/S FILL
XDFFSR_145 DFFSR_145/Q CLKBUF1_12/Y DFFSR_145/R DFFSR_186/S DFFSR_145/D INVX1_23/gnd
+ DFFSR_186/S DFFSR
XFILL_13_DFFPOSX1_23 INVX1_23/gnd DFFSR_91/S FILL
XFILL_2_NAND2X1_100 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_8_OAI21X1_203 BUFX2_35/A DFFSR_14/S FILL
XFILL_3_NAND3X1_27 BUFX2_37/A DFFSR_81/S FILL
XFILL_2_NAND3X1_30 INVX1_94/gnd DFFSR_52/S FILL
XFILL_14_DFFSR_37 INVX1_89/gnd DFFSR_2/S FILL
XFILL_3_OAI22X1_12 INVX1_4/gnd DFFSR_51/S FILL
XFILL_2_INVX1_406 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_45_DFFSR_173 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_4_DFFSR_142 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_1_NAND3X1_33 INVX1_8/gnd DFFSR_7/S FILL
XFILL_2_OAI22X1_15 INVX1_4/gnd DFFSR_4/S FILL
XFILL_0_NAND3X1_36 BUFX2_35/A DFFSR_97/S FILL
XFILL_1_OAI22X1_18 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_35_DFFSR_176 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_23_DFFPOSX1_12 INVX1_8/gnd DFFSR_5/S FILL
XFILL_45_DFFSR_4 INVX1_4/gnd DFFSR_4/S FILL
XFILL_0_OAI22X1_21 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_1_INVX1_226 BUFX2_35/A DFFSR_14/S FILL
XFILL_49_DFFSR_54 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_25_DFFSR_179 INVX1_2/gnd DFFSR_1/S FILL
XFILL_38_DFFSR_94 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_15_DFFSR_182 INVX1_89/gnd DFFSR_36/S FILL
XDFFSR_91 DFFSR_91/Q INVX1_172/A DFFSR_89/R DFFSR_91/S DFFSR_91/D BUFX2_6/gnd DFFSR_91/S
+ DFFSR
XFILL_0_NAND2X1_196 BUFX2_7/gnd DFFSR_54/S FILL
XINVX1_38 DFFSR_33/Q INVX1_94/gnd INVX1_38/Y DFFSR_52/S INVX1
XFILL_22_DFFSR_44 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_5_DFFSR_51 INVX1_2/gnd DFFSR_51/S FILL
XFILL_48_DFFSR_100 INVX1_23/gnd DFFSR_186/S FILL
XFILL_11_DFFSR_84 BUFX2_43/A DFFSR_23/S FILL
XFILL_2_OAI21X1_9 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_38_DFFSR_103 INVX1_8/gnd DFFSR_7/S FILL
XFILL_0_INVX1_6 INVX1_8/gnd DFFSR_5/S FILL
XFILL_28_DFFSR_106 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_1_DFFSR_179 INVX1_2/gnd DFFSR_1/S FILL
XINVX1_156 INVX1_156/A DFFSR_73/gnd INVX1_156/Y DFFSR_57/S INVX1
XFILL_7_OAI21X1_233 BUFX2_36/A DFFSR_8/S FILL
XFILL_1_NAND2X1_130 INVX1_4/gnd DFFSR_4/S FILL
XFILL_18_DFFSR_109 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_2_INVX1_45 INVX1_8/gnd DFFSR_5/S FILL
XFILL_41_DFFSR_11 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_19_DFFSR_91 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_2_DFFSR_98 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_30_DFFSR_51 INVX1_2/gnd DFFSR_51/S FILL
XDFFSR_109 DFFSR_109/Q CLKBUF1_7/Y DFFSR_105/R DFFSR_14/S DFFSR_109/D BUFX2_6/gnd
+ DFFSR_14/S DFFSR
XFILL_2_INVX1_370 BUFX2_36/A DFFSR_8/S FILL
XFILL_8_OAI21X1_167 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_1_BUFX2_36 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_4_DFFSR_106 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_45_DFFSR_137 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_35_DFFSR_140 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_25_DFFSR_143 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_11_DFFSR_2 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_9_OAI21X1_101 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_15_DFFSR_146 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_1_INVX1_190 BUFX2_43/A DFFSR_97/S FILL
XFILL_27_DFFSR_98 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_49_DFFSR_18 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_38_DFFSR_58 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_40_4 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_0_NOR2X1_25 DFFSR_71/gnd DFFSR_45/S FILL
XDFFSR_55 DFFSR_55/Q DFFSR_28/CLK DFFSR_54/R DFFSR_36/S DFFSR_55/D INVX1_89/gnd DFFSR_36/S
+ DFFSR
XFILL_6_OAI21X1_263 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_0_NAND2X1_160 INVX1_8/gnd DFFSR_5/S FILL
XFILL_5_DFFSR_15 INVX1_8/gnd DFFSR_7/S FILL
XFILL_11_DFFSR_48 INVX1_4/gnd DFFSR_4/S FILL
XFILL_8_NAND3X1_113 BUFX2_8/gnd DFFSR_10/S FILL
XINVX1_120 INVX1_342/A DFFSR_1/gnd INVX1_120/Y DFFSR_1/S INVX1
XFILL_42_DFFSR_174 BUFX2_43/A DFFSR_97/S FILL
XFILL_12_DFFPOSX1_17 BUFX2_37/A DFFSR_8/S FILL
XFILL_1_DFFSR_143 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_7_OAI21X1_197 INVX1_8/gnd DFFSR_7/S FILL
XFILL_46_DFFSR_65 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_32_DFFSR_177 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_2_DFFSR_62 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_19_DFFSR_55 INVX1_89/gnd DFFSR_36/S FILL
XFILL_30_DFFSR_15 INVX1_8/gnd DFFSR_7/S FILL
XFILL_22_DFFSR_180 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_12_DFFSR_183 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_8_OAI21X1_131 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_2_INVX1_334 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_9_OAI21X1_7 INVX1_8/gnd DFFSR_5/S FILL
XFILL_32_5_0 INVX1_8/gnd DFFSR_5/S FILL
XFILL_45_DFFSR_101 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_8_DFFSR_177 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_35_DFFSR_104 INVX1_4/gnd DFFSR_4/S FILL
XFILL_2_DFFPOSX1_28 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_25_DFFSR_107 BUFX2_36/A DFFSR_8/S FILL
XFILL_27_DFFSR_62 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_38_DFFSR_22 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_1_INVX1_154 INVX1_8/gnd DFFSR_7/S FILL
XFILL_15_DFFSR_110 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_6_OAI21X1_227 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_0_NAND2X1_124 DFFSR_79/gnd DFFSR_36/S FILL
XDFFSR_19 INVX1_22/A DFFSR_15/CLK DFFSR_20/R DFFSR_9/S DFFSR_19/D DFFSR_1/gnd DFFSR_9/S
+ DFFSR
XFILL_11_DFFSR_12 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_1_DFFSR_107 BUFX2_36/A DFFSR_8/S FILL
XOAI21X1_263 NOR2X1_53/Y NOR2X1_52/A INVX1_434/Y DFFSR_5/gnd OAI21X1_263/Y DFFSR_5/S
+ OAI21X1
XFILL_7_OAI21X1_161 INVX1_23/gnd DFFSR_186/S FILL
XFILL_35_DFFSR_69 BUFX2_43/A DFFSR_23/S FILL
XFILL_46_DFFSR_29 INVX1_4/gnd DFFSR_4/S FILL
XFILL_42_DFFSR_138 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_32_DFFSR_141 INVX1_94/gnd DFFSR_25/S FILL
XFILL_22_DFFSR_144 INVX1_8/gnd DFFSR_5/S FILL
XFILL_8_CLKBUF1_9 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_2_DFFSR_26 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_12_DFFSR_147 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_19_DFFSR_19 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_42_0_0 INVX1_4/gnd DFFSR_4/S FILL
XFILL_2_INVX1_298 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_1_NOR2X1_7 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_19_CLKBUF1_12 BUFX2_43/A DFFSR_23/S FILL
XFILL_43_DFFSR_76 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_49_DFFSR_172 BUFX2_37/A DFFSR_8/S FILL
XFILL_8_DFFSR_141 INVX1_94/gnd DFFSR_25/S FILL
XFILL_18_CLKBUF1_15 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_5_OAI21X1_257 INVX1_2/gnd DFFSR_51/S FILL
XFILL_40_2_1 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_39_DFFSR_175 INVX1_23/gnd DFFSR_91/S FILL
XFILL_17_CLKBUF1_18 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_7_NAND3X1_107 BUFX2_43/A DFFSR_97/S FILL
XFILL_1_INVX1_118 BUFX2_37/A DFFSR_8/S FILL
XFILL_27_DFFSR_26 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_16_DFFSR_66 INVX1_2/gnd DFFSR_51/S FILL
XFILL_38_4_2 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_16_CLKBUF1_21 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_29_DFFSR_178 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_11_DFFPOSX1_11 INVX1_4/gnd DFFSR_4/S FILL
XFILL_15_CLKBUF1_24 INVX1_23/gnd DFFSR_186/S FILL
XFILL_19_DFFSR_181 INVX1_23/gnd DFFSR_186/S FILL
XFILL_6_OAI21X1_191 BUFX2_37/A DFFSR_8/S FILL
XFILL_3_XOR2X1_3 BUFX2_17/gnd DFFSR_7/S FILL
XOAI21X1_227 AOI21X1_25/C AOI21X1_22/Y AOI21X1_25/A BUFX2_5/gnd AOI21X1_26/A DFFSR_23/S
+ OAI21X1
XFILL_6_OAI21X1_8 BUFX2_36/A DFFSR_6/S FILL
XFILL_23_DFFSR_5 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_42_DFFSR_102 INVX1_8/gnd DFFSR_7/S FILL
XFILL_32_DFFSR_105 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_7_OAI21X1_125 BUFX2_35/A DFFSR_14/S FILL
XFILL_35_DFFSR_33 INVX1_94/gnd DFFSR_52/S FILL
XFILL_5_DFFSR_178 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_7_DFFSR_80 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_24_DFFSR_73 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_22_DFFSR_108 INVX1_89/gnd DFFSR_2/S FILL
XFILL_1_DFFPOSX1_22 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_12_DFFSR_111 INVX1_8/gnd DFFSR_5/S FILL
XFILL_6_BUFX2_18 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_2_INVX1_262 INVX1_2/gnd DFFSR_1/S FILL
XFILL_44_DFFSR_1 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_8_DFFSR_105 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_5_OAI21X1_221 BUFX2_35/A DFFSR_14/S FILL
XFILL_43_DFFSR_40 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_4_INVX1_74 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_32_DFFSR_80 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_49_DFFSR_136 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_22_1 INVX1_94/gnd DFFSR_25/S FILL
XFILL_16_DFFSR_30 INVX1_89/gnd DFFSR_36/S FILL
XFILL_39_DFFSR_139 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_29_DFFSR_142 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_19_DFFSR_145 INVX1_23/gnd DFFSR_186/S FILL
XFILL_20_DFFPOSX1_30 BUFX2_43/A DFFSR_97/S FILL
XFILL_6_OAI21X1_155 BUFX2_7/gnd DFFSR_81/S FILL
XNOR2X1_27 NOR2X1_27/A NOR2X1_27/B BUFX2_17/gnd NOR2X1_27/Y DFFSR_57/S NOR2X1
XFILL_4_NOR2X1_24 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_40_DFFSR_87 DFFSR_3/gnd DFFSR_4/S FILL
XOAI21X1_191 INVX1_224/A OAI21X1_201/C OAI21X1_190/Y BUFX2_37/A INVX1_233/A DFFSR_8/S
+ OAI21X1
XFILL_7_DFFSR_44 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_24_DFFSR_37 INVX1_89/gnd DFFSR_2/S FILL
XFILL_13_DFFSR_77 INVX1_89/gnd DFFSR_2/S FILL
XFILL_6_NAND2X1_269 INVX1_4/gnd DFFSR_4/S FILL
XFILL_3_INVX1_406 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_46_DFFSR_173 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_14_0_1 BUFX2_37/A DFFSR_8/S FILL
XFILL_5_DFFSR_142 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_4_OAI21X1_251 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_36_DFFSR_176 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_2_INVX1_226 BUFX2_35/A DFFSR_14/S FILL
XFILL_12_2_2 BUFX2_36/A DFFSR_6/S FILL
XFILL_26_DFFSR_179 INVX1_2/gnd DFFSR_1/S FILL
XFILL_48_DFFSR_94 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_6_NAND3X1_101 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_16_DFFSR_182 INVX1_89/gnd DFFSR_36/S FILL
XFILL_4_DFFSR_91 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_7_CLKBUF1_12 BUFX2_43/A DFFSR_23/S FILL
XFILL_49_DFFSR_100 INVX1_23/gnd DFFSR_186/S FILL
XFILL_21_DFFSR_84 BUFX2_43/A DFFSR_23/S FILL
XFILL_5_OAI21X1_185 BUFX2_36/A DFFSR_8/S FILL
XFILL_32_DFFSR_44 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_6_CLKBUF1_15 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_3_OAI21X1_9 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_5_CLKBUF1_18 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_39_DFFSR_103 INVX1_8/gnd DFFSR_7/S FILL
XFILL_5_5 BUFX2_6/gnd DFFSR_91/S FILL
XCLKBUF1_15 clk BUFX2_17/gnd CLKBUF1_15/Y DFFSR_7/S CLKBUF1
XFILL_4_CLKBUF1_21 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_2_DFFSR_179 INVX1_2/gnd DFFSR_1/S FILL
XFILL_3_BUFX2_29 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_3_CLKBUF1_24 INVX1_23/gnd DFFSR_186/S FILL
XFILL_29_DFFSR_106 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_19_DFFSR_109 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_6_OAI21X1_119 BUFX2_37/A DFFSR_8/S FILL
XFILL_0_DFFPOSX1_16 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_29_DFFSR_91 BUFX2_6/gnd DFFSR_91/S FILL
XOAI21X1_155 DFFSR_81/S INVX1_184/Y NAND2X1_155/Y BUFX2_7/gnd DFFSR_155/D DFFSR_81/S
+ OAI21X1
XFILL_40_DFFSR_51 INVX1_2/gnd DFFSR_51/S FILL
XFILL_1_INVX1_85 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_39_5_0 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_3_INVX1_370 BUFX2_36/A DFFSR_8/S FILL
XFILL_6_NAND2X1_233 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_13_DFFSR_41 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_5_DFFSR_106 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_5_NAND3X1_131 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_46_DFFSR_137 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_36_DFFSR_140 DFFSR_71/gnd DFFSR_10/S FILL
XNAND2X1_269 DFFSR_4/S INVX1_200/A INVX1_4/gnd NAND2X1_269/Y DFFSR_4/S NAND2X1
XFILL_4_OAI21X1_215 BUFX2_43/A DFFSR_97/S FILL
XFILL_35_DFFSR_8 BUFX2_36/A DFFSR_8/S FILL
XFILL_26_DFFSR_143 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_16_DFFSR_146 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_2_INVX1_190 BUFX2_43/A DFFSR_97/S FILL
XFILL_37_DFFSR_98 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_44_1 INVX1_4/gnd DFFSR_51/S FILL
XFILL_48_DFFSR_58 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_5_OAI21X1_149 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_19_DFFPOSX1_24 BUFX2_43/A DFFSR_23/S FILL
XFILL_1_NOR2X1_25 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_4_DFFSR_55 INVX1_89/gnd DFFSR_36/S FILL
XFILL_21_DFFSR_48 INVX1_4/gnd DFFSR_4/S FILL
XFILL_10_DFFSR_88 DFFSR_3/gnd DFFSR_4/S FILL
XNAND3X1_101 XOR2X1_6/Y AOI21X1_31/B AOI21X1_31/A DFFSR_89/gnd NAND3X1_101/Y DFFSR_186/S
+ NAND3X1
XFILL_0_INVX1_407 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_43_DFFSR_174 BUFX2_43/A DFFSR_97/S FILL
XFILL_2_DFFSR_143 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_5_NAND2X1_263 INVX1_2/gnd DFFSR_51/S FILL
XFILL_33_DFFSR_177 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_1_INVX1_49 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_18_DFFSR_95 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_29_DFFSR_55 INVX1_89/gnd DFFSR_36/S FILL
XFILL_40_DFFSR_15 INVX1_8/gnd DFFSR_7/S FILL
XFILL_23_DFFSR_180 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_13_DFFSR_183 DFFSR_89/gnd DFFSR_186/S FILL
XOAI21X1_119 BUFX2_20/Y INVX1_134/Y OAI21X1_119/C BUFX2_37/A DFFSR_119/D DFFSR_8/S
+ OAI21X1
XFILL_3_OAI21X1_245 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_47_2_1 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_3_INVX1_334 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_6_NAND2X1_197 INVX1_8/gnd DFFSR_5/S FILL
XFILL_0_BUFX2_40 BUFX2_35/A DFFSR_14/S FILL
XFILL_45_4_2 INVX1_2/gnd DFFSR_1/S FILL
XFILL_46_DFFSR_101 DFFSR_73/gnd DFFSR_57/S FILL
XNAND2X1_233 OAI22X1_4/Y NAND2X1_233/B BUFX2_7/gnd DFFPOSX1_9/D DFFSR_81/S NAND2X1
XFILL_9_DFFSR_177 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_36_DFFSR_104 INVX1_4/gnd DFFSR_4/S FILL
XFILL_4_OAI21X1_179 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_26_DFFSR_107 BUFX2_36/A DFFSR_8/S FILL
XFILL_37_DFFSR_62 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_48_DFFSR_22 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_2_INVX1_154 INVX1_8/gnd DFFSR_7/S FILL
XFILL_16_DFFSR_110 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_4_DFFSR_19 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_5_OAI21X1_113 INVX1_23/gnd DFFSR_91/S FILL
XFILL_21_DFFSR_12 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_10_DFFSR_52 INVX1_94/gnd DFFSR_52/S FILL
XFILL_0_INVX1_371 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_13_3_0 BUFX2_36/A DFFSR_8/S FILL
XFILL_2_DFFSR_107 BUFX2_36/A DFFSR_8/S FILL
XFILL_5_NAND2X1_227 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_45_DFFSR_69 BUFX2_43/A DFFSR_23/S FILL
XFILL_11_5_1 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_22_DFFSR_2 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_43_DFFSR_138 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_33_DFFSR_141 INVX1_94/gnd DFFSR_25/S FILL
XFILL_23_DFFSR_144 INVX1_8/gnd DFFSR_5/S FILL
XFILL_4_NAND3X1_125 INVX1_8/gnd DFFSR_5/S FILL
XFILL_9_CLKBUF1_9 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_13_DFFSR_147 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_6_BUFX2_3 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_29_DFFSR_19 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_1_DFFSR_66 INVX1_2/gnd DFFSR_51/S FILL
XFILL_18_DFFSR_59 INVX1_4/gnd DFFSR_51/S FILL
XFILL_1_INVX1_13 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_6_NAND2X1_161 INVX1_23/gnd DFFSR_186/S FILL
XFILL_3_OAI21X1_209 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_3_INVX1_298 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_50_DFFSR_172 BUFX2_37/A DFFSR_8/S FILL
XFILL_18_DFFPOSX1_18 BUFX2_37/A DFFSR_8/S FILL
XFILL_9_DFFSR_141 INVX1_94/gnd DFFSR_25/S FILL
XNAND2X1_197 AOI21X1_13/B NAND3X1_58/A INVX1_8/gnd NAND2X1_197/Y DFFSR_5/S NAND2X1
XFILL_4_OAI21X1_143 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_40_DFFSR_175 INVX1_23/gnd DFFSR_91/S FILL
XFILL_2_INVX1_118 BUFX2_37/A DFFSR_8/S FILL
XFILL_18_DFFPOSX1_3 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_37_DFFSR_26 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_26_DFFSR_66 INVX1_2/gnd DFFSR_51/S FILL
XFILL_9_DFFSR_73 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_30_DFFSR_178 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_17_DFFPOSX1_6 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_20_DFFSR_181 INVX1_23/gnd DFFSR_186/S FILL
XFILL_16_DFFPOSX1_9 BUFX2_37/A DFFSR_8/S FILL
XFILL_10_DFFSR_16 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_4_NAND2X1_257 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_10_DFFSR_184 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_7_OAI21X1_8 BUFX2_36/A DFFSR_6/S FILL
XFILL_0_INVX1_335 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_21_0_1 INVX1_94/gnd DFFSR_25/S FILL
XFILL_43_DFFSR_102 INVX1_8/gnd DFFSR_7/S FILL
XFILL_8_DFFPOSX1_29 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_2_OAI21X1_239 INVX1_4/gnd DFFSR_4/S FILL
XFILL_5_NAND2X1_191 BUFX2_37/A DFFSR_8/S FILL
XFILL_19_2_2 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_45_DFFSR_33 INVX1_94/gnd DFFSR_52/S FILL
XFILL_6_DFFSR_178 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_34_DFFSR_73 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_1_1_1 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_33_DFFSR_105 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_18_DFFSR_23 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_1_DFFSR_30 INVX1_89/gnd DFFSR_36/S FILL
XFILL_23_DFFSR_108 INVX1_89/gnd DFFSR_2/S FILL
XFILL_3_OAI21X1_173 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_10_OAI22X1_4 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_13_DFFSR_111 INVX1_8/gnd DFFSR_5/S FILL
XFILL_6_NAND2X1_125 BUFX2_35/A DFFSR_14/S FILL
XFILL_3_INVX1_262 INVX1_2/gnd DFFSR_1/S FILL
XFILL_9_DFFSR_105 DFFSR_89/gnd DFFSR_186/S FILL
XNAND2X1_161 BUFX2_2/Y INVX1_218/A INVX1_23/gnd NAND2X1_161/Y DFFSR_186/S NAND2X1
XFILL_42_DFFSR_80 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_4_OAI21X1_107 BUFX2_36/A DFFSR_6/S FILL
XFILL_50_DFFSR_136 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_26_DFFSR_30 INVX1_89/gnd DFFSR_36/S FILL
XFILL_9_DFFSR_37 INVX1_89/gnd DFFSR_2/S FILL
XFILL_15_DFFSR_70 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_40_DFFSR_139 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_30_DFFSR_142 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_46_5_0 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_20_DFFSR_145 INVX1_23/gnd DFFSR_186/S FILL
XFILL_10_DFFSR_148 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_4_NAND2X1_221 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_2_XOR2X1_7 INVX1_23/gnd DFFSR_91/S FILL
XFILL_5_NOR2X1_24 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_0_INVX1_299 INVX1_89/gnd DFFSR_36/S FILL
XFILL_3_NAND3X1_119 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_13_DFFSR_9 DFFSR_9/gnd DFFSR_9/S FILL
XINVX1_409 NAND2X1_4/B INVX1_2/gnd INVX1_409/Y DFFSR_51/S INVX1
XFILL_50_DFFSR_87 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_2_OAI21X1_203 BUFX2_35/A DFFSR_14/S FILL
XFILL_6_DFFSR_84 BUFX2_43/A DFFSR_23/S FILL
XFILL_5_NAND2X1_155 BUFX2_37/A DFFSR_81/S FILL
XFILL_34_DFFSR_37 INVX1_89/gnd DFFSR_2/S FILL
XFILL_47_DFFSR_173 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_6_DFFSR_142 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_23_DFFSR_77 INVX1_89/gnd DFFSR_2/S FILL
XFILL_8_OR2X2_1 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_5_BUFX2_22 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_17_DFFPOSX1_12 INVX1_8/gnd DFFSR_5/S FILL
XFILL_37_DFFSR_176 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_3_INVX1_226 BUFX2_35/A DFFSR_14/S FILL
XFILL_3_OAI21X1_137 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_9_OAI21X1_98 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_27_DFFSR_179 INVX1_2/gnd DFFSR_1/S FILL
XFILL_15_NOR3X1_1 INVX1_94/gnd DFFSR_52/S FILL
XFILL_17_DFFSR_182 INVX1_89/gnd DFFSR_36/S FILL
XFILL_34_DFFSR_5 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_50_DFFSR_100 INVX1_23/gnd DFFSR_186/S FILL
XNAND2X1_125 BUFX2_21/Y DFFSR_117/Q BUFX2_35/A OAI21X1_125/C DFFSR_14/S NAND2X1
XFILL_3_NAND2X1_251 BUFX2_35/A DFFSR_97/S FILL
XFILL_31_DFFSR_84 BUFX2_43/A DFFSR_23/S FILL
XFILL_3_INVX1_78 BUFX2_36/A DFFSR_8/S FILL
XFILL_42_DFFSR_44 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_8_AOI21X1_17 INVX1_8/gnd DFFSR_5/S FILL
XFILL_40_DFFSR_103 INVX1_8/gnd DFFSR_7/S FILL
XFILL_4_OAI21X1_9 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_9_2 BUFX2_43/A DFFSR_97/S FILL
XFILL_7_AOI21X1_20 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_6_DFFPOSX1_3 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_15_DFFSR_34 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_3_DFFSR_179 INVX1_2/gnd DFFSR_1/S FILL
XFILL_6_AOI21X1_23 BUFX2_5/gnd DFFSR_6/S FILL
XDFFPOSX1_3 INVX1_218/A CLKBUF1_15/Y DFFPOSX1_3/D DFFSR_71/gnd DFFSR_45/S DFFPOSX1
XFILL_30_DFFSR_106 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_5_DFFPOSX1_6 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_7_DFFPOSX1_23 INVX1_23/gnd DFFSR_91/S FILL
XFILL_20_DFFSR_109 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_5_AOI21X1_26 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_1_OAI21X1_233 BUFX2_36/A DFFSR_8/S FILL
XFILL_4_DFFPOSX1_9 BUFX2_37/A DFFSR_8/S FILL
XFILL_4_NAND2X1_185 BUFX2_19/gnd DFFSR_52/S FILL
XAOI21X1_23 AOI21X1_23/A NAND3X1_62/Y AOI21X1_23/C BUFX2_5/gnd AOI21X1_23/Y DFFSR_6/S
+ AOI21X1
XFILL_4_AOI21X1_29 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_10_DFFSR_112 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_39_DFFSR_91 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_3_AOI21X1_32 BUFX2_43/A DFFSR_23/S FILL
XFILL_50_DFFSR_51 INVX1_2/gnd DFFSR_51/S FILL
XINVX1_373 INVX1_88/A DFFSR_3/gnd INVX1_373/Y DFFSR_65/S INVX1
XFILL_0_INVX1_263 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_4_INVX1_370 BUFX2_36/A DFFSR_8/S FILL
XFILL_2_AOI21X1_35 INVX1_94/gnd DFFSR_25/S FILL
XFILL_2_OAI21X1_167 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_1_AOI21X1_38 BUFX2_36/A DFFSR_8/S FILL
XFILL_5_NAND2X1_119 BUFX2_37/A DFFSR_8/S FILL
XFILL_12_DFFSR_81 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_23_DFFSR_41 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_6_DFFSR_106 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_6_DFFSR_48 INVX1_4/gnd DFFSR_4/S FILL
XFILL_0_AOI21X1_41 BUFX2_35/A DFFSR_14/S FILL
XFILL_47_DFFSR_137 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_37_DFFSR_140 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_9_OAI21X1_62 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_27_DFFSR_143 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_2_NAND2X1_281 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_3_OAI21X1_101 BUFX2_17/gnd DFFSR_7/S FILL
XBUFX2_26 BUFX2_26/A DFFSR_9/gnd dout[0] DFFSR_9/S BUFX2
XFILL_17_DFFSR_146 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_3_INVX1_190 BUFX2_43/A DFFSR_97/S FILL
XFILL_20_3_0 INVX1_94/gnd DFFSR_52/S FILL
XFILL_26_DFFPOSX1_31 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_47_DFFSR_98 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_8_OAI21X1_65 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_7_OAI21X1_68 BUFX2_37/A DFFSR_81/S FILL
XFILL_8_AND2X2_7 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_18_5_1 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_2_NOR2X1_25 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_3_DFFSR_95 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_3_INVX1_42 INVX1_89/gnd DFFSR_36/S FILL
XFILL_0_OAI21X1_263 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_6_NAND2X1_86 INVX1_4/gnd DFFSR_51/S FILL
XFILL_31_DFFSR_48 INVX1_4/gnd DFFSR_4/S FILL
XFILL_20_DFFSR_88 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_0_4_0 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_3_NAND2X1_215 BUFX2_43/A DFFSR_23/S FILL
XFILL_5_NAND2X1_89 BUFX2_37/A DFFSR_8/S FILL
XFILL_6_OAI21X1_71 BUFX2_8/gnd DFFSR_10/S FILL
XNAND2X1_86 BUFX2_15/Y INVX1_88/A INVX1_4/gnd NAND2X1_86/Y DFFSR_51/S NAND2X1
XFILL_4_NAND2X1_92 BUFX2_5/gnd DFFSR_23/S FILL
XOAI21X1_71 BUFX2_19/Y INVX1_80/Y OAI21X1_71/C BUFX2_8/gnd DFFSR_71/D DFFSR_10/S OAI21X1
XFILL_1_INVX1_407 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_5_OAI21X1_74 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_2_BUFX2_33 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_3_DFFSR_143 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_2_NAND3X1_113 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_4_OAI21X1_77 INVX1_89/gnd DFFSR_36/S FILL
XFILL_3_NAND2X1_95 INVX1_89/gnd DFFSR_36/S FILL
XFILL_44_DFFSR_174 BUFX2_43/A DFFSR_97/S FILL
XFILL_1_DFFSR_8 BUFX2_36/A DFFSR_8/S FILL
XFILL_1_OAI21X1_197 INVX1_8/gnd DFFSR_7/S FILL
XFILL_2_NAND2X1_98 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_3_OAI21X1_80 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_4_NAND2X1_149 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_2_OAI21X1_83 INVX1_94/gnd DFFSR_52/S FILL
XFILL_34_DFFSR_177 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_0_INVX1_227 BUFX2_5/gnd DFFSR_6/S FILL
XINVX1_337 DFFSR_89/Q BUFX2_36/A INVX1_337/Y DFFSR_8/S INVX1
XFILL_28_DFFSR_95 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_39_DFFSR_55 INVX1_89/gnd DFFSR_36/S FILL
XFILL_0_INVX1_89 INVX1_89/gnd DFFSR_2/S FILL
XFILL_50_DFFSR_15 INVX1_8/gnd DFFSR_7/S FILL
XFILL_24_DFFSR_180 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_1_OAI21X1_86 INVX1_4/gnd DFFSR_51/S FILL
XFILL_14_DFFSR_183 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_0_OAI21X1_89 BUFX2_35/A DFFSR_14/S FILL
XFILL_6_DFFSR_12 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_4_INVX1_334 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_2_OAI21X1_131 DFFSR_9/gnd DFFSR_9/S FILL
XBUFX2_4 BUFX2_2/A BUFX2_8/gnd BUFX2_4/Y DFFSR_25/S BUFX2
XFILL_12_DFFSR_45 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_47_DFFSR_101 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_2_NAND2X1_245 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_0_DFFSR_180 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_37_DFFSR_104 INVX1_4/gnd DFFSR_4/S FILL
XFILL_27_DFFSR_107 BUFX2_36/A DFFSR_8/S FILL
XFILL_47_DFFSR_62 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_3_INVX1_154 INVX1_8/gnd DFFSR_7/S FILL
XFILL_28_0_1 INVX1_89/gnd DFFSR_36/S FILL
XFILL_8_OAI21X1_29 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_17_DFFSR_110 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_6_NAND2X1_50 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_0_NAND2X1_1 INVX1_2/gnd DFFSR_51/S FILL
XFILL_7_OAI21X1_32 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_31_DFFSR_12 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_0_OAI21X1_227 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_6_DFFPOSX1_17 BUFX2_37/A DFFSR_8/S FILL
XFILL_20_DFFSR_52 INVX1_94/gnd DFFSR_52/S FILL
XFILL_3_NAND2X1_179 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_5_NAND2X1_53 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_26_2_2 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_6_OAI21X1_35 INVX1_8/gnd DFFSR_5/S FILL
XFILL_3_DFFSR_59 INVX1_4/gnd DFFSR_51/S FILL
XFILL_1_INVX1_371 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_5_OAI21X1_38 DFFSR_5/gnd DFFSR_5/S FILL
XNAND2X1_50 DFFSR_5/S INVX1_48/A BUFX2_17/gnd NAND2X1_50/Y DFFSR_7/S NAND2X1
XFILL_4_NAND2X1_56 INVX1_4/gnd DFFSR_51/S FILL
XFILL_8_1_1 BUFX2_43/A DFFSR_97/S FILL
XFILL_3_DFFSR_107 BUFX2_36/A DFFSR_8/S FILL
XOAI21X1_35 DFFSR_5/S INVX1_40/Y OAI21X1_35/C INVX1_8/gnd DFFSR_35/D DFFSR_5/S OAI21X1
XFILL_4_OAI21X1_41 INVX1_8/gnd DFFSR_7/S FILL
XFILL_3_NAND2X1_59 INVX1_2/gnd DFFSR_1/S FILL
XFILL_46_DFFSR_8 BUFX2_36/A DFFSR_8/S FILL
XFILL_2_NAND2X1_62 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_3_OAI21X1_44 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_44_DFFSR_138 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_1_OAI21X1_161 INVX1_23/gnd DFFSR_186/S FILL
XFILL_4_NAND2X1_113 INVX1_23/gnd DFFSR_91/S FILL
XFILL_6_3_2 BUFX2_35/A DFFSR_14/S FILL
XFILL_34_DFFSR_141 INVX1_94/gnd DFFSR_25/S FILL
XFILL_2_OAI21X1_47 INVX1_89/gnd DFFSR_2/S FILL
XFILL_1_NAND2X1_65 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_0_NAND2X1_68 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_24_DFFSR_144 INVX1_8/gnd DFFSR_5/S FILL
XFILL_1_OAI21X1_50 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_14_DFFSR_147 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_17_DFFSR_99 BUFX2_35/A DFFSR_97/S FILL
XFILL_0_INVX1_191 BUFX2_5/gnd DFFSR_23/S FILL
XINVX1_301 INVX1_42/A INVX1_89/gnd INVX1_301/Y DFFSR_2/S INVX1
XFILL_0_INVX1_53 INVX1_89/gnd DFFSR_2/S FILL
XFILL_39_DFFSR_19 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_28_DFFSR_59 INVX1_4/gnd DFFSR_51/S FILL
XFILL_0_OAI21X1_53 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_1_NAND2X1_275 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_4_INVX1_298 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_25_DFFPOSX1_25 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_2_NAND2X1_209 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_0_DFFSR_144 INVX1_8/gnd DFFSR_5/S FILL
XFILL_41_DFFSR_175 INVX1_23/gnd DFFSR_91/S FILL
XFILL_3_INVX1_118 BUFX2_37/A DFFSR_8/S FILL
XFILL_47_DFFSR_26 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_36_DFFSR_66 INVX1_2/gnd DFFSR_51/S FILL
XFILL_1_NAND3X1_107 BUFX2_43/A DFFSR_97/S FILL
XFILL_31_DFFSR_178 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_21_DFFSR_181 INVX1_23/gnd DFFSR_186/S FILL
XFILL_6_NAND2X1_14 BUFX2_43/A DFFSR_23/S FILL
XFILL_3_DFFSR_23 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_0_OAI21X1_191 BUFX2_37/A DFFSR_8/S FILL
XFILL_20_DFFSR_16 DFFSR_71/gnd DFFSR_45/S FILL
XNAND2X1_14 DFFSR_97/S DFFSR_6/Q BUFX2_43/A OAI21X1_14/C DFFSR_23/S NAND2X1
XFILL_3_NAND2X1_143 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_5_NAND2X1_17 INVX1_8/gnd DFFSR_7/S FILL
XFILL_11_DFFSR_184 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_9_OAI21X1_246 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_4_NAND2X1_20 INVX1_23/gnd DFFSR_186/S FILL
XFILL_1_INVX1_335 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_11_OAI22X1_61 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_3_NAND2X1_23 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_8_OAI21X1_8 BUFX2_36/A DFFSR_6/S FILL
XDFFPOSX1_17 NAND2X1_168/A CLKBUF1_16/Y INVX1_403/Y BUFX2_37/A DFFSR_8/S DFFPOSX1
XFILL_2_NOR2X1_4 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_44_DFFSR_102 INVX1_8/gnd DFFSR_7/S FILL
XFILL_1_OAI21X1_125 BUFX2_35/A DFFSR_14/S FILL
XFILL_12_DFFSR_6 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_10_OAI22X1_64 INVX1_94/gnd DFFSR_25/S FILL
XFILL_7_DFFSR_178 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_2_NAND2X1_26 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_44_DFFSR_73 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_34_DFFSR_105 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_9_NAND3X1_82 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_1_NAND2X1_29 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_2_OAI21X1_11 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_1_OAI21X1_14 BUFX2_43/A DFFSR_23/S FILL
XFILL_28_DFFSR_23 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_17_DFFSR_63 INVX1_94/gnd DFFSR_52/S FILL
XFILL_0_INVX1_155 INVX1_94/gnd DFFSR_52/S FILL
XFILL_8_NAND3X1_85 BUFX2_8/gnd DFFSR_10/S FILL
XINVX1_265 NOR2X1_2/A DFFSR_71/gnd INVX1_265/Y DFFSR_10/S INVX1
XFILL_24_DFFSR_108 INVX1_89/gnd DFFSR_2/S FILL
XFILL_0_INVX1_17 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_0_DFFSR_70 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_9_OAI22X1_67 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_0_NAND2X1_32 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_11_OAI22X1_4 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_7_NAND3X1_88 INVX1_94/gnd DFFSR_52/S FILL
XFILL_0_OAI21X1_17 INVX1_8/gnd DFFSR_5/S FILL
XFILL_14_DFFSR_111 INVX1_8/gnd DFFSR_5/S FILL
XFILL_6_NAND3X1_91 BUFX2_43/A DFFSR_97/S FILL
XFILL_1_NAND2X1_239 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_4_INVX1_262 INVX1_2/gnd DFFSR_1/S FILL
XFILL_5_NAND3X1_94 BUFX2_35/A DFFSR_97/S FILL
XFILL_4_NAND3X1_97 BUFX2_35/A DFFSR_97/S FILL
XNAND3X1_91 NAND3X1_97/B NAND3X1_97/C INVX1_259/Y BUFX2_43/A NAND3X1_95/B DFFSR_97/S
+ NAND3X1
XFILL_33_DFFSR_2 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_2_NAND2X1_173 BUFX2_35/A DFFSR_14/S FILL
XFILL_0_DFFSR_108 INVX1_89/gnd DFFSR_2/S FILL
XFILL_5_DFFPOSX1_11 INVX1_4/gnd DFFSR_4/S FILL
XFILL_36_DFFSR_30 INVX1_89/gnd DFFSR_36/S FILL
XFILL_8_DFFSR_77 INVX1_89/gnd DFFSR_2/S FILL
XFILL_25_DFFSR_70 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_41_DFFSR_139 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_31_DFFSR_142 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_21_DFFSR_145 INVX1_23/gnd DFFSR_186/S FILL
XFILL_11_DFFSR_148 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_14_DFFPOSX1_30 BUFX2_43/A DFFSR_97/S FILL
XFILL_3_NAND2X1_107 BUFX2_36/A DFFSR_6/S FILL
XFILL_0_OAI21X1_155 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_9_OAI21X1_210 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_6_NOR2X1_24 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_1_INVX1_299 INVX1_89/gnd DFFSR_36/S FILL
XFILL_0_NOR3X1_1 INVX1_94/gnd DFFSR_52/S FILL
XFILL_0_AOI22X1_10 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_10_OAI22X1_28 INVX1_94/gnd DFFSR_25/S FILL
XFILL_44_DFFSR_37 INVX1_89/gnd DFFSR_2/S FILL
XFILL_0_NAND2X1_269 INVX1_4/gnd DFFSR_4/S FILL
XFILL_7_DFFSR_142 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_27_3_0 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_33_DFFSR_77 INVX1_89/gnd DFFSR_2/S FILL
XFILL_24_DFFPOSX1_19 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_48_DFFSR_173 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_8_NAND3X1_49 BUFX2_37/A DFFSR_8/S FILL
XFILL_9_OAI22X1_31 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_0_INVX1_119 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_7_NAND3X1_52 BUFX2_36/A DFFSR_8/S FILL
XFILL_25_5_1 DFFSR_71/gnd DFFSR_45/S FILL
XINVX1_229 INVX1_229/A DFFSR_5/gnd INVX1_229/Y DFFSR_2/S INVX1
XFILL_17_DFFSR_27 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_0_DFFSR_34 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_38_DFFSR_176 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_8_OAI22X1_34 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_4_INVX1_226 BUFX2_35/A DFFSR_14/S FILL
XFILL_1_NAND2X1_203 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_6_NAND3X1_55 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_7_OAI22X1_37 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_28_DFFSR_179 INVX1_2/gnd DFFSR_1/S FILL
XFILL_7_4_0 BUFX2_35/A DFFSR_97/S FILL
XFILL_6_OAI22X1_40 BUFX2_37/A DFFSR_8/S FILL
XFILL_5_NAND3X1_58 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_18_DFFSR_182 INVX1_89/gnd DFFSR_36/S FILL
XFILL_0_NAND3X1_101 DFFSR_89/gnd DFFSR_186/S FILL
XNAND3X1_55 NOR3X1_1/Y NAND3X1_51/Y NAND3X1_54/Y BUFX2_7/gnd NAND3X1_55/Y DFFSR_54/S
+ NAND3X1
XFILL_4_NAND3X1_61 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_51_DFFSR_100 INVX1_23/gnd DFFSR_186/S FILL
XFILL_41_DFFSR_84 BUFX2_43/A DFFSR_23/S FILL
XOAI22X1_40 INVX1_338/Y OAI22X1_40/B INVX1_339/Y OAI22X1_40/D BUFX2_37/A NOR2X1_29/A
+ DFFSR_8/S OAI22X1
XFILL_5_OAI22X1_43 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_3_NAND3X1_64 BUFX2_35/A DFFSR_14/S FILL
XFILL_2_NAND2X1_137 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_4_OAI22X1_46 BUFX2_19/gnd DFFSR_52/S FILL
XDFFSR_182 INVX1_412/A DFFSR_3/CLK DFFSR_183/R DFFSR_36/S DFFSR_182/D INVX1_89/gnd
+ DFFSR_36/S DFFSR
XFILL_8_OAI21X1_240 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_5_OAI21X1_9 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_2_NAND3X1_67 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_3_OAI22X1_49 INVX1_94/gnd DFFSR_25/S FILL
XFILL_41_DFFSR_103 INVX1_8/gnd DFFSR_7/S FILL
XFILL_8_DFFSR_41 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_25_DFFSR_34 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_14_DFFSR_74 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_4_DFFSR_179 INVX1_2/gnd DFFSR_1/S FILL
XFILL_1_NAND3X1_70 BUFX2_35/A DFFSR_14/S FILL
XFILL_2_OAI22X1_52 INVX1_94/gnd DFFSR_25/S FILL
XFILL_31_DFFSR_106 DFFSR_1/gnd DFFSR_1/S FILL
XNAND2X1_3 DFFSR_51/S NAND2X1_3/B INVX1_4/gnd NAND2X1_3/Y DFFSR_51/S NAND2X1
XFILL_21_DFFSR_109 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_0_NAND3X1_73 BUFX2_43/A DFFSR_23/S FILL
XFILL_0_OAI21X1_119 BUFX2_37/A DFFSR_8/S FILL
XFILL_1_OAI22X1_55 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_9_OAI21X1_174 BUFX2_43/A DFFSR_23/S FILL
XFILL_0_DFFSR_5 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_0_OAI22X1_58 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_11_DFFSR_112 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_49_DFFSR_91 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_1_INVX1_263 BUFX2_16/gnd DFFSR_65/S FILL
XOAI22X1_2 OAI22X1_2/A NOR2X1_8/A OAI22X1_2/C OAI22X1_2/D BUFX2_36/A OAI22X1_2/Y DFFSR_8/S
+ OAI22X1
XFILL_0_NAND2X1_233 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_22_DFFSR_81 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_33_DFFSR_41 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_7_DFFSR_106 DFFSR_1/gnd DFFSR_1/S FILL
XINVX1_75 INVX1_75/A INVX1_4/gnd INVX1_75/Y DFFSR_51/S INVX1
XFILL_5_DFFSR_88 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_48_DFFSR_137 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_35_0_1 BUFX2_17/gnd DFFSR_57/S FILL
XINVX1_193 BUFX2_7/Y BUFX2_36/A DFFSR_159/R DFFSR_6/S INVX1
XFILL_8_NAND3X1_13 INVX1_94/gnd DFFSR_25/S FILL
XFILL_38_DFFSR_140 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_7_NAND3X1_16 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_28_DFFSR_143 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_4_BUFX2_26 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_18_DFFSR_146 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_4_INVX1_190 BUFX2_43/A DFFSR_97/S FILL
XFILL_6_NAND3X1_19 INVX1_8/gnd DFFSR_5/S FILL
XFILL_33_2_2 INVX1_8/gnd DFFSR_7/S FILL
XFILL_1_NAND2X1_167 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_5_NAND3X1_22 BUFX2_37/A DFFSR_81/S FILL
XFILL_24_DFFSR_9 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_2_INVX1_82 BUFX2_35/A DFFSR_97/S FILL
XFILL_4_NAND3X1_25 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_3_NOR2X1_25 DFFSR_71/gnd DFFSR_45/S FILL
XNAND3X1_19 BUFX2_3/Y NOR3X1_1/A INVX1_228/Y INVX1_8/gnd NAND3X1_19/Y DFFSR_5/S NAND3X1
XFILL_41_DFFSR_48 INVX1_4/gnd DFFSR_4/S FILL
XFILL_30_DFFSR_88 DFFSR_3/gnd DFFSR_4/S FILL
XDFFSR_146 DFFSR_146/Q CLKBUF1_12/Y DFFSR_146/R DFFSR_92/S DFFSR_146/D DFFSR_89/gnd
+ DFFSR_92/S DFFSR
XFILL_13_DFFPOSX1_24 BUFX2_43/A DFFSR_23/S FILL
XFILL_3_NAND3X1_28 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_2_NAND2X1_101 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_4_OAI22X1_10 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_8_OAI21X1_204 BUFX2_36/A DFFSR_6/S FILL
XFILL_2_NAND3X1_31 INVX1_94/gnd DFFSR_52/S FILL
XFILL_2_INVX1_407 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_3_OAI22X1_13 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_4_DFFSR_143 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_14_DFFSR_38 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_1_NAND3X1_34 INVX1_2/gnd DFFSR_1/S FILL
XFILL_2_OAI22X1_16 INVX1_4/gnd DFFSR_4/S FILL
XFILL_0_NAND3X1_37 BUFX2_43/A DFFSR_97/S FILL
XFILL_45_DFFSR_174 BUFX2_43/A DFFSR_97/S FILL
XFILL_1_OAI22X1_19 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_23_DFFPOSX1_13 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_35_DFFSR_177 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_0_OAI22X1_22 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_1_INVX1_227 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_38_DFFSR_95 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_49_DFFSR_55 INVX1_89/gnd DFFSR_36/S FILL
XFILL_45_DFFSR_5 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_25_DFFSR_180 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_15_DFFSR_183 DFFSR_89/gnd DFFSR_186/S FILL
XDFFSR_92 DFFSR_92/Q INVX1_172/A DFFSR_89/R DFFSR_92/S DFFSR_92/D DFFSR_89/gnd DFFSR_92/S
+ DFFSR
XFILL_5_DFFSR_52 INVX1_94/gnd DFFSR_52/S FILL
XFILL_0_NAND2X1_197 INVX1_8/gnd DFFSR_5/S FILL
XINVX1_39 INVX1_39/A DFFSR_1/gnd INVX1_39/Y DFFSR_1/S INVX1
XFILL_11_DFFSR_85 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_22_DFFSR_45 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_48_DFFSR_101 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_0_INVX1_7 BUFX2_36/A DFFSR_8/S FILL
XFILL_1_DFFSR_180 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_38_DFFSR_104 INVX1_4/gnd DFFSR_4/S FILL
XINVX1_157 XOR2X1_11/B BUFX2_16/gnd INVX1_157/Y DFFSR_65/S INVX1
XFILL_7_OAI21X1_234 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_28_DFFSR_107 BUFX2_36/A DFFSR_8/S FILL
XFILL_1_NAND2X1_131 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_18_DFFSR_110 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_1_NAND2X1_1 INVX1_2/gnd DFFSR_51/S FILL
XFILL_19_DFFSR_92 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_41_DFFSR_12 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_2_DFFSR_99 BUFX2_35/A DFFSR_97/S FILL
XFILL_30_DFFSR_52 INVX1_94/gnd DFFSR_52/S FILL
XFILL_2_INVX1_46 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_2_INVX1_371 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_8_OAI21X1_168 BUFX2_36/A DFFSR_6/S FILL
XDFFSR_110 DFFSR_110/Q CLKBUF1_3/Y DFFSR_105/R DFFSR_57/S DFFSR_110/D DFFSR_73/gnd
+ DFFSR_57/S DFFSR
XFILL_4_DFFSR_107 BUFX2_36/A DFFSR_8/S FILL
XFILL_1_BUFX2_37 BUFX2_37/A DFFSR_81/S FILL
XFILL_45_DFFSR_138 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_35_DFFSR_141 INVX1_94/gnd DFFSR_25/S FILL
XFILL_25_DFFSR_144 INVX1_8/gnd DFFSR_5/S FILL
XFILL_9_OAI21X1_102 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_11_DFFSR_3 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_15_DFFSR_147 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_27_DFFSR_99 BUFX2_35/A DFFSR_97/S FILL
XFILL_1_INVX1_191 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_49_DFFSR_19 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_38_DFFSR_59 INVX1_4/gnd DFFSR_51/S FILL
XFILL_0_NAND2X1_161 INVX1_23/gnd DFFSR_186/S FILL
XFILL_5_DFFSR_16 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_6_OAI21X1_264 DFFSR_5/gnd DFFSR_5/S FILL
XDFFSR_56 DFFSR_56/Q DFFSR_24/CLK DFFSR_54/R DFFSR_1/S DFFSR_56/D INVX1_2/gnd DFFSR_51/S
+ DFFSR
XFILL_0_NOR2X1_26 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_11_DFFSR_49 DFFSR_73/gnd DFFSR_11/S FILL
XINVX1_121 INVX1_121/A BUFX2_36/A INVX1_121/Y DFFSR_6/S INVX1
XFILL_8_NAND3X1_114 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_12_DFFPOSX1_18 BUFX2_37/A DFFSR_8/S FILL
XFILL_1_DFFSR_144 INVX1_8/gnd DFFSR_5/S FILL
XFILL_42_DFFSR_175 INVX1_23/gnd DFFSR_91/S FILL
XFILL_7_OAI21X1_198 INVX1_8/gnd DFFSR_7/S FILL
XFILL_46_DFFSR_66 INVX1_2/gnd DFFSR_51/S FILL
XFILL_32_DFFSR_178 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_22_DFFSR_181 INVX1_23/gnd DFFSR_186/S FILL
XFILL_2_INVX1_10 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_2_DFFSR_63 INVX1_94/gnd DFFSR_52/S FILL
XFILL_30_DFFSR_16 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_19_DFFSR_56 INVX1_2/gnd DFFSR_51/S FILL
XFILL_34_3_0 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_12_DFFSR_184 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_8_OAI21X1_132 INVX1_4/gnd DFFSR_4/S FILL
XFILL_2_INVX1_335 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_9_OAI21X1_8 BUFX2_36/A DFFSR_6/S FILL
XFILL_32_5_1 INVX1_8/gnd DFFSR_5/S FILL
XFILL_45_DFFSR_102 INVX1_8/gnd DFFSR_7/S FILL
XFILL_8_DFFSR_178 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_2_DFFPOSX1_29 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_35_DFFSR_105 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_38_DFFSR_23 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_27_DFFSR_63 INVX1_94/gnd DFFSR_52/S FILL
XFILL_1_INVX1_155 INVX1_94/gnd DFFSR_52/S FILL
XFILL_25_DFFSR_108 INVX1_89/gnd DFFSR_2/S FILL
XFILL_15_DFFSR_111 INVX1_8/gnd DFFSR_5/S FILL
XDFFSR_20 DFFSR_20/Q DFFSR_20/CLK DFFSR_20/R DFFSR_92/S DFFSR_20/D DFFSR_89/gnd DFFSR_92/S
+ DFFSR
XFILL_0_NAND2X1_125 BUFX2_35/A DFFSR_14/S FILL
XFILL_6_OAI21X1_228 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_11_DFFSR_13 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_1_DFFSR_108 INVX1_89/gnd DFFSR_2/S FILL
XOAI21X1_264 INVX1_436/Y AOI21X1_46/Y NOR2X1_51/A DFFSR_5/gnd OAI21X1_264/Y DFFSR_5/S
+ OAI21X1
XFILL_7_OAI21X1_162 INVX1_23/gnd DFFSR_91/S FILL
XFILL_46_DFFSR_30 INVX1_89/gnd DFFSR_36/S FILL
XFILL_42_DFFSR_139 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_32_DFFSR_142 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_35_DFFSR_70 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_22_DFFSR_145 INVX1_23/gnd DFFSR_186/S FILL
XFILL_19_DFFSR_20 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_12_DFFSR_148 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_2_DFFSR_27 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_2_INVX1_299 INVX1_89/gnd DFFSR_36/S FILL
XFILL_1_NOR2X1_8 BUFX2_43/A DFFSR_23/S FILL
XFILL_20_CLKBUF1_10 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_42_0_1 INVX1_4/gnd DFFSR_4/S FILL
XFILL_8_DFFSR_142 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_43_DFFSR_77 INVX1_89/gnd DFFSR_2/S FILL
XFILL_5_OAI21X1_258 INVX1_2/gnd DFFSR_51/S FILL
XFILL_19_CLKBUF1_13 INVX1_4/gnd DFFSR_51/S FILL
XFILL_40_2_2 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_49_DFFSR_173 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_18_CLKBUF1_16 BUFX2_36/A DFFSR_6/S FILL
XFILL_1_INVX1_119 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_7_NAND3X1_108 BUFX2_37/A DFFSR_81/S FILL
XFILL_27_DFFSR_27 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_17_CLKBUF1_19 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_16_DFFSR_67 INVX1_2/gnd DFFSR_51/S FILL
XFILL_39_DFFSR_176 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_16_CLKBUF1_22 INVX1_94/gnd DFFSR_25/S FILL
XFILL_11_DFFPOSX1_12 INVX1_8/gnd DFFSR_5/S FILL
XFILL_29_DFFSR_179 INVX1_2/gnd DFFSR_1/S FILL
XFILL_15_CLKBUF1_25 INVX1_23/gnd DFFSR_186/S FILL
XFILL_6_OAI21X1_192 BUFX2_37/A DFFSR_81/S FILL
XFILL_19_DFFSR_182 INVX1_89/gnd DFFSR_36/S FILL
XFILL_3_XOR2X1_4 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_51_DFFSR_84 BUFX2_43/A DFFSR_23/S FILL
XFILL_23_DFFSR_6 BUFX2_5/gnd DFFSR_6/S FILL
XOAI21X1_228 AOI21X1_18/Y AOI21X1_17/Y INVX1_244/A DFFSR_71/gnd AOI21X1_35/A DFFSR_10/S
+ OAI21X1
XFILL_6_OAI21X1_9 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_7_DFFSR_81 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_42_DFFSR_103 INVX1_8/gnd DFFSR_7/S FILL
XFILL_7_OAI21X1_126 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_35_DFFSR_34 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_24_DFFSR_74 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_5_DFFSR_179 INVX1_2/gnd DFFSR_1/S FILL
XFILL_32_DFFSR_106 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_1_DFFPOSX1_23 INVX1_23/gnd DFFSR_91/S FILL
XFILL_22_DFFSR_109 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_6_BUFX2_19 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_12_DFFSR_112 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_2_INVX1_263 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_44_DFFSR_2 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_32_DFFSR_81 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_43_DFFSR_41 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_8_DFFSR_106 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_4_INVX1_75 INVX1_4/gnd DFFSR_51/S FILL
XFILL_5_OAI21X1_222 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_49_DFFSR_137 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_16_DFFSR_31 BUFX2_35/A DFFSR_97/S FILL
XFILL_39_DFFSR_140 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_22_2 INVX1_94/gnd DFFSR_25/S FILL
XFILL_29_DFFSR_143 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_19_DFFSR_146 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_6_OAI21X1_156 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_20_DFFPOSX1_31 BUFX2_17/gnd DFFSR_57/S FILL
XNOR2X1_28 NOR2X1_28/A NOR2X1_28/B INVX1_94/gnd NOR2X1_28/Y DFFSR_52/S NOR2X1
XFILL_4_NOR2X1_25 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_51_DFFSR_48 INVX1_4/gnd DFFSR_4/S FILL
XFILL_40_DFFSR_88 DFFSR_3/gnd DFFSR_4/S FILL
XOAI21X1_192 NAND3X1_8/A AOI22X1_2/Y NAND3X1_7/C BUFX2_37/A AOI21X1_5/C DFFSR_81/S
+ OAI21X1
XFILL_6_NAND2X1_270 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_7_DFFSR_45 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_3_INVX1_407 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_5_DFFSR_143 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_24_DFFSR_38 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_13_DFFSR_78 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_46_DFFSR_174 BUFX2_43/A DFFSR_97/S FILL
XFILL_14_0_2 BUFX2_37/A DFFSR_8/S FILL
XFILL_36_DFFSR_177 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_4_OAI21X1_252 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_2_INVX1_227 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_48_DFFSR_95 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_26_DFFSR_180 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_16_DFFSR_183 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_6_NAND3X1_102 INVX1_23/gnd DFFSR_186/S FILL
XFILL_8_CLKBUF1_10 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_7_CLKBUF1_13 INVX1_4/gnd DFFSR_51/S FILL
XFILL_4_DFFSR_92 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_6_CLKBUF1_16 BUFX2_36/A DFFSR_6/S FILL
XFILL_5_OAI21X1_186 BUFX2_36/A DFFSR_8/S FILL
XFILL_21_DFFSR_85 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_32_DFFSR_45 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_5_CLKBUF1_19 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_49_DFFSR_101 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_5_6 BUFX2_6/gnd DFFSR_91/S FILL
XCLKBUF1_16 clk BUFX2_36/A CLKBUF1_16/Y DFFSR_6/S CLKBUF1
XFILL_4_CLKBUF1_22 INVX1_94/gnd DFFSR_25/S FILL
XFILL_2_DFFSR_180 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_3_BUFX2_30 INVX1_4/gnd DFFSR_51/S FILL
XFILL_39_DFFSR_104 INVX1_4/gnd DFFSR_4/S FILL
XFILL_3_CLKBUF1_25 INVX1_23/gnd DFFSR_186/S FILL
XFILL_29_DFFSR_107 BUFX2_36/A DFFSR_8/S FILL
XFILL_41_3_0 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_6_OAI21X1_120 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_19_DFFSR_110 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_2_NAND2X1_1 INVX1_2/gnd DFFSR_51/S FILL
XFILL_29_DFFSR_92 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_51_DFFSR_12 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_0_DFFPOSX1_17 BUFX2_37/A DFFSR_8/S FILL
XFILL_1_INVX1_86 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_40_DFFSR_52 INVX1_94/gnd DFFSR_52/S FILL
XFILL_39_5_1 BUFX2_16/gnd DFFSR_65/S FILL
XOAI21X1_156 DFFSR_91/S INVX1_186/Y OAI21X1_156/C BUFX2_6/gnd DFFSR_156/D DFFSR_14/S
+ OAI21X1
XFILL_3_INVX1_371 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_6_NAND2X1_234 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_5_DFFSR_107 BUFX2_36/A DFFSR_8/S FILL
XFILL_13_DFFSR_42 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_5_NAND3X1_132 INVX1_8/gnd DFFSR_7/S FILL
XFILL_46_DFFSR_138 DFFSR_73/gnd DFFSR_11/S FILL
XNAND2X1_270 DFFSR_52/S INVX1_201/A BUFX2_19/gnd OAI21X1_259/C DFFSR_52/S NAND2X1
XFILL_36_DFFSR_141 INVX1_94/gnd DFFSR_25/S FILL
XFILL_4_OAI21X1_216 BUFX2_35/A DFFSR_14/S FILL
XFILL_26_DFFSR_144 INVX1_8/gnd DFFSR_5/S FILL
XFILL_35_DFFSR_9 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_16_DFFSR_147 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_37_DFFSR_99 BUFX2_35/A DFFSR_97/S FILL
XFILL_2_INVX1_191 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_48_DFFSR_59 INVX1_4/gnd DFFSR_51/S FILL
XFILL_44_2 INVX1_4/gnd DFFSR_51/S FILL
XFILL_10_DFFSR_89 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_19_DFFPOSX1_25 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_4_DFFSR_56 INVX1_2/gnd DFFSR_51/S FILL
XFILL_21_DFFSR_49 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_5_OAI21X1_150 INVX1_94/gnd DFFSR_52/S FILL
XFILL_1_NOR2X1_26 DFFSR_73/gnd DFFSR_11/S FILL
XNAND3X1_102 INVX1_254/Y AOI21X1_30/B AOI21X1_30/A INVX1_23/gnd NAND3X1_102/Y DFFSR_186/S
+ NAND3X1
XFILL_0_INVX1_408 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_2_DFFSR_144 INVX1_8/gnd DFFSR_5/S FILL
XFILL_5_NAND2X1_264 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_43_DFFSR_175 INVX1_23/gnd DFFSR_91/S FILL
XFILL_33_DFFSR_178 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_23_DFFSR_181 INVX1_23/gnd DFFSR_186/S FILL
XFILL_1_INVX1_50 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_40_DFFSR_16 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_18_DFFSR_96 INVX1_2/gnd DFFSR_1/S FILL
XFILL_29_DFFSR_56 INVX1_2/gnd DFFSR_51/S FILL
XFILL_13_DFFSR_184 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_47_2_2 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_3_OAI21X1_246 DFFSR_9/gnd DFFSR_9/S FILL
XOAI21X1_120 BUFX2_16/Y INVX1_135/Y OAI21X1_120/C BUFX2_16/gnd DFFSR_120/D DFFSR_65/S
+ OAI21X1
XFILL_3_INVX1_335 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_6_NAND2X1_198 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_0_BUFX2_41 BUFX2_37/A DFFSR_81/S FILL
XFILL_46_DFFSR_102 INVX1_8/gnd DFFSR_7/S FILL
XFILL_9_DFFSR_178 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_36_DFFSR_105 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_4_OAI21X1_180 DFFSR_71/gnd DFFSR_10/S FILL
XNAND2X1_234 NOR2X1_13/Y NOR2X1_12/Y BUFX2_16/gnd NAND2X1_65/A DFFSR_65/S NAND2X1
XFILL_48_DFFSR_23 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_37_DFFSR_63 INVX1_94/gnd DFFSR_52/S FILL
XFILL_2_INVX1_155 INVX1_94/gnd DFFSR_52/S FILL
XFILL_26_DFFSR_108 INVX1_89/gnd DFFSR_2/S FILL
XFILL_15_1_0 BUFX2_37/A DFFSR_81/S FILL
XFILL_16_DFFSR_111 INVX1_8/gnd DFFSR_5/S FILL
XFILL_4_DFFSR_20 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_10_DFFSR_53 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_5_OAI21X1_114 INVX1_89/gnd DFFSR_36/S FILL
XFILL_21_DFFSR_13 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_13_3_1 BUFX2_36/A DFFSR_8/S FILL
XFILL_0_INVX1_372 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_3_NOR2X1_1 BUFX2_36/A DFFSR_6/S FILL
XFILL_2_DFFSR_108 INVX1_89/gnd DFFSR_2/S FILL
XFILL_11_5_2 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_43_DFFSR_139 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_22_DFFSR_3 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_5_NAND2X1_228 INVX1_23/gnd DFFSR_91/S FILL
XFILL_33_DFFSR_142 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_45_DFFSR_70 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_23_DFFSR_145 INVX1_23/gnd DFFSR_186/S FILL
XFILL_4_NAND3X1_126 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_29_DFFSR_20 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_13_DFFSR_148 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_1_INVX1_14 BUFX2_35/A DFFSR_14/S FILL
XFILL_18_DFFSR_60 BUFX2_37/A DFFSR_8/S FILL
XFILL_1_DFFSR_67 INVX1_2/gnd DFFSR_51/S FILL
XFILL_6_BUFX2_4 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_6_NAND2X1_162 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_3_OAI21X1_210 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_3_INVX1_299 INVX1_89/gnd DFFSR_36/S FILL
XFILL_9_DFFSR_142 BUFX2_19/gnd DFFSR_54/S FILL
XNAND2X1_198 INVX1_235/Y NAND2X1_197/Y BUFX2_17/gnd AOI21X1_17/B DFFSR_57/S NAND2X1
XFILL_18_DFFPOSX1_19 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_50_DFFSR_173 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_19_DFFPOSX1_1 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_4_OAI21X1_144 INVX1_8/gnd DFFSR_7/S FILL
XFILL_2_INVX1_119 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_18_DFFPOSX1_4 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_37_DFFSR_27 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_9_DFFSR_74 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_26_DFFSR_67 INVX1_2/gnd DFFSR_51/S FILL
XFILL_40_DFFSR_176 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_17_DFFPOSX1_7 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_30_DFFSR_179 INVX1_2/gnd DFFSR_1/S FILL
XFILL_20_DFFSR_182 INVX1_89/gnd DFFSR_36/S FILL
XFILL_10_DFFSR_17 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_4_NAND2X1_258 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_10_DFFSR_185 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_0_INVX1_336 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_21_0_2 INVX1_94/gnd DFFSR_25/S FILL
XFILL_7_OAI21X1_9 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_8_DFFPOSX1_30 BUFX2_43/A DFFSR_97/S FILL
XFILL_5_NAND2X1_192 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_2_OAI21X1_240 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_43_DFFSR_103 INVX1_8/gnd DFFSR_7/S FILL
XFILL_45_DFFSR_34 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_34_DFFSR_74 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_6_DFFSR_179 INVX1_2/gnd DFFSR_1/S FILL
XFILL_1_1_2 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_33_DFFSR_106 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_23_DFFSR_109 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_1_DFFSR_31 BUFX2_35/A DFFSR_97/S FILL
XFILL_18_DFFSR_24 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_3_OAI21X1_174 BUFX2_43/A DFFSR_23/S FILL
XFILL_13_DFFSR_112 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_10_OAI22X1_5 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_6_NAND2X1_126 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_3_INVX1_263 BUFX2_16/gnd DFFSR_65/S FILL
XXOR2X1_1 XOR2X1_1/A NOR2X1_4/A DFFSR_79/gnd XOR2X1_1/Y DFFSR_45/S XOR2X1
XFILL_42_DFFSR_81 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_9_DFFSR_106 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_50_DFFSR_137 BUFX2_7/gnd DFFSR_54/S FILL
XNAND2X1_162 BUFX2_4/Y AOI21X1_1/C BUFX2_8/gnd OAI21X1_162/C DFFSR_25/S NAND2X1
XFILL_4_OAI21X1_108 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_48_3_0 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_26_DFFSR_31 BUFX2_35/A DFFSR_97/S FILL
XFILL_40_DFFSR_140 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_9_DFFSR_38 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_30_DFFSR_143 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_15_DFFSR_71 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_46_5_1 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_20_DFFSR_146 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_4_NAND2X1_222 INVX1_23/gnd DFFSR_186/S FILL
XFILL_10_DFFSR_149 INVX1_23/gnd DFFSR_91/S FILL
XFILL_2_XOR2X1_8 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_50_DFFSR_88 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_0_INVX1_300 BUFX2_16/gnd DFFSR_11/S FILL
XINVX1_410 NAND2X1_5/B DFFSR_73/gnd INVX1_410/Y DFFSR_11/S INVX1
XFILL_5_NOR2X1_25 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_3_NAND3X1_120 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_5_NAND2X1_156 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_2_OAI21X1_204 BUFX2_36/A DFFSR_6/S FILL
XFILL_6_DFFSR_143 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_6_DFFSR_85 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_34_DFFSR_38 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_23_DFFSR_78 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_47_DFFSR_174 BUFX2_43/A DFFSR_97/S FILL
XFILL_8_OR2X2_2 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_5_BUFX2_23 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_37_DFFSR_177 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_17_DFFPOSX1_13 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_9_OAI21X1_99 BUFX2_43/A DFFSR_97/S FILL
XFILL_3_INVX1_227 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_27_DFFSR_180 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_3_OAI21X1_138 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_17_DFFSR_183 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_34_DFFSR_6 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_15_NOR3X1_2 INVX1_89/gnd DFFSR_2/S FILL
XFILL_3_NAND2X1_252 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_31_DFFSR_85 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_42_DFFSR_45 DFFSR_79/gnd DFFSR_45/S FILL
XNAND2X1_126 BUFX2_16/Y INVX1_374/A BUFX2_17/gnd OAI21X1_126/C DFFSR_7/S NAND2X1
XFILL_3_INVX1_79 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_7_DFFPOSX1_1 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_8_AOI21X1_18 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_50_DFFSR_101 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_9_3 BUFX2_43/A DFFSR_97/S FILL
XFILL_7_AOI21X1_21 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_15_DFFSR_35 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_3_DFFSR_180 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_6_DFFPOSX1_4 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_40_DFFSR_104 INVX1_4/gnd DFFSR_4/S FILL
XFILL_6_AOI21X1_24 BUFX2_43/A DFFSR_97/S FILL
XFILL_30_DFFSR_107 BUFX2_36/A DFFSR_8/S FILL
XFILL_5_DFFPOSX1_7 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_1_OAI21X1_234 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_7_DFFPOSX1_24 BUFX2_43/A DFFSR_23/S FILL
XFILL_5_AOI21X1_27 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_4_NAND2X1_186 BUFX2_37/A DFFSR_81/S FILL
XDFFPOSX1_4 AOI21X1_1/C CLKBUF1_10/Y DFFPOSX1_4/D BUFX2_17/gnd DFFSR_7/S DFFPOSX1
XFILL_20_DFFSR_110 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_10_DFFSR_113 INVX1_23/gnd DFFSR_186/S FILL
XFILL_4_AOI21X1_30 INVX1_23/gnd DFFSR_91/S FILL
XAOI21X1_24 INVX1_241/Y NAND3X1_37/B NOR2X1_8/Y BUFX2_43/A NAND3X1_69/C DFFSR_97/S
+ AOI21X1
XFILL_3_NAND2X1_1 INVX1_2/gnd DFFSR_51/S FILL
XFILL_39_DFFSR_92 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_3_AOI21X1_33 BUFX2_35/A DFFSR_14/S FILL
XFILL_50_DFFSR_52 INVX1_94/gnd DFFSR_52/S FILL
XFILL_0_INVX1_264 DFFSR_71/gnd DFFSR_10/S FILL
XINVX1_374 INVX1_374/A BUFX2_17/gnd INVX1_374/Y DFFSR_7/S INVX1
XFILL_2_AOI21X1_36 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_0_AND2X2_1 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_2_OAI21X1_168 BUFX2_36/A DFFSR_6/S FILL
XFILL_6_DFFSR_107 BUFX2_36/A DFFSR_8/S FILL
XFILL_1_AOI21X1_39 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_12_DFFSR_82 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_23_DFFSR_42 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_5_NAND2X1_120 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_6_DFFSR_49 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_0_AOI21X1_42 INVX1_23/gnd DFFSR_91/S FILL
XFILL_47_DFFSR_138 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_37_DFFSR_141 INVX1_94/gnd DFFSR_25/S FILL
XFILL_22_1_0 BUFX2_8/gnd DFFSR_25/S FILL
XBUFX2_27 BUFX2_27/A DFFSR_89/gnd dout[1] DFFSR_186/S BUFX2
XFILL_2_NAND2X1_282 INVX1_89/gnd DFFSR_2/S FILL
XFILL_27_DFFSR_144 INVX1_8/gnd DFFSR_5/S FILL
XFILL_3_OAI21X1_102 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_17_DFFSR_147 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_47_DFFSR_99 BUFX2_35/A DFFSR_97/S FILL
XFILL_3_INVX1_191 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_20_3_1 INVX1_94/gnd DFFSR_52/S FILL
XFILL_9_OAI21X1_63 INVX1_94/gnd DFFSR_25/S FILL
XFILL_2_2_0 INVX1_23/gnd DFFSR_186/S FILL
XFILL_8_OAI21X1_66 INVX1_4/gnd DFFSR_51/S FILL
XFILL_20_DFFSR_89 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_8_AND2X2_8 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_7_OAI21X1_69 BUFX2_37/A DFFSR_8/S FILL
XFILL_18_5_2 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_6_NAND2X1_87 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_3_INVX1_43 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_0_OAI21X1_264 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_3_DFFSR_96 INVX1_2/gnd DFFSR_1/S FILL
XFILL_31_DFFSR_49 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_3_NAND2X1_216 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_6_OAI21X1_72 DFFSR_5/gnd DFFSR_2/S FILL
XNAND2X1_87 BUFX2_22/Y DFFSR_79/Q DFFSR_5/gnd NAND2X1_87/Y DFFSR_2/S NAND2X1
XFILL_5_NAND2X1_90 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_2_NOR2X1_26 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_0_4_1 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_1_INVX1_408 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_5_OAI21X1_75 INVX1_4/gnd DFFSR_4/S FILL
XFILL_4_NAND2X1_93 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_2_BUFX2_34 BUFX2_37/A DFFSR_81/S FILL
XFILL_2_NAND3X1_114 DFFSR_71/gnd DFFSR_10/S FILL
XOAI21X1_72 BUFX2_17/Y INVX1_81/Y OAI21X1_72/C DFFSR_5/gnd DFFSR_72/D DFFSR_2/S OAI21X1
XFILL_3_DFFSR_144 INVX1_8/gnd DFFSR_5/S FILL
XFILL_4_OAI21X1_78 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_3_NAND2X1_96 INVX1_4/gnd DFFSR_51/S FILL
XFILL_44_DFFSR_175 INVX1_23/gnd DFFSR_91/S FILL
XFILL_2_NAND2X1_99 BUFX2_43/A DFFSR_97/S FILL
XFILL_3_OAI21X1_81 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_1_OAI21X1_198 INVX1_8/gnd DFFSR_7/S FILL
XFILL_1_DFFSR_9 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_2_OAI21X1_84 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_4_NAND2X1_150 BUFX2_37/A DFFSR_81/S FILL
XFILL_34_DFFSR_178 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_24_DFFSR_181 INVX1_23/gnd DFFSR_186/S FILL
XINVX1_338 DFFSR_121/Q BUFX2_36/A INVX1_338/Y DFFSR_8/S INVX1
XFILL_50_DFFSR_16 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_0_INVX1_228 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_28_DFFSR_96 INVX1_2/gnd DFFSR_1/S FILL
XFILL_39_DFFSR_56 INVX1_2/gnd DFFSR_51/S FILL
XFILL_1_OAI21X1_87 INVX1_4/gnd DFFSR_4/S FILL
XFILL_0_INVX1_90 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_0_OAI21X1_90 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_14_DFFSR_184 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_2_OAI21X1_132 INVX1_4/gnd DFFSR_4/S FILL
XBUFX2_5 rst BUFX2_5/gnd BUFX2_5/Y DFFSR_23/S BUFX2
XFILL_12_DFFSR_46 BUFX2_36/A DFFSR_6/S FILL
XFILL_5_BUFX2_1 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_6_DFFSR_13 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_47_DFFSR_102 INVX1_8/gnd DFFSR_7/S FILL
XFILL_37_DFFSR_105 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_0_DFFSR_181 INVX1_23/gnd DFFSR_186/S FILL
XFILL_47_DFFSR_63 INVX1_94/gnd DFFSR_52/S FILL
XFILL_3_INVX1_155 INVX1_94/gnd DFFSR_52/S FILL
XFILL_2_NAND2X1_246 INVX1_94/gnd DFFSR_25/S FILL
XFILL_27_DFFSR_108 INVX1_89/gnd DFFSR_2/S FILL
XFILL_8_OAI21X1_30 INVX1_89/gnd DFFSR_36/S FILL
XFILL_28_0_2 INVX1_89/gnd DFFSR_36/S FILL
XFILL_17_DFFSR_111 INVX1_8/gnd DFFSR_5/S FILL
XFILL_7_OAI21X1_33 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_0_NAND2X1_2 INVX1_8/gnd DFFSR_5/S FILL
XFILL_6_NAND2X1_51 INVX1_2/gnd DFFSR_51/S FILL
XFILL_6_DFFPOSX1_18 BUFX2_37/A DFFSR_8/S FILL
XFILL_3_DFFSR_60 BUFX2_37/A DFFSR_8/S FILL
XFILL_5_NAND2X1_54 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_3_NAND2X1_180 INVX1_94/gnd DFFSR_52/S FILL
XFILL_0_OAI21X1_228 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_20_DFFSR_53 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_6_OAI21X1_36 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_31_DFFSR_13 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_5_OAI21X1_39 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_4_NAND2X1_57 BUFX2_17/gnd DFFSR_57/S FILL
XNAND2X1_51 DFFSR_1/S DFFSR_43/Q INVX1_2/gnd OAI21X1_51/C DFFSR_51/S NAND2X1
XFILL_1_INVX1_372 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_8_1_2 BUFX2_43/A DFFSR_97/S FILL
XFILL_3_NAND2X1_60 BUFX2_7/gnd DFFSR_54/S FILL
XOAI21X1_36 DFFSR_45/S INVX1_41/Y NAND2X1_36/Y DFFSR_79/gnd DFFSR_36/D DFFSR_45/S
+ OAI21X1
XFILL_3_DFFSR_108 INVX1_89/gnd DFFSR_2/S FILL
XFILL_4_OAI21X1_42 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_0_OAI22X1_1 BUFX2_36/A DFFSR_8/S FILL
XFILL_2_NAND2X1_63 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_44_DFFSR_139 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_1_OAI21X1_162 INVX1_23/gnd DFFSR_91/S FILL
XFILL_34_DFFSR_142 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_3_OAI21X1_45 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_4_NAND2X1_114 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_46_DFFSR_9 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_24_DFFSR_145 INVX1_23/gnd DFFSR_186/S FILL
XFILL_11_AOI22X1_14 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_1_NAND2X1_66 INVX1_4/gnd DFFSR_51/S FILL
XFILL_2_OAI21X1_48 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_39_DFFSR_20 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_14_DFFSR_148 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_0_INVX1_192 BUFX2_35/A DFFSR_14/S FILL
XFILL_28_DFFSR_60 BUFX2_37/A DFFSR_8/S FILL
XFILL_0_NAND2X1_69 BUFX2_19/gnd DFFSR_54/S FILL
XINVX1_302 INVX1_33/A INVX1_8/gnd INVX1_302/Y DFFSR_7/S INVX1
XFILL_1_OAI21X1_51 INVX1_2/gnd DFFSR_51/S FILL
XFILL_0_INVX1_54 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_0_OAI21X1_54 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_1_NAND2X1_276 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_4_INVX1_299 INVX1_89/gnd DFFSR_36/S FILL
XFILL_25_DFFPOSX1_26 BUFX2_37/A DFFSR_81/S FILL
XFILL_12_DFFSR_10 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_0_DFFSR_145 INVX1_23/gnd DFFSR_186/S FILL
XFILL_2_NAND2X1_210 BUFX2_35/A DFFSR_97/S FILL
XFILL_3_INVX1_119 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_47_DFFSR_27 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_36_DFFSR_67 INVX1_2/gnd DFFSR_51/S FILL
XFILL_41_DFFSR_176 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_1_NAND3X1_108 BUFX2_37/A DFFSR_81/S FILL
XFILL_31_DFFSR_179 INVX1_2/gnd DFFSR_1/S FILL
XFILL_0_OAI21X1_192 BUFX2_37/A DFFSR_81/S FILL
XFILL_21_DFFSR_182 INVX1_89/gnd DFFSR_36/S FILL
XFILL_20_DFFSR_17 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_6_NAND2X1_15 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_3_DFFSR_24 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_11_DFFSR_185 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_3_NAND2X1_144 INVX1_8/gnd DFFSR_7/S FILL
XNAND2X1_15 DFFSR_15/S INVX1_8/A BUFX2_17/gnd NAND2X1_15/Y DFFSR_7/S NAND2X1
XFILL_9_OAI21X1_247 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_5_NAND2X1_18 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_1_INVX1_336 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_4_NAND2X1_21 INVX1_4/gnd DFFSR_4/S FILL
XDFFPOSX1_18 NAND2X1_169/B CLKBUF1_16/Y XOR2X1_9/Y BUFX2_37/A DFFSR_8/S DFFPOSX1
XFILL_11_OAI22X1_62 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_2_NOR2X1_5 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_3_NAND2X1_24 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_8_OAI21X1_9 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_12_DFFSR_7 INVX1_8/gnd DFFSR_7/S FILL
XFILL_44_DFFSR_103 INVX1_8/gnd DFFSR_7/S FILL
XFILL_1_OAI21X1_126 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_2_NAND2X1_27 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_44_DFFSR_74 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_7_DFFSR_179 INVX1_2/gnd DFFSR_1/S FILL
XFILL_10_OAI22X1_65 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_2_OAI21X1_12 BUFX2_35/A DFFSR_14/S FILL
XFILL_1_NAND2X1_30 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_34_DFFSR_106 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_24_DFFSR_109 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_8_NAND3X1_86 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_0_NAND2X1_33 BUFX2_19/gnd DFFSR_52/S FILL
XINVX1_266 NOR2X1_1/B BUFX2_8/gnd INVX1_266/Y DFFSR_10/S INVX1
XFILL_0_DFFSR_71 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_0_INVX1_18 INVX1_89/gnd DFFSR_2/S FILL
XFILL_9_OAI22X1_68 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_1_OAI21X1_15 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_28_DFFSR_24 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_0_INVX1_156 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_7_NAND3X1_89 BUFX2_43/A DFFSR_23/S FILL
XFILL_0_OAI21X1_18 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_14_DFFSR_112 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_11_OAI22X1_5 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_17_DFFSR_64 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_6_NAND3X1_92 BUFX2_43/A DFFSR_23/S FILL
XFILL_1_NAND2X1_240 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_5_NAND3X1_95 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_4_NAND3X1_98 BUFX2_35/A DFFSR_14/S FILL
XNAND3X1_92 NAND3X1_92/A INVX1_258/A NAND3X1_92/C BUFX2_43/A NAND3X1_94/B DFFSR_23/S
+ NAND3X1
XFILL_4_XOR2X1_1 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_33_DFFSR_3 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_0_DFFSR_109 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_13_1 BUFX2_36/A DFFSR_6/S FILL
XFILL_5_DFFPOSX1_12 INVX1_8/gnd DFFSR_5/S FILL
XFILL_2_NAND2X1_174 BUFX2_43/A DFFSR_97/S FILL
XFILL_41_DFFSR_140 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_8_DFFSR_78 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_36_DFFSR_31 BUFX2_35/A DFFSR_97/S FILL
XFILL_31_DFFSR_143 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_25_DFFSR_71 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_21_DFFSR_146 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_11_DFFSR_149 INVX1_23/gnd DFFSR_91/S FILL
XFILL_0_OAI21X1_156 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_3_NAND2X1_108 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_14_DFFPOSX1_31 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_1_INVX1_300 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_6_NOR2X1_25 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_0_NOR3X1_2 INVX1_89/gnd DFFSR_2/S FILL
XFILL_29_1_0 INVX1_89/gnd DFFSR_2/S FILL
XFILL_0_AOI22X1_11 INVX1_23/gnd DFFSR_91/S FILL
XFILL_0_NAND2X1_270 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_10_OAI22X1_29 INVX1_8/gnd DFFSR_5/S FILL
XFILL_24_DFFPOSX1_20 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_7_DFFSR_143 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_27_3_1 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_44_DFFSR_38 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_33_DFFSR_78 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_48_DFFSR_174 BUFX2_43/A DFFSR_97/S FILL
XFILL_8_NAND3X1_50 BUFX2_37/A DFFSR_81/S FILL
XFILL_9_OAI22X1_32 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_9_2_0 BUFX2_43/A DFFSR_23/S FILL
XFILL_7_NAND3X1_53 BUFX2_37/A DFFSR_81/S FILL
XFILL_17_DFFSR_28 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_25_5_2 DFFSR_71/gnd DFFSR_45/S FILL
XINVX1_230 NOR3X1_1/A DFFSR_79/gnd INVX1_230/Y DFFSR_45/S INVX1
XFILL_0_DFFSR_35 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_38_DFFSR_177 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_8_OAI22X1_35 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_0_INVX1_120 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_4_INVX1_227 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_1_NAND2X1_204 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_6_NAND3X1_56 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_28_DFFSR_180 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_18_DFFSR_183 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_7_4_1 BUFX2_35/A DFFSR_97/S FILL
XFILL_7_OAI22X1_38 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_0_NAND3X1_102 INVX1_23/gnd DFFSR_186/S FILL
XNAND3X1_56 NAND3X1_56/A NAND3X1_49/Y NAND3X1_50/Y BUFX2_7/gnd NAND3X1_56/Y DFFSR_81/S
+ NAND3X1
XFILL_5_NAND3X1_59 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_6_OAI22X1_41 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_4_NAND3X1_62 BUFX2_43/A DFFSR_23/S FILL
XFILL_41_DFFSR_85 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_5_OAI22X1_44 BUFX2_16/gnd DFFSR_11/S FILL
XOAI22X1_41 INVX1_341/Y OAI22X1_49/D INVX1_340/Y OAI22X1_52/D DFFSR_73/gnd NOR2X1_30/B
+ DFFSR_57/S OAI22X1
XDFFSR_183 INVX1_413/A DFFSR_20/CLK DFFSR_183/R DFFSR_186/S DFFSR_183/D DFFSR_89/gnd
+ DFFSR_186/S DFFSR
XFILL_3_NAND3X1_65 BUFX2_35/A DFFSR_14/S FILL
XFILL_8_OAI21X1_241 BUFX2_35/A DFFSR_97/S FILL
XFILL_4_OAI22X1_47 BUFX2_37/A DFFSR_8/S FILL
XFILL_2_NAND2X1_138 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_2_NAND3X1_68 BUFX2_35/A DFFSR_14/S FILL
XFILL_3_OAI22X1_50 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_25_DFFSR_35 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_4_DFFSR_180 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_14_DFFSR_75 INVX1_4/gnd DFFSR_51/S FILL
XFILL_41_DFFSR_104 INVX1_4/gnd DFFSR_4/S FILL
XFILL_8_DFFSR_42 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_1_NAND3X1_71 BUFX2_35/A DFFSR_14/S FILL
XFILL_31_DFFSR_107 BUFX2_36/A DFFSR_8/S FILL
XFILL_2_OAI22X1_53 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_0_NAND3X1_74 BUFX2_35/A DFFSR_14/S FILL
XFILL_1_OAI22X1_56 BUFX2_37/A DFFSR_8/S FILL
XNAND2X1_4 DFFSR_1/S NAND2X1_4/B INVX1_2/gnd OAI21X1_4/C DFFSR_51/S NAND2X1
XFILL_0_OAI21X1_120 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_21_DFFSR_110 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_11_DFFSR_113 INVX1_23/gnd DFFSR_186/S FILL
XFILL_9_OAI21X1_175 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_0_OAI22X1_59 INVX1_8/gnd DFFSR_7/S FILL
XFILL_4_NAND2X1_1 INVX1_2/gnd DFFSR_51/S FILL
XFILL_49_DFFSR_92 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_0_DFFSR_6 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_1_INVX1_264 DFFSR_71/gnd DFFSR_10/S FILL
XOAI22X1_3 NAND3X1_2/A OAI22X1_3/B OAI22X1_3/C OAI22X1_3/D DFFSR_79/gnd OAI22X1_3/Y
+ DFFSR_45/S OAI22X1
XFILL_5_DFFSR_89 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_7_DFFSR_107 BUFX2_36/A DFFSR_8/S FILL
XFILL_22_DFFSR_82 DFFSR_1/gnd DFFSR_9/S FILL
XINVX1_76 DFFSR_67/Q INVX1_2/gnd INVX1_76/Y DFFSR_1/S INVX1
XFILL_33_DFFSR_42 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_0_NAND2X1_234 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_9_NAND3X1_11 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_35_0_2 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_48_DFFSR_138 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_8_NAND3X1_14 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_38_DFFSR_141 INVX1_94/gnd DFFSR_25/S FILL
XINVX1_194 DFFSR_160/Q DFFSR_73/gnd INVX1_194/Y DFFSR_57/S INVX1
XFILL_4_BUFX2_27 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_7_NAND3X1_17 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_28_DFFSR_144 INVX1_8/gnd DFFSR_5/S FILL
XFILL_35_1 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_18_DFFSR_147 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_4_INVX1_191 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_1_NAND2X1_168 BUFX2_36/A DFFSR_6/S FILL
XFILL_6_NAND3X1_20 BUFX2_37/A DFFSR_8/S FILL
XFILL_5_NAND3X1_23 BUFX2_37/A DFFSR_81/S FILL
XFILL_30_DFFSR_89 DFFSR_89/gnd DFFSR_92/S FILL
XNAND3X1_20 AOI22X1_5/D AOI22X1_5/C NAND3X1_24/C BUFX2_37/A AOI21X1_5/A DFFSR_8/S
+ NAND3X1
XFILL_4_NAND3X1_26 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_9_NAND3X1_121 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_2_INVX1_83 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_41_DFFSR_49 DFFSR_73/gnd DFFSR_11/S FILL
XDFFSR_147 INVX1_168/A CLKBUF1_12/Y DFFSR_147/R DFFSR_186/S DFFSR_147/D DFFSR_89/gnd
+ DFFSR_186/S DFFSR
XFILL_3_NAND3X1_29 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_13_DFFPOSX1_25 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_2_NAND2X1_102 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_4_OAI22X1_11 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_3_NOR2X1_26 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_8_OAI21X1_205 BUFX2_36/A DFFSR_8/S FILL
XFILL_2_NAND3X1_32 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_2_INVX1_408 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_3_OAI22X1_14 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_1_NAND3X1_35 BUFX2_35/A DFFSR_97/S FILL
XFILL_2_OAI22X1_17 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_14_DFFSR_39 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_4_DFFSR_144 INVX1_8/gnd DFFSR_5/S FILL
XFILL_45_DFFSR_175 INVX1_23/gnd DFFSR_91/S FILL
XFILL_0_NAND3X1_38 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_1_OAI22X1_20 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_23_DFFPOSX1_14 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_0_OAI22X1_23 INVX1_89/gnd DFFSR_2/S FILL
XFILL_35_DFFSR_178 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_25_DFFSR_181 INVX1_23/gnd DFFSR_186/S FILL
XFILL_45_DFFSR_6 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_1_INVX1_228 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_49_DFFSR_56 INVX1_2/gnd DFFSR_51/S FILL
XFILL_38_DFFSR_96 INVX1_2/gnd DFFSR_1/S FILL
XFILL_15_DFFSR_184 DFFSR_1/gnd DFFSR_9/S FILL
XINVX1_40 DFFSR_35/Q INVX1_8/gnd INVX1_40/Y DFFSR_5/S INVX1
XFILL_0_NAND2X1_198 BUFX2_17/gnd DFFSR_57/S FILL
XDFFSR_93 DFFSR_93/Q CLKBUF1_5/Y DFFSR_89/R DFFSR_51/S DFFSR_93/D INVX1_2/gnd DFFSR_51/S
+ DFFSR
XFILL_22_DFFSR_46 BUFX2_36/A DFFSR_6/S FILL
XFILL_5_DFFSR_53 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_11_DFFSR_86 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_48_DFFSR_102 INVX1_8/gnd DFFSR_7/S FILL
XFILL_38_DFFSR_105 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_1_DFFSR_181 INVX1_23/gnd DFFSR_186/S FILL
XINVX1_158 DFFSR_140/Q DFFSR_79/gnd INVX1_158/Y DFFSR_36/S INVX1
XFILL_0_INVX1_8 INVX1_8/gnd DFFSR_5/S FILL
XFILL_7_OAI21X1_235 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_4_INVX1_155 INVX1_94/gnd DFFSR_52/S FILL
XFILL_28_DFFSR_108 INVX1_89/gnd DFFSR_2/S FILL
XFILL_1_NAND2X1_132 INVX1_8/gnd DFFSR_5/S FILL
XFILL_18_DFFSR_111 INVX1_8/gnd DFFSR_5/S FILL
XFILL_1_NAND2X1_2 INVX1_8/gnd DFFSR_5/S FILL
XFILL_30_DFFSR_53 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_2_INVX1_47 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_19_DFFSR_93 INVX1_2/gnd DFFSR_51/S FILL
XFILL_41_DFFSR_13 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_8_OAI21X1_169 BUFX2_36/A DFFSR_8/S FILL
XDFFSR_111 INVX1_387/A CLKBUF1_4/Y DFFSR_105/R DFFSR_5/S DFFSR_111/D INVX1_8/gnd DFFSR_5/S
+ DFFSR
XFILL_4_DFFSR_108 INVX1_89/gnd DFFSR_2/S FILL
XFILL_2_INVX1_372 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_1_OAI22X1_1 BUFX2_36/A DFFSR_8/S FILL
XFILL_1_BUFX2_38 BUFX2_37/A DFFSR_81/S FILL
XFILL_45_DFFSR_139 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_35_DFFSR_142 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_25_DFFSR_145 INVX1_23/gnd DFFSR_186/S FILL
XFILL_9_OAI21X1_103 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_11_DFFSR_4 INVX1_4/gnd DFFSR_4/S FILL
XFILL_49_DFFSR_20 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_15_DFFSR_148 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_1_INVX1_192 BUFX2_35/A DFFSR_14/S FILL
XFILL_38_DFFSR_60 BUFX2_37/A DFFSR_8/S FILL
XFILL_6_OAI21X1_265 BUFX2_43/A DFFSR_97/S FILL
XFILL_0_NAND2X1_162 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_22_DFFSR_10 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_5_DFFSR_17 DFFSR_5/gnd DFFSR_5/S FILL
XDFFSR_57 DFFSR_57/Q DFFSR_2/CLK DFFSR_61/R DFFSR_57/S DFFSR_57/D DFFSR_73/gnd DFFSR_57/S
+ DFFSR
XFILL_11_DFFSR_50 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_0_NOR2X1_27 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_8_NAND3X1_115 BUFX2_8/gnd DFFSR_10/S FILL
XINVX1_122 INVX1_122/A DFFSR_71/gnd INVX1_122/Y DFFSR_10/S INVX1
XFILL_1_DFFSR_145 INVX1_23/gnd DFFSR_186/S FILL
XFILL_12_DFFPOSX1_19 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_4_INVX1_119 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_7_OAI21X1_199 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_46_DFFSR_67 INVX1_2/gnd DFFSR_51/S FILL
XFILL_42_DFFSR_176 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_32_DFFSR_179 INVX1_2/gnd DFFSR_1/S FILL
XFILL_36_1_0 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_22_DFFSR_182 INVX1_89/gnd DFFSR_36/S FILL
XFILL_30_DFFSR_17 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_19_DFFSR_57 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_2_INVX1_11 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_2_DFFSR_64 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_12_DFFSR_185 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_34_3_1 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_2_INVX1_336 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_8_OAI21X1_133 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_9_OAI21X1_9 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_2_DFFPOSX1_30 BUFX2_43/A DFFSR_97/S FILL
XFILL_32_5_2 INVX1_8/gnd DFFSR_5/S FILL
XFILL_45_DFFSR_103 INVX1_8/gnd DFFSR_7/S FILL
XFILL_8_DFFSR_179 INVX1_2/gnd DFFSR_1/S FILL
XFILL_35_DFFSR_106 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_25_DFFSR_109 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_38_DFFSR_24 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_1_INVX1_156 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_15_DFFSR_112 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_27_DFFSR_64 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_0_NAND2X1_126 BUFX2_17/gnd DFFSR_7/S FILL
XDFFSR_21 INVX1_24/A DFFSR_1/CLK DFFSR_20/R DFFSR_1/S DFFSR_21/D INVX1_2/gnd DFFSR_1/S
+ DFFSR
XFILL_11_DFFSR_14 BUFX2_35/A DFFSR_14/S FILL
XFILL_6_OAI21X1_229 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_1_DFFSR_109 BUFX2_6/gnd DFFSR_14/S FILL
XOAI21X1_265 NOR2X1_1/B NOR2X1_1/A INVX1_437/Y BUFX2_43/A AOI21X1_47/C DFFSR_97/S
+ OAI21X1
XFILL_42_DFFSR_140 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_7_OAI21X1_163 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_46_DFFSR_31 BUFX2_35/A DFFSR_97/S FILL
XFILL_32_DFFSR_143 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_35_DFFSR_71 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_22_DFFSR_146 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_12_DFFSR_149 INVX1_23/gnd DFFSR_91/S FILL
XFILL_2_DFFSR_28 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_19_DFFSR_21 INVX1_2/gnd DFFSR_1/S FILL
XFILL_2_INVX1_300 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_1_NOR2X1_9 BUFX2_43/A DFFSR_97/S FILL
XFILL_42_0_2 INVX1_4/gnd DFFSR_4/S FILL
XFILL_20_CLKBUF1_11 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_5_OAI21X1_259 INVX1_23/gnd DFFSR_186/S FILL
XFILL_19_CLKBUF1_14 BUFX2_43/A DFFSR_23/S FILL
XFILL_8_DFFSR_143 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_43_DFFSR_78 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_49_DFFSR_174 BUFX2_43/A DFFSR_97/S FILL
XFILL_18_CLKBUF1_17 INVX1_94/gnd DFFSR_25/S FILL
XFILL_16_DFFSR_68 BUFX2_35/A DFFSR_14/S FILL
XFILL_7_NAND3X1_109 BUFX2_36/A DFFSR_8/S FILL
XFILL_27_DFFSR_28 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_39_DFFSR_177 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_1_INVX1_120 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_17_CLKBUF1_20 INVX1_4/gnd DFFSR_51/S FILL
XFILL_11_DFFPOSX1_13 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_16_CLKBUF1_23 INVX1_89/gnd DFFSR_2/S FILL
XFILL_29_DFFSR_180 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_19_DFFSR_183 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_6_OAI21X1_193 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_3_XOR2X1_5 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_23_DFFSR_7 INVX1_8/gnd DFFSR_7/S FILL
XOAI21X1_229 AOI21X1_29/Y OAI21X1_229/B NAND3X1_2/A DFFSR_71/gnd OAI22X1_3/D DFFSR_45/S
+ OAI21X1
XFILL_7_OAI21X1_127 BUFX2_43/A DFFSR_23/S FILL
XFILL_35_DFFSR_35 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_5_DFFSR_180 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_7_DFFSR_82 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_24_DFFSR_75 INVX1_4/gnd DFFSR_51/S FILL
XFILL_42_DFFSR_104 INVX1_4/gnd DFFSR_4/S FILL
XFILL_32_DFFSR_107 BUFX2_36/A DFFSR_8/S FILL
XFILL_1_DFFPOSX1_24 BUFX2_43/A DFFSR_23/S FILL
XFILL_22_DFFSR_110 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_12_DFFSR_113 INVX1_23/gnd DFFSR_186/S FILL
XFILL_6_BUFX2_20 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_5_NAND2X1_1 INVX1_2/gnd DFFSR_51/S FILL
XFILL_2_INVX1_264 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_44_DFFSR_3 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_8_DFFSR_107 BUFX2_36/A DFFSR_8/S FILL
XFILL_32_DFFSR_82 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_4_INVX1_76 INVX1_2/gnd DFFSR_1/S FILL
XFILL_43_DFFSR_42 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_5_OAI21X1_223 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_49_DFFSR_138 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_39_DFFSR_141 INVX1_94/gnd DFFSR_25/S FILL
XFILL_22_3 INVX1_94/gnd DFFSR_25/S FILL
XFILL_29_DFFSR_144 INVX1_8/gnd DFFSR_5/S FILL
XFILL_16_DFFSR_32 INVX1_2/gnd DFFSR_1/S FILL
XFILL_19_DFFSR_147 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_6_OAI21X1_157 BUFX2_35/A DFFSR_97/S FILL
XNOR2X1_29 NOR2X1_29/A NOR2X1_29/B BUFX2_37/A NOR2X1_29/Y DFFSR_81/S NOR2X1
XFILL_40_DFFSR_89 DFFSR_89/gnd DFFSR_92/S FILL
XOAI21X1_193 AOI21X1_5/Y AOI21X1_4/Y INVX1_233/Y BUFX2_7/gnd AOI22X1_4/C DFFSR_54/S
+ OAI21X1
XFILL_4_NOR2X1_26 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_6_NAND2X1_271 INVX1_89/gnd DFFSR_2/S FILL
XFILL_3_INVX1_408 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_7_DFFSR_46 BUFX2_36/A DFFSR_6/S FILL
XFILL_24_DFFSR_39 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_13_DFFSR_79 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_5_DFFSR_144 INVX1_8/gnd DFFSR_5/S FILL
XFILL_46_DFFSR_175 INVX1_23/gnd DFFSR_91/S FILL
XFILL_4_OAI21X1_253 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_36_DFFSR_178 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_26_DFFSR_181 INVX1_23/gnd DFFSR_186/S FILL
XFILL_2_INVX1_228 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_8_CLKBUF1_11 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_48_DFFSR_96 INVX1_2/gnd DFFSR_1/S FILL
XFILL_10_DFFSR_1 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_16_DFFSR_184 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_6_NAND3X1_103 INVX1_23/gnd DFFSR_186/S FILL
XFILL_7_CLKBUF1_14 BUFX2_43/A DFFSR_23/S FILL
XFILL_32_DFFSR_46 BUFX2_36/A DFFSR_6/S FILL
XFILL_5_OAI21X1_187 BUFX2_37/A DFFSR_8/S FILL
XFILL_6_CLKBUF1_17 INVX1_94/gnd DFFSR_25/S FILL
XFILL_21_DFFSR_86 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_4_DFFSR_93 INVX1_2/gnd DFFSR_51/S FILL
XFILL_49_DFFSR_102 INVX1_8/gnd DFFSR_7/S FILL
XFILL_43_1_0 INVX1_4/gnd DFFSR_51/S FILL
XFILL_5_CLKBUF1_20 INVX1_4/gnd DFFSR_51/S FILL
XFILL_39_DFFSR_105 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_2_DFFSR_181 INVX1_23/gnd DFFSR_186/S FILL
XFILL_5_7 BUFX2_6/gnd DFFSR_91/S FILL
XCLKBUF1_17 INVX1_402/Y INVX1_94/gnd DFFSR_52/CLK DFFSR_25/S CLKBUF1
XFILL_4_CLKBUF1_23 INVX1_89/gnd DFFSR_2/S FILL
XFILL_29_DFFSR_108 INVX1_89/gnd DFFSR_2/S FILL
XFILL_3_BUFX2_31 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_6_OAI21X1_121 BUFX2_36/A DFFSR_8/S FILL
XFILL_19_DFFSR_111 INVX1_8/gnd DFFSR_5/S FILL
XFILL_41_3_1 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_2_NAND2X1_2 INVX1_8/gnd DFFSR_5/S FILL
XFILL_40_DFFSR_53 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_1_INVX1_87 INVX1_89/gnd DFFSR_36/S FILL
XFILL_29_DFFSR_93 INVX1_2/gnd DFFSR_51/S FILL
XFILL_39_5_2 BUFX2_16/gnd DFFSR_65/S FILL
XOAI21X1_157 DFFSR_23/S INVX1_188/Y OAI21X1_157/C BUFX2_35/A DFFSR_157/D DFFSR_97/S
+ OAI21X1
XFILL_0_DFFPOSX1_18 BUFX2_37/A DFFSR_8/S FILL
XFILL_6_NAND2X1_235 INVX1_4/gnd DFFSR_51/S FILL
XFILL_13_DFFSR_43 INVX1_94/gnd DFFSR_25/S FILL
XFILL_7_DFFSR_10 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_5_DFFSR_108 INVX1_89/gnd DFFSR_2/S FILL
XFILL_3_INVX1_372 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_2_OAI22X1_1 BUFX2_36/A DFFSR_8/S FILL
XFILL_5_NAND3X1_133 INVX1_8/gnd DFFSR_5/S FILL
XFILL_46_DFFSR_139 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_36_DFFSR_142 BUFX2_19/gnd DFFSR_54/S FILL
XNAND2X1_271 XOR2X1_17/A DFFSR_137/Q INVX1_89/gnd XOR2X1_10/B DFFSR_2/S NAND2X1
XFILL_26_DFFSR_145 INVX1_23/gnd DFFSR_186/S FILL
XFILL_4_OAI21X1_217 INVX1_23/gnd DFFSR_91/S FILL
XFILL_16_DFFSR_148 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_2_INVX1_192 BUFX2_35/A DFFSR_14/S FILL
XFILL_48_DFFSR_60 BUFX2_37/A DFFSR_8/S FILL
XFILL_44_3 INVX1_4/gnd DFFSR_51/S FILL
XFILL_19_DFFPOSX1_26 BUFX2_37/A DFFSR_81/S FILL
XFILL_32_DFFSR_10 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_4_DFFSR_57 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_10_DFFSR_90 INVX1_2/gnd DFFSR_1/S FILL
XFILL_21_DFFSR_50 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_5_OAI21X1_151 BUFX2_37/A DFFSR_81/S FILL
XFILL_1_NOR2X1_27 BUFX2_17/gnd DFFSR_57/S FILL
XNAND3X1_103 NAND3X1_101/Y NAND3X1_102/Y INVX1_260/Y INVX1_23/gnd AOI21X1_32/A DFFSR_186/S
+ NAND3X1
XFILL_0_INVX1_409 INVX1_2/gnd DFFSR_51/S FILL
XFILL_2_DFFSR_145 INVX1_23/gnd DFFSR_186/S FILL
XFILL_5_NAND2X1_265 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_43_DFFSR_176 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_33_DFFSR_179 INVX1_2/gnd DFFSR_1/S FILL
XFILL_1_INVX1_51 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_23_DFFSR_182 INVX1_89/gnd DFFSR_36/S FILL
XFILL_40_DFFSR_17 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_29_DFFSR_57 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_13_DFFSR_185 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_18_DFFSR_97 BUFX2_35/A DFFSR_97/S FILL
XOAI21X1_121 BUFX2_20/Y INVX1_137/Y NAND2X1_121/Y BUFX2_36/A DFFSR_121/D DFFSR_8/S
+ OAI21X1
XFILL_3_INVX1_336 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_6_NAND2X1_199 BUFX2_36/A DFFSR_8/S FILL
XFILL_3_OAI21X1_247 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_0_BUFX2_42 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_46_DFFSR_103 INVX1_8/gnd DFFSR_7/S FILL
XFILL_9_DFFSR_179 INVX1_2/gnd DFFSR_1/S FILL
XFILL_4_OAI21X1_181 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_36_DFFSR_106 DFFSR_1/gnd DFFSR_1/S FILL
XNAND2X1_235 NOR2X1_15/Y NOR2X1_14/Y INVX1_4/gnd NAND2X1_66/B DFFSR_51/S NAND2X1
XFILL_26_DFFSR_109 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_2_INVX1_156 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_16_DFFSR_112 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_48_DFFSR_24 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_37_DFFSR_64 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_15_1_1 BUFX2_37/A DFFSR_81/S FILL
XFILL_21_DFFSR_14 BUFX2_35/A DFFSR_14/S FILL
XFILL_5_OAI21X1_115 BUFX2_36/A DFFSR_6/S FILL
XFILL_10_DFFSR_54 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_4_DFFSR_21 INVX1_2/gnd DFFSR_1/S FILL
XFILL_13_3_2 BUFX2_36/A DFFSR_8/S FILL
XFILL_2_DFFSR_109 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_3_NOR2X1_2 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_0_INVX1_373 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_43_DFFSR_140 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_22_DFFSR_4 INVX1_4/gnd DFFSR_4/S FILL
XFILL_5_NAND2X1_229 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_33_DFFSR_143 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_45_DFFSR_71 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_23_DFFSR_146 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_4_NAND3X1_127 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_13_DFFSR_149 INVX1_23/gnd DFFSR_91/S FILL
XFILL_1_DFFSR_68 BUFX2_35/A DFFSR_14/S FILL
XFILL_18_DFFSR_61 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_29_DFFSR_21 INVX1_2/gnd DFFSR_1/S FILL
XFILL_1_INVX1_15 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_6_BUFX2_5 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_3_OAI21X1_211 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_6_NAND2X1_163 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_3_INVX1_300 BUFX2_16/gnd DFFSR_11/S FILL
XNAND2X1_199 AND2X2_8/Y INVX1_224/Y BUFX2_36/A INVX1_238/A DFFSR_8/S NAND2X1
XFILL_9_DFFSR_143 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_4_OAI21X1_145 INVX1_23/gnd DFFSR_91/S FILL
XFILL_50_DFFSR_174 BUFX2_43/A DFFSR_97/S FILL
XFILL_18_DFFPOSX1_20 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_19_DFFPOSX1_2 INVX1_89/gnd DFFSR_36/S FILL
XFILL_26_DFFSR_68 BUFX2_35/A DFFSR_14/S FILL
XFILL_37_DFFSR_28 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_40_DFFSR_177 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_2_INVX1_120 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_9_DFFSR_75 INVX1_4/gnd DFFSR_51/S FILL
XFILL_30_DFFSR_180 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_18_DFFPOSX1_5 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_20_DFFSR_183 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_17_DFFPOSX1_8 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_10_DFFSR_18 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_4_NAND2X1_259 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_10_DFFSR_186 INVX1_23/gnd DFFSR_186/S FILL
XFILL_0_INVX1_337 BUFX2_36/A DFFSR_8/S FILL
XFILL_2_OAI21X1_241 BUFX2_35/A DFFSR_97/S FILL
XFILL_5_NAND2X1_193 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_45_DFFSR_35 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_6_DFFSR_180 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_8_DFFPOSX1_31 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_34_DFFSR_75 INVX1_4/gnd DFFSR_51/S FILL
XFILL_43_DFFSR_104 INVX1_4/gnd DFFSR_4/S FILL
XFILL_33_DFFSR_107 BUFX2_36/A DFFSR_8/S FILL
XFILL_1_DFFSR_32 INVX1_2/gnd DFFSR_1/S FILL
XFILL_23_DFFSR_110 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_13_DFFSR_113 INVX1_23/gnd DFFSR_186/S FILL
XFILL_18_DFFSR_25 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_6_NAND2X1_1 INVX1_2/gnd DFFSR_51/S FILL
XFILL_3_OAI21X1_175 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_6_NAND2X1_127 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_3_INVX1_264 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_10_OAI22X1_6 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_9_DFFSR_107 BUFX2_36/A DFFSR_8/S FILL
XXOR2X1_2 XOR2X1_2/A XOR2X1_2/B BUFX2_8/gnd OR2X2_1/A DFFSR_10/S XOR2X1
XFILL_42_DFFSR_82 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_4_OAI21X1_109 BUFX2_5/gnd DFFSR_6/S FILL
XNAND2X1_163 BUFX2_1/Y INVX1_229/A DFFSR_73/gnd NAND2X1_163/Y DFFSR_57/S NAND2X1
XFILL_48_3_1 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_50_DFFSR_138 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_40_DFFSR_141 INVX1_94/gnd DFFSR_25/S FILL
XFILL_9_DFFSR_39 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_30_DFFSR_144 INVX1_8/gnd DFFSR_5/S FILL
XFILL_15_DFFSR_72 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_46_5_2 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_26_DFFSR_32 INVX1_2/gnd DFFSR_1/S FILL
XFILL_20_DFFSR_147 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_4_NAND2X1_223 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_50_DFFSR_89 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_2_XOR2X1_9 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_10_DFFSR_150 BUFX2_8/gnd DFFSR_25/S FILL
XINVX1_411 INVX1_411/A DFFSR_89/gnd INVX1_411/Y DFFSR_186/S INVX1
XFILL_0_INVX1_301 INVX1_89/gnd DFFSR_2/S FILL
XFILL_3_NAND3X1_121 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_5_NOR2X1_26 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_2_OAI21X1_205 BUFX2_36/A DFFSR_8/S FILL
XFILL_5_NAND2X1_157 BUFX2_35/A DFFSR_97/S FILL
XFILL_34_DFFSR_39 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_23_DFFSR_79 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_6_DFFSR_144 INVX1_8/gnd DFFSR_5/S FILL
XFILL_6_DFFSR_86 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_47_DFFSR_175 INVX1_23/gnd DFFSR_91/S FILL
XFILL_14_4_0 BUFX2_37/A DFFSR_8/S FILL
XFILL_8_OR2X2_3 BUFX2_43/A DFFSR_23/S FILL
XFILL_37_DFFSR_178 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_27_DFFSR_181 INVX1_23/gnd DFFSR_186/S FILL
XFILL_17_DFFPOSX1_14 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_3_OAI21X1_139 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_5_BUFX2_24 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_3_INVX1_228 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_34_DFFSR_7 INVX1_8/gnd DFFSR_7/S FILL
XFILL_17_DFFSR_184 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_9_AOI21X1_16 BUFX2_43/A DFFSR_23/S FILL
XNAND2X1_127 BUFX2_20/Y INVX1_134/A BUFX2_5/gnd OAI21X1_127/C DFFSR_6/S NAND2X1
XFILL_42_DFFSR_46 BUFX2_36/A DFFSR_6/S FILL
XFILL_3_INVX1_80 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_31_DFFSR_86 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_3_NAND2X1_253 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_8_AOI21X1_19 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_7_DFFPOSX1_2 INVX1_89/gnd DFFSR_36/S FILL
XFILL_50_DFFSR_102 INVX1_8/gnd DFFSR_7/S FILL
XFILL_40_DFFSR_105 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_9_4 BUFX2_43/A DFFSR_97/S FILL
XFILL_7_AOI21X1_22 BUFX2_43/A DFFSR_97/S FILL
XFILL_15_DFFSR_36 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_6_DFFPOSX1_5 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_3_DFFSR_181 INVX1_23/gnd DFFSR_186/S FILL
XFILL_6_AOI21X1_25 BUFX2_43/A DFFSR_97/S FILL
XFILL_5_DFFPOSX1_8 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_30_DFFSR_108 INVX1_89/gnd DFFSR_2/S FILL
XFILL_1_OAI21X1_235 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_4_NAND2X1_187 BUFX2_37/A DFFSR_8/S FILL
XFILL_7_DFFPOSX1_25 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_5_AOI21X1_28 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_20_DFFSR_111 INVX1_8/gnd DFFSR_5/S FILL
XDFFPOSX1_5 INVX1_229/A CLKBUF1_10/Y DFFPOSX1_5/D DFFSR_73/gnd DFFSR_11/S DFFPOSX1
XFILL_4_AOI21X1_31 INVX1_23/gnd DFFSR_186/S FILL
XAOI21X1_25 AOI21X1_25/A AOI22X1_8/D AOI21X1_25/C BUFX2_43/A AOI21X1_25/Y DFFSR_97/S
+ AOI21X1
XFILL_10_DFFSR_114 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_3_NAND2X1_2 INVX1_8/gnd DFFSR_5/S FILL
XFILL_3_AOI21X1_34 INVX1_94/gnd DFFSR_25/S FILL
XFILL_50_DFFSR_53 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_0_INVX1_265 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_39_DFFSR_93 INVX1_2/gnd DFFSR_51/S FILL
XINVX1_375 DFFSR_110/Q DFFSR_73/gnd INVX1_375/Y DFFSR_57/S INVX1
XFILL_2_AOI21X1_37 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_2_OAI21X1_169 BUFX2_36/A DFFSR_8/S FILL
XFILL_5_NAND2X1_121 BUFX2_36/A DFFSR_8/S FILL
XFILL_0_AND2X2_2 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_12_DFFSR_83 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_23_DFFSR_43 INVX1_94/gnd DFFSR_25/S FILL
XFILL_6_DFFSR_108 INVX1_89/gnd DFFSR_2/S FILL
XFILL_6_DFFSR_50 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_4_INVX1_372 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_3_OAI22X1_1 BUFX2_36/A DFFSR_8/S FILL
XFILL_1_AOI21X1_40 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_47_DFFSR_139 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_37_DFFSR_142 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_22_1_1 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_0_AOI21X1_43 BUFX2_17/gnd DFFSR_7/S FILL
XBUFX2_28 BUFX2_28/A DFFSR_89/gnd dout[2] DFFSR_186/S BUFX2
XFILL_27_DFFSR_145 INVX1_23/gnd DFFSR_186/S FILL
XFILL_4_0_0 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_2_NAND2X1_283 INVX1_89/gnd DFFSR_36/S FILL
XFILL_17_DFFSR_148 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_3_INVX1_192 BUFX2_35/A DFFSR_14/S FILL
XFILL_20_3_2 INVX1_94/gnd DFFSR_52/S FILL
XFILL_3_OAI21X1_103 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_9_OAI21X1_64 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_2_2_1 INVX1_23/gnd DFFSR_186/S FILL
XFILL_8_OAI21X1_67 INVX1_2/gnd DFFSR_1/S FILL
XFILL_8_AND2X2_9 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_3_DFFSR_97 BUFX2_35/A DFFSR_97/S FILL
XFILL_42_DFFSR_10 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_3_INVX1_44 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_6_NAND2X1_88 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_31_DFFSR_50 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_7_OAI21X1_70 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_0_OAI21X1_265 BUFX2_43/A DFFSR_97/S FILL
XFILL_5_NAND2X1_91 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_3_NAND2X1_217 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_2_NOR2X1_27 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_20_DFFSR_90 INVX1_2/gnd DFFSR_1/S FILL
XFILL_6_OAI21X1_73 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_0_4_2 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_5_OAI21X1_76 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_1_INVX1_409 INVX1_2/gnd DFFSR_51/S FILL
XNAND2X1_88 BUFX2_18/Y INVX1_90/A DFFSR_3/gnd NAND2X1_88/Y DFFSR_65/S NAND2X1
XFILL_4_NAND2X1_94 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_3_DFFSR_145 INVX1_23/gnd DFFSR_186/S FILL
XFILL_2_BUFX2_35 BUFX2_35/A DFFSR_14/S FILL
XFILL_3_NAND2X1_97 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_2_NAND3X1_115 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_4_OAI21X1_79 INVX1_89/gnd DFFSR_36/S FILL
XOAI21X1_73 BUFX2_16/Y INVX1_83/Y OAI21X1_73/C DFFSR_73/gnd DFFSR_73/D DFFSR_11/S
+ OAI21X1
XFILL_1_OAI21X1_199 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_3_OAI21X1_82 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_44_DFFSR_176 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_4_NAND2X1_151 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_2_OAI21X1_85 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_21_DFFSR_1 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_34_DFFSR_179 INVX1_2/gnd DFFSR_1/S FILL
XFILL_24_DFFSR_182 INVX1_89/gnd DFFSR_36/S FILL
XFILL_50_DFFSR_17 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_1_OAI21X1_88 INVX1_4/gnd DFFSR_4/S FILL
XFILL_14_DFFSR_185 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_28_DFFSR_97 BUFX2_35/A DFFSR_97/S FILL
XFILL_0_OAI21X1_91 BUFX2_43/A DFFSR_97/S FILL
XINVX1_339 DFFSR_105/Q BUFX2_36/A INVX1_339/Y DFFSR_8/S INVX1
XFILL_0_INVX1_91 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_0_INVX1_229 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_39_DFFSR_57 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_2_OAI21X1_133 BUFX2_7/gnd DFFSR_81/S FILL
XBUFX2_6 rst BUFX2_6/gnd BUFX2_6/Y DFFSR_14/S BUFX2
XFILL_6_DFFSR_14 BUFX2_35/A DFFSR_14/S FILL
XFILL_5_BUFX2_2 BUFX2_43/A DFFSR_23/S FILL
XFILL_12_DFFSR_47 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_47_DFFSR_103 INVX1_8/gnd DFFSR_7/S FILL
XFILL_37_DFFSR_106 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_27_DFFSR_109 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_0_DFFSR_182 INVX1_89/gnd DFFSR_36/S FILL
XFILL_2_NAND2X1_247 INVX1_8/gnd DFFSR_5/S FILL
XFILL_3_INVX1_156 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_8_OAI21X1_31 BUFX2_35/A DFFSR_97/S FILL
XFILL_17_DFFSR_112 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_47_DFFSR_64 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_6_NAND2X1_52 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_7_OAI21X1_34 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_0_NAND2X1_3 INVX1_4/gnd DFFSR_51/S FILL
XFILL_31_DFFSR_14 BUFX2_35/A DFFSR_14/S FILL
XFILL_3_DFFSR_61 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_20_DFFSR_54 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_0_OAI21X1_229 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_6_OAI21X1_37 INVX1_89/gnd DFFSR_2/S FILL
XFILL_5_NAND2X1_55 INVX1_89/gnd DFFSR_2/S FILL
XFILL_6_DFFPOSX1_19 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_3_NAND2X1_181 BUFX2_19/gnd DFFSR_52/S FILL
XNAND2X1_52 DFFSR_45/S INVX1_50/A DFFSR_71/gnd OAI21X1_52/C DFFSR_10/S NAND2X1
XFILL_4_NAND2X1_58 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_3_DFFSR_109 BUFX2_6/gnd DFFSR_14/S FILL
XOAI21X1_37 DFFSR_2/S INVX1_42/Y OAI21X1_37/C INVX1_89/gnd DFFSR_37/D DFFSR_2/S OAI21X1
XFILL_5_OAI21X1_40 INVX1_8/gnd DFFSR_7/S FILL
XFILL_1_INVX1_373 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_0_OAI22X1_2 BUFX2_36/A DFFSR_8/S FILL
XFILL_3_NAND2X1_61 BUFX2_37/A DFFSR_81/S FILL
XFILL_4_OAI21X1_43 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_44_DFFSR_140 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_4_NAND2X1_115 BUFX2_36/A DFFSR_6/S FILL
XFILL_3_OAI21X1_46 BUFX2_37/A DFFSR_81/S FILL
XFILL_34_DFFSR_143 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_1_OAI21X1_163 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_2_NAND2X1_64 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_24_DFFSR_146 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_1_NAND2X1_67 INVX1_2/gnd DFFSR_1/S FILL
XFILL_2_OAI21X1_49 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_28_DFFSR_61 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_0_INVX1_193 BUFX2_36/A DFFSR_6/S FILL
XFILL_0_INVX1_55 BUFX2_36/A DFFSR_8/S FILL
XFILL_1_OAI21X1_52 INVX1_94/gnd DFFSR_25/S FILL
XINVX1_303 DFFSR_61/Q INVX1_94/gnd INVX1_303/Y DFFSR_25/S INVX1
XFILL_0_NAND2X1_70 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_39_DFFSR_21 INVX1_2/gnd DFFSR_1/S FILL
XFILL_14_DFFSR_149 INVX1_23/gnd DFFSR_91/S FILL
XFILL_1_NAND2X1_277 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_0_OAI21X1_55 INVX1_89/gnd DFFSR_2/S FILL
XFILL_25_DFFPOSX1_27 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_4_INVX1_300 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_12_DFFSR_11 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_0_DFFSR_146 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_2_NAND2X1_211 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_51_DFFSR_174 BUFX2_43/A DFFSR_97/S FILL
XFILL_36_DFFSR_68 BUFX2_35/A DFFSR_14/S FILL
XFILL_47_DFFSR_28 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_41_DFFSR_177 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_3_INVX1_120 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_1_NAND3X1_109 BUFX2_36/A DFFSR_8/S FILL
XFILL_31_DFFSR_180 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_21_DFFSR_183 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_3_DFFSR_25 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_6_NAND2X1_16 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_20_DFFSR_18 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_11_DFFSR_186 INVX1_23/gnd DFFSR_186/S FILL
XFILL_3_NAND2X1_145 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_0_OAI21X1_193 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_9_OAI21X1_248 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_5_NAND2X1_19 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_1_INVX1_337 BUFX2_36/A DFFSR_8/S FILL
XFILL_4_NAND2X1_22 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_21_4_0 INVX1_94/gnd DFFSR_25/S FILL
XNAND2X1_16 DFFSR_45/S INVX1_9/A DFFSR_79/gnd NAND2X1_16/Y DFFSR_36/S NAND2X1
XFILL_11_OAI22X1_63 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_3_NAND2X1_25 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_2_NOR2X1_6 BUFX2_17/gnd DFFSR_57/S FILL
XDFFPOSX1_19 NAND2X1_170/B CLKBUF1_10/Y NAND2X1_254/Y BUFX2_16/gnd DFFSR_65/S DFFPOSX1
XFILL_1_OAI21X1_127 BUFX2_43/A DFFSR_23/S FILL
XFILL_12_DFFSR_8 BUFX2_36/A DFFSR_8/S FILL
XFILL_2_NAND2X1_28 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_3_OAI21X1_10 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_10_OAI22X1_66 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_44_DFFSR_75 INVX1_4/gnd DFFSR_51/S FILL
XFILL_44_DFFSR_104 INVX1_4/gnd DFFSR_4/S FILL
XFILL_1_5_0 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_1_NAND2X1_31 BUFX2_43/A DFFSR_97/S FILL
XFILL_34_DFFSR_107 BUFX2_36/A DFFSR_8/S FILL
XFILL_7_DFFSR_180 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_2_OAI21X1_13 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_8_NAND3X1_87 INVX1_94/gnd DFFSR_52/S FILL
XFILL_1_OAI21X1_16 INVX1_89/gnd DFFSR_36/S FILL
XFILL_0_NAND2X1_34 INVX1_2/gnd DFFSR_1/S FILL
XFILL_0_INVX1_19 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_24_DFFSR_110 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_14_DFFSR_113 INVX1_23/gnd DFFSR_186/S FILL
XFILL_7_NAND3X1_90 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_28_DFFSR_25 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_0_DFFSR_72 BUFX2_17/gnd DFFSR_7/S FILL
XINVX1_267 DFFSR_49/Q BUFX2_17/gnd INVX1_267/Y DFFSR_57/S INVX1
XFILL_0_OAI21X1_19 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_17_DFFSR_65 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_0_INVX1_157 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_6_NAND3X1_93 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_4_INVX1_264 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_1_NAND2X1_241 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_5_NAND3X1_96 BUFX2_43/A DFFSR_97/S FILL
XFILL_4_NAND3X1_99 BUFX2_6/gnd DFFSR_14/S FILL
XNAND3X1_93 INVX1_258/Y NAND3X1_90/B NAND3X1_90/C BUFX2_5/gnd NAND3X1_94/C DFFSR_23/S
+ NAND3X1
XFILL_4_XOR2X1_2 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_5_DFFPOSX1_13 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_33_DFFSR_4 INVX1_4/gnd DFFSR_4/S FILL
XFILL_2_NAND2X1_175 BUFX2_35/A DFFSR_14/S FILL
XFILL_13_2 BUFX2_36/A DFFSR_6/S FILL
XFILL_41_DFFSR_141 INVX1_94/gnd DFFSR_25/S FILL
XFILL_0_DFFSR_110 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_8_DFFSR_79 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_31_DFFSR_144 INVX1_8/gnd DFFSR_5/S FILL
XFILL_25_DFFSR_72 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_36_DFFSR_32 INVX1_2/gnd DFFSR_1/S FILL
XFILL_21_DFFSR_147 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_0_OAI21X1_157 BUFX2_35/A DFFSR_97/S FILL
XFILL_3_NAND2X1_109 INVX1_94/gnd DFFSR_25/S FILL
XFILL_11_DFFSR_150 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_1_INVX1_301 INVX1_89/gnd DFFSR_2/S FILL
XFILL_29_1_1 INVX1_89/gnd DFFSR_2/S FILL
XFILL_6_NOR2X1_26 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_0_AOI22X1_12 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_10_OAI22X1_30 INVX1_94/gnd DFFSR_25/S FILL
XFILL_9_NAND3X1_48 BUFX2_43/A DFFSR_23/S FILL
XFILL_24_DFFPOSX1_21 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_44_DFFSR_39 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_27_3_2 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_33_DFFSR_79 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_0_NAND2X1_271 INVX1_89/gnd DFFSR_2/S FILL
XFILL_7_DFFSR_144 INVX1_8/gnd DFFSR_5/S FILL
XFILL_48_DFFSR_175 INVX1_23/gnd DFFSR_91/S FILL
XINVX1_231 AND2X2_8/B BUFX2_43/A INVX1_231/Y DFFSR_23/S INVX1
XFILL_9_2_1 BUFX2_43/A DFFSR_23/S FILL
XFILL_0_INVX1_121 BUFX2_36/A DFFSR_6/S FILL
XFILL_8_NAND3X1_51 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_0_DFFSR_36 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_9_OAI22X1_33 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_38_DFFSR_178 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_17_DFFSR_29 INVX1_4/gnd DFFSR_4/S FILL
XFILL_28_DFFSR_181 INVX1_23/gnd DFFSR_186/S FILL
XFILL_1_NAND2X1_205 BUFX2_36/A DFFSR_6/S FILL
XFILL_7_NAND3X1_54 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_8_OAI22X1_36 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_7_4_2 BUFX2_35/A DFFSR_97/S FILL
XFILL_7_OAI22X1_39 BUFX2_37/A DFFSR_8/S FILL
XFILL_6_NAND3X1_57 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_18_DFFSR_184 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_0_NAND3X1_103 INVX1_23/gnd DFFSR_186/S FILL
XNAND3X1_57 NOR3X1_1/B NAND3X1_52/Y NAND3X1_53/Y BUFX2_19/gnd NAND3X1_57/Y DFFSR_54/S
+ NAND3X1
XFILL_5_NAND3X1_60 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_6_OAI22X1_42 INVX1_8/gnd DFFSR_7/S FILL
XFILL_4_NAND3X1_63 BUFX2_43/A DFFSR_23/S FILL
XFILL_5_OAI22X1_45 INVX1_89/gnd DFFSR_2/S FILL
XOAI22X1_42 INVX1_342/Y OAI22X1_40/D INVX1_343/Y OAI22X1_38/D INVX1_8/gnd NOR2X1_30/A
+ DFFSR_7/S OAI22X1
XFILL_41_DFFSR_86 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_3_NAND3X1_66 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_8_OAI21X1_242 BUFX2_35/A DFFSR_97/S FILL
XFILL_4_OAI22X1_48 BUFX2_37/A DFFSR_81/S FILL
XFILL_2_NAND2X1_139 BUFX2_17/gnd DFFSR_57/S FILL
XDFFSR_184 BUFX2_26/A DFFSR_1/CLK DFFSR_185/R DFFSR_9/S DFFSR_184/D DFFSR_1/gnd DFFSR_9/S
+ DFFSR
XFILL_41_DFFSR_105 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_2_NAND3X1_69 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_3_OAI22X1_51 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_14_DFFSR_76 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_8_DFFSR_43 INVX1_94/gnd DFFSR_25/S FILL
XFILL_25_DFFSR_36 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_4_DFFSR_181 INVX1_23/gnd DFFSR_186/S FILL
XFILL_1_NAND3X1_72 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_2_OAI22X1_54 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_31_DFFSR_108 INVX1_89/gnd DFFSR_2/S FILL
XFILL_0_NAND3X1_75 BUFX2_35/A DFFSR_97/S FILL
XFILL_21_DFFSR_111 INVX1_8/gnd DFFSR_5/S FILL
XNAND2X1_5 DFFSR_5/S NAND2X1_5/B INVX1_8/gnd OAI21X1_5/C DFFSR_7/S NAND2X1
XFILL_1_OAI22X1_57 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_0_OAI21X1_121 BUFX2_36/A DFFSR_8/S FILL
XFILL_9_OAI21X1_176 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_11_DFFSR_114 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_4_NAND2X1_2 INVX1_8/gnd DFFSR_5/S FILL
XFILL_0_OAI22X1_60 INVX1_8/gnd DFFSR_5/S FILL
XFILL_1_INVX1_265 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_0_DFFSR_7 INVX1_8/gnd DFFSR_7/S FILL
XFILL_49_DFFSR_93 INVX1_2/gnd DFFSR_51/S FILL
XINVX1_77 DFFSR_68/Q BUFX2_37/A INVX1_77/Y DFFSR_81/S INVX1
XOAI22X1_4 OAI22X1_4/A OAI22X1_4/B OAI22X1_4/C OAI22X1_4/D BUFX2_7/gnd OAI22X1_4/Y
+ DFFSR_54/S OAI22X1
XFILL_22_DFFSR_83 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_33_DFFSR_43 INVX1_94/gnd DFFSR_25/S FILL
XFILL_7_DFFSR_108 INVX1_89/gnd DFFSR_2/S FILL
XFILL_5_DFFSR_90 INVX1_2/gnd DFFSR_1/S FILL
XFILL_0_NAND2X1_235 INVX1_4/gnd DFFSR_51/S FILL
XFILL_4_OAI22X1_1 BUFX2_36/A DFFSR_8/S FILL
XFILL_48_DFFSR_139 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_38_DFFSR_142 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_8_NAND3X1_15 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_4_BUFX2_28 DFFSR_89/gnd DFFSR_186/S FILL
XINVX1_195 DFFSR_161/Q INVX1_23/gnd INVX1_195/Y DFFSR_186/S INVX1
XFILL_28_DFFSR_145 INVX1_23/gnd DFFSR_186/S FILL
XFILL_7_NAND3X1_18 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_4_INVX1_192 BUFX2_35/A DFFSR_14/S FILL
XFILL_1_NAND2X1_169 BUFX2_36/A DFFSR_8/S FILL
XFILL_6_NAND3X1_21 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_35_2 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_18_DFFSR_148 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_5_NAND3X1_24 BUFX2_37/A DFFSR_8/S FILL
XFILL_4_NAND3X1_27 BUFX2_37/A DFFSR_81/S FILL
XNAND3X1_21 BUFX2_14/Y AND2X2_6/B NAND3X1_21/C BUFX2_7/gnd NAND3X1_22/B DFFSR_81/S
+ NAND3X1
XFILL_2_INVX1_84 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_41_DFFSR_50 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_13_DFFPOSX1_26 BUFX2_37/A DFFSR_81/S FILL
XFILL_3_NAND3X1_30 INVX1_94/gnd DFFSR_52/S FILL
XFILL_3_NOR2X1_27 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_30_DFFSR_90 INVX1_2/gnd DFFSR_1/S FILL
XFILL_4_OAI22X1_12 INVX1_4/gnd DFFSR_51/S FILL
XDFFSR_148 DFFSR_148/Q CLKBUF1_12/Y DFFSR_148/R DFFSR_92/S DFFSR_148/D DFFSR_89/gnd
+ DFFSR_92/S DFFSR
XFILL_8_OAI21X1_206 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_2_NAND2X1_103 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_2_NAND3X1_33 INVX1_8/gnd DFFSR_7/S FILL
XFILL_2_INVX1_409 INVX1_2/gnd DFFSR_51/S FILL
XFILL_3_OAI22X1_15 INVX1_4/gnd DFFSR_4/S FILL
XFILL_4_DFFSR_145 INVX1_23/gnd DFFSR_186/S FILL
XFILL_1_NAND3X1_36 BUFX2_35/A DFFSR_97/S FILL
XFILL_14_DFFSR_40 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_2_OAI22X1_18 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_45_DFFSR_176 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_23_DFFPOSX1_15 BUFX2_35/A DFFSR_14/S FILL
XFILL_0_NAND3X1_39 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_35_DFFSR_179 INVX1_2/gnd DFFSR_1/S FILL
XFILL_1_OAI22X1_21 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_0_OAI22X1_24 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_25_DFFSR_182 INVX1_89/gnd DFFSR_36/S FILL
XFILL_45_DFFSR_7 INVX1_8/gnd DFFSR_7/S FILL
XFILL_15_DFFSR_185 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_38_DFFSR_97 BUFX2_35/A DFFSR_97/S FILL
XFILL_1_INVX1_229 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_49_DFFSR_57 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_0_NAND2X1_199 BUFX2_36/A DFFSR_8/S FILL
XFILL_5_DFFSR_54 BUFX2_7/gnd DFFSR_81/S FILL
XINVX1_41 INVX1_41/A DFFSR_79/gnd INVX1_41/Y DFFSR_45/S INVX1
XFILL_22_DFFSR_47 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_11_DFFSR_87 DFFSR_3/gnd DFFSR_4/S FILL
XDFFSR_94 DFFSR_94/Q CLKBUF1_5/Y DFFSR_89/R DFFSR_4/S DFFSR_94/D BUFX2_16/gnd DFFSR_65/S
+ DFFSR
XFILL_48_DFFSR_103 INVX1_8/gnd DFFSR_7/S FILL
XFILL_0_INVX1_9 BUFX2_36/A DFFSR_6/S FILL
XINVX1_159 INVX1_159/A INVX1_94/gnd INVX1_159/Y DFFSR_52/S INVX1
XFILL_38_DFFSR_106 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_28_DFFSR_109 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_1_NAND2X1_133 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_1_DFFSR_182 INVX1_89/gnd DFFSR_36/S FILL
XFILL_7_OAI21X1_236 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_28_4_0 INVX1_89/gnd DFFSR_36/S FILL
XFILL_18_DFFSR_112 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_4_INVX1_156 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_1_NAND2X1_3 INVX1_4/gnd DFFSR_51/S FILL
XFILL_41_DFFSR_14 BUFX2_35/A DFFSR_14/S FILL
XFILL_30_DFFSR_54 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_19_DFFSR_94 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_2_INVX1_48 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_8_OAI21X1_170 INVX1_94/gnd DFFSR_25/S FILL
XDFFSR_112 INVX1_391/A CLKBUF1_4/Y DFFSR_105/R DFFSR_65/S DFFSR_112/D DFFSR_3/gnd
+ DFFSR_65/S DFFSR
XFILL_8_5_0 BUFX2_43/A DFFSR_97/S FILL
XFILL_2_INVX1_373 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_4_DFFSR_109 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_1_BUFX2_39 BUFX2_43/A DFFSR_97/S FILL
XFILL_1_OAI22X1_2 BUFX2_36/A DFFSR_8/S FILL
XFILL_45_DFFSR_140 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_35_DFFSR_143 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_25_DFFSR_146 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_11_DFFSR_5 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_9_OAI21X1_104 INVX1_4/gnd DFFSR_51/S FILL
XFILL_38_DFFSR_61 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_1_INVX1_193 BUFX2_36/A DFFSR_6/S FILL
XFILL_49_DFFSR_21 INVX1_2/gnd DFFSR_1/S FILL
XFILL_15_DFFSR_149 INVX1_23/gnd DFFSR_91/S FILL
XFILL_0_NAND2X1_163 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_5_DFFSR_18 DFFSR_9/gnd DFFSR_9/S FILL
XDFFSR_58 INVX1_66/A DFFSR_15/CLK DFFSR_61/R DFFSR_4/S DFFSR_58/D DFFSR_3/gnd DFFSR_4/S
+ DFFSR
XFILL_22_DFFSR_11 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_0_NOR2X1_28 INVX1_94/gnd DFFSR_52/S FILL
XFILL_11_DFFSR_51 INVX1_2/gnd DFFSR_51/S FILL
XFILL_8_NAND3X1_116 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_1_DFFSR_146 DFFSR_89/gnd DFFSR_92/S FILL
XINVX1_123 DFFSR_109/Q BUFX2_5/gnd INVX1_123/Y DFFSR_6/S INVX1
XFILL_12_DFFPOSX1_20 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_46_DFFSR_68 BUFX2_35/A DFFSR_14/S FILL
XFILL_7_OAI21X1_200 BUFX2_37/A DFFSR_8/S FILL
XFILL_42_DFFSR_177 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_32_DFFSR_1 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_4_INVX1_120 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_32_DFFSR_180 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_36_1_1 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_22_DFFSR_183 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_2_INVX1_12 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_2_DFFSR_65 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_12_DFFSR_186 INVX1_23/gnd DFFSR_186/S FILL
XFILL_30_DFFSR_18 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_19_DFFSR_58 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_2_INVX1_337 BUFX2_36/A DFFSR_8/S FILL
XFILL_8_OAI21X1_134 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_34_3_2 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_2_DFFPOSX1_31 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_45_DFFSR_104 INVX1_4/gnd DFFSR_4/S FILL
XFILL_35_DFFSR_107 BUFX2_36/A DFFSR_8/S FILL
XFILL_8_DFFSR_180 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_25_DFFSR_110 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_15_DFFSR_113 INVX1_23/gnd DFFSR_186/S FILL
XFILL_38_DFFSR_25 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_27_DFFSR_65 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_1_INVX1_157 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_6_OAI21X1_230 INVX1_23/gnd DFFSR_186/S FILL
XFILL_0_NAND2X1_127 BUFX2_5/gnd DFFSR_6/S FILL
XDFFSR_22 INVX1_25/A DFFSR_28/CLK DFFSR_20/R DFFSR_10/S DFFSR_22/D BUFX2_8/gnd DFFSR_10/S
+ DFFSR
XFILL_11_DFFSR_15 INVX1_8/gnd DFFSR_7/S FILL
XFILL_42_DFFSR_141 INVX1_94/gnd DFFSR_25/S FILL
XFILL_7_OAI21X1_164 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_1_DFFSR_110 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_32_DFFSR_144 INVX1_8/gnd DFFSR_5/S FILL
XFILL_35_DFFSR_72 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_46_DFFSR_32 INVX1_2/gnd DFFSR_1/S FILL
XFILL_22_DFFSR_147 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_19_DFFSR_22 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_2_DFFSR_29 INVX1_4/gnd DFFSR_4/S FILL
XFILL_12_DFFSR_150 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_2_INVX1_301 INVX1_89/gnd DFFSR_2/S FILL
XFILL_20_CLKBUF1_12 BUFX2_43/A DFFSR_23/S FILL
XFILL_43_DFFSR_79 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_8_DFFSR_144 INVX1_8/gnd DFFSR_5/S FILL
XFILL_19_CLKBUF1_15 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_5_OAI21X1_260 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_49_DFFSR_175 INVX1_23/gnd DFFSR_91/S FILL
XFILL_18_CLKBUF1_18 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_16_DFFSR_69 BUFX2_43/A DFFSR_23/S FILL
XFILL_1_INVX1_121 BUFX2_36/A DFFSR_6/S FILL
XFILL_17_CLKBUF1_21 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_39_DFFSR_178 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_27_DFFSR_29 INVX1_4/gnd DFFSR_4/S FILL
XFILL_16_CLKBUF1_24 INVX1_23/gnd DFFSR_186/S FILL
XFILL_29_DFFSR_181 INVX1_23/gnd DFFSR_186/S FILL
XFILL_11_DFFPOSX1_14 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_7_NAND3X1_110 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_6_OAI21X1_194 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_19_DFFSR_184 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_3_XOR2X1_6 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_23_DFFSR_8 BUFX2_36/A DFFSR_8/S FILL
XOAI21X1_230 INVX1_247/Y XNOR2X1_3/A AOI22X1_13/A INVX1_23/gnd XOR2X1_6/A DFFSR_186/S
+ OAI21X1
XFILL_42_DFFSR_105 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_24_DFFSR_76 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_7_DFFSR_83 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_7_OAI21X1_128 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_35_DFFSR_36 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_5_DFFSR_181 INVX1_23/gnd DFFSR_186/S FILL
XFILL_32_DFFSR_108 INVX1_89/gnd DFFSR_2/S FILL
XFILL_22_DFFSR_111 INVX1_8/gnd DFFSR_5/S FILL
XFILL_6_BUFX2_21 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_1_DFFPOSX1_25 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_12_DFFSR_114 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_5_NAND2X1_2 INVX1_8/gnd DFFSR_5/S FILL
XFILL_2_INVX1_265 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_44_DFFSR_4 INVX1_4/gnd DFFSR_4/S FILL
XFILL_4_INVX1_77 BUFX2_37/A DFFSR_81/S FILL
XFILL_32_DFFSR_83 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_43_DFFSR_43 INVX1_94/gnd DFFSR_25/S FILL
XFILL_5_OAI21X1_224 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_5_OAI22X1_1 BUFX2_36/A DFFSR_8/S FILL
XFILL_8_DFFSR_108 INVX1_89/gnd DFFSR_2/S FILL
XFILL_35_4_0 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_49_DFFSR_139 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_39_DFFSR_142 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_29_DFFSR_145 INVX1_23/gnd DFFSR_186/S FILL
XFILL_16_DFFSR_33 INVX1_94/gnd DFFSR_52/S FILL
XFILL_22_4 INVX1_94/gnd DFFSR_25/S FILL
XFILL_19_DFFSR_148 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_6_OAI21X1_158 BUFX2_43/A DFFSR_97/S FILL
XNOR2X1_30 NOR2X1_30/A NOR2X1_30/B DFFSR_73/gnd NOR2X1_30/Y DFFSR_57/S NOR2X1
XOAI21X1_194 INVX1_224/A AOI21X1_6/Y NAND3X1_9/Y BUFX2_19/gnd AOI21X1_7/C DFFSR_54/S
+ OAI21X1
XFILL_4_NOR2X1_27 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_40_DFFSR_90 INVX1_2/gnd DFFSR_1/S FILL
XFILL_51_DFFSR_50 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_3_INVX1_409 INVX1_2/gnd DFFSR_51/S FILL
XFILL_6_NAND2X1_272 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_5_DFFSR_145 INVX1_23/gnd DFFSR_186/S FILL
XFILL_7_DFFSR_47 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_24_DFFSR_40 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_13_DFFSR_80 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_46_DFFSR_176 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_36_DFFSR_179 INVX1_2/gnd DFFSR_1/S FILL
XFILL_4_OAI21X1_254 INVX1_23/gnd DFFSR_91/S FILL
XFILL_26_DFFSR_182 INVX1_89/gnd DFFSR_36/S FILL
XFILL_16_DFFSR_185 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_48_DFFSR_97 BUFX2_35/A DFFSR_97/S FILL
XFILL_8_CLKBUF1_12 BUFX2_43/A DFFSR_23/S FILL
XFILL_2_INVX1_229 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_10_DFFSR_2 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_6_NAND3X1_104 INVX1_23/gnd DFFSR_186/S FILL
XFILL_7_CLKBUF1_15 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_6_CLKBUF1_18 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_5_OAI21X1_188 INVX1_89/gnd DFFSR_2/S FILL
XFILL_32_DFFSR_47 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_21_DFFSR_87 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_4_DFFSR_94 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_49_DFFSR_103 INVX1_8/gnd DFFSR_7/S FILL
XFILL_5_CLKBUF1_21 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_4_CLKBUF1_24 INVX1_23/gnd DFFSR_186/S FILL
XFILL_5_8 BUFX2_6/gnd DFFSR_91/S FILL
XCLKBUF1_18 INVX1_402/Y BUFX2_8/gnd DFFSR_3/CLK DFFSR_25/S CLKBUF1
XFILL_39_DFFSR_106 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_43_1_1 INVX1_4/gnd DFFSR_51/S FILL
XFILL_29_DFFSR_109 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_2_DFFSR_182 INVX1_89/gnd DFFSR_36/S FILL
XFILL_3_BUFX2_32 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_6_OAI21X1_122 INVX1_94/gnd DFFSR_25/S FILL
XFILL_41_3_2 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_19_DFFSR_112 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_2_NAND2X1_3 INVX1_4/gnd DFFSR_51/S FILL
XFILL_40_DFFSR_54 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_1_INVX1_88 INVX1_2/gnd DFFSR_1/S FILL
XFILL_29_DFFSR_94 BUFX2_16/gnd DFFSR_65/S FILL
XOAI21X1_158 DFFSR_158/S INVX1_190/Y NAND2X1_158/Y BUFX2_43/A DFFSR_158/D DFFSR_97/S
+ OAI21X1
XFILL_0_DFFPOSX1_19 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_13_DFFSR_44 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_3_INVX1_373 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_7_DFFSR_11 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_5_DFFSR_109 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_2_OAI22X1_2 BUFX2_36/A DFFSR_8/S FILL
XFILL_5_NAND3X1_134 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_46_DFFSR_140 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_36_DFFSR_143 BUFX2_8/gnd DFFSR_25/S FILL
XNAND2X1_272 NOR2X1_46/A INVX1_156/A BUFX2_16/gnd NAND2X1_272/Y DFFSR_11/S NAND2X1
XFILL_4_OAI21X1_218 INVX1_23/gnd DFFSR_186/S FILL
XFILL_26_DFFSR_146 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_48_DFFSR_61 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_2_INVX1_193 BUFX2_36/A DFFSR_6/S FILL
XFILL_16_DFFSR_149 INVX1_23/gnd DFFSR_91/S FILL
XFILL_44_4 INVX1_4/gnd DFFSR_51/S FILL
XFILL_4_DFFSR_58 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_32_DFFSR_11 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_10_DFFSR_91 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_5_OAI21X1_152 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_1_NOR2X1_28 INVX1_94/gnd DFFSR_52/S FILL
XFILL_19_DFFPOSX1_27 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_21_DFFSR_51 INVX1_2/gnd DFFSR_51/S FILL
XNAND3X1_104 INVX1_260/A NAND3X1_101/Y NAND3X1_102/Y INVX1_23/gnd AOI21X1_33/B DFFSR_186/S
+ NAND3X1
XFILL_0_INVX1_410 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_2_DFFSR_146 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_43_DFFSR_177 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_5_NAND2X1_266 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_33_DFFSR_180 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_23_DFFSR_183 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_13_DFFSR_186 INVX1_23/gnd DFFSR_186/S FILL
XFILL_1_INVX1_52 BUFX2_37/A DFFSR_81/S FILL
XOAI21X1_122 BUFX2_19/Y INVX1_138/Y NAND2X1_122/Y INVX1_94/gnd DFFSR_122/D DFFSR_25/S
+ OAI21X1
XFILL_18_DFFSR_98 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_40_DFFSR_18 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_29_DFFSR_58 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_6_NAND2X1_200 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_3_INVX1_337 BUFX2_36/A DFFSR_8/S FILL
XFILL_3_OAI21X1_248 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_0_BUFX2_43 BUFX2_35/A DFFSR_97/S FILL
XFILL_46_DFFSR_104 INVX1_4/gnd DFFSR_4/S FILL
XFILL_36_DFFSR_107 BUFX2_36/A DFFSR_8/S FILL
XFILL_9_DFFSR_180 BUFX2_17/gnd DFFSR_7/S FILL
XNAND2X1_236 NOR2X1_17/Y NOR2X1_16/Y INVX1_2/gnd NAND2X1_67/B DFFSR_1/S NAND2X1
XFILL_4_OAI21X1_182 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_26_DFFSR_110 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_16_DFFSR_113 INVX1_23/gnd DFFSR_186/S FILL
XFILL_48_DFFSR_25 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_37_DFFSR_65 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_2_INVX1_157 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_15_1_2 BUFX2_37/A DFFSR_81/S FILL
XFILL_4_DFFSR_22 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_10_DFFSR_55 INVX1_89/gnd DFFSR_36/S FILL
XFILL_5_OAI21X1_116 INVX1_89/gnd DFFSR_2/S FILL
XFILL_21_DFFSR_15 INVX1_8/gnd DFFSR_7/S FILL
XFILL_0_INVX1_374 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_3_NOR2X1_3 INVX1_94/gnd DFFSR_25/S FILL
XFILL_43_DFFSR_141 INVX1_94/gnd DFFSR_25/S FILL
XFILL_22_DFFSR_5 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_2_DFFSR_110 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_5_NAND2X1_230 BUFX2_36/A DFFSR_6/S FILL
XFILL_33_DFFSR_144 INVX1_8/gnd DFFSR_5/S FILL
XFILL_45_DFFSR_72 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_23_DFFSR_147 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_1_INVX1_16 BUFX2_43/A DFFSR_23/S FILL
XFILL_1_DFFSR_69 BUFX2_43/A DFFSR_23/S FILL
XFILL_18_DFFSR_62 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_29_DFFSR_22 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_4_NAND3X1_128 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_6_BUFX2_6 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_3_OAI21X1_212 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_13_DFFSR_150 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_3_INVX1_301 INVX1_89/gnd DFFSR_2/S FILL
XFILL_6_NAND2X1_164 INVX1_8/gnd DFFSR_5/S FILL
XFILL_42_4_0 INVX1_4/gnd DFFSR_4/S FILL
XNAND2X1_200 AND2X2_11/A INVX1_246/A BUFX2_6/gnd INVX1_239/A DFFSR_14/S NAND2X1
XFILL_9_DFFSR_144 INVX1_8/gnd DFFSR_5/S FILL
XFILL_43_DFFSR_1 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_4_OAI21X1_146 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_50_DFFSR_175 INVX1_23/gnd DFFSR_91/S FILL
XFILL_18_DFFPOSX1_21 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_26_DFFSR_69 BUFX2_43/A DFFSR_23/S FILL
XFILL_2_INVX1_121 BUFX2_36/A DFFSR_6/S FILL
XFILL_9_DFFSR_76 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_19_DFFPOSX1_3 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_40_DFFSR_178 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_37_DFFSR_29 INVX1_4/gnd DFFSR_4/S FILL
XFILL_30_DFFSR_181 INVX1_23/gnd DFFSR_186/S FILL
XFILL_18_DFFPOSX1_6 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_17_DFFPOSX1_9 BUFX2_37/A DFFSR_8/S FILL
XFILL_20_DFFSR_184 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_4_NAND2X1_260 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_10_DFFSR_19 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_10_DFFSR_187 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_0_INVX1_338 BUFX2_36/A DFFSR_8/S FILL
XFILL_43_DFFSR_105 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_2_OAI21X1_242 BUFX2_35/A DFFSR_97/S FILL
XFILL_5_NAND2X1_194 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_34_DFFSR_76 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_45_DFFSR_36 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_6_DFFSR_181 INVX1_23/gnd DFFSR_186/S FILL
XFILL_33_DFFSR_108 INVX1_89/gnd DFFSR_2/S FILL
XFILL_23_DFFSR_111 INVX1_8/gnd DFFSR_5/S FILL
XFILL_1_DFFSR_33 INVX1_94/gnd DFFSR_52/S FILL
XFILL_13_DFFSR_114 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_6_NAND2X1_2 INVX1_8/gnd DFFSR_5/S FILL
XFILL_18_DFFSR_26 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_3_OAI21X1_176 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_3_INVX1_265 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_6_NAND2X1_128 INVX1_89/gnd DFFSR_2/S FILL
XFILL_10_OAI22X1_7 DFFSR_5/gnd DFFSR_5/S FILL
XXOR2X1_3 XOR2X1_3/A XOR2X1_3/B BUFX2_17/gnd XOR2X1_3/Y DFFSR_7/S XOR2X1
XFILL_6_OAI22X1_1 BUFX2_36/A DFFSR_8/S FILL
XFILL_42_DFFSR_83 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_9_DFFSR_108 INVX1_89/gnd DFFSR_2/S FILL
XNAND2X1_164 BUFX2_3/Y INVX1_235/A INVX1_8/gnd OAI21X1_164/C DFFSR_5/S NAND2X1
XFILL_48_3_2 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_50_DFFSR_139 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_4_OAI21X1_110 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_40_DFFSR_142 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_26_DFFSR_33 INVX1_94/gnd DFFSR_52/S FILL
XFILL_26_1 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_9_DFFSR_40 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_15_DFFSR_73 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_30_DFFSR_145 INVX1_23/gnd DFFSR_186/S FILL
XFILL_20_DFFSR_148 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_4_NAND2X1_224 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_10_DFFSR_151 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_16_2_0 BUFX2_7/gnd DFFSR_81/S FILL
XINVX1_412 INVX1_412/A DFFSR_79/gnd INVX1_412/Y DFFSR_36/S INVX1
XFILL_3_NAND3X1_122 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_0_INVX1_302 INVX1_8/gnd DFFSR_7/S FILL
XFILL_5_NOR2X1_27 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_50_DFFSR_90 INVX1_2/gnd DFFSR_1/S FILL
XFILL_2_OAI21X1_206 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_6_DFFSR_145 INVX1_23/gnd DFFSR_186/S FILL
XFILL_5_NAND2X1_158 BUFX2_35/A DFFSR_97/S FILL
XFILL_34_DFFSR_40 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_6_DFFSR_87 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_23_DFFSR_80 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_14_4_1 BUFX2_37/A DFFSR_8/S FILL
XFILL_47_DFFSR_176 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_37_DFFSR_179 INVX1_2/gnd DFFSR_1/S FILL
XFILL_17_DFFPOSX1_15 BUFX2_35/A DFFSR_14/S FILL
XFILL_5_BUFX2_25 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_3_OAI21X1_140 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_27_DFFSR_182 INVX1_89/gnd DFFSR_36/S FILL
XFILL_17_DFFSR_185 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_3_INVX1_229 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_34_DFFSR_8 BUFX2_36/A DFFSR_8/S FILL
XNAND2X1_128 BUFX2_22/Y INVX1_390/A INVX1_89/gnd OAI21X1_128/C DFFSR_2/S NAND2X1
XFILL_42_DFFSR_47 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_3_INVX1_81 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_31_DFFSR_87 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_8_AOI21X1_20 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_3_NAND2X1_254 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_7_DFFPOSX1_3 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_50_DFFSR_103 INVX1_8/gnd DFFSR_7/S FILL
XFILL_7_AOI21X1_23 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_15_DFFSR_37 INVX1_89/gnd DFFSR_2/S FILL
XFILL_40_DFFSR_106 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_6_DFFPOSX1_6 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_30_DFFSR_109 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_6_AOI21X1_26 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_5_DFFPOSX1_9 BUFX2_37/A DFFSR_8/S FILL
XFILL_3_DFFSR_182 INVX1_89/gnd DFFSR_36/S FILL
XFILL_1_OAI21X1_236 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_7_DFFPOSX1_26 BUFX2_37/A DFFSR_81/S FILL
XFILL_5_AOI21X1_29 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_4_NAND2X1_188 INVX1_8/gnd DFFSR_7/S FILL
XFILL_20_DFFSR_112 DFFSR_3/gnd DFFSR_65/S FILL
XDFFPOSX1_6 INVX1_235/A CLKBUF1_10/Y DFFPOSX1_6/D DFFSR_3/gnd DFFSR_65/S DFFPOSX1
XFILL_10_DFFSR_115 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_4_AOI21X1_32 BUFX2_43/A DFFSR_23/S FILL
XAOI21X1_26 AOI21X1_26/A NAND3X1_73/Y AOI21X1_26/C BUFX2_5/gnd AOI21X1_26/Y DFFSR_23/S
+ AOI21X1
XFILL_3_NAND2X1_3 INVX1_4/gnd DFFSR_51/S FILL
XFILL_50_DFFSR_54 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_0_INVX1_266 BUFX2_8/gnd DFFSR_10/S FILL
XINVX1_376 INVX1_376/A INVX1_8/gnd INVX1_376/Y DFFSR_7/S INVX1
XFILL_39_DFFSR_94 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_3_AOI21X1_35 INVX1_94/gnd DFFSR_25/S FILL
XFILL_2_AOI21X1_38 BUFX2_36/A DFFSR_8/S FILL
XFILL_2_OAI21X1_170 INVX1_94/gnd DFFSR_25/S FILL
XFILL_5_NAND2X1_122 INVX1_94/gnd DFFSR_25/S FILL
XFILL_23_DFFSR_44 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_0_AND2X2_3 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_6_DFFSR_51 INVX1_2/gnd DFFSR_51/S FILL
XFILL_6_DFFSR_109 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_1_AOI21X1_41 BUFX2_35/A DFFSR_14/S FILL
XFILL_12_DFFSR_84 BUFX2_43/A DFFSR_23/S FILL
XFILL_3_OAI22X1_2 BUFX2_36/A DFFSR_8/S FILL
XFILL_47_DFFSR_140 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_37_DFFSR_143 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_22_1_2 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_0_AOI21X1_44 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_4_0_1 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_2_NAND2X1_284 INVX1_8/gnd DFFSR_5/S FILL
XBUFX2_29 BUFX2_29/A BUFX2_16/gnd dout[3] DFFSR_65/S BUFX2
XFILL_27_DFFSR_146 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_3_INVX1_193 BUFX2_36/A DFFSR_6/S FILL
XFILL_3_OAI21X1_104 INVX1_4/gnd DFFSR_51/S FILL
XFILL_17_DFFSR_149 INVX1_23/gnd DFFSR_91/S FILL
XFILL_8_OAI21X1_68 BUFX2_37/A DFFSR_81/S FILL
XFILL_48_1 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_2_2_2 INVX1_23/gnd DFFSR_186/S FILL
XFILL_6_NAND2X1_89 BUFX2_37/A DFFSR_8/S FILL
XFILL_7_OAI21X1_71 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_3_INVX1_45 INVX1_8/gnd DFFSR_5/S FILL
XFILL_42_DFFSR_11 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_20_DFFSR_91 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_5_NAND2X1_92 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_2_NOR2X1_28 INVX1_94/gnd DFFSR_52/S FILL
XFILL_3_NAND2X1_218 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_6_OAI21X1_74 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_3_DFFSR_98 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_31_DFFSR_51 INVX1_2/gnd DFFSR_51/S FILL
XNAND2X1_89 DFFSR_81/Q BUFX2_20/Y BUFX2_37/A OAI21X1_89/C DFFSR_8/S NAND2X1
XFILL_5_OAI21X1_77 INVX1_89/gnd DFFSR_36/S FILL
XFILL_4_NAND2X1_95 INVX1_89/gnd DFFSR_36/S FILL
XFILL_1_INVX1_410 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_3_DFFSR_146 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_2_BUFX2_36 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_2_NAND3X1_116 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_3_NAND2X1_98 DFFSR_1/gnd DFFSR_9/S FILL
XOAI21X1_74 BUFX2_18/Y INVX1_84/Y NAND2X1_74/Y DFFSR_9/gnd DFFSR_74/D DFFSR_9/S OAI21X1
XFILL_4_OAI21X1_80 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_3_OAI21X1_83 INVX1_94/gnd DFFSR_52/S FILL
XFILL_44_DFFSR_177 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_4_NAND2X1_152 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_1_OAI21X1_200 BUFX2_37/A DFFSR_8/S FILL
XFILL_34_DFFSR_180 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_2_OAI21X1_86 INVX1_4/gnd DFFSR_51/S FILL
XFILL_24_DFFSR_183 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_1_OAI21X1_89 BUFX2_35/A DFFSR_14/S FILL
XFILL_21_DFFSR_2 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_14_DFFSR_186 INVX1_23/gnd DFFSR_186/S FILL
XFILL_0_INVX1_92 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_0_INVX1_230 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_28_DFFSR_98 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_50_DFFSR_18 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_39_DFFSR_58 DFFSR_3/gnd DFFSR_4/S FILL
XINVX1_340 INVX1_75/A DFFSR_3/gnd INVX1_340/Y DFFSR_65/S INVX1
XFILL_0_OAI21X1_92 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_4_INVX1_337 BUFX2_36/A DFFSR_8/S FILL
XFILL_2_OAI21X1_134 DFFSR_79/gnd DFFSR_36/S FILL
XBUFX2_7 rst BUFX2_7/gnd BUFX2_7/Y DFFSR_81/S BUFX2
XFILL_5_BUFX2_3 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_6_DFFSR_15 INVX1_8/gnd DFFSR_7/S FILL
XFILL_12_DFFSR_48 INVX1_4/gnd DFFSR_4/S FILL
XFILL_47_DFFSR_104 INVX1_4/gnd DFFSR_4/S FILL
XFILL_37_DFFSR_107 BUFX2_36/A DFFSR_8/S FILL
XFILL_0_DFFSR_183 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_2_NAND2X1_248 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_27_DFFSR_110 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_17_DFFSR_113 INVX1_23/gnd DFFSR_186/S FILL
XFILL_8_OAI21X1_32 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_47_DFFSR_65 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_3_INVX1_157 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_0_NAND2X1_4 INVX1_2/gnd DFFSR_51/S FILL
XFILL_0_OAI21X1_230 INVX1_23/gnd DFFSR_186/S FILL
XFILL_6_DFFPOSX1_20 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_3_DFFSR_62 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_6_NAND2X1_53 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_20_DFFSR_55 INVX1_89/gnd DFFSR_36/S FILL
XFILL_7_OAI21X1_35 INVX1_8/gnd DFFSR_5/S FILL
XFILL_31_DFFSR_15 INVX1_8/gnd DFFSR_7/S FILL
XFILL_3_NAND2X1_182 BUFX2_8/gnd DFFSR_25/S FILL
XNAND2X1_53 DFFSR_45/S DFFSR_45/Q DFFSR_79/gnd OAI21X1_53/C DFFSR_45/S NAND2X1
XFILL_6_OAI21X1_38 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_5_NAND2X1_56 INVX1_4/gnd DFFSR_51/S FILL
XOAI21X1_38 DFFSR_5/S INVX1_43/Y OAI21X1_38/C DFFSR_5/gnd DFFSR_38/D DFFSR_5/S OAI21X1
XFILL_5_OAI21X1_41 INVX1_8/gnd DFFSR_7/S FILL
XFILL_1_INVX1_374 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_4_NAND2X1_59 INVX1_2/gnd DFFSR_1/S FILL
XFILL_3_NAND2X1_62 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_44_DFFSR_141 INVX1_94/gnd DFFSR_25/S FILL
XFILL_4_OAI21X1_44 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_0_OAI22X1_3 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_3_DFFSR_110 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_4_NAND2X1_116 INVX1_89/gnd DFFSR_36/S FILL
XFILL_3_OAI21X1_47 INVX1_89/gnd DFFSR_2/S FILL
XFILL_1_OAI21X1_164 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_2_NAND2X1_65 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_1_NAND2X1_68 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_34_DFFSR_144 INVX1_8/gnd DFFSR_5/S FILL
XFILL_2_OAI21X1_50 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_24_DFFSR_147 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_28_DFFSR_62 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_39_DFFSR_22 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_0_NAND2X1_71 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_1_OAI21X1_53 DFFSR_71/gnd DFFSR_45/S FILL
XINVX1_304 DFFSR_45/Q DFFSR_79/gnd INVX1_304/Y DFFSR_36/S INVX1
XFILL_0_INVX1_194 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_0_INVX1_56 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_14_DFFSR_150 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_0_OAI21X1_56 INVX1_2/gnd DFFSR_51/S FILL
XFILL_1_NAND2X1_278 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_4_INVX1_301 INVX1_89/gnd DFFSR_2/S FILL
XFILL_25_DFFPOSX1_28 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_12_DFFSR_12 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_0_DFFSR_147 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_2_NAND2X1_212 INVX1_23/gnd DFFSR_186/S FILL
XFILL_36_DFFSR_69 BUFX2_43/A DFFSR_23/S FILL
XFILL_3_INVX1_121 BUFX2_36/A DFFSR_6/S FILL
XFILL_41_DFFSR_178 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_47_DFFSR_29 INVX1_4/gnd DFFSR_4/S FILL
XFILL_31_DFFSR_181 INVX1_23/gnd DFFSR_186/S FILL
XFILL_1_NAND3X1_110 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_23_2_0 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_6_NAND2X1_17 INVX1_8/gnd DFFSR_7/S FILL
XFILL_21_DFFSR_184 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_3_DFFSR_26 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_9_OAI21X1_249 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_5_NAND2X1_20 INVX1_23/gnd DFFSR_186/S FILL
XFILL_3_NAND2X1_146 INVX1_23/gnd DFFSR_91/S FILL
XFILL_0_OAI21X1_194 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_20_DFFSR_19 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_11_DFFSR_187 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_4_NAND2X1_23 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_1_INVX1_338 BUFX2_36/A DFFSR_8/S FILL
XFILL_21_4_1 INVX1_94/gnd DFFSR_25/S FILL
XNAND2X1_17 DFFSR_9/Q DFFSR_57/S INVX1_8/gnd OAI21X1_17/C DFFSR_7/S NAND2X1
XFILL_2_NOR2X1_7 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_3_3_0 INVX1_23/gnd DFFSR_91/S FILL
XFILL_11_OAI22X1_64 INVX1_94/gnd DFFSR_25/S FILL
XFILL_9_DFFSR_1 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_3_NAND2X1_26 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_44_DFFSR_105 DFFSR_89/gnd DFFSR_186/S FILL
XDFFPOSX1_20 DFFPOSX1_20/Q CLKBUF1_16/Y INVX1_405/Y BUFX2_7/gnd DFFSR_54/S DFFPOSX1
XFILL_44_DFFSR_76 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_12_DFFSR_9 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_2_NAND2X1_29 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_10_OAI22X1_67 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_3_OAI21X1_11 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_7_DFFSR_181 INVX1_23/gnd DFFSR_186/S FILL
XFILL_2_OAI21X1_14 BUFX2_43/A DFFSR_23/S FILL
XFILL_1_OAI21X1_128 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_34_DFFSR_108 INVX1_89/gnd DFFSR_2/S FILL
XFILL_1_NAND2X1_32 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_1_5_1 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_8_NAND3X1_88 INVX1_94/gnd DFFSR_52/S FILL
XFILL_1_OAI21X1_17 INVX1_8/gnd DFFSR_5/S FILL
XFILL_24_DFFSR_111 INVX1_8/gnd DFFSR_5/S FILL
XFILL_0_NAND2X1_35 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_7_NAND3X1_91 BUFX2_43/A DFFSR_97/S FILL
XFILL_14_DFFSR_114 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_0_INVX1_158 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_0_INVX1_20 INVX1_8/gnd DFFSR_5/S FILL
XINVX1_268 DFFSR_17/Q INVX1_8/gnd INVX1_268/Y DFFSR_7/S INVX1
XFILL_28_DFFSR_26 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_17_DFFSR_66 INVX1_2/gnd DFFSR_51/S FILL
XFILL_0_DFFSR_73 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_0_OAI21X1_20 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_6_NAND3X1_94 BUFX2_35/A DFFSR_97/S FILL
XFILL_1_NAND2X1_242 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_4_INVX1_265 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_11_OAI22X1_7 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_5_NAND3X1_97 BUFX2_35/A DFFSR_97/S FILL
XFILL_7_OR2X2_1 BUFX2_8/gnd DFFSR_10/S FILL
XNAND3X1_94 XOR2X1_7/Y NAND3X1_94/B NAND3X1_94/C BUFX2_35/A NAND3X1_95/A DFFSR_97/S
+ NAND3X1
XFILL_4_XOR2X1_3 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_5_DFFPOSX1_14 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_7_OAI22X1_1 BUFX2_36/A DFFSR_8/S FILL
XFILL_33_DFFSR_5 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_51_DFFSR_139 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_2_NAND2X1_176 INVX1_94/gnd DFFSR_25/S FILL
XFILL_0_DFFSR_111 INVX1_8/gnd DFFSR_5/S FILL
XFILL_41_DFFSR_142 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_36_DFFSR_33 INVX1_94/gnd DFFSR_52/S FILL
XFILL_8_DFFSR_80 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_25_DFFSR_73 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_31_DFFSR_145 INVX1_23/gnd DFFSR_186/S FILL
XFILL_21_DFFSR_148 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_0_OAI21X1_158 BUFX2_43/A DFFSR_97/S FILL
XFILL_11_DFFSR_151 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_3_NAND2X1_110 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_1_AOI22X1_10 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_29_1_2 INVX1_89/gnd DFFSR_2/S FILL
XFILL_1_INVX1_302 INVX1_8/gnd DFFSR_7/S FILL
XFILL_6_NOR2X1_27 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_10_OAI22X1_31 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_0_AOI22X1_13 INVX1_23/gnd DFFSR_186/S FILL
XFILL_7_DFFSR_145 INVX1_23/gnd DFFSR_186/S FILL
XFILL_44_DFFSR_40 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_33_DFFSR_80 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_0_NAND2X1_272 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_24_DFFPOSX1_22 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_48_DFFSR_176 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_9_2_2 BUFX2_43/A DFFSR_23/S FILL
XFILL_8_NAND3X1_52 BUFX2_36/A DFFSR_8/S FILL
XINVX1_232 OAI22X1_2/C BUFX2_37/A AOI22X1_5/D DFFSR_8/S INVX1
XFILL_0_INVX1_122 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_17_DFFSR_30 INVX1_89/gnd DFFSR_36/S FILL
XFILL_0_DFFSR_37 INVX1_89/gnd DFFSR_2/S FILL
XFILL_38_DFFSR_179 INVX1_2/gnd DFFSR_1/S FILL
XFILL_9_OAI22X1_34 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_7_NAND3X1_55 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_8_OAI22X1_37 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_28_DFFSR_182 INVX1_89/gnd DFFSR_36/S FILL
XFILL_18_DFFSR_185 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_1_NAND2X1_206 BUFX2_43/A DFFSR_97/S FILL
XFILL_7_OAI22X1_40 BUFX2_37/A DFFSR_8/S FILL
XFILL_6_NAND3X1_58 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_4_INVX1_229 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_0_NAND3X1_104 INVX1_23/gnd DFFSR_186/S FILL
XFILL_6_OAI22X1_43 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_5_NAND3X1_61 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_4_NAND3X1_64 BUFX2_35/A DFFSR_14/S FILL
XNAND3X1_58 NAND3X1_58/A NAND3X1_56/Y NAND3X1_57/Y BUFX2_19/gnd NAND3X1_58/Y DFFSR_54/S
+ NAND3X1
XFILL_5_OAI22X1_46 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_41_DFFSR_87 DFFSR_3/gnd DFFSR_4/S FILL
XDFFSR_185 BUFX2_27/A DFFSR_20/CLK DFFSR_185/R DFFSR_92/S DFFSR_185/D DFFSR_89/gnd
+ DFFSR_92/S DFFSR
XFILL_3_NAND3X1_67 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_8_OAI21X1_243 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_4_OAI22X1_49 INVX1_94/gnd DFFSR_25/S FILL
XOAI22X1_43 INVX1_345/Y OAI22X1_40/B INVX1_344/Y OAI22X1_38/B BUFX2_8/gnd NOR2X1_31/A
+ DFFSR_25/S OAI22X1
XFILL_2_NAND2X1_140 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_51_DFFSR_103 INVX1_8/gnd DFFSR_7/S FILL
XFILL_2_NAND3X1_70 BUFX2_35/A DFFSR_14/S FILL
XFILL_3_OAI22X1_52 INVX1_94/gnd DFFSR_25/S FILL
XFILL_8_DFFSR_44 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_25_DFFSR_37 INVX1_89/gnd DFFSR_2/S FILL
XFILL_14_DFFSR_77 INVX1_89/gnd DFFSR_2/S FILL
XFILL_41_DFFSR_106 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_31_DFFSR_109 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_1_NAND3X1_73 BUFX2_43/A DFFSR_23/S FILL
XFILL_2_OAI22X1_55 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_4_DFFSR_182 INVX1_89/gnd DFFSR_36/S FILL
XNAND2X1_6 DFFSR_186/S INVX1_411/A INVX1_23/gnd NAND2X1_6/Y DFFSR_186/S NAND2X1
XFILL_0_NAND3X1_76 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_1_OAI22X1_58 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_21_DFFSR_112 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_11_DFFSR_115 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_0_OAI21X1_122 INVX1_94/gnd DFFSR_25/S FILL
XFILL_9_OAI21X1_177 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_0_OAI22X1_61 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_4_NAND2X1_3 INVX1_4/gnd DFFSR_51/S FILL
XFILL_0_DFFSR_8 BUFX2_36/A DFFSR_8/S FILL
XFILL_1_INVX1_266 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_49_DFFSR_94 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_5_DFFSR_91 BUFX2_6/gnd DFFSR_91/S FILL
XINVX1_78 DFFSR_69/Q BUFX2_36/A INVX1_78/Y DFFSR_8/S INVX1
XFILL_0_NAND2X1_236 INVX1_2/gnd DFFSR_1/S FILL
XOAI22X1_5 OAI22X1_5/A OAI22X1_9/B OAI22X1_5/C OAI22X1_9/D BUFX2_16/gnd NOR2X1_12/B
+ DFFSR_65/S OAI22X1
XFILL_7_DFFSR_109 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_22_DFFSR_84 BUFX2_43/A DFFSR_23/S FILL
XFILL_4_OAI22X1_2 BUFX2_36/A DFFSR_8/S FILL
XFILL_33_DFFSR_44 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_48_DFFSR_140 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_8_NAND3X1_16 BUFX2_19/gnd DFFSR_52/S FILL
XINVX1_196 DFFSR_162/Q DFFSR_89/gnd INVX1_196/Y DFFSR_186/S INVX1
XFILL_38_DFFSR_143 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_7_NAND3X1_19 INVX1_8/gnd DFFSR_5/S FILL
XFILL_4_BUFX2_29 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_28_DFFSR_146 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_4_INVX1_193 BUFX2_36/A DFFSR_6/S FILL
XFILL_6_NAND3X1_22 BUFX2_37/A DFFSR_81/S FILL
XFILL_35_3 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_1_NAND2X1_170 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_18_DFFSR_149 INVX1_23/gnd DFFSR_91/S FILL
XFILL_5_NAND3X1_25 BUFX2_7/gnd DFFSR_81/S FILL
XNAND3X1_22 OAI22X1_2/C NAND3X1_22/B NAND3X1_22/C BUFX2_37/A AOI21X1_5/B DFFSR_81/S
+ NAND3X1
XFILL_4_NAND3X1_28 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_5_OAI22X1_10 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_30_DFFSR_91 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_3_NAND3X1_31 INVX1_94/gnd DFFSR_52/S FILL
XFILL_3_NOR2X1_28 INVX1_94/gnd DFFSR_52/S FILL
XFILL_13_DFFPOSX1_27 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_41_DFFSR_51 INVX1_2/gnd DFFSR_51/S FILL
XFILL_2_INVX1_85 DFFSR_3/gnd DFFSR_65/S FILL
XDFFSR_149 DFFSR_149/Q CLKBUF1_12/Y DFFSR_149/R DFFSR_91/S DFFSR_149/D INVX1_23/gnd
+ DFFSR_91/S DFFSR
XFILL_8_OAI21X1_207 BUFX2_37/A DFFSR_8/S FILL
XFILL_2_NAND2X1_104 INVX1_4/gnd DFFSR_51/S FILL
XFILL_4_OAI22X1_13 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_2_INVX1_410 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_4_DFFSR_146 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_14_DFFSR_41 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_2_NAND3X1_34 INVX1_2/gnd DFFSR_1/S FILL
XFILL_3_OAI22X1_16 INVX1_4/gnd DFFSR_4/S FILL
XFILL_1_NAND3X1_37 BUFX2_43/A DFFSR_97/S FILL
XFILL_2_OAI22X1_19 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_45_DFFSR_177 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_0_NAND3X1_40 BUFX2_43/A DFFSR_23/S FILL
XFILL_35_DFFSR_180 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_1_OAI22X1_22 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_25_DFFSR_183 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_23_DFFPOSX1_16 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_45_DFFSR_8 BUFX2_36/A DFFSR_8/S FILL
XFILL_0_OAI22X1_25 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_15_DFFSR_186 INVX1_23/gnd DFFSR_186/S FILL
XFILL_1_INVX1_230 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_38_DFFSR_98 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_49_DFFSR_58 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_0_NAND2X1_200 BUFX2_6/gnd DFFSR_14/S FILL
XDFFSR_95 DFFSR_95/Q CLKBUF1_1/Y DFFSR_89/R DFFSR_45/S DFFSR_95/D DFFSR_79/gnd DFFSR_45/S
+ DFFSR
XINVX1_42 INVX1_42/A INVX1_89/gnd INVX1_42/Y DFFSR_36/S INVX1
XFILL_5_DFFSR_55 INVX1_89/gnd DFFSR_36/S FILL
XFILL_22_DFFSR_48 INVX1_4/gnd DFFSR_4/S FILL
XFILL_11_DFFSR_88 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_48_DFFSR_104 INVX1_4/gnd DFFSR_4/S FILL
XFILL_38_DFFSR_107 BUFX2_36/A DFFSR_8/S FILL
XINVX1_160 DFFSR_142/Q BUFX2_19/gnd INVX1_160/Y DFFSR_52/S INVX1
XFILL_30_2_0 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_1_DFFSR_183 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_1_NAND2X1_134 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_28_DFFSR_110 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_18_DFFSR_113 INVX1_23/gnd DFFSR_186/S FILL
XFILL_7_OAI21X1_237 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_28_4_1 INVX1_89/gnd DFFSR_36/S FILL
XFILL_4_INVX1_157 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_1_NAND2X1_4 INVX1_2/gnd DFFSR_51/S FILL
XFILL_2_INVX1_49 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_19_DFFSR_95 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_30_DFFSR_55 INVX1_89/gnd DFFSR_36/S FILL
XFILL_41_DFFSR_15 INVX1_8/gnd DFFSR_7/S FILL
XDFFSR_113 DFFSR_113/Q CLKBUF1_7/Y DFFSR_113/R DFFSR_186/S DFFSR_113/D INVX1_23/gnd
+ DFFSR_186/S DFFSR
XFILL_8_OAI21X1_171 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_8_5_1 BUFX2_43/A DFFSR_97/S FILL
XFILL_2_INVX1_374 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_1_BUFX2_40 BUFX2_35/A DFFSR_14/S FILL
XFILL_1_OAI22X1_3 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_4_DFFSR_110 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_45_DFFSR_141 INVX1_94/gnd DFFSR_25/S FILL
XFILL_11_DFFSR_6 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_35_DFFSR_144 INVX1_8/gnd DFFSR_5/S FILL
XFILL_25_DFFSR_147 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_38_DFFSR_62 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_49_DFFSR_22 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_1_INVX1_194 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_15_DFFSR_150 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_0_NAND2X1_164 INVX1_8/gnd DFFSR_5/S FILL
XFILL_5_DFFSR_19 DFFSR_1/gnd DFFSR_9/S FILL
XDFFSR_59 INVX1_67/A DFFSR_15/CLK DFFSR_61/R DFFSR_51/S DFFSR_59/D INVX1_4/gnd DFFSR_51/S
+ DFFSR
XFILL_22_DFFSR_12 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_0_NOR2X1_29 BUFX2_37/A DFFSR_81/S FILL
XFILL_11_DFFSR_52 INVX1_94/gnd DFFSR_52/S FILL
XFILL_1_DFFSR_147 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_12_DFFPOSX1_21 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_8_NAND3X1_117 INVX1_94/gnd DFFSR_25/S FILL
XINVX1_124 DFFSR_110/Q DFFSR_73/gnd INVX1_124/Y DFFSR_57/S INVX1
XFILL_7_OAI21X1_201 BUFX2_35/A DFFSR_97/S FILL
XFILL_46_DFFSR_69 BUFX2_43/A DFFSR_23/S FILL
XFILL_4_INVX1_121 BUFX2_36/A DFFSR_6/S FILL
XFILL_32_DFFSR_2 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_42_DFFSR_178 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_32_DFFSR_181 INVX1_23/gnd DFFSR_186/S FILL
XFILL_22_DFFSR_184 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_36_1_2 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_30_DFFSR_19 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_2_DFFSR_66 INVX1_2/gnd DFFSR_51/S FILL
XFILL_19_DFFSR_59 INVX1_4/gnd DFFSR_51/S FILL
XFILL_2_INVX1_13 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_12_DFFSR_187 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_8_OAI21X1_135 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_2_INVX1_338 BUFX2_36/A DFFSR_8/S FILL
XFILL_22_DFFPOSX1_10 INVX1_8/gnd DFFSR_5/S FILL
XFILL_45_DFFSR_105 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_8_DFFSR_181 INVX1_23/gnd DFFSR_186/S FILL
XFILL_35_DFFSR_108 INVX1_89/gnd DFFSR_2/S FILL
XFILL_25_DFFSR_111 INVX1_8/gnd DFFSR_5/S FILL
XFILL_15_DFFSR_114 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_1_INVX1_158 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_38_DFFSR_26 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_27_DFFSR_66 INVX1_2/gnd DFFSR_51/S FILL
XDFFSR_23 INVX1_26/A DFFSR_20/CLK DFFSR_20/R DFFSR_23/S DFFSR_23/D BUFX2_5/gnd DFFSR_23/S
+ DFFSR
XFILL_6_OAI21X1_231 BUFX2_36/A DFFSR_6/S FILL
XFILL_11_DFFSR_16 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_0_NAND2X1_128 INVX1_89/gnd DFFSR_2/S FILL
XFILL_8_OAI22X1_1 BUFX2_36/A DFFSR_8/S FILL
XFILL_1_DFFSR_111 INVX1_8/gnd DFFSR_5/S FILL
XFILL_7_OAI21X1_165 BUFX2_35/A DFFSR_97/S FILL
XFILL_42_DFFSR_142 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_46_DFFSR_33 INVX1_94/gnd DFFSR_52/S FILL
XFILL_35_DFFSR_73 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_32_DFFSR_145 INVX1_23/gnd DFFSR_186/S FILL
XFILL_22_DFFSR_148 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_19_DFFSR_23 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_2_DFFSR_30 INVX1_89/gnd DFFSR_36/S FILL
XFILL_12_DFFSR_151 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_2_INVX1_302 INVX1_8/gnd DFFSR_7/S FILL
XFILL_20_CLKBUF1_13 INVX1_4/gnd DFFSR_51/S FILL
XFILL_8_DFFSR_145 INVX1_23/gnd DFFSR_186/S FILL
XFILL_19_CLKBUF1_16 BUFX2_36/A DFFSR_6/S FILL
XFILL_43_DFFSR_80 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_5_OAI21X1_261 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_18_CLKBUF1_19 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_49_DFFSR_176 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_17_CLKBUF1_22 INVX1_94/gnd DFFSR_25/S FILL
XFILL_1_INVX1_122 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_27_DFFSR_30 INVX1_89/gnd DFFSR_36/S FILL
XFILL_16_DFFSR_70 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_39_DFFSR_179 INVX1_2/gnd DFFSR_1/S FILL
XFILL_16_CLKBUF1_25 INVX1_23/gnd DFFSR_186/S FILL
XFILL_7_NAND3X1_111 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_29_DFFSR_182 INVX1_89/gnd DFFSR_36/S FILL
XFILL_19_DFFSR_185 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_11_DFFPOSX1_15 BUFX2_35/A DFFSR_14/S FILL
XFILL_6_OAI21X1_195 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_3_XOR2X1_7 INVX1_23/gnd DFFSR_91/S FILL
XFILL_23_DFFSR_9 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_51_DFFSR_87 DFFSR_3/gnd DFFSR_4/S FILL
XOAI21X1_231 NOR2X1_10/A NOR2X1_10/B XNOR2X1_2/Y BUFX2_36/A NAND3X1_92/A DFFSR_6/S
+ OAI21X1
XFILL_7_DFFSR_84 BUFX2_43/A DFFSR_23/S FILL
XFILL_35_DFFSR_37 INVX1_89/gnd DFFSR_2/S FILL
XFILL_42_DFFSR_106 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_7_OAI21X1_129 INVX1_4/gnd DFFSR_4/S FILL
XFILL_32_DFFSR_109 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_5_DFFSR_182 INVX1_89/gnd DFFSR_36/S FILL
XFILL_24_DFFSR_77 INVX1_89/gnd DFFSR_2/S FILL
XFILL_22_DFFSR_112 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_12_DFFSR_115 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_1_DFFPOSX1_26 BUFX2_37/A DFFSR_81/S FILL
XFILL_6_BUFX2_22 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_5_NAND2X1_3 INVX1_4/gnd DFFSR_51/S FILL
XFILL_2_INVX1_266 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_16_NOR3X1_1 INVX1_94/gnd DFFSR_52/S FILL
XFILL_44_DFFSR_5 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_37_2_0 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_5_OAI21X1_225 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_8_DFFSR_109 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_32_DFFSR_84 BUFX2_43/A DFFSR_23/S FILL
XFILL_5_OAI22X1_2 BUFX2_36/A DFFSR_8/S FILL
XFILL_4_INVX1_78 BUFX2_36/A DFFSR_8/S FILL
XFILL_43_DFFSR_44 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_49_DFFSR_140 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_35_4_1 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_22_5 INVX1_94/gnd DFFSR_25/S FILL
XFILL_39_DFFSR_143 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_16_DFFSR_34 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_29_DFFSR_146 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_19_DFFSR_149 INVX1_23/gnd DFFSR_91/S FILL
XFILL_6_OAI21X1_159 BUFX2_43/A DFFSR_97/S FILL
XNOR2X1_31 NOR2X1_31/A NOR2X1_31/B DFFSR_73/gnd NOR2X1_31/Y DFFSR_11/S NOR2X1
XFILL_40_DFFSR_91 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_4_NOR2X1_28 INVX1_94/gnd DFFSR_52/S FILL
XOAI21X1_195 AOI21X1_5/Y AOI21X1_4/Y INVX1_233/A BUFX2_7/gnd AOI21X1_7/B DFFSR_81/S
+ OAI21X1
XFILL_6_NAND2X1_273 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_3_INVX1_410 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_5_DFFSR_146 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_13_DFFSR_81 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_24_DFFSR_41 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_7_DFFSR_48 INVX1_4/gnd DFFSR_4/S FILL
XFILL_46_DFFSR_177 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_36_DFFSR_180 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_26_DFFSR_183 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_9_CLKBUF1_10 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_4_OAI21X1_255 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_16_DFFSR_186 INVX1_23/gnd DFFSR_186/S FILL
XFILL_2_INVX1_230 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_48_DFFSR_98 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_8_CLKBUF1_13 INVX1_4/gnd DFFSR_51/S FILL
XFILL_10_DFFSR_3 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_6_NAND3X1_105 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_7_CLKBUF1_16 BUFX2_36/A DFFSR_6/S FILL
XFILL_4_DFFSR_95 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_32_DFFSR_48 INVX1_4/gnd DFFSR_4/S FILL
XFILL_21_DFFSR_88 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_5_OAI21X1_189 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_6_CLKBUF1_19 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_49_DFFSR_104 INVX1_4/gnd DFFSR_4/S FILL
XFILL_39_DFFSR_107 BUFX2_36/A DFFSR_8/S FILL
XFILL_5_CLKBUF1_22 INVX1_94/gnd DFFSR_25/S FILL
XCLKBUF1_19 INVX1_402/Y DFFSR_9/gnd DFFSR_1/CLK DFFSR_9/S CLKBUF1
XFILL_43_1_2 INVX1_4/gnd DFFSR_51/S FILL
XFILL_3_BUFX2_33 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_2_DFFSR_183 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_4_CLKBUF1_25 INVX1_23/gnd DFFSR_186/S FILL
XFILL_29_DFFSR_110 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_19_DFFSR_113 INVX1_23/gnd DFFSR_186/S FILL
XFILL_6_OAI21X1_123 INVX1_23/gnd DFFSR_91/S FILL
XFILL_2_NAND2X1_4 INVX1_2/gnd DFFSR_51/S FILL
XFILL_29_DFFSR_95 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_40_DFFSR_55 INVX1_89/gnd DFFSR_36/S FILL
XFILL_1_INVX1_89 INVX1_89/gnd DFFSR_2/S FILL
XFILL_51_DFFSR_15 INVX1_8/gnd DFFSR_7/S FILL
XOAI21X1_159 DFFSR_23/S INVX1_192/Y NAND2X1_159/Y BUFX2_43/A DFFSR_159/D DFFSR_97/S
+ OAI21X1
XFILL_0_DFFPOSX1_20 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_7_DFFSR_12 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_11_0_0 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_6_NAND2X1_237 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_3_INVX1_374 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_2_OAI22X1_3 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_13_DFFSR_45 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_5_DFFSR_110 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_46_DFFSR_141 INVX1_94/gnd DFFSR_25/S FILL
XFILL_4_OAI21X1_219 BUFX2_35/A DFFSR_97/S FILL
XFILL_36_DFFSR_144 INVX1_8/gnd DFFSR_5/S FILL
XNAND2X1_273 NAND2X1_272/Y INVX1_424/Y BUFX2_16/gnd XOR2X1_10/A DFFSR_65/S NAND2X1
XFILL_26_DFFSR_147 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_48_DFFSR_62 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_2_INVX1_194 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_16_DFFSR_150 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_44_5 INVX1_4/gnd DFFSR_51/S FILL
XFILL_10_DFFSR_92 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_32_DFFSR_12 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_5_OAI21X1_153 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_1_NOR2X1_29 BUFX2_37/A DFFSR_81/S FILL
XFILL_21_DFFSR_52 INVX1_94/gnd DFFSR_52/S FILL
XFILL_4_DFFSR_59 INVX1_4/gnd DFFSR_51/S FILL
XFILL_19_DFFPOSX1_28 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_0_INVX1_411 DFFSR_89/gnd DFFSR_186/S FILL
XNAND3X1_105 INVX1_253/A AOI21X1_33/B AOI21X1_33/A BUFX2_6/gnd NAND3X1_105/Y DFFSR_14/S
+ NAND3X1
XFILL_2_DFFSR_147 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_43_DFFSR_178 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_5_NAND2X1_267 INVX1_4/gnd DFFSR_4/S FILL
XFILL_33_DFFSR_181 INVX1_23/gnd DFFSR_186/S FILL
XFILL_23_DFFSR_184 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_18_DFFSR_99 BUFX2_35/A DFFSR_97/S FILL
XFILL_1_INVX1_53 INVX1_89/gnd DFFSR_2/S FILL
XFILL_40_DFFSR_19 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_29_DFFSR_59 INVX1_4/gnd DFFSR_51/S FILL
XFILL_13_DFFSR_187 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_3_OAI21X1_249 DFFSR_89/gnd DFFSR_186/S FILL
XOAI21X1_123 BUFX2_21/Y INVX1_139/Y OAI21X1_123/C INVX1_23/gnd DFFSR_123/D DFFSR_91/S
+ OAI21X1
XFILL_6_NAND2X1_201 BUFX2_35/A DFFSR_14/S FILL
XFILL_3_INVX1_338 BUFX2_36/A DFFSR_8/S FILL
XFILL_46_DFFSR_105 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_9_DFFSR_181 INVX1_23/gnd DFFSR_186/S FILL
XNAND2X1_237 NOR2X1_18/Y NOR2X1_19/Y BUFX2_8/gnd NAND2X1_68/B DFFSR_10/S NAND2X1
XFILL_36_DFFSR_108 INVX1_89/gnd DFFSR_2/S FILL
XFILL_26_DFFSR_111 INVX1_8/gnd DFFSR_5/S FILL
XFILL_4_OAI21X1_183 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_16_DFFSR_114 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_2_INVX1_158 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_48_DFFSR_26 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_37_DFFSR_66 INVX1_2/gnd DFFSR_51/S FILL
XFILL_5_OAI21X1_117 BUFX2_35/A DFFSR_97/S FILL
XFILL_4_DFFSR_23 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_21_DFFSR_16 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_10_DFFSR_56 INVX1_2/gnd DFFSR_51/S FILL
XFILL_9_OAI22X1_1 BUFX2_36/A DFFSR_8/S FILL
XFILL_0_INVX1_375 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_3_NOR2X1_4 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_2_DFFSR_111 INVX1_8/gnd DFFSR_5/S FILL
XFILL_22_DFFSR_6 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_5_NAND2X1_231 BUFX2_37/A DFFSR_81/S FILL
XFILL_43_DFFSR_142 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_45_DFFSR_73 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_33_DFFSR_145 INVX1_23/gnd DFFSR_186/S FILL
XFILL_23_DFFSR_148 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_4_NAND3X1_129 BUFX2_35/A DFFSR_14/S FILL
XFILL_29_DFFSR_23 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_18_DFFSR_63 INVX1_94/gnd DFFSR_52/S FILL
XFILL_1_INVX1_17 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_1_DFFSR_70 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_44_2_0 INVX1_2/gnd DFFSR_51/S FILL
XFILL_3_OAI21X1_213 BUFX2_36/A DFFSR_6/S FILL
XFILL_6_BUFX2_7 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_13_DFFSR_151 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_6_NAND2X1_165 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_3_INVX1_302 INVX1_8/gnd DFFSR_7/S FILL
XFILL_42_4_1 INVX1_4/gnd DFFSR_4/S FILL
XFILL_9_DFFSR_145 INVX1_23/gnd DFFSR_186/S FILL
XFILL_43_DFFSR_2 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_4_OAI21X1_147 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_20_DFFPOSX1_1 BUFX2_6/gnd DFFSR_14/S FILL
XNAND2X1_201 AND2X2_8/Y AND2X2_9/Y BUFX2_35/A NAND3X1_35/C DFFSR_14/S NAND2X1
XFILL_50_DFFSR_176 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_18_DFFPOSX1_22 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_2_INVX1_122 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_37_DFFSR_30 INVX1_89/gnd DFFSR_36/S FILL
XFILL_9_DFFSR_77 INVX1_89/gnd DFFSR_2/S FILL
XFILL_19_DFFPOSX1_4 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_26_DFFSR_70 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_40_DFFSR_179 INVX1_2/gnd DFFSR_1/S FILL
XFILL_18_DFFPOSX1_7 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_30_DFFSR_182 INVX1_89/gnd DFFSR_36/S FILL
XFILL_20_DFFSR_185 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_10_DFFSR_20 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_4_NAND2X1_261 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_10_DFFSR_188 INVX1_2/gnd DFFSR_1/S FILL
XFILL_0_INVX1_339 BUFX2_36/A DFFSR_8/S FILL
XFILL_4_1 INVX1_23/gnd DFFSR_91/S FILL
XFILL_1_NOR3X1_1 INVX1_94/gnd DFFSR_52/S FILL
XFILL_2_OAI21X1_243 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_5_NAND2X1_195 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_45_DFFSR_37 INVX1_89/gnd DFFSR_2/S FILL
XFILL_43_DFFSR_106 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_33_DFFSR_109 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_6_DFFSR_182 INVX1_89/gnd DFFSR_36/S FILL
XFILL_34_DFFSR_77 INVX1_89/gnd DFFSR_2/S FILL
XFILL_23_DFFSR_112 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_13_DFFSR_115 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_18_DFFSR_27 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_1_DFFSR_34 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_6_NAND2X1_3 INVX1_4/gnd DFFSR_51/S FILL
XFILL_3_INVX1_266 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_3_OAI21X1_177 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_10_OAI22X1_8 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_6_NAND2X1_129 INVX1_4/gnd DFFSR_4/S FILL
XXOR2X1_4 XOR2X1_4/A XOR2X1_4/B DFFSR_89/gnd XOR2X1_4/Y DFFSR_186/S XOR2X1
XFILL_9_DFFSR_109 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_42_DFFSR_84 BUFX2_43/A DFFSR_23/S FILL
XFILL_6_OAI22X1_2 BUFX2_36/A DFFSR_8/S FILL
XNAND2X1_165 BUFX2_4/Y INVX1_243/A BUFX2_8/gnd OAI21X1_165/C DFFSR_25/S NAND2X1
XFILL_50_DFFSR_140 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_4_OAI21X1_111 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_40_DFFSR_143 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_26_2 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_9_DFFSR_41 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_26_DFFSR_34 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_15_DFFSR_74 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_30_DFFSR_146 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_20_DFFSR_149 INVX1_23/gnd DFFSR_91/S FILL
XFILL_4_NAND2X1_225 BUFX2_36/A DFFSR_8/S FILL
XFILL_18_0_0 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_10_DFFSR_152 BUFX2_5/gnd DFFSR_23/S FILL
XINVX1_413 INVX1_413/A DFFSR_89/gnd INVX1_413/Y DFFSR_92/S INVX1
XFILL_50_DFFSR_91 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_5_NOR2X1_28 INVX1_94/gnd DFFSR_52/S FILL
XFILL_0_INVX1_303 INVX1_94/gnd DFFSR_25/S FILL
XFILL_3_NAND3X1_123 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_16_2_1 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_6_DFFSR_146 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_5_NAND2X1_159 BUFX2_43/A DFFSR_97/S FILL
XFILL_2_OAI21X1_207 BUFX2_37/A DFFSR_8/S FILL
XFILL_23_DFFSR_81 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_34_DFFSR_41 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_6_DFFSR_88 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_14_4_2 BUFX2_37/A DFFSR_8/S FILL
XFILL_47_DFFSR_177 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_37_DFFSR_180 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_27_DFFSR_183 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_17_DFFPOSX1_16 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_3_OAI21X1_141 INVX1_94/gnd DFFSR_52/S FILL
XFILL_5_BUFX2_26 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_17_DFFSR_186 INVX1_23/gnd DFFSR_186/S FILL
XFILL_3_INVX1_230 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_34_DFFSR_9 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_8_DFFPOSX1_1 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_3_INVX1_82 BUFX2_35/A DFFSR_97/S FILL
XFILL_42_DFFSR_48 INVX1_4/gnd DFFSR_4/S FILL
XFILL_31_DFFSR_88 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_8_AOI21X1_21 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_7_DFFPOSX1_4 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_50_DFFSR_104 INVX1_4/gnd DFFSR_4/S FILL
XNAND2X1_129 NAND2X1_65/A DFFSR_1/S INVX1_4/gnd OAI21X1_129/C DFFSR_4/S NAND2X1
XFILL_3_NAND2X1_255 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_7_AOI21X1_24 BUFX2_43/A DFFSR_97/S FILL
XFILL_40_DFFSR_107 BUFX2_36/A DFFSR_8/S FILL
XFILL_6_DFFPOSX1_7 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_3_DFFSR_183 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_6_AOI21X1_27 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_15_DFFSR_38 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_30_DFFSR_110 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_20_DFFSR_113 INVX1_23/gnd DFFSR_186/S FILL
XFILL_1_OAI21X1_237 BUFX2_8/gnd DFFSR_10/S FILL
XDFFPOSX1_7 INVX1_243/A CLKBUF1_15/Y DFFPOSX1_7/D DFFSR_71/gnd DFFSR_45/S DFFPOSX1
XFILL_7_DFFPOSX1_27 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_5_AOI21X1_30 INVX1_23/gnd DFFSR_91/S FILL
XAOI21X1_27 INVX1_238/Y AOI21X1_27/B AOI21X1_26/Y BUFX2_5/gnd AOI21X1_27/Y DFFSR_6/S
+ AOI21X1
XFILL_4_NAND2X1_189 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_10_DFFSR_116 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_3_NAND2X1_4 INVX1_2/gnd DFFSR_51/S FILL
XFILL_4_AOI21X1_33 BUFX2_35/A DFFSR_14/S FILL
XFILL_39_DFFSR_95 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_50_DFFSR_55 INVX1_89/gnd DFFSR_36/S FILL
XFILL_0_INVX1_267 BUFX2_17/gnd DFFSR_57/S FILL
XINVX1_377 DFFSR_94/Q DFFSR_73/gnd INVX1_377/Y DFFSR_57/S INVX1
XFILL_3_AOI21X1_36 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_5_NAND2X1_123 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_2_AOI21X1_39 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_0_AND2X2_4 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_2_OAI21X1_171 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_6_DFFSR_52 INVX1_94/gnd DFFSR_52/S FILL
XFILL_4_INVX1_374 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_1_AOI21X1_42 INVX1_23/gnd DFFSR_91/S FILL
XFILL_12_DFFSR_85 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_3_OAI22X1_3 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_23_DFFSR_45 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_6_DFFSR_110 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_47_DFFSR_141 INVX1_94/gnd DFFSR_25/S FILL
XFILL_0_AOI21X1_45 INVX1_89/gnd DFFSR_36/S FILL
XFILL_4_0_2 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_37_DFFSR_144 INVX1_8/gnd DFFSR_5/S FILL
XBUFX2_30 BUFX2_30/A INVX1_4/gnd dout[4] DFFSR_51/S BUFX2
XFILL_27_DFFSR_147 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_3_OAI21X1_105 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_2_NAND2X1_285 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_3_INVX1_194 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_8_OAI21X1_69 BUFX2_37/A DFFSR_8/S FILL
XFILL_17_DFFSR_150 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_48_2 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_7_OAI21X1_72 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_6_NAND2X1_90 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_20_DFFSR_92 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_42_DFFSR_12 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_3_DFFSR_99 BUFX2_35/A DFFSR_97/S FILL
XFILL_2_NOR2X1_29 BUFX2_37/A DFFSR_81/S FILL
XFILL_3_NAND2X1_219 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_31_DFFSR_52 INVX1_94/gnd DFFSR_52/S FILL
XFILL_3_INVX1_46 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_6_OAI21X1_75 INVX1_4/gnd DFFSR_4/S FILL
XFILL_5_NAND2X1_93 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_1_INVX1_411 DFFSR_89/gnd DFFSR_186/S FILL
XNAND2X1_90 BUFX2_18/Y DFFSR_82/Q DFFSR_1/gnd NAND2X1_90/Y DFFSR_1/S NAND2X1
XFILL_5_OAI21X1_78 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_4_NAND2X1_96 INVX1_4/gnd DFFSR_51/S FILL
XFILL_3_DFFSR_147 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_3_NAND2X1_99 BUFX2_43/A DFFSR_97/S FILL
XFILL_4_OAI21X1_81 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_2_NAND3X1_117 INVX1_94/gnd DFFSR_25/S FILL
XOAI21X1_75 BUFX2_18/Y INVX1_85/Y OAI21X1_75/C INVX1_4/gnd DFFSR_75/D DFFSR_4/S OAI21X1
XFILL_3_OAI21X1_84 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_2_BUFX2_37 BUFX2_37/A DFFSR_81/S FILL
XFILL_44_DFFSR_178 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_34_DFFSR_181 INVX1_23/gnd DFFSR_186/S FILL
XFILL_1_OAI21X1_201 BUFX2_35/A DFFSR_97/S FILL
XFILL_4_NAND2X1_153 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_24_DFFSR_184 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_2_OAI21X1_87 INVX1_4/gnd DFFSR_4/S FILL
XFILL_21_DFFSR_3 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_28_DFFSR_99 BUFX2_35/A DFFSR_97/S FILL
XFILL_0_INVX1_231 BUFX2_43/A DFFSR_23/S FILL
XFILL_1_OAI21X1_90 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_50_DFFSR_19 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_0_INVX1_93 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_39_DFFSR_59 INVX1_4/gnd DFFSR_51/S FILL
XINVX1_341 DFFSR_74/Q DFFSR_3/gnd INVX1_341/Y DFFSR_65/S INVX1
XFILL_14_DFFSR_187 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_4_INVX1_338 BUFX2_36/A DFFSR_8/S FILL
XFILL_16_DFFPOSX1_10 INVX1_8/gnd DFFSR_5/S FILL
XFILL_0_OAI21X1_93 INVX1_4/gnd DFFSR_51/S FILL
XFILL_2_OAI21X1_135 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_5_BUFX2_4 BUFX2_8/gnd DFFSR_25/S FILL
XBUFX2_8 rst BUFX2_8/gnd BUFX2_8/Y DFFSR_10/S BUFX2
XFILL_6_DFFSR_16 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_12_DFFSR_49 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_47_DFFSR_105 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_37_DFFSR_108 INVX1_89/gnd DFFSR_2/S FILL
XFILL_27_DFFSR_111 INVX1_8/gnd DFFSR_5/S FILL
XFILL_2_NAND2X1_249 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_0_DFFSR_184 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_17_DFFSR_114 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_3_INVX1_158 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_47_DFFSR_66 INVX1_2/gnd DFFSR_51/S FILL
XFILL_15_5_0 BUFX2_37/A DFFSR_81/S FILL
XFILL_8_OAI21X1_33 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_6_DFFPOSX1_21 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_0_OAI21X1_231 BUFX2_36/A DFFSR_6/S FILL
XFILL_3_INVX1_10 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_6_NAND2X1_54 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_3_DFFSR_63 INVX1_94/gnd DFFSR_52/S FILL
XFILL_31_DFFSR_16 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_7_OAI21X1_36 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_0_NAND2X1_5 INVX1_8/gnd DFFSR_7/S FILL
XFILL_20_DFFSR_56 INVX1_2/gnd DFFSR_51/S FILL
XNAND2X1_54 DFFSR_8/S DFFSR_46/Q BUFX2_7/gnd OAI21X1_54/C DFFSR_54/S NAND2X1
XFILL_6_OAI21X1_39 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_3_NAND2X1_183 INVX1_8/gnd DFFSR_7/S FILL
XFILL_5_NAND2X1_57 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_4_NAND2X1_60 BUFX2_7/gnd DFFSR_54/S FILL
XOAI21X1_39 DFFSR_36/S INVX1_44/Y NAND2X1_39/Y DFFSR_71/gnd DFFSR_39/D DFFSR_45/S
+ OAI21X1
XFILL_5_OAI21X1_42 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_1_INVX1_375 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_0_OAI22X1_4 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_3_NAND2X1_63 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_4_OAI21X1_45 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_3_DFFSR_111 INVX1_8/gnd DFFSR_5/S FILL
XFILL_1_OAI21X1_165 BUFX2_35/A DFFSR_97/S FILL
XFILL_44_DFFSR_142 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_2_NAND2X1_66 INVX1_4/gnd DFFSR_51/S FILL
XFILL_3_OAI21X1_48 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_34_DFFSR_145 INVX1_23/gnd DFFSR_186/S FILL
XFILL_4_NAND2X1_117 BUFX2_35/A DFFSR_14/S FILL
XFILL_1_NAND2X1_69 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_2_OAI21X1_51 INVX1_2/gnd DFFSR_51/S FILL
XFILL_24_DFFSR_148 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_0_INVX1_195 INVX1_23/gnd DFFSR_186/S FILL
XFILL_39_DFFSR_23 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_1_OAI21X1_54 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_28_DFFSR_63 INVX1_94/gnd DFFSR_52/S FILL
XINVX1_305 INVX1_25/A BUFX2_8/gnd INVX1_305/Y DFFSR_25/S INVX1
XFILL_0_NAND2X1_72 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_0_INVX1_57 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_14_DFFSR_151 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_0_OAI21X1_57 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_1_NAND2X1_279 INVX1_89/gnd DFFSR_2/S FILL
XFILL_4_INVX1_302 INVX1_8/gnd DFFSR_7/S FILL
XFILL_25_DFFPOSX1_29 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_12_DFFSR_13 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_0_DFFSR_148 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_2_NAND2X1_213 BUFX2_35/A DFFSR_97/S FILL
XNOR2X1_1 NOR2X1_1/A NOR2X1_1/B BUFX2_36/A AND2X2_1/A DFFSR_6/S NOR2X1
XFILL_51_DFFSR_176 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_3_INVX1_122 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_25_0_0 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_47_DFFSR_30 INVX1_89/gnd DFFSR_36/S FILL
XFILL_41_DFFSR_179 INVX1_2/gnd DFFSR_1/S FILL
XFILL_1_NAND3X1_111 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_31_DFFSR_182 INVX1_89/gnd DFFSR_36/S FILL
XFILL_36_DFFSR_70 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_21_DFFSR_185 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_23_2_1 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_6_NAND2X1_18 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_20_DFFSR_20 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_3_NAND2X1_147 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_5_1_0 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_0_OAI21X1_195 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_9_OAI21X1_250 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_3_DFFSR_27 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_11_DFFSR_188 INVX1_2/gnd DFFSR_1/S FILL
XFILL_5_NAND2X1_21 INVX1_4/gnd DFFSR_4/S FILL
XFILL_1_INVX1_339 BUFX2_36/A DFFSR_8/S FILL
XFILL_21_4_2 INVX1_94/gnd DFFSR_25/S FILL
XFILL_4_NAND2X1_24 DFFSR_73/gnd DFFSR_57/S FILL
XNAND2X1_18 DFFSR_9/S DFFSR_10/Q DFFSR_1/gnd NAND2X1_18/Y DFFSR_9/S NAND2X1
XFILL_3_3_1 INVX1_23/gnd DFFSR_91/S FILL
XFILL_2_NOR2X1_8 BUFX2_43/A DFFSR_23/S FILL
XFILL_9_DFFSR_2 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_3_NAND2X1_27 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_11_OAI22X1_65 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_3_OAI21X1_12 BUFX2_35/A DFFSR_14/S FILL
XDFFPOSX1_21 AND2X2_11/A CLKBUF1_11/Y XOR2X1_17/Y BUFX2_5/gnd DFFSR_23/S DFFPOSX1
XFILL_2_NAND2X1_30 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_10_OAI22X1_68 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_44_DFFSR_106 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_34_DFFSR_109 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_1_NAND2X1_33 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_7_DFFSR_182 INVX1_89/gnd DFFSR_36/S FILL
XFILL_44_DFFSR_77 INVX1_89/gnd DFFSR_2/S FILL
XFILL_1_OAI21X1_129 INVX1_4/gnd DFFSR_4/S FILL
XFILL_1_5_2 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_8_NAND3X1_89 BUFX2_43/A DFFSR_23/S FILL
XFILL_2_OAI21X1_15 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_24_DFFSR_112 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_14_DFFSR_115 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_7_NAND3X1_92 BUFX2_43/A DFFSR_23/S FILL
XFILL_0_INVX1_159 INVX1_94/gnd DFFSR_52/S FILL
XFILL_0_NAND2X1_36 DFFSR_71/gnd DFFSR_45/S FILL
XINVX1_269 DFFSR_33/Q DFFSR_5/gnd INVX1_269/Y DFFSR_5/S INVX1
XFILL_28_DFFSR_27 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_0_INVX1_21 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_0_DFFSR_74 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_1_OAI21X1_18 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_17_DFFSR_67 INVX1_2/gnd DFFSR_51/S FILL
XFILL_6_NAND3X1_95 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_4_INVX1_266 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_11_OAI22X1_8 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_0_OAI21X1_21 INVX1_2/gnd DFFSR_51/S FILL
XFILL_1_NAND2X1_243 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_7_OR2X2_2 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_4_XOR2X1_4 DFFSR_89/gnd DFFSR_186/S FILL
XNAND3X1_95 NAND3X1_95/A NAND3X1_95/B OR2X2_2/Y BUFX2_6/gnd AOI21X1_30/A DFFSR_91/S
+ NAND3X1
XFILL_5_NAND3X1_98 BUFX2_35/A DFFSR_14/S FILL
XFILL_33_DFFSR_6 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_7_OAI22X1_2 BUFX2_36/A DFFSR_8/S FILL
XFILL_5_DFFPOSX1_15 BUFX2_35/A DFFSR_14/S FILL
XFILL_2_NAND2X1_177 INVX1_89/gnd DFFSR_36/S FILL
XFILL_0_DFFSR_112 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_8_DFFSR_81 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_41_DFFSR_143 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_36_DFFSR_34 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_25_DFFSR_74 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_31_DFFSR_146 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_21_DFFSR_149 INVX1_23/gnd DFFSR_91/S FILL
XFILL_0_OAI21X1_159 BUFX2_43/A DFFSR_97/S FILL
XFILL_9_OAI21X1_214 BUFX2_35/A DFFSR_97/S FILL
XFILL_11_DFFSR_152 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_3_NAND2X1_111 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_6_NOR2X1_28 INVX1_94/gnd DFFSR_52/S FILL
XFILL_1_INVX1_303 INVX1_94/gnd DFFSR_25/S FILL
XFILL_1_AOI22X1_11 INVX1_23/gnd DFFSR_91/S FILL
XFILL_7_DFFSR_146 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_33_DFFSR_81 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_10_OAI22X1_32 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_0_AOI22X1_14 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_44_DFFSR_41 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_0_NAND2X1_273 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_24_DFFPOSX1_23 INVX1_23/gnd DFFSR_91/S FILL
XFILL_48_DFFSR_177 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_17_DFFSR_31 BUFX2_35/A DFFSR_97/S FILL
XFILL_0_INVX1_123 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_8_NAND3X1_53 BUFX2_37/A DFFSR_81/S FILL
XINVX1_233 INVX1_233/A BUFX2_7/gnd INVX1_233/Y DFFSR_54/S INVX1
XFILL_38_DFFSR_180 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_9_OAI22X1_35 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_0_DFFSR_38 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_28_DFFSR_183 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_7_NAND3X1_56 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_8_OAI22X1_38 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_18_DFFSR_186 INVX1_23/gnd DFFSR_186/S FILL
XFILL_1_NAND2X1_207 BUFX2_43/A DFFSR_97/S FILL
XFILL_6_NAND3X1_59 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_7_OAI22X1_41 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_0_NAND3X1_105 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_5_NAND3X1_62 BUFX2_43/A DFFSR_23/S FILL
XFILL_6_OAI22X1_44 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_4_NAND3X1_65 BUFX2_35/A DFFSR_14/S FILL
XFILL_5_OAI22X1_47 BUFX2_37/A DFFSR_8/S FILL
XNAND3X1_59 INVX1_243/A NAND3X1_55/Y NAND3X1_58/Y BUFX2_8/gnd INVX1_244/A DFFSR_25/S
+ NAND3X1
XFILL_10_XOR2X1_1 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_41_DFFSR_88 DFFSR_3/gnd DFFSR_4/S FILL
XDFFSR_186 BUFX2_28/A DFFSR_20/CLK DFFSR_185/R DFFSR_186/S DFFSR_186/D INVX1_23/gnd
+ DFFSR_186/S DFFSR
XFILL_3_NAND3X1_68 BUFX2_35/A DFFSR_14/S FILL
XFILL_2_NAND2X1_141 INVX1_94/gnd DFFSR_25/S FILL
XFILL_4_OAI22X1_50 DFFSR_79/gnd DFFSR_36/S FILL
XOAI22X1_44 INVX1_347/Y OAI22X1_39/B INVX1_346/Y OAI22X1_39/D BUFX2_16/gnd NOR2X1_31/B
+ DFFSR_11/S OAI22X1
XFILL_2_NAND3X1_71 BUFX2_35/A DFFSR_14/S FILL
XFILL_41_DFFSR_107 BUFX2_36/A DFFSR_8/S FILL
XFILL_3_OAI22X1_53 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_8_DFFSR_45 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_8_OAI21X1_244 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_4_DFFSR_183 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_1_NAND3X1_74 BUFX2_35/A DFFSR_14/S FILL
XFILL_2_OAI22X1_56 BUFX2_37/A DFFSR_8/S FILL
XFILL_25_DFFSR_38 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_14_DFFSR_78 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_31_DFFSR_110 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_21_DFFSR_113 INVX1_23/gnd DFFSR_186/S FILL
XFILL_0_NAND3X1_77 BUFX2_37/A DFFSR_81/S FILL
XNAND2X1_7 DFFSR_36/S INVX1_412/A INVX1_89/gnd NAND2X1_7/Y DFFSR_36/S NAND2X1
XFILL_1_OAI22X1_59 INVX1_8/gnd DFFSR_7/S FILL
XFILL_0_OAI21X1_123 INVX1_23/gnd DFFSR_91/S FILL
XFILL_0_OAI22X1_62 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_11_DFFSR_116 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_49_DFFSR_95 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_1_INVX1_267 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_0_DFFSR_9 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_4_NAND2X1_4 INVX1_2/gnd DFFSR_51/S FILL
XFILL_0_NAND2X1_237 BUFX2_8/gnd DFFSR_10/S FILL
XOAI22X1_6 INVX1_267/Y OAI22X1_6/B INVX1_268/Y OAI22X1_6/D DFFSR_73/gnd OAI22X1_6/Y
+ DFFSR_11/S OAI22X1
XINVX1_79 DFFSR_70/Q DFFSR_73/gnd INVX1_79/Y DFFSR_57/S INVX1
XFILL_5_DFFSR_92 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_9_NAND3X1_14 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_22_DFFSR_85 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_4_OAI22X1_3 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_33_DFFSR_45 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_7_DFFSR_110 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_48_DFFSR_141 INVX1_94/gnd DFFSR_25/S FILL
XFILL_22_5_0 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_8_NAND3X1_17 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_4_BUFX2_1 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_7_NAND3X1_20 BUFX2_37/A DFFSR_8/S FILL
XFILL_38_DFFSR_144 INVX1_8/gnd DFFSR_5/S FILL
XFILL_4_BUFX2_30 INVX1_4/gnd DFFSR_51/S FILL
XINVX1_197 DFFSR_163/Q DFFSR_3/gnd INVX1_197/Y DFFSR_4/S INVX1
XFILL_28_DFFSR_147 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_6_NAND3X1_23 BUFX2_37/A DFFSR_81/S FILL
XFILL_1_NAND2X1_171 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_35_4 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_4_INVX1_194 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_18_DFFSR_150 BUFX2_8/gnd DFFSR_25/S FILL
XNAND3X1_23 AOI21X1_5/C AOI21X1_5/A AOI21X1_5/B BUFX2_37/A NAND3X1_23/Y DFFSR_81/S
+ NAND3X1
XFILL_5_NAND3X1_26 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_30_DFFSR_92 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_3_NOR2X1_29 BUFX2_37/A DFFSR_81/S FILL
XFILL_4_NAND3X1_29 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_2_INVX1_86 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_41_DFFSR_52 INVX1_94/gnd DFFSR_52/S FILL
XFILL_9_NAND3X1_124 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_5_OAI22X1_11 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_13_DFFPOSX1_28 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_2_INVX1_411 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_2_NAND2X1_105 BUFX2_35/A DFFSR_14/S FILL
XFILL_8_OAI21X1_208 BUFX2_5/gnd DFFSR_6/S FILL
XDFFSR_150 INVX1_174/A CLKBUF1_9/Y INVX1_175/Y DFFSR_25/S DFFSR_150/D BUFX2_8/gnd
+ DFFSR_25/S DFFSR
XFILL_3_NAND3X1_32 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_4_OAI22X1_14 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_4_DFFSR_147 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_2_NAND3X1_35 BUFX2_35/A DFFSR_97/S FILL
XFILL_3_OAI22X1_17 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_14_DFFSR_42 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_1_NAND3X1_38 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_2_OAI22X1_20 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_45_DFFSR_178 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_35_DFFSR_181 INVX1_23/gnd DFFSR_186/S FILL
XFILL_0_NAND3X1_41 BUFX2_43/A DFFSR_23/S FILL
XFILL_1_OAI22X1_23 INVX1_89/gnd DFFSR_2/S FILL
XFILL_23_DFFPOSX1_17 BUFX2_37/A DFFSR_8/S FILL
XFILL_0_OAI22X1_26 INVX1_94/gnd DFFSR_52/S FILL
XFILL_25_DFFSR_184 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_45_DFFSR_9 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_38_DFFSR_99 BUFX2_35/A DFFSR_97/S FILL
XFILL_1_INVX1_231 BUFX2_43/A DFFSR_23/S FILL
XFILL_49_DFFSR_59 INVX1_4/gnd DFFSR_51/S FILL
XFILL_15_DFFSR_187 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_11_DFFSR_89 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_0_NAND2X1_201 BUFX2_35/A DFFSR_14/S FILL
XINVX1_43 INVX1_43/A DFFSR_5/gnd INVX1_43/Y DFFSR_5/S INVX1
XFILL_32_0_0 INVX1_8/gnd DFFSR_5/S FILL
XDFFSR_96 DFFSR_96/Q CLKBUF1_5/Y DFFSR_89/R DFFSR_1/S DFFSR_96/D INVX1_2/gnd DFFSR_1/S
+ DFFSR
XFILL_5_DFFSR_56 INVX1_2/gnd DFFSR_51/S FILL
XFILL_22_DFFSR_49 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_48_DFFSR_105 DFFSR_89/gnd DFFSR_186/S FILL
XINVX1_161 DFFSR_143/Q BUFX2_8/gnd INVX1_161/Y DFFSR_10/S INVX1
XFILL_38_DFFSR_108 INVX1_89/gnd DFFSR_2/S FILL
XFILL_30_2_1 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_28_DFFSR_111 INVX1_8/gnd DFFSR_5/S FILL
XFILL_1_DFFSR_184 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_1_NAND2X1_135 BUFX2_36/A DFFSR_6/S FILL
XFILL_7_OAI21X1_238 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_18_DFFSR_114 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_4_INVX1_158 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_28_4_2 INVX1_89/gnd DFFSR_36/S FILL
XFILL_2_INVX1_50 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_41_DFFSR_16 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_1_NAND2X1_5 INVX1_8/gnd DFFSR_7/S FILL
XFILL_19_DFFSR_96 INVX1_2/gnd DFFSR_1/S FILL
XFILL_30_DFFSR_56 INVX1_2/gnd DFFSR_51/S FILL
XDFFSR_114 INVX1_344/A CLKBUF1_1/Y DFFSR_113/R DFFSR_45/S DFFSR_114/D DFFSR_71/gnd
+ DFFSR_45/S DFFSR
XFILL_8_5_2 BUFX2_43/A DFFSR_97/S FILL
XFILL_8_OAI21X1_172 BUFX2_36/A DFFSR_6/S FILL
XFILL_2_INVX1_375 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_1_BUFX2_41 BUFX2_37/A DFFSR_81/S FILL
XFILL_1_OAI22X1_4 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_4_DFFSR_111 INVX1_8/gnd DFFSR_5/S FILL
XFILL_45_DFFSR_142 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_35_DFFSR_145 INVX1_23/gnd DFFSR_186/S FILL
XFILL_11_DFFSR_7 INVX1_8/gnd DFFSR_7/S FILL
XFILL_25_DFFSR_148 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_1_INVX1_195 INVX1_23/gnd DFFSR_186/S FILL
XFILL_49_DFFSR_23 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_38_DFFSR_63 INVX1_94/gnd DFFSR_52/S FILL
XFILL_15_DFFSR_151 BUFX2_7/gnd DFFSR_81/S FILL
XDFFSR_60 DFFSR_60/Q INVX1_1/A DFFSR_61/R DFFSR_8/S DFFSR_60/D BUFX2_37/A DFFSR_8/S
+ DFFSR
XFILL_0_NAND2X1_165 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_5_DFFSR_20 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_11_DFFSR_53 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_22_DFFSR_13 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_0_NOR2X1_30 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_1_DFFSR_148 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_4_NOR2X1_1 BUFX2_36/A DFFSR_6/S FILL
XFILL_8_NAND3X1_118 DFFSR_79/gnd DFFSR_45/S FILL
XINVX1_125 INVX1_387/A DFFSR_5/gnd INVX1_125/Y DFFSR_5/S INVX1
XFILL_12_DFFPOSX1_22 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_7_OAI21X1_202 BUFX2_35/A DFFSR_14/S FILL
XFILL_4_INVX1_122 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_42_DFFSR_179 INVX1_2/gnd DFFSR_1/S FILL
XFILL_32_DFFSR_3 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_32_DFFSR_182 INVX1_89/gnd DFFSR_36/S FILL
XFILL_46_DFFSR_70 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_22_DFFSR_185 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_30_DFFSR_20 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_2_INVX1_14 BUFX2_35/A DFFSR_14/S FILL
XFILL_19_DFFSR_60 BUFX2_37/A DFFSR_8/S FILL
XFILL_12_DFFSR_188 INVX1_2/gnd DFFSR_1/S FILL
XFILL_2_DFFSR_67 INVX1_2/gnd DFFSR_51/S FILL
XFILL_2_INVX1_339 BUFX2_36/A DFFSR_8/S FILL
XFILL_8_OAI21X1_136 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_22_DFFPOSX1_11 INVX1_4/gnd DFFSR_4/S FILL
XFILL_45_DFFSR_106 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_35_DFFSR_109 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_8_DFFSR_182 INVX1_89/gnd DFFSR_36/S FILL
XFILL_25_DFFSR_112 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_15_DFFSR_115 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_1_INVX1_159 INVX1_94/gnd DFFSR_52/S FILL
XFILL_38_DFFSR_27 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_27_DFFSR_67 INVX1_2/gnd DFFSR_51/S FILL
XFILL_6_OAI21X1_232 BUFX2_35/A DFFSR_97/S FILL
XFILL_11_DFFSR_17 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_0_NAND2X1_129 INVX1_4/gnd DFFSR_4/S FILL
XDFFSR_24 INVX1_27/A DFFSR_24/CLK DFFSR_20/R DFFSR_65/S DFFSR_24/D BUFX2_16/gnd DFFSR_65/S
+ DFFSR
XFILL_8_OAI22X1_2 BUFX2_36/A DFFSR_8/S FILL
XFILL_17_1 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_1_DFFSR_112 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_42_DFFSR_143 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_46_DFFSR_34 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_35_DFFSR_74 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_7_OAI21X1_166 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_32_DFFSR_146 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_22_DFFSR_149 INVX1_23/gnd DFFSR_91/S FILL
XFILL_2_DFFSR_31 BUFX2_35/A DFFSR_97/S FILL
XFILL_19_DFFSR_24 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_12_DFFSR_152 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_8_OAI21X1_100 INVX1_23/gnd DFFSR_91/S FILL
XFILL_2_INVX1_303 INVX1_94/gnd DFFSR_25/S FILL
XFILL_29_5_0 INVX1_89/gnd DFFSR_2/S FILL
XFILL_8_DFFSR_146 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_43_DFFSR_81 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_19_CLKBUF1_17 INVX1_94/gnd DFFSR_25/S FILL
XFILL_5_OAI21X1_262 INVX1_89/gnd DFFSR_36/S FILL
XFILL_49_DFFSR_177 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_18_CLKBUF1_20 INVX1_4/gnd DFFSR_51/S FILL
XFILL_1_INVX1_123 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_17_CLKBUF1_23 INVX1_89/gnd DFFSR_2/S FILL
XFILL_39_DFFSR_180 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_29_DFFSR_183 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_27_DFFSR_31 BUFX2_35/A DFFSR_97/S FILL
XFILL_7_NAND3X1_112 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_16_DFFSR_71 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_19_DFFSR_186 INVX1_23/gnd DFFSR_186/S FILL
XFILL_11_DFFPOSX1_16 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_6_OAI21X1_196 INVX1_94/gnd DFFSR_25/S FILL
XFILL_3_XOR2X1_8 BUFX2_5/gnd DFFSR_6/S FILL
XOAI21X1_232 INVX1_248/A INVX1_249/A NAND3X1_66/C BUFX2_35/A INVX1_258/A DFFSR_97/S
+ OAI21X1
XFILL_42_DFFSR_107 BUFX2_36/A DFFSR_8/S FILL
XFILL_7_OAI21X1_130 INVX1_4/gnd DFFSR_4/S FILL
XFILL_5_DFFSR_183 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_7_DFFSR_85 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_35_DFFSR_38 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_24_DFFSR_78 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_32_DFFSR_110 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_22_DFFSR_113 INVX1_23/gnd DFFSR_186/S FILL
XFILL_6_BUFX2_23 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_1_DFFPOSX1_27 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_12_DFFSR_116 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_39_0_0 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_2_INVX1_267 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_5_NAND2X1_4 INVX1_2/gnd DFFSR_51/S FILL
XFILL_44_DFFSR_6 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_16_NOR3X1_2 INVX1_89/gnd DFFSR_2/S FILL
XFILL_37_2_1 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_5_OAI21X1_226 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_32_DFFSR_85 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_5_OAI22X1_3 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_43_DFFSR_45 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_4_INVX1_79 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_8_DFFSR_110 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_49_DFFSR_141 INVX1_94/gnd DFFSR_25/S FILL
XFILL_35_4_2 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_22_6 INVX1_94/gnd DFFSR_25/S FILL
XFILL_16_DFFSR_35 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_39_DFFSR_144 INVX1_8/gnd DFFSR_5/S FILL
XFILL_29_DFFSR_147 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_39_1 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_19_DFFSR_150 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_6_OAI21X1_160 DFFSR_73/gnd DFFSR_57/S FILL
XNOR2X1_32 NOR2X1_32/A NOR2X1_32/B INVX1_94/gnd NOR2X1_32/Y DFFSR_52/S NOR2X1
XFILL_40_DFFSR_92 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_4_NOR2X1_29 BUFX2_37/A DFFSR_81/S FILL
XOAI21X1_196 NOR3X1_1/B NOR3X1_1/C NOR3X1_1/A INVX1_94/gnd AOI21X1_13/B DFFSR_25/S
+ OAI21X1
XFILL_6_NAND2X1_274 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_5_DFFSR_147 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_3_INVX1_411 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_1_AND2X2_1 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_13_DFFSR_82 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_24_DFFSR_42 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_7_DFFSR_49 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_46_DFFSR_178 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_36_DFFSR_181 INVX1_23/gnd DFFSR_186/S FILL
XFILL_9_CLKBUF1_11 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_26_DFFSR_184 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_4_OAI21X1_256 INVX1_2/gnd DFFSR_51/S FILL
XFILL_48_DFFSR_99 BUFX2_35/A DFFSR_97/S FILL
XFILL_2_INVX1_231 BUFX2_43/A DFFSR_23/S FILL
XFILL_10_DFFSR_4 INVX1_4/gnd DFFSR_4/S FILL
XFILL_16_DFFSR_187 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_8_CLKBUF1_14 BUFX2_43/A DFFSR_23/S FILL
XFILL_6_NAND3X1_106 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_21_DFFSR_89 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_9_AND2X2_8 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_7_CLKBUF1_17 INVX1_94/gnd DFFSR_25/S FILL
XFILL_10_DFFPOSX1_10 INVX1_8/gnd DFFSR_5/S FILL
XFILL_4_DFFSR_96 INVX1_2/gnd DFFSR_1/S FILL
XFILL_32_DFFSR_49 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_49_DFFSR_105 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_5_OAI21X1_190 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_6_CLKBUF1_20 INVX1_4/gnd DFFSR_51/S FILL
XFILL_5_CLKBUF1_23 INVX1_89/gnd DFFSR_2/S FILL
XFILL_39_DFFSR_108 INVX1_89/gnd DFFSR_2/S FILL
XCLKBUF1_20 INVX1_402/Y INVX1_4/gnd DFFSR_24/CLK DFFSR_51/S CLKBUF1
XFILL_3_BUFX2_34 BUFX2_37/A DFFSR_81/S FILL
XFILL_29_DFFSR_111 INVX1_8/gnd DFFSR_5/S FILL
XFILL_2_DFFSR_184 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_19_DFFSR_114 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_6_OAI21X1_124 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_2_NAND2X1_5 INVX1_8/gnd DFFSR_7/S FILL
XFILL_29_DFFSR_96 INVX1_2/gnd DFFSR_1/S FILL
XFILL_40_DFFSR_56 INVX1_2/gnd DFFSR_51/S FILL
XFILL_1_INVX1_90 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_0_DFFPOSX1_21 BUFX2_5/gnd DFFSR_23/S FILL
XOAI21X1_160 BUFX2_1/Y INVX1_194/Y NAND2X1_160/Y DFFSR_73/gnd DFFSR_160/D DFFSR_57/S
+ OAI21X1
XFILL_11_0_1 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_6_NAND2X1_238 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_3_INVX1_375 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_13_DFFSR_46 BUFX2_36/A DFFSR_6/S FILL
XFILL_2_OAI22X1_4 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_5_DFFSR_111 INVX1_8/gnd DFFSR_5/S FILL
XFILL_7_DFFSR_13 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_46_DFFSR_142 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_36_DFFSR_145 INVX1_23/gnd DFFSR_186/S FILL
XFILL_4_OAI21X1_220 BUFX2_43/A DFFSR_97/S FILL
XNAND2X1_274 NOR2X1_47/A INVX1_426/Y BUFX2_17/gnd AOI21X1_44/B DFFSR_57/S NAND2X1
XFILL_26_DFFSR_148 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_2_INVX1_195 INVX1_23/gnd DFFSR_186/S FILL
XFILL_48_DFFSR_63 INVX1_94/gnd DFFSR_52/S FILL
XFILL_16_DFFSR_151 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_4_DFFSR_60 BUFX2_37/A DFFSR_8/S FILL
XFILL_5_OAI21X1_154 BUFX2_37/A DFFSR_8/S FILL
XFILL_21_DFFSR_53 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_19_DFFPOSX1_29 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_10_DFFSR_93 INVX1_2/gnd DFFSR_51/S FILL
XFILL_32_DFFSR_13 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_1_NOR2X1_30 DFFSR_73/gnd DFFSR_57/S FILL
XNAND3X1_106 XOR2X1_8/B AOI21X1_32/B AOI21X1_32/A BUFX2_5/gnd NAND3X1_107/C DFFSR_6/S
+ NAND3X1
XFILL_2_DFFSR_148 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_0_INVX1_412 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_43_DFFSR_179 INVX1_2/gnd DFFSR_1/S FILL
XFILL_5_NAND2X1_268 BUFX2_37/A DFFSR_8/S FILL
XFILL_33_DFFSR_182 INVX1_89/gnd DFFSR_36/S FILL
XFILL_36_5_0 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_23_DFFSR_185 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_40_DFFSR_20 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_29_DFFSR_60 BUFX2_37/A DFFSR_8/S FILL
XFILL_13_DFFSR_188 INVX1_2/gnd DFFSR_1/S FILL
XFILL_1_INVX1_54 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_6_NAND2X1_202 BUFX2_35/A DFFSR_97/S FILL
XFILL_3_OAI21X1_250 DFFSR_79/gnd DFFSR_36/S FILL
XOAI21X1_124 BUFX2_23/Y INVX1_140/Y NAND2X1_124/Y DFFSR_79/gnd DFFSR_124/D DFFSR_36/S
+ OAI21X1
XFILL_3_INVX1_339 BUFX2_36/A DFFSR_8/S FILL
XFILL_13_DFFSR_10 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_5_NAND3X1_100 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_46_DFFSR_106 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_36_DFFSR_109 BUFX2_6/gnd DFFSR_14/S FILL
XNAND2X1_238 NOR2X1_21/Y NOR2X1_20/Y DFFSR_79/gnd NAND2X1_69/B DFFSR_36/S NAND2X1
XFILL_9_DFFSR_182 INVX1_89/gnd DFFSR_36/S FILL
XFILL_4_OAI21X1_184 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_26_DFFSR_112 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_16_DFFSR_115 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_2_INVX1_159 INVX1_94/gnd DFFSR_52/S FILL
XFILL_48_DFFSR_27 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_37_DFFSR_67 INVX1_2/gnd DFFSR_51/S FILL
XFILL_21_DFFSR_17 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_10_DFFSR_57 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_4_DFFSR_24 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_5_OAI21X1_118 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_9_OAI22X1_2 BUFX2_36/A DFFSR_8/S FILL
XFILL_0_INVX1_376 INVX1_8/gnd DFFSR_7/S FILL
XFILL_3_NOR2X1_5 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_46_0_0 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_2_DFFSR_112 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_5_NAND2X1_232 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_43_DFFSR_143 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_22_DFFSR_7 INVX1_8/gnd DFFSR_7/S FILL
XFILL_45_DFFSR_74 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_33_DFFSR_146 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_23_DFFSR_149 INVX1_23/gnd DFFSR_91/S FILL
XFILL_4_NAND3X1_130 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_1_DFFSR_71 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_1_INVX1_18 INVX1_89/gnd DFFSR_2/S FILL
XFILL_44_2_1 INVX1_2/gnd DFFSR_51/S FILL
XFILL_29_DFFSR_24 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_13_DFFSR_152 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_6_BUFX2_8 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_18_DFFSR_64 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_3_OAI21X1_214 BUFX2_35/A DFFSR_97/S FILL
XFILL_3_INVX1_303 INVX1_94/gnd DFFSR_25/S FILL
XFILL_42_4_2 INVX1_4/gnd DFFSR_4/S FILL
XFILL_6_NAND2X1_166 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_9_DFFSR_146 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_5_XOR2X1_1 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_43_DFFSR_3 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_4_OAI21X1_148 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_18_DFFPOSX1_23 INVX1_23/gnd DFFSR_91/S FILL
XNAND2X1_202 INVX1_256/A AND2X2_5/B BUFX2_35/A INVX1_241/A DFFSR_97/S NAND2X1
XFILL_20_DFFPOSX1_2 INVX1_89/gnd DFFSR_36/S FILL
XFILL_50_DFFSR_177 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_2_INVX1_123 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_40_DFFSR_180 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_9_DFFSR_78 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_19_DFFPOSX1_5 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_30_DFFSR_183 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_37_DFFSR_31 BUFX2_35/A DFFSR_97/S FILL
XFILL_26_DFFSR_71 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_18_DFFPOSX1_8 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_20_DFFSR_186 INVX1_23/gnd DFFSR_186/S FILL
XFILL_10_3_0 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_4_NAND2X1_262 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_10_DFFSR_189 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_10_DFFSR_21 INVX1_2/gnd DFFSR_1/S FILL
XFILL_4_2 INVX1_23/gnd DFFSR_91/S FILL
XFILL_1_NOR3X1_2 INVX1_89/gnd DFFSR_2/S FILL
XFILL_0_INVX1_340 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_43_DFFSR_107 BUFX2_36/A DFFSR_8/S FILL
XFILL_2_OAI21X1_244 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_6_DFFSR_183 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_5_NAND2X1_196 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_45_DFFSR_38 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_34_DFFSR_78 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_33_DFFSR_110 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_23_DFFSR_113 INVX1_23/gnd DFFSR_186/S FILL
XFILL_18_DFFSR_28 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_1_DFFSR_35 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_13_DFFSR_116 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_3_OAI21X1_178 INVX1_94/gnd DFFSR_25/S FILL
XFILL_10_OAI22X1_9 INVX1_8/gnd DFFSR_5/S FILL
XFILL_3_INVX1_267 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_6_NAND2X1_4 INVX1_2/gnd DFFSR_51/S FILL
XFILL_6_NAND2X1_130 INVX1_4/gnd DFFSR_4/S FILL
XXOR2X1_5 XOR2X1_5/A XOR2X1_5/B DFFSR_89/gnd XOR2X1_5/Y DFFSR_186/S XOR2X1
XFILL_42_DFFSR_85 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_6_OAI22X1_3 DFFSR_79/gnd DFFSR_45/S FILL
XNAND2X1_166 BUFX2_1/Y INVX1_250/A DFFSR_3/gnd NAND2X1_166/Y DFFSR_65/S NAND2X1
XFILL_9_DFFSR_110 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_50_DFFSR_141 INVX1_94/gnd DFFSR_25/S FILL
XFILL_4_OAI21X1_112 INVX1_4/gnd DFFSR_4/S FILL
XFILL_26_3 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_26_DFFSR_35 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_40_DFFSR_144 INVX1_8/gnd DFFSR_5/S FILL
XFILL_15_DFFSR_75 INVX1_4/gnd DFFSR_51/S FILL
XFILL_9_DFFSR_42 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_30_DFFSR_147 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_4_NAND2X1_226 BUFX2_36/A DFFSR_6/S FILL
XFILL_18_0_1 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_20_DFFSR_150 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_10_DFFSR_153 BUFX2_36/A DFFSR_8/S FILL
XFILL_50_DFFSR_92 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_5_NOR2X1_29 BUFX2_37/A DFFSR_81/S FILL
XFILL_0_INVX1_304 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_3_NAND3X1_124 DFFSR_5/gnd DFFSR_5/S FILL
XINVX1_414 BUFX2_8/Y INVX1_2/gnd DFFSR_183/R DFFSR_1/S INVX1
XFILL_16_2_2 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_6_DFFSR_89 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_6_DFFSR_147 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_2_OAI21X1_208 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_5_NAND2X1_160 INVX1_8/gnd DFFSR_5/S FILL
XFILL_23_DFFSR_82 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_34_DFFSR_42 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_47_DFFSR_178 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_37_DFFSR_181 INVX1_23/gnd DFFSR_186/S FILL
XFILL_5_BUFX2_27 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_17_DFFPOSX1_17 BUFX2_37/A DFFSR_8/S FILL
XFILL_3_OAI21X1_142 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_27_DFFSR_184 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_3_INVX1_231 BUFX2_43/A DFFSR_23/S FILL
XFILL_17_DFFSR_187 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_31_DFFSR_89 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_9_AOI21X1_19 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_8_DFFPOSX1_2 INVX1_89/gnd DFFSR_36/S FILL
XFILL_3_INVX1_83 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_42_DFFSR_49 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_50_DFFSR_105 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_8_AOI21X1_22 BUFX2_43/A DFFSR_97/S FILL
XFILL_3_NAND2X1_256 DFFSR_5/gnd DFFSR_2/S FILL
XNAND2X1_130 DFFSR_4/S NAND2X1_66/B INVX1_4/gnd OAI21X1_130/C DFFSR_4/S NAND2X1
XFILL_7_DFFPOSX1_5 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_6_DFFPOSX1_8 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_40_DFFSR_108 INVX1_89/gnd DFFSR_2/S FILL
XFILL_43_5_0 INVX1_4/gnd DFFSR_51/S FILL
XFILL_7_AOI21X1_25 BUFX2_43/A DFFSR_97/S FILL
XFILL_15_DFFSR_39 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_30_DFFSR_111 INVX1_8/gnd DFFSR_5/S FILL
XFILL_3_DFFSR_184 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_1_OAI21X1_238 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_6_AOI21X1_28 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_20_DFFSR_114 DFFSR_71/gnd DFFSR_45/S FILL
XDFFPOSX1_8 INVX1_250/A CLKBUF1_15/Y OAI22X1_3/Y DFFSR_79/gnd DFFSR_36/S DFFPOSX1
XFILL_7_DFFPOSX1_28 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_5_AOI21X1_31 INVX1_23/gnd DFFSR_186/S FILL
XFILL_10_DFFSR_117 INVX1_23/gnd DFFSR_91/S FILL
XFILL_4_NAND2X1_190 BUFX2_35/A DFFSR_97/S FILL
XAOI21X1_28 NAND3X1_85/Y NAND3X1_88/Y AOI21X1_35/A DFFSR_71/gnd OAI22X1_3/C DFFSR_10/S
+ AOI21X1
XFILL_4_AOI21X1_34 INVX1_94/gnd DFFSR_25/S FILL
XFILL_3_NAND2X1_5 INVX1_8/gnd DFFSR_7/S FILL
XFILL_50_DFFSR_56 INVX1_2/gnd DFFSR_51/S FILL
XFILL_3_AOI21X1_37 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_0_INVX1_268 INVX1_8/gnd DFFSR_7/S FILL
XINVX1_378 INVX1_378/A INVX1_8/gnd INVX1_378/Y DFFSR_7/S INVX1
XFILL_39_DFFSR_96 INVX1_2/gnd DFFSR_1/S FILL
XFILL_2_OAI21X1_172 BUFX2_36/A DFFSR_6/S FILL
XFILL_0_AND2X2_5 BUFX2_37/A DFFSR_81/S FILL
XFILL_2_AOI21X1_40 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_23_DFFSR_46 BUFX2_36/A DFFSR_6/S FILL
XFILL_3_OAI22X1_4 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_6_DFFSR_53 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_5_NAND2X1_124 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_6_DFFSR_111 INVX1_8/gnd DFFSR_5/S FILL
XFILL_1_AOI21X1_43 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_12_DFFSR_86 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_47_DFFSR_142 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_0_AOI21X1_46 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_37_DFFSR_145 INVX1_23/gnd DFFSR_186/S FILL
XBUFX2_31 BUFX2_31/A DFFSR_1/gnd dout[5] DFFSR_9/S BUFX2
XFILL_27_DFFSR_148 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_3_INVX1_195 INVX1_23/gnd DFFSR_186/S FILL
XFILL_2_NAND2X1_286 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_3_OAI21X1_106 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_17_DFFSR_151 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_48_3 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_8_OAI21X1_70 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_6_NAND2X1_91 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_7_OAI21X1_73 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_3_NAND2X1_220 BUFX2_35/A DFFSR_14/S FILL
XFILL_6_OAI21X1_76 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_31_DFFSR_53 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_3_INVX1_47 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_20_DFFSR_93 INVX1_2/gnd DFFSR_51/S FILL
XFILL_42_DFFSR_13 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_5_NAND2X1_94 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_2_NOR2X1_30 DFFSR_73/gnd DFFSR_57/S FILL
XNAND2X1_91 BUFX2_25/Y DFFSR_83/Q BUFX2_5/gnd OAI21X1_91/C DFFSR_23/S NAND2X1
XFILL_4_NAND2X1_97 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_5_OAI21X1_79 INVX1_89/gnd DFFSR_36/S FILL
XFILL_3_DFFSR_148 DFFSR_89/gnd DFFSR_92/S FILL
XOAI21X1_76 BUFX2_19/Y INVX1_86/Y OAI21X1_76/C BUFX2_19/gnd DFFSR_76/D DFFSR_54/S
+ OAI21X1
XFILL_2_NAND3X1_118 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_1_INVX1_412 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_2_BUFX2_38 BUFX2_37/A DFFSR_81/S FILL
XFILL_4_OAI21X1_82 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_44_DFFSR_179 INVX1_2/gnd DFFSR_1/S FILL
XFILL_1_OAI21X1_202 BUFX2_35/A DFFSR_14/S FILL
XFILL_4_NAND2X1_154 BUFX2_37/A DFFSR_8/S FILL
XFILL_3_OAI21X1_85 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_34_DFFSR_182 INVX1_89/gnd DFFSR_36/S FILL
XFILL_24_DFFSR_185 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_2_OAI21X1_88 INVX1_4/gnd DFFSR_4/S FILL
XFILL_21_DFFSR_4 INVX1_4/gnd DFFSR_4/S FILL
XFILL_50_DFFSR_20 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_1_OAI21X1_91 BUFX2_43/A DFFSR_97/S FILL
XFILL_0_INVX1_232 BUFX2_37/A DFFSR_8/S FILL
XFILL_39_DFFSR_60 BUFX2_37/A DFFSR_8/S FILL
XFILL_0_INVX1_94 INVX1_94/gnd DFFSR_52/S FILL
XINVX1_342 INVX1_342/A INVX1_8/gnd INVX1_342/Y DFFSR_7/S INVX1
XFILL_14_DFFSR_188 INVX1_2/gnd DFFSR_1/S FILL
XFILL_16_DFFPOSX1_11 INVX1_4/gnd DFFSR_4/S FILL
XFILL_0_OAI21X1_94 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_5_BUFX2_5 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_4_INVX1_339 BUFX2_36/A DFFSR_8/S FILL
XBUFX2_9 rst BUFX2_37/A BUFX2_9/Y DFFSR_8/S BUFX2
XFILL_23_DFFSR_10 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_2_OAI21X1_136 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_6_DFFSR_17 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_12_DFFSR_50 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_47_DFFSR_106 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_37_DFFSR_109 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_0_AOI21X1_10 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_0_DFFSR_185 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_17_3_0 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_2_NAND2X1_250 INVX1_8/gnd DFFSR_5/S FILL
XFILL_27_DFFSR_112 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_17_DFFSR_115 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_3_INVX1_159 INVX1_94/gnd DFFSR_52/S FILL
XFILL_47_DFFSR_67 INVX1_2/gnd DFFSR_51/S FILL
XFILL_15_5_1 BUFX2_37/A DFFSR_81/S FILL
XFILL_8_OAI21X1_34 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_0_NAND2X1_6 INVX1_23/gnd DFFSR_186/S FILL
XFILL_7_OAI21X1_37 INVX1_89/gnd DFFSR_2/S FILL
XFILL_6_NAND2X1_55 INVX1_89/gnd DFFSR_2/S FILL
XFILL_31_DFFSR_17 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_20_DFFSR_57 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_3_INVX1_11 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_3_DFFSR_64 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_0_OAI21X1_232 BUFX2_35/A DFFSR_97/S FILL
XFILL_3_NAND2X1_184 BUFX2_37/A DFFSR_8/S FILL
XFILL_6_OAI21X1_40 INVX1_8/gnd DFFSR_7/S FILL
XFILL_5_NAND2X1_58 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_6_DFFPOSX1_22 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_4_NAND2X1_61 BUFX2_37/A DFFSR_81/S FILL
XFILL_5_OAI21X1_43 BUFX2_8/gnd DFFSR_10/S FILL
XNAND2X1_55 DFFSR_36/S INVX1_53/A INVX1_89/gnd OAI21X1_55/C DFFSR_2/S NAND2X1
XFILL_1_INVX1_376 INVX1_8/gnd DFFSR_7/S FILL
XFILL_4_OAI21X1_46 BUFX2_37/A DFFSR_81/S FILL
XOAI21X1_40 DFFSR_7/S INVX1_45/Y OAI21X1_40/C INVX1_8/gnd DFFSR_40/D DFFSR_7/S OAI21X1
XFILL_3_DFFSR_112 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_3_NAND2X1_64 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_0_OAI22X1_5 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_44_DFFSR_143 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_2_NAND2X1_67 INVX1_2/gnd DFFSR_1/S FILL
XFILL_1_OAI21X1_166 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_3_OAI21X1_49 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_34_DFFSR_146 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_2_OAI21X1_52 INVX1_94/gnd DFFSR_25/S FILL
XFILL_1_NAND2X1_70 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_4_NAND2X1_118 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_0_INVX1_196 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_24_DFFSR_149 INVX1_23/gnd DFFSR_91/S FILL
XFILL_1_OAI21X1_55 INVX1_89/gnd DFFSR_2/S FILL
XFILL_39_DFFSR_24 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_0_INVX1_58 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_0_NAND2X1_73 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_14_DFFSR_152 BUFX2_5/gnd DFFSR_23/S FILL
XINVX1_306 DFFSR_14/Q INVX1_94/gnd INVX1_306/Y DFFSR_25/S INVX1
XFILL_0_OAI21X1_58 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_28_DFFSR_64 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_2_OAI21X1_100 INVX1_23/gnd DFFSR_91/S FILL
XFILL_25_DFFPOSX1_30 BUFX2_43/A DFFSR_97/S FILL
XFILL_4_INVX1_303 INVX1_94/gnd DFFSR_25/S FILL
XFILL_1_NAND2X1_280 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_12_DFFSR_14 BUFX2_35/A DFFSR_14/S FILL
XFILL_0_DFFSR_149 INVX1_23/gnd DFFSR_91/S FILL
XNOR2X1_2 NOR2X1_2/A BUFX2_7/Y BUFX2_7/gnd AND2X2_1/B DFFSR_81/S NOR2X1
XFILL_2_NAND2X1_214 BUFX2_35/A DFFSR_97/S FILL
XFILL_3_INVX1_123 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_25_0_1 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_41_DFFSR_180 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_31_DFFSR_183 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_47_DFFSR_31 BUFX2_35/A DFFSR_97/S FILL
XFILL_1_NAND3X1_112 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_36_DFFSR_71 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_21_DFFSR_186 INVX1_23/gnd DFFSR_186/S FILL
XFILL_23_2_2 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_6_NAND2X1_19 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_3_NAND2X1_148 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_5_1_1 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_3_DFFSR_28 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_5_NAND2X1_22 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_0_OAI21X1_196 INVX1_94/gnd DFFSR_25/S FILL
XFILL_20_DFFSR_21 INVX1_2/gnd DFFSR_1/S FILL
XFILL_9_OAI21X1_251 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_4_NAND2X1_25 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_11_DFFSR_189 DFFSR_1/gnd DFFSR_1/S FILL
XNAND2X1_19 DFFSR_1/S DFFSR_11/Q DFFSR_1/gnd OAI21X1_19/C DFFSR_1/S NAND2X1
XFILL_2_NOR2X1_9 BUFX2_43/A DFFSR_97/S FILL
XFILL_11_OAI22X1_66 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_1_INVX1_340 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_3_3_2 INVX1_23/gnd DFFSR_91/S FILL
XFILL_44_DFFSR_107 BUFX2_36/A DFFSR_8/S FILL
XFILL_3_NAND2X1_28 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_4_OAI21X1_10 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_9_DFFSR_3 DFFSR_3/gnd DFFSR_4/S FILL
XDFFPOSX1_22 AND2X2_8/A CLKBUF1_13/Y XOR2X1_10/Y BUFX2_16/gnd DFFSR_11/S DFFPOSX1
XFILL_7_DFFSR_183 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_2_NAND2X1_31 BUFX2_43/A DFFSR_97/S FILL
XFILL_44_DFFSR_78 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_1_OAI21X1_130 INVX1_4/gnd DFFSR_4/S FILL
XFILL_3_OAI21X1_13 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_34_DFFSR_110 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_24_DFFSR_113 INVX1_23/gnd DFFSR_186/S FILL
XFILL_8_NAND3X1_90 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_2_OAI21X1_16 INVX1_89/gnd DFFSR_36/S FILL
XFILL_1_NAND2X1_34 INVX1_2/gnd DFFSR_1/S FILL
XFILL_17_DFFSR_68 BUFX2_35/A DFFSR_14/S FILL
XFILL_28_DFFSR_28 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_0_INVX1_160 BUFX2_19/gnd DFFSR_52/S FILL
XINVX1_270 DFFSR_25/Q DFFSR_79/gnd INVX1_270/Y DFFSR_36/S INVX1
XFILL_14_DFFSR_116 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_0_NAND2X1_37 INVX1_8/gnd DFFSR_5/S FILL
XFILL_1_OAI21X1_19 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_0_INVX1_22 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_0_DFFSR_75 INVX1_4/gnd DFFSR_51/S FILL
XFILL_7_NAND3X1_93 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_1_NAND2X1_244 INVX1_94/gnd DFFSR_52/S FILL
XFILL_0_OAI21X1_22 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_11_OAI22X1_9 INVX1_8/gnd DFFSR_5/S FILL
XFILL_6_NAND3X1_96 BUFX2_43/A DFFSR_97/S FILL
XFILL_7_OR2X2_3 BUFX2_43/A DFFSR_23/S FILL
XFILL_4_XOR2X1_5 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_5_NAND3X1_99 BUFX2_6/gnd DFFSR_14/S FILL
XNAND3X1_96 NAND3X1_94/B NAND3X1_94/C INVX1_259/Y BUFX2_43/A NAND3X1_98/C DFFSR_97/S
+ NAND3X1
XFILL_7_OAI22X1_3 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_33_DFFSR_7 INVX1_8/gnd DFFSR_7/S FILL
XFILL_0_DFFSR_113 INVX1_23/gnd DFFSR_186/S FILL
XFILL_5_DFFPOSX1_16 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_2_NAND2X1_178 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_36_DFFSR_35 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_41_DFFSR_144 INVX1_8/gnd DFFSR_5/S FILL
XFILL_8_DFFSR_82 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_25_DFFSR_75 INVX1_4/gnd DFFSR_51/S FILL
XFILL_31_DFFSR_147 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_21_DFFSR_150 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_11_DFFSR_153 BUFX2_36/A DFFSR_8/S FILL
XFILL_0_OAI21X1_160 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_3_NAND2X1_112 INVX1_4/gnd DFFSR_4/S FILL
XFILL_6_NOR2X1_29 BUFX2_37/A DFFSR_81/S FILL
XFILL_1_INVX1_304 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_1_AOI22X1_12 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_7_DFFSR_147 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_0_NAND2X1_274 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_10_OAI22X1_33 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_33_DFFSR_82 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_44_DFFSR_42 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_24_DFFPOSX1_24 BUFX2_43/A DFFSR_23/S FILL
XFILL_9_NAND3X1_51 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_48_DFFSR_178 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_38_DFFSR_181 INVX1_23/gnd DFFSR_186/S FILL
XFILL_8_NAND3X1_54 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_0_DFFSR_39 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_9_OAI22X1_36 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_0_INVX1_124 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_8_OAI22X1_39 BUFX2_37/A DFFSR_8/S FILL
XFILL_7_NAND3X1_57 BUFX2_19/gnd DFFSR_54/S FILL
XINVX1_234 NOR2X1_5/A BUFX2_17/gnd INVX1_234/Y DFFSR_57/S INVX1
XFILL_28_DFFSR_184 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_17_DFFSR_32 INVX1_2/gnd DFFSR_1/S FILL
XFILL_1_NAND2X1_208 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_6_NAND3X1_60 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_7_OAI22X1_42 INVX1_8/gnd DFFSR_7/S FILL
XFILL_18_DFFSR_187 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_5_NAND3X1_63 BUFX2_43/A DFFSR_23/S FILL
XFILL_6_OAI22X1_45 INVX1_89/gnd DFFSR_2/S FILL
XFILL_41_DFFSR_89 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_4_NAND3X1_66 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_0_NAND3X1_106 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_5_OAI22X1_48 BUFX2_37/A DFFSR_81/S FILL
XFILL_10_XOR2X1_2 BUFX2_8/gnd DFFSR_10/S FILL
XNAND3X1_60 INVX1_244/A NAND3X1_60/B NAND3X1_60/C DFFSR_71/gnd NAND3X1_60/Y DFFSR_10/S
+ NAND3X1
XFILL_3_NAND3X1_69 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_4_OAI22X1_51 BUFX2_7/gnd DFFSR_81/S FILL
XOAI22X1_45 INVX1_349/Y OAI22X1_49/D INVX1_348/Y OAI22X1_52/D INVX1_89/gnd NOR2X1_32/B
+ DFFSR_2/S OAI22X1
XFILL_2_NAND3X1_72 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_3_OAI22X1_54 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_2_NAND2X1_142 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_41_DFFSR_108 INVX1_89/gnd DFFSR_2/S FILL
XFILL_8_OAI21X1_245 DFFSR_5/gnd DFFSR_2/S FILL
XDFFSR_187 BUFX2_29/A DFFSR_3/CLK DFFSR_185/R DFFSR_11/S DFFSR_187/D BUFX2_16/gnd
+ DFFSR_11/S DFFSR
XFILL_1_NAND3X1_75 BUFX2_35/A DFFSR_97/S FILL
XFILL_8_DFFSR_46 BUFX2_36/A DFFSR_6/S FILL
XFILL_25_DFFSR_39 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_14_DFFSR_79 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_31_DFFSR_111 INVX1_8/gnd DFFSR_5/S FILL
XFILL_2_OAI22X1_57 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_4_DFFSR_184 DFFSR_1/gnd DFFSR_9/S FILL
XNAND2X1_8 DFFSR_6/S INVX1_413/A BUFX2_5/gnd NAND2X1_8/Y DFFSR_6/S NAND2X1
XFILL_21_DFFSR_114 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_0_NAND3X1_78 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_0_OAI21X1_124 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_1_OAI22X1_60 INVX1_8/gnd DFFSR_5/S FILL
XFILL_11_DFFSR_117 INVX1_23/gnd DFFSR_91/S FILL
XFILL_0_OAI22X1_63 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_4_NAND2X1_5 INVX1_8/gnd DFFSR_7/S FILL
XFILL_1_INVX1_268 INVX1_8/gnd DFFSR_7/S FILL
XFILL_49_DFFSR_96 INVX1_2/gnd DFFSR_1/S FILL
XFILL_20_DFFSR_1 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_24_3_0 DFFSR_71/gnd DFFSR_10/S FILL
XOAI22X1_7 INVX1_270/Y OAI22X1_7/B INVX1_269/Y OAI22X1_7/D DFFSR_5/gnd OAI22X1_7/Y
+ DFFSR_5/S OAI22X1
XFILL_33_DFFSR_46 BUFX2_36/A DFFSR_6/S FILL
XINVX1_80 INVX1_80/A BUFX2_8/gnd INVX1_80/Y DFFSR_10/S INVX1
XFILL_0_NAND2X1_238 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_7_DFFSR_111 INVX1_8/gnd DFFSR_5/S FILL
XFILL_22_DFFSR_86 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_5_DFFSR_93 INVX1_2/gnd DFFSR_51/S FILL
XFILL_4_OAI22X1_4 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_48_DFFSR_142 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_22_5_1 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_8_NAND3X1_18 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_38_DFFSR_145 INVX1_23/gnd DFFSR_186/S FILL
XFILL_4_4_0 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_4_BUFX2_2 BUFX2_43/A DFFSR_23/S FILL
XINVX1_198 DFFSR_164/Q DFFSR_5/gnd INVX1_198/Y DFFSR_2/S INVX1
XFILL_28_DFFSR_148 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_4_INVX1_195 INVX1_23/gnd DFFSR_186/S FILL
XFILL_1_NAND2X1_172 BUFX2_36/A DFFSR_6/S FILL
XFILL_7_NAND3X1_21 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_4_DFFPOSX1_10 INVX1_8/gnd DFFSR_5/S FILL
XFILL_35_5 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_4_BUFX2_31 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_6_NAND3X1_24 BUFX2_37/A DFFSR_8/S FILL
XFILL_18_DFFSR_151 BUFX2_7/gnd DFFSR_81/S FILL
XNAND3X1_24 OAI22X1_2/C AOI22X1_5/C NAND3X1_24/C BUFX2_37/A AOI21X1_4/A DFFSR_8/S
+ NAND3X1
XFILL_5_NAND3X1_27 BUFX2_37/A DFFSR_81/S FILL
XFILL_4_NAND3X1_30 INVX1_94/gnd DFFSR_52/S FILL
XFILL_41_DFFSR_53 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_2_INVX1_87 INVX1_89/gnd DFFSR_36/S FILL
XFILL_13_DFFPOSX1_29 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_30_DFFSR_93 INVX1_2/gnd DFFSR_51/S FILL
XFILL_5_OAI22X1_12 INVX1_4/gnd DFFSR_51/S FILL
XFILL_3_NOR2X1_30 DFFSR_73/gnd DFFSR_57/S FILL
XDFFSR_151 INVX1_176/A CLKBUF1_11/Y INVX1_177/Y DFFSR_81/S DFFSR_151/D BUFX2_7/gnd
+ DFFSR_81/S DFFSR
XFILL_3_NAND3X1_33 INVX1_8/gnd DFFSR_7/S FILL
XFILL_8_OAI21X1_209 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_2_NAND2X1_106 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_4_OAI22X1_15 INVX1_4/gnd DFFSR_4/S FILL
XFILL_4_DFFSR_148 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_2_NAND3X1_36 BUFX2_35/A DFFSR_97/S FILL
XFILL_14_DFFSR_43 INVX1_94/gnd DFFSR_25/S FILL
XFILL_3_OAI22X1_18 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_8_DFFSR_10 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_2_INVX1_412 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_1_NAND3X1_39 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_45_DFFSR_179 INVX1_2/gnd DFFSR_1/S FILL
XFILL_2_OAI22X1_21 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_0_NAND3X1_42 BUFX2_43/A DFFSR_23/S FILL
XFILL_1_OAI22X1_24 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_35_DFFSR_182 INVX1_89/gnd DFFSR_36/S FILL
XFILL_25_DFFSR_185 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_23_DFFPOSX1_18 BUFX2_37/A DFFSR_8/S FILL
XFILL_0_OAI22X1_27 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_1_INVX1_232 BUFX2_37/A DFFSR_8/S FILL
XFILL_49_DFFSR_60 BUFX2_37/A DFFSR_8/S FILL
XFILL_15_DFFSR_188 INVX1_2/gnd DFFSR_1/S FILL
XFILL_0_NAND2X1_202 BUFX2_35/A DFFSR_97/S FILL
XDFFSR_97 DFFSR_97/Q CLKBUF1_7/Y DFFSR_97/R DFFSR_97/S DFFSR_97/D BUFX2_35/A DFFSR_97/S
+ DFFSR
XFILL_33_DFFSR_10 DFFSR_71/gnd DFFSR_10/S FILL
XINVX1_44 DFFSR_39/Q DFFSR_79/gnd INVX1_44/Y DFFSR_36/S INVX1
XFILL_32_0_1 INVX1_8/gnd DFFSR_5/S FILL
XFILL_5_DFFSR_57 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_11_DFFSR_90 INVX1_2/gnd DFFSR_1/S FILL
XFILL_22_DFFSR_50 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_48_DFFSR_106 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_38_DFFSR_109 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_30_2_2 DFFSR_5/gnd DFFSR_2/S FILL
XINVX1_162 DFFSR_144/Q INVX1_8/gnd INVX1_162/Y DFFSR_7/S INVX1
XFILL_1_DFFSR_185 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_28_DFFSR_112 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_18_DFFSR_115 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_4_INVX1_159 INVX1_94/gnd DFFSR_52/S FILL
XFILL_1_NAND2X1_136 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_7_OAI21X1_239 INVX1_4/gnd DFFSR_4/S FILL
XFILL_1_NAND2X1_6 INVX1_23/gnd DFFSR_186/S FILL
XFILL_2_INVX1_51 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_41_DFFSR_17 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_30_DFFSR_57 DFFSR_73/gnd DFFSR_57/S FILL
XDFFSR_115 DFFSR_115/Q INVX1_172/A DFFSR_113/R DFFSR_14/S DFFSR_115/D BUFX2_6/gnd
+ DFFSR_14/S DFFSR
XFILL_19_DFFSR_97 BUFX2_35/A DFFSR_97/S FILL
XFILL_8_OAI21X1_173 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_2_INVX1_376 INVX1_8/gnd DFFSR_7/S FILL
XFILL_1_BUFX2_42 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_4_DFFSR_112 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_45_DFFSR_143 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_1_OAI22X1_5 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_35_DFFSR_146 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_11_DFFSR_8 BUFX2_36/A DFFSR_8/S FILL
XFILL_25_DFFSR_149 INVX1_23/gnd DFFSR_91/S FILL
XFILL_1_INVX1_196 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_15_DFFSR_152 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_49_DFFSR_24 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_38_DFFSR_64 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_0_NAND2X1_166 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_22_DFFSR_14 BUFX2_35/A DFFSR_14/S FILL
XDFFSR_61 DFFSR_61/Q DFFSR_20/CLK DFFSR_61/R DFFSR_6/S DFFSR_61/D BUFX2_5/gnd DFFSR_6/S
+ DFFSR
XFILL_11_DFFSR_54 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_5_DFFSR_21 INVX1_2/gnd DFFSR_1/S FILL
XFILL_0_NOR2X1_31 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_4_NOR2X1_2 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_8_NAND3X1_119 DFFSR_5/gnd DFFSR_2/S FILL
XINVX1_126 INVX1_391/A BUFX2_16/gnd INVX1_126/Y DFFSR_65/S INVX1
XFILL_12_DFFPOSX1_23 INVX1_23/gnd DFFSR_91/S FILL
XFILL_1_DFFSR_149 INVX1_23/gnd DFFSR_91/S FILL
XFILL_1_NAND2X1_100 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_7_OAI21X1_203 BUFX2_35/A DFFSR_14/S FILL
XFILL_4_INVX1_123 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_42_DFFSR_180 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_32_DFFSR_4 INVX1_4/gnd DFFSR_4/S FILL
XFILL_32_DFFSR_183 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_46_DFFSR_71 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_22_DFFSR_186 INVX1_23/gnd DFFSR_186/S FILL
XFILL_2_DFFSR_68 BUFX2_35/A DFFSR_14/S FILL
XFILL_19_DFFSR_61 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_30_DFFSR_21 INVX1_2/gnd DFFSR_1/S FILL
XFILL_2_INVX1_15 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_8_OAI21X1_137 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_22_DFFPOSX1_12 INVX1_8/gnd DFFSR_5/S FILL
XFILL_12_DFFSR_189 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_2_INVX1_340 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_45_DFFSR_107 BUFX2_36/A DFFSR_8/S FILL
XFILL_8_DFFSR_183 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_35_DFFSR_110 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_25_DFFSR_113 INVX1_23/gnd DFFSR_186/S FILL
XFILL_27_DFFSR_68 BUFX2_35/A DFFSR_14/S FILL
XFILL_38_DFFSR_28 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_1_INVX1_160 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_15_DFFSR_116 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_6_OAI21X1_233 BUFX2_36/A DFFSR_8/S FILL
XDFFSR_25 DFFSR_25/Q DFFSR_52/CLK DFFSR_31/R DFFSR_25/S DFFSR_25/D BUFX2_8/gnd DFFSR_25/S
+ DFFSR
XFILL_11_DFFSR_18 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_0_NAND2X1_130 INVX1_4/gnd DFFSR_4/S FILL
XFILL_1_DFFSR_113 INVX1_23/gnd DFFSR_186/S FILL
XFILL_17_2 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_8_OAI22X1_3 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_7_OAI21X1_167 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_46_DFFSR_35 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_42_DFFSR_144 INVX1_8/gnd DFFSR_5/S FILL
XFILL_35_DFFSR_75 INVX1_4/gnd DFFSR_51/S FILL
XFILL_32_DFFSR_147 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_22_DFFSR_150 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_31_3_0 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_2_DFFSR_32 INVX1_2/gnd DFFSR_1/S FILL
XFILL_12_DFFSR_153 BUFX2_36/A DFFSR_8/S FILL
XFILL_19_DFFSR_25 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_21_CLKBUF1_12 BUFX2_43/A DFFSR_23/S FILL
XFILL_2_INVX1_304 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_29_5_1 INVX1_89/gnd DFFSR_2/S FILL
XFILL_8_OAI21X1_101 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_20_CLKBUF1_15 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_8_DFFSR_147 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_19_CLKBUF1_18 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_43_DFFSR_82 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_5_OAI21X1_263 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_18_CLKBUF1_21 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_49_DFFSR_178 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_17_CLKBUF1_24 INVX1_23/gnd DFFSR_186/S FILL
XFILL_39_DFFSR_181 INVX1_23/gnd DFFSR_186/S FILL
XFILL_1_INVX1_124 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_7_NAND3X1_113 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_16_DFFSR_72 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_29_DFFSR_184 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_27_DFFSR_32 INVX1_2/gnd DFFSR_1/S FILL
XFILL_11_DFFPOSX1_17 BUFX2_37/A DFFSR_8/S FILL
XFILL_6_OAI21X1_197 INVX1_8/gnd DFFSR_7/S FILL
XFILL_19_DFFSR_187 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_3_XOR2X1_9 BUFX2_19/gnd DFFSR_52/S FILL
XOAI21X1_233 NOR2X1_10/A NOR2X1_10/B INVX1_257/Y BUFX2_36/A NAND3X1_90/C DFFSR_8/S
+ OAI21X1
XFILL_42_DFFSR_108 INVX1_89/gnd DFFSR_2/S FILL
XFILL_7_OAI21X1_131 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_35_DFFSR_39 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_24_DFFSR_79 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_32_DFFSR_111 INVX1_8/gnd DFFSR_5/S FILL
XFILL_5_DFFSR_184 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_7_DFFSR_86 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_22_DFFSR_114 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_1_DFFPOSX1_28 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_39_0_1 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_12_DFFSR_117 INVX1_23/gnd DFFSR_91/S FILL
XFILL_5_NAND2X1_5 INVX1_8/gnd DFFSR_7/S FILL
XFILL_6_BUFX2_24 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_44_DFFSR_7 INVX1_8/gnd DFFSR_7/S FILL
XFILL_2_INVX1_268 INVX1_8/gnd DFFSR_7/S FILL
XFILL_37_2_2 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_5_OAI21X1_227 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_43_DFFSR_46 BUFX2_36/A DFFSR_6/S FILL
XFILL_4_INVX1_80 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_8_DFFSR_111 INVX1_8/gnd DFFSR_5/S FILL
XFILL_32_DFFSR_86 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_5_OAI22X1_4 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_49_DFFSR_142 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_39_DFFSR_145 INVX1_23/gnd DFFSR_186/S FILL
XFILL_22_7 INVX1_94/gnd DFFSR_25/S FILL
XFILL_16_DFFSR_36 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_29_DFFSR_148 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_39_2 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_6_OAI21X1_161 INVX1_23/gnd DFFSR_186/S FILL
XFILL_19_DFFSR_151 BUFX2_7/gnd DFFSR_81/S FILL
XNOR2X1_33 NOR2X1_33/A NOR2X1_33/B BUFX2_37/A NOR2X1_33/Y DFFSR_81/S NOR2X1
XFILL_51_DFFSR_53 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_40_DFFSR_93 INVX1_2/gnd DFFSR_51/S FILL
XFILL_4_NOR2X1_30 DFFSR_73/gnd DFFSR_57/S FILL
XOAI21X1_197 AOI21X1_10/Y AOI21X1_11/Y INVX1_236/A INVX1_8/gnd AOI21X1_17/A DFFSR_7/S
+ OAI21X1
XFILL_1_AND2X2_2 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_13_DFFSR_83 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_24_DFFSR_43 INVX1_94/gnd DFFSR_25/S FILL
XFILL_3_INVX1_412 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_6_NAND2X1_275 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_7_DFFSR_50 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_5_DFFSR_148 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_46_DFFSR_179 INVX1_2/gnd DFFSR_1/S FILL
XFILL_36_DFFSR_182 INVX1_89/gnd DFFSR_36/S FILL
XFILL_4_OAI21X1_257 INVX1_2/gnd DFFSR_51/S FILL
XFILL_26_DFFSR_185 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_9_CLKBUF1_12 BUFX2_43/A DFFSR_23/S FILL
XFILL_2_INVX1_232 BUFX2_37/A DFFSR_8/S FILL
XFILL_6_NAND3X1_107 BUFX2_43/A DFFSR_97/S FILL
XFILL_10_DFFSR_5 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_8_CLKBUF1_15 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_16_DFFSR_188 INVX1_2/gnd DFFSR_1/S FILL
XFILL_9_AND2X2_9 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_4_DFFSR_97 BUFX2_35/A DFFSR_97/S FILL
XFILL_7_CLKBUF1_18 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_43_DFFSR_10 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_10_DFFPOSX1_11 INVX1_4/gnd DFFSR_4/S FILL
XFILL_32_DFFSR_50 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_5_OAI21X1_191 BUFX2_37/A DFFSR_8/S FILL
XFILL_6_CLKBUF1_21 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_49_DFFSR_106 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_21_DFFSR_90 INVX1_2/gnd DFFSR_1/S FILL
XFILL_5_CLKBUF1_24 INVX1_23/gnd DFFSR_186/S FILL
XFILL_39_DFFSR_109 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_2_DFFSR_185 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_3_BUFX2_35 BUFX2_35/A DFFSR_14/S FILL
XOR2X2_1 OR2X2_1/A OR2X2_1/B BUFX2_8/gnd OR2X2_1/Y DFFSR_10/S OR2X2
XCLKBUF1_21 INVX1_402/Y BUFX2_17/gnd DFFSR_15/CLK DFFSR_7/S CLKBUF1
XFILL_29_DFFSR_112 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_19_DFFSR_115 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_6_OAI21X1_125 BUFX2_35/A DFFSR_14/S FILL
XFILL_31_DFFSR_1 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_2_NAND2X1_6 INVX1_23/gnd DFFSR_186/S FILL
XOAI21X1_161 BUFX2_2/Y INVX1_195/Y NAND2X1_161/Y INVX1_23/gnd DFFSR_161/D DFFSR_186/S
+ OAI21X1
XFILL_29_DFFSR_97 BUFX2_35/A DFFSR_97/S FILL
XFILL_1_INVX1_91 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_40_DFFSR_57 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_0_DFFPOSX1_22 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_11_0_2 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_6_NAND2X1_239 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_3_INVX1_376 INVX1_8/gnd DFFSR_7/S FILL
XFILL_7_DFFSR_14 BUFX2_35/A DFFSR_14/S FILL
XFILL_13_DFFSR_47 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_5_DFFSR_112 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_46_DFFSR_143 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_2_OAI22X1_5 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_36_DFFSR_146 DFFSR_89/gnd DFFSR_92/S FILL
XNAND2X1_275 AND2X2_17/B AND2X2_17/A DFFSR_5/gnd XOR2X1_14/A DFFSR_5/S NAND2X1
XFILL_26_DFFSR_149 INVX1_23/gnd DFFSR_91/S FILL
XFILL_4_OAI21X1_221 BUFX2_35/A DFFSR_14/S FILL
XFILL_2_INVX1_196 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_16_DFFSR_152 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_48_DFFSR_64 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_32_DFFSR_14 BUFX2_35/A DFFSR_14/S FILL
XFILL_19_DFFPOSX1_30 BUFX2_43/A DFFSR_97/S FILL
XFILL_4_DFFSR_61 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_21_DFFSR_54 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_5_OAI21X1_155 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_10_DFFSR_94 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_1_NOR2X1_31 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_0_INVX1_413 DFFSR_89/gnd DFFSR_92/S FILL
XNAND3X1_107 XOR2X1_8/A NAND3X1_105/Y NAND3X1_107/C BUFX2_43/A AOI21X1_39/B DFFSR_97/S
+ NAND3X1
XFILL_38_3_0 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_2_DFFSR_149 INVX1_23/gnd DFFSR_91/S FILL
XFILL_43_DFFSR_180 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_33_DFFSR_183 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_5_NAND2X1_269 INVX1_4/gnd DFFSR_4/S FILL
XFILL_36_5_1 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_23_DFFSR_186 INVX1_23/gnd DFFSR_186/S FILL
XFILL_29_DFFSR_61 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_1_INVX1_55 BUFX2_36/A DFFSR_8/S FILL
XFILL_40_DFFSR_21 INVX1_2/gnd DFFSR_1/S FILL
XFILL_3_OAI21X1_251 DFFSR_89/gnd DFFSR_92/S FILL
XOAI21X1_125 BUFX2_21/Y INVX1_141/Y OAI21X1_125/C BUFX2_35/A DFFSR_125/D DFFSR_14/S
+ OAI21X1
XFILL_13_DFFSR_189 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_6_NAND2X1_203 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_3_INVX1_340 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_13_DFFSR_11 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_5_NAND3X1_101 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_46_DFFSR_107 BUFX2_36/A DFFSR_8/S FILL
XFILL_9_DFFSR_183 DFFSR_89/gnd DFFSR_186/S FILL
XNAND2X1_239 NOR2X1_22/Y NOR2X1_23/Y DFFSR_79/gnd NAND2X1_70/B DFFSR_45/S NAND2X1
XFILL_36_DFFSR_110 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_26_DFFSR_113 INVX1_23/gnd DFFSR_186/S FILL
XFILL_4_OAI21X1_185 BUFX2_36/A DFFSR_8/S FILL
XFILL_37_DFFSR_68 BUFX2_35/A DFFSR_14/S FILL
XFILL_48_DFFSR_28 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_2_INVX1_160 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_16_DFFSR_116 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_4_DFFSR_25 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_21_DFFSR_18 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_5_OAI21X1_119 BUFX2_37/A DFFSR_8/S FILL
XFILL_10_DFFSR_58 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_0_INVX1_377 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_2_DFFSR_113 INVX1_23/gnd DFFSR_186/S FILL
XFILL_9_OAI22X1_3 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_3_NOR2X1_6 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_22_DFFSR_8 BUFX2_36/A DFFSR_8/S FILL
XFILL_5_NAND2X1_233 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_43_DFFSR_144 INVX1_8/gnd DFFSR_5/S FILL
XFILL_46_0_1 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_45_DFFSR_75 INVX1_4/gnd DFFSR_51/S FILL
XFILL_33_DFFSR_147 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_4_NAND3X1_131 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_23_DFFSR_150 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_44_2_2 INVX1_2/gnd DFFSR_51/S FILL
XFILL_1_INVX1_19 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_13_DFFSR_153 BUFX2_36/A DFFSR_8/S FILL
XFILL_6_BUFX2_9 BUFX2_37/A DFFSR_8/S FILL
XFILL_29_DFFSR_25 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_1_DFFSR_72 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_18_DFFSR_65 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_3_OAI21X1_215 BUFX2_43/A DFFSR_97/S FILL
XFILL_3_INVX1_304 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_6_NAND2X1_167 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_0_BUFX2_10 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_5_XOR2X1_2 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_9_DFFSR_147 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_4_OAI21X1_149 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_18_DFFPOSX1_24 BUFX2_43/A DFFSR_23/S FILL
XNAND2X1_203 AND2X2_6/Y AND2X2_10/Y BUFX2_5/gnd NAND3X1_37/C DFFSR_23/S NAND2X1
XFILL_20_DFFPOSX1_3 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_50_DFFSR_178 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_43_DFFSR_4 INVX1_4/gnd DFFSR_4/S FILL
XFILL_40_DFFSR_181 INVX1_23/gnd DFFSR_186/S FILL
XFILL_12_1_0 BUFX2_36/A DFFSR_6/S FILL
XFILL_19_DFFPOSX1_6 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_18_DFFPOSX1_9 BUFX2_37/A DFFSR_8/S FILL
XFILL_9_DFFSR_79 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_26_DFFSR_72 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_37_DFFSR_32 INVX1_2/gnd DFFSR_1/S FILL
XFILL_2_INVX1_124 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_10_3_1 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_30_DFFSR_184 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_10_DFFSR_22 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_4_NAND2X1_263 INVX1_2/gnd DFFSR_51/S FILL
XFILL_20_DFFSR_187 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_10_DFFSR_190 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_4_3 INVX1_23/gnd DFFSR_91/S FILL
XFILL_0_INVX1_341 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_43_DFFSR_108 INVX1_89/gnd DFFSR_2/S FILL
XFILL_2_OAI21X1_245 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_45_DFFSR_39 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_34_DFFSR_79 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_5_NAND2X1_197 INVX1_8/gnd DFFSR_5/S FILL
XFILL_33_DFFSR_111 INVX1_8/gnd DFFSR_5/S FILL
XFILL_6_DFFSR_184 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_23_DFFSR_114 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_1_DFFSR_36 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_18_DFFSR_29 INVX1_4/gnd DFFSR_4/S FILL
XFILL_13_DFFSR_117 INVX1_23/gnd DFFSR_91/S FILL
XFILL_3_OAI21X1_179 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_6_NAND2X1_5 INVX1_8/gnd DFFSR_7/S FILL
XFILL_3_INVX1_268 INVX1_8/gnd DFFSR_7/S FILL
XFILL_6_NAND2X1_131 DFFSR_9/gnd DFFSR_9/S FILL
XXOR2X1_6 XOR2X1_6/A XOR2X1_5/Y DFFSR_89/gnd XOR2X1_6/Y DFFSR_186/S XOR2X1
XFILL_9_DFFSR_111 INVX1_8/gnd DFFSR_5/S FILL
XFILL_42_DFFSR_86 DFFSR_1/gnd DFFSR_9/S FILL
XNAND2X1_167 BUFX2_4/Y INVX1_261/A DFFSR_9/gnd OAI21X1_167/C DFFSR_9/S NAND2X1
XFILL_4_OAI21X1_113 INVX1_23/gnd DFFSR_91/S FILL
XFILL_6_OAI22X1_4 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_50_DFFSR_142 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_40_DFFSR_145 INVX1_23/gnd DFFSR_186/S FILL
XFILL_15_DFFSR_76 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_9_DFFSR_43 INVX1_94/gnd DFFSR_25/S FILL
XFILL_26_4 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_26_DFFSR_36 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_30_DFFSR_148 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_4_NAND2X1_227 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_20_DFFSR_151 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_10_DFFSR_154 BUFX2_36/A DFFSR_6/S FILL
XFILL_18_0_2 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_0_INVX1_305 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_3_NAND3X1_125 INVX1_8/gnd DFFSR_5/S FILL
XINVX1_415 BUFX2_26/A DFFSR_9/gnd INVX1_415/Y DFFSR_9/S INVX1
XFILL_50_DFFSR_93 INVX1_2/gnd DFFSR_51/S FILL
XFILL_5_NOR2X1_30 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_5_NAND2X1_161 INVX1_23/gnd DFFSR_186/S FILL
XFILL_23_DFFSR_83 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_34_DFFSR_43 INVX1_94/gnd DFFSR_25/S FILL
XFILL_2_OAI21X1_209 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_6_DFFSR_90 INVX1_2/gnd DFFSR_1/S FILL
XFILL_6_DFFSR_148 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_47_DFFSR_179 INVX1_2/gnd DFFSR_1/S FILL
XFILL_37_DFFSR_182 INVX1_89/gnd DFFSR_36/S FILL
XFILL_5_BUFX2_28 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_17_DFFPOSX1_18 BUFX2_37/A DFFSR_8/S FILL
XFILL_27_DFFSR_185 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_3_INVX1_232 BUFX2_37/A DFFSR_8/S FILL
XFILL_3_OAI21X1_143 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_17_DFFSR_188 INVX1_2/gnd DFFSR_1/S FILL
XFILL_8_DFFPOSX1_3 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_3_INVX1_84 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_45_3_0 INVX1_2/gnd DFFSR_1/S FILL
XFILL_42_DFFSR_50 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_50_DFFSR_106 DFFSR_1/gnd DFFSR_1/S FILL
XNAND2X1_131 DFFSR_9/S NAND2X1_67/B DFFSR_9/gnd NAND2X1_131/Y DFFSR_9/S NAND2X1
XFILL_3_NAND2X1_257 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_31_DFFSR_90 INVX1_2/gnd DFFSR_1/S FILL
XFILL_40_DFFSR_109 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_8_AOI21X1_23 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_43_5_1 INVX1_4/gnd DFFSR_51/S FILL
XFILL_7_DFFPOSX1_6 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_3_DFFSR_185 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_7_AOI21X1_26 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_6_DFFPOSX1_9 BUFX2_37/A DFFSR_8/S FILL
XFILL_15_DFFSR_40 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_30_DFFSR_112 DFFSR_3/gnd DFFSR_65/S FILL
XDFFPOSX1_9 INVX1_261/A CLKBUF1_15/Y DFFPOSX1_9/D BUFX2_37/A DFFSR_8/S DFFPOSX1
XFILL_6_AOI21X1_29 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_20_DFFSR_115 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_5_AOI21X1_32 BUFX2_43/A DFFSR_23/S FILL
XFILL_4_NAND2X1_191 BUFX2_37/A DFFSR_8/S FILL
XFILL_7_DFFPOSX1_29 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_1_OAI21X1_239 INVX1_4/gnd DFFSR_4/S FILL
XFILL_3_NAND2X1_6 INVX1_23/gnd DFFSR_186/S FILL
XFILL_4_AOI21X1_35 INVX1_94/gnd DFFSR_25/S FILL
XAOI21X1_29 NAND3X1_60/C NAND3X1_60/B INVX1_244/Y DFFSR_71/gnd AOI21X1_29/Y DFFSR_45/S
+ AOI21X1
XFILL_10_DFFSR_118 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_39_DFFSR_97 BUFX2_35/A DFFSR_97/S FILL
XFILL_3_AOI21X1_38 BUFX2_36/A DFFSR_8/S FILL
XFILL_0_INVX1_269 DFFSR_5/gnd DFFSR_5/S FILL
XINVX1_379 DFFSR_70/Q BUFX2_17/gnd INVX1_379/Y DFFSR_57/S INVX1
XFILL_50_DFFSR_57 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_2_OAI21X1_173 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_2_AOI21X1_41 BUFX2_35/A DFFSR_14/S FILL
XFILL_0_AND2X2_6 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_4_INVX1_376 INVX1_8/gnd DFFSR_7/S FILL
XFILL_5_NAND2X1_125 BUFX2_35/A DFFSR_14/S FILL
XFILL_6_DFFSR_54 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_23_DFFSR_47 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_1_AOI21X1_44 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_12_DFFSR_87 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_6_DFFSR_112 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_0_AOI21X1_47 BUFX2_43/A DFFSR_23/S FILL
XFILL_47_DFFSR_143 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_3_OAI22X1_5 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_37_DFFSR_146 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_27_DFFSR_149 INVX1_23/gnd DFFSR_91/S FILL
XFILL_3_OAI21X1_107 BUFX2_36/A DFFSR_6/S FILL
XBUFX2_32 BUFX2_32/A DFFSR_9/gnd dout[6] DFFSR_9/S BUFX2
XFILL_3_INVX1_196 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_17_DFFSR_152 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_8_OAI21X1_71 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_48_4 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_6_NAND2X1_92 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_42_DFFSR_14 BUFX2_35/A DFFSR_14/S FILL
XFILL_31_DFFSR_54 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_7_OAI21X1_74 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_20_DFFSR_94 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_3_INVX1_48 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_2_NOR2X1_31 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_3_NAND2X1_221 BUFX2_6/gnd DFFSR_14/S FILL
XNAND2X1_92 BUFX2_20/Y DFFSR_84/Q BUFX2_5/gnd NAND2X1_92/Y DFFSR_23/S NAND2X1
XFILL_6_OAI21X1_77 INVX1_89/gnd DFFSR_36/S FILL
XFILL_5_NAND2X1_95 INVX1_89/gnd DFFSR_36/S FILL
XFILL_1_INVX1_413 DFFSR_89/gnd DFFSR_92/S FILL
XOAI21X1_77 BUFX2_17/Y INVX1_87/Y NAND2X1_77/Y INVX1_89/gnd DFFSR_77/D DFFSR_36/S
+ OAI21X1
XFILL_2_NAND3X1_119 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_4_NAND2X1_98 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_5_OAI21X1_80 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_3_DFFSR_149 INVX1_23/gnd DFFSR_91/S FILL
XFILL_2_BUFX2_39 BUFX2_43/A DFFSR_97/S FILL
XFILL_4_OAI21X1_83 INVX1_94/gnd DFFSR_52/S FILL
XFILL_44_DFFSR_180 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_1_OAI21X1_203 BUFX2_35/A DFFSR_14/S FILL
XFILL_4_NAND2X1_155 BUFX2_37/A DFFSR_81/S FILL
XFILL_3_OAI21X1_86 INVX1_4/gnd DFFSR_51/S FILL
XFILL_34_DFFSR_183 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_2_OAI21X1_89 BUFX2_35/A DFFSR_14/S FILL
XFILL_21_DFFSR_5 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_24_DFFSR_186 INVX1_23/gnd DFFSR_186/S FILL
XFILL_1_OAI21X1_92 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_39_DFFSR_61 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_0_INVX1_95 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_0_INVX1_233 BUFX2_7/gnd DFFSR_54/S FILL
XINVX1_343 DFFSR_82/Q DFFSR_1/gnd INVX1_343/Y DFFSR_1/S INVX1
XFILL_50_DFFSR_21 INVX1_2/gnd DFFSR_1/S FILL
XFILL_0_OAI21X1_95 INVX1_89/gnd DFFSR_36/S FILL
XFILL_14_DFFSR_189 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_19_1_0 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_2_OAI21X1_137 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_16_DFFPOSX1_12 INVX1_8/gnd DFFSR_5/S FILL
XFILL_6_DFFSR_18 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_4_INVX1_340 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_23_DFFSR_11 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_5_BUFX2_6 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_47_DFFSR_107 BUFX2_36/A DFFSR_8/S FILL
XFILL_12_DFFSR_51 INVX1_2/gnd DFFSR_51/S FILL
XFILL_0_AOI21X1_11 INVX1_8/gnd DFFSR_5/S FILL
XFILL_37_DFFSR_110 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_0_DFFSR_186 INVX1_23/gnd DFFSR_186/S FILL
XFILL_2_NAND2X1_251 BUFX2_35/A DFFSR_97/S FILL
XFILL_17_3_1 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_27_DFFSR_113 INVX1_23/gnd DFFSR_186/S FILL
XFILL_47_DFFSR_68 BUFX2_35/A DFFSR_14/S FILL
XFILL_3_INVX1_160 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_42_DFFSR_1 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_15_5_2 BUFX2_37/A DFFSR_81/S FILL
XFILL_17_DFFSR_116 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_8_OAI21X1_35 INVX1_8/gnd DFFSR_5/S FILL
XFILL_3_INVX1_12 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_0_NAND2X1_7 INVX1_89/gnd DFFSR_36/S FILL
XFILL_7_OAI21X1_38 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_6_NAND2X1_56 INVX1_4/gnd DFFSR_51/S FILL
XFILL_3_DFFSR_65 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_6_DFFPOSX1_23 INVX1_23/gnd DFFSR_91/S FILL
XFILL_0_OAI21X1_233 BUFX2_36/A DFFSR_8/S FILL
XFILL_3_NAND2X1_185 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_6_OAI21X1_41 INVX1_8/gnd DFFSR_7/S FILL
XFILL_31_DFFSR_18 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_5_NAND2X1_59 INVX1_2/gnd DFFSR_1/S FILL
XFILL_20_DFFSR_58 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_4_NAND2X1_62 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_5_OAI21X1_44 DFFSR_71/gnd DFFSR_45/S FILL
XNAND2X1_56 DFFSR_1/S INVX1_54/A INVX1_4/gnd NAND2X1_56/Y DFFSR_51/S NAND2X1
XFILL_1_INVX1_377 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_3_DFFSR_113 INVX1_23/gnd DFFSR_186/S FILL
XFILL_4_OAI21X1_47 INVX1_89/gnd DFFSR_2/S FILL
XOAI21X1_41 DFFSR_57/S INVX1_47/Y NAND2X1_41/Y INVX1_8/gnd DFFSR_41/D DFFSR_7/S OAI21X1
XFILL_3_NAND2X1_65 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_2_NAND2X1_68 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_44_DFFSR_144 INVX1_8/gnd DFFSR_5/S FILL
XFILL_3_OAI21X1_50 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_0_OAI22X1_6 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_34_DFFSR_147 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_4_NAND2X1_119 BUFX2_37/A DFFSR_8/S FILL
XFILL_1_OAI21X1_167 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_1_NAND2X1_71 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_2_OAI21X1_53 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_24_DFFSR_150 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_0_NAND2X1_74 INVX1_2/gnd DFFSR_1/S FILL
XFILL_1_OAI21X1_56 INVX1_2/gnd DFFSR_51/S FILL
XFILL_14_DFFSR_153 BUFX2_36/A DFFSR_8/S FILL
XINVX1_307 DFFSR_54/Q BUFX2_19/gnd INVX1_307/Y DFFSR_54/S INVX1
XFILL_0_INVX1_59 INVX1_94/gnd DFFSR_25/S FILL
XFILL_39_DFFSR_25 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_0_OAI21X1_59 INVX1_4/gnd DFFSR_51/S FILL
XFILL_0_INVX1_197 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_28_DFFSR_65 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_1_NAND2X1_281 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_4_INVX1_304 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_2_OAI21X1_101 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_12_DFFSR_15 INVX1_8/gnd DFFSR_7/S FILL
XFILL_25_DFFPOSX1_31 BUFX2_17/gnd DFFSR_57/S FILL
XNOR2X1_3 NOR2X1_3/A NOR2X1_3/B INVX1_94/gnd NOR2X1_3/Y DFFSR_25/S NOR2X1
XFILL_41_DFFSR_181 INVX1_23/gnd DFFSR_186/S FILL
XFILL_2_NAND2X1_215 BUFX2_43/A DFFSR_23/S FILL
XFILL_0_DFFSR_150 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_25_0_2 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_36_DFFSR_72 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_47_DFFSR_32 INVX1_2/gnd DFFSR_1/S FILL
XFILL_3_INVX1_124 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_6_NAND2X1_20 INVX1_23/gnd DFFSR_186/S FILL
XFILL_1_NAND3X1_113 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_31_DFFSR_184 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_20_DFFSR_22 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_0_OAI21X1_197 INVX1_8/gnd DFFSR_7/S FILL
XFILL_3_DFFSR_29 INVX1_4/gnd DFFSR_4/S FILL
XFILL_21_DFFSR_187 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_3_NAND2X1_149 DFFSR_89/gnd DFFSR_186/S FILL
XNAND2X1_20 DFFSR_91/S DFFSR_12/Q INVX1_23/gnd OAI21X1_20/C DFFSR_186/S NAND2X1
XFILL_5_1_2 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_5_NAND2X1_23 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_11_DFFSR_190 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_4_NAND2X1_26 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_11_OAI22X1_67 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_1_INVX1_341 DFFSR_3/gnd DFFSR_65/S FILL
XDFFPOSX1_23 AND2X2_9/A CLKBUF1_14/Y XOR2X1_12/Y INVX1_23/gnd DFFSR_91/S DFFPOSX1
XFILL_44_DFFSR_108 INVX1_89/gnd DFFSR_2/S FILL
XFILL_9_DFFSR_4 INVX1_4/gnd DFFSR_4/S FILL
XFILL_3_NAND2X1_29 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_4_OAI21X1_11 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_3_OAI21X1_14 BUFX2_43/A DFFSR_23/S FILL
XFILL_44_DFFSR_79 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_34_DFFSR_111 INVX1_8/gnd DFFSR_5/S FILL
XFILL_7_DFFSR_184 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_1_OAI21X1_131 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_2_NAND2X1_32 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_9_NAND3X1_88 INVX1_94/gnd DFFSR_52/S FILL
XFILL_2_OAI21X1_17 INVX1_8/gnd DFFSR_5/S FILL
XFILL_1_NAND2X1_35 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_1_OAI21X1_20 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_0_INVX1_23 INVX1_23/gnd DFFSR_91/S FILL
XFILL_8_NAND3X1_91 BUFX2_43/A DFFSR_97/S FILL
XFILL_17_DFFSR_69 BUFX2_43/A DFFSR_23/S FILL
XFILL_0_DFFSR_76 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_0_INVX1_161 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_24_DFFSR_114 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_0_NAND2X1_38 DFFSR_5/gnd DFFSR_5/S FILL
XINVX1_271 DFFSR_57/Q DFFSR_73/gnd OAI22X1_8/A DFFSR_57/S INVX1
XFILL_28_DFFSR_29 INVX1_4/gnd DFFSR_4/S FILL
XFILL_14_DFFSR_117 INVX1_23/gnd DFFSR_91/S FILL
XFILL_7_NAND3X1_94 BUFX2_35/A DFFSR_97/S FILL
XFILL_0_OAI21X1_23 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_1_NAND2X1_245 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_6_NAND3X1_97 BUFX2_35/A DFFSR_97/S FILL
XFILL_4_INVX1_268 INVX1_8/gnd DFFSR_7/S FILL
XFILL_4_XOR2X1_6 DFFSR_89/gnd DFFSR_186/S FILL
XNAND3X1_97 XOR2X1_7/Y NAND3X1_97/B NAND3X1_97/C BUFX2_35/A NAND3X1_98/B DFFSR_97/S
+ NAND3X1
XFILL_33_DFFSR_8 BUFX2_36/A DFFSR_8/S FILL
XFILL_5_DFFPOSX1_17 BUFX2_37/A DFFSR_8/S FILL
XFILL_7_OAI22X1_4 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_51_DFFSR_142 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_2_NAND2X1_179 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_0_DFFSR_114 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_41_DFFSR_145 INVX1_23/gnd DFFSR_186/S FILL
XFILL_25_DFFSR_76 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_8_DFFSR_83 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_36_DFFSR_36 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_30_1 INVX1_89/gnd DFFSR_2/S FILL
XFILL_31_DFFSR_148 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_21_DFFSR_151 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_0_OAI21X1_161 INVX1_23/gnd DFFSR_186/S FILL
XFILL_3_NAND2X1_113 INVX1_23/gnd DFFSR_91/S FILL
XFILL_11_DFFSR_154 BUFX2_36/A DFFSR_6/S FILL
XFILL_2_AOI22X1_10 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_1_INVX1_305 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_6_NOR2X1_30 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_1_AOI22X1_13 INVX1_23/gnd DFFSR_186/S FILL
XFILL_33_DFFSR_83 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_44_DFFSR_43 INVX1_94/gnd DFFSR_25/S FILL
XFILL_0_NAND2X1_275 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_10_OAI22X1_34 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_7_DFFSR_148 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_24_DFFPOSX1_25 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_48_DFFSR_179 INVX1_2/gnd DFFSR_1/S FILL
XFILL_8_NAND3X1_55 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_9_OAI22X1_37 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_8_OAI22X1_40 BUFX2_37/A DFFSR_8/S FILL
XFILL_7_NAND3X1_58 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_17_DFFSR_33 INVX1_94/gnd DFFSR_52/S FILL
XFILL_38_DFFSR_182 INVX1_89/gnd DFFSR_36/S FILL
XFILL_0_DFFSR_40 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_0_INVX1_125 DFFSR_5/gnd DFFSR_5/S FILL
XINVX1_235 INVX1_235/A INVX1_4/gnd INVX1_235/Y DFFSR_51/S INVX1
XFILL_28_DFFSR_185 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_4_INVX1_232 BUFX2_37/A DFFSR_8/S FILL
XFILL_7_OAI22X1_43 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_1_NAND2X1_209 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_6_NAND3X1_61 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_5_NAND3X1_64 BUFX2_35/A DFFSR_14/S FILL
XFILL_6_OAI22X1_46 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_18_DFFSR_188 INVX1_2/gnd DFFSR_1/S FILL
XFILL_4_NAND3X1_67 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_0_NAND3X1_107 BUFX2_43/A DFFSR_97/S FILL
XFILL_5_OAI22X1_49 INVX1_94/gnd DFFSR_25/S FILL
XNAND3X1_61 NAND3X1_2/A NAND3X1_60/Y NAND3X1_61/C DFFSR_79/gnd NAND3X1_61/Y DFFSR_45/S
+ NAND3X1
XFILL_10_XOR2X1_3 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_3_NAND3X1_70 BUFX2_35/A DFFSR_14/S FILL
XOAI22X1_46 INVX1_350/Y OAI22X1_38/B INVX1_351/Y OAI22X1_38/D BUFX2_19/gnd NOR2X1_32/A
+ DFFSR_52/S OAI22X1
XFILL_41_DFFSR_90 INVX1_2/gnd DFFSR_1/S FILL
XFILL_41_DFFSR_109 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_4_OAI22X1_52 INVX1_94/gnd DFFSR_25/S FILL
XFILL_2_NAND2X1_143 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_8_OAI21X1_246 DFFSR_9/gnd DFFSR_9/S FILL
XDFFSR_188 BUFX2_30/A DFFSR_1/CLK DFFSR_185/R DFFSR_1/S DFFSR_188/D INVX1_2/gnd DFFSR_1/S
+ DFFSR
XFILL_4_DFFSR_185 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_2_NAND3X1_73 BUFX2_43/A DFFSR_23/S FILL
XFILL_3_OAI22X1_55 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_8_DFFSR_47 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_25_DFFSR_40 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_14_DFFSR_80 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_1_NAND3X1_76 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_2_OAI22X1_58 BUFX2_17/gnd DFFSR_7/S FILL
XNAND2X1_9 INVX1_2/A DFFSR_1/S DFFSR_1/gnd NAND2X1_9/Y DFFSR_1/S NAND2X1
XFILL_31_DFFSR_112 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_21_DFFSR_115 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_0_OAI21X1_125 BUFX2_35/A DFFSR_14/S FILL
XFILL_0_NAND3X1_79 BUFX2_36/A DFFSR_6/S FILL
XFILL_1_OAI22X1_61 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_4_NAND2X1_6 INVX1_23/gnd DFFSR_186/S FILL
XFILL_0_OAI22X1_64 INVX1_94/gnd DFFSR_25/S FILL
XFILL_26_1_0 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_11_DFFSR_118 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_49_DFFSR_97 BUFX2_35/A DFFSR_97/S FILL
XFILL_20_DFFSR_2 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_1_INVX1_269 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_24_3_1 DFFSR_71/gnd DFFSR_10/S FILL
XOAI22X1_8 OAI22X1_8/A OAI22X1_8/B OAI22X1_8/C OAI22X1_8/D DFFSR_73/gnd NOR2X1_13/A
+ DFFSR_57/S OAI22X1
XFILL_6_2_0 BUFX2_35/A DFFSR_14/S FILL
XFILL_0_NAND2X1_239 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_33_DFFSR_47 DFFSR_5/gnd DFFSR_2/S FILL
XINVX1_81 INVX1_81/A DFFSR_5/gnd INVX1_81/Y DFFSR_2/S INVX1
XFILL_22_DFFSR_87 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_7_DFFSR_112 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_5_DFFSR_94 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_22_5_2 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_48_DFFSR_143 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_4_OAI22X1_5 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_38_DFFSR_146 DFFSR_89/gnd DFFSR_92/S FILL
XINVX1_199 DFFSR_165/Q BUFX2_35/A INVX1_199/Y DFFSR_97/S INVX1
XFILL_4_BUFX2_3 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_8_NAND3X1_19 INVX1_8/gnd DFFSR_5/S FILL
XFILL_28_DFFSR_149 INVX1_23/gnd DFFSR_91/S FILL
XFILL_4_4_1 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_1_NAND2X1_173 BUFX2_35/A DFFSR_14/S FILL
XFILL_7_NAND3X1_22 BUFX2_37/A DFFSR_81/S FILL
XFILL_35_6 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_4_BUFX2_32 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_4_DFFPOSX1_11 INVX1_4/gnd DFFSR_4/S FILL
XFILL_4_INVX1_196 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_18_DFFSR_152 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_6_NAND3X1_25 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_5_NAND3X1_28 BUFX2_7/gnd DFFSR_81/S FILL
XNAND3X1_25 AOI22X1_5/D NAND3X1_22/B NAND3X1_22/C BUFX2_7/gnd AOI21X1_4/B DFFSR_81/S
+ NAND3X1
XFILL_6_OAI22X1_10 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_41_DFFSR_54 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_4_NAND3X1_31 INVX1_94/gnd DFFSR_52/S FILL
XFILL_2_INVX1_88 INVX1_2/gnd DFFSR_1/S FILL
XFILL_5_OAI22X1_13 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_30_DFFSR_94 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_3_NOR2X1_31 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_13_DFFPOSX1_30 BUFX2_43/A DFFSR_97/S FILL
XDFFSR_152 DFFSR_152/Q CLKBUF1_11/Y DFFSR_152/R DFFSR_23/S DFFSR_152/D BUFX2_5/gnd
+ DFFSR_23/S DFFSR
XFILL_2_NAND2X1_107 BUFX2_36/A DFFSR_6/S FILL
XFILL_8_OAI21X1_210 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_3_NAND3X1_34 INVX1_2/gnd DFFSR_1/S FILL
XFILL_4_OAI22X1_16 INVX1_4/gnd DFFSR_4/S FILL
XOAI22X1_10 INVX1_275/Y OAI22X1_8/D INVX1_276/Y OAI22X1_6/D DFFSR_3/gnd NOR2X1_14/A
+ DFFSR_4/S OAI22X1
XFILL_2_INVX1_413 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_2_NAND3X1_37 BUFX2_43/A DFFSR_97/S FILL
XFILL_14_DFFSR_44 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_3_OAI22X1_19 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_8_DFFSR_11 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_4_DFFSR_149 INVX1_23/gnd DFFSR_91/S FILL
XFILL_1_NAND3X1_40 BUFX2_43/A DFFSR_23/S FILL
XFILL_45_DFFSR_180 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_2_OAI22X1_22 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_0_NAND3X1_43 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_1_OAI22X1_25 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_35_DFFSR_183 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_0_OAI22X1_28 INVX1_94/gnd DFFSR_25/S FILL
XFILL_23_DFFPOSX1_19 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_25_DFFSR_186 INVX1_23/gnd DFFSR_186/S FILL
XFILL_49_DFFSR_61 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_1_INVX1_233 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_15_DFFSR_189 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_0_NAND2X1_203 BUFX2_5/gnd DFFSR_23/S FILL
XINVX1_45 DFFSR_40/Q INVX1_8/gnd INVX1_45/Y DFFSR_5/S INVX1
XFILL_32_0_2 INVX1_8/gnd DFFSR_5/S FILL
XDFFSR_98 DFFSR_98/Q CLKBUF1_2/Y DFFSR_97/R DFFSR_9/S DFFSR_98/D DFFSR_9/gnd DFFSR_9/S
+ DFFSR
XFILL_5_DFFSR_58 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_33_DFFSR_11 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_11_DFFSR_91 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_48_DFFSR_107 BUFX2_36/A DFFSR_8/S FILL
XFILL_22_DFFSR_51 INVX1_2/gnd DFFSR_51/S FILL
XFILL_38_DFFSR_110 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_1_DFFSR_186 INVX1_23/gnd DFFSR_186/S FILL
XINVX1_163 BUFX2_10/Y INVX1_94/gnd DFFSR_137/R DFFSR_52/S INVX1
XFILL_28_DFFSR_113 INVX1_23/gnd DFFSR_186/S FILL
XFILL_4_INVX1_160 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_1_NAND2X1_137 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_7_OAI21X1_240 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_18_DFFSR_116 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_1_NAND2X1_7 INVX1_89/gnd DFFSR_36/S FILL
XFILL_2_INVX1_52 BUFX2_37/A DFFSR_81/S FILL
XFILL_19_DFFSR_98 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_41_DFFSR_18 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_30_DFFSR_58 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_8_OAI21X1_174 BUFX2_43/A DFFSR_23/S FILL
XDFFSR_116 INVX1_131/A CLKBUF1_1/Y DFFSR_113/R DFFSR_2/S DFFSR_116/D DFFSR_5/gnd DFFSR_2/S
+ DFFSR
XFILL_2_INVX1_377 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_4_DFFSR_113 INVX1_23/gnd DFFSR_186/S FILL
XFILL_1_BUFX2_43 BUFX2_35/A DFFSR_97/S FILL
XFILL_45_DFFSR_144 INVX1_8/gnd DFFSR_5/S FILL
XFILL_1_OAI22X1_6 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_35_DFFSR_147 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_8_DFFSR_1 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_25_DFFSR_150 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_11_DFFSR_9 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_15_DFFSR_153 BUFX2_36/A DFFSR_8/S FILL
XFILL_49_DFFSR_25 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_1_INVX1_197 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_38_DFFSR_65 DFFSR_3/gnd DFFSR_65/S FILL
XDFFSR_62 INVX1_70/A DFFSR_28/CLK DFFSR_61/R DFFSR_52/S DFFSR_62/D BUFX2_19/gnd DFFSR_52/S
+ DFFSR
XFILL_0_NOR2X1_32 INVX1_94/gnd DFFSR_52/S FILL
XFILL_5_DFFSR_22 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_11_DFFSR_55 INVX1_89/gnd DFFSR_36/S FILL
XFILL_22_DFFSR_15 INVX1_8/gnd DFFSR_7/S FILL
XFILL_0_NAND2X1_167 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_6_OR2X2_1 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_8_NAND3X1_120 DFFSR_5/gnd DFFSR_5/S FILL
XINVX1_127 BUFX2_8/Y INVX1_2/gnd DFFSR_105/R DFFSR_1/S INVX1
XFILL_12_DFFPOSX1_24 BUFX2_43/A DFFSR_23/S FILL
XFILL_4_NOR2X1_3 INVX1_94/gnd DFFSR_25/S FILL
XFILL_1_DFFSR_150 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_32_DFFSR_5 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_1_NAND2X1_101 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_42_DFFSR_181 INVX1_23/gnd DFFSR_186/S FILL
XFILL_7_OAI21X1_204 BUFX2_36/A DFFSR_6/S FILL
XFILL_46_DFFSR_72 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_4_INVX1_124 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_32_DFFSR_184 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_2_INVX1_16 BUFX2_43/A DFFSR_23/S FILL
XFILL_2_DFFSR_69 BUFX2_43/A DFFSR_23/S FILL
XFILL_19_DFFSR_62 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_30_DFFSR_22 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_22_DFFSR_187 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_22_DFFPOSX1_13 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_12_DFFSR_190 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_8_OAI21X1_138 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_2_INVX1_341 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_45_DFFSR_108 INVX1_89/gnd DFFSR_2/S FILL
XFILL_8_DFFSR_184 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_35_DFFSR_111 INVX1_8/gnd DFFSR_5/S FILL
XFILL_27_DFFSR_69 BUFX2_43/A DFFSR_23/S FILL
XFILL_1_INVX1_161 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_25_DFFSR_114 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_38_DFFSR_29 INVX1_4/gnd DFFSR_4/S FILL
XFILL_15_DFFSR_117 INVX1_23/gnd DFFSR_91/S FILL
XFILL_6_OAI21X1_234 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_0_NAND2X1_131 DFFSR_9/gnd DFFSR_9/S FILL
XDFFSR_26 INVX1_30/A DFFSR_24/CLK DFFSR_31/R DFFSR_9/S DFFSR_26/D DFFSR_9/gnd DFFSR_9/S
+ DFFSR
XFILL_11_DFFSR_19 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_17_3 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_8_OAI22X1_4 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_1_DFFSR_114 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_42_DFFSR_145 INVX1_23/gnd DFFSR_186/S FILL
XFILL_7_OAI21X1_168 BUFX2_36/A DFFSR_6/S FILL
XFILL_35_DFFSR_76 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_46_DFFSR_36 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_33_1_0 INVX1_8/gnd DFFSR_7/S FILL
XFILL_32_DFFSR_148 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_22_DFFSR_151 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_31_3_1 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_12_DFFSR_154 BUFX2_36/A DFFSR_6/S FILL
XFILL_2_DFFSR_33 INVX1_94/gnd DFFSR_52/S FILL
XFILL_19_DFFSR_26 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_2_INVX1_305 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_8_OAI21X1_102 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_20_CLKBUF1_16 BUFX2_36/A DFFSR_6/S FILL
XFILL_29_5_2 INVX1_89/gnd DFFSR_2/S FILL
XFILL_19_CLKBUF1_19 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_8_DFFSR_148 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_43_DFFSR_83 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_18_CLKBUF1_22 INVX1_94/gnd DFFSR_25/S FILL
XFILL_5_OAI21X1_264 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_49_DFFSR_179 INVX1_2/gnd DFFSR_1/S FILL
XFILL_17_CLKBUF1_25 INVX1_23/gnd DFFSR_186/S FILL
XFILL_27_DFFSR_33 INVX1_94/gnd DFFSR_52/S FILL
XFILL_7_NAND3X1_114 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_39_DFFSR_182 INVX1_89/gnd DFFSR_36/S FILL
XFILL_1_INVX1_125 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_16_DFFSR_73 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_29_DFFSR_185 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_11_DFFPOSX1_18 BUFX2_37/A DFFSR_8/S FILL
XFILL_6_OAI21X1_198 INVX1_8/gnd DFFSR_7/S FILL
XFILL_19_DFFSR_188 INVX1_2/gnd DFFSR_1/S FILL
XOAI21X1_234 AOI21X1_30/Y AOI21X1_31/Y INVX1_260/A BUFX2_6/gnd AOI21X1_32/B DFFSR_91/S
+ OAI21X1
XFILL_42_DFFSR_109 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_5_DFFSR_185 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_35_DFFSR_40 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_7_OAI21X1_132 INVX1_4/gnd DFFSR_4/S FILL
XFILL_7_DFFSR_87 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_24_DFFSR_80 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_32_DFFSR_112 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_22_DFFSR_115 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_1_DFFPOSX1_29 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_39_0_2 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_5_NAND2X1_6 INVX1_23/gnd DFFSR_186/S FILL
XFILL_6_BUFX2_25 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_12_DFFSR_118 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_2_INVX1_269 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_44_DFFSR_8 BUFX2_36/A DFFSR_8/S FILL
XFILL_5_OAI21X1_228 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_43_DFFSR_47 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_4_INVX1_81 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_32_DFFSR_87 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_8_DFFSR_112 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_49_DFFSR_143 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_5_OAI22X1_5 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_39_DFFSR_146 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_22_8 INVX1_94/gnd DFFSR_25/S FILL
XFILL_16_DFFSR_37 INVX1_89/gnd DFFSR_2/S FILL
XFILL_29_DFFSR_149 INVX1_23/gnd DFFSR_91/S FILL
XFILL_39_3 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_6_OAI21X1_162 INVX1_23/gnd DFFSR_91/S FILL
XFILL_19_DFFSR_152 BUFX2_5/gnd DFFSR_23/S FILL
XNOR2X1_34 NOR2X1_34/A NOR2X1_34/B DFFSR_71/gnd NOR2X1_34/Y DFFSR_10/S NOR2X1
XFILL_40_DFFSR_94 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_4_NOR2X1_31 DFFSR_73/gnd DFFSR_11/S FILL
XOAI21X1_198 AOI21X1_13/Y INVX1_237/Y AOI21X1_12/Y INVX1_8/gnd NAND3X1_34/C DFFSR_7/S
+ OAI21X1
XFILL_3_INVX1_413 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_24_DFFSR_44 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_6_NAND2X1_276 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_1_AND2X2_3 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_7_DFFSR_51 INVX1_2/gnd DFFSR_51/S FILL
XFILL_5_DFFSR_149 INVX1_23/gnd DFFSR_91/S FILL
XFILL_13_DFFSR_84 BUFX2_43/A DFFSR_23/S FILL
XFILL_46_DFFSR_180 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_10_CLKBUF1_10 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_36_DFFSR_183 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_4_OAI21X1_258 INVX1_2/gnd DFFSR_51/S FILL
XFILL_26_DFFSR_186 INVX1_23/gnd DFFSR_186/S FILL
XFILL_2_INVX1_233 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_9_CLKBUF1_13 INVX1_4/gnd DFFSR_51/S FILL
XFILL_10_DFFSR_6 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_8_CLKBUF1_16 BUFX2_36/A DFFSR_6/S FILL
XFILL_6_NAND3X1_108 BUFX2_37/A DFFSR_81/S FILL
XFILL_16_DFFSR_189 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_10_DFFPOSX1_12 INVX1_8/gnd DFFSR_5/S FILL
XFILL_7_CLKBUF1_19 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_21_DFFSR_91 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_49_DFFSR_107 BUFX2_36/A DFFSR_8/S FILL
XFILL_5_OAI21X1_192 BUFX2_37/A DFFSR_81/S FILL
XFILL_6_CLKBUF1_22 INVX1_94/gnd DFFSR_25/S FILL
XFILL_4_DFFSR_98 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_32_DFFSR_51 INVX1_2/gnd DFFSR_51/S FILL
XFILL_43_DFFSR_11 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_5_CLKBUF1_25 INVX1_23/gnd DFFSR_186/S FILL
XFILL_2_DFFSR_186 INVX1_23/gnd DFFSR_186/S FILL
XOR2X2_2 OR2X2_2/A OR2X2_2/B BUFX2_6/gnd OR2X2_2/Y DFFSR_91/S OR2X2
XFILL_3_BUFX2_36 BUFX2_5/gnd DFFSR_23/S FILL
XCLKBUF1_22 INVX1_402/Y INVX1_94/gnd DFFSR_28/CLK DFFSR_25/S CLKBUF1
XFILL_39_DFFSR_110 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_29_DFFSR_113 INVX1_23/gnd DFFSR_186/S FILL
XFILL_19_DFFSR_116 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_6_OAI21X1_126 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_2_NAND2X1_7 INVX1_89/gnd DFFSR_36/S FILL
XFILL_31_DFFSR_2 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_0_DFFPOSX1_23 INVX1_23/gnd DFFSR_91/S FILL
XFILL_1_INVX1_92 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_29_DFFSR_98 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_40_DFFSR_58 DFFSR_3/gnd DFFSR_4/S FILL
XOAI21X1_162 BUFX2_2/Y INVX1_196/Y OAI21X1_162/C INVX1_23/gnd DFFSR_162/D DFFSR_91/S
+ OAI21X1
XFILL_6_NAND2X1_240 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_3_INVX1_377 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_5_DFFSR_113 INVX1_23/gnd DFFSR_186/S FILL
XFILL_7_DFFSR_15 INVX1_8/gnd DFFSR_7/S FILL
XFILL_13_DFFSR_48 INVX1_4/gnd DFFSR_4/S FILL
XFILL_46_DFFSR_144 INVX1_8/gnd DFFSR_5/S FILL
XFILL_2_OAI22X1_6 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_36_DFFSR_147 DFFSR_89/gnd DFFSR_186/S FILL
XNAND2X1_276 INVX1_427/Y INVX1_428/Y DFFSR_71/gnd AND2X2_16/A DFFSR_10/S NAND2X1
XFILL_4_OAI21X1_222 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_26_DFFSR_150 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_16_DFFSR_153 BUFX2_36/A DFFSR_8/S FILL
XFILL_2_INVX1_197 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_48_DFFSR_65 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_5_OAI21X1_156 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_4_DFFSR_62 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_1_NOR2X1_32 INVX1_94/gnd DFFSR_52/S FILL
XFILL_10_DFFSR_95 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_21_DFFSR_55 INVX1_89/gnd DFFSR_36/S FILL
XFILL_32_DFFSR_15 INVX1_8/gnd DFFSR_7/S FILL
XFILL_19_DFFPOSX1_31 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_40_1_0 DFFSR_3/gnd DFFSR_65/S FILL
XNAND3X1_108 INVX1_251/Y AOI21X1_39/B AOI21X1_39/A BUFX2_37/A NAND2X1_231/B DFFSR_81/S
+ NAND3X1
XFILL_0_INVX1_414 INVX1_2/gnd DFFSR_1/S FILL
XFILL_38_3_1 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_2_DFFSR_150 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_43_DFFSR_181 INVX1_23/gnd DFFSR_186/S FILL
XFILL_5_NAND2X1_270 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_36_5_2 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_33_DFFSR_184 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_29_DFFSR_62 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_40_DFFSR_22 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_23_DFFSR_187 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_1_INVX1_56 DFFSR_73/gnd DFFSR_11/S FILL
XOAI21X1_126 BUFX2_16/Y INVX1_142/Y OAI21X1_126/C BUFX2_17/gnd DFFSR_126/D DFFSR_7/S
+ OAI21X1
XFILL_3_OAI21X1_252 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_13_DFFSR_190 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_6_NAND2X1_204 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_3_INVX1_341 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_13_DFFSR_12 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_46_DFFSR_108 INVX1_89/gnd DFFSR_2/S FILL
XFILL_5_NAND3X1_102 INVX1_23/gnd DFFSR_186/S FILL
XFILL_9_DFFSR_184 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_4_OAI21X1_186 BUFX2_36/A DFFSR_8/S FILL
XNAND2X1_240 NOR2X1_25/Y NOR2X1_24/Y BUFX2_8/gnd NAND2X1_71/B DFFSR_10/S NAND2X1
XFILL_36_DFFSR_111 INVX1_8/gnd DFFSR_5/S FILL
XFILL_37_DFFSR_69 BUFX2_43/A DFFSR_23/S FILL
XFILL_2_INVX1_161 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_26_DFFSR_114 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_48_DFFSR_29 INVX1_4/gnd DFFSR_4/S FILL
XFILL_16_DFFSR_117 INVX1_23/gnd DFFSR_91/S FILL
XFILL_4_DFFSR_26 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_21_DFFSR_19 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_10_DFFSR_59 INVX1_4/gnd DFFSR_51/S FILL
XFILL_5_OAI21X1_120 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_0_INVX1_378 INVX1_8/gnd DFFSR_7/S FILL
XFILL_3_NOR2X1_7 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_9_OAI22X1_4 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_2_DFFSR_114 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_43_DFFSR_145 INVX1_23/gnd DFFSR_186/S FILL
XFILL_45_DFFSR_76 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_46_0_2 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_22_DFFSR_9 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_5_NAND2X1_234 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_33_DFFSR_148 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_23_DFFSR_151 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_4_NAND3X1_132 INVX1_8/gnd DFFSR_7/S FILL
XFILL_13_DFFSR_154 BUFX2_36/A DFFSR_6/S FILL
XFILL_1_INVX1_20 INVX1_8/gnd DFFSR_5/S FILL
XFILL_29_DFFSR_26 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_18_DFFSR_66 INVX1_2/gnd DFFSR_51/S FILL
XFILL_1_DFFSR_73 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_3_OAI21X1_216 BUFX2_35/A DFFSR_14/S FILL
XFILL_6_NAND2X1_168 BUFX2_36/A DFFSR_6/S FILL
XFILL_3_INVX1_305 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_21_DFFPOSX1_1 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_0_BUFX2_11 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_5_XOR2X1_3 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_9_DFFSR_148 DFFSR_89/gnd DFFSR_92/S FILL
XNAND2X1_204 AND2X2_6/A AND2X2_6/B BUFX2_5/gnd NOR2X1_8/A DFFSR_6/S NAND2X1
XFILL_18_DFFPOSX1_25 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_43_DFFSR_5 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_20_DFFPOSX1_4 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_12_1_1 BUFX2_36/A DFFSR_6/S FILL
XFILL_4_OAI21X1_150 INVX1_94/gnd DFFSR_52/S FILL
XFILL_19_DFFPOSX1_7 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_50_DFFSR_179 INVX1_2/gnd DFFSR_1/S FILL
XFILL_37_DFFSR_33 INVX1_94/gnd DFFSR_52/S FILL
XFILL_40_DFFSR_182 INVX1_89/gnd DFFSR_36/S FILL
XFILL_2_INVX1_125 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_9_DFFSR_80 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_26_DFFSR_73 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_30_DFFSR_185 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_4_NAND2X1_264 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_10_3_2 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_10_DFFSR_23 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_20_DFFSR_188 INVX1_2/gnd DFFSR_1/S FILL
XFILL_10_DFFSR_191 INVX1_23/gnd DFFSR_91/S FILL
XFILL_0_INVX1_342 INVX1_8/gnd DFFSR_7/S FILL
XFILL_4_4 INVX1_23/gnd DFFSR_91/S FILL
XFILL_6_DFFSR_185 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_43_DFFSR_109 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_45_DFFSR_40 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_5_NAND2X1_198 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_2_OAI21X1_246 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_34_DFFSR_80 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_33_DFFSR_112 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_23_DFFSR_115 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_18_DFFSR_30 INVX1_89/gnd DFFSR_36/S FILL
XFILL_1_DFFSR_37 INVX1_89/gnd DFFSR_2/S FILL
XFILL_6_NAND2X1_6 INVX1_23/gnd DFFSR_186/S FILL
XFILL_3_OAI21X1_180 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_13_DFFSR_118 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_3_INVX1_269 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_6_NAND2X1_132 INVX1_8/gnd DFFSR_5/S FILL
XXOR2X1_7 XOR2X1_7/A XOR2X1_7/B INVX1_23/gnd XOR2X1_7/Y DFFSR_91/S XOR2X1
XNAND2X1_168 NAND2X1_168/A DFFSR_6/S BUFX2_36/A NAND2X1_168/Y DFFSR_6/S NAND2X1
XFILL_42_DFFSR_87 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_9_DFFSR_112 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_50_DFFSR_143 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_4_OAI21X1_114 INVX1_89/gnd DFFSR_36/S FILL
XFILL_6_OAI22X1_5 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_40_DFFSR_146 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_9_DFFSR_44 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_26_5 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_26_DFFSR_37 INVX1_89/gnd DFFSR_2/S FILL
XFILL_30_DFFSR_149 INVX1_23/gnd DFFSR_91/S FILL
XFILL_15_DFFSR_77 INVX1_89/gnd DFFSR_2/S FILL
XFILL_20_DFFSR_152 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_4_NAND2X1_228 INVX1_23/gnd DFFSR_91/S FILL
XFILL_10_DFFSR_155 BUFX2_7/gnd DFFSR_54/S FILL
XINVX1_416 BUFX2_27/A DFFSR_89/gnd INVX1_416/Y DFFSR_92/S INVX1
XFILL_0_INVX1_306 INVX1_94/gnd DFFSR_25/S FILL
XFILL_3_NAND3X1_126 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_50_DFFSR_94 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_5_NOR2X1_31 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_6_DFFSR_91 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_5_NAND2X1_162 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_2_OAI21X1_210 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_6_DFFSR_149 INVX1_23/gnd DFFSR_91/S FILL
XFILL_23_DFFSR_84 BUFX2_43/A DFFSR_23/S FILL
XFILL_34_DFFSR_44 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_47_DFFSR_180 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_37_DFFSR_183 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_47_1_0 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_5_BUFX2_29 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_27_DFFSR_186 INVX1_23/gnd DFFSR_186/S FILL
XFILL_3_INVX1_233 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_3_OAI21X1_144 INVX1_8/gnd DFFSR_7/S FILL
XFILL_17_DFFPOSX1_19 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_17_DFFSR_189 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_9_DFFPOSX1_1 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_45_3_1 INVX1_2/gnd DFFSR_1/S FILL
XFILL_31_DFFSR_91 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_9_AOI21X1_21 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_50_DFFSR_107 BUFX2_36/A DFFSR_8/S FILL
XNAND2X1_132 DFFSR_7/S NAND2X1_68/B INVX1_8/gnd NAND2X1_132/Y DFFSR_5/S NAND2X1
XFILL_8_DFFPOSX1_4 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_3_NAND2X1_258 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_42_DFFSR_51 INVX1_2/gnd DFFSR_51/S FILL
XFILL_3_INVX1_85 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_8_AOI21X1_24 BUFX2_43/A DFFSR_97/S FILL
XFILL_7_DFFPOSX1_7 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_43_5_2 INVX1_4/gnd DFFSR_51/S FILL
XFILL_3_DFFSR_186 INVX1_23/gnd DFFSR_186/S FILL
XFILL_7_AOI21X1_27 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_15_DFFSR_41 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_40_DFFSR_110 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_30_DFFSR_113 INVX1_23/gnd DFFSR_186/S FILL
XFILL_6_AOI21X1_30 INVX1_23/gnd DFFSR_91/S FILL
XFILL_5_AOI21X1_33 BUFX2_35/A DFFSR_14/S FILL
XFILL_7_DFFPOSX1_30 BUFX2_43/A DFFSR_97/S FILL
XFILL_4_NAND2X1_192 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_20_DFFSR_116 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_1_OAI21X1_240 DFFSR_5/gnd DFFSR_5/S FILL
XAOI21X1_30 AOI21X1_30/A AOI21X1_30/B INVX1_254/Y INVX1_23/gnd AOI21X1_30/Y DFFSR_91/S
+ AOI21X1
XFILL_10_DFFSR_119 BUFX2_37/A DFFSR_81/S FILL
XFILL_4_AOI21X1_36 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_3_NAND2X1_7 INVX1_89/gnd DFFSR_36/S FILL
XFILL_3_AOI21X1_39 BUFX2_7/gnd DFFSR_81/S FILL
XINVX1_380 INVX1_80/A DFFSR_79/gnd INVX1_380/Y DFFSR_45/S INVX1
XFILL_0_INVX1_270 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_39_DFFSR_98 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_50_DFFSR_58 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_2_AOI21X1_42 INVX1_23/gnd DFFSR_91/S FILL
XFILL_2_OAI21X1_174 BUFX2_43/A DFFSR_23/S FILL
XFILL_11_4_0 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_6_DFFSR_113 INVX1_23/gnd DFFSR_186/S FILL
XFILL_0_AND2X2_7 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_6_DFFSR_55 INVX1_89/gnd DFFSR_36/S FILL
XFILL_1_AOI21X1_45 INVX1_89/gnd DFFSR_36/S FILL
XFILL_5_NAND2X1_126 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_23_DFFSR_48 INVX1_4/gnd DFFSR_4/S FILL
XFILL_12_DFFSR_88 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_0_AOI21X1_48 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_47_DFFSR_144 INVX1_8/gnd DFFSR_5/S FILL
XFILL_3_OAI22X1_6 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_37_DFFSR_147 DFFSR_89/gnd DFFSR_186/S FILL
XBUFX2_33 BUFX2_33/A DFFSR_89/gnd dout[7] DFFSR_186/S BUFX2
XFILL_27_DFFSR_150 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_3_OAI21X1_108 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_17_DFFSR_153 BUFX2_36/A DFFSR_8/S FILL
XFILL_48_5 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_3_INVX1_197 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_8_OAI21X1_72 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_2_NOR2X1_32 INVX1_94/gnd DFFSR_52/S FILL
XFILL_3_INVX1_49 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_20_DFFSR_95 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_31_DFFSR_55 INVX1_89/gnd DFFSR_36/S FILL
XFILL_42_DFFSR_15 INVX1_8/gnd DFFSR_7/S FILL
XFILL_7_OAI21X1_75 INVX1_4/gnd DFFSR_4/S FILL
XFILL_6_NAND2X1_93 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_3_NAND2X1_222 INVX1_23/gnd DFFSR_186/S FILL
XFILL_6_OAI21X1_78 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_5_NAND2X1_96 INVX1_4/gnd DFFSR_51/S FILL
XNAND2X1_93 BUFX2_18/Y DFFSR_85/Q DFFSR_3/gnd NAND2X1_93/Y DFFSR_65/S NAND2X1
XFILL_4_NAND2X1_99 BUFX2_43/A DFFSR_97/S FILL
XFILL_5_OAI21X1_81 BUFX2_19/gnd DFFSR_54/S FILL
XOAI21X1_78 BUFX2_18/Y INVX1_88/Y NAND2X1_78/Y DFFSR_1/gnd DFFSR_78/D DFFSR_1/S OAI21X1
XFILL_1_INVX1_414 INVX1_2/gnd DFFSR_1/S FILL
XFILL_2_BUFX2_40 BUFX2_35/A DFFSR_14/S FILL
XFILL_4_OAI21X1_84 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_3_DFFSR_150 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_2_NAND3X1_120 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_44_DFFSR_181 INVX1_23/gnd DFFSR_186/S FILL
XFILL_1_OAI21X1_204 BUFX2_36/A DFFSR_6/S FILL
XFILL_3_OAI21X1_87 INVX1_4/gnd DFFSR_4/S FILL
XFILL_21_DFFSR_6 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_4_NAND2X1_156 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_2_OAI21X1_90 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_34_DFFSR_184 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_39_DFFSR_62 BUFX2_19/gnd DFFSR_52/S FILL
XINVX1_344 INVX1_344/A BUFX2_8/gnd INVX1_344/Y DFFSR_25/S INVX1
XFILL_50_DFFSR_22 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_0_INVX1_96 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_0_INVX1_234 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_1_OAI21X1_93 INVX1_4/gnd DFFSR_51/S FILL
XFILL_24_DFFSR_187 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_14_DFFSR_190 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_0_OAI21X1_96 INVX1_4/gnd DFFSR_51/S FILL
XFILL_16_DFFPOSX1_13 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_6_DFFSR_19 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_2_OAI21X1_138 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_23_DFFSR_12 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_5_BUFX2_7 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_19_1_1 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_12_DFFSR_52 INVX1_94/gnd DFFSR_52/S FILL
XFILL_1_0_0 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_47_DFFSR_108 INVX1_89/gnd DFFSR_2/S FILL
XFILL_0_AOI21X1_12 INVX1_8/gnd DFFSR_7/S FILL
XFILL_17_3_2 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_2_NAND2X1_252 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_37_DFFSR_111 INVX1_8/gnd DFFSR_5/S FILL
XFILL_0_DFFSR_187 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_47_DFFSR_69 BUFX2_43/A DFFSR_23/S FILL
XFILL_9_OAI21X1_33 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_3_INVX1_161 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_27_DFFSR_114 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_42_DFFSR_2 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_17_DFFSR_117 INVX1_23/gnd DFFSR_91/S FILL
XFILL_8_OAI21X1_36 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_0_NAND2X1_8 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_7_OAI21X1_39 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_6_NAND2X1_57 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_0_OAI21X1_234 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_6_DFFPOSX1_24 BUFX2_43/A DFFSR_23/S FILL
XFILL_3_NAND2X1_186 BUFX2_37/A DFFSR_81/S FILL
XFILL_5_NAND2X1_60 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_31_DFFSR_19 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_3_DFFSR_66 INVX1_2/gnd DFFSR_51/S FILL
XFILL_20_DFFSR_59 INVX1_4/gnd DFFSR_51/S FILL
XFILL_6_OAI21X1_42 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_3_INVX1_13 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_4_NAND2X1_63 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_5_OAI21X1_45 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_1_INVX1_378 INVX1_8/gnd DFFSR_7/S FILL
XNAND2X1_57 DFFSR_49/Q DFFSR_17/S BUFX2_17/gnd NAND2X1_57/Y DFFSR_57/S NAND2X1
XFILL_3_DFFSR_114 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_3_NAND2X1_66 INVX1_4/gnd DFFSR_51/S FILL
XFILL_4_OAI21X1_48 DFFSR_3/gnd DFFSR_4/S FILL
XOAI21X1_42 DFFSR_11/S INVX1_48/Y OAI21X1_42/C BUFX2_16/gnd DFFSR_42/D DFFSR_65/S
+ OAI21X1
XFILL_44_DFFSR_145 INVX1_23/gnd DFFSR_186/S FILL
XFILL_2_NAND2X1_69 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_0_OAI22X1_7 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_3_OAI21X1_51 INVX1_2/gnd DFFSR_51/S FILL
XFILL_34_DFFSR_148 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_1_OAI21X1_168 BUFX2_36/A DFFSR_6/S FILL
XFILL_2_OAI21X1_54 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_1_NAND2X1_72 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_4_NAND2X1_120 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_24_DFFSR_151 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_14_DFFSR_154 BUFX2_36/A DFFSR_6/S FILL
XINVX1_308 DFFSR_46/Q BUFX2_7/gnd INVX1_308/Y DFFSR_54/S INVX1
XFILL_0_INVX1_60 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_0_INVX1_198 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_39_DFFSR_26 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_28_DFFSR_66 INVX1_2/gnd DFFSR_51/S FILL
XFILL_0_NAND2X1_75 INVX1_4/gnd DFFSR_4/S FILL
XFILL_1_OAI21X1_57 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_0_OAI21X1_60 BUFX2_37/A DFFSR_81/S FILL
XFILL_4_INVX1_305 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_1_NAND2X1_282 INVX1_89/gnd DFFSR_2/S FILL
XFILL_2_OAI21X1_102 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_12_DFFSR_16 DFFSR_71/gnd DFFSR_45/S FILL
XNOR2X1_4 NOR2X1_4/A NOR2X1_3/A BUFX2_8/gnd NOR2X1_4/Y DFFSR_10/S NOR2X1
XFILL_2_NAND2X1_216 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_0_DFFSR_151 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_51_DFFSR_179 INVX1_2/gnd DFFSR_1/S FILL
XFILL_47_DFFSR_33 INVX1_94/gnd DFFSR_52/S FILL
XFILL_41_DFFSR_182 INVX1_89/gnd DFFSR_36/S FILL
XFILL_3_INVX1_125 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_36_DFFSR_73 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_31_DFFSR_185 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_1_NAND3X1_114 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_20_DFFSR_23 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_3_DFFSR_30 INVX1_89/gnd DFFSR_36/S FILL
XFILL_0_OAI21X1_198 INVX1_8/gnd DFFSR_7/S FILL
XFILL_21_DFFSR_188 INVX1_2/gnd DFFSR_1/S FILL
XFILL_6_NAND2X1_21 INVX1_4/gnd DFFSR_4/S FILL
XFILL_11_DFFSR_191 INVX1_23/gnd DFFSR_91/S FILL
XFILL_3_NAND2X1_150 BUFX2_37/A DFFSR_81/S FILL
XFILL_5_NAND2X1_24 DFFSR_73/gnd DFFSR_57/S FILL
XNAND2X1_21 DFFSR_3/S DFFSR_13/Q INVX1_4/gnd NAND2X1_21/Y DFFSR_4/S NAND2X1
XFILL_8_1 BUFX2_35/A DFFSR_97/S FILL
XFILL_1_INVX1_342 INVX1_8/gnd DFFSR_7/S FILL
XFILL_4_NAND2X1_27 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_4_OAI21X1_12 BUFX2_35/A DFFSR_14/S FILL
XDFFPOSX1_24 AND2X2_5/B CLKBUF1_16/Y XNOR2X1_4/Y BUFX2_43/A DFFSR_23/S DFFPOSX1
XFILL_3_NAND2X1_30 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_9_DFFSR_5 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_11_OAI22X1_68 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_7_DFFSR_185 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_44_DFFSR_109 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_2_NAND2X1_33 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_3_OAI21X1_15 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_1_OAI21X1_132 INVX1_4/gnd DFFSR_4/S FILL
XFILL_44_DFFSR_80 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_1_NAND2X1_36 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_2_OAI21X1_18 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_34_DFFSR_112 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_24_DFFSR_115 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_8_NAND3X1_92 BUFX2_43/A DFFSR_23/S FILL
XFILL_0_NAND2X1_39 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_28_DFFSR_30 INVX1_89/gnd DFFSR_36/S FILL
XFILL_0_DFFSR_77 INVX1_89/gnd DFFSR_2/S FILL
XFILL_0_INVX1_162 INVX1_8/gnd DFFSR_7/S FILL
XFILL_17_DFFSR_70 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_0_INVX1_24 INVX1_2/gnd DFFSR_51/S FILL
XFILL_1_OAI21X1_21 INVX1_2/gnd DFFSR_51/S FILL
XINVX1_272 INVX1_47/A DFFSR_73/gnd OAI22X1_8/C DFFSR_11/S INVX1
XFILL_7_NAND3X1_95 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_14_DFFSR_118 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_0_OAI21X1_24 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_6_NAND3X1_98 BUFX2_35/A DFFSR_14/S FILL
XFILL_1_NAND2X1_246 INVX1_94/gnd DFFSR_25/S FILL
XFILL_4_INVX1_269 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_4_XOR2X1_7 INVX1_23/gnd DFFSR_91/S FILL
XNAND3X1_98 NOR2X1_11/Y NAND3X1_98/B NAND3X1_98/C BUFX2_35/A AOI21X1_30/B DFFSR_14/S
+ NAND3X1
XFILL_33_DFFSR_9 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_0_DFFSR_115 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_5_DFFPOSX1_18 BUFX2_37/A DFFSR_8/S FILL
XFILL_2_NAND2X1_180 INVX1_94/gnd DFFSR_52/S FILL
XFILL_7_OAI22X1_5 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_41_DFFSR_146 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_8_DFFSR_84 BUFX2_43/A DFFSR_23/S FILL
XFILL_30_2 INVX1_89/gnd DFFSR_2/S FILL
XFILL_36_DFFSR_37 INVX1_89/gnd DFFSR_2/S FILL
XFILL_31_DFFSR_149 INVX1_23/gnd DFFSR_91/S FILL
XFILL_25_DFFSR_77 INVX1_89/gnd DFFSR_2/S FILL
XFILL_21_DFFSR_152 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_0_OAI21X1_162 INVX1_23/gnd DFFSR_91/S FILL
XFILL_11_DFFSR_155 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_18_4_0 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_3_NAND2X1_114 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_2_AOI22X1_11 INVX1_23/gnd DFFSR_91/S FILL
XFILL_1_INVX1_306 INVX1_94/gnd DFFSR_25/S FILL
XFILL_6_NOR2X1_31 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_17_NOR3X1_1 INVX1_94/gnd DFFSR_52/S FILL
XFILL_1_AOI22X1_14 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_0_NAND2X1_276 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_10_OAI22X1_35 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_7_DFFSR_149 INVX1_23/gnd DFFSR_91/S FILL
XFILL_33_DFFSR_84 BUFX2_43/A DFFSR_23/S FILL
XFILL_24_DFFPOSX1_26 BUFX2_37/A DFFSR_81/S FILL
XFILL_44_DFFSR_44 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_8_NAND3X1_56 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_9_OAI22X1_38 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_48_DFFSR_180 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_38_DFFSR_183 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_7_NAND3X1_59 BUFX2_8/gnd DFFSR_25/S FILL
XINVX1_236 INVX1_236/A INVX1_8/gnd INVX1_236/Y DFFSR_7/S INVX1
XFILL_0_DFFSR_41 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_17_DFFSR_34 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_0_INVX1_126 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_8_OAI22X1_41 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_28_DFFSR_186 INVX1_23/gnd DFFSR_186/S FILL
XFILL_1_NAND2X1_210 BUFX2_35/A DFFSR_97/S FILL
XFILL_6_NAND3X1_62 BUFX2_43/A DFFSR_23/S FILL
XFILL_7_OAI22X1_44 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_5_NAND3X1_65 BUFX2_35/A DFFSR_14/S FILL
XFILL_18_DFFSR_189 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_10_XOR2X1_4 DFFSR_89/gnd DFFSR_186/S FILL
XNAND3X1_62 AOI22X1_8/C AOI22X1_8/D AOI21X1_25/A BUFX2_43/A NAND3X1_62/Y DFFSR_23/S
+ NAND3X1
XFILL_6_OAI22X1_47 BUFX2_37/A DFFSR_8/S FILL
XFILL_0_NAND3X1_108 BUFX2_37/A DFFSR_81/S FILL
XFILL_41_DFFSR_91 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_4_NAND3X1_68 BUFX2_35/A DFFSR_14/S FILL
XOAI22X1_47 INVX1_353/Y OAI22X1_39/B INVX1_352/Y OAI22X1_39/D BUFX2_37/A NOR2X1_33/B
+ DFFSR_8/S OAI22X1
XFILL_5_OAI22X1_50 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_3_NAND3X1_71 BUFX2_35/A DFFSR_14/S FILL
XFILL_51_DFFSR_107 BUFX2_36/A DFFSR_8/S FILL
XFILL_4_OAI22X1_53 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_2_NAND2X1_144 INVX1_8/gnd DFFSR_7/S FILL
XDFFSR_189 BUFX2_31/A DFFSR_1/CLK DFFSR_185/R DFFSR_1/S DFFSR_189/D DFFSR_1/gnd DFFSR_1/S
+ DFFSR
XFILL_8_OAI21X1_247 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_4_DFFSR_186 INVX1_23/gnd DFFSR_186/S FILL
XFILL_2_NAND3X1_74 BUFX2_35/A DFFSR_14/S FILL
XFILL_3_OAI22X1_56 BUFX2_37/A DFFSR_8/S FILL
XFILL_14_DFFSR_81 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_25_DFFSR_41 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_8_DFFSR_48 INVX1_4/gnd DFFSR_4/S FILL
XFILL_41_DFFSR_110 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_31_DFFSR_113 INVX1_23/gnd DFFSR_186/S FILL
XFILL_1_NAND3X1_77 BUFX2_37/A DFFSR_81/S FILL
XFILL_2_OAI22X1_59 INVX1_8/gnd DFFSR_7/S FILL
XFILL_0_NAND3X1_80 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_1_OAI22X1_62 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_21_DFFSR_116 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_0_OAI21X1_126 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_11_DFFSR_119 BUFX2_37/A DFFSR_81/S FILL
XFILL_26_1_1 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_4_NAND2X1_7 INVX1_89/gnd DFFSR_36/S FILL
XFILL_9_OAI21X1_181 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_0_OAI22X1_65 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_8_0_0 BUFX2_43/A DFFSR_97/S FILL
XFILL_1_INVX1_270 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_49_DFFSR_98 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_20_DFFSR_3 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_24_3_2 DFFSR_71/gnd DFFSR_10/S FILL
XOAI22X1_9 INVX1_274/Y OAI22X1_9/B OAI22X1_9/C OAI22X1_9/D INVX1_8/gnd OAI22X1_9/Y
+ DFFSR_5/S OAI22X1
XFILL_7_DFFSR_113 INVX1_23/gnd DFFSR_186/S FILL
XFILL_6_2_1 BUFX2_35/A DFFSR_14/S FILL
XINVX1_82 BUFX2_5/Y BUFX2_35/A DFFSR_68/R DFFSR_97/S INVX1
XFILL_0_NAND2X1_240 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_5_DFFSR_95 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_33_DFFSR_48 INVX1_4/gnd DFFSR_4/S FILL
XFILL_22_DFFSR_88 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_9_NAND3X1_17 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_48_DFFSR_144 INVX1_8/gnd DFFSR_5/S FILL
XFILL_4_OAI22X1_6 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_38_DFFSR_147 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_8_NAND3X1_20 BUFX2_37/A DFFSR_8/S FILL
XFILL_4_BUFX2_4 BUFX2_8/gnd DFFSR_25/S FILL
XINVX1_200 INVX1_200/A INVX1_4/gnd INVX1_200/Y DFFSR_4/S INVX1
XFILL_4_BUFX2_33 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_4_4_2 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_7_NAND3X1_23 BUFX2_37/A DFFSR_81/S FILL
XFILL_28_DFFSR_150 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_4_DFFPOSX1_12 INVX1_8/gnd DFFSR_5/S FILL
XFILL_35_7 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_1_NAND2X1_174 BUFX2_43/A DFFSR_97/S FILL
XFILL_18_DFFSR_153 BUFX2_36/A DFFSR_8/S FILL
XFILL_6_NAND3X1_26 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_4_INVX1_197 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_5_NAND3X1_29 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_6_OAI22X1_11 DFFSR_3/gnd DFFSR_4/S FILL
XNAND3X1_26 AOI21X1_4/B AOI21X1_4/A AOI21X1_4/C BUFX2_7/gnd NAND3X1_27/C DFFSR_81/S
+ NAND3X1
XFILL_30_DFFSR_95 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_41_DFFSR_55 INVX1_89/gnd DFFSR_36/S FILL
XFILL_2_INVX1_89 INVX1_89/gnd DFFSR_2/S FILL
XFILL_4_NAND3X1_32 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_5_OAI22X1_14 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_3_NAND3X1_35 BUFX2_35/A DFFSR_97/S FILL
XDFFSR_153 DFFSR_153/Q CLKBUF1_11/Y DFFSR_153/R DFFSR_8/S DFFSR_153/D BUFX2_36/A DFFSR_8/S
+ DFFSR
XFILL_2_NAND2X1_108 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_3_NOR2X1_32 INVX1_94/gnd DFFSR_52/S FILL
XFILL_4_OAI22X1_17 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_13_DFFPOSX1_31 BUFX2_17/gnd DFFSR_57/S FILL
XOAI22X1_11 INVX1_278/Y OAI22X1_8/B INVX1_277/Y OAI22X1_6/B DFFSR_3/gnd NOR2X1_15/A
+ DFFSR_4/S OAI22X1
XFILL_8_DFFSR_12 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_2_NAND3X1_38 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_3_OAI22X1_20 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_8_OAI21X1_211 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_2_INVX1_414 INVX1_2/gnd DFFSR_1/S FILL
XFILL_1_NAND3X1_41 BUFX2_43/A DFFSR_23/S FILL
XFILL_4_DFFSR_150 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_14_DFFSR_45 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_2_OAI22X1_23 INVX1_89/gnd DFFSR_2/S FILL
XFILL_45_DFFSR_181 INVX1_23/gnd DFFSR_186/S FILL
XFILL_0_NAND3X1_44 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_1_OAI22X1_26 INVX1_94/gnd DFFSR_52/S FILL
XFILL_23_DFFPOSX1_20 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_0_OAI22X1_29 INVX1_8/gnd DFFSR_5/S FILL
XFILL_35_DFFSR_184 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_49_DFFSR_62 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_1_INVX1_234 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_25_DFFSR_187 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_15_DFFSR_190 DFFSR_9/gnd DFFSR_9/S FILL
XDFFSR_99 DFFSR_99/Q INVX1_172/A DFFSR_97/R DFFSR_97/S DFFSR_99/D BUFX2_35/A DFFSR_97/S
+ DFFSR
XFILL_0_NAND2X1_204 BUFX2_5/gnd DFFSR_6/S FILL
XINVX1_46 BUFX2_10/Y DFFSR_71/gnd DFFSR_33/R DFFSR_45/S INVX1
XFILL_11_DFFSR_92 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_33_DFFSR_12 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_22_DFFSR_52 INVX1_94/gnd DFFSR_52/S FILL
XFILL_5_DFFSR_59 INVX1_4/gnd DFFSR_51/S FILL
XFILL_48_DFFSR_108 INVX1_89/gnd DFFSR_2/S FILL
XINVX1_164 DFFSR_145/Q INVX1_23/gnd INVX1_164/Y DFFSR_91/S INVX1
XFILL_38_DFFSR_111 INVX1_8/gnd DFFSR_5/S FILL
XFILL_1_DFFSR_187 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_7_OAI21X1_241 BUFX2_35/A DFFSR_97/S FILL
XFILL_4_INVX1_161 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_28_DFFSR_114 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_1_NAND2X1_138 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_18_DFFSR_117 INVX1_23/gnd DFFSR_91/S FILL
XFILL_1_NAND2X1_8 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_19_DFFSR_99 BUFX2_35/A DFFSR_97/S FILL
XFILL_2_INVX1_53 INVX1_89/gnd DFFSR_2/S FILL
XFILL_41_DFFSR_19 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_30_DFFSR_59 INVX1_4/gnd DFFSR_51/S FILL
XDFFSR_117 DFFSR_117/Q CLKBUF1_7/Y DFFSR_113/R DFFSR_91/S DFFSR_117/D INVX1_23/gnd
+ DFFSR_91/S DFFSR
XFILL_8_OAI21X1_175 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_2_INVX1_378 INVX1_8/gnd DFFSR_7/S FILL
XFILL_4_DFFSR_114 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_45_DFFSR_145 INVX1_23/gnd DFFSR_186/S FILL
XFILL_1_OAI22X1_7 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_35_DFFSR_148 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_8_DFFSR_2 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_25_DFFSR_151 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_15_DFFSR_154 BUFX2_36/A DFFSR_6/S FILL
XFILL_1_INVX1_198 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_49_DFFSR_26 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_38_DFFSR_66 INVX1_2/gnd DFFSR_51/S FILL
XFILL_5_DFFSR_23 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_0_NAND2X1_168 BUFX2_36/A DFFSR_6/S FILL
XINVX1_10 BUFX2_10/Y BUFX2_7/gnd DFFSR_6/R DFFSR_81/S INVX1
XDFFSR_63 DFFSR_63/Q DFFSR_28/CLK DFFSR_61/R DFFSR_52/S DFFSR_63/D INVX1_94/gnd DFFSR_52/S
+ DFFSR
XFILL_22_DFFSR_16 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_11_DFFSR_56 INVX1_2/gnd DFFSR_51/S FILL
XFILL_6_OR2X2_2 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_0_NOR2X1_33 BUFX2_37/A DFFSR_81/S FILL
XINVX1_128 DFFSR_113/Q INVX1_23/gnd INVX1_128/Y DFFSR_91/S INVX1
XFILL_8_NAND3X1_121 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_1_DFFSR_151 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_12_DFFPOSX1_25 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_4_NOR2X1_4 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_25_4_0 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_32_DFFSR_6 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_7_OAI21X1_205 BUFX2_36/A DFFSR_8/S FILL
XFILL_42_DFFSR_182 INVX1_89/gnd DFFSR_36/S FILL
XFILL_4_INVX1_125 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_1_NAND2X1_102 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_46_DFFSR_73 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_32_DFFSR_185 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_5_5_0 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_30_DFFSR_23 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_19_DFFSR_63 INVX1_94/gnd DFFSR_52/S FILL
XFILL_2_INVX1_17 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_2_DFFSR_70 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_22_DFFSR_188 INVX1_2/gnd DFFSR_1/S FILL
XFILL_12_DFFSR_191 INVX1_23/gnd DFFSR_91/S FILL
XFILL_22_DFFPOSX1_14 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_2_INVX1_342 INVX1_8/gnd DFFSR_7/S FILL
XFILL_8_OAI21X1_139 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_8_DFFSR_185 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_45_DFFSR_109 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_35_DFFSR_112 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_25_DFFSR_115 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_38_DFFSR_30 INVX1_89/gnd DFFSR_36/S FILL
XFILL_1_INVX1_162 INVX1_8/gnd DFFSR_7/S FILL
XFILL_27_DFFSR_70 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_15_DFFSR_118 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_6_OAI21X1_235 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_0_NAND2X1_132 INVX1_8/gnd DFFSR_5/S FILL
XDFFSR_27 INVX1_31/A DFFSR_24/CLK DFFSR_31/R DFFSR_1/S DFFSR_27/D DFFSR_1/gnd DFFSR_1/S
+ DFFSR
XFILL_11_DFFSR_20 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_1_DFFSR_115 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_17_4 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_2_NOR3X1_1 INVX1_94/gnd DFFSR_52/S FILL
XFILL_8_OAI22X1_5 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_42_DFFSR_146 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_7_OAI21X1_169 BUFX2_36/A DFFSR_8/S FILL
XFILL_46_DFFSR_37 INVX1_89/gnd DFFSR_2/S FILL
XFILL_33_1_1 INVX1_8/gnd DFFSR_7/S FILL
XFILL_32_DFFSR_149 INVX1_23/gnd DFFSR_91/S FILL
XFILL_35_DFFSR_77 INVX1_89/gnd DFFSR_2/S FILL
XFILL_22_DFFSR_152 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_31_3_2 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_12_DFFSR_155 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_19_DFFSR_27 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_2_DFFSR_34 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_2_INVX1_306 INVX1_94/gnd DFFSR_25/S FILL
XFILL_8_OAI21X1_103 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_20_CLKBUF1_17 INVX1_94/gnd DFFSR_25/S FILL
XFILL_8_DFFSR_149 INVX1_23/gnd DFFSR_91/S FILL
XFILL_5_OAI21X1_265 BUFX2_43/A DFFSR_97/S FILL
XFILL_43_DFFSR_84 BUFX2_43/A DFFSR_23/S FILL
XFILL_19_CLKBUF1_20 INVX1_4/gnd DFFSR_51/S FILL
XFILL_18_CLKBUF1_23 INVX1_89/gnd DFFSR_2/S FILL
XFILL_49_DFFSR_180 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_39_DFFSR_183 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_7_NAND3X1_115 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_27_DFFSR_34 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_16_DFFSR_74 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_1_INVX1_126 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_29_DFFSR_186 INVX1_23/gnd DFFSR_186/S FILL
XFILL_3_BUFX2_1 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_11_DFFPOSX1_19 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_6_OAI21X1_199 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_19_DFFSR_189 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_51_DFFSR_91 BUFX2_6/gnd DFFSR_91/S FILL
XOAI21X1_235 AOI21X1_30/Y AOI21X1_31/Y INVX1_260/Y BUFX2_6/gnd AOI21X1_33/A DFFSR_91/S
+ OAI21X1
XFILL_5_DFFSR_186 INVX1_23/gnd DFFSR_186/S FILL
XFILL_7_OAI21X1_133 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_24_DFFSR_81 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_35_DFFSR_41 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_7_DFFSR_88 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_42_DFFSR_110 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_32_DFFSR_113 INVX1_23/gnd DFFSR_186/S FILL
XFILL_1_DFFPOSX1_30 BUFX2_43/A DFFSR_97/S FILL
XFILL_22_DFFSR_116 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_12_DFFSR_119 BUFX2_37/A DFFSR_81/S FILL
XFILL_5_NAND2X1_7 INVX1_89/gnd DFFSR_36/S FILL
XFILL_6_BUFX2_26 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_2_INVX1_270 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_44_DFFSR_9 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_8_DFFSR_113 INVX1_23/gnd DFFSR_186/S FILL
XFILL_4_INVX1_82 BUFX2_35/A DFFSR_97/S FILL
XFILL_43_DFFSR_48 INVX1_4/gnd DFFSR_4/S FILL
XFILL_32_DFFSR_88 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_5_OAI21X1_229 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_49_DFFSR_144 INVX1_8/gnd DFFSR_5/S FILL
XFILL_5_OAI22X1_6 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_39_DFFSR_147 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_29_DFFSR_150 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_16_DFFSR_38 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_39_4 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_19_DFFSR_153 BUFX2_36/A DFFSR_8/S FILL
XFILL_6_OAI21X1_163 DFFSR_3/gnd DFFSR_4/S FILL
XNOR2X1_35 NOR2X1_35/A NOR2X1_35/B INVX1_94/gnd NOR2X1_35/Y DFFSR_52/S NOR2X1
XFILL_40_DFFSR_95 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_4_NOR2X1_32 INVX1_94/gnd DFFSR_52/S FILL
XOAI21X1_199 NAND3X1_2/A NAND2X1_197/Y NAND3X1_34/Y DFFSR_73/gnd DFFPOSX1_6/D DFFSR_57/S
+ OAI21X1
XFILL_1_AND2X2_4 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_7_DFFSR_52 INVX1_94/gnd DFFSR_52/S FILL
XFILL_6_NAND2X1_277 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_3_INVX1_414 INVX1_2/gnd DFFSR_1/S FILL
XFILL_5_DFFSR_150 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_13_DFFSR_85 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_24_DFFSR_45 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_46_DFFSR_181 INVX1_23/gnd DFFSR_186/S FILL
XFILL_10_CLKBUF1_11 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_4_OAI21X1_259 INVX1_23/gnd DFFSR_186/S FILL
XFILL_36_DFFSR_184 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_9_CLKBUF1_14 BUFX2_43/A DFFSR_23/S FILL
XFILL_2_INVX1_234 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_26_DFFSR_187 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_8_CLKBUF1_17 INVX1_94/gnd DFFSR_25/S FILL
XFILL_10_DFFSR_7 INVX1_8/gnd DFFSR_7/S FILL
XFILL_16_DFFSR_190 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_10_DFFPOSX1_13 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_6_NAND3X1_109 BUFX2_36/A DFFSR_8/S FILL
XFILL_32_4_0 INVX1_8/gnd DFFSR_5/S FILL
XFILL_7_CLKBUF1_20 INVX1_4/gnd DFFSR_51/S FILL
XFILL_21_DFFSR_92 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_43_DFFSR_12 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_4_DFFSR_99 BUFX2_35/A DFFSR_97/S FILL
XFILL_5_OAI21X1_193 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_32_DFFSR_52 INVX1_94/gnd DFFSR_52/S FILL
XFILL_6_CLKBUF1_23 INVX1_89/gnd DFFSR_2/S FILL
XFILL_49_DFFSR_108 INVX1_89/gnd DFFSR_2/S FILL
XOR2X2_3 OR2X2_3/A OR2X2_3/B BUFX2_43/A OR2X2_3/Y DFFSR_23/S OR2X2
XCLKBUF1_23 INVX1_402/Y INVX1_89/gnd DFFSR_2/CLK DFFSR_2/S CLKBUF1
XFILL_39_DFFSR_111 INVX1_8/gnd DFFSR_5/S FILL
XFILL_2_DFFSR_187 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_3_BUFX2_37 BUFX2_37/A DFFSR_81/S FILL
XFILL_29_DFFSR_114 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_19_DFFSR_117 INVX1_23/gnd DFFSR_91/S FILL
XFILL_6_OAI21X1_127 BUFX2_43/A DFFSR_23/S FILL
XFILL_2_NAND2X1_8 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_31_DFFSR_3 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_29_DFFSR_99 BUFX2_35/A DFFSR_97/S FILL
XFILL_0_DFFPOSX1_24 BUFX2_43/A DFFSR_23/S FILL
XFILL_51_DFFSR_19 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_1_INVX1_93 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_40_DFFSR_59 INVX1_4/gnd DFFSR_51/S FILL
XFILL_3_INVX1_378 INVX1_8/gnd DFFSR_7/S FILL
XFILL_6_NAND2X1_241 BUFX2_17/gnd DFFSR_57/S FILL
XOAI21X1_163 BUFX2_1/Y INVX1_197/Y NAND2X1_163/Y DFFSR_3/gnd DFFSR_163/D DFFSR_4/S
+ OAI21X1
XFILL_7_DFFSR_16 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_5_DFFSR_114 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_13_DFFSR_49 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_46_DFFSR_145 INVX1_23/gnd DFFSR_186/S FILL
XFILL_2_OAI22X1_7 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_36_DFFSR_148 DFFSR_89/gnd DFFSR_92/S FILL
XNAND2X1_277 DFFSR_133/Q INVX1_159/A DFFSR_71/gnd AND2X2_16/B DFFSR_10/S NAND2X1
XFILL_4_OAI21X1_223 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_26_DFFSR_151 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_16_DFFSR_154 BUFX2_36/A DFFSR_6/S FILL
XFILL_2_INVX1_198 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_48_DFFSR_66 INVX1_2/gnd DFFSR_51/S FILL
XFILL_4_DFFSR_63 INVX1_94/gnd DFFSR_52/S FILL
XFILL_32_DFFSR_16 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_10_DFFSR_96 INVX1_2/gnd DFFSR_1/S FILL
XFILL_21_DFFSR_56 INVX1_2/gnd DFFSR_51/S FILL
XFILL_40_1_1 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_5_OAI21X1_157 BUFX2_35/A DFFSR_97/S FILL
XFILL_1_NOR2X1_33 BUFX2_37/A DFFSR_81/S FILL
XNAND3X1_109 INVX1_251/A AOI21X1_38/B OR2X2_3/Y BUFX2_36/A NAND3X1_109/Y DFFSR_8/S
+ NAND3X1
XFILL_0_INVX1_415 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_2_DFFSR_151 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_38_3_2 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_43_DFFSR_182 INVX1_89/gnd DFFSR_36/S FILL
XFILL_5_NAND2X1_271 INVX1_89/gnd DFFSR_2/S FILL
XFILL_33_DFFSR_185 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_40_DFFSR_23 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_29_DFFSR_63 INVX1_94/gnd DFFSR_52/S FILL
XFILL_1_INVX1_57 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_23_DFFSR_188 INVX1_2/gnd DFFSR_1/S FILL
XFILL_3_OAI21X1_253 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_13_DFFSR_191 INVX1_23/gnd DFFSR_91/S FILL
XOAI21X1_127 BUFX2_21/Y INVX1_143/Y OAI21X1_127/C BUFX2_43/A DFFSR_127/D DFFSR_23/S
+ OAI21X1
XFILL_6_NAND2X1_205 BUFX2_36/A DFFSR_6/S FILL
XFILL_3_INVX1_342 INVX1_8/gnd DFFSR_7/S FILL
XFILL_13_DFFSR_13 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_9_DFFSR_185 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_5_NAND3X1_103 INVX1_23/gnd DFFSR_186/S FILL
XFILL_46_DFFSR_109 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_4_OAI21X1_187 BUFX2_37/A DFFSR_8/S FILL
XNAND2X1_241 NOR2X1_26/Y NOR2X1_27/Y BUFX2_17/gnd NAND2X1_72/B DFFSR_57/S NAND2X1
XFILL_36_DFFSR_112 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_26_DFFSR_115 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_48_DFFSR_30 INVX1_89/gnd DFFSR_36/S FILL
XFILL_2_INVX1_162 INVX1_8/gnd DFFSR_7/S FILL
XFILL_37_DFFSR_70 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_16_DFFSR_118 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_21_DFFSR_20 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_5_OAI21X1_121 BUFX2_36/A DFFSR_8/S FILL
XFILL_10_DFFSR_60 BUFX2_37/A DFFSR_8/S FILL
XFILL_4_DFFSR_27 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_2_DFFSR_115 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_3_NOR2X1_8 BUFX2_43/A DFFSR_23/S FILL
XFILL_21_1 INVX1_94/gnd DFFSR_52/S FILL
XFILL_0_INVX1_379 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_9_OAI22X1_5 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_43_DFFSR_146 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_33_DFFSR_149 INVX1_23/gnd DFFSR_91/S FILL
XFILL_45_DFFSR_77 INVX1_89/gnd DFFSR_2/S FILL
XFILL_5_NAND2X1_235 INVX1_4/gnd DFFSR_51/S FILL
XFILL_23_DFFSR_152 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_4_NAND3X1_133 INVX1_8/gnd DFFSR_5/S FILL
XFILL_13_DFFSR_155 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_29_DFFSR_27 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_1_INVX1_21 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_1_DFFSR_74 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_18_DFFSR_67 INVX1_2/gnd DFFSR_51/S FILL
XFILL_3_OAI21X1_217 INVX1_23/gnd DFFSR_91/S FILL
XFILL_6_NAND2X1_169 BUFX2_36/A DFFSR_8/S FILL
XFILL_3_INVX1_306 INVX1_94/gnd DFFSR_25/S FILL
XFILL_5_XOR2X1_4 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_0_BUFX2_12 BUFX2_37/A DFFSR_81/S FILL
XFILL_21_DFFPOSX1_2 INVX1_89/gnd DFFSR_36/S FILL
XFILL_9_DFFSR_149 INVX1_23/gnd DFFSR_91/S FILL
XFILL_43_DFFSR_6 BUFX2_5/gnd DFFSR_6/S FILL
XNAND2X1_205 BUFX2_13/Y AND2X2_10/B BUFX2_36/A NOR2X1_9/A DFFSR_6/S NAND2X1
XFILL_20_DFFPOSX1_5 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_12_1_2 BUFX2_36/A DFFSR_6/S FILL
XFILL_18_DFFPOSX1_26 BUFX2_37/A DFFSR_81/S FILL
XFILL_4_OAI21X1_151 BUFX2_37/A DFFSR_81/S FILL
XFILL_19_DFFPOSX1_8 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_50_DFFSR_180 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_40_DFFSR_183 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_9_DFFSR_81 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_37_DFFSR_34 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_26_DFFSR_74 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_2_INVX1_126 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_30_DFFSR_186 INVX1_23/gnd DFFSR_186/S FILL
XFILL_4_NAND2X1_265 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_20_DFFSR_189 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_10_DFFSR_24 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_0_INVX1_343 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_4_5 INVX1_23/gnd DFFSR_91/S FILL
XFILL_6_DFFSR_186 INVX1_23/gnd DFFSR_186/S FILL
XFILL_5_NAND2X1_199 BUFX2_36/A DFFSR_8/S FILL
XFILL_34_DFFSR_81 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_45_DFFSR_41 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_2_OAI21X1_247 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_43_DFFSR_110 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_33_DFFSR_113 INVX1_23/gnd DFFSR_186/S FILL
XFILL_18_DFFSR_31 BUFX2_35/A DFFSR_97/S FILL
XFILL_23_DFFSR_116 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_1_DFFSR_38 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_39_4_0 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_13_DFFSR_119 BUFX2_37/A DFFSR_81/S FILL
XFILL_6_NAND2X1_7 INVX1_89/gnd DFFSR_36/S FILL
XFILL_3_OAI21X1_181 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_6_NAND2X1_133 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_3_INVX1_270 DFFSR_79/gnd DFFSR_36/S FILL
XXOR2X1_8 XOR2X1_8/A XOR2X1_8/B BUFX2_5/gnd OR2X2_3/B DFFSR_6/S XOR2X1
XFILL_9_DFFSR_113 INVX1_23/gnd DFFSR_186/S FILL
XFILL_11_XOR2X1_1 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_42_DFFSR_88 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_4_OAI21X1_115 BUFX2_36/A DFFSR_6/S FILL
XNAND2X1_169 DFFSR_8/S NAND2X1_169/B BUFX2_36/A NAND2X1_169/Y DFFSR_8/S NAND2X1
XFILL_50_DFFSR_144 INVX1_8/gnd DFFSR_5/S FILL
XFILL_6_OAI22X1_6 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_40_DFFSR_147 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_26_6 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_9_DFFSR_45 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_30_DFFSR_150 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_26_DFFSR_38 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_15_DFFSR_78 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_43_1 INVX1_4/gnd DFFSR_4/S FILL
XFILL_20_DFFSR_153 BUFX2_36/A DFFSR_8/S FILL
XFILL_10_DFFSR_156 INVX1_23/gnd DFFSR_91/S FILL
XFILL_4_NAND2X1_229 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_0_INVX1_307 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_50_DFFSR_95 DFFSR_79/gnd DFFSR_45/S FILL
XINVX1_417 BUFX2_28/A INVX1_23/gnd INVX1_417/Y DFFSR_91/S INVX1
XFILL_5_NOR2X1_32 INVX1_94/gnd DFFSR_52/S FILL
XFILL_3_NAND3X1_127 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_2_OAI21X1_211 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_6_DFFSR_92 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_6_DFFSR_150 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_23_DFFSR_85 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_34_DFFSR_45 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_5_NAND2X1_163 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_47_DFFSR_181 INVX1_23/gnd DFFSR_186/S FILL
XFILL_37_DFFSR_184 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_3_OAI21X1_145 INVX1_23/gnd DFFSR_91/S FILL
XFILL_17_DFFPOSX1_20 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_3_INVX1_234 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_47_1_1 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_5_BUFX2_30 INVX1_4/gnd DFFSR_51/S FILL
XFILL_27_DFFSR_187 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_17_DFFSR_190 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_9_DFFPOSX1_2 INVX1_89/gnd DFFSR_36/S FILL
XFILL_45_3_2 INVX1_2/gnd DFFSR_1/S FILL
XFILL_31_DFFSR_92 DFFSR_89/gnd DFFSR_92/S FILL
XNAND2X1_133 DFFSR_54/S NAND2X1_69/B BUFX2_19/gnd OAI21X1_133/C DFFSR_54/S NAND2X1
XFILL_3_INVX1_86 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_42_DFFSR_52 INVX1_94/gnd DFFSR_52/S FILL
XFILL_8_DFFPOSX1_5 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_3_NAND2X1_259 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_8_AOI21X1_25 BUFX2_43/A DFFSR_97/S FILL
XFILL_7_DFFPOSX1_8 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_50_DFFSR_108 INVX1_89/gnd DFFSR_2/S FILL
XFILL_7_AOI21X1_28 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_40_DFFSR_111 INVX1_8/gnd DFFSR_5/S FILL
XFILL_15_DFFSR_42 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_3_DFFSR_187 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_6_AOI21X1_31 INVX1_23/gnd DFFSR_186/S FILL
XFILL_30_DFFSR_114 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_20_DFFSR_117 INVX1_23/gnd DFFSR_91/S FILL
XFILL_1_OAI21X1_241 BUFX2_35/A DFFSR_97/S FILL
XFILL_4_NAND2X1_193 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_5_AOI21X1_34 INVX1_94/gnd DFFSR_25/S FILL
XFILL_7_DFFPOSX1_31 BUFX2_17/gnd DFFSR_57/S FILL
XAOI21X1_31 AOI21X1_31/A AOI21X1_31/B XOR2X1_6/Y INVX1_23/gnd AOI21X1_31/Y DFFSR_186/S
+ AOI21X1
XFILL_3_NAND2X1_8 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_13_2_0 BUFX2_36/A DFFSR_8/S FILL
XFILL_4_AOI21X1_37 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_10_DFFSR_120 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_39_DFFSR_99 BUFX2_35/A DFFSR_97/S FILL
XINVX1_381 DFFSR_79/Q DFFSR_79/gnd INVX1_381/Y DFFSR_45/S INVX1
XFILL_0_INVX1_271 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_50_DFFSR_59 INVX1_4/gnd DFFSR_51/S FILL
XFILL_3_AOI21X1_40 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_11_4_1 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_2_AOI21X1_43 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_12_DFFSR_89 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_2_OAI21X1_175 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_0_AND2X2_8 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_5_NAND2X1_127 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_6_DFFSR_114 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_1_AOI21X1_46 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_4_INVX1_378 INVX1_8/gnd DFFSR_7/S FILL
XFILL_6_DFFSR_56 INVX1_2/gnd DFFSR_51/S FILL
XFILL_23_DFFSR_49 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_47_DFFSR_145 INVX1_23/gnd DFFSR_186/S FILL
XFILL_3_OAI22X1_7 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_37_DFFSR_148 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_3_OAI21X1_109 BUFX2_5/gnd DFFSR_6/S FILL
XBUFX2_34 BUFX2_37/A BUFX2_37/A BUFX2_34/Y DFFSR_81/S BUFX2
XFILL_27_DFFSR_151 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_17_DFFSR_154 BUFX2_36/A DFFSR_6/S FILL
XFILL_3_INVX1_198 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_48_6 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_8_OAI21X1_73 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_7_OAI21X1_76 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_3_INVX1_50 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_42_DFFSR_16 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_20_DFFSR_96 INVX1_2/gnd DFFSR_1/S FILL
XFILL_31_DFFSR_56 INVX1_2/gnd DFFSR_51/S FILL
XFILL_6_NAND2X1_94 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_3_NAND2X1_223 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_5_NAND2X1_97 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_2_NOR2X1_33 BUFX2_37/A DFFSR_81/S FILL
XFILL_6_OAI21X1_79 INVX1_89/gnd DFFSR_36/S FILL
XFILL_1_INVX1_415 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_5_OAI21X1_82 DFFSR_9/gnd DFFSR_9/S FILL
XNAND2X1_94 BUFX2_16/Y INVX1_97/A BUFX2_16/gnd NAND2X1_94/Y DFFSR_11/S NAND2X1
XFILL_2_BUFX2_41 BUFX2_37/A DFFSR_81/S FILL
XFILL_3_DFFSR_151 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_4_OAI21X1_85 DFFSR_79/gnd DFFSR_45/S FILL
XOAI21X1_79 BUFX2_22/Y INVX1_89/Y NAND2X1_79/Y INVX1_89/gnd DFFSR_79/D DFFSR_36/S
+ OAI21X1
XFILL_2_NAND3X1_121 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_1_OAI21X1_205 BUFX2_36/A DFFSR_8/S FILL
XFILL_44_DFFSR_182 INVX1_89/gnd DFFSR_36/S FILL
XFILL_3_OAI21X1_88 INVX1_4/gnd DFFSR_4/S FILL
XFILL_34_DFFSR_185 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_4_NAND2X1_157 BUFX2_35/A DFFSR_97/S FILL
XFILL_2_OAI21X1_91 BUFX2_43/A DFFSR_97/S FILL
XFILL_21_DFFSR_7 INVX1_8/gnd DFFSR_7/S FILL
XFILL_50_DFFSR_23 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_39_DFFSR_63 INVX1_94/gnd DFFSR_52/S FILL
XFILL_24_DFFSR_188 INVX1_2/gnd DFFSR_1/S FILL
XFILL_0_INVX1_235 INVX1_4/gnd DFFSR_51/S FILL
XFILL_0_INVX1_97 INVX1_4/gnd DFFSR_4/S FILL
XFILL_1_OAI21X1_94 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_14_DFFSR_191 INVX1_23/gnd DFFSR_91/S FILL
XFILL_0_OAI21X1_97 BUFX2_5/gnd DFFSR_23/S FILL
XINVX1_345 DFFSR_122/Q INVX1_94/gnd INVX1_345/Y DFFSR_52/S INVX1
XFILL_16_DFFPOSX1_14 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_4_INVX1_342 INVX1_8/gnd DFFSR_7/S FILL
XFILL_2_OAI21X1_139 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_6_DFFSR_20 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_19_1_2 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_5_BUFX2_8 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_12_DFFSR_53 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_1_AOI21X1_10 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_23_DFFSR_13 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_1_0_1 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_47_DFFSR_109 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_0_AOI21X1_13 INVX1_8/gnd DFFSR_7/S FILL
XFILL_5_NOR2X1_1 BUFX2_36/A DFFSR_6/S FILL
XFILL_0_DFFSR_188 INVX1_2/gnd DFFSR_1/S FILL
XFILL_37_DFFSR_112 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_27_DFFSR_115 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_2_NAND2X1_253 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_3_INVX1_162 INVX1_8/gnd DFFSR_7/S FILL
XFILL_9_OAI21X1_34 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_42_DFFSR_3 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_8_OAI21X1_37 INVX1_89/gnd DFFSR_2/S FILL
XFILL_47_DFFSR_70 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_17_DFFSR_118 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_7_OAI21X1_40 INVX1_8/gnd DFFSR_7/S FILL
XFILL_0_NAND2X1_9 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_6_NAND2X1_58 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_31_DFFSR_20 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_0_OAI21X1_235 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_3_INVX1_14 BUFX2_35/A DFFSR_14/S FILL
XFILL_3_NAND2X1_187 BUFX2_37/A DFFSR_8/S FILL
XFILL_20_DFFSR_60 BUFX2_37/A DFFSR_8/S FILL
XFILL_5_NAND2X1_61 BUFX2_37/A DFFSR_81/S FILL
XFILL_6_DFFPOSX1_25 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_6_OAI21X1_43 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_3_DFFSR_67 INVX1_2/gnd DFFSR_51/S FILL
XFILL_5_OAI21X1_46 BUFX2_37/A DFFSR_81/S FILL
XNAND2X1_58 DFFSR_65/S INVX1_57/A DFFSR_3/gnd NAND2X1_58/Y DFFSR_65/S NAND2X1
XFILL_4_NAND2X1_64 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_3_DFFSR_115 BUFX2_6/gnd DFFSR_14/S FILL
XOAI21X1_43 DFFSR_25/S INVX1_49/Y OAI21X1_43/C BUFX2_8/gnd DFFSR_43/D DFFSR_10/S OAI21X1
XFILL_1_INVX1_379 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_3_NAND2X1_67 INVX1_2/gnd DFFSR_1/S FILL
XFILL_44_DFFSR_146 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_0_OAI22X1_8 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_46_4_0 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_4_OAI21X1_49 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_34_DFFSR_149 INVX1_23/gnd DFFSR_91/S FILL
XFILL_1_OAI21X1_169 BUFX2_36/A DFFSR_8/S FILL
XFILL_4_NAND2X1_121 BUFX2_36/A DFFSR_8/S FILL
XFILL_3_OAI21X1_52 INVX1_94/gnd DFFSR_25/S FILL
XFILL_2_NAND2X1_70 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_24_DFFSR_152 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_2_OAI21X1_55 INVX1_89/gnd DFFSR_2/S FILL
XFILL_1_NAND2X1_73 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_0_INVX1_199 BUFX2_35/A DFFSR_97/S FILL
XFILL_0_INVX1_61 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_14_DFFSR_155 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_0_NAND2X1_76 BUFX2_19/gnd DFFSR_52/S FILL
XINVX1_309 INVX1_43/A DFFSR_79/gnd INVX1_309/Y DFFSR_36/S INVX1
XFILL_39_DFFSR_27 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_28_DFFSR_67 INVX1_2/gnd DFFSR_51/S FILL
XFILL_1_OAI21X1_58 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_0_OAI21X1_61 BUFX2_36/A DFFSR_8/S FILL
XFILL_4_INVX1_306 INVX1_94/gnd DFFSR_25/S FILL
XFILL_1_NAND2X1_283 INVX1_89/gnd DFFSR_36/S FILL
XFILL_12_DFFSR_17 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_2_OAI21X1_103 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_0_DFFSR_152 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_2_NAND2X1_217 BUFX2_8/gnd DFFSR_10/S FILL
XNOR2X1_5 NOR2X1_5/A NOR2X1_5/B BUFX2_17/gnd AND2X2_3/A DFFSR_57/S NOR2X1
XFILL_41_DFFSR_183 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_47_DFFSR_34 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_36_DFFSR_74 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_3_INVX1_126 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_31_DFFSR_186 INVX1_23/gnd DFFSR_186/S FILL
XFILL_1_NAND3X1_115 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_3_DFFSR_31 BUFX2_35/A DFFSR_97/S FILL
XFILL_6_NAND2X1_22 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_21_DFFSR_189 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_20_DFFSR_24 BUFX2_16/gnd DFFSR_65/S FILL
XNAND2X1_22 DFFSR_54/S DFFSR_14/Q BUFX2_19/gnd NAND2X1_22/Y DFFSR_52/S NAND2X1
XFILL_3_NAND2X1_151 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_5_NAND2X1_25 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_0_OAI21X1_199 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_8_2 BUFX2_35/A DFFSR_97/S FILL
XFILL_4_NAND2X1_28 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_5_OAI21X1_10 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_1_INVX1_343 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_3_NAND2X1_31 BUFX2_43/A DFFSR_97/S FILL
XFILL_9_DFFSR_6 BUFX2_5/gnd DFFSR_6/S FILL
XDFFPOSX1_25 AND2X2_6/B CLKBUF1_16/Y XOR2X1_14/Y BUFX2_19/gnd DFFSR_54/S DFFPOSX1
XFILL_4_OAI21X1_13 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_7_DFFSR_186 INVX1_23/gnd DFFSR_186/S FILL
XFILL_1_OAI21X1_133 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_44_DFFSR_81 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_3_OAI21X1_16 INVX1_89/gnd DFFSR_36/S FILL
XFILL_2_NAND2X1_34 INVX1_2/gnd DFFSR_1/S FILL
XFILL_44_DFFSR_110 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_34_DFFSR_113 INVX1_23/gnd DFFSR_186/S FILL
XFILL_1_NAND2X1_37 INVX1_8/gnd DFFSR_5/S FILL
XFILL_2_OAI21X1_19 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_8_NAND3X1_93 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_0_INVX1_163 INVX1_94/gnd DFFSR_52/S FILL
XFILL_0_INVX1_25 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_1_OAI21X1_22 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_24_DFFSR_116 DFFSR_5/gnd DFFSR_2/S FILL
XAOI21X1_1 AOI21X1_1/A INVX1_223/A AOI21X1_1/C INVX1_8/gnd NOR2X1_5/A DFFSR_5/S AOI21X1
XINVX1_273 DFFSR_2/Q INVX1_8/gnd OAI22X1_9/C DFFSR_5/S INVX1
XFILL_0_DFFSR_78 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_0_NAND2X1_40 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_28_DFFSR_31 BUFX2_35/A DFFSR_97/S FILL
XFILL_7_NAND3X1_96 BUFX2_43/A DFFSR_97/S FILL
XFILL_14_DFFSR_119 BUFX2_37/A DFFSR_81/S FILL
XFILL_0_OAI21X1_25 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_17_DFFSR_71 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_6_NAND3X1_99 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_4_INVX1_270 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_1_NAND2X1_247 INVX1_8/gnd DFFSR_5/S FILL
XNAND3X1_99 NOR2X1_11/Y NAND3X1_95/A NAND3X1_95/B BUFX2_6/gnd AOI21X1_31/B DFFSR_14/S
+ NAND3X1
XFILL_4_XOR2X1_8 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_0_DFFSR_116 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_5_DFFPOSX1_19 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_7_OAI22X1_6 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_41_DFFSR_147 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_2_NAND2X1_181 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_20_2_0 INVX1_94/gnd DFFSR_52/S FILL
XFILL_30_3 INVX1_89/gnd DFFSR_2/S FILL
XFILL_31_DFFSR_150 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_8_DFFSR_85 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_36_DFFSR_38 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_25_DFFSR_78 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_21_DFFSR_153 BUFX2_36/A DFFSR_8/S FILL
XFILL_11_DFFSR_156 INVX1_23/gnd DFFSR_91/S FILL
XFILL_3_NAND2X1_115 BUFX2_36/A DFFSR_6/S FILL
XFILL_18_4_1 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_0_OAI21X1_163 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_0_3_0 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_9_OAI21X1_218 INVX1_23/gnd DFFSR_186/S FILL
XFILL_2_AOI22X1_12 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_1_INVX1_307 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_6_NOR2X1_32 INVX1_94/gnd DFFSR_52/S FILL
XFILL_17_NOR3X1_2 INVX1_89/gnd DFFSR_2/S FILL
XFILL_0_NAND2X1_277 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_10_OAI22X1_36 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_9_NAND3X1_54 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_7_DFFSR_150 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_24_DFFPOSX1_27 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_33_DFFSR_85 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_44_DFFSR_45 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_48_DFFSR_181 INVX1_23/gnd DFFSR_186/S FILL
XFILL_9_OAI22X1_39 BUFX2_37/A DFFSR_8/S FILL
XFILL_8_NAND3X1_57 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_17_DFFSR_35 DFFSR_5/gnd DFFSR_2/S FILL
XINVX1_237 INVX1_237/A INVX1_8/gnd INVX1_237/Y DFFSR_7/S INVX1
XFILL_38_DFFSR_184 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_0_INVX1_127 INVX1_2/gnd DFFSR_1/S FILL
XFILL_0_DFFSR_42 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_1_NAND2X1_211 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_7_NAND3X1_60 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_8_OAI22X1_42 INVX1_8/gnd DFFSR_7/S FILL
XFILL_28_DFFSR_187 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_6_NAND3X1_63 BUFX2_43/A DFFSR_23/S FILL
XFILL_7_OAI22X1_45 INVX1_89/gnd DFFSR_2/S FILL
XFILL_18_DFFSR_190 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_10_XOR2X1_5 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_5_NAND3X1_66 BUFX2_6/gnd DFFSR_14/S FILL
XNAND3X1_63 AND2X2_6/A AOI22X1_9/B AND2X2_10/Y BUFX2_43/A NAND3X1_66/C DFFSR_23/S
+ NAND3X1
XFILL_0_NAND3X1_109 BUFX2_36/A DFFSR_8/S FILL
XFILL_6_OAI22X1_48 BUFX2_37/A DFFSR_81/S FILL
XFILL_41_DFFSR_92 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_4_NAND3X1_69 BUFX2_6/gnd DFFSR_14/S FILL
XOAI22X1_48 INVX1_354/Y OAI22X1_40/B INVX1_355/Y OAI22X1_40/D BUFX2_37/A NOR2X1_33/A
+ DFFSR_81/S OAI22X1
XFILL_5_OAI22X1_51 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_2_NAND2X1_145 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_3_NAND3X1_72 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_4_OAI22X1_54 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_8_OAI21X1_248 DFFSR_73/gnd DFFSR_57/S FILL
XDFFSR_190 BUFX2_32/A DFFSR_1/CLK DFFSR_185/R DFFSR_9/S DFFSR_190/D DFFSR_9/gnd DFFSR_9/S
+ DFFSR
XFILL_2_NAND3X1_75 BUFX2_35/A DFFSR_97/S FILL
XFILL_2_AND2X2_1 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_41_DFFSR_111 INVX1_8/gnd DFFSR_5/S FILL
XFILL_3_OAI22X1_57 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_14_DFFSR_82 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_25_DFFSR_42 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_4_DFFSR_187 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_8_DFFSR_49 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_1_NAND3X1_78 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_31_DFFSR_114 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_2_OAI22X1_60 INVX1_8/gnd DFFSR_5/S FILL
XFILL_21_DFFSR_117 INVX1_23/gnd DFFSR_91/S FILL
XFILL_0_OAI21X1_127 BUFX2_43/A DFFSR_23/S FILL
XFILL_0_NAND3X1_81 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_1_OAI22X1_63 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_4_NAND2X1_8 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_26_1_2 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_0_OAI22X1_66 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_11_DFFSR_120 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_49_DFFSR_99 BUFX2_35/A DFFSR_97/S FILL
XFILL_8_0_1 BUFX2_43/A DFFSR_97/S FILL
XFILL_1_INVX1_271 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_20_DFFSR_4 INVX1_4/gnd DFFSR_4/S FILL
XFILL_22_DFFSR_89 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_7_DFFSR_114 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_0_NAND2X1_241 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_5_DFFSR_96 INVX1_2/gnd DFFSR_1/S FILL
XINVX1_83 DFFSR_73/Q DFFSR_73/gnd INVX1_83/Y DFFSR_11/S INVX1
XFILL_33_DFFSR_49 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_48_DFFSR_145 INVX1_23/gnd DFFSR_186/S FILL
XFILL_6_2_2 BUFX2_35/A DFFSR_14/S FILL
XFILL_4_OAI22X1_7 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_38_DFFSR_148 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_4_BUFX2_5 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_8_NAND3X1_21 BUFX2_7/gnd DFFSR_81/S FILL
XINVX1_201 INVX1_201/A BUFX2_8/gnd INVX1_201/Y DFFSR_25/S INVX1
XFILL_4_DFFPOSX1_13 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_7_NAND3X1_24 BUFX2_37/A DFFSR_8/S FILL
XFILL_4_BUFX2_34 BUFX2_37/A DFFSR_81/S FILL
XFILL_28_DFFSR_151 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_1_NAND2X1_175 BUFX2_35/A DFFSR_14/S FILL
XFILL_18_DFFSR_154 BUFX2_36/A DFFSR_6/S FILL
XFILL_6_NAND3X1_27 BUFX2_37/A DFFSR_81/S FILL
XFILL_4_INVX1_198 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_35_8 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_5_NAND3X1_30 INVX1_94/gnd DFFSR_52/S FILL
XFILL_6_OAI22X1_12 INVX1_4/gnd DFFSR_51/S FILL
XNAND3X1_27 INVX1_233/A NAND3X1_23/Y NAND3X1_27/C BUFX2_37/A AOI22X1_4/D DFFSR_81/S
+ NAND3X1
XFILL_4_NAND3X1_33 INVX1_8/gnd DFFSR_7/S FILL
XFILL_30_DFFSR_96 INVX1_2/gnd DFFSR_1/S FILL
XFILL_41_DFFSR_56 INVX1_2/gnd DFFSR_51/S FILL
XFILL_5_OAI22X1_15 INVX1_4/gnd DFFSR_4/S FILL
XFILL_2_INVX1_90 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_3_NAND3X1_36 BUFX2_35/A DFFSR_97/S FILL
XDFFSR_154 DFFSR_154/Q CLKBUF1_11/Y DFFSR_154/R DFFSR_6/S DFFSR_154/D BUFX2_36/A DFFSR_6/S
+ DFFSR
XFILL_3_NOR2X1_33 BUFX2_37/A DFFSR_81/S FILL
XFILL_4_OAI22X1_18 BUFX2_8/gnd DFFSR_10/S FILL
XOAI22X1_12 INVX1_280/Y OAI22X1_7/B INVX1_279/Y OAI22X1_7/D INVX1_4/gnd NOR2X1_15/B
+ DFFSR_51/S OAI22X1
XFILL_8_OAI21X1_212 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_2_NAND3X1_39 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_2_NAND2X1_109 INVX1_94/gnd DFFSR_25/S FILL
XFILL_2_INVX1_415 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_3_OAI22X1_21 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_1_NAND3X1_42 BUFX2_43/A DFFSR_23/S FILL
XFILL_14_DFFSR_46 BUFX2_36/A DFFSR_6/S FILL
XFILL_4_DFFSR_151 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_2_OAI22X1_24 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_8_DFFSR_13 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_0_NAND3X1_45 BUFX2_35/A DFFSR_97/S FILL
XFILL_1_OAI22X1_27 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_45_DFFSR_182 INVX1_89/gnd DFFSR_36/S FILL
XFILL_35_DFFSR_185 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_23_DFFPOSX1_21 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_49_DFFSR_63 INVX1_94/gnd DFFSR_52/S FILL
XFILL_0_OAI22X1_30 INVX1_94/gnd DFFSR_25/S FILL
XFILL_25_DFFSR_188 INVX1_2/gnd DFFSR_1/S FILL
XFILL_1_INVX1_235 INVX1_4/gnd DFFSR_51/S FILL
XFILL_15_DFFSR_191 INVX1_23/gnd DFFSR_91/S FILL
XFILL_0_NAND2X1_205 BUFX2_36/A DFFSR_6/S FILL
XFILL_5_DFFSR_60 BUFX2_37/A DFFSR_8/S FILL
XFILL_22_DFFSR_53 DFFSR_71/gnd DFFSR_10/S FILL
XINVX1_47 INVX1_47/A BUFX2_17/gnd INVX1_47/Y DFFSR_7/S INVX1
XFILL_11_DFFSR_93 INVX1_2/gnd DFFSR_51/S FILL
XFILL_33_DFFSR_13 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_48_DFFSR_109 BUFX2_6/gnd DFFSR_14/S FILL
XINVX1_165 BUFX2_6/Y INVX1_23/gnd DFFSR_145/R DFFSR_186/S INVX1
XFILL_38_DFFSR_112 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_28_DFFSR_115 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_7_OAI21X1_242 BUFX2_35/A DFFSR_97/S FILL
XFILL_4_INVX1_162 INVX1_8/gnd DFFSR_7/S FILL
XFILL_1_NAND2X1_139 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_1_DFFSR_188 INVX1_2/gnd DFFSR_1/S FILL
XFILL_18_DFFSR_118 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_1_NAND2X1_9 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_41_DFFSR_20 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_30_DFFSR_60 BUFX2_37/A DFFSR_8/S FILL
XFILL_2_INVX1_54 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_8_OAI21X1_176 BUFX2_8/gnd DFFSR_25/S FILL
XDFFSR_118 INVX1_374/A CLKBUF1_3/Y DFFSR_113/R DFFSR_11/S DFFSR_118/D BUFX2_16/gnd
+ DFFSR_11/S DFFSR
XFILL_4_DFFSR_115 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_14_DFFSR_10 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_2_INVX1_379 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_45_DFFSR_146 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_1_OAI22X1_8 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_35_DFFSR_149 INVX1_23/gnd DFFSR_91/S FILL
XFILL_8_DFFSR_3 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_25_DFFSR_152 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_1_INVX1_199 BUFX2_35/A DFFSR_97/S FILL
XFILL_15_DFFSR_155 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_49_DFFSR_27 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_38_DFFSR_67 INVX1_2/gnd DFFSR_51/S FILL
XFILL_0_NAND2X1_169 BUFX2_36/A DFFSR_8/S FILL
XFILL_22_DFFSR_17 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_11_DFFSR_57 DFFSR_73/gnd DFFSR_57/S FILL
XINVX1_11 DFFSR_9/Q DFFSR_1/gnd INVX1_11/Y DFFSR_1/S INVX1
XFILL_5_DFFSR_24 BUFX2_16/gnd DFFSR_65/S FILL
XDFFSR_64 DFFSR_64/Q DFFSR_15/CLK DFFSR_61/R DFFSR_11/S DFFSR_64/D BUFX2_16/gnd DFFSR_11/S
+ DFFSR
XFILL_6_OR2X2_3 BUFX2_43/A DFFSR_23/S FILL
XFILL_0_NOR2X1_34 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_27_2_0 DFFSR_79/gnd DFFSR_36/S FILL
XINVX1_129 INVX1_344/A INVX1_89/gnd INVX1_129/Y DFFSR_36/S INVX1
XFILL_8_NAND3X1_122 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_1_DFFSR_152 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_12_DFFPOSX1_26 BUFX2_37/A DFFSR_81/S FILL
XFILL_25_4_1 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_4_NOR2X1_5 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_42_DFFSR_183 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_7_3_0 BUFX2_35/A DFFSR_97/S FILL
XFILL_7_OAI21X1_206 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_1_NAND2X1_103 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_32_DFFSR_7 INVX1_8/gnd DFFSR_7/S FILL
XFILL_46_DFFSR_74 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_4_INVX1_126 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_32_DFFSR_186 INVX1_23/gnd DFFSR_186/S FILL
XFILL_2_DFFSR_71 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_2_INVX1_18 INVX1_89/gnd DFFSR_2/S FILL
XFILL_22_DFFSR_189 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_30_DFFSR_24 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_5_5_1 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_22_DFFPOSX1_15 BUFX2_35/A DFFSR_14/S FILL
XFILL_19_DFFSR_64 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_8_OAI21X1_140 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_2_INVX1_343 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_8_DFFSR_186 INVX1_23/gnd DFFSR_186/S FILL
XFILL_6_XOR2X1_1 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_45_DFFSR_110 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_35_DFFSR_113 INVX1_23/gnd DFFSR_186/S FILL
XFILL_1_INVX1_163 INVX1_94/gnd DFFSR_52/S FILL
XFILL_25_DFFSR_116 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_38_DFFSR_31 BUFX2_35/A DFFSR_97/S FILL
XFILL_15_DFFSR_119 BUFX2_37/A DFFSR_81/S FILL
XFILL_27_DFFSR_71 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_0_NAND2X1_133 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_6_OAI21X1_236 BUFX2_5/gnd DFFSR_23/S FILL
XDFFSR_28 INVX1_32/A DFFSR_28/CLK DFFSR_31/R DFFSR_54/S DFFSR_28/D BUFX2_19/gnd DFFSR_54/S
+ DFFSR
XFILL_11_DFFSR_21 INVX1_2/gnd DFFSR_1/S FILL
XFILL_17_5 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_2_NOR3X1_2 INVX1_89/gnd DFFSR_2/S FILL
XFILL_1_DFFSR_116 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_8_OAI22X1_6 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_42_DFFSR_147 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_7_OAI21X1_170 INVX1_94/gnd DFFSR_25/S FILL
XFILL_33_1_2 INVX1_8/gnd DFFSR_7/S FILL
XFILL_32_DFFSR_150 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_46_DFFSR_38 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_35_DFFSR_78 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_22_DFFSR_153 BUFX2_36/A DFFSR_8/S FILL
XFILL_19_DFFSR_28 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_2_DFFSR_35 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_12_DFFSR_156 INVX1_23/gnd DFFSR_91/S FILL
XFILL_8_OAI21X1_104 INVX1_4/gnd DFFSR_51/S FILL
XFILL_2_INVX1_307 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_20_CLKBUF1_18 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_8_DFFSR_150 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_43_DFFSR_85 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_19_CLKBUF1_21 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_19_DFFSR_1 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_18_CLKBUF1_24 INVX1_23/gnd DFFSR_186/S FILL
XFILL_49_DFFSR_181 INVX1_23/gnd DFFSR_186/S FILL
XFILL_27_DFFSR_35 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_39_DFFSR_184 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_1_INVX1_127 INVX1_2/gnd DFFSR_1/S FILL
XFILL_16_DFFSR_75 INVX1_4/gnd DFFSR_51/S FILL
XFILL_3_BUFX2_2 BUFX2_43/A DFFSR_23/S FILL
XFILL_11_DFFPOSX1_20 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_7_NAND3X1_116 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_29_DFFSR_187 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_6_OAI21X1_200 BUFX2_37/A DFFSR_8/S FILL
XFILL_19_DFFSR_190 DFFSR_9/gnd DFFSR_9/S FILL
XOAI21X1_236 AOI21X1_33/Y AOI21X1_32/Y INVX1_252/Y BUFX2_5/gnd AOI21X1_39/A DFFSR_23/S
+ OAI21X1
XFILL_7_DFFSR_89 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_7_OAI21X1_134 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_42_DFFSR_111 INVX1_8/gnd DFFSR_5/S FILL
XFILL_24_DFFSR_82 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_35_DFFSR_42 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_32_DFFSR_114 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_5_DFFSR_187 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_22_DFFSR_117 INVX1_23/gnd DFFSR_91/S FILL
XFILL_1_DFFPOSX1_31 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_6_BUFX2_27 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_5_NAND2X1_8 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_12_DFFSR_120 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_2_INVX1_271 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_32_DFFSR_89 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_8_DFFSR_114 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_4_INVX1_83 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_43_DFFSR_49 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_5_OAI21X1_230 INVX1_23/gnd DFFSR_186/S FILL
XFILL_49_DFFSR_145 INVX1_23/gnd DFFSR_186/S FILL
XFILL_5_OAI22X1_7 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_39_DFFSR_148 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_29_DFFSR_151 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_16_DFFSR_39 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_39_5 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_19_DFFSR_154 BUFX2_36/A DFFSR_6/S FILL
XNAND3X1_1 BUFX2_14/Y AND2X2_11/A NAND3X1_1/C INVX1_94/gnd NAND3X1_1/Y DFFSR_25/S
+ NAND3X1
XNOR2X1_36 NOR2X1_36/A NOR2X1_36/B BUFX2_8/gnd NOR2X1_36/Y DFFSR_10/S NOR2X1
XFILL_6_OAI21X1_164 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_51_DFFSR_56 INVX1_2/gnd DFFSR_51/S FILL
XOAI21X1_200 INVX1_233/A AOI21X1_5/Y NAND3X1_23/Y BUFX2_37/A AOI21X1_23/C DFFSR_8/S
+ OAI21X1
XFILL_4_NOR2X1_33 BUFX2_37/A DFFSR_81/S FILL
XFILL_40_DFFSR_96 INVX1_2/gnd DFFSR_1/S FILL
XFILL_1_AND2X2_5 BUFX2_37/A DFFSR_81/S FILL
XFILL_6_NAND2X1_278 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_3_INVX1_415 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_24_DFFSR_46 BUFX2_36/A DFFSR_6/S FILL
XFILL_5_DFFSR_151 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_7_DFFSR_53 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_13_DFFSR_86 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_10_CLKBUF1_12 BUFX2_43/A DFFSR_23/S FILL
XFILL_46_DFFSR_182 INVX1_89/gnd DFFSR_36/S FILL
XFILL_36_DFFSR_185 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_4_OAI21X1_260 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_9_CLKBUF1_15 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_34_2_0 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_26_DFFSR_188 INVX1_2/gnd DFFSR_1/S FILL
XFILL_16_DFFSR_191 INVX1_23/gnd DFFSR_91/S FILL
XFILL_10_DFFSR_8 BUFX2_36/A DFFSR_8/S FILL
XFILL_8_CLKBUF1_18 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_2_INVX1_235 INVX1_4/gnd DFFSR_51/S FILL
XFILL_10_DFFPOSX1_14 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_6_NAND3X1_110 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_32_4_1 INVX1_8/gnd DFFSR_5/S FILL
XFILL_7_CLKBUF1_21 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_6_CLKBUF1_24 INVX1_23/gnd DFFSR_186/S FILL
XFILL_5_OAI21X1_194 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_32_DFFSR_53 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_4_INVX1_47 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_21_DFFSR_93 INVX1_2/gnd DFFSR_51/S FILL
XFILL_43_DFFSR_13 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_49_DFFSR_109 BUFX2_6/gnd DFFSR_14/S FILL
XCLKBUF1_24 INVX1_402/Y INVX1_23/gnd DFFSR_20/CLK DFFSR_186/S CLKBUF1
XFILL_39_DFFSR_112 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_29_DFFSR_115 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_3_BUFX2_38 BUFX2_37/A DFFSR_81/S FILL
XFILL_2_DFFSR_188 INVX1_2/gnd DFFSR_1/S FILL
XFILL_6_OAI21X1_128 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_19_DFFSR_118 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_2_NAND2X1_9 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_31_DFFSR_4 INVX1_4/gnd DFFSR_4/S FILL
XFILL_40_DFFSR_60 BUFX2_37/A DFFSR_8/S FILL
XFILL_1_INVX1_94 INVX1_94/gnd DFFSR_52/S FILL
XFILL_0_DFFPOSX1_25 BUFX2_19/gnd DFFSR_54/S FILL
XOAI21X1_164 BUFX2_3/Y INVX1_198/Y OAI21X1_164/C DFFSR_5/gnd DFFSR_164/D DFFSR_2/S
+ OAI21X1
XFILL_5_DFFSR_115 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_6_NAND2X1_242 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_24_DFFSR_10 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_7_DFFSR_17 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_3_INVX1_379 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_13_DFFSR_50 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_46_DFFSR_146 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_2_OAI22X1_8 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_36_DFFSR_149 INVX1_23/gnd DFFSR_91/S FILL
XNAND2X1_278 AND2X2_16/B AND2X2_16/A DFFSR_79/gnd NOR3X1_2/C DFFSR_45/S NAND2X1
XFILL_4_OAI21X1_224 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_26_DFFSR_152 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_2_INVX1_199 BUFX2_35/A DFFSR_97/S FILL
XFILL_48_DFFSR_67 INVX1_2/gnd DFFSR_51/S FILL
XFILL_16_DFFSR_155 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_32_DFFSR_17 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_21_DFFSR_57 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_4_DFFSR_64 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_10_DFFSR_97 BUFX2_35/A DFFSR_97/S FILL
XFILL_5_OAI21X1_158 BUFX2_43/A DFFSR_97/S FILL
XFILL_1_NOR2X1_34 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_40_1_2 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_0_INVX1_416 DFFSR_89/gnd DFFSR_92/S FILL
XNAND3X1_110 NAND2X1_231/Y NAND3X1_110/B AOI21X1_37/Y BUFX2_7/gnd NAND2X1_233/B DFFSR_54/S
+ NAND3X1
XFILL_2_DFFSR_152 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_43_DFFSR_183 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_5_NAND2X1_272 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_33_DFFSR_186 INVX1_23/gnd DFFSR_186/S FILL
XFILL_23_DFFSR_189 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_40_DFFSR_24 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_1_INVX1_58 BUFX2_16/gnd DFFSR_65/S FILL
XOAI21X1_128 BUFX2_19/Y INVX1_144/Y OAI21X1_128/C BUFX2_8/gnd DFFSR_128/D DFFSR_25/S
+ OAI21X1
XFILL_29_DFFSR_64 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_3_OAI21X1_254 INVX1_23/gnd DFFSR_91/S FILL
XFILL_6_NAND2X1_206 BUFX2_43/A DFFSR_97/S FILL
XFILL_3_INVX1_343 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_13_DFFSR_14 BUFX2_35/A DFFSR_14/S FILL
XFILL_5_NAND3X1_104 INVX1_23/gnd DFFSR_186/S FILL
XFILL_46_DFFSR_110 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_9_DFFSR_186 INVX1_23/gnd DFFSR_186/S FILL
XFILL_36_DFFSR_113 INVX1_23/gnd DFFSR_186/S FILL
XNAND2X1_242 NOR2X1_29/Y NOR2X1_28/Y BUFX2_19/gnd NAND2X1_242/Y DFFSR_52/S NAND2X1
XFILL_4_OAI21X1_188 INVX1_89/gnd DFFSR_2/S FILL
XFILL_26_DFFSR_116 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_48_DFFSR_31 BUFX2_35/A DFFSR_97/S FILL
XFILL_16_DFFSR_119 BUFX2_37/A DFFSR_81/S FILL
XFILL_2_INVX1_163 INVX1_94/gnd DFFSR_52/S FILL
XFILL_37_DFFSR_71 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_10_DFFSR_61 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_4_DFFSR_28 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_5_OAI21X1_122 INVX1_94/gnd DFFSR_25/S FILL
XFILL_21_DFFSR_21 INVX1_2/gnd DFFSR_1/S FILL
XFILL_3_NOR2X1_9 BUFX2_43/A DFFSR_97/S FILL
XFILL_21_2 INVX1_94/gnd DFFSR_52/S FILL
XFILL_0_INVX1_380 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_9_OAI22X1_6 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_43_DFFSR_147 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_2_DFFSR_116 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_33_DFFSR_150 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_45_DFFSR_78 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_5_NAND2X1_236 INVX1_2/gnd DFFSR_1/S FILL
XFILL_23_DFFSR_153 BUFX2_36/A DFFSR_8/S FILL
XFILL_18_DFFSR_68 BUFX2_35/A DFFSR_14/S FILL
XFILL_29_DFFSR_28 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_4_NAND3X1_134 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_1_INVX1_22 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_1_DFFSR_75 INVX1_4/gnd DFFSR_51/S FILL
XFILL_3_OAI21X1_218 INVX1_23/gnd DFFSR_186/S FILL
XFILL_13_DFFSR_156 INVX1_23/gnd DFFSR_91/S FILL
XFILL_3_INVX1_307 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_6_NAND2X1_170 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_5_XOR2X1_5 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_0_BUFX2_13 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_21_DFFPOSX1_3 DFFSR_71/gnd DFFSR_45/S FILL
XNAND2X1_206 AOI22X1_7/A AOI22X1_7/B BUFX2_43/A NAND3X1_73/B DFFSR_97/S NAND2X1
XFILL_9_DFFSR_150 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_43_DFFSR_7 INVX1_8/gnd DFFSR_7/S FILL
XFILL_20_DFFPOSX1_6 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_50_DFFSR_181 INVX1_23/gnd DFFSR_186/S FILL
XFILL_4_OAI21X1_152 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_18_DFFPOSX1_27 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_19_DFFPOSX1_9 BUFX2_37/A DFFSR_8/S FILL
XFILL_37_DFFSR_35 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_40_DFFSR_184 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_9_DFFSR_82 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_2_INVX1_127 INVX1_2/gnd DFFSR_1/S FILL
XFILL_26_DFFSR_75 INVX1_4/gnd DFFSR_51/S FILL
XFILL_30_DFFSR_187 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_20_DFFSR_190 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_4_NAND2X1_266 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_10_DFFSR_25 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_0_INVX1_344 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_4_6 INVX1_23/gnd DFFSR_91/S FILL
XFILL_5_NAND2X1_200 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_43_DFFSR_111 INVX1_8/gnd DFFSR_5/S FILL
XFILL_2_OAI21X1_248 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_34_DFFSR_82 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_41_2_0 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_45_DFFSR_42 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_33_DFFSR_114 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_6_DFFSR_187 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_23_DFFSR_117 INVX1_23/gnd DFFSR_91/S FILL
XFILL_1_DFFSR_39 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_6_NAND2X1_8 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_18_DFFSR_32 INVX1_2/gnd DFFSR_1/S FILL
XFILL_39_4_1 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_13_DFFSR_120 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_6_NAND2X1_134 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_3_OAI21X1_182 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_3_INVX1_271 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_42_DFFSR_89 DFFSR_89/gnd DFFSR_92/S FILL
XXOR2X1_9 NOR2X1_1/B NOR2X1_1/A BUFX2_19/gnd XOR2X1_9/Y DFFSR_52/S XOR2X1
XFILL_11_XOR2X1_2 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_9_DFFSR_114 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_50_DFFSR_145 INVX1_23/gnd DFFSR_186/S FILL
XFILL_4_OAI21X1_116 INVX1_89/gnd DFFSR_2/S FILL
XFILL_6_OAI22X1_7 DFFSR_5/gnd DFFSR_5/S FILL
XNAND2X1_170 DFFSR_11/S NAND2X1_170/B BUFX2_16/gnd OAI21X1_170/C DFFSR_11/S NAND2X1
XFILL_40_DFFSR_148 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_9_DFFSR_46 BUFX2_36/A DFFSR_6/S FILL
XFILL_30_DFFSR_151 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_26_DFFSR_39 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_15_DFFSR_79 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_43_2 INVX1_4/gnd DFFSR_4/S FILL
XFILL_4_NAND2X1_230 BUFX2_36/A DFFSR_6/S FILL
XFILL_20_DFFSR_154 BUFX2_36/A DFFSR_6/S FILL
XFILL_10_DFFSR_157 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_5_NOR2X1_33 BUFX2_37/A DFFSR_81/S FILL
XFILL_0_INVX1_308 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_3_NAND3X1_128 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_50_DFFSR_96 INVX1_2/gnd DFFSR_1/S FILL
XFILL_30_DFFSR_1 DFFSR_1/gnd DFFSR_1/S FILL
XINVX1_418 BUFX2_29/A DFFSR_3/gnd INVX1_418/Y DFFSR_4/S INVX1
XFILL_2_OAI21X1_212 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_4_INVX1_415 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_34_DFFSR_46 BUFX2_36/A DFFSR_6/S FILL
XFILL_6_DFFSR_151 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_5_NAND2X1_164 INVX1_8/gnd DFFSR_5/S FILL
XFILL_23_DFFSR_86 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_6_DFFSR_93 INVX1_2/gnd DFFSR_51/S FILL
XFILL_47_DFFSR_182 INVX1_89/gnd DFFSR_36/S FILL
XFILL_37_DFFSR_185 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_3_OAI21X1_146 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_17_DFFPOSX1_21 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_5_BUFX2_31 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_47_1_2 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_27_DFFSR_188 INVX1_2/gnd DFFSR_1/S FILL
XFILL_17_DFFSR_191 INVX1_23/gnd DFFSR_91/S FILL
XFILL_3_INVX1_235 INVX1_4/gnd DFFSR_51/S FILL
XFILL_9_DFFPOSX1_3 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_9_AOI21X1_23 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_42_DFFSR_53 DFFSR_71/gnd DFFSR_10/S FILL
XNAND2X1_134 DFFSR_45/S NAND2X1_70/B DFFSR_79/gnd OAI21X1_134/C DFFSR_36/S NAND2X1
XFILL_3_INVX1_87 INVX1_89/gnd DFFSR_36/S FILL
XFILL_31_DFFSR_93 INVX1_2/gnd DFFSR_51/S FILL
XFILL_8_DFFPOSX1_6 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_3_NAND2X1_260 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_50_DFFSR_109 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_8_AOI21X1_26 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_7_DFFPOSX1_9 BUFX2_37/A DFFSR_8/S FILL
XFILL_27_DFFPOSX1_10 INVX1_8/gnd DFFSR_5/S FILL
XFILL_15_DFFSR_43 INVX1_94/gnd DFFSR_25/S FILL
XFILL_9_DFFSR_10 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_7_AOI21X1_29 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_40_DFFSR_112 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_30_DFFSR_115 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_6_AOI21X1_32 BUFX2_43/A DFFSR_23/S FILL
XFILL_15_0_0 BUFX2_37/A DFFSR_81/S FILL
XFILL_3_DFFSR_188 INVX1_2/gnd DFFSR_1/S FILL
XFILL_1_OAI21X1_242 BUFX2_35/A DFFSR_97/S FILL
XFILL_4_NAND2X1_194 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_5_AOI21X1_35 INVX1_94/gnd DFFSR_25/S FILL
XFILL_20_DFFSR_118 BUFX2_16/gnd DFFSR_11/S FILL
XAOI21X1_32 AOI21X1_32/A AOI21X1_32/B XOR2X1_8/B BUFX2_43/A AOI21X1_32/Y DFFSR_23/S
+ AOI21X1
XFILL_10_DFFSR_121 BUFX2_36/A DFFSR_6/S FILL
XFILL_4_AOI21X1_38 BUFX2_36/A DFFSR_8/S FILL
XFILL_13_2_1 BUFX2_36/A DFFSR_8/S FILL
XFILL_3_NAND2X1_9 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_3_AOI21X1_41 BUFX2_35/A DFFSR_14/S FILL
XFILL_50_DFFSR_60 BUFX2_37/A DFFSR_8/S FILL
XINVX1_382 INVX1_134/A BUFX2_19/gnd INVX1_382/Y DFFSR_54/S INVX1
XFILL_0_INVX1_272 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_0_AND2X2_9 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_11_4_2 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_2_OAI21X1_176 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_34_DFFSR_10 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_5_NAND2X1_128 INVX1_89/gnd DFFSR_2/S FILL
XFILL_2_AOI21X1_44 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_6_DFFSR_57 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_12_DFFSR_90 INVX1_2/gnd DFFSR_1/S FILL
XFILL_23_DFFSR_50 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_47_DFFSR_146 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_6_DFFSR_115 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_1_AOI21X1_47 BUFX2_43/A DFFSR_23/S FILL
XFILL_3_OAI22X1_8 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_37_DFFSR_149 INVX1_23/gnd DFFSR_91/S FILL
XBUFX2_35 BUFX2_35/A BUFX2_35/A BUFX2_35/Y DFFSR_14/S BUFX2
XFILL_27_DFFSR_152 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_3_INVX1_199 BUFX2_35/A DFFSR_97/S FILL
XFILL_3_OAI21X1_110 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_17_DFFSR_155 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_48_7 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_8_OAI21X1_74 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_3_INVX1_51 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_7_OAI21X1_77 INVX1_89/gnd DFFSR_36/S FILL
XFILL_6_NAND2X1_95 INVX1_89/gnd DFFSR_36/S FILL
XFILL_42_DFFSR_17 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_20_DFFSR_97 BUFX2_35/A DFFSR_97/S FILL
XFILL_3_NAND2X1_224 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_2_NOR2X1_34 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_31_DFFSR_57 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_5_NAND2X1_98 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_6_OAI21X1_80 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_1_INVX1_416 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_5_OAI21X1_83 INVX1_94/gnd DFFSR_52/S FILL
XNAND2X1_95 BUFX2_22/Y DFFSR_87/Q INVX1_89/gnd NAND2X1_95/Y DFFSR_36/S NAND2X1
XFILL_2_BUFX2_42 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_3_DFFSR_152 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_2_NAND3X1_122 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_4_OAI21X1_86 INVX1_4/gnd DFFSR_51/S FILL
XOAI21X1_80 BUFX2_17/Y INVX1_90/Y NAND2X1_80/Y DFFSR_73/gnd DFFSR_80/D DFFSR_11/S
+ OAI21X1
XFILL_44_DFFSR_183 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_3_OAI21X1_89 BUFX2_35/A DFFSR_14/S FILL
XFILL_1_OAI21X1_206 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_34_DFFSR_186 INVX1_23/gnd DFFSR_186/S FILL
XFILL_4_NAND2X1_158 BUFX2_35/A DFFSR_97/S FILL
XFILL_2_OAI21X1_92 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_21_DFFSR_8 BUFX2_36/A DFFSR_8/S FILL
XFILL_1_OAI21X1_95 INVX1_89/gnd DFFSR_36/S FILL
XFILL_24_DFFSR_189 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_0_INVX1_236 INVX1_8/gnd DFFSR_7/S FILL
XINVX1_346 DFFSR_98/Q DFFSR_1/gnd INVX1_346/Y DFFSR_1/S INVX1
XFILL_0_OAI21X1_98 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_0_INVX1_98 INVX1_4/gnd DFFSR_4/S FILL
XFILL_50_DFFSR_24 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_39_DFFSR_64 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_16_DFFPOSX1_15 BUFX2_35/A DFFSR_14/S FILL
XFILL_2_OAI21X1_140 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_23_DFFSR_14 BUFX2_35/A DFFSR_14/S FILL
XFILL_5_BUFX2_9 BUFX2_37/A DFFSR_8/S FILL
XFILL_12_DFFSR_54 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_1_AOI21X1_11 INVX1_8/gnd DFFSR_5/S FILL
XFILL_6_DFFSR_21 INVX1_2/gnd DFFSR_1/S FILL
XFILL_1_0_2 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_0_AOI21X1_14 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_47_DFFSR_110 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_37_DFFSR_113 INVX1_23/gnd DFFSR_186/S FILL
XFILL_5_NOR2X1_2 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_2_NAND2X1_254 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_27_DFFSR_116 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_9_OAI21X1_35 INVX1_8/gnd DFFSR_5/S FILL
XFILL_0_DFFSR_189 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_42_DFFSR_4 INVX1_4/gnd DFFSR_4/S FILL
XFILL_17_DFFSR_119 BUFX2_37/A DFFSR_81/S FILL
XFILL_3_INVX1_163 INVX1_94/gnd DFFSR_52/S FILL
XFILL_47_DFFSR_71 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_8_OAI21X1_38 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_7_OAI21X1_41 INVX1_8/gnd DFFSR_7/S FILL
XFILL_6_NAND2X1_59 INVX1_2/gnd DFFSR_1/S FILL
XFILL_3_DFFSR_68 BUFX2_35/A DFFSR_14/S FILL
XFILL_0_OAI21X1_236 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_20_DFFSR_61 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_6_DFFPOSX1_26 BUFX2_37/A DFFSR_81/S FILL
XFILL_5_NAND2X1_62 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_31_DFFSR_21 INVX1_2/gnd DFFSR_1/S FILL
XFILL_3_INVX1_15 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_6_OAI21X1_44 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_3_NAND2X1_188 INVX1_8/gnd DFFSR_7/S FILL
XFILL_48_2_0 DFFSR_9/gnd DFFSR_9/S FILL
XNAND2X1_59 DFFSR_1/S INVX1_58/A INVX1_2/gnd OAI21X1_59/C DFFSR_1/S NAND2X1
XOAI21X1_44 DFFSR_45/S INVX1_50/Y OAI21X1_44/C DFFSR_71/gnd DFFSR_44/D DFFSR_45/S
+ OAI21X1
XFILL_1_INVX1_380 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_5_OAI21X1_47 INVX1_89/gnd DFFSR_2/S FILL
XFILL_4_NAND2X1_65 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_44_DFFSR_147 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_3_NAND2X1_68 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_3_DFFSR_116 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_0_OAI22X1_9 INVX1_8/gnd DFFSR_5/S FILL
XFILL_4_OAI21X1_50 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_46_4_1 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_1_OAI21X1_170 INVX1_94/gnd DFFSR_25/S FILL
XFILL_4_NAND2X1_122 INVX1_94/gnd DFFSR_25/S FILL
XFILL_34_DFFSR_150 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_2_NAND2X1_71 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_3_OAI21X1_53 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_1_NAND2X1_74 INVX1_2/gnd DFFSR_1/S FILL
XFILL_2_OAI21X1_56 INVX1_2/gnd DFFSR_51/S FILL
XFILL_28_DFFSR_68 BUFX2_35/A DFFSR_14/S FILL
XFILL_24_DFFSR_153 BUFX2_36/A DFFSR_8/S FILL
XFILL_39_DFFSR_28 BUFX2_19/gnd DFFSR_54/S FILL
XINVX1_310 DFFSR_30/Q DFFSR_79/gnd INVX1_310/Y DFFSR_36/S INVX1
XFILL_0_NAND2X1_77 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_0_INVX1_62 INVX1_89/gnd DFFSR_2/S FILL
XFILL_1_OAI21X1_59 INVX1_4/gnd DFFSR_51/S FILL
XFILL_0_INVX1_200 INVX1_4/gnd DFFSR_4/S FILL
XFILL_14_DFFSR_156 INVX1_23/gnd DFFSR_91/S FILL
XFILL_0_OAI21X1_62 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_1_NAND2X1_284 INVX1_8/gnd DFFSR_5/S FILL
XFILL_4_INVX1_307 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_12_DFFSR_18 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_2_OAI21X1_104 INVX1_4/gnd DFFSR_51/S FILL
XFILL_12_5_0 BUFX2_36/A DFFSR_6/S FILL
XFILL_0_DFFSR_153 BUFX2_36/A DFFSR_8/S FILL
XNOR2X1_6 AND2X2_3/B AND2X2_3/A BUFX2_17/gnd NOR2X1_6/Y DFFSR_57/S NOR2X1
XFILL_2_NAND2X1_218 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_47_DFFSR_35 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_41_DFFSR_184 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_3_INVX1_127 INVX1_2/gnd DFFSR_1/S FILL
XFILL_36_DFFSR_75 INVX1_4/gnd DFFSR_51/S FILL
XFILL_1_NAND3X1_116 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_31_DFFSR_187 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_6_NAND2X1_23 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_21_DFFSR_190 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_3_DFFSR_32 INVX1_2/gnd DFFSR_1/S FILL
XFILL_3_NAND2X1_152 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_0_OAI21X1_200 BUFX2_37/A DFFSR_8/S FILL
XFILL_20_DFFSR_25 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_5_NAND2X1_26 DFFSR_1/gnd DFFSR_9/S FILL
XNAND2X1_23 DFFSR_6/S DFFSR_15/Q BUFX2_5/gnd OAI21X1_23/C DFFSR_6/S NAND2X1
XFILL_1_INVX1_344 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_4_NAND2X1_29 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_5_OAI21X1_11 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_4_OAI21X1_14 BUFX2_43/A DFFSR_23/S FILL
XDFFPOSX1_26 AND2X2_10/B CLKBUF1_16/Y XOR2X1_15/Y BUFX2_37/A DFFSR_81/S DFFPOSX1
XFILL_9_DFFSR_7 INVX1_8/gnd DFFSR_7/S FILL
XFILL_3_NAND2X1_32 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_1_OAI21X1_134 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_3_OAI21X1_17 INVX1_8/gnd DFFSR_5/S FILL
XFILL_44_DFFSR_111 INVX1_8/gnd DFFSR_5/S FILL
XFILL_2_NAND2X1_35 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_44_DFFSR_82 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_2_OAI21X1_20 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_9_NAND3X1_91 BUFX2_43/A DFFSR_97/S FILL
XFILL_34_DFFSR_114 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_1_NAND2X1_38 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_7_DFFSR_187 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_24_DFFSR_117 INVX1_23/gnd DFFSR_91/S FILL
XFILL_8_NAND3X1_94 BUFX2_35/A DFFSR_97/S FILL
XFILL_1_OAI21X1_23 BUFX2_5/gnd DFFSR_23/S FILL
XAOI21X1_2 NAND3X1_4/B NAND3X1_4/A NOR2X1_3/Y INVX1_94/gnd AOI21X1_2/Y DFFSR_52/S
+ AOI21X1
XFILL_0_NAND2X1_41 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_0_INVX1_164 INVX1_23/gnd DFFSR_91/S FILL
XFILL_7_NAND3X1_97 BUFX2_35/A DFFSR_97/S FILL
XFILL_0_INVX1_26 BUFX2_43/A DFFSR_23/S FILL
XFILL_0_DFFSR_79 DFFSR_79/gnd DFFSR_36/S FILL
XINVX1_274 DFFSR_10/Q INVX1_8/gnd INVX1_274/Y DFFSR_5/S INVX1
XFILL_17_DFFSR_72 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_0_OAI21X1_26 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_28_DFFSR_32 INVX1_2/gnd DFFSR_1/S FILL
XFILL_14_DFFSR_120 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_1_NAND2X1_248 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_4_INVX1_271 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_4_XOR2X1_9 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_22_0_0 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_5_DFFPOSX1_20 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_7_OAI22X1_7 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_41_DFFSR_148 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_0_DFFSR_117 INVX1_23/gnd DFFSR_91/S FILL
XFILL_2_NAND2X1_182 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_31_DFFSR_151 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_20_2_1 INVX1_94/gnd DFFSR_52/S FILL
XFILL_36_DFFSR_39 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_25_DFFSR_79 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_8_DFFSR_86 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_2_1_0 INVX1_23/gnd DFFSR_186/S FILL
XFILL_3_AOI22X1_10 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_21_DFFSR_154 BUFX2_36/A DFFSR_6/S FILL
XFILL_18_4_2 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_0_OAI21X1_164 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_0_3_1 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_2_AOI22X1_13 INVX1_23/gnd DFFSR_186/S FILL
XFILL_11_DFFSR_157 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_3_NAND2X1_116 INVX1_89/gnd DFFSR_36/S FILL
XFILL_6_NOR2X1_33 BUFX2_37/A DFFSR_81/S FILL
XFILL_1_INVX1_308 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_10_OAI22X1_37 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_44_DFFSR_46 BUFX2_36/A DFFSR_6/S FILL
XFILL_7_DFFSR_151 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_0_NAND2X1_278 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_33_DFFSR_86 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_24_DFFPOSX1_28 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_48_DFFSR_182 INVX1_89/gnd DFFSR_36/S FILL
XFILL_38_DFFSR_185 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_0_INVX1_128 INVX1_23/gnd DFFSR_91/S FILL
XFILL_9_OAI22X1_40 BUFX2_37/A DFFSR_8/S FILL
XINVX1_238 INVX1_238/A BUFX2_37/A INVX1_238/Y DFFSR_81/S INVX1
XFILL_8_NAND3X1_58 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_0_DFFSR_43 INVX1_94/gnd DFFSR_25/S FILL
XFILL_17_DFFSR_36 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_1_NAND2X1_212 INVX1_23/gnd DFFSR_186/S FILL
XFILL_8_OAI22X1_43 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_7_NAND3X1_61 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_28_DFFSR_188 INVX1_2/gnd DFFSR_1/S FILL
XFILL_18_DFFSR_191 INVX1_23/gnd DFFSR_91/S FILL
XFILL_6_NAND3X1_64 BUFX2_35/A DFFSR_14/S FILL
XFILL_7_OAI22X1_46 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_5_NAND3X1_67 BUFX2_6/gnd DFFSR_14/S FILL
XNAND3X1_64 INVX1_249/Y INVX1_248/Y NAND3X1_66/C BUFX2_35/A NAND3X1_64/Y DFFSR_14/S
+ NAND3X1
XFILL_0_NAND3X1_110 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_6_OAI22X1_49 INVX1_94/gnd DFFSR_25/S FILL
XFILL_10_XOR2X1_6 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_4_NAND3X1_70 BUFX2_35/A DFFSR_14/S FILL
XFILL_5_OAI22X1_52 INVX1_94/gnd DFFSR_25/S FILL
XFILL_41_DFFSR_93 INVX1_2/gnd DFFSR_51/S FILL
XFILL_8_OAI21X1_249 DFFSR_89/gnd DFFSR_186/S FILL
XDFFSR_191 BUFX2_33/A DFFSR_20/CLK DFFSR_185/R DFFSR_91/S DFFSR_191/D INVX1_23/gnd
+ DFFSR_91/S DFFSR
XFILL_2_NAND2X1_146 INVX1_23/gnd DFFSR_91/S FILL
XFILL_3_NAND3X1_73 BUFX2_43/A DFFSR_23/S FILL
XOAI22X1_49 INVX1_356/Y OAI22X1_38/D INVX1_357/Y OAI22X1_49/D INVX1_94/gnd NOR2X1_34/B
+ DFFSR_25/S OAI22X1
XFILL_4_OAI22X1_55 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_2_NAND3X1_76 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_2_AND2X2_2 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_14_DFFSR_83 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_25_DFFSR_43 INVX1_94/gnd DFFSR_25/S FILL
XFILL_3_OAI22X1_58 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_41_DFFSR_112 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_8_DFFSR_50 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_31_DFFSR_115 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_1_NAND3X1_79 BUFX2_36/A DFFSR_6/S FILL
XFILL_2_OAI22X1_61 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_4_DFFSR_188 INVX1_2/gnd DFFSR_1/S FILL
XFILL_0_NAND3X1_82 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_1_OAI22X1_64 INVX1_94/gnd DFFSR_25/S FILL
XFILL_21_DFFSR_118 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_11_DFFSR_121 BUFX2_36/A DFFSR_6/S FILL
XFILL_0_OAI21X1_128 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_4_NAND2X1_9 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_0_OAI22X1_67 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_8_0_2 BUFX2_43/A DFFSR_97/S FILL
XFILL_1_INVX1_272 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_20_DFFSR_5 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_5_DFFSR_97 BUFX2_35/A DFFSR_97/S FILL
XFILL_0_NAND2X1_242 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_44_DFFSR_10 DFFSR_71/gnd DFFSR_10/S FILL
XINVX1_84 DFFSR_74/Q DFFSR_9/gnd INVX1_84/Y DFFSR_9/S INVX1
XFILL_33_DFFSR_50 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_48_DFFSR_146 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_7_DFFSR_115 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_4_OAI22X1_8 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_22_DFFSR_90 INVX1_2/gnd DFFSR_1/S FILL
XFILL_38_DFFSR_149 INVX1_23/gnd DFFSR_91/S FILL
XFILL_4_BUFX2_6 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_8_NAND3X1_22 BUFX2_37/A DFFSR_81/S FILL
XFILL_4_BUFX2_35 BUFX2_35/A DFFSR_14/S FILL
XINVX1_202 BUFX2_7/Y BUFX2_37/A DFFSR_162/R DFFSR_81/S INVX1
XFILL_7_NAND3X1_25 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_4_DFFPOSX1_14 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_4_INVX1_199 BUFX2_35/A DFFSR_97/S FILL
XFILL_28_DFFSR_152 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_6_NAND3X1_28 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_1_NAND2X1_176 INVX1_94/gnd DFFSR_25/S FILL
XFILL_7_OAI22X1_10 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_18_DFFSR_155 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_5_NAND3X1_31 INVX1_94/gnd DFFSR_52/S FILL
XFILL_41_DFFSR_1 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_6_OAI22X1_13 DFFSR_3/gnd DFFSR_65/S FILL
XNAND3X1_28 INVX1_233/Y NAND3X1_23/Y NAND3X1_27/C BUFX2_7/gnd AOI21X1_7/A DFFSR_81/S
+ NAND3X1
XFILL_4_NAND3X1_34 INVX1_2/gnd DFFSR_1/S FILL
XFILL_5_OAI22X1_16 INVX1_4/gnd DFFSR_4/S FILL
XFILL_30_DFFSR_97 BUFX2_35/A DFFSR_97/S FILL
XFILL_3_NAND3X1_37 BUFX2_43/A DFFSR_97/S FILL
XFILL_2_INVX1_91 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_3_NOR2X1_34 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_4_OAI22X1_19 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_41_DFFSR_57 DFFSR_73/gnd DFFSR_57/S FILL
XOAI22X1_13 INVX1_282/Y OAI22X1_9/B INVX1_281/Y OAI22X1_9/D DFFSR_3/gnd NOR2X1_16/B
+ DFFSR_65/S OAI22X1
XFILL_2_INVX1_416 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_2_NAND3X1_40 BUFX2_43/A DFFSR_23/S FILL
XFILL_8_OAI21X1_213 BUFX2_36/A DFFSR_6/S FILL
XDFFSR_155 INVX1_184/A CLKBUF1_11/Y DFFSR_155/R DFFSR_54/S DFFSR_155/D BUFX2_7/gnd
+ DFFSR_54/S DFFSR
XFILL_2_NAND2X1_110 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_8_DFFSR_14 BUFX2_35/A DFFSR_14/S FILL
XFILL_4_DFFSR_152 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_14_DFFSR_47 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_3_OAI22X1_22 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_45_DFFSR_183 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_1_NAND3X1_43 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_2_OAI22X1_25 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_35_DFFSR_186 INVX1_23/gnd DFFSR_186/S FILL
XFILL_0_NAND3X1_46 BUFX2_35/A DFFSR_97/S FILL
XFILL_1_OAI22X1_28 INVX1_94/gnd DFFSR_25/S FILL
XFILL_23_DFFPOSX1_22 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_0_OAI22X1_31 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_25_DFFSR_189 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_1_INVX1_236 INVX1_8/gnd DFFSR_7/S FILL
XFILL_49_DFFSR_64 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_33_DFFSR_14 BUFX2_35/A DFFSR_14/S FILL
XFILL_0_NAND2X1_206 BUFX2_43/A DFFSR_97/S FILL
XFILL_5_DFFSR_61 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_22_DFFSR_54 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_19_5_0 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_11_DFFSR_94 BUFX2_16/gnd DFFSR_65/S FILL
XINVX1_48 INVX1_48/A BUFX2_16/gnd INVX1_48/Y DFFSR_65/S INVX1
XFILL_48_DFFSR_110 DFFSR_73/gnd DFFSR_57/S FILL
XINVX1_166 DFFSR_146/Q DFFSR_89/gnd INVX1_166/Y DFFSR_92/S INVX1
XFILL_38_DFFSR_113 INVX1_23/gnd DFFSR_186/S FILL
XFILL_1_NAND2X1_140 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_28_DFFSR_116 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_1_DFFSR_189 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_7_OAI21X1_243 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_18_DFFSR_119 BUFX2_37/A DFFSR_81/S FILL
XFILL_4_INVX1_163 INVX1_94/gnd DFFSR_52/S FILL
XFILL_30_DFFSR_61 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_2_INVX1_55 BUFX2_36/A DFFSR_8/S FILL
XFILL_41_DFFSR_21 INVX1_2/gnd DFFSR_1/S FILL
XDFFSR_119 INVX1_134/A CLKBUF1_6/Y DFFSR_113/R DFFSR_81/S DFFSR_119/D BUFX2_37/A DFFSR_81/S
+ DFFSR
XFILL_8_OAI21X1_177 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_2_INVX1_380 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_14_DFFSR_11 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_45_DFFSR_147 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_4_DFFSR_116 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_1_OAI22X1_9 INVX1_8/gnd DFFSR_5/S FILL
XFILL_0_NAND3X1_10 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_35_DFFSR_150 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_8_DFFSR_4 INVX1_4/gnd DFFSR_4/S FILL
XFILL_38_DFFSR_68 BUFX2_35/A DFFSR_14/S FILL
XFILL_25_DFFSR_153 BUFX2_36/A DFFSR_8/S FILL
XFILL_49_DFFSR_28 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_1_INVX1_200 INVX1_4/gnd DFFSR_4/S FILL
XFILL_15_DFFSR_156 INVX1_23/gnd DFFSR_91/S FILL
XFILL_29_0_0 INVX1_89/gnd DFFSR_2/S FILL
XFILL_5_DFFSR_25 BUFX2_8/gnd DFFSR_25/S FILL
XINVX1_12 DFFSR_10/Q DFFSR_71/gnd INVX1_12/Y DFFSR_45/S INVX1
XFILL_22_DFFSR_18 DFFSR_9/gnd DFFSR_9/S FILL
XDFFSR_65 DFFSR_65/Q CLKBUF1_3/Y DFFSR_68/R DFFSR_65/S DFFSR_65/D DFFSR_3/gnd DFFSR_65/S
+ DFFSR
XFILL_0_NAND2X1_170 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_0_NOR2X1_35 INVX1_94/gnd DFFSR_52/S FILL
XFILL_27_2_1 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_11_DFFSR_58 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_9_1_0 BUFX2_43/A DFFSR_23/S FILL
XINVX1_130 DFFSR_115/Q BUFX2_36/A INVX1_130/Y DFFSR_6/S INVX1
XFILL_1_DFFSR_153 BUFX2_36/A DFFSR_8/S FILL
XFILL_25_4_2 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_12_DFFPOSX1_27 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_8_NAND3X1_123 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_4_NOR2X1_6 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_32_DFFSR_8 BUFX2_36/A DFFSR_8/S FILL
XFILL_7_OAI21X1_207 BUFX2_37/A DFFSR_8/S FILL
XFILL_42_DFFSR_184 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_4_INVX1_127 INVX1_2/gnd DFFSR_1/S FILL
XFILL_1_NAND2X1_104 INVX1_4/gnd DFFSR_51/S FILL
XFILL_46_DFFSR_75 INVX1_4/gnd DFFSR_51/S FILL
XFILL_7_3_1 BUFX2_35/A DFFSR_97/S FILL
XFILL_32_DFFSR_187 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_22_DFFSR_190 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_2_INVX1_19 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_5_5_2 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_30_DFFSR_25 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_2_DFFSR_72 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_19_DFFSR_65 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_22_DFFPOSX1_16 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_8_OAI21X1_141 INVX1_94/gnd DFFSR_52/S FILL
XFILL_2_INVX1_344 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_1_BUFX2_10 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_6_XOR2X1_2 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_45_DFFSR_111 INVX1_8/gnd DFFSR_5/S FILL
XFILL_35_DFFSR_114 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_8_DFFSR_187 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_25_DFFSR_117 INVX1_23/gnd DFFSR_91/S FILL
XFILL_1_INVX1_164 INVX1_23/gnd DFFSR_91/S FILL
XFILL_27_DFFSR_72 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_38_DFFSR_32 INVX1_2/gnd DFFSR_1/S FILL
XFILL_15_DFFSR_120 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_6_OAI21X1_237 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_11_DFFSR_22 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_0_NAND2X1_134 DFFSR_79/gnd DFFSR_36/S FILL
XDFFSR_29 INVX1_33/A DFFSR_15/CLK DFFSR_31/R DFFSR_4/S DFFSR_29/D INVX1_4/gnd DFFSR_4/S
+ DFFSR
XFILL_8_OAI22X1_7 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_42_DFFSR_148 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_1_DFFSR_117 INVX1_23/gnd DFFSR_91/S FILL
XFILL_17_6 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_34_1 INVX1_8/gnd DFFSR_7/S FILL
XFILL_7_OAI21X1_171 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_46_DFFSR_39 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_35_DFFSR_79 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_32_DFFSR_151 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_22_DFFSR_154 BUFX2_36/A DFFSR_6/S FILL
XFILL_2_DFFSR_36 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_19_DFFSR_29 INVX1_4/gnd DFFSR_4/S FILL
XFILL_12_DFFSR_157 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_8_OAI21X1_105 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_2_INVX1_308 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_20_CLKBUF1_19 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_8_DFFSR_151 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_19_CLKBUF1_22 INVX1_94/gnd DFFSR_25/S FILL
XFILL_19_DFFSR_2 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_43_DFFSR_86 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_18_CLKBUF1_25 INVX1_23/gnd DFFSR_186/S FILL
XFILL_49_DFFSR_182 INVX1_89/gnd DFFSR_36/S FILL
XFILL_39_DFFSR_185 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_1_INVX1_128 INVX1_23/gnd DFFSR_91/S FILL
XFILL_16_DFFSR_76 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_27_DFFSR_36 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_11_DFFPOSX1_21 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_7_NAND3X1_117 INVX1_94/gnd DFFSR_25/S FILL
XFILL_3_BUFX2_3 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_29_DFFSR_188 INVX1_2/gnd DFFSR_1/S FILL
XFILL_19_DFFSR_191 INVX1_23/gnd DFFSR_91/S FILL
XFILL_6_OAI21X1_201 BUFX2_35/A DFFSR_97/S FILL
XFILL_51_DFFSR_93 INVX1_2/gnd DFFSR_51/S FILL
XOAI21X1_237 AOI21X1_36/Y AOI21X1_29/Y NAND3X1_85/Y BUFX2_8/gnd AOI21X1_37/A DFFSR_10/S
+ OAI21X1
XFILL_7_OAI21X1_135 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_24_DFFSR_83 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_35_DFFSR_43 INVX1_94/gnd DFFSR_25/S FILL
XFILL_21_DFFPOSX1_10 INVX1_8/gnd DFFSR_5/S FILL
XFILL_7_DFFSR_90 INVX1_2/gnd DFFSR_1/S FILL
XFILL_42_DFFSR_112 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_32_DFFSR_115 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_5_DFFSR_188 INVX1_2/gnd DFFSR_1/S FILL
XFILL_22_DFFSR_118 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_6_BUFX2_28 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_12_DFFSR_121 BUFX2_36/A DFFSR_6/S FILL
XFILL_26_5_0 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_5_NAND2X1_9 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_2_INVX1_272 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_4_INVX1_84 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_43_DFFSR_50 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_49_DFFSR_146 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_8_DFFSR_115 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_5_OAI21X1_231 BUFX2_36/A DFFSR_6/S FILL
XFILL_5_OAI22X1_8 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_32_DFFSR_90 INVX1_2/gnd DFFSR_1/S FILL
XFILL_39_DFFSR_149 INVX1_23/gnd DFFSR_91/S FILL
XFILL_16_DFFSR_40 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_29_DFFSR_152 BUFX2_5/gnd DFFSR_23/S FILL
XNAND3X1_2 NAND3X1_2/A NAND3X1_2/B OR2X2_1/Y BUFX2_8/gnd NAND3X1_2/Y DFFSR_10/S NAND3X1
XFILL_39_6 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_6_OAI21X1_165 BUFX2_35/A DFFSR_97/S FILL
XFILL_19_DFFSR_155 BUFX2_7/gnd DFFSR_54/S FILL
XNOR2X1_37 NOR2X1_37/A NOR2X1_37/B INVX1_94/gnd NOR2X1_37/Y DFFSR_25/S NOR2X1
XFILL_40_DFFSR_97 BUFX2_35/A DFFSR_97/S FILL
XFILL_4_NOR2X1_34 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_51_DFFSR_57 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_3_INVX1_416 DFFSR_89/gnd DFFSR_92/S FILL
XOAI21X1_201 INVX1_226/Y INVX1_240/Y OAI21X1_201/C BUFX2_35/A NAND3X1_35/A DFFSR_97/S
+ OAI21X1
XFILL_1_AND2X2_6 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_6_NAND2X1_279 INVX1_89/gnd DFFSR_2/S FILL
XFILL_5_DFFSR_152 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_7_DFFSR_54 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_24_DFFSR_47 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_11_CLKBUF1_10 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_13_DFFSR_87 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_46_DFFSR_183 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_10_CLKBUF1_13 INVX1_4/gnd DFFSR_51/S FILL
XFILL_36_0_0 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_36_DFFSR_186 INVX1_23/gnd DFFSR_186/S FILL
XFILL_9_CLKBUF1_16 BUFX2_36/A DFFSR_6/S FILL
XFILL_4_OAI21X1_261 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_34_2_1 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_26_DFFSR_189 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_2_INVX1_236 INVX1_8/gnd DFFSR_7/S FILL
XFILL_7_DFFSR_1 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_10_DFFSR_9 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_8_CLKBUF1_19 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_7_CLKBUF1_22 INVX1_94/gnd DFFSR_25/S FILL
XFILL_6_NAND3X1_111 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_32_4_2 INVX1_8/gnd DFFSR_5/S FILL
XFILL_6_CLKBUF1_25 INVX1_23/gnd DFFSR_186/S FILL
XFILL_10_DFFPOSX1_15 BUFX2_35/A DFFSR_14/S FILL
XFILL_43_DFFSR_14 BUFX2_35/A DFFSR_14/S FILL
XFILL_5_OAI21X1_195 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_32_DFFSR_54 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_21_DFFSR_94 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_4_INVX1_48 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_49_DFFSR_110 DFFSR_73/gnd DFFSR_57/S FILL
XCLKBUF1_25 INVX1_402/Y INVX1_23/gnd INVX1_1/A DFFSR_186/S CLKBUF1
XFILL_39_DFFSR_113 INVX1_23/gnd DFFSR_186/S FILL
XFILL_3_BUFX2_39 BUFX2_43/A DFFSR_97/S FILL
XFILL_5_OR2X2_1 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_29_DFFSR_116 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_2_DFFSR_189 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_19_DFFSR_119 BUFX2_37/A DFFSR_81/S FILL
XFILL_6_OAI21X1_129 INVX1_4/gnd DFFSR_4/S FILL
XFILL_31_DFFSR_5 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_40_DFFSR_61 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_1_INVX1_95 BUFX2_5/gnd DFFSR_6/S FILL
XOAI21X1_165 BUFX2_2/Y INVX1_199/Y OAI21X1_165/C BUFX2_35/A DFFSR_165/D DFFSR_97/S
+ OAI21X1
XFILL_0_DFFPOSX1_26 BUFX2_37/A DFFSR_81/S FILL
XFILL_3_INVX1_380 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_7_DFFSR_18 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_24_DFFSR_11 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_6_NAND2X1_243 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_46_DFFSR_147 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_5_DFFSR_116 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_2_OAI22X1_9 INVX1_8/gnd DFFSR_5/S FILL
XFILL_13_DFFSR_51 INVX1_2/gnd DFFSR_51/S FILL
XFILL_4_OAI21X1_225 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_36_DFFSR_150 BUFX2_8/gnd DFFSR_25/S FILL
XNAND2X1_279 NOR3X1_2/Y XOR2X1_14/A INVX1_89/gnd AOI22X1_14/C DFFSR_2/S NAND2X1
XFILL_48_DFFSR_68 BUFX2_35/A DFFSR_14/S FILL
XFILL_26_DFFSR_153 BUFX2_36/A DFFSR_8/S FILL
XFILL_2_INVX1_200 INVX1_4/gnd DFFSR_4/S FILL
XFILL_16_DFFSR_156 INVX1_23/gnd DFFSR_91/S FILL
XFILL_4_DFFSR_65 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_5_OAI21X1_159 BUFX2_43/A DFFSR_97/S FILL
XFILL_1_NOR2X1_35 INVX1_94/gnd DFFSR_52/S FILL
XFILL_10_DFFSR_98 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_32_DFFSR_18 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_21_DFFSR_58 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_0_INVX1_417 INVX1_23/gnd DFFSR_91/S FILL
XNAND3X1_111 NOR2X1_1/B INVX1_264/Y INVX1_265/Y DFFSR_71/gnd OAI22X1_9/B DFFSR_45/S
+ NAND3X1
XFILL_2_DFFSR_153 BUFX2_36/A DFFSR_8/S FILL
XFILL_43_DFFSR_184 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_5_NAND2X1_273 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_33_DFFSR_187 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_23_DFFSR_190 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_1_INVX1_59 INVX1_94/gnd DFFSR_25/S FILL
XFILL_40_DFFSR_25 BUFX2_8/gnd DFFSR_25/S FILL
XOAI21X1_129 DFFSR_51/S INVX1_146/Y OAI21X1_129/C INVX1_4/gnd DFFSR_129/D DFFSR_4/S
+ OAI21X1
XFILL_29_DFFSR_65 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_6_NAND2X1_207 BUFX2_43/A DFFSR_97/S FILL
XFILL_3_INVX1_344 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_3_OAI21X1_255 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_13_DFFSR_15 INVX1_8/gnd DFFSR_7/S FILL
XFILL_5_NAND3X1_105 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_46_DFFSR_111 INVX1_8/gnd DFFSR_5/S FILL
XFILL_36_DFFSR_114 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_9_DFFSR_187 BUFX2_16/gnd DFFSR_11/S FILL
XNAND2X1_243 NOR2X1_31/Y NOR2X1_30/Y DFFSR_73/gnd NAND2X1_243/Y DFFSR_57/S NAND2X1
XFILL_26_DFFSR_117 INVX1_23/gnd DFFSR_91/S FILL
XFILL_4_OAI21X1_189 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_2_INVX1_164 INVX1_23/gnd DFFSR_91/S FILL
XFILL_37_DFFSR_72 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_48_DFFSR_32 INVX1_2/gnd DFFSR_1/S FILL
XFILL_16_DFFSR_120 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_5_OAI21X1_123 INVX1_23/gnd DFFSR_91/S FILL
XFILL_10_DFFSR_62 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_21_DFFSR_22 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_4_DFFSR_29 INVX1_4/gnd DFFSR_4/S FILL
XFILL_21_3 INVX1_94/gnd DFFSR_52/S FILL
XFILL_0_INVX1_381 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_9_OAI22X1_7 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_43_DFFSR_148 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_2_DFFSR_117 INVX1_23/gnd DFFSR_91/S FILL
XFILL_33_5_0 INVX1_8/gnd DFFSR_7/S FILL
XFILL_5_NAND2X1_237 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_45_DFFSR_79 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_33_DFFSR_151 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_1_INVX1_23 INVX1_23/gnd DFFSR_91/S FILL
XFILL_18_DFFSR_69 BUFX2_43/A DFFSR_23/S FILL
XFILL_23_DFFSR_154 BUFX2_36/A DFFSR_6/S FILL
XFILL_1_DFFSR_76 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_29_DFFSR_29 INVX1_4/gnd DFFSR_4/S FILL
XFILL_13_DFFSR_157 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_3_OAI21X1_219 BUFX2_35/A DFFSR_97/S FILL
XFILL_3_INVX1_308 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_6_NAND2X1_171 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_5_XOR2X1_6 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_22_DFFPOSX1_1 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_0_BUFX2_14 BUFX2_37/A DFFSR_81/S FILL
XNAND2X1_207 AOI22X1_8/A AOI22X1_8/B BUFX2_43/A AOI21X1_25/A DFFSR_97/S NAND2X1
XFILL_43_DFFSR_8 BUFX2_36/A DFFSR_8/S FILL
XFILL_9_DFFSR_151 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_21_DFFPOSX1_4 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_4_OAI21X1_153 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_20_DFFPOSX1_7 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_50_DFFSR_182 INVX1_89/gnd DFFSR_36/S FILL
XFILL_18_DFFPOSX1_28 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_40_DFFSR_185 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_2_INVX1_128 INVX1_23/gnd DFFSR_91/S FILL
XFILL_26_DFFSR_76 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_9_DFFSR_83 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_37_DFFSR_36 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_30_DFFSR_188 INVX1_2/gnd DFFSR_1/S FILL
XFILL_20_DFFSR_191 INVX1_23/gnd DFFSR_91/S FILL
XFILL_10_DFFSR_26 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_4_NAND2X1_267 INVX1_4/gnd DFFSR_4/S FILL
XFILL_0_INVX1_345 INVX1_94/gnd DFFSR_52/S FILL
XFILL_43_0_0 INVX1_4/gnd DFFSR_51/S FILL
XFILL_4_7 INVX1_23/gnd DFFSR_91/S FILL
XFILL_2_OAI21X1_249 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_5_NAND2X1_201 BUFX2_35/A DFFSR_14/S FILL
XFILL_34_DFFSR_83 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_45_DFFSR_43 INVX1_94/gnd DFFSR_25/S FILL
XFILL_41_2_1 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_43_DFFSR_112 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_33_DFFSR_115 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_6_DFFSR_188 INVX1_2/gnd DFFSR_1/S FILL
XFILL_23_DFFSR_118 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_13_DFFSR_121 BUFX2_36/A DFFSR_6/S FILL
XFILL_18_DFFSR_33 INVX1_94/gnd DFFSR_52/S FILL
XFILL_1_DFFSR_40 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_6_NAND2X1_9 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_39_4_2 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_6_NAND2X1_135 BUFX2_36/A DFFSR_6/S FILL
XFILL_3_OAI21X1_183 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_3_INVX1_272 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_11_XOR2X1_3 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_50_DFFSR_146 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_9_DFFSR_115 BUFX2_6/gnd DFFSR_14/S FILL
XNAND2X1_171 DFFSR_25/S DFFPOSX1_20/Q BUFX2_19/gnd NAND2X1_171/Y DFFSR_54/S NAND2X1
XFILL_6_OAI22X1_8 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_42_DFFSR_90 INVX1_2/gnd DFFSR_1/S FILL
XFILL_4_OAI21X1_117 BUFX2_35/A DFFSR_97/S FILL
XFILL_40_DFFSR_149 INVX1_23/gnd DFFSR_91/S FILL
XFILL_9_DFFSR_47 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_26_DFFSR_40 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_43_3 INVX1_4/gnd DFFSR_4/S FILL
XFILL_15_DFFSR_80 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_30_DFFSR_152 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_4_NAND2X1_231 BUFX2_37/A DFFSR_81/S FILL
XFILL_20_DFFSR_155 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_10_DFFSR_158 BUFX2_43/A DFFSR_23/S FILL
XFILL_3_NAND3X1_129 BUFX2_35/A DFFSR_14/S FILL
XFILL_50_DFFSR_97 BUFX2_35/A DFFSR_97/S FILL
XFILL_5_NOR2X1_34 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_0_INVX1_309 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_30_DFFSR_2 DFFSR_5/gnd DFFSR_2/S FILL
XINVX1_419 BUFX2_30/A INVX1_2/gnd INVX1_419/Y DFFSR_51/S INVX1
XFILL_4_INVX1_416 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_2_OAI21X1_213 BUFX2_36/A DFFSR_6/S FILL
XFILL_6_DFFSR_152 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_5_NAND2X1_165 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_34_DFFSR_47 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_23_DFFSR_87 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_6_DFFSR_94 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_47_DFFSR_183 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_37_DFFSR_186 INVX1_23/gnd DFFSR_186/S FILL
XFILL_3_OAI21X1_147 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_10_DFFPOSX1_1 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_27_DFFSR_189 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_5_BUFX2_32 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_17_DFFPOSX1_22 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_3_INVX1_236 INVX1_8/gnd DFFSR_7/S FILL
XFILL_9_DFFPOSX1_4 BUFX2_17/gnd DFFSR_7/S FILL
XNAND2X1_135 DFFSR_8/S NAND2X1_71/B BUFX2_36/A OAI21X1_135/C DFFSR_6/S NAND2X1
XFILL_42_DFFSR_54 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_8_DFFPOSX1_7 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_3_INVX1_88 INVX1_2/gnd DFFSR_1/S FILL
XFILL_31_DFFSR_94 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_8_AOI21X1_27 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_3_NAND2X1_261 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_27_DFFPOSX1_11 INVX1_4/gnd DFFSR_4/S FILL
XFILL_50_DFFSR_110 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_40_DFFSR_113 INVX1_23/gnd DFFSR_186/S FILL
XFILL_7_AOI21X1_30 INVX1_23/gnd DFFSR_91/S FILL
XFILL_15_DFFSR_44 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_9_DFFSR_11 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_6_AOI21X1_33 BUFX2_35/A DFFSR_14/S FILL
XFILL_15_0_1 BUFX2_37/A DFFSR_81/S FILL
XFILL_30_DFFSR_116 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_3_DFFSR_189 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_1_OAI21X1_243 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_20_DFFSR_119 BUFX2_37/A DFFSR_81/S FILL
XFILL_5_AOI21X1_36 BUFX2_8/gnd DFFSR_25/S FILL
XAOI21X1_33 AOI21X1_33/A AOI21X1_33/B INVX1_253/A BUFX2_35/A AOI21X1_33/Y DFFSR_14/S
+ AOI21X1
XFILL_13_2_2 BUFX2_36/A DFFSR_8/S FILL
XFILL_4_NAND2X1_195 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_10_DFFSR_122 INVX1_94/gnd DFFSR_52/S FILL
XFILL_50_DFFSR_61 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_4_AOI21X1_39 BUFX2_7/gnd DFFSR_81/S FILL
XINVX1_383 DFFSR_87/Q INVX1_89/gnd INVX1_383/Y DFFSR_2/S INVX1
XFILL_0_AOI21X1_1 INVX1_8/gnd DFFSR_5/S FILL
XFILL_0_INVX1_273 INVX1_8/gnd DFFSR_5/S FILL
XFILL_3_AOI21X1_42 INVX1_23/gnd DFFSR_91/S FILL
XFILL_2_OAI21X1_177 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_4_INVX1_380 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_2_AOI21X1_45 INVX1_89/gnd DFFSR_36/S FILL
XFILL_5_NAND2X1_129 INVX1_4/gnd DFFSR_4/S FILL
XFILL_6_DFFSR_58 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_34_DFFSR_11 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_12_DFFSR_91 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_1_AOI21X1_48 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_6_DFFSR_116 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_3_OAI22X1_9 INVX1_8/gnd DFFSR_5/S FILL
XFILL_23_DFFSR_51 INVX1_2/gnd DFFSR_51/S FILL
XFILL_47_DFFSR_147 DFFSR_89/gnd DFFSR_186/S FILL
XBUFX2_36 BUFX2_36/A BUFX2_5/gnd BUFX2_36/Y DFFSR_23/S BUFX2
XFILL_37_DFFSR_150 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_27_DFFSR_153 BUFX2_36/A DFFSR_8/S FILL
XFILL_3_OAI21X1_111 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_3_INVX1_200 INVX1_4/gnd DFFSR_4/S FILL
XFILL_17_DFFSR_156 INVX1_23/gnd DFFSR_91/S FILL
XFILL_48_8 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_8_OAI21X1_75 INVX1_4/gnd DFFSR_4/S FILL
XFILL_7_OAI21X1_78 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_6_NAND2X1_96 INVX1_4/gnd DFFSR_51/S FILL
XFILL_40_5_0 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_5_NAND2X1_99 BUFX2_43/A DFFSR_97/S FILL
XFILL_3_NAND2X1_225 BUFX2_36/A DFFSR_8/S FILL
XFILL_3_INVX1_52 BUFX2_37/A DFFSR_81/S FILL
XFILL_6_OAI21X1_81 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_2_NOR2X1_35 INVX1_94/gnd DFFSR_52/S FILL
XFILL_20_DFFSR_98 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_42_DFFSR_18 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_31_DFFSR_58 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_1_INVX1_417 INVX1_23/gnd DFFSR_91/S FILL
XFILL_5_OAI21X1_84 BUFX2_5/gnd DFFSR_6/S FILL
XNAND2X1_96 BUFX2_15/Y DFFSR_88/Q INVX1_4/gnd OAI21X1_96/C DFFSR_51/S NAND2X1
XFILL_2_BUFX2_43 BUFX2_35/A DFFSR_97/S FILL
XFILL_3_DFFSR_153 BUFX2_36/A DFFSR_8/S FILL
XOAI21X1_81 BUFX2_19/Y INVX1_92/Y OAI21X1_81/C BUFX2_19/gnd DFFSR_81/D DFFSR_54/S
+ OAI21X1
XFILL_2_NAND3X1_123 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_4_OAI21X1_87 INVX1_4/gnd DFFSR_4/S FILL
XFILL_3_OAI21X1_90 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_44_DFFSR_184 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_4_NAND2X1_159 BUFX2_43/A DFFSR_97/S FILL
XFILL_1_OAI21X1_207 BUFX2_37/A DFFSR_8/S FILL
XFILL_2_OAI21X1_93 INVX1_4/gnd DFFSR_51/S FILL
XFILL_34_DFFSR_187 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_24_DFFSR_190 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_21_DFFSR_9 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_50_DFFSR_25 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_0_INVX1_237 INVX1_8/gnd DFFSR_7/S FILL
XFILL_1_OAI21X1_96 INVX1_4/gnd DFFSR_51/S FILL
XFILL_0_INVX1_99 INVX1_4/gnd DFFSR_4/S FILL
XINVX1_347 DFFSR_90/Q INVX1_4/gnd INVX1_347/Y DFFSR_4/S INVX1
XFILL_39_DFFSR_65 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_16_DFFPOSX1_16 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_0_OAI21X1_99 BUFX2_43/A DFFSR_97/S FILL
XFILL_2_OAI21X1_141 INVX1_94/gnd DFFSR_52/S FILL
XFILL_4_INVX1_344 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_6_DFFSR_22 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_12_DFFSR_55 INVX1_89/gnd DFFSR_36/S FILL
XFILL_1_AOI21X1_12 INVX1_8/gnd DFFSR_7/S FILL
XFILL_23_DFFSR_15 INVX1_8/gnd DFFSR_7/S FILL
XFILL_0_AOI21X1_15 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_47_DFFSR_111 INVX1_8/gnd DFFSR_5/S FILL
XFILL_37_DFFSR_114 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_27_DFFSR_117 INVX1_23/gnd DFFSR_91/S FILL
XFILL_5_NOR2X1_3 INVX1_94/gnd DFFSR_25/S FILL
XFILL_9_OAI21X1_36 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_42_DFFSR_5 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_0_DFFSR_190 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_2_NAND2X1_255 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_3_INVX1_164 INVX1_23/gnd DFFSR_91/S FILL
XFILL_47_DFFSR_72 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_17_DFFSR_120 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_8_OAI21X1_39 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_3_INVX1_16 BUFX2_43/A DFFSR_23/S FILL
XFILL_3_DFFSR_69 BUFX2_43/A DFFSR_23/S FILL
XFILL_6_NAND2X1_60 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_20_DFFSR_62 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_0_OAI21X1_237 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_31_DFFSR_22 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_6_DFFPOSX1_27 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_7_OAI21X1_42 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_3_NAND2X1_189 BUFX2_5/gnd DFFSR_6/S FILL
XNAND2X1_60 DFFSR_54/S DFFSR_52/Q BUFX2_7/gnd OAI21X1_60/C DFFSR_54/S NAND2X1
XFILL_5_NAND2X1_63 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_6_OAI21X1_45 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_48_2_1 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_1_INVX1_381 DFFSR_79/gnd DFFSR_45/S FILL
XOAI21X1_45 DFFSR_36/S INVX1_51/Y OAI21X1_45/C DFFSR_79/gnd DFFSR_45/D DFFSR_36/S
+ OAI21X1
XFILL_4_NAND2X1_66 INVX1_4/gnd DFFSR_51/S FILL
XFILL_5_OAI21X1_48 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_3_DFFSR_117 INVX1_23/gnd DFFSR_91/S FILL
XFILL_3_NAND2X1_69 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_46_4_2 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_4_OAI21X1_51 INVX1_2/gnd DFFSR_51/S FILL
XFILL_44_DFFSR_148 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_3_OAI21X1_54 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_1_OAI21X1_171 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_2_NAND2X1_72 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_4_NAND2X1_123 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_34_DFFSR_151 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_1_NAND2X1_75 INVX1_4/gnd DFFSR_4/S FILL
XFILL_2_OAI21X1_57 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_28_DFFSR_69 BUFX2_43/A DFFSR_23/S FILL
XFILL_24_DFFSR_154 BUFX2_36/A DFFSR_6/S FILL
XFILL_1_OAI21X1_60 BUFX2_37/A DFFSR_81/S FILL
XINVX1_311 INVX1_70/A INVX1_94/gnd INVX1_311/Y DFFSR_52/S INVX1
XFILL_0_INVX1_201 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_0_INVX1_63 INVX1_2/gnd DFFSR_51/S FILL
XFILL_39_DFFSR_29 INVX1_4/gnd DFFSR_4/S FILL
XFILL_0_NAND2X1_78 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_14_DFFSR_157 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_0_OAI21X1_63 INVX1_94/gnd DFFSR_25/S FILL
XFILL_2_OAI21X1_105 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_4_INVX1_308 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_1_NAND2X1_285 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_14_3_0 BUFX2_37/A DFFSR_8/S FILL
XFILL_12_DFFSR_19 DFFSR_1/gnd DFFSR_9/S FILL
XNOR2X1_7 NOR2X1_7/A NOR2X1_7/B DFFSR_89/gnd NOR2X1_7/Y DFFSR_92/S NOR2X1
XFILL_0_DFFSR_154 BUFX2_36/A DFFSR_6/S FILL
XFILL_2_NAND2X1_219 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_51_DFFSR_182 INVX1_89/gnd DFFSR_36/S FILL
XFILL_41_DFFSR_185 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_3_INVX1_128 INVX1_23/gnd DFFSR_91/S FILL
XFILL_12_5_1 BUFX2_36/A DFFSR_6/S FILL
XFILL_36_DFFSR_76 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_47_DFFSR_36 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_1_NAND3X1_117 INVX1_94/gnd DFFSR_25/S FILL
XFILL_31_DFFSR_188 INVX1_2/gnd DFFSR_1/S FILL
XFILL_21_DFFSR_191 INVX1_23/gnd DFFSR_91/S FILL
XFILL_6_NAND2X1_24 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_0_OAI21X1_201 BUFX2_35/A DFFSR_97/S FILL
XFILL_3_NAND2X1_153 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_3_DFFSR_33 INVX1_94/gnd DFFSR_52/S FILL
XFILL_5_NAND2X1_27 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_20_DFFSR_26 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_5_OAI21X1_12 BUFX2_35/A DFFSR_14/S FILL
XFILL_1_INVX1_345 INVX1_94/gnd DFFSR_52/S FILL
XFILL_4_NAND2X1_30 DFFSR_79/gnd DFFSR_36/S FILL
XNAND2X1_24 DFFSR_57/S DFFSR_16/Q DFFSR_73/gnd NAND2X1_24/Y DFFSR_57/S NAND2X1
XFILL_9_DFFSR_8 BUFX2_36/A DFFSR_8/S FILL
XFILL_3_NAND2X1_33 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_4_OAI21X1_15 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_2_NAND2X1_36 DFFSR_71/gnd DFFSR_45/S FILL
XDFFPOSX1_27 AOI22X1_9/B CLKBUF1_15/Y NOR2X1_52/Y DFFSR_71/gnd DFFSR_45/S DFFPOSX1
XFILL_15_DFFPOSX1_10 INVX1_8/gnd DFFSR_5/S FILL
XFILL_3_OAI21X1_18 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_44_DFFSR_112 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_34_DFFSR_115 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_1_OAI21X1_135 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_44_DFFSR_83 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_1_NAND2X1_39 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_7_DFFSR_188 INVX1_2/gnd DFFSR_1/S FILL
XFILL_2_OAI21X1_21 INVX1_2/gnd DFFSR_51/S FILL
XFILL_8_NAND3X1_95 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_0_NAND2X1_42 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_24_DFFSR_118 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_0_INVX1_165 INVX1_23/gnd DFFSR_186/S FILL
XFILL_7_NAND3X1_98 BUFX2_35/A DFFSR_14/S FILL
XFILL_14_DFFSR_121 BUFX2_36/A DFFSR_6/S FILL
XFILL_28_DFFSR_33 INVX1_94/gnd DFFSR_52/S FILL
XAOI21X1_3 AOI22X1_4/B AOI21X1_3/B INVX1_223/Y DFFSR_79/gnd AOI21X1_3/Y DFFSR_45/S
+ AOI21X1
XFILL_0_DFFSR_80 BUFX2_16/gnd DFFSR_65/S FILL
XINVX1_275 INVX1_48/A BUFX2_16/gnd INVX1_275/Y DFFSR_11/S INVX1
XFILL_17_DFFSR_73 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_1_OAI21X1_24 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_0_INVX1_27 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_1_NAND2X1_249 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_0_OAI21X1_27 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_22_0_1 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_7_OAI22X1_8 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_5_DFFPOSX1_21 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_2_NAND2X1_183 INVX1_8/gnd DFFSR_7/S FILL
XFILL_0_DFFSR_118 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_41_DFFSR_149 INVX1_23/gnd DFFSR_91/S FILL
XFILL_20_2_2 INVX1_94/gnd DFFSR_52/S FILL
XFILL_36_DFFSR_40 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_8_DFFSR_87 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_25_DFFSR_80 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_2_1_1 INVX1_23/gnd DFFSR_186/S FILL
XFILL_31_DFFSR_152 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_3_AOI22X1_11 INVX1_23/gnd DFFSR_91/S FILL
XFILL_0_OAI21X1_165 BUFX2_35/A DFFSR_97/S FILL
XFILL_21_DFFSR_155 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_0_3_2 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_3_NAND2X1_117 BUFX2_35/A DFFSR_14/S FILL
XFILL_11_DFFSR_158 BUFX2_43/A DFFSR_23/S FILL
XFILL_2_AOI22X1_14 DFFSR_79/gnd DFFSR_36/S FILL
XINVX1_1 INVX1_1/A BUFX2_37/A INVX1_1/Y DFFSR_81/S INVX1
XFILL_6_NOR2X1_34 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_1_INVX1_309 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_7_DFFSR_152 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_10_OAI22X1_38 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_0_NAND2X1_279 INVX1_89/gnd DFFSR_2/S FILL
XFILL_44_DFFSR_47 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_24_DFFPOSX1_29 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_33_DFFSR_87 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_48_DFFSR_183 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_38_DFFSR_186 INVX1_23/gnd DFFSR_186/S FILL
XINVX1_239 INVX1_239/A BUFX2_35/A INVX1_239/Y DFFSR_97/S INVX1
XFILL_8_NAND3X1_59 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_0_DFFSR_44 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_0_INVX1_129 INVX1_89/gnd DFFSR_36/S FILL
XFILL_17_DFFSR_37 INVX1_89/gnd DFFSR_2/S FILL
XFILL_9_OAI22X1_41 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_7_NAND3X1_62 BUFX2_43/A DFFSR_23/S FILL
XFILL_28_DFFSR_189 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_47_5_0 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_8_OAI22X1_44 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_6_NAND3X1_65 BUFX2_35/A DFFSR_14/S FILL
XFILL_1_NAND2X1_213 BUFX2_35/A DFFSR_97/S FILL
XFILL_7_OAI22X1_47 BUFX2_37/A DFFSR_8/S FILL
XFILL_5_NAND3X1_68 BUFX2_35/A DFFSR_14/S FILL
XFILL_0_NAND3X1_111 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_6_OAI22X1_50 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_10_XOR2X1_7 INVX1_23/gnd DFFSR_91/S FILL
XFILL_4_NAND3X1_71 BUFX2_35/A DFFSR_14/S FILL
XNAND3X1_65 NAND3X1_64/Y NAND3X1_68/B NAND3X1_69/C BUFX2_35/A AOI22X1_10/C DFFSR_14/S
+ NAND3X1
XFILL_5_OAI22X1_53 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_41_DFFSR_94 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_2_NAND2X1_147 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_3_NAND3X1_74 BUFX2_35/A DFFSR_14/S FILL
XFILL_4_OAI22X1_56 BUFX2_37/A DFFSR_8/S FILL
XOAI22X1_50 INVX1_358/Y OAI22X1_38/B INVX1_359/Y OAI22X1_40/D DFFSR_79/gnd NOR2X1_34/A
+ DFFSR_36/S OAI22X1
XFILL_41_DFFSR_113 INVX1_23/gnd DFFSR_186/S FILL
XFILL_2_NAND3X1_77 BUFX2_37/A DFFSR_81/S FILL
XFILL_25_DFFSR_44 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_8_OAI21X1_250 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_3_OAI22X1_59 INVX1_8/gnd DFFSR_7/S FILL
XFILL_2_AND2X2_3 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_8_DFFSR_51 INVX1_2/gnd DFFSR_51/S FILL
XFILL_14_DFFSR_84 BUFX2_43/A DFFSR_23/S FILL
XFILL_1_NAND3X1_80 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_2_OAI22X1_62 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_31_DFFSR_116 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_4_DFFSR_189 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_0_NAND3X1_83 BUFX2_37/A DFFSR_81/S FILL
XFILL_21_DFFSR_119 BUFX2_37/A DFFSR_81/S FILL
XFILL_1_OAI22X1_65 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_11_DFFSR_122 INVX1_94/gnd DFFSR_52/S FILL
XFILL_0_OAI22X1_68 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_0_OAI21X1_129 INVX1_4/gnd DFFSR_4/S FILL
XFILL_1_AOI21X1_1 INVX1_8/gnd DFFSR_5/S FILL
XFILL_1_INVX1_273 INVX1_8/gnd DFFSR_5/S FILL
XFILL_20_DFFSR_6 BUFX2_5/gnd DFFSR_6/S FILL
XINVX1_85 INVX1_85/A DFFSR_3/gnd INVX1_85/Y DFFSR_65/S INVX1
XFILL_0_NAND2X1_243 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_22_DFFSR_91 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_7_DFFSR_116 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_4_OAI22X1_9 INVX1_8/gnd DFFSR_5/S FILL
XFILL_5_DFFSR_98 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_33_DFFSR_51 INVX1_2/gnd DFFSR_51/S FILL
XFILL_44_DFFSR_11 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_48_DFFSR_147 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_8_NAND3X1_23 BUFX2_37/A DFFSR_81/S FILL
XFILL_4_BUFX2_7 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_4_BUFX2_36 BUFX2_5/gnd DFFSR_23/S FILL
XINVX1_203 BUFX2_11/Y BUFX2_36/A INVX1_203/Y DFFSR_6/S INVX1
XFILL_7_NAND3X1_26 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_38_DFFSR_150 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_4_DFFPOSX1_15 BUFX2_35/A DFFSR_14/S FILL
XFILL_28_DFFSR_153 BUFX2_36/A DFFSR_8/S FILL
XFILL_6_NAND3X1_29 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_1_NAND2X1_177 INVX1_89/gnd DFFSR_36/S FILL
XFILL_4_INVX1_200 INVX1_4/gnd DFFSR_4/S FILL
XFILL_7_OAI22X1_11 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_18_DFFSR_156 INVX1_23/gnd DFFSR_91/S FILL
XFILL_5_NAND3X1_32 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_6_OAI22X1_14 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_4_NAND3X1_35 BUFX2_35/A DFFSR_97/S FILL
XNAND3X1_29 AOI21X1_7/A AOI21X1_7/B AOI21X1_7/C BUFX2_7/gnd NAND3X1_56/A DFFSR_54/S
+ NAND3X1
XFILL_41_DFFSR_2 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_2_INVX1_92 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_3_NOR2X1_35 INVX1_94/gnd DFFSR_52/S FILL
XFILL_5_OAI22X1_17 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_30_DFFSR_98 DFFSR_9/gnd DFFSR_9/S FILL
XOAI22X1_14 INVX1_283/Y OAI22X1_6/B INVX1_284/Y OAI22X1_6/D DFFSR_3/gnd NOR2X1_16/A
+ DFFSR_4/S OAI22X1
XFILL_41_DFFSR_58 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_2_INVX1_417 INVX1_23/gnd DFFSR_91/S FILL
XDFFSR_156 DFFSR_156/Q CLKBUF1_12/Y INVX1_187/Y DFFSR_91/S DFFSR_156/D INVX1_23/gnd
+ DFFSR_91/S DFFSR
XFILL_8_OAI21X1_214 BUFX2_35/A DFFSR_97/S FILL
XFILL_3_NAND3X1_38 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_4_OAI22X1_20 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_2_NAND2X1_111 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_2_NAND3X1_41 BUFX2_43/A DFFSR_23/S FILL
XFILL_4_DFFSR_153 BUFX2_36/A DFFSR_8/S FILL
XFILL_3_OAI22X1_23 INVX1_89/gnd DFFSR_2/S FILL
XFILL_8_DFFSR_15 INVX1_8/gnd DFFSR_7/S FILL
XFILL_14_DFFSR_48 INVX1_4/gnd DFFSR_4/S FILL
XFILL_1_NAND3X1_44 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_2_OAI22X1_26 INVX1_94/gnd DFFSR_52/S FILL
XFILL_45_DFFSR_184 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_0_NAND3X1_47 BUFX2_43/A DFFSR_97/S FILL
XFILL_1_OAI22X1_29 INVX1_8/gnd DFFSR_5/S FILL
XFILL_35_DFFSR_187 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_23_DFFPOSX1_23 INVX1_23/gnd DFFSR_91/S FILL
XFILL_0_OAI22X1_32 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_25_DFFSR_190 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_21_3_0 INVX1_94/gnd DFFSR_25/S FILL
XFILL_1_INVX1_237 INVX1_8/gnd DFFSR_7/S FILL
XFILL_49_DFFSR_65 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_0_NAND2X1_207 BUFX2_43/A DFFSR_97/S FILL
XFILL_19_5_1 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_5_DFFSR_62 BUFX2_19/gnd DFFSR_52/S FILL
XINVX1_49 DFFSR_43/Q BUFX2_8/gnd INVX1_49/Y DFFSR_10/S INVX1
XFILL_11_DFFSR_95 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_22_DFFSR_55 INVX1_89/gnd DFFSR_36/S FILL
XFILL_33_DFFSR_15 INVX1_8/gnd DFFSR_7/S FILL
XFILL_1_4_0 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_48_DFFSR_111 INVX1_8/gnd DFFSR_5/S FILL
XINVX1_167 BUFX2_6/Y DFFSR_89/gnd DFFSR_146/R DFFSR_92/S INVX1
XFILL_38_DFFSR_114 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_28_DFFSR_117 INVX1_23/gnd DFFSR_91/S FILL
XFILL_1_DFFSR_190 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_4_INVX1_164 INVX1_23/gnd DFFSR_91/S FILL
XFILL_1_NAND2X1_141 INVX1_94/gnd DFFSR_25/S FILL
XFILL_7_OAI21X1_244 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_18_DFFSR_120 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_30_DFFSR_62 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_41_DFFSR_22 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_2_INVX1_56 DFFSR_73/gnd DFFSR_11/S FILL
XDFFSR_120 INVX1_390/A CLKBUF1_4/Y DFFSR_113/R DFFSR_11/S DFFSR_120/D BUFX2_16/gnd
+ DFFSR_11/S DFFSR
XFILL_8_OAI21X1_178 INVX1_94/gnd DFFSR_25/S FILL
XFILL_2_INVX1_381 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_4_DFFSR_117 INVX1_23/gnd DFFSR_91/S FILL
XFILL_14_DFFSR_12 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_45_DFFSR_148 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_0_NAND3X1_11 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_35_DFFSR_151 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_8_DFFSR_5 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_38_DFFSR_69 BUFX2_43/A DFFSR_23/S FILL
XFILL_25_DFFSR_154 BUFX2_36/A DFFSR_6/S FILL
XFILL_1_INVX1_201 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_49_DFFSR_29 INVX1_4/gnd DFFSR_4/S FILL
XFILL_15_DFFSR_157 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_29_0_1 INVX1_89/gnd DFFSR_2/S FILL
XFILL_0_NAND2X1_171 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_0_NAND3X1_1 INVX1_94/gnd DFFSR_25/S FILL
XDFFSR_66 INVX1_75/A CLKBUF1_5/Y DFFSR_68/R DFFSR_66/S DFFSR_66/D INVX1_2/gnd DFFSR_51/S
+ DFFSR
XINVX1_13 DFFSR_11/Q BUFX2_16/gnd INVX1_13/Y DFFSR_11/S INVX1
XFILL_0_NOR2X1_36 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_27_2_2 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_22_DFFSR_19 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_5_DFFSR_26 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_11_DFFSR_59 INVX1_4/gnd DFFSR_51/S FILL
XFILL_9_1_1 BUFX2_43/A DFFSR_23/S FILL
XFILL_4_NOR2X1_7 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_1_DFFSR_154 BUFX2_36/A DFFSR_6/S FILL
XINVX1_131 INVX1_131/A INVX1_89/gnd INVX1_131/Y DFFSR_36/S INVX1
XFILL_8_NAND3X1_124 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_12_DFFPOSX1_28 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_42_DFFSR_185 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_4_INVX1_128 INVX1_23/gnd DFFSR_91/S FILL
XFILL_1_NAND2X1_105 BUFX2_35/A DFFSR_14/S FILL
XFILL_7_OAI21X1_208 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_46_DFFSR_76 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_32_DFFSR_9 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_7_3_2 BUFX2_35/A DFFSR_97/S FILL
XFILL_32_DFFSR_188 INVX1_2/gnd DFFSR_1/S FILL
XFILL_22_DFFSR_191 INVX1_23/gnd DFFSR_91/S FILL
XFILL_2_INVX1_20 INVX1_8/gnd DFFSR_5/S FILL
XFILL_30_DFFSR_26 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_19_DFFSR_66 INVX1_2/gnd DFFSR_51/S FILL
XFILL_2_DFFSR_73 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_22_DFFPOSX1_17 BUFX2_37/A DFFSR_8/S FILL
XFILL_8_OAI21X1_142 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_2_INVX1_345 INVX1_94/gnd DFFSR_52/S FILL
XFILL_1_BUFX2_11 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_6_XOR2X1_3 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_45_DFFSR_112 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_35_DFFSR_115 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_8_DFFSR_188 INVX1_2/gnd DFFSR_1/S FILL
XFILL_25_DFFSR_118 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_1_INVX1_165 INVX1_23/gnd DFFSR_186/S FILL
XFILL_15_DFFSR_121 BUFX2_36/A DFFSR_6/S FILL
XFILL_38_DFFSR_33 INVX1_94/gnd DFFSR_52/S FILL
XFILL_27_DFFSR_73 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_11_DFFSR_23 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_0_NAND2X1_135 BUFX2_36/A DFFSR_6/S FILL
XFILL_6_OAI21X1_238 BUFX2_19/gnd DFFSR_52/S FILL
XDFFSR_30 DFFSR_30/Q DFFSR_52/CLK DFFSR_31/R DFFSR_36/S DFFSR_30/D INVX1_89/gnd DFFSR_36/S
+ DFFSR
XFILL_8_OAI22X1_8 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_17_7 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_34_2 INVX1_8/gnd DFFSR_7/S FILL
XFILL_1_DFFSR_118 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_42_DFFSR_149 INVX1_23/gnd DFFSR_91/S FILL
XFILL_7_OAI21X1_172 BUFX2_36/A DFFSR_6/S FILL
XFILL_46_DFFSR_40 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_35_DFFSR_80 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_32_DFFSR_152 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_22_DFFSR_155 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_19_DFFSR_30 INVX1_89/gnd DFFSR_36/S FILL
XFILL_2_DFFSR_37 INVX1_89/gnd DFFSR_2/S FILL
XFILL_12_DFFSR_158 BUFX2_43/A DFFSR_23/S FILL
XFILL_2_INVX1_309 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_8_OAI21X1_106 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_20_CLKBUF1_20 INVX1_4/gnd DFFSR_51/S FILL
XFILL_8_DFFSR_152 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_19_CLKBUF1_23 INVX1_89/gnd DFFSR_2/S FILL
XFILL_43_DFFSR_87 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_19_DFFSR_3 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_49_DFFSR_183 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_39_DFFSR_186 INVX1_23/gnd DFFSR_186/S FILL
XFILL_1_INVX1_129 INVX1_89/gnd DFFSR_36/S FILL
XFILL_27_DFFSR_37 INVX1_89/gnd DFFSR_2/S FILL
XFILL_3_BUFX2_4 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_7_NAND3X1_118 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_16_DFFSR_77 INVX1_89/gnd DFFSR_2/S FILL
XFILL_29_DFFSR_189 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_6_OAI21X1_202 BUFX2_35/A DFFSR_14/S FILL
XFILL_11_DFFPOSX1_22 BUFX2_16/gnd DFFSR_11/S FILL
XOAI21X1_238 AND2X2_13/B AND2X2_13/A NAND3X1_2/A BUFX2_19/gnd OAI22X1_4/C DFFSR_52/S
+ OAI21X1
XFILL_42_DFFSR_113 INVX1_23/gnd DFFSR_186/S FILL
XFILL_7_DFFSR_91 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_7_OAI21X1_136 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_21_DFFPOSX1_11 INVX1_4/gnd DFFSR_4/S FILL
XFILL_24_DFFSR_84 BUFX2_43/A DFFSR_23/S FILL
XFILL_35_DFFSR_44 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_28_3_0 INVX1_89/gnd DFFSR_36/S FILL
XFILL_32_DFFSR_116 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_5_DFFSR_189 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_22_DFFSR_119 BUFX2_37/A DFFSR_81/S FILL
XFILL_12_DFFSR_122 INVX1_94/gnd DFFSR_52/S FILL
XFILL_26_5_1 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_6_BUFX2_29 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_8_4_0 BUFX2_43/A DFFSR_97/S FILL
XFILL_2_AOI21X1_1 INVX1_8/gnd DFFSR_5/S FILL
XFILL_2_INVX1_273 INVX1_8/gnd DFFSR_5/S FILL
XFILL_32_DFFSR_91 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_5_OAI21X1_232 BUFX2_35/A DFFSR_97/S FILL
XFILL_8_DFFSR_116 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_5_OAI22X1_9 INVX1_8/gnd DFFSR_5/S FILL
XFILL_43_DFFSR_51 INVX1_2/gnd DFFSR_51/S FILL
XFILL_4_INVX1_85 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_49_DFFSR_147 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_39_DFFSR_150 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_16_DFFSR_41 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_29_DFFSR_153 BUFX2_36/A DFFSR_8/S FILL
XNAND3X1_3 AND2X2_8/A AND2X2_6/A AND2X2_2/Y BUFX2_19/gnd NAND3X1_3/Y DFFSR_54/S NAND3X1
XFILL_39_7 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_19_DFFSR_156 INVX1_23/gnd DFFSR_91/S FILL
XFILL_6_OAI21X1_166 DFFSR_3/gnd DFFSR_4/S FILL
XNOR2X1_38 NOR2X1_38/A NOR2X1_38/B BUFX2_17/gnd NOR2X1_38/Y DFFSR_7/S NOR2X1
XFILL_4_NOR2X1_35 INVX1_94/gnd DFFSR_52/S FILL
XFILL_40_DFFSR_98 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_3_INVX1_417 INVX1_23/gnd DFFSR_91/S FILL
XOAI21X1_202 NOR2X1_7/A INVX1_231/Y AND2X2_9/Y BUFX2_35/A NAND3X1_36/B DFFSR_14/S
+ OAI21X1
XFILL_6_NAND2X1_280 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_7_OAI21X1_100 INVX1_23/gnd DFFSR_91/S FILL
XFILL_5_DFFSR_153 BUFX2_36/A DFFSR_8/S FILL
XFILL_1_AND2X2_7 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_11_CLKBUF1_11 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_7_DFFSR_55 INVX1_89/gnd DFFSR_36/S FILL
XFILL_24_DFFSR_48 INVX1_4/gnd DFFSR_4/S FILL
XFILL_13_DFFSR_88 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_10_CLKBUF1_14 BUFX2_43/A DFFSR_23/S FILL
XFILL_46_DFFSR_184 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_36_0_1 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_36_DFFSR_187 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_9_CLKBUF1_17 INVX1_94/gnd DFFSR_25/S FILL
XFILL_4_OAI21X1_262 INVX1_89/gnd DFFSR_36/S FILL
XFILL_34_2_2 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_26_DFFSR_190 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_7_DFFSR_2 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_2_INVX1_237 INVX1_8/gnd DFFSR_7/S FILL
XFILL_8_CLKBUF1_20 INVX1_4/gnd DFFSR_51/S FILL
XFILL_6_NAND3X1_112 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_10_DFFPOSX1_16 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_4_INVX1_49 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_21_DFFSR_95 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_32_DFFSR_55 INVX1_89/gnd DFFSR_36/S FILL
XFILL_7_CLKBUF1_23 INVX1_89/gnd DFFSR_2/S FILL
XFILL_43_DFFSR_15 INVX1_8/gnd DFFSR_7/S FILL
XFILL_5_OAI21X1_196 INVX1_94/gnd DFFSR_25/S FILL
XFILL_49_DFFSR_111 INVX1_8/gnd DFFSR_5/S FILL
XFILL_39_DFFSR_114 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_29_DFFSR_117 INVX1_23/gnd DFFSR_91/S FILL
XFILL_5_OR2X2_2 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_3_BUFX2_40 BUFX2_35/A DFFSR_14/S FILL
XFILL_2_DFFSR_190 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_6_OAI21X1_130 INVX1_4/gnd DFFSR_4/S FILL
XFILL_19_DFFSR_120 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_31_DFFSR_6 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_40_DFFSR_62 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_51_DFFSR_22 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_1_INVX1_96 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_0_DFFPOSX1_27 DFFSR_71/gnd DFFSR_45/S FILL
XOAI21X1_166 BUFX2_1/Y INVX1_200/Y NAND2X1_166/Y DFFSR_3/gnd DFFSR_166/D DFFSR_4/S
+ OAI21X1
XFILL_6_NAND2X1_244 INVX1_94/gnd DFFSR_52/S FILL
XFILL_3_INVX1_381 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_7_DFFSR_19 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_5_DFFSR_117 INVX1_23/gnd DFFSR_91/S FILL
XFILL_24_DFFSR_12 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_13_DFFSR_52 INVX1_94/gnd DFFSR_52/S FILL
XFILL_46_DFFSR_148 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_4_OAI21X1_226 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_36_DFFSR_151 BUFX2_7/gnd DFFSR_81/S FILL
XNAND2X1_280 DFFSR_143/Q INVX1_432/Y DFFSR_79/gnd AOI22X1_14/A DFFSR_45/S NAND2X1
XFILL_48_DFFSR_69 BUFX2_43/A DFFSR_23/S FILL
XFILL_26_DFFSR_154 BUFX2_36/A DFFSR_6/S FILL
XFILL_2_INVX1_201 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_16_DFFSR_157 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_1_NAND3X1_1 INVX1_94/gnd DFFSR_25/S FILL
XFILL_10_DFFSR_99 BUFX2_35/A DFFSR_97/S FILL
XFILL_1_NOR2X1_36 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_5_OAI21X1_160 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_32_DFFSR_19 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_4_DFFSR_66 INVX1_2/gnd DFFSR_51/S FILL
XFILL_21_DFFSR_59 INVX1_4/gnd DFFSR_51/S FILL
XNAND3X1_112 INVX1_266/Y INVX1_264/Y INVX1_265/Y DFFSR_71/gnd OAI22X1_9/D DFFSR_10/S
+ NAND3X1
XFILL_0_INVX1_418 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_2_DFFSR_154 BUFX2_36/A DFFSR_6/S FILL
XFILL_43_DFFSR_185 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_5_NAND2X1_274 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_33_DFFSR_188 INVX1_2/gnd DFFSR_1/S FILL
XFILL_23_DFFSR_191 INVX1_23/gnd DFFSR_91/S FILL
XFILL_1_INVX1_60 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_40_DFFSR_26 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_29_DFFSR_66 INVX1_2/gnd DFFSR_51/S FILL
XFILL_3_INVX1_345 INVX1_94/gnd DFFSR_52/S FILL
XFILL_6_NAND2X1_208 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_3_OAI21X1_256 INVX1_2/gnd DFFSR_51/S FILL
XOAI21X1_130 DFFSR_51/S INVX1_147/Y OAI21X1_130/C INVX1_4/gnd DFFSR_130/D DFFSR_4/S
+ OAI21X1
XFILL_13_DFFSR_16 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_5_NAND3X1_106 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_46_DFFSR_112 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_36_DFFSR_115 BUFX2_6/gnd DFFSR_14/S FILL
XNAND2X1_244 NOR2X1_33/Y NOR2X1_32/Y INVX1_94/gnd NAND2X1_244/Y DFFSR_52/S NAND2X1
XFILL_9_DFFSR_188 INVX1_2/gnd DFFSR_1/S FILL
XFILL_4_OAI21X1_190 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_26_DFFSR_118 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_2_INVX1_165 INVX1_23/gnd DFFSR_186/S FILL
XFILL_16_DFFSR_121 BUFX2_36/A DFFSR_6/S FILL
XFILL_48_DFFSR_33 INVX1_94/gnd DFFSR_52/S FILL
XFILL_37_DFFSR_73 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_21_DFFSR_23 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_10_DFFSR_63 INVX1_94/gnd DFFSR_52/S FILL
XFILL_4_DFFSR_30 INVX1_89/gnd DFFSR_36/S FILL
XFILL_5_OAI21X1_124 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_2_BUFX2_1 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_35_3_0 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_0_INVX1_382 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_21_4 INVX1_94/gnd DFFSR_52/S FILL
XFILL_9_OAI22X1_8 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_33_5_1 INVX1_8/gnd DFFSR_7/S FILL
XFILL_2_DFFSR_118 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_43_DFFSR_149 INVX1_23/gnd DFFSR_91/S FILL
XFILL_5_NAND2X1_238 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_45_DFFSR_80 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_33_DFFSR_152 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_23_DFFSR_155 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_29_DFFSR_30 INVX1_89/gnd DFFSR_36/S FILL
XFILL_1_DFFSR_77 INVX1_89/gnd DFFSR_2/S FILL
XFILL_18_DFFSR_70 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_1_INVX1_24 INVX1_2/gnd DFFSR_51/S FILL
XFILL_3_OAI21X1_220 BUFX2_43/A DFFSR_97/S FILL
XFILL_13_DFFSR_158 BUFX2_43/A DFFSR_23/S FILL
XFILL_9_DFFPOSX1_10 INVX1_8/gnd DFFSR_5/S FILL
XFILL_6_NAND2X1_172 BUFX2_36/A DFFSR_6/S FILL
XFILL_3_INVX1_309 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_22_DFFPOSX1_2 INVX1_89/gnd DFFSR_36/S FILL
XFILL_0_BUFX2_15 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_5_XOR2X1_7 INVX1_23/gnd DFFSR_91/S FILL
XFILL_9_DFFSR_152 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_43_DFFSR_9 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_21_DFFPOSX1_5 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_50_DFFSR_183 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_4_OAI21X1_154 BUFX2_37/A DFFSR_8/S FILL
XNAND2X1_208 NAND3X1_55/Y NAND3X1_58/Y BUFX2_8/gnd NAND2X1_208/Y DFFSR_10/S NAND2X1
XFILL_20_DFFPOSX1_8 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_18_DFFPOSX1_29 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_40_DFFSR_186 INVX1_23/gnd DFFSR_186/S FILL
XFILL_9_DFFSR_84 BUFX2_43/A DFFSR_23/S FILL
XFILL_2_INVX1_129 INVX1_89/gnd DFFSR_36/S FILL
XFILL_37_DFFSR_37 INVX1_89/gnd DFFSR_2/S FILL
XFILL_26_DFFSR_77 INVX1_89/gnd DFFSR_2/S FILL
XFILL_30_DFFSR_189 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_4_NAND2X1_268 BUFX2_37/A DFFSR_8/S FILL
XFILL_10_DFFSR_27 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_0_INVX1_346 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_43_0_1 INVX1_4/gnd DFFSR_51/S FILL
XFILL_43_DFFSR_113 INVX1_23/gnd DFFSR_186/S FILL
XFILL_2_OAI21X1_250 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_5_NAND2X1_202 BUFX2_35/A DFFSR_97/S FILL
XFILL_34_DFFSR_84 BUFX2_43/A DFFSR_23/S FILL
XFILL_45_DFFSR_44 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_33_DFFSR_116 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_6_DFFSR_189 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_41_2_2 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_4_NAND3X1_100 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_23_DFFSR_119 BUFX2_37/A DFFSR_81/S FILL
XFILL_13_DFFSR_122 INVX1_94/gnd DFFSR_52/S FILL
XFILL_1_DFFSR_41 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_18_DFFSR_34 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_3_OAI21X1_184 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_6_NAND2X1_136 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_3_AOI21X1_1 INVX1_8/gnd DFFSR_5/S FILL
XFILL_3_INVX1_273 INVX1_8/gnd DFFSR_5/S FILL
XFILL_11_XOR2X1_4 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_42_DFFSR_91 BUFX2_6/gnd DFFSR_91/S FILL
XNAND2X1_172 NAND2X1_172/A BUFX2_36/A BUFX2_36/A NAND2X1_172/Y DFFSR_6/S NAND2X1
XFILL_9_DFFSR_116 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_6_OAI22X1_9 INVX1_8/gnd DFFSR_5/S FILL
XFILL_50_DFFSR_147 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_4_OAI21X1_118 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_15_DFFSR_81 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_40_DFFSR_150 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_26_DFFSR_41 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_9_DFFSR_48 INVX1_4/gnd DFFSR_4/S FILL
XFILL_43_4 INVX1_4/gnd DFFSR_4/S FILL
XFILL_30_DFFSR_153 BUFX2_36/A DFFSR_8/S FILL
XFILL_20_DFFSR_156 INVX1_23/gnd DFFSR_91/S FILL
XFILL_4_NAND2X1_232 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_10_DFFSR_159 BUFX2_36/A DFFSR_6/S FILL
XFILL_3_NAND3X1_130 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_5_NOR2X1_35 INVX1_94/gnd DFFSR_52/S FILL
XFILL_0_INVX1_310 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_50_DFFSR_98 DFFSR_9/gnd DFFSR_9/S FILL
XINVX1_420 BUFX2_31/A INVX1_2/gnd INVX1_420/Y DFFSR_51/S INVX1
XFILL_30_DFFSR_3 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_4_INVX1_417 INVX1_23/gnd DFFSR_91/S FILL
XFILL_2_OAI21X1_214 BUFX2_35/A DFFSR_97/S FILL
XFILL_6_DFFSR_153 BUFX2_36/A DFFSR_8/S FILL
XFILL_6_DFFSR_95 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_34_DFFSR_48 INVX1_4/gnd DFFSR_4/S FILL
XFILL_23_DFFSR_88 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_5_NAND2X1_166 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_47_DFFSR_184 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_37_DFFSR_187 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_5_BUFX2_33 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_3_OAI21X1_148 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_17_DFFPOSX1_23 INVX1_23/gnd DFFSR_91/S FILL
XFILL_10_DFFPOSX1_2 INVX1_89/gnd DFFSR_36/S FILL
XFILL_27_DFFSR_190 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_6_NAND2X1_100 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_3_INVX1_237 INVX1_8/gnd DFFSR_7/S FILL
XFILL_9_DFFPOSX1_5 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_31_DFFSR_95 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_8_DFFPOSX1_8 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_42_DFFSR_55 INVX1_89/gnd DFFSR_36/S FILL
XFILL_3_INVX1_89 INVX1_89/gnd DFFSR_2/S FILL
XFILL_3_NAND2X1_262 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_8_AOI21X1_28 DFFSR_71/gnd DFFSR_10/S FILL
XNAND2X1_136 DFFSR_5/S NAND2X1_72/B DFFSR_5/gnd NAND2X1_136/Y DFFSR_2/S NAND2X1
XFILL_50_DFFSR_111 INVX1_8/gnd DFFSR_5/S FILL
XFILL_7_AOI21X1_31 INVX1_23/gnd DFFSR_186/S FILL
XFILL_9_DFFSR_12 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_40_DFFSR_114 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_27_DFFPOSX1_12 INVX1_8/gnd DFFSR_5/S FILL
XFILL_30_DFFSR_117 INVX1_23/gnd DFFSR_91/S FILL
XFILL_15_0_2 BUFX2_37/A DFFSR_81/S FILL
XFILL_15_DFFSR_45 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_3_DFFSR_190 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_6_AOI21X1_34 INVX1_94/gnd DFFSR_25/S FILL
XFILL_1_OAI21X1_244 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_20_DFFSR_120 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_10_DFFSR_123 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_4_NAND2X1_196 BUFX2_7/gnd DFFSR_54/S FILL
XAOI21X1_34 NAND3X1_86/Y NAND3X1_87/Y INVX1_250/Y INVX1_94/gnd AOI21X1_35/C DFFSR_25/S
+ AOI21X1
XFILL_5_AOI21X1_37 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_50_DFFSR_62 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_0_AOI21X1_2 INVX1_94/gnd DFFSR_52/S FILL
XINVX1_384 INVX1_116/A DFFSR_5/gnd INVX1_384/Y DFFSR_5/S INVX1
XFILL_0_INVX1_274 INVX1_8/gnd DFFSR_5/S FILL
XFILL_4_AOI21X1_40 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_3_AOI21X1_43 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_2_OAI21X1_178 INVX1_94/gnd DFFSR_25/S FILL
XFILL_2_AOI21X1_46 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_12_DFFSR_92 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_6_DFFSR_117 INVX1_23/gnd DFFSR_91/S FILL
XFILL_34_DFFSR_12 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_23_DFFSR_52 INVX1_94/gnd DFFSR_52/S FILL
XFILL_6_DFFSR_59 INVX1_4/gnd DFFSR_51/S FILL
XFILL_5_NAND2X1_130 INVX1_4/gnd DFFSR_4/S FILL
XFILL_47_DFFSR_148 DFFSR_89/gnd DFFSR_92/S FILL
XBUFX2_37 BUFX2_37/A BUFX2_37/A BUFX2_37/Y DFFSR_81/S BUFX2
XFILL_37_DFFSR_151 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_27_DFFSR_154 BUFX2_36/A DFFSR_6/S FILL
XFILL_3_INVX1_201 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_3_OAI21X1_112 INVX1_4/gnd DFFSR_4/S FILL
XFILL_42_3_0 INVX1_4/gnd DFFSR_4/S FILL
XFILL_17_DFFSR_157 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_8_OAI21X1_76 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_48_9 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_6_NAND2X1_97 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_2_NAND3X1_1 INVX1_94/gnd DFFSR_25/S FILL
XFILL_7_OAI21X1_79 INVX1_89/gnd DFFSR_36/S FILL
XNAND2X1_100 BUFX2_25/Y DFFSR_92/Q BUFX2_6/gnd OAI21X1_100/C DFFSR_14/S NAND2X1
XFILL_20_DFFSR_99 BUFX2_35/A DFFSR_97/S FILL
XFILL_3_NAND2X1_226 BUFX2_36/A DFFSR_6/S FILL
XFILL_2_NOR2X1_36 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_3_INVX1_53 INVX1_89/gnd DFFSR_2/S FILL
XFILL_42_DFFSR_19 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_6_OAI21X1_82 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_31_DFFSR_59 INVX1_4/gnd DFFSR_51/S FILL
XFILL_40_5_1 DFFSR_3/gnd DFFSR_65/S FILL
XNAND2X1_97 DFFSR_89/Q BUFX2_20/Y BUFX2_5/gnd OAI21X1_97/C DFFSR_23/S NAND2X1
XFILL_5_OAI21X1_85 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_3_DFFSR_154 BUFX2_36/A DFFSR_6/S FILL
XFILL_2_NAND3X1_124 DFFSR_5/gnd DFFSR_5/S FILL
XOAI21X1_82 BUFX2_18/Y INVX1_93/Y NAND2X1_82/Y DFFSR_9/gnd DFFSR_82/D DFFSR_9/S OAI21X1
XFILL_4_OAI21X1_88 INVX1_4/gnd DFFSR_4/S FILL
XFILL_1_INVX1_418 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_44_DFFSR_185 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_3_OAI21X1_91 BUFX2_43/A DFFSR_97/S FILL
XFILL_1_OAI21X1_208 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_4_NAND2X1_160 INVX1_8/gnd DFFSR_5/S FILL
XFILL_34_DFFSR_188 INVX1_2/gnd DFFSR_1/S FILL
XFILL_24_DFFSR_191 INVX1_23/gnd DFFSR_91/S FILL
XFILL_2_OAI21X1_94 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_1_OAI21X1_97 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_0_INVX1_238 BUFX2_37/A DFFSR_81/S FILL
XFILL_50_DFFSR_26 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_39_DFFSR_66 INVX1_2/gnd DFFSR_51/S FILL
XINVX1_348 DFFSR_67/Q INVX1_4/gnd INVX1_348/Y DFFSR_4/S INVX1
XFILL_16_DFFPOSX1_17 BUFX2_37/A DFFSR_8/S FILL
XFILL_2_AOI21X1_10 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_6_DFFSR_23 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_2_OAI21X1_142 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_23_DFFSR_16 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_1_AOI21X1_13 INVX1_8/gnd DFFSR_7/S FILL
XFILL_12_DFFSR_56 INVX1_2/gnd DFFSR_51/S FILL
XFILL_0_AOI21X1_16 BUFX2_43/A DFFSR_23/S FILL
XFILL_47_DFFSR_112 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_37_DFFSR_115 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_0_DFFSR_191 INVX1_23/gnd DFFSR_91/S FILL
XFILL_5_NOR2X1_4 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_2_NAND2X1_256 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_27_DFFSR_118 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_3_INVX1_165 INVX1_23/gnd DFFSR_186/S FILL
XFILL_42_DFFSR_6 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_17_DFFSR_121 BUFX2_36/A DFFSR_6/S FILL
XFILL_9_OAI21X1_37 INVX1_89/gnd DFFSR_2/S FILL
XFILL_47_DFFSR_73 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_8_OAI21X1_40 INVX1_8/gnd DFFSR_7/S FILL
XFILL_31_DFFSR_23 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_6_NAND2X1_61 BUFX2_37/A DFFSR_81/S FILL
XFILL_0_OAI21X1_238 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_20_DFFSR_63 INVX1_94/gnd DFFSR_52/S FILL
XFILL_7_OAI21X1_43 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_3_INVX1_17 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_3_DFFSR_70 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_3_NAND2X1_190 BUFX2_35/A DFFSR_97/S FILL
XNAND2X1_61 DFFSR_81/S DFFSR_53/Q BUFX2_37/A OAI21X1_61/C DFFSR_81/S NAND2X1
XFILL_6_OAI21X1_46 BUFX2_37/A DFFSR_81/S FILL
XFILL_48_2_2 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_6_DFFPOSX1_28 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_5_NAND2X1_64 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_1_INVX1_382 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_25_1 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_4_NAND2X1_67 INVX1_2/gnd DFFSR_1/S FILL
XFILL_5_OAI21X1_49 DFFSR_73/gnd DFFSR_11/S FILL
XOAI21X1_46 DFFSR_81/S INVX1_52/Y OAI21X1_46/C BUFX2_37/A DFFSR_46/D DFFSR_81/S OAI21X1
XFILL_4_OAI21X1_52 INVX1_94/gnd DFFSR_25/S FILL
XFILL_3_NAND2X1_70 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_3_DFFSR_118 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_44_DFFSR_149 INVX1_23/gnd DFFSR_91/S FILL
XFILL_1_OAI21X1_172 BUFX2_36/A DFFSR_6/S FILL
XFILL_3_OAI21X1_55 INVX1_89/gnd DFFSR_2/S FILL
XFILL_2_NAND2X1_73 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_34_DFFSR_152 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_1_NAND2X1_76 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_4_NAND2X1_124 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_2_OAI21X1_58 DFFSR_3/gnd DFFSR_65/S FILL
XINVX1_312 DFFSR_6/Q BUFX2_36/A INVX1_312/Y DFFSR_6/S INVX1
XFILL_1_OAI21X1_61 BUFX2_36/A DFFSR_8/S FILL
XFILL_0_INVX1_202 BUFX2_37/A DFFSR_81/S FILL
XFILL_0_INVX1_64 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_24_DFFSR_155 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_39_DFFSR_30 INVX1_89/gnd DFFSR_36/S FILL
XFILL_0_NAND2X1_79 INVX1_89/gnd DFFSR_36/S FILL
XFILL_28_DFFSR_70 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_14_DFFSR_158 BUFX2_43/A DFFSR_23/S FILL
XFILL_16_1_0 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_0_OAI21X1_64 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_1_NAND2X1_286 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_4_INVX1_309 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_2_OAI21X1_106 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_12_DFFSR_20 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_14_3_1 BUFX2_37/A DFFSR_8/S FILL
XNOR2X1_8 NOR2X1_8/A NOR2X1_9/A BUFX2_43/A NOR2X1_8/Y DFFSR_23/S NOR2X1
XFILL_0_DFFSR_155 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_3_NOR3X1_1 INVX1_94/gnd DFFSR_52/S FILL
XFILL_41_DFFSR_186 INVX1_23/gnd DFFSR_186/S FILL
XFILL_2_NAND2X1_220 BUFX2_35/A DFFSR_14/S FILL
XFILL_12_5_2 BUFX2_36/A DFFSR_6/S FILL
XFILL_3_INVX1_129 INVX1_89/gnd DFFSR_36/S FILL
XFILL_1_NAND3X1_118 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_47_DFFSR_37 INVX1_89/gnd DFFSR_2/S FILL
XFILL_36_DFFSR_77 INVX1_89/gnd DFFSR_2/S FILL
XFILL_31_DFFSR_189 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_6_NAND2X1_25 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_0_OAI21X1_202 BUFX2_35/A DFFSR_14/S FILL
XFILL_3_NAND2X1_154 BUFX2_37/A DFFSR_8/S FILL
XFILL_5_NAND2X1_28 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_6_OAI21X1_10 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_20_DFFSR_27 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_3_DFFSR_34 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_4_NAND2X1_31 BUFX2_43/A DFFSR_97/S FILL
XNAND2X1_25 DFFSR_17/Q DFFSR_45/S DFFSR_79/gnd OAI21X1_25/C DFFSR_45/S NAND2X1
XFILL_1_INVX1_346 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_5_OAI21X1_13 BUFX2_16/gnd DFFSR_65/S FILL
XOAI21X1_10 DFFSR_44/S INVX1_12/Y OAI21X1_10/C DFFSR_71/gnd DFFSR_10/D DFFSR_45/S
+ OAI21X1
XFILL_4_OAI21X1_16 INVX1_89/gnd DFFSR_36/S FILL
XFILL_3_NAND2X1_34 INVX1_2/gnd DFFSR_1/S FILL
XFILL_44_DFFSR_113 INVX1_23/gnd DFFSR_186/S FILL
XFILL_2_NAND2X1_37 INVX1_8/gnd DFFSR_5/S FILL
XFILL_9_DFFSR_9 DFFSR_9/gnd DFFSR_9/S FILL
XDFFPOSX1_28 NAND2X1_224/B CLKBUF1_10/Y NAND2X1_284/Y DFFSR_3/gnd DFFSR_65/S DFFPOSX1
XFILL_44_DFFSR_84 BUFX2_43/A DFFSR_23/S FILL
XFILL_1_OAI21X1_136 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_34_DFFSR_116 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_7_DFFSR_189 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_3_OAI21X1_19 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_15_DFFPOSX1_11 INVX1_4/gnd DFFSR_4/S FILL
XFILL_8_NAND3X1_96 BUFX2_43/A DFFSR_97/S FILL
XFILL_24_DFFSR_119 BUFX2_37/A DFFSR_81/S FILL
XFILL_2_OAI21X1_22 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_1_NAND2X1_40 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_0_INVX1_166 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_7_NAND3X1_99 BUFX2_6/gnd DFFSR_14/S FILL
XAOI21X1_4 AOI21X1_4/A AOI21X1_4/B AOI21X1_4/C BUFX2_7/gnd AOI21X1_4/Y DFFSR_81/S
+ AOI21X1
XFILL_0_DFFSR_81 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_0_INVX1_28 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_14_DFFSR_122 INVX1_94/gnd DFFSR_52/S FILL
XFILL_1_OAI21X1_25 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_0_NAND2X1_43 INVX1_89/gnd DFFSR_2/S FILL
XINVX1_276 INVX1_21/A DFFSR_1/gnd INVX1_276/Y DFFSR_1/S INVX1
XFILL_28_DFFSR_34 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_17_DFFSR_74 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_0_OAI21X1_28 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_4_AOI21X1_1 INVX1_8/gnd DFFSR_5/S FILL
XFILL_1_NAND2X1_250 INVX1_8/gnd DFFSR_5/S FILL
XFILL_22_0_2 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_7_OAI22X1_9 INVX1_8/gnd DFFSR_5/S FILL
XFILL_2_NAND2X1_184 BUFX2_37/A DFFSR_8/S FILL
XFILL_0_DFFSR_119 BUFX2_37/A DFFSR_81/S FILL
XFILL_5_DFFPOSX1_22 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_25_DFFSR_81 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_41_DFFSR_150 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_36_DFFSR_41 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_47_1 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_8_DFFSR_88 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_2_1_2 INVX1_23/gnd DFFSR_186/S FILL
XFILL_31_DFFSR_153 BUFX2_36/A DFFSR_8/S FILL
XFILL_21_DFFSR_156 INVX1_23/gnd DFFSR_91/S FILL
XFILL_0_OAI21X1_166 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_3_AOI22X1_12 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_9_OAI21X1_221 BUFX2_35/A DFFSR_14/S FILL
XFILL_11_DFFSR_159 BUFX2_36/A DFFSR_6/S FILL
XFILL_3_NAND2X1_118 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_6_NOR2X1_35 INVX1_94/gnd DFFSR_52/S FILL
XFILL_1_INVX1_310 DFFSR_79/gnd DFFSR_36/S FILL
XINVX1_2 INVX1_2/A INVX1_2/gnd INVX1_2/Y DFFSR_51/S INVX1
XFILL_1_OAI21X1_100 INVX1_23/gnd DFFSR_91/S FILL
XFILL_7_DFFSR_153 BUFX2_36/A DFFSR_8/S FILL
XFILL_10_OAI22X1_39 BUFX2_37/A DFFSR_8/S FILL
XFILL_0_NAND2X1_280 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_44_DFFSR_48 INVX1_4/gnd DFFSR_4/S FILL
XFILL_33_DFFSR_88 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_24_DFFPOSX1_30 BUFX2_43/A DFFSR_97/S FILL
XFILL_9_NAND3X1_57 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_48_DFFSR_184 DFFSR_1/gnd DFFSR_9/S FILL
XINVX1_240 AND2X2_9/B BUFX2_35/A INVX1_240/Y DFFSR_14/S INVX1
XFILL_0_INVX1_130 BUFX2_36/A DFFSR_6/S FILL
XFILL_8_NAND3X1_60 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_0_DFFSR_45 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_9_OAI22X1_42 INVX1_8/gnd DFFSR_7/S FILL
XFILL_38_DFFSR_187 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_7_NAND3X1_63 BUFX2_43/A DFFSR_23/S FILL
XFILL_8_OAI22X1_45 INVX1_89/gnd DFFSR_2/S FILL
XFILL_17_DFFSR_38 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_47_5_1 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_28_DFFSR_190 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_6_NAND3X1_66 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_1_NAND2X1_214 BUFX2_35/A DFFSR_97/S FILL
XFILL_7_OAI22X1_48 BUFX2_37/A DFFSR_81/S FILL
XFILL_5_NAND3X1_69 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_6_OAI22X1_51 BUFX2_7/gnd DFFSR_81/S FILL
XNAND3X1_66 INVX1_248/A INVX1_249/Y NAND3X1_66/C BUFX2_6/gnd NAND3X1_66/Y DFFSR_14/S
+ NAND3X1
XFILL_4_NAND3X1_72 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_10_XOR2X1_8 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_5_OAI22X1_54 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_0_NAND3X1_112 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_41_DFFSR_95 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_3_NAND3X1_75 BUFX2_35/A DFFSR_97/S FILL
XOAI22X1_51 INVX1_361/Y OAI22X1_39/B INVX1_360/Y OAI22X1_39/D BUFX2_7/gnd NOR2X1_35/A
+ DFFSR_81/S OAI22X1
XFILL_51_DFFSR_111 INVX1_8/gnd DFFSR_5/S FILL
XFILL_4_OAI22X1_57 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_8_OAI21X1_251 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_2_NAND2X1_148 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_2_NAND3X1_78 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_2_AND2X2_4 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_8_DFFSR_52 INVX1_94/gnd DFFSR_52/S FILL
XFILL_41_DFFSR_114 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_3_OAI22X1_60 INVX1_8/gnd DFFSR_5/S FILL
XFILL_31_DFFSR_117 INVX1_23/gnd DFFSR_91/S FILL
XFILL_1_NAND3X1_81 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_2_OAI22X1_63 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_14_DFFSR_85 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_25_DFFSR_45 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_4_DFFSR_190 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_0_NAND3X1_84 INVX1_94/gnd DFFSR_25/S FILL
XFILL_1_OAI22X1_66 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_21_DFFSR_120 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_11_DFFSR_123 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_0_OAI21X1_130 INVX1_4/gnd DFFSR_4/S FILL
XFILL_1_AOI21X1_2 INVX1_94/gnd DFFSR_52/S FILL
XFILL_1_INVX1_274 INVX1_8/gnd DFFSR_5/S FILL
XFILL_20_DFFSR_7 INVX1_8/gnd DFFSR_7/S FILL
XINVX1_86 DFFSR_76/Q BUFX2_19/gnd INVX1_86/Y DFFSR_52/S INVX1
XFILL_0_NAND2X1_244 INVX1_94/gnd DFFSR_52/S FILL
XFILL_22_DFFSR_92 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_7_DFFSR_117 INVX1_23/gnd DFFSR_91/S FILL
XFILL_44_DFFSR_12 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_5_DFFSR_99 BUFX2_35/A DFFSR_97/S FILL
XFILL_9_NAND3X1_21 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_33_DFFSR_52 INVX1_94/gnd DFFSR_52/S FILL
XFILL_48_DFFSR_148 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_8_NAND3X1_24 BUFX2_37/A DFFSR_8/S FILL
XFILL_4_BUFX2_8 BUFX2_8/gnd DFFSR_10/S FILL
XINVX1_204 AND2X2_6/A BUFX2_36/A INVX1_204/Y DFFSR_8/S INVX1
XFILL_7_NAND3X1_27 BUFX2_37/A DFFSR_81/S FILL
XFILL_38_DFFSR_151 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_4_DFFPOSX1_16 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_28_DFFSR_154 BUFX2_36/A DFFSR_6/S FILL
XFILL_4_BUFX2_37 BUFX2_37/A DFFSR_81/S FILL
XFILL_4_INVX1_201 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_1_NAND2X1_178 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_18_DFFSR_157 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_6_NAND3X1_30 INVX1_94/gnd DFFSR_52/S FILL
XFILL_7_OAI22X1_12 INVX1_4/gnd DFFSR_51/S FILL
XNAND3X1_30 AOI22X1_4/D AOI22X1_4/C AOI21X1_9/Y INVX1_94/gnd NAND3X1_30/Y DFFSR_52/S
+ NAND3X1
XFILL_3_NAND3X1_1 INVX1_94/gnd DFFSR_25/S FILL
XFILL_5_NAND3X1_33 INVX1_8/gnd DFFSR_7/S FILL
XFILL_6_OAI22X1_15 INVX1_4/gnd DFFSR_4/S FILL
XFILL_41_DFFSR_3 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_4_NAND3X1_36 BUFX2_35/A DFFSR_97/S FILL
XFILL_30_DFFSR_99 BUFX2_35/A DFFSR_97/S FILL
XFILL_9_NAND3X1_131 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_5_OAI22X1_18 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_3_NOR2X1_36 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_2_INVX1_93 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_41_DFFSR_59 INVX1_4/gnd DFFSR_51/S FILL
XOAI22X1_15 INVX1_286/Y OAI22X1_7/B INVX1_285/Y OAI22X1_7/D INVX1_4/gnd NOR2X1_17/B
+ DFFSR_4/S OAI22X1
XDFFSR_157 DFFSR_157/Q CLKBUF1_12/Y DFFSR_157/R DFFSR_91/S DFFSR_157/D BUFX2_6/gnd
+ DFFSR_91/S DFFSR
XFILL_8_OAI21X1_215 BUFX2_43/A DFFSR_97/S FILL
XFILL_3_NAND3X1_39 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_2_NAND2X1_112 INVX1_4/gnd DFFSR_4/S FILL
XFILL_4_OAI22X1_21 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_2_NAND3X1_42 BUFX2_43/A DFFSR_23/S FILL
XFILL_4_DFFSR_154 BUFX2_36/A DFFSR_6/S FILL
XFILL_8_DFFSR_16 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_3_OAI22X1_24 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_2_INVX1_418 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_14_DFFSR_49 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_45_DFFSR_185 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_1_NAND3X1_45 BUFX2_35/A DFFSR_97/S FILL
XFILL_23_1_0 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_2_OAI22X1_27 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_0_NAND3X1_48 BUFX2_43/A DFFSR_23/S FILL
XFILL_1_OAI22X1_30 INVX1_94/gnd DFFSR_25/S FILL
XFILL_35_DFFSR_188 INVX1_2/gnd DFFSR_1/S FILL
XFILL_25_DFFSR_191 INVX1_23/gnd DFFSR_91/S FILL
XFILL_23_DFFPOSX1_24 BUFX2_43/A DFFSR_23/S FILL
XFILL_0_OAI22X1_33 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_1_INVX1_238 BUFX2_37/A DFFSR_81/S FILL
XFILL_21_3_1 INVX1_94/gnd DFFSR_25/S FILL
XFILL_49_DFFSR_66 INVX1_2/gnd DFFSR_51/S FILL
XFILL_3_2_0 INVX1_23/gnd DFFSR_91/S FILL
XFILL_19_5_2 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_5_DFFSR_63 INVX1_94/gnd DFFSR_52/S FILL
XINVX1_50 INVX1_50/A BUFX2_8/gnd INVX1_50/Y DFFSR_25/S INVX1
XFILL_0_NAND2X1_208 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_33_DFFSR_16 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_11_DFFSR_96 INVX1_2/gnd DFFSR_1/S FILL
XFILL_22_DFFSR_56 INVX1_2/gnd DFFSR_51/S FILL
XFILL_1_4_1 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_48_DFFSR_112 DFFSR_3/gnd DFFSR_65/S FILL
XINVX1_168 INVX1_168/A DFFSR_89/gnd INVX1_168/Y DFFSR_92/S INVX1
XFILL_38_DFFSR_115 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_1_DFFSR_191 INVX1_23/gnd DFFSR_91/S FILL
XFILL_28_DFFSR_118 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_4_INVX1_165 INVX1_23/gnd DFFSR_186/S FILL
XFILL_18_DFFSR_121 BUFX2_36/A DFFSR_6/S FILL
XFILL_1_NAND2X1_142 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_7_OAI21X1_245 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_41_DFFSR_23 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_30_DFFSR_63 INVX1_94/gnd DFFSR_52/S FILL
XFILL_2_INVX1_57 BUFX2_17/gnd DFFSR_57/S FILL
XDFFSR_121 DFFSR_121/Q CLKBUF1_6/Y DFFSR_123/R DFFSR_6/S DFFSR_121/D BUFX2_36/A DFFSR_6/S
+ DFFSR
XFILL_2_INVX1_382 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_8_OAI21X1_179 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_14_DFFSR_13 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_4_DFFSR_118 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_45_DFFSR_149 INVX1_23/gnd DFFSR_91/S FILL
XFILL_0_NAND3X1_12 INVX1_94/gnd DFFSR_52/S FILL
XFILL_35_DFFSR_152 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_8_DFFSR_6 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_1_INVX1_202 BUFX2_37/A DFFSR_81/S FILL
XFILL_25_DFFSR_155 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_49_DFFSR_30 INVX1_89/gnd DFFSR_36/S FILL
XFILL_15_DFFSR_158 BUFX2_43/A DFFSR_23/S FILL
XFILL_29_0_2 INVX1_89/gnd DFFSR_2/S FILL
XFILL_38_DFFSR_70 BUFX2_17/gnd DFFSR_57/S FILL
XINVX1_14 DFFSR_12/Q BUFX2_35/A INVX1_14/Y DFFSR_14/S INVX1
XFILL_0_NAND2X1_172 BUFX2_36/A DFFSR_6/S FILL
XFILL_0_NAND3X1_2 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_3_DFFPOSX1_10 INVX1_8/gnd DFFSR_5/S FILL
XDFFSR_67 DFFSR_67/Q CLKBUF1_2/Y DFFSR_68/R DFFSR_51/S DFFSR_67/D INVX1_2/gnd DFFSR_51/S
+ DFFSR
XFILL_22_DFFSR_20 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_11_DFFSR_60 BUFX2_37/A DFFSR_8/S FILL
XFILL_0_NOR2X1_37 INVX1_94/gnd DFFSR_25/S FILL
XFILL_5_DFFSR_27 DFFSR_1/gnd DFFSR_1/S FILL
XINVX1_132 DFFSR_117/Q BUFX2_35/A INVX1_132/Y DFFSR_97/S INVX1
XFILL_4_NOR2X1_8 BUFX2_43/A DFFSR_23/S FILL
XFILL_9_1_2 BUFX2_43/A DFFSR_23/S FILL
XFILL_1_DFFSR_155 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_8_NAND3X1_125 INVX1_8/gnd DFFSR_5/S FILL
XFILL_42_DFFSR_186 INVX1_23/gnd DFFSR_186/S FILL
XFILL_4_INVX1_129 INVX1_89/gnd DFFSR_36/S FILL
XFILL_7_OAI21X1_209 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_12_DFFPOSX1_29 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_1_NAND2X1_106 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_46_DFFSR_77 INVX1_89/gnd DFFSR_2/S FILL
XFILL_32_DFFSR_189 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_30_DFFSR_27 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_2_INVX1_21 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_2_DFFSR_74 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_19_DFFSR_67 INVX1_2/gnd DFFSR_51/S FILL
XFILL_22_DFFPOSX1_18 BUFX2_37/A DFFSR_8/S FILL
XFILL_8_OAI21X1_143 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_2_INVX1_346 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_6_XOR2X1_4 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_45_DFFSR_113 INVX1_23/gnd DFFSR_186/S FILL
XFILL_1_BUFX2_12 BUFX2_37/A DFFSR_81/S FILL
XFILL_35_DFFSR_116 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_8_DFFSR_189 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_25_DFFSR_119 BUFX2_37/A DFFSR_81/S FILL
XFILL_1_INVX1_166 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_15_DFFSR_122 INVX1_94/gnd DFFSR_52/S FILL
XFILL_38_DFFSR_34 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_27_DFFSR_74 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_5_AOI21X1_1 INVX1_8/gnd DFFSR_5/S FILL
XDFFSR_31 INVX1_35/A DFFSR_20/CLK DFFSR_31/R DFFSR_97/S DFFSR_31/D BUFX2_35/A DFFSR_97/S
+ DFFSR
XFILL_0_NAND2X1_136 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_6_OAI21X1_239 INVX1_4/gnd DFFSR_4/S FILL
XFILL_11_DFFSR_24 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_8_OAI22X1_9 INVX1_8/gnd DFFSR_5/S FILL
XFILL_1_DFFSR_119 BUFX2_37/A DFFSR_81/S FILL
XFILL_34_3 INVX1_8/gnd DFFSR_7/S FILL
XFILL_7_OAI21X1_173 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_35_DFFSR_81 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_42_DFFSR_150 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_46_DFFSR_41 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_32_DFFSR_153 BUFX2_36/A DFFSR_8/S FILL
XFILL_22_DFFSR_156 INVX1_23/gnd DFFSR_91/S FILL
XFILL_19_DFFSR_31 BUFX2_35/A DFFSR_97/S FILL
XFILL_2_DFFSR_38 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_12_DFFSR_159 BUFX2_36/A DFFSR_6/S FILL
XFILL_8_OAI21X1_107 BUFX2_36/A DFFSR_6/S FILL
XFILL_2_INVX1_310 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_20_CLKBUF1_21 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_19_CLKBUF1_24 INVX1_23/gnd DFFSR_186/S FILL
XFILL_8_DFFSR_153 BUFX2_36/A DFFSR_8/S FILL
XFILL_12_XOR2X1_1 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_19_DFFSR_4 INVX1_4/gnd DFFSR_4/S FILL
XFILL_43_DFFSR_88 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_49_DFFSR_184 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_1_INVX1_130 BUFX2_36/A DFFSR_6/S FILL
XFILL_39_DFFSR_187 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_7_NAND3X1_119 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_27_DFFSR_38 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_16_DFFSR_78 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_29_DFFSR_190 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_11_DFFPOSX1_23 INVX1_23/gnd DFFSR_91/S FILL
XFILL_0_NAND2X1_100 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_3_BUFX2_5 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_6_OAI21X1_203 BUFX2_35/A DFFSR_14/S FILL
XFILL_30_1_0 DFFSR_5/gnd DFFSR_2/S FILL
XOAI21X1_239 INVX1_397/A INVX1_331/A AOI21X1_40/Y INVX1_4/gnd DFFPOSX1_11/D DFFSR_4/S
+ OAI21X1
XFILL_7_OAI21X1_137 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_42_DFFSR_114 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_21_DFFPOSX1_12 INVX1_8/gnd DFFSR_5/S FILL
XFILL_7_DFFSR_92 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_32_DFFSR_117 INVX1_23/gnd DFFSR_91/S FILL
XFILL_24_DFFSR_85 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_35_DFFSR_45 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_28_3_1 INVX1_89/gnd DFFSR_36/S FILL
XFILL_5_DFFSR_190 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_22_DFFSR_120 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_12_DFFSR_123 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_26_5_2 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_2_AOI21X1_2 INVX1_94/gnd DFFSR_52/S FILL
XFILL_6_BUFX2_30 INVX1_4/gnd DFFSR_51/S FILL
XFILL_8_4_1 BUFX2_43/A DFFSR_97/S FILL
XFILL_2_INVX1_274 INVX1_8/gnd DFFSR_5/S FILL
XFILL_32_DFFSR_92 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_8_DFFSR_117 INVX1_23/gnd DFFSR_91/S FILL
XFILL_5_OAI21X1_233 BUFX2_36/A DFFSR_8/S FILL
XFILL_4_INVX1_86 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_43_DFFSR_52 INVX1_94/gnd DFFSR_52/S FILL
XFILL_49_DFFSR_148 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_39_DFFSR_151 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_16_DFFSR_42 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_29_DFFSR_154 BUFX2_36/A DFFSR_6/S FILL
XNAND3X1_4 NAND3X1_4/A NAND3X1_4/B NAND3X1_3/Y INVX1_94/gnd NAND3X1_4/Y DFFSR_52/S
+ NAND3X1
XFILL_19_DFFSR_157 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_6_OAI21X1_167 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_4_NAND3X1_1 INVX1_94/gnd DFFSR_25/S FILL
XNOR2X1_39 NOR2X1_39/A NOR2X1_39/B INVX1_8/gnd NOR2X1_39/Y DFFSR_5/S NOR2X1
XFILL_40_DFFSR_99 BUFX2_35/A DFFSR_97/S FILL
XFILL_4_NOR2X1_36 BUFX2_8/gnd DFFSR_10/S FILL
XOAI21X1_203 INVX1_226/Y INVX1_240/Y AND2X2_8/Y BUFX2_35/A NAND3X1_36/C DFFSR_14/S
+ OAI21X1
XFILL_13_DFFSR_89 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_11_CLKBUF1_12 BUFX2_43/A DFFSR_23/S FILL
XFILL_1_AND2X2_8 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_5_DFFSR_154 BUFX2_36/A DFFSR_6/S FILL
XFILL_6_NAND2X1_281 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_7_OAI21X1_101 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_7_DFFSR_56 INVX1_2/gnd DFFSR_51/S FILL
XFILL_3_INVX1_418 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_24_DFFSR_49 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_46_DFFSR_185 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_10_CLKBUF1_15 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_36_0_2 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_36_DFFSR_188 INVX1_2/gnd DFFSR_1/S FILL
XFILL_26_DFFSR_191 INVX1_23/gnd DFFSR_91/S FILL
XFILL_4_OAI21X1_263 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_2_INVX1_238 BUFX2_37/A DFFSR_81/S FILL
XFILL_9_CLKBUF1_18 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_7_DFFSR_3 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_6_NAND3X1_113 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_8_CLKBUF1_21 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_7_CLKBUF1_24 INVX1_23/gnd DFFSR_186/S FILL
XFILL_10_DFFPOSX1_17 BUFX2_37/A DFFSR_8/S FILL
XFILL_4_INVX1_50 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_43_DFFSR_16 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_21_DFFSR_96 INVX1_2/gnd DFFSR_1/S FILL
XFILL_32_DFFSR_56 INVX1_2/gnd DFFSR_51/S FILL
XFILL_5_OAI21X1_197 INVX1_8/gnd DFFSR_7/S FILL
XFILL_49_DFFSR_112 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_39_DFFSR_115 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_2_DFFSR_191 INVX1_23/gnd DFFSR_91/S FILL
XFILL_5_OR2X2_3 BUFX2_43/A DFFSR_23/S FILL
XFILL_3_BUFX2_41 BUFX2_37/A DFFSR_81/S FILL
XFILL_29_DFFSR_118 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_19_DFFSR_121 BUFX2_36/A DFFSR_6/S FILL
XFILL_31_DFFSR_7 INVX1_8/gnd DFFSR_7/S FILL
XFILL_6_OAI21X1_131 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_40_DFFSR_63 INVX1_94/gnd DFFSR_52/S FILL
XFILL_1_INVX1_97 INVX1_4/gnd DFFSR_4/S FILL
XOAI21X1_167 BUFX2_4/Y INVX1_201/Y OAI21X1_167/C BUFX2_8/gnd DFFSR_167/D DFFSR_25/S
+ OAI21X1
XFILL_0_DFFPOSX1_28 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_3_INVX1_382 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_6_NAND2X1_245 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_7_DFFSR_20 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_13_DFFSR_53 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_24_DFFSR_13 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_5_DFFSR_118 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_46_DFFSR_149 INVX1_23/gnd DFFSR_91/S FILL
XFILL_4_OAI21X1_227 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_36_DFFSR_152 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_6_NOR2X1_1 BUFX2_36/A DFFSR_6/S FILL
XNAND2X1_281 DFFSR_135/Q NOR2X1_53/B DFFSR_79/gnd AOI22X1_14/B DFFSR_45/S NAND2X1
XFILL_2_INVX1_202 BUFX2_37/A DFFSR_81/S FILL
XFILL_26_DFFSR_155 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_16_DFFSR_158 BUFX2_43/A DFFSR_23/S FILL
XFILL_48_DFFSR_70 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_1_NAND3X1_2 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_32_DFFSR_20 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_5_OAI21X1_161 INVX1_23/gnd DFFSR_186/S FILL
XFILL_21_DFFSR_60 BUFX2_37/A DFFSR_8/S FILL
XFILL_1_NOR2X1_37 INVX1_94/gnd DFFSR_25/S FILL
XFILL_4_DFFSR_67 INVX1_2/gnd DFFSR_51/S FILL
XNAND3X1_113 NOR2X1_1/A INVX1_266/Y INVX1_265/Y BUFX2_8/gnd OAI22X1_6/D DFFSR_10/S
+ NAND3X1
XFILL_2_DFFSR_155 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_0_INVX1_419 INVX1_2/gnd DFFSR_51/S FILL
XFILL_43_DFFSR_186 INVX1_23/gnd DFFSR_186/S FILL
XFILL_5_NAND2X1_275 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_33_DFFSR_189 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_1_INVX1_61 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_40_DFFSR_27 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_29_DFFSR_67 INVX1_2/gnd DFFSR_51/S FILL
XOAI21X1_131 DFFSR_9/S INVX1_148/Y NAND2X1_131/Y DFFSR_9/gnd DFFSR_131/D DFFSR_9/S
+ OAI21X1
XFILL_3_OAI21X1_257 INVX1_2/gnd DFFSR_51/S FILL
XFILL_6_NAND2X1_209 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_13_DFFSR_17 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_3_INVX1_346 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_46_DFFSR_113 INVX1_23/gnd DFFSR_186/S FILL
XFILL_5_NAND3X1_107 BUFX2_43/A DFFSR_97/S FILL
XNAND2X1_245 NOR2X1_34/Y NOR2X1_35/Y DFFSR_71/gnd NAND2X1_245/Y DFFSR_10/S NAND2X1
XFILL_36_DFFSR_116 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_9_DFFSR_189 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_4_OAI21X1_191 BUFX2_37/A DFFSR_8/S FILL
XFILL_26_DFFSR_119 BUFX2_37/A DFFSR_81/S FILL
XFILL_18_DFFSR_1 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_2_INVX1_166 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_16_DFFSR_122 INVX1_94/gnd DFFSR_52/S FILL
XFILL_48_DFFSR_34 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_37_DFFSR_74 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_6_AOI21X1_1 INVX1_8/gnd DFFSR_5/S FILL
XFILL_37_1_0 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_4_DFFSR_31 BUFX2_35/A DFFSR_97/S FILL
XFILL_21_DFFSR_24 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_10_DFFSR_64 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_5_OAI21X1_125 BUFX2_35/A DFFSR_14/S FILL
XFILL_2_BUFX2_2 BUFX2_43/A DFFSR_23/S FILL
XFILL_35_3_1 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_0_INVX1_383 INVX1_89/gnd DFFSR_2/S FILL
XFILL_9_OAI22X1_9 INVX1_8/gnd DFFSR_5/S FILL
XFILL_2_DFFSR_119 BUFX2_37/A DFFSR_81/S FILL
XFILL_21_5 INVX1_94/gnd DFFSR_52/S FILL
XFILL_45_DFFSR_81 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_43_DFFSR_150 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_5_NAND2X1_239 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_33_5_2 INVX1_8/gnd DFFSR_7/S FILL
XFILL_33_DFFSR_153 BUFX2_36/A DFFSR_8/S FILL
XFILL_23_DFFSR_156 INVX1_23/gnd DFFSR_91/S FILL
XFILL_1_INVX1_25 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_1_DFFSR_78 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_29_DFFSR_31 BUFX2_35/A DFFSR_97/S FILL
XFILL_13_DFFSR_159 BUFX2_36/A DFFSR_6/S FILL
XFILL_18_DFFSR_71 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_3_OAI21X1_221 BUFX2_35/A DFFSR_14/S FILL
XFILL_6_NAND2X1_173 BUFX2_35/A DFFSR_14/S FILL
XFILL_3_INVX1_310 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_9_DFFPOSX1_11 INVX1_4/gnd DFFSR_4/S FILL
XFILL_22_DFFPOSX1_3 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_0_BUFX2_16 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_5_XOR2X1_8 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_9_DFFSR_153 BUFX2_36/A DFFSR_8/S FILL
XFILL_21_DFFPOSX1_6 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_18_DFFPOSX1_30 BUFX2_43/A DFFSR_97/S FILL
XFILL_20_DFFPOSX1_9 BUFX2_37/A DFFSR_8/S FILL
XFILL_4_OAI21X1_155 BUFX2_7/gnd DFFSR_81/S FILL
XNAND2X1_209 INVX1_243/Y NAND2X1_208/Y DFFSR_71/gnd NAND3X1_60/B DFFSR_10/S NAND2X1
XFILL_50_DFFSR_184 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_2_INVX1_130 BUFX2_36/A DFFSR_6/S FILL
XFILL_40_DFFSR_187 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_9_DFFSR_85 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_37_DFFSR_38 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_26_DFFSR_78 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_30_DFFSR_190 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_10_DFFSR_28 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_4_NAND2X1_269 INVX1_4/gnd DFFSR_4/S FILL
XFILL_43_0_2 INVX1_4/gnd DFFSR_51/S FILL
XFILL_18_NOR3X1_2 INVX1_89/gnd DFFSR_2/S FILL
XFILL_0_INVX1_347 INVX1_4/gnd DFFSR_4/S FILL
XFILL_2_OAI21X1_251 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_43_DFFSR_114 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_33_DFFSR_117 INVX1_23/gnd DFFSR_91/S FILL
XFILL_5_NAND2X1_203 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_34_DFFSR_85 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_45_DFFSR_45 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_6_DFFSR_190 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_23_DFFSR_120 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_4_NAND3X1_101 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_13_DFFSR_123 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_18_DFFSR_35 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_1_DFFSR_42 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_3_OAI21X1_185 BUFX2_36/A DFFSR_8/S FILL
XFILL_6_NAND2X1_137 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_3_AOI21X1_2 INVX1_94/gnd DFFSR_52/S FILL
XFILL_3_INVX1_274 INVX1_8/gnd DFFSR_5/S FILL
XFILL_11_XOR2X1_5 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_42_DFFSR_92 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_9_DFFSR_117 INVX1_23/gnd DFFSR_91/S FILL
XNAND2X1_173 DFFSR_12/S BUFX2_35/A BUFX2_35/A OAI21X1_173/C DFFSR_14/S NAND2X1
XFILL_50_DFFSR_148 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_4_OAI21X1_119 BUFX2_37/A DFFSR_8/S FILL
XFILL_3_AND2X2_1 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_40_DFFSR_151 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_15_DFFSR_82 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_26_DFFSR_42 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_9_DFFSR_49 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_30_DFFSR_154 BUFX2_36/A DFFSR_6/S FILL
XFILL_43_5 INVX1_4/gnd DFFSR_4/S FILL
XFILL_20_DFFSR_157 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_4_NAND2X1_233 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_5_NAND3X1_1 INVX1_94/gnd DFFSR_25/S FILL
XFILL_10_DFFSR_160 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_50_DFFSR_99 BUFX2_35/A DFFSR_97/S FILL
XFILL_3_NAND3X1_131 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_0_INVX1_311 INVX1_94/gnd DFFSR_52/S FILL
XFILL_5_NOR2X1_36 BUFX2_8/gnd DFFSR_10/S FILL
XINVX1_421 BUFX2_32/A DFFSR_1/gnd INVX1_421/Y DFFSR_9/S INVX1
XFILL_30_DFFSR_4 INVX1_4/gnd DFFSR_4/S FILL
XFILL_23_DFFSR_89 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_2_OAI21X1_215 BUFX2_43/A DFFSR_97/S FILL
XFILL_6_DFFSR_154 BUFX2_36/A DFFSR_6/S FILL
XFILL_6_DFFSR_96 INVX1_2/gnd DFFSR_1/S FILL
XFILL_5_NAND2X1_167 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_4_INVX1_418 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_34_DFFSR_49 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_47_DFFSR_185 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_37_DFFSR_188 INVX1_2/gnd DFFSR_1/S FILL
XFILL_27_DFFSR_191 INVX1_23/gnd DFFSR_91/S FILL
XFILL_17_DFFPOSX1_24 BUFX2_43/A DFFSR_23/S FILL
XFILL_5_BUFX2_34 BUFX2_37/A DFFSR_81/S FILL
XFILL_10_DFFPOSX1_3 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_3_OAI21X1_149 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_3_INVX1_238 BUFX2_37/A DFFSR_81/S FILL
XFILL_6_NAND2X1_101 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_9_DFFPOSX1_6 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_8_DFFPOSX1_9 BUFX2_37/A DFFSR_8/S FILL
XFILL_31_DFFSR_96 INVX1_2/gnd DFFSR_1/S FILL
XFILL_42_DFFSR_56 INVX1_2/gnd DFFSR_51/S FILL
XFILL_3_INVX1_90 DFFSR_73/gnd DFFSR_11/S FILL
XNAND2X1_137 NAND2X1_242/Y DFFSR_25/S BUFX2_19/gnd NAND2X1_137/Y DFFSR_52/S NAND2X1
XFILL_3_NAND2X1_263 INVX1_2/gnd DFFSR_51/S FILL
XFILL_50_DFFSR_112 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_27_DFFPOSX1_13 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_40_DFFSR_115 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_8_AOI21X1_29 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_3_DFFSR_191 INVX1_23/gnd DFFSR_91/S FILL
XFILL_7_AOI21X1_32 BUFX2_43/A DFFSR_23/S FILL
XFILL_15_DFFSR_46 BUFX2_36/A DFFSR_6/S FILL
XFILL_9_DFFSR_13 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_30_DFFSR_118 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_20_DFFSR_121 BUFX2_36/A DFFSR_6/S FILL
XFILL_6_AOI21X1_35 INVX1_94/gnd DFFSR_25/S FILL
XFILL_1_OAI21X1_245 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_5_AOI21X1_38 BUFX2_36/A DFFSR_8/S FILL
XAOI21X1_35 AOI21X1_35/A NAND3X1_88/Y AOI21X1_35/C INVX1_94/gnd AND2X2_13/A DFFSR_25/S
+ AOI21X1
XFILL_4_NAND2X1_197 INVX1_8/gnd DFFSR_5/S FILL
XFILL_4_AOI21X1_41 BUFX2_35/A DFFSR_14/S FILL
XFILL_50_DFFSR_63 INVX1_94/gnd DFFSR_52/S FILL
XFILL_0_AOI21X1_3 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_10_DFFSR_124 INVX1_89/gnd DFFSR_36/S FILL
XINVX1_385 DFFSR_95/Q BUFX2_8/gnd INVX1_385/Y DFFSR_10/S INVX1
XFILL_3_AOI21X1_44 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_0_INVX1_275 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_2_AOI21X1_47 BUFX2_43/A DFFSR_23/S FILL
XFILL_4_INVX1_382 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_2_OAI21X1_179 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_6_DFFSR_60 BUFX2_37/A DFFSR_8/S FILL
XFILL_23_DFFSR_53 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_5_NAND2X1_131 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_12_DFFSR_93 INVX1_2/gnd DFFSR_51/S FILL
XFILL_34_DFFSR_13 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_6_DFFSR_118 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_47_DFFSR_149 INVX1_23/gnd DFFSR_91/S FILL
XFILL_44_1_0 INVX1_2/gnd DFFSR_51/S FILL
XFILL_37_DFFSR_152 BUFX2_5/gnd DFFSR_23/S FILL
XBUFX2_38 BUFX2_37/A BUFX2_37/A BUFX2_38/Y DFFSR_81/S BUFX2
XFILL_3_OAI21X1_113 INVX1_23/gnd DFFSR_91/S FILL
XFILL_27_DFFSR_155 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_17_DFFSR_158 BUFX2_43/A DFFSR_23/S FILL
XFILL_3_INVX1_202 BUFX2_37/A DFFSR_81/S FILL
XFILL_8_OAI21X1_77 INVX1_89/gnd DFFSR_36/S FILL
XFILL_42_3_1 INVX1_4/gnd DFFSR_4/S FILL
XFILL_2_NAND3X1_2 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_6_NAND2X1_98 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_7_OAI21X1_80 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_42_DFFSR_20 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_31_DFFSR_60 BUFX2_37/A DFFSR_8/S FILL
XFILL_6_OAI21X1_83 INVX1_94/gnd DFFSR_52/S FILL
XFILL_2_NOR2X1_37 INVX1_94/gnd DFFSR_25/S FILL
XNAND2X1_101 BUFX2_16/Y DFFSR_93/Q BUFX2_17/gnd NAND2X1_101/Y DFFSR_7/S NAND2X1
XFILL_3_INVX1_54 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_40_5_2 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_3_NAND2X1_227 BUFX2_6/gnd DFFSR_91/S FILL
XNAND2X1_98 BUFX2_18/Y DFFSR_90/Q DFFSR_1/gnd NAND2X1_98/Y DFFSR_9/S NAND2X1
XOAI21X1_83 BUFX2_19/Y INVX1_94/Y OAI21X1_83/C INVX1_94/gnd DFFSR_83/D DFFSR_52/S
+ OAI21X1
XFILL_15_DFFSR_10 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_2_NAND3X1_125 INVX1_8/gnd DFFSR_5/S FILL
XFILL_1_INVX1_419 INVX1_2/gnd DFFSR_51/S FILL
XFILL_5_OAI21X1_86 INVX1_4/gnd DFFSR_51/S FILL
XFILL_44_DFFSR_186 INVX1_23/gnd DFFSR_186/S FILL
XFILL_4_OAI21X1_89 BUFX2_35/A DFFSR_14/S FILL
XFILL_3_DFFSR_155 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_4_NAND2X1_161 INVX1_23/gnd DFFSR_186/S FILL
XFILL_3_OAI21X1_92 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_1_OAI21X1_209 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_34_DFFSR_189 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_2_OAI21X1_95 INVX1_89/gnd DFFSR_36/S FILL
XFILL_0_INVX1_239 BUFX2_35/A DFFSR_97/S FILL
XINVX1_349 INVX1_85/A INVX1_89/gnd INVX1_349/Y DFFSR_2/S INVX1
XFILL_50_DFFSR_27 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_1_OAI21X1_98 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_39_DFFSR_67 INVX1_2/gnd DFFSR_51/S FILL
XFILL_3_1 INVX1_23/gnd DFFSR_186/S FILL
XFILL_16_DFFPOSX1_18 BUFX2_37/A DFFSR_8/S FILL
XFILL_2_AOI21X1_11 INVX1_8/gnd DFFSR_5/S FILL
XFILL_2_OAI21X1_143 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_23_DFFSR_17 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_12_DFFSR_57 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_4_INVX1_346 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_6_DFFSR_24 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_47_DFFSR_113 INVX1_23/gnd DFFSR_186/S FILL
XFILL_1_AOI21X1_14 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_37_DFFSR_116 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_0_AOI21X1_17 INVX1_8/gnd DFFSR_5/S FILL
XFILL_27_DFFSR_119 BUFX2_37/A DFFSR_81/S FILL
XFILL_5_NOR2X1_5 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_2_NAND2X1_257 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_3_INVX1_166 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_9_OAI21X1_38 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_42_DFFSR_7 INVX1_8/gnd DFFSR_7/S FILL
XFILL_47_DFFSR_74 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_17_DFFSR_122 INVX1_94/gnd DFFSR_52/S FILL
XFILL_7_AOI21X1_1 INVX1_8/gnd DFFSR_5/S FILL
XFILL_8_OAI21X1_41 INVX1_8/gnd DFFSR_7/S FILL
XFILL_6_NAND2X1_62 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_3_DFFSR_71 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_7_OAI21X1_44 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_3_INVX1_18 INVX1_89/gnd DFFSR_2/S FILL
XFILL_31_DFFSR_24 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_3_NAND2X1_191 BUFX2_37/A DFFSR_8/S FILL
XFILL_6_OAI21X1_47 INVX1_89/gnd DFFSR_2/S FILL
XFILL_6_DFFPOSX1_29 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_0_OAI21X1_239 INVX1_4/gnd DFFSR_4/S FILL
XFILL_5_NAND2X1_65 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_20_DFFSR_64 BUFX2_16/gnd DFFSR_11/S FILL
XNAND2X1_62 DFFSR_52/S DFFSR_54/Q BUFX2_19/gnd NAND2X1_62/Y DFFSR_54/S NAND2X1
XFILL_4_NAND2X1_68 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_25_2 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_1_INVX1_383 INVX1_89/gnd DFFSR_2/S FILL
XFILL_5_OAI21X1_50 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_3_DFFSR_119 BUFX2_37/A DFFSR_81/S FILL
XFILL_3_NAND2X1_71 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_4_OAI21X1_53 DFFSR_71/gnd DFFSR_45/S FILL
XOAI21X1_47 DFFSR_2/S INVX1_53/Y NAND2X1_47/Y INVX1_89/gnd DFFSR_47/D DFFSR_2/S OAI21X1
XFILL_1_OAI21X1_173 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_44_DFFSR_150 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_7_XOR2X1_1 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_2_NAND2X1_74 INVX1_2/gnd DFFSR_1/S FILL
XFILL_3_OAI21X1_56 INVX1_2/gnd DFFSR_51/S FILL
XFILL_4_NAND2X1_125 BUFX2_35/A DFFSR_14/S FILL
XFILL_34_DFFSR_153 BUFX2_36/A DFFSR_8/S FILL
XFILL_1_NAND2X1_77 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_2_OAI21X1_59 INVX1_4/gnd DFFSR_51/S FILL
XFILL_24_DFFSR_156 INVX1_23/gnd DFFSR_91/S FILL
XFILL_1_OAI21X1_62 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_0_NAND2X1_80 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_39_DFFSR_31 BUFX2_35/A DFFSR_97/S FILL
XFILL_14_DFFSR_159 BUFX2_36/A DFFSR_6/S FILL
XFILL_0_INVX1_203 BUFX2_36/A DFFSR_6/S FILL
XFILL_16_1_1 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_28_DFFSR_71 DFFSR_71/gnd DFFSR_10/S FILL
XINVX1_313 INVX1_8/A INVX1_8/gnd INVX1_313/Y DFFSR_5/S INVX1
XFILL_0_OAI21X1_65 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_0_INVX1_65 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_2_OAI21X1_107 BUFX2_36/A DFFSR_6/S FILL
XFILL_4_INVX1_310 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_12_DFFSR_21 INVX1_2/gnd DFFSR_1/S FILL
XFILL_14_3_2 BUFX2_37/A DFFSR_8/S FILL
XNOR2X1_9 NOR2X1_9/A NOR2X1_9/B BUFX2_43/A NOR2X1_9/Y DFFSR_97/S NOR2X1
XFILL_3_NOR3X1_2 INVX1_89/gnd DFFSR_2/S FILL
XDFFSR_1 INVX1_2/A DFFSR_1/CLK DFFSR_6/R DFFSR_1/S DFFSR_1/D DFFSR_1/gnd DFFSR_1/S
+ DFFSR
XFILL_0_DFFSR_156 INVX1_23/gnd DFFSR_91/S FILL
XFILL_2_NAND2X1_221 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_3_INVX1_130 BUFX2_36/A DFFSR_6/S FILL
XFILL_41_DFFSR_187 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_47_DFFSR_38 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_36_DFFSR_78 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_31_DFFSR_190 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_1_NAND3X1_119 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_6_NAND2X1_26 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_0_OAI21X1_203 BUFX2_35/A DFFSR_14/S FILL
XFILL_20_DFFSR_28 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_3_DFFSR_35 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_5_NAND2X1_29 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_6_OAI21X1_11 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_3_NAND2X1_155 BUFX2_37/A DFFSR_81/S FILL
XNAND2X1_26 DFFSR_9/S INVX1_21/A DFFSR_1/gnd OAI21X1_26/C DFFSR_9/S NAND2X1
XFILL_5_OAI21X1_14 BUFX2_43/A DFFSR_23/S FILL
XFILL_1_INVX1_347 INVX1_4/gnd DFFSR_4/S FILL
XFILL_4_NAND2X1_32 DFFSR_3/gnd DFFSR_65/S FILL
XOAI21X1_11 DFFSR_49/S INVX1_13/Y OAI21X1_11/C BUFX2_16/gnd DFFSR_11/D DFFSR_11/S
+ OAI21X1
XFILL_44_DFFSR_114 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_4_OAI21X1_17 INVX1_8/gnd DFFSR_5/S FILL
XFILL_3_NAND2X1_35 BUFX2_17/gnd DFFSR_7/S FILL
XDFFPOSX1_29 NOR2X1_1/B CLKBUF1_13/Y NOR2X1_54/Y DFFSR_1/gnd DFFSR_9/S DFFPOSX1
XFILL_3_OAI21X1_20 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_34_DFFSR_117 INVX1_23/gnd DFFSR_91/S FILL
XFILL_9_NAND3X1_94 BUFX2_35/A DFFSR_97/S FILL
XFILL_1_OAI21X1_137 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_44_DFFSR_85 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_2_NAND2X1_38 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_15_DFFPOSX1_12 INVX1_8/gnd DFFSR_5/S FILL
XFILL_29_DFFSR_1 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_7_DFFSR_190 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_2_OAI21X1_23 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_1_NAND2X1_41 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_24_DFFSR_120 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_0_INVX1_167 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_8_NAND3X1_97 BUFX2_35/A DFFSR_97/S FILL
XAOI21X1_5 AOI21X1_5/A AOI21X1_5/B AOI21X1_5/C BUFX2_37/A AOI21X1_5/Y DFFSR_81/S AOI21X1
XFILL_0_INVX1_29 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_0_NAND2X1_44 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_28_DFFSR_35 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_1_OAI21X1_26 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_0_DFFSR_82 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_17_DFFSR_75 INVX1_4/gnd DFFSR_51/S FILL
XINVX1_277 INVX1_57/A DFFSR_3/gnd INVX1_277/Y DFFSR_4/S INVX1
XFILL_14_DFFSR_123 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_1_NAND2X1_251 BUFX2_35/A DFFSR_97/S FILL
XFILL_4_AOI21X1_2 INVX1_94/gnd DFFSR_52/S FILL
XFILL_0_OAI21X1_29 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_4_INVX1_274 INVX1_8/gnd DFFSR_5/S FILL
XFILL_5_DFFPOSX1_23 INVX1_23/gnd DFFSR_91/S FILL
XFILL_2_NAND2X1_185 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_0_DFFSR_120 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_8_DFFSR_89 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_41_DFFSR_151 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_47_2 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_25_DFFSR_82 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_36_DFFSR_42 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_31_DFFSR_154 BUFX2_36/A DFFSR_6/S FILL
XFILL_4_AOI22X1_10 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_21_DFFSR_157 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_3_AOI22X1_13 INVX1_23/gnd DFFSR_186/S FILL
XFILL_3_NAND2X1_119 BUFX2_37/A DFFSR_8/S FILL
XFILL_6_NAND3X1_1 INVX1_94/gnd DFFSR_25/S FILL
XFILL_0_OAI21X1_167 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_11_DFFSR_160 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_1_INVX1_311 INVX1_94/gnd DFFSR_52/S FILL
XFILL_6_NOR2X1_36 BUFX2_8/gnd DFFSR_10/S FILL
XINVX1_3 DFFSR_2/Q INVX1_8/gnd INVX1_3/Y DFFSR_5/S INVX1
XFILL_11_OAI22X1_37 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_33_DFFSR_89 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_10_OAI22X1_40 BUFX2_37/A DFFSR_8/S FILL
XFILL_0_NAND2X1_281 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_1_OAI21X1_101 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_44_DFFSR_49 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_48_DFFSR_185 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_7_DFFSR_154 BUFX2_36/A DFFSR_6/S FILL
XFILL_24_DFFPOSX1_31 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_9_OAI22X1_43 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_8_NAND3X1_61 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_38_DFFSR_188 INVX1_2/gnd DFFSR_1/S FILL
XFILL_28_DFFSR_191 INVX1_23/gnd DFFSR_91/S FILL
XFILL_7_NAND3X1_64 BUFX2_35/A DFFSR_14/S FILL
XINVX1_241 INVX1_241/A BUFX2_43/A INVX1_241/Y DFFSR_23/S INVX1
XFILL_0_DFFSR_46 BUFX2_36/A DFFSR_6/S FILL
XFILL_8_OAI22X1_46 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_17_DFFSR_39 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_0_INVX1_131 INVX1_89/gnd DFFSR_36/S FILL
XFILL_47_5_2 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_6_NAND3X1_67 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_1_NAND2X1_215 BUFX2_43/A DFFSR_23/S FILL
XFILL_7_OAI22X1_49 INVX1_94/gnd DFFSR_25/S FILL
XFILL_5_NAND3X1_70 BUFX2_35/A DFFSR_14/S FILL
XFILL_6_OAI22X1_52 INVX1_94/gnd DFFSR_25/S FILL
XNAND3X1_67 NAND3X1_66/Y NAND3X1_67/B NAND3X1_67/C BUFX2_6/gnd AOI22X1_10/D DFFSR_14/S
+ NAND3X1
XFILL_4_NAND3X1_73 BUFX2_43/A DFFSR_23/S FILL
XFILL_10_XOR2X1_9 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_0_NAND3X1_113 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_5_OAI22X1_55 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_3_NAND3X1_76 BUFX2_5/gnd DFFSR_6/S FILL
XOAI22X1_52 INVX1_362/Y OAI22X1_40/B INVX1_363/Y OAI22X1_52/D INVX1_94/gnd NOR2X1_35/B
+ DFFSR_25/S OAI22X1
XFILL_4_OAI22X1_58 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_41_DFFSR_96 INVX1_2/gnd DFFSR_1/S FILL
XFILL_2_NAND2X1_149 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_41_DFFSR_115 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_2_NAND3X1_79 BUFX2_36/A DFFSR_6/S FILL
XFILL_2_AND2X2_5 BUFX2_37/A DFFSR_81/S FILL
XFILL_3_OAI22X1_61 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_8_OAI21X1_252 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_4_DFFSR_191 INVX1_23/gnd DFFSR_91/S FILL
XFILL_25_DFFSR_46 BUFX2_36/A DFFSR_6/S FILL
XFILL_15_4_0 BUFX2_37/A DFFSR_81/S FILL
XFILL_8_DFFSR_53 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_14_DFFSR_86 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_31_DFFSR_118 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_1_NAND3X1_82 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_2_OAI22X1_64 INVX1_94/gnd DFFSR_25/S FILL
XFILL_21_DFFSR_121 BUFX2_36/A DFFSR_6/S FILL
XFILL_0_NAND3X1_85 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_0_OAI21X1_131 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_1_OAI22X1_67 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_1_AOI21X1_3 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_11_DFFSR_124 INVX1_89/gnd DFFSR_36/S FILL
XFILL_20_DFFSR_8 BUFX2_36/A DFFSR_8/S FILL
XFILL_1_INVX1_275 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_33_DFFSR_53 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_0_NAND2X1_245 DFFSR_71/gnd DFFSR_10/S FILL
XINVX1_87 INVX1_87/A INVX1_89/gnd INVX1_87/Y DFFSR_36/S INVX1
XFILL_22_DFFSR_93 INVX1_2/gnd DFFSR_51/S FILL
XFILL_44_DFFSR_13 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_7_DFFSR_118 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_48_DFFSR_149 INVX1_23/gnd DFFSR_91/S FILL
XFILL_38_DFFSR_152 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_4_BUFX2_9 BUFX2_37/A DFFSR_8/S FILL
XFILL_8_NAND3X1_25 BUFX2_7/gnd DFFSR_81/S FILL
XINVX1_205 INVX1_256/A INVX1_94/gnd INVX1_205/Y DFFSR_25/S INVX1
XFILL_0_DFFSR_10 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_4_DFFPOSX1_17 BUFX2_37/A DFFSR_8/S FILL
XFILL_4_BUFX2_38 BUFX2_37/A DFFSR_81/S FILL
XFILL_7_NAND3X1_28 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_28_DFFSR_155 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_1_NAND2X1_179 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_8_OAI22X1_10 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_18_DFFSR_158 BUFX2_43/A DFFSR_23/S FILL
XFILL_4_INVX1_202 BUFX2_37/A DFFSR_81/S FILL
XFILL_6_NAND3X1_31 INVX1_94/gnd DFFSR_52/S FILL
XFILL_7_OAI22X1_13 DFFSR_3/gnd DFFSR_65/S FILL
XNAND3X1_31 NAND3X1_56/A NAND3X1_30/Y INVX1_230/Y INVX1_94/gnd NAND3X1_58/A DFFSR_52/S
+ NAND3X1
XFILL_3_NAND3X1_2 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_5_NAND3X1_34 INVX1_2/gnd DFFSR_1/S FILL
XFILL_6_OAI22X1_16 INVX1_4/gnd DFFSR_4/S FILL
XFILL_41_DFFSR_4 INVX1_4/gnd DFFSR_4/S FILL
XFILL_4_NAND3X1_37 BUFX2_43/A DFFSR_97/S FILL
XFILL_41_DFFSR_60 BUFX2_37/A DFFSR_8/S FILL
XFILL_2_INVX1_94 INVX1_94/gnd DFFSR_52/S FILL
XFILL_3_NOR2X1_37 INVX1_94/gnd DFFSR_25/S FILL
XFILL_5_OAI22X1_19 DFFSR_71/gnd DFFSR_45/S FILL
XOAI22X1_16 INVX1_287/Y OAI22X1_8/B INVX1_288/Y OAI22X1_8/D INVX1_4/gnd NOR2X1_17/A
+ DFFSR_4/S OAI22X1
XFILL_2_NAND2X1_113 INVX1_23/gnd DFFSR_91/S FILL
XFILL_8_OAI21X1_216 BUFX2_35/A DFFSR_14/S FILL
XFILL_3_NAND3X1_40 BUFX2_43/A DFFSR_23/S FILL
XDFFSR_158 INVX1_190/A CLKBUF1_14/Y DFFSR_158/R DFFSR_158/S DFFSR_158/D BUFX2_43/A
+ DFFSR_23/S DFFSR
XFILL_4_OAI22X1_22 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_2_NAND3X1_43 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_3_OAI22X1_25 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_25_DFFSR_10 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_8_DFFSR_17 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_2_INVX1_419 INVX1_2/gnd DFFSR_51/S FILL
XFILL_14_DFFSR_50 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_45_DFFSR_186 INVX1_23/gnd DFFSR_186/S FILL
XFILL_1_NAND3X1_46 BUFX2_35/A DFFSR_97/S FILL
XFILL_4_DFFSR_155 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_2_OAI22X1_28 INVX1_94/gnd DFFSR_25/S FILL
XFILL_0_NAND3X1_49 BUFX2_37/A DFFSR_8/S FILL
XFILL_23_1_1 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_1_OAI22X1_31 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_35_DFFSR_189 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_5_0_0 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_23_DFFPOSX1_25 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_0_OAI22X1_34 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_1_INVX1_239 BUFX2_35/A DFFSR_97/S FILL
XFILL_21_3_2 INVX1_94/gnd DFFSR_25/S FILL
XFILL_49_DFFSR_67 INVX1_2/gnd DFFSR_51/S FILL
XFILL_3_2_1 INVX1_23/gnd DFFSR_91/S FILL
XFILL_0_NAND2X1_209 DFFSR_71/gnd DFFSR_10/S FILL
XINVX1_51 DFFSR_45/Q DFFSR_79/gnd INVX1_51/Y DFFSR_36/S INVX1
XFILL_33_DFFSR_17 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_22_DFFSR_57 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_5_DFFSR_64 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_1_4_2 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_48_DFFSR_113 INVX1_23/gnd DFFSR_186/S FILL
XFILL_11_DFFSR_97 BUFX2_35/A DFFSR_97/S FILL
XFILL_38_DFFSR_116 DFFSR_5/gnd DFFSR_2/S FILL
XINVX1_169 BUFX2_6/Y DFFSR_89/gnd DFFSR_147/R DFFSR_186/S INVX1
XFILL_28_DFFSR_119 BUFX2_37/A DFFSR_81/S FILL
XFILL_4_INVX1_166 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_1_NAND2X1_143 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_7_OAI21X1_246 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_18_DFFSR_122 INVX1_94/gnd DFFSR_52/S FILL
XFILL_8_AOI21X1_1 INVX1_8/gnd DFFSR_5/S FILL
XFILL_41_DFFSR_24 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_2_INVX1_58 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_30_DFFSR_64 BUFX2_16/gnd DFFSR_11/S FILL
XDFFSR_122 DFFSR_122/Q CLKBUF1_1/Y DFFSR_123/R DFFSR_52/S DFFSR_122/D INVX1_94/gnd
+ DFFSR_52/S DFFSR
XFILL_8_OAI21X1_180 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_2_INVX1_383 INVX1_89/gnd DFFSR_2/S FILL
XFILL_14_DFFSR_14 BUFX2_35/A DFFSR_14/S FILL
XFILL_4_DFFSR_119 BUFX2_37/A DFFSR_81/S FILL
XFILL_1_NAND3X1_10 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_45_DFFSR_150 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_35_DFFSR_153 BUFX2_36/A DFFSR_8/S FILL
XFILL_0_NAND3X1_13 INVX1_94/gnd DFFSR_25/S FILL
XFILL_8_DFFSR_7 INVX1_8/gnd DFFSR_7/S FILL
XFILL_25_DFFSR_156 INVX1_23/gnd DFFSR_91/S FILL
XFILL_49_DFFSR_31 BUFX2_35/A DFFSR_97/S FILL
XFILL_15_DFFSR_159 BUFX2_36/A DFFSR_6/S FILL
XFILL_1_INVX1_203 BUFX2_36/A DFFSR_6/S FILL
XFILL_38_DFFSR_71 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_0_NAND3X1_3 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_3_DFFPOSX1_11 INVX1_4/gnd DFFSR_4/S FILL
XFILL_0_NAND2X1_173 BUFX2_35/A DFFSR_14/S FILL
XDFFSR_68 DFFSR_68/Q INVX1_172/A DFFSR_68/R DFFSR_14/S DFFSR_68/D BUFX2_35/A DFFSR_14/S
+ DFFSR
XFILL_11_DFFSR_61 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_5_DFFSR_28 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_0_NOR2X1_38 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_22_DFFSR_21 INVX1_2/gnd DFFSR_1/S FILL
XINVX1_15 DFFSR_13/Q DFFSR_3/gnd INVX1_15/Y DFFSR_65/S INVX1
XFILL_4_NOR2X1_9 BUFX2_43/A DFFSR_97/S FILL
XFILL_8_NAND3X1_126 DFFSR_5/gnd DFFSR_5/S FILL
XINVX1_133 INVX1_374/A DFFSR_73/gnd INVX1_133/Y DFFSR_11/S INVX1
XFILL_1_DFFSR_156 INVX1_23/gnd DFFSR_91/S FILL
XFILL_12_DFFPOSX1_30 BUFX2_43/A DFFSR_97/S FILL
XFILL_1_NAND2X1_107 BUFX2_36/A DFFSR_6/S FILL
XFILL_42_DFFSR_187 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_4_INVX1_130 BUFX2_36/A DFFSR_6/S FILL
XFILL_7_OAI21X1_210 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_46_DFFSR_78 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_32_DFFSR_190 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_19_DFFSR_68 BUFX2_35/A DFFSR_14/S FILL
XFILL_30_DFFSR_28 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_2_INVX1_22 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_2_DFFSR_75 INVX1_4/gnd DFFSR_51/S FILL
XFILL_8_OAI21X1_144 INVX1_8/gnd DFFSR_7/S FILL
XFILL_22_DFFPOSX1_19 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_2_INVX1_347 INVX1_4/gnd DFFSR_4/S FILL
XFILL_6_XOR2X1_5 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_1_BUFX2_13 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_45_DFFSR_114 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_35_DFFSR_117 INVX1_23/gnd DFFSR_91/S FILL
XFILL_8_DFFSR_190 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_1_INVX1_167 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_38_DFFSR_35 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_27_DFFSR_75 INVX1_4/gnd DFFSR_51/S FILL
XFILL_25_DFFSR_120 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_15_DFFSR_123 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_5_AOI21X1_2 INVX1_94/gnd DFFSR_52/S FILL
XFILL_0_NAND2X1_137 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_6_OAI21X1_240 DFFSR_5/gnd DFFSR_5/S FILL
XDFFSR_32 INVX1_36/A DFFSR_24/CLK DFFSR_31/R DFFSR_1/S DFFSR_32/D INVX1_2/gnd DFFSR_1/S
+ DFFSR
XFILL_11_DFFSR_25 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_22_4_0 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_1_DFFSR_120 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_7_OAI21X1_174 BUFX2_43/A DFFSR_23/S FILL
XFILL_42_DFFSR_151 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_34_4 INVX1_8/gnd DFFSR_7/S FILL
XFILL_35_DFFSR_82 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_46_DFFSR_42 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_2_5_0 INVX1_23/gnd DFFSR_186/S FILL
XFILL_32_DFFSR_154 BUFX2_36/A DFFSR_6/S FILL
XFILL_22_DFFSR_157 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_2_DFFSR_39 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_7_NAND3X1_1 INVX1_94/gnd DFFSR_25/S FILL
XFILL_12_DFFSR_160 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_19_DFFSR_32 INVX1_2/gnd DFFSR_1/S FILL
XFILL_2_INVX1_311 INVX1_94/gnd DFFSR_52/S FILL
XFILL_8_OAI21X1_108 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_20_CLKBUF1_22 INVX1_94/gnd DFFSR_25/S FILL
XFILL_43_DFFSR_89 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_19_CLKBUF1_25 INVX1_23/gnd DFFSR_186/S FILL
XFILL_12_XOR2X1_2 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_19_DFFSR_5 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_49_DFFSR_185 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_8_DFFSR_154 BUFX2_36/A DFFSR_6/S FILL
XFILL_39_DFFSR_188 INVX1_2/gnd DFFSR_1/S FILL
XFILL_27_DFFSR_39 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_16_DFFSR_79 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_1_INVX1_131 INVX1_89/gnd DFFSR_36/S FILL
XFILL_7_NAND3X1_120 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_29_DFFSR_191 INVX1_23/gnd DFFSR_91/S FILL
XFILL_3_BUFX2_6 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_11_DFFPOSX1_24 BUFX2_43/A DFFSR_23/S FILL
XFILL_6_OAI21X1_204 BUFX2_36/A DFFSR_6/S FILL
XFILL_0_NAND2X1_101 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_30_1_1 DFFSR_5/gnd DFFSR_2/S FILL
XOAI21X1_240 INVX1_397/A INVX1_331/A INVX1_332/A DFFSR_5/gnd NAND3X1_128/B DFFSR_5/S
+ OAI21X1
XFILL_51_DFFSR_96 INVX1_2/gnd DFFSR_1/S FILL
XFILL_40_DFFSR_1 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_21_DFFPOSX1_13 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_42_DFFSR_115 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_5_DFFSR_191 INVX1_23/gnd DFFSR_91/S FILL
XFILL_35_DFFSR_46 BUFX2_36/A DFFSR_6/S FILL
XFILL_28_3_2 INVX1_89/gnd DFFSR_36/S FILL
XFILL_24_DFFSR_86 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_7_DFFSR_93 INVX1_2/gnd DFFSR_51/S FILL
XFILL_32_DFFSR_118 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_7_OAI21X1_138 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_22_DFFSR_121 BUFX2_36/A DFFSR_6/S FILL
XFILL_2_AOI21X1_3 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_12_DFFSR_124 INVX1_89/gnd DFFSR_36/S FILL
XFILL_6_BUFX2_31 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_8_4_2 BUFX2_43/A DFFSR_97/S FILL
XFILL_2_INVX1_275 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_5_OAI21X1_234 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_43_DFFSR_53 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_4_INVX1_87 INVX1_89/gnd DFFSR_36/S FILL
XFILL_32_DFFSR_93 INVX1_2/gnd DFFSR_51/S FILL
XFILL_8_DFFSR_118 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_49_DFFSR_149 INVX1_23/gnd DFFSR_91/S FILL
XFILL_39_DFFSR_152 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_16_DFFSR_43 INVX1_94/gnd DFFSR_25/S FILL
XFILL_29_DFFSR_155 BUFX2_7/gnd DFFSR_54/S FILL
XNAND3X1_5 NOR2X1_4/Y NAND3X1_4/Y NAND3X1_5/C BUFX2_8/gnd INVX1_223/A DFFSR_10/S NAND3X1
XFILL_19_DFFSR_158 BUFX2_43/A DFFSR_23/S FILL
XFILL_6_OAI21X1_168 BUFX2_36/A DFFSR_6/S FILL
XFILL_4_NAND3X1_2 BUFX2_8/gnd DFFSR_10/S FILL
XNOR2X1_40 NOR2X1_40/A NOR2X1_40/B BUFX2_8/gnd NOR2X1_40/Y DFFSR_10/S NOR2X1
XFILL_51_DFFSR_60 BUFX2_37/A DFFSR_8/S FILL
XFILL_4_NOR2X1_37 INVX1_94/gnd DFFSR_25/S FILL
XOAI21X1_204 INVX1_213/Y NOR2X1_10/B NOR2X1_8/A BUFX2_36/A NAND3X1_37/B DFFSR_6/S
+ OAI21X1
XFILL_12_CLKBUF1_10 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_1_AND2X2_9 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_35_DFFSR_10 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_6_NAND2X1_282 INVX1_89/gnd DFFSR_2/S FILL
XFILL_7_OAI21X1_102 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_7_DFFSR_57 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_13_DFFSR_90 INVX1_2/gnd DFFSR_1/S FILL
XFILL_3_INVX1_419 INVX1_2/gnd DFFSR_51/S FILL
XFILL_11_CLKBUF1_13 INVX1_4/gnd DFFSR_51/S FILL
XFILL_24_DFFSR_50 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_46_DFFSR_186 INVX1_23/gnd DFFSR_186/S FILL
XFILL_10_CLKBUF1_16 BUFX2_36/A DFFSR_6/S FILL
XFILL_5_DFFSR_155 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_4_OAI21X1_264 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_36_DFFSR_189 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_2_INVX1_239 BUFX2_35/A DFFSR_97/S FILL
XFILL_9_CLKBUF1_19 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_7_DFFSR_4 INVX1_4/gnd DFFSR_4/S FILL
XFILL_8_CLKBUF1_22 INVX1_94/gnd DFFSR_25/S FILL
XFILL_6_NAND3X1_114 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_7_CLKBUF1_25 INVX1_23/gnd DFFSR_186/S FILL
XFILL_10_DFFPOSX1_18 BUFX2_37/A DFFSR_8/S FILL
XFILL_4_INVX1_51 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_43_DFFSR_17 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_49_DFFSR_113 INVX1_23/gnd DFFSR_186/S FILL
XFILL_21_DFFSR_97 BUFX2_35/A DFFSR_97/S FILL
XFILL_5_OAI21X1_198 INVX1_8/gnd DFFSR_7/S FILL
XFILL_32_DFFSR_57 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_39_DFFSR_116 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_3_BUFX2_42 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_29_DFFSR_119 BUFX2_37/A DFFSR_81/S FILL
XFILL_31_DFFSR_8 BUFX2_36/A DFFSR_8/S FILL
XFILL_19_DFFSR_122 INVX1_94/gnd DFFSR_52/S FILL
XFILL_6_OAI21X1_132 INVX1_4/gnd DFFSR_4/S FILL
XOAI21X1_168 DFFSR_23/S INVX1_203/Y NAND2X1_168/Y BUFX2_36/A DFFSR_168/D DFFSR_6/S
+ OAI21X1
XFILL_16_1 BUFX2_37/A DFFSR_81/S FILL
XFILL_0_DFFPOSX1_29 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_1_INVX1_98 INVX1_4/gnd DFFSR_4/S FILL
XFILL_40_DFFSR_64 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_6_NAND2X1_246 INVX1_94/gnd DFFSR_25/S FILL
XFILL_3_INVX1_383 INVX1_89/gnd DFFSR_2/S FILL
XFILL_24_DFFSR_14 BUFX2_35/A DFFSR_14/S FILL
XFILL_5_DFFSR_119 BUFX2_37/A DFFSR_81/S FILL
XFILL_13_DFFSR_54 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_7_DFFSR_21 INVX1_2/gnd DFFSR_1/S FILL
XFILL_46_DFFSR_150 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_36_DFFSR_153 BUFX2_36/A DFFSR_8/S FILL
XFILL_6_NOR2X1_2 BUFX2_7/gnd DFFSR_81/S FILL
XNAND2X1_282 AND2X2_16/Y XOR2X1_15/B INVX1_89/gnd AOI21X1_46/C DFFSR_2/S NAND2X1
XFILL_26_DFFSR_156 INVX1_23/gnd DFFSR_91/S FILL
XFILL_4_OAI21X1_228 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_16_DFFSR_159 BUFX2_36/A DFFSR_6/S FILL
XFILL_2_INVX1_203 BUFX2_36/A DFFSR_6/S FILL
XFILL_48_DFFSR_71 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_29_4_0 INVX1_89/gnd DFFSR_2/S FILL
XFILL_1_NAND3X1_3 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_5_OAI21X1_162 INVX1_23/gnd DFFSR_91/S FILL
XFILL_4_DFFSR_68 BUFX2_35/A DFFSR_14/S FILL
XFILL_21_DFFSR_61 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_1_NOR2X1_38 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_32_DFFSR_21 INVX1_2/gnd DFFSR_1/S FILL
XFILL_9_5_0 BUFX2_43/A DFFSR_23/S FILL
XNAND3X1_114 NOR2X1_1/A NOR2X1_2/A INVX1_266/Y DFFSR_71/gnd OAI22X1_6/B DFFSR_10/S
+ NAND3X1
XFILL_0_INVX1_420 INVX1_2/gnd DFFSR_51/S FILL
XFILL_2_DFFSR_156 INVX1_23/gnd DFFSR_91/S FILL
XFILL_43_DFFSR_187 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_5_NAND2X1_276 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_33_DFFSR_190 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_29_DFFSR_68 BUFX2_35/A DFFSR_14/S FILL
XFILL_40_DFFSR_28 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_1_INVX1_62 INVX1_89/gnd DFFSR_2/S FILL
XFILL_0_CLKBUF1_10 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_3_OAI21X1_258 INVX1_2/gnd DFFSR_51/S FILL
XOAI21X1_132 DFFSR_51/S INVX1_149/Y NAND2X1_132/Y INVX1_4/gnd DFFSR_132/D DFFSR_4/S
+ OAI21X1
XFILL_6_NAND2X1_210 BUFX2_35/A DFFSR_97/S FILL
XFILL_13_DFFSR_18 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_3_INVX1_347 INVX1_4/gnd DFFSR_4/S FILL
XFILL_5_NAND3X1_108 BUFX2_37/A DFFSR_81/S FILL
XFILL_46_DFFSR_114 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_36_DFFSR_117 INVX1_23/gnd DFFSR_91/S FILL
XNAND2X1_246 NOR2X1_37/Y NOR2X1_36/Y INVX1_94/gnd NAND2X1_246/Y DFFSR_25/S NAND2X1
XFILL_9_DFFSR_190 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_4_OAI21X1_192 BUFX2_37/A DFFSR_81/S FILL
XFILL_18_DFFSR_2 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_2_INVX1_167 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_48_DFFSR_35 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_37_DFFSR_75 INVX1_4/gnd DFFSR_51/S FILL
XFILL_26_DFFSR_120 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_16_DFFSR_123 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_6_AOI21X1_2 INVX1_94/gnd DFFSR_52/S FILL
XFILL_37_1_1 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_4_DFFSR_32 INVX1_2/gnd DFFSR_1/S FILL
XFILL_21_DFFSR_25 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_2_BUFX2_3 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_5_OAI21X1_126 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_35_3_2 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_10_DFFSR_65 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_0_INVX1_384 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_21_6 INVX1_94/gnd DFFSR_52/S FILL
XFILL_2_DFFSR_120 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_38_1 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_43_DFFSR_151 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_5_NAND2X1_240 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_45_DFFSR_82 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_33_DFFSR_154 BUFX2_36/A DFFSR_6/S FILL
XFILL_23_DFFSR_157 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_1_INVX1_26 BUFX2_43/A DFFSR_23/S FILL
XFILL_8_NAND3X1_1 INVX1_94/gnd DFFSR_25/S FILL
XFILL_1_DFFSR_79 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_18_DFFSR_72 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_13_DFFSR_160 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_29_DFFSR_32 INVX1_2/gnd DFFSR_1/S FILL
XFILL_3_OAI21X1_222 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_23_DFFPOSX1_1 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_6_NAND2X1_174 BUFX2_43/A DFFSR_97/S FILL
XFILL_3_INVX1_311 INVX1_94/gnd DFFSR_52/S FILL
XFILL_9_DFFPOSX1_12 INVX1_8/gnd DFFSR_5/S FILL
XFILL_22_DFFPOSX1_4 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_0_BUFX2_17 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_5_XOR2X1_9 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_21_DFFPOSX1_7 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_50_DFFSR_185 DFFSR_89/gnd DFFSR_92/S FILL
XNAND2X1_210 AND2X2_9/A AND2X2_8/B BUFX2_35/A XOR2X1_4/A DFFSR_97/S NAND2X1
XFILL_9_DFFSR_154 BUFX2_36/A DFFSR_6/S FILL
XFILL_18_DFFPOSX1_31 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_4_OAI21X1_156 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_37_DFFSR_39 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_26_DFFSR_79 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_2_INVX1_131 INVX1_89/gnd DFFSR_36/S FILL
XFILL_9_DFFSR_86 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_40_DFFSR_188 INVX1_2/gnd DFFSR_1/S FILL
XFILL_30_DFFSR_191 INVX1_23/gnd DFFSR_91/S FILL
XFILL_4_NAND2X1_270 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_10_DFFSR_29 INVX1_4/gnd DFFSR_4/S FILL
XFILL_0_INVX1_348 INVX1_4/gnd DFFSR_4/S FILL
XFILL_43_DFFSR_115 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_2_OAI21X1_252 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_6_DFFSR_191 INVX1_23/gnd DFFSR_91/S FILL
XFILL_5_NAND2X1_204 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_45_DFFSR_46 BUFX2_36/A DFFSR_6/S FILL
XFILL_34_DFFSR_86 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_33_DFFSR_118 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_4_NAND3X1_102 INVX1_23/gnd DFFSR_186/S FILL
XFILL_23_DFFSR_121 BUFX2_36/A DFFSR_6/S FILL
XFILL_1_DFFSR_43 INVX1_94/gnd DFFSR_25/S FILL
XFILL_18_DFFSR_36 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_3_OAI21X1_186 BUFX2_36/A DFFSR_8/S FILL
XFILL_13_DFFSR_124 INVX1_89/gnd DFFSR_36/S FILL
XFILL_3_AOI21X1_3 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_3_INVX1_275 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_6_NAND2X1_138 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_6_DFFSR_1 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_11_XOR2X1_6 DFFSR_89/gnd DFFSR_186/S FILL
XNAND2X1_174 DFFSR_6/S BUFX2_43/A BUFX2_43/A NAND2X1_174/Y DFFSR_97/S NAND2X1
XFILL_42_DFFSR_93 INVX1_2/gnd DFFSR_51/S FILL
XFILL_9_DFFSR_118 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_50_DFFSR_149 INVX1_23/gnd DFFSR_91/S FILL
XFILL_4_OAI21X1_120 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_40_DFFSR_152 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_3_AND2X2_2 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_15_DFFSR_83 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_26_DFFSR_43 INVX1_94/gnd DFFSR_25/S FILL
XFILL_9_DFFSR_50 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_30_DFFSR_155 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_43_6 INVX1_4/gnd DFFSR_4/S FILL
XFILL_20_DFFSR_158 BUFX2_43/A DFFSR_23/S FILL
XFILL_4_OR2X2_1 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_10_DFFSR_161 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_5_NAND3X1_2 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_4_NAND2X1_234 BUFX2_16/gnd DFFSR_65/S FILL
XINVX1_422 BUFX2_33/A INVX1_23/gnd INVX1_422/Y DFFSR_186/S INVX1
XFILL_0_INVX1_312 BUFX2_36/A DFFSR_6/S FILL
XFILL_5_NOR2X1_37 INVX1_94/gnd DFFSR_25/S FILL
XFILL_3_NAND3X1_132 INVX1_8/gnd DFFSR_7/S FILL
XFILL_30_DFFSR_5 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_2_OAI21X1_216 BUFX2_35/A DFFSR_14/S FILL
XFILL_6_DFFSR_97 BUFX2_35/A DFFSR_97/S FILL
XFILL_5_NAND2X1_168 BUFX2_36/A DFFSR_6/S FILL
XFILL_45_DFFSR_10 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_4_INVX1_419 INVX1_2/gnd DFFSR_51/S FILL
XFILL_34_DFFSR_50 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_47_DFFSR_186 INVX1_23/gnd DFFSR_186/S FILL
XFILL_6_DFFSR_155 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_36_4_0 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_23_DFFSR_90 INVX1_2/gnd DFFSR_1/S FILL
XFILL_11_DFFPOSX1_1 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_5_BUFX2_35 BUFX2_35/A DFFSR_14/S FILL
XFILL_17_DFFPOSX1_25 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_10_DFFPOSX1_4 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_37_DFFSR_189 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_3_INVX1_239 BUFX2_35/A DFFSR_97/S FILL
XFILL_3_OAI21X1_150 INVX1_94/gnd DFFSR_52/S FILL
XFILL_6_NAND2X1_102 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_51_DFFSR_1 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_9_DFFPOSX1_7 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_3_NAND2X1_264 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_50_DFFSR_113 INVX1_23/gnd DFFSR_186/S FILL
XFILL_31_DFFSR_97 BUFX2_35/A DFFSR_97/S FILL
XFILL_9_AOI21X1_27 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_3_INVX1_91 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_42_DFFSR_57 DFFSR_73/gnd DFFSR_57/S FILL
XNAND2X1_138 DFFSR_11/S NAND2X1_243/Y DFFSR_73/gnd NAND2X1_138/Y DFFSR_57/S NAND2X1
XFILL_8_AOI21X1_30 INVX1_23/gnd DFFSR_91/S FILL
XFILL_27_DFFPOSX1_14 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_40_DFFSR_116 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_7_AOI21X1_33 BUFX2_35/A DFFSR_14/S FILL
XFILL_9_DFFSR_14 BUFX2_35/A DFFSR_14/S FILL
XFILL_15_DFFSR_47 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_30_DFFSR_119 BUFX2_37/A DFFSR_81/S FILL
XFILL_6_AOI21X1_36 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_5_AOI21X1_39 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_20_DFFSR_122 INVX1_94/gnd DFFSR_52/S FILL
XFILL_4_NAND2X1_198 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_1_OAI21X1_246 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_4_AOI21X1_42 INVX1_23/gnd DFFSR_91/S FILL
XFILL_10_DFFSR_125 BUFX2_6/gnd DFFSR_91/S FILL
XAOI21X1_36 NAND3X1_81/Y NAND3X1_84/Y INVX1_250/A BUFX2_8/gnd AOI21X1_36/Y DFFSR_25/S
+ AOI21X1
XFILL_0_AOI21X1_4 BUFX2_7/gnd DFFSR_81/S FILL
XINVX1_386 DFFSR_127/Q INVX1_94/gnd INVX1_386/Y DFFSR_52/S INVX1
XFILL_3_AOI21X1_45 INVX1_89/gnd DFFSR_36/S FILL
XFILL_0_INVX1_276 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_50_DFFSR_64 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_2_OAI21X1_180 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_2_AOI21X1_48 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_34_DFFSR_14 BUFX2_35/A DFFSR_14/S FILL
XFILL_6_DFFSR_61 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_6_DFFSR_119 BUFX2_37/A DFFSR_81/S FILL
XFILL_23_DFFSR_54 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_5_NAND2X1_132 INVX1_8/gnd DFFSR_5/S FILL
XFILL_12_DFFSR_94 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_47_DFFSR_150 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_44_1_1 INVX1_2/gnd DFFSR_51/S FILL
XFILL_37_DFFSR_153 BUFX2_36/A DFFSR_8/S FILL
XFILL_27_DFFSR_156 INVX1_23/gnd DFFSR_91/S FILL
XBUFX2_39 BUFX2_35/A BUFX2_43/A BUFX2_39/Y DFFSR_97/S BUFX2
XFILL_3_OAI21X1_114 INVX1_89/gnd DFFSR_36/S FILL
XFILL_17_DFFSR_159 BUFX2_36/A DFFSR_6/S FILL
XFILL_3_INVX1_203 BUFX2_36/A DFFSR_6/S FILL
XFILL_42_3_2 INVX1_4/gnd DFFSR_4/S FILL
XFILL_2_NAND3X1_3 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_8_OAI21X1_78 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_6_NAND2X1_99 BUFX2_43/A DFFSR_97/S FILL
XFILL_31_DFFSR_61 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_3_INVX1_55 BUFX2_36/A DFFSR_8/S FILL
XFILL_7_OAI21X1_81 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_2_NOR2X1_38 BUFX2_17/gnd DFFSR_7/S FILL
XNAND2X1_102 BUFX2_16/Y DFFSR_94/Q BUFX2_17/gnd NAND2X1_102/Y DFFSR_57/S NAND2X1
XFILL_42_DFFSR_21 INVX1_2/gnd DFFSR_1/S FILL
XFILL_3_NAND2X1_228 INVX1_23/gnd DFFSR_91/S FILL
XNAND2X1_99 BUFX2_25/Y DFFSR_91/Q BUFX2_43/A NAND2X1_99/Y DFFSR_97/S NAND2X1
XFILL_6_OAI21X1_84 BUFX2_5/gnd DFFSR_6/S FILL
XOAI21X1_84 BUFX2_20/Y INVX1_95/Y OAI21X1_84/C BUFX2_5/gnd DFFSR_84/D DFFSR_6/S OAI21X1
XFILL_1_INVX1_420 INVX1_2/gnd DFFSR_51/S FILL
XFILL_5_OAI21X1_87 INVX1_4/gnd DFFSR_4/S FILL
XFILL_15_DFFSR_11 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_3_DFFSR_156 INVX1_23/gnd DFFSR_91/S FILL
XFILL_2_NAND3X1_126 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_4_OAI21X1_90 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_10_2_0 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_1_OAI21X1_210 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_3_OAI21X1_93 INVX1_4/gnd DFFSR_51/S FILL
XFILL_44_DFFSR_187 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_4_NAND2X1_162 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_34_DFFSR_190 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_2_OAI21X1_96 INVX1_4/gnd DFFSR_51/S FILL
XFILL_0_INVX1_240 BUFX2_35/A DFFSR_14/S FILL
XFILL_39_DFFSR_68 BUFX2_35/A DFFSR_14/S FILL
XFILL_1_OAI21X1_99 BUFX2_43/A DFFSR_97/S FILL
XINVX1_350 DFFSR_115/Q BUFX2_7/gnd INVX1_350/Y DFFSR_81/S INVX1
XFILL_50_DFFSR_28 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_3_2 INVX1_23/gnd DFFSR_186/S FILL
XFILL_6_DFFSR_25 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_2_AOI21X1_12 INVX1_8/gnd DFFSR_7/S FILL
XFILL_2_OAI21X1_144 INVX1_8/gnd DFFSR_7/S FILL
XFILL_23_DFFSR_18 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_16_DFFPOSX1_19 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_1_AOI21X1_15 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_47_DFFSR_114 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_12_DFFSR_58 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_0_AOI21X1_18 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_37_DFFSR_117 INVX1_23/gnd DFFSR_91/S FILL
XFILL_5_NOR2X1_6 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_2_NAND2X1_258 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_3_INVX1_167 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_42_DFFSR_8 BUFX2_36/A DFFSR_8/S FILL
XFILL_9_OAI21X1_39 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_47_DFFSR_75 INVX1_4/gnd DFFSR_51/S FILL
XFILL_27_DFFSR_120 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_17_DFFSR_123 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_8_OAI21X1_42 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_7_AOI21X1_2 INVX1_94/gnd DFFSR_52/S FILL
XFILL_6_NAND2X1_63 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_7_OAI21X1_45 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_6_DFFPOSX1_30 BUFX2_43/A DFFSR_97/S FILL
XFILL_3_NAND2X1_192 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_31_DFFSR_25 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_0_OAI21X1_240 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_3_DFFSR_72 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_5_NAND2X1_66 INVX1_4/gnd DFFSR_51/S FILL
XFILL_6_OAI21X1_48 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_20_DFFSR_65 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_3_INVX1_19 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_4_NAND2X1_69 BUFX2_19/gnd DFFSR_54/S FILL
XNAND2X1_63 DFFSR_25/S DFFSR_55/Q BUFX2_8/gnd OAI21X1_63/C DFFSR_25/S NAND2X1
XFILL_1_INVX1_384 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_5_OAI21X1_51 INVX1_2/gnd DFFSR_51/S FILL
XFILL_2_BUFX2_10 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_4_OAI21X1_54 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_25_3 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_3_NAND2X1_72 DFFSR_5/gnd DFFSR_2/S FILL
XOAI21X1_48 DFFSR_1/S INVX1_54/Y NAND2X1_48/Y DFFSR_3/gnd DFFSR_48/D DFFSR_4/S OAI21X1
XFILL_3_DFFSR_120 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_44_DFFSR_151 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_7_XOR2X1_2 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_2_NAND2X1_75 INVX1_4/gnd DFFSR_4/S FILL
XFILL_3_OAI21X1_57 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_1_OAI21X1_174 BUFX2_43/A DFFSR_23/S FILL
XFILL_34_DFFSR_154 BUFX2_36/A DFFSR_6/S FILL
XFILL_2_OAI21X1_60 BUFX2_37/A DFFSR_81/S FILL
XFILL_4_NAND2X1_126 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_1_NAND2X1_78 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_24_DFFSR_157 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_1_OAI21X1_63 INVX1_94/gnd DFFSR_25/S FILL
XFILL_0_NAND2X1_81 INVX1_94/gnd DFFSR_25/S FILL
XFILL_0_INVX1_204 BUFX2_36/A DFFSR_8/S FILL
XFILL_16_1_2 BUFX2_7/gnd DFFSR_81/S FILL
XINVX1_314 DFFSR_15/Q INVX1_8/gnd INVX1_314/Y DFFSR_5/S INVX1
XFILL_28_DFFSR_72 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_14_DFFSR_160 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_39_DFFSR_32 INVX1_2/gnd DFFSR_1/S FILL
XFILL_0_INVX1_66 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_4_INVX1_311 INVX1_94/gnd DFFSR_52/S FILL
XFILL_2_OAI21X1_108 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_0_OAI21X1_66 INVX1_4/gnd DFFSR_51/S FILL
XFILL_12_DFFSR_22 BUFX2_8/gnd DFFSR_10/S FILL
XDFFSR_2 DFFSR_2/Q DFFSR_2/CLK DFFSR_6/R DFFSR_2/S DFFSR_2/D DFFSR_5/gnd DFFSR_2/S
+ DFFSR
XFILL_2_NAND2X1_222 INVX1_23/gnd DFFSR_186/S FILL
XFILL_0_DFFSR_157 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_47_DFFSR_39 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_36_DFFSR_79 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_3_INVX1_131 INVX1_89/gnd DFFSR_36/S FILL
XFILL_41_DFFSR_188 INVX1_2/gnd DFFSR_1/S FILL
XFILL_31_DFFSR_191 INVX1_23/gnd DFFSR_91/S FILL
XFILL_1_NAND3X1_120 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_0_OAI21X1_204 BUFX2_36/A DFFSR_6/S FILL
XFILL_3_DFFSR_36 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_6_NAND2X1_27 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_20_DFFSR_29 INVX1_4/gnd DFFSR_4/S FILL
XFILL_6_OAI21X1_12 BUFX2_35/A DFFSR_14/S FILL
XFILL_3_NAND2X1_156 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_5_NAND2X1_30 DFFSR_79/gnd DFFSR_36/S FILL
XNAND2X1_27 DFFSR_1/S INVX1_22/A DFFSR_1/gnd OAI21X1_27/C DFFSR_1/S NAND2X1
XFILL_43_4_0 INVX1_4/gnd DFFSR_51/S FILL
XOAI21X1_12 DFFSR_12/S INVX1_14/Y OAI21X1_12/C BUFX2_35/A DFFSR_12/D DFFSR_14/S OAI21X1
XFILL_4_NAND2X1_33 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_5_OAI21X1_15 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_1_INVX1_348 INVX1_4/gnd DFFSR_4/S FILL
XFILL_44_DFFSR_115 BUFX2_6/gnd DFFSR_14/S FILL
XDFFPOSX1_30 NOR2X1_1/A CLKBUF1_11/Y AOI21X1_47/Y BUFX2_43/A DFFSR_97/S DFFPOSX1
XFILL_3_NAND2X1_36 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_4_OAI21X1_18 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_7_DFFSR_191 INVX1_23/gnd DFFSR_91/S FILL
XFILL_15_DFFPOSX1_13 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_2_NAND2X1_39 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_29_DFFSR_2 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_44_DFFSR_86 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_3_OAI21X1_21 INVX1_2/gnd DFFSR_51/S FILL
XFILL_1_OAI21X1_138 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_1_NAND2X1_42 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_34_DFFSR_118 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_2_OAI21X1_24 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_0_INVX1_168 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_8_NAND3X1_98 BUFX2_35/A DFFSR_14/S FILL
XFILL_24_DFFSR_121 BUFX2_36/A DFFSR_6/S FILL
XFILL_17_DFFSR_76 BUFX2_7/gnd DFFSR_54/S FILL
XAOI21X1_6 NAND3X1_8/Y NAND3X1_7/Y AOI21X1_6/C BUFX2_19/gnd AOI21X1_6/Y DFFSR_54/S
+ AOI21X1
XFILL_0_DFFSR_83 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_28_DFFSR_36 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_0_NAND2X1_45 INVX1_89/gnd DFFSR_36/S FILL
XFILL_1_OAI21X1_27 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_0_INVX1_30 DFFSR_1/gnd DFFSR_9/S FILL
XINVX1_278 INVX1_66/A DFFSR_3/gnd INVX1_278/Y DFFSR_4/S INVX1
XFILL_0_OAI21X1_30 INVX1_89/gnd DFFSR_36/S FILL
XFILL_14_DFFSR_124 INVX1_89/gnd DFFSR_36/S FILL
XFILL_1_NAND2X1_252 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_4_AOI21X1_3 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_5_DFFPOSX1_24 BUFX2_43/A DFFSR_23/S FILL
XFILL_0_DFFSR_121 BUFX2_36/A DFFSR_6/S FILL
XFILL_2_NAND2X1_186 BUFX2_37/A DFFSR_81/S FILL
XFILL_41_DFFSR_152 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_25_DFFSR_83 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_36_DFFSR_43 INVX1_94/gnd DFFSR_25/S FILL
XFILL_8_DFFSR_90 INVX1_2/gnd DFFSR_1/S FILL
XFILL_31_DFFSR_155 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_4_AOI22X1_11 INVX1_23/gnd DFFSR_91/S FILL
XFILL_21_DFFSR_158 BUFX2_43/A DFFSR_23/S FILL
XFILL_11_DFFSR_161 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_9_OAI21X1_223 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_0_OAI21X1_168 BUFX2_36/A DFFSR_6/S FILL
XFILL_6_NAND3X1_2 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_3_AOI22X1_14 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_3_NAND2X1_120 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_1_INVX1_312 BUFX2_36/A DFFSR_6/S FILL
XFILL_6_NOR2X1_37 INVX1_94/gnd DFFSR_25/S FILL
XINVX1_4 DFFSR_3/Q INVX1_4/gnd INVX1_4/Y DFFSR_4/S INVX1
XFILL_11_OAI22X1_38 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_0_NAND2X1_282 INVX1_89/gnd DFFSR_2/S FILL
XFILL_44_DFFSR_50 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_10_OAI22X1_41 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_7_DFFSR_155 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_1_OAI21X1_102 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_33_DFFSR_90 INVX1_2/gnd DFFSR_1/S FILL
XFILL_48_DFFSR_186 INVX1_23/gnd DFFSR_186/S FILL
XFILL_8_NAND3X1_62 BUFX2_43/A DFFSR_23/S FILL
XFILL_9_OAI22X1_44 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_7_NAND3X1_65 BUFX2_35/A DFFSR_14/S FILL
XFILL_0_INVX1_132 BUFX2_35/A DFFSR_97/S FILL
XINVX1_242 AND2X2_10/B BUFX2_36/A NOR2X1_10/B DFFSR_6/S INVX1
XFILL_8_OAI22X1_47 BUFX2_37/A DFFSR_8/S FILL
XFILL_0_DFFSR_47 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_17_DFFSR_40 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_38_DFFSR_189 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_6_NAND3X1_68 BUFX2_35/A DFFSR_14/S FILL
XFILL_1_NAND2X1_216 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_7_OAI22X1_50 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_5_NAND3X1_71 BUFX2_35/A DFFSR_14/S FILL
XFILL_6_OAI22X1_53 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_4_NAND3X1_74 BUFX2_35/A DFFSR_14/S FILL
XNAND3X1_68 NAND3X1_64/Y NAND3X1_68/B NAND3X1_67/C BUFX2_35/A INVX1_255/A DFFSR_14/S
+ NAND3X1
XFILL_0_NAND3X1_114 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_41_DFFSR_97 BUFX2_35/A DFFSR_97/S FILL
XFILL_5_OAI22X1_56 BUFX2_37/A DFFSR_8/S FILL
XFILL_17_2_0 BUFX2_7/gnd DFFSR_54/S FILL
XOAI22X1_53 INVX1_365/Y OAI22X1_49/D INVX1_364/Y OAI22X1_52/D DFFSR_71/gnd NOR2X1_36/B
+ DFFSR_10/S OAI22X1
XFILL_8_OAI21X1_253 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_2_AND2X2_6 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_3_NAND3X1_77 BUFX2_37/A DFFSR_81/S FILL
XFILL_2_NAND2X1_150 BUFX2_37/A DFFSR_81/S FILL
XFILL_4_OAI22X1_59 INVX1_8/gnd DFFSR_7/S FILL
XFILL_15_4_1 BUFX2_37/A DFFSR_81/S FILL
XFILL_8_DFFSR_54 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_2_NAND3X1_80 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_3_OAI22X1_62 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_25_DFFSR_47 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_41_DFFSR_116 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_14_DFFSR_87 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_1_NAND3X1_83 BUFX2_37/A DFFSR_81/S FILL
XFILL_31_DFFSR_119 BUFX2_37/A DFFSR_81/S FILL
XFILL_2_OAI22X1_65 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_0_NAND3X1_86 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_21_DFFSR_122 INVX1_94/gnd DFFSR_52/S FILL
XFILL_1_OAI22X1_68 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_0_OAI21X1_132 INVX1_4/gnd DFFSR_4/S FILL
XFILL_11_DFFSR_125 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_1_AOI21X1_4 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_1_INVX1_276 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_20_DFFSR_9 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_44_DFFSR_14 BUFX2_35/A DFFSR_14/S FILL
XFILL_7_DFFSR_119 BUFX2_37/A DFFSR_81/S FILL
XFILL_33_DFFSR_54 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_0_NAND2X1_246 INVX1_94/gnd DFFSR_25/S FILL
XINVX1_88 INVX1_88/A INVX1_2/gnd INVX1_88/Y DFFSR_1/S INVX1
XFILL_22_DFFSR_94 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_9_NAND3X1_23 BUFX2_37/A DFFSR_81/S FILL
XFILL_48_DFFSR_150 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_38_DFFSR_153 BUFX2_36/A DFFSR_8/S FILL
XFILL_8_NAND3X1_26 BUFX2_7/gnd DFFSR_81/S FILL
XINVX1_206 AND2X2_9/B BUFX2_19/gnd INVX1_206/Y DFFSR_54/S INVX1
XFILL_0_DFFSR_11 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_28_DFFSR_156 INVX1_23/gnd DFFSR_91/S FILL
XFILL_4_BUFX2_39 BUFX2_43/A DFFSR_97/S FILL
XFILL_4_DFFPOSX1_18 BUFX2_37/A DFFSR_8/S FILL
XFILL_7_NAND3X1_29 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_8_OAI22X1_11 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_18_DFFSR_159 BUFX2_36/A DFFSR_6/S FILL
XFILL_1_NAND2X1_180 INVX1_94/gnd DFFSR_52/S FILL
XFILL_6_NAND3X1_32 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_7_OAI22X1_14 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_5_NAND3X1_35 BUFX2_35/A DFFSR_97/S FILL
XFILL_3_NAND3X1_3 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_6_OAI22X1_17 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_41_DFFSR_5 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_4_NAND3X1_38 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_41_DFFSR_61 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_2_INVX1_95 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_5_OAI22X1_20 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_9_NAND3X1_133 INVX1_8/gnd DFFSR_5/S FILL
XFILL_3_NOR2X1_38 BUFX2_17/gnd DFFSR_7/S FILL
XNAND3X1_32 INVX1_235/A AOI21X1_13/B NAND3X1_58/A DFFSR_73/gnd INVX1_237/A DFFSR_57/S
+ NAND3X1
XFILL_3_NAND3X1_41 BUFX2_43/A DFFSR_23/S FILL
XDFFSR_159 BUFX2_2/A CLKBUF1_15/Y DFFSR_159/R DFFSR_8/S DFFSR_159/D BUFX2_36/A DFFSR_6/S
+ DFFSR
XOAI22X1_17 INVX1_289/Y OAI22X1_6/D INVX1_290/Y OAI22X1_9/B BUFX2_8/gnd NOR2X1_18/B
+ DFFSR_25/S OAI22X1
XFILL_4_OAI22X1_23 INVX1_89/gnd DFFSR_2/S FILL
XFILL_2_NAND2X1_114 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_8_OAI21X1_217 INVX1_23/gnd DFFSR_91/S FILL
XFILL_2_NAND3X1_44 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_3_OAI22X1_26 INVX1_94/gnd DFFSR_52/S FILL
XFILL_8_DFFSR_18 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_2_INVX1_420 INVX1_2/gnd DFFSR_51/S FILL
XFILL_25_DFFSR_11 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_4_DFFSR_156 INVX1_23/gnd DFFSR_91/S FILL
XFILL_1_NAND3X1_47 BUFX2_43/A DFFSR_97/S FILL
XFILL_2_OAI22X1_29 INVX1_8/gnd DFFSR_5/S FILL
XFILL_14_DFFSR_51 INVX1_2/gnd DFFSR_51/S FILL
XFILL_0_NAND3X1_50 BUFX2_37/A DFFSR_81/S FILL
XFILL_23_1_2 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_1_OAI22X1_32 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_45_DFFSR_187 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_5_0_1 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_23_DFFPOSX1_26 BUFX2_37/A DFFSR_81/S FILL
XFILL_0_OAI22X1_35 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_35_DFFSR_190 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_1_INVX1_240 BUFX2_35/A DFFSR_14/S FILL
XFILL_49_DFFSR_68 BUFX2_35/A DFFSR_14/S FILL
XFILL_3_2_2 INVX1_23/gnd DFFSR_91/S FILL
XFILL_0_NAND2X1_210 BUFX2_35/A DFFSR_97/S FILL
XINVX1_52 DFFSR_46/Q BUFX2_37/A INVX1_52/Y DFFSR_81/S INVX1
XFILL_5_DFFSR_65 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_48_DFFSR_114 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_11_DFFSR_98 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_33_DFFSR_18 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_22_DFFSR_58 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_38_DFFSR_117 INVX1_23/gnd DFFSR_91/S FILL
XINVX1_170 DFFSR_148/Q BUFX2_6/gnd INVX1_170/Y DFFSR_91/S INVX1
XFILL_4_INVX1_167 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_1_NAND2X1_144 INVX1_8/gnd DFFSR_7/S FILL
XFILL_7_OAI21X1_247 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_28_DFFSR_120 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_18_DFFSR_123 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_8_AOI21X1_2 INVX1_94/gnd DFFSR_52/S FILL
XFILL_2_INVX1_59 INVX1_94/gnd DFFSR_25/S FILL
XFILL_41_DFFSR_25 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_30_DFFSR_65 DFFSR_3/gnd DFFSR_65/S FILL
XDFFSR_123 DFFSR_123/Q CLKBUF1_7/Y DFFSR_123/R DFFSR_186/S DFFSR_123/D DFFSR_89/gnd
+ DFFSR_186/S DFFSR
XFILL_2_INVX1_384 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_8_OAI21X1_181 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_14_DFFSR_15 INVX1_8/gnd DFFSR_7/S FILL
XFILL_4_DFFSR_120 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_45_DFFSR_151 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_1_NAND3X1_11 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_35_DFFSR_154 BUFX2_36/A DFFSR_6/S FILL
XFILL_8_DFFSR_8 BUFX2_36/A DFFSR_8/S FILL
XFILL_0_NAND3X1_14 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_25_DFFSR_157 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_1_INVX1_204 BUFX2_36/A DFFSR_8/S FILL
XFILL_38_DFFSR_72 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_15_DFFSR_160 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_49_DFFSR_32 INVX1_2/gnd DFFSR_1/S FILL
XFILL_0_NAND3X1_4 INVX1_94/gnd DFFSR_52/S FILL
XFILL_3_DFFPOSX1_12 INVX1_8/gnd DFFSR_5/S FILL
XFILL_0_NAND2X1_174 BUFX2_43/A DFFSR_97/S FILL
XINVX1_16 DFFSR_14/Q BUFX2_43/A INVX1_16/Y DFFSR_23/S INVX1
XDFFSR_69 DFFSR_69/Q INVX1_172/A DFFSR_68/R DFFSR_23/S DFFSR_69/D BUFX2_43/A DFFSR_23/S
+ DFFSR
XFILL_11_DFFSR_62 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_22_DFFSR_22 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_0_NOR2X1_39 INVX1_8/gnd DFFSR_5/S FILL
XFILL_5_DFFSR_29 INVX1_4/gnd DFFSR_4/S FILL
XINVX1_134 INVX1_134/A BUFX2_37/A INVX1_134/Y DFFSR_8/S INVX1
XFILL_8_NAND3X1_127 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_1_DFFSR_157 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_12_DFFPOSX1_31 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_1_NAND2X1_108 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_7_OAI21X1_211 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_46_DFFSR_79 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_4_INVX1_131 INVX1_89/gnd DFFSR_36/S FILL
XFILL_42_DFFSR_188 INVX1_2/gnd DFFSR_1/S FILL
XFILL_32_DFFSR_191 INVX1_23/gnd DFFSR_91/S FILL
XFILL_2_INVX1_23 INVX1_23/gnd DFFSR_91/S FILL
XFILL_19_DFFSR_69 BUFX2_43/A DFFSR_23/S FILL
XFILL_2_DFFSR_76 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_30_DFFSR_29 INVX1_4/gnd DFFSR_4/S FILL
XFILL_8_OAI21X1_145 INVX1_23/gnd DFFSR_91/S FILL
XFILL_22_DFFPOSX1_20 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_2_INVX1_348 INVX1_4/gnd DFFSR_4/S FILL
XFILL_6_XOR2X1_6 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_1_BUFX2_14 BUFX2_37/A DFFSR_81/S FILL
XFILL_8_DFFSR_191 INVX1_23/gnd DFFSR_91/S FILL
XFILL_45_DFFSR_115 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_35_DFFSR_118 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_1_INVX1_168 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_25_DFFSR_121 BUFX2_36/A DFFSR_6/S FILL
XFILL_27_DFFSR_76 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_38_DFFSR_36 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_24_2_0 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_15_DFFSR_124 INVX1_89/gnd DFFSR_36/S FILL
XFILL_6_OAI21X1_241 BUFX2_35/A DFFSR_97/S FILL
XDFFSR_33 DFFSR_33/Q DFFSR_28/CLK DFFSR_33/R DFFSR_52/S DFFSR_33/D INVX1_94/gnd DFFSR_52/S
+ DFFSR
XFILL_5_AOI21X1_3 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_0_NAND2X1_138 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_11_DFFSR_26 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_22_4_1 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_4_3_0 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_1_DFFSR_121 BUFX2_36/A DFFSR_6/S FILL
XFILL_7_OAI21X1_175 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_42_DFFSR_152 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_35_DFFSR_83 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_46_DFFSR_43 INVX1_94/gnd DFFSR_25/S FILL
XFILL_34_5 INVX1_8/gnd DFFSR_7/S FILL
XFILL_2_5_1 INVX1_23/gnd DFFSR_186/S FILL
XFILL_32_DFFSR_155 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_22_DFFSR_158 BUFX2_43/A DFFSR_23/S FILL
XFILL_12_DFFSR_161 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_19_DFFSR_33 INVX1_94/gnd DFFSR_52/S FILL
XFILL_7_NAND3X1_2 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_2_DFFSR_40 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_8_OAI21X1_109 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_2_INVX1_312 BUFX2_36/A DFFSR_6/S FILL
XFILL_20_CLKBUF1_23 INVX1_89/gnd DFFSR_2/S FILL
XFILL_19_DFFSR_6 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_12_XOR2X1_3 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_8_DFFSR_155 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_43_DFFSR_90 INVX1_2/gnd DFFSR_1/S FILL
XFILL_49_DFFSR_186 INVX1_23/gnd DFFSR_186/S FILL
XFILL_1_INVX1_132 BUFX2_35/A DFFSR_97/S FILL
XFILL_27_DFFSR_40 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_7_NAND3X1_121 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_39_DFFSR_189 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_16_DFFSR_80 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_3_BUFX2_7 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_11_DFFPOSX1_25 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_6_OAI21X1_205 BUFX2_36/A DFFSR_8/S FILL
XFILL_0_NAND2X1_102 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_51_DFFSR_97 BUFX2_35/A DFFSR_97/S FILL
XFILL_40_DFFSR_2 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_30_1_2 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_21_DFFPOSX1_14 BUFX2_6/gnd DFFSR_14/S FILL
XOAI21X1_241 NOR2X1_44/A AND2X2_14/B INVX1_400/Y BUFX2_35/A NOR2X1_45/B DFFSR_97/S
+ OAI21X1
XFILL_35_DFFSR_47 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_42_DFFSR_116 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_24_DFFSR_87 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_7_OAI21X1_139 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_7_DFFSR_94 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_32_DFFSR_119 BUFX2_37/A DFFSR_81/S FILL
XFILL_22_DFFSR_122 INVX1_94/gnd DFFSR_52/S FILL
XFILL_12_DFFSR_125 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_6_BUFX2_32 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_2_AOI21X1_4 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_2_INVX1_276 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_8_DFFSR_119 BUFX2_37/A DFFSR_81/S FILL
XFILL_43_DFFSR_54 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_4_INVX1_88 INVX1_2/gnd DFFSR_1/S FILL
XFILL_32_DFFSR_94 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_5_OAI21X1_235 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_49_DFFSR_150 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_39_DFFSR_153 BUFX2_36/A DFFSR_8/S FILL
XFILL_16_DFFSR_44 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_29_DFFSR_156 INVX1_23/gnd DFFSR_91/S FILL
XFILL_19_DFFSR_159 BUFX2_36/A DFFSR_6/S FILL
XFILL_6_OAI21X1_169 BUFX2_36/A DFFSR_8/S FILL
XNAND3X1_6 AOI21X1_1/C INVX1_223/A AOI21X1_1/A INVX1_8/gnd NAND3X1_6/Y DFFSR_7/S NAND3X1
XFILL_4_NAND3X1_3 BUFX2_19/gnd DFFSR_54/S FILL
XNOR2X1_41 NOR2X1_41/A NOR2X1_41/B BUFX2_8/gnd NOR2X1_41/Y DFFSR_10/S NOR2X1
XFILL_4_NOR2X1_38 BUFX2_17/gnd DFFSR_7/S FILL
XOAI21X1_205 AOI22X1_7/Y AOI22X1_8/Y AOI21X1_23/C BUFX2_36/A NAND3X1_52/B DFFSR_8/S
+ OAI21X1
XFILL_12_CLKBUF1_11 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_6_NAND2X1_283 INVX1_89/gnd DFFSR_36/S FILL
XFILL_7_OAI21X1_103 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_3_INVX1_420 INVX1_2/gnd DFFSR_51/S FILL
XFILL_7_DFFSR_58 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_35_DFFSR_11 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_5_DFFSR_156 INVX1_23/gnd DFFSR_91/S FILL
XFILL_13_DFFSR_91 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_11_CLKBUF1_14 BUFX2_43/A DFFSR_23/S FILL
XFILL_24_DFFSR_51 INVX1_2/gnd DFFSR_51/S FILL
XFILL_10_CLKBUF1_17 INVX1_94/gnd DFFSR_25/S FILL
XFILL_46_DFFSR_187 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_4_OAI21X1_265 BUFX2_43/A DFFSR_97/S FILL
XFILL_36_DFFSR_190 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_2_INVX1_240 BUFX2_35/A DFFSR_14/S FILL
XFILL_7_DFFSR_5 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_9_CLKBUF1_20 INVX1_4/gnd DFFSR_51/S FILL
XFILL_6_NAND3X1_115 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_8_CLKBUF1_23 INVX1_89/gnd DFFSR_2/S FILL
XFILL_10_DFFPOSX1_19 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_4_INVX1_52 BUFX2_37/A DFFSR_81/S FILL
XFILL_5_OAI21X1_199 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_21_DFFSR_98 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_43_DFFSR_18 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_32_DFFSR_58 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_49_DFFSR_114 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_39_DFFSR_117 INVX1_23/gnd DFFSR_91/S FILL
XFILL_3_BUFX2_43 BUFX2_35/A DFFSR_97/S FILL
XFILL_29_DFFSR_120 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_19_DFFSR_123 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_6_OAI21X1_133 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_31_DFFSR_9 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_0_DFFPOSX1_30 BUFX2_43/A DFFSR_97/S FILL
XFILL_1_INVX1_99 INVX1_4/gnd DFFSR_4/S FILL
XFILL_40_DFFSR_65 DFFSR_3/gnd DFFSR_65/S FILL
XOAI21X1_169 DFFSR_8/S INVX1_204/Y NAND2X1_169/Y BUFX2_36/A DFFSR_169/D DFFSR_8/S
+ OAI21X1
XFILL_16_2 BUFX2_37/A DFFSR_81/S FILL
XFILL_3_INVX1_384 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_6_NAND2X1_247 INVX1_8/gnd DFFSR_5/S FILL
XFILL_7_DFFSR_22 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_13_DFFSR_55 INVX1_89/gnd DFFSR_36/S FILL
XFILL_24_DFFSR_15 INVX1_8/gnd DFFSR_7/S FILL
XFILL_5_DFFSR_120 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_46_DFFSR_151 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_36_DFFSR_154 BUFX2_36/A DFFSR_6/S FILL
XNAND2X1_283 AOI22X1_14/A AOI22X1_14/B INVX1_89/gnd NOR2X1_51/A DFFSR_36/S NAND2X1
XFILL_31_2_0 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_26_DFFSR_157 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_6_NOR2X1_3 INVX1_94/gnd DFFSR_25/S FILL
XFILL_4_OAI21X1_229 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_2_INVX1_204 BUFX2_36/A DFFSR_8/S FILL
XFILL_29_4_1 INVX1_89/gnd DFFSR_2/S FILL
XFILL_48_DFFSR_72 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_16_DFFSR_160 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_1_NAND3X1_4 INVX1_94/gnd DFFSR_52/S FILL
XFILL_4_DFFSR_69 BUFX2_43/A DFFSR_23/S FILL
XFILL_21_DFFSR_62 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_32_DFFSR_22 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_1_NOR2X1_39 INVX1_8/gnd DFFSR_5/S FILL
XFILL_5_OAI21X1_163 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_9_5_1 BUFX2_43/A DFFSR_23/S FILL
XNAND3X1_115 NOR2X1_1/B NOR2X1_1/A INVX1_265/Y BUFX2_8/gnd OAI22X1_7/B DFFSR_10/S
+ NAND3X1
XFILL_0_INVX1_421 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_2_DFFSR_157 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_5_NAND2X1_277 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_43_DFFSR_188 INVX1_2/gnd DFFSR_1/S FILL
XFILL_33_DFFSR_191 INVX1_23/gnd DFFSR_91/S FILL
XFILL_29_DFFSR_69 BUFX2_43/A DFFSR_23/S FILL
XFILL_1_INVX1_63 INVX1_2/gnd DFFSR_51/S FILL
XFILL_40_DFFSR_29 INVX1_4/gnd DFFSR_4/S FILL
XFILL_3_OAI21X1_259 INVX1_23/gnd DFFSR_186/S FILL
XOAI21X1_133 DFFSR_81/S INVX1_150/Y OAI21X1_133/C BUFX2_7/gnd DFFSR_133/D DFFSR_81/S
+ OAI21X1
XFILL_0_CLKBUF1_11 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_6_NAND2X1_211 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_3_INVX1_348 INVX1_4/gnd DFFSR_4/S FILL
XFILL_13_DFFSR_19 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_9_DFFSR_191 INVX1_23/gnd DFFSR_91/S FILL
XFILL_46_DFFSR_115 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_5_NAND3X1_109 BUFX2_36/A DFFSR_8/S FILL
XFILL_4_OAI21X1_193 BUFX2_7/gnd DFFSR_54/S FILL
XNAND2X1_247 NOR2X1_38/Y NOR2X1_39/Y INVX1_8/gnd NAND2X1_142/B DFFSR_5/S NAND2X1
XFILL_18_DFFSR_3 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_36_DFFSR_118 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_2_INVX1_168 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_26_DFFSR_121 BUFX2_36/A DFFSR_6/S FILL
XFILL_37_DFFSR_76 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_48_DFFSR_36 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_16_DFFSR_124 INVX1_89/gnd DFFSR_36/S FILL
XFILL_37_1_2 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_6_AOI21X1_3 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_5_OAI21X1_127 BUFX2_43/A DFFSR_23/S FILL
XFILL_4_DFFSR_33 INVX1_94/gnd DFFSR_52/S FILL
XFILL_2_BUFX2_4 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_21_DFFSR_26 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_10_DFFSR_66 INVX1_2/gnd DFFSR_51/S FILL
XFILL_0_INVX1_385 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_2_DFFSR_121 BUFX2_36/A DFFSR_6/S FILL
XFILL_21_7 INVX1_94/gnd DFFSR_52/S FILL
XFILL_43_DFFSR_152 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_38_2 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_33_DFFSR_155 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_45_DFFSR_83 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_5_NAND2X1_241 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_23_DFFSR_158 BUFX2_43/A DFFSR_23/S FILL
XFILL_13_DFFSR_161 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_29_DFFSR_33 INVX1_94/gnd DFFSR_52/S FILL
XFILL_8_NAND3X1_2 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_1_DFFSR_80 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_18_DFFSR_73 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_1_INVX1_27 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_3_OAI21X1_223 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_9_DFFPOSX1_13 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_6_NAND2X1_175 BUFX2_35/A DFFSR_14/S FILL
XFILL_3_INVX1_312 BUFX2_36/A DFFSR_6/S FILL
XFILL_23_DFFPOSX1_2 INVX1_89/gnd DFFSR_36/S FILL
XFILL_22_DFFPOSX1_5 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_21_DFFPOSX1_8 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_0_BUFX2_18 DFFSR_3/gnd DFFSR_65/S FILL
XNAND2X1_211 AND2X2_5/B AND2X2_9/B BUFX2_6/gnd XOR2X1_4/B DFFSR_91/S NAND2X1
XFILL_9_DFFSR_155 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_50_DFFSR_186 INVX1_23/gnd DFFSR_186/S FILL
XFILL_4_OAI21X1_157 BUFX2_35/A DFFSR_97/S FILL
XFILL_2_INVX1_132 BUFX2_35/A DFFSR_97/S FILL
XFILL_37_DFFSR_40 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_40_DFFSR_189 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_9_DFFSR_87 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_26_DFFSR_80 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_10_DFFSR_30 INVX1_89/gnd DFFSR_36/S FILL
XFILL_4_NAND2X1_271 INVX1_89/gnd DFFSR_2/S FILL
XFILL_0_INVX1_349 INVX1_89/gnd DFFSR_2/S FILL
XFILL_2_OAI21X1_253 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_5_NAND2X1_205 BUFX2_36/A DFFSR_6/S FILL
XFILL_45_DFFSR_47 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_43_DFFSR_116 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_34_DFFSR_87 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_33_DFFSR_119 BUFX2_37/A DFFSR_81/S FILL
XFILL_4_NAND3X1_103 INVX1_23/gnd DFFSR_186/S FILL
XFILL_23_DFFSR_122 INVX1_94/gnd DFFSR_52/S FILL
XFILL_1_DFFSR_44 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_18_DFFSR_37 INVX1_89/gnd DFFSR_2/S FILL
XFILL_13_DFFSR_125 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_3_OAI21X1_187 BUFX2_37/A DFFSR_8/S FILL
XFILL_3_AOI21X1_4 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_6_NAND2X1_139 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_3_INVX1_276 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_6_DFFSR_2 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_11_XOR2X1_7 INVX1_23/gnd DFFSR_91/S FILL
XFILL_9_DFFSR_119 BUFX2_37/A DFFSR_81/S FILL
XFILL_42_DFFSR_94 BUFX2_16/gnd DFFSR_65/S FILL
XNAND2X1_175 DFFSR_12/S BUFX2_35/A BUFX2_35/A OAI21X1_175/C DFFSR_14/S NAND2X1
XFILL_4_OAI21X1_121 BUFX2_36/A DFFSR_8/S FILL
XFILL_50_DFFSR_150 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_40_DFFSR_153 BUFX2_36/A DFFSR_8/S FILL
XFILL_26_DFFSR_44 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_3_AND2X2_3 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_9_DFFSR_51 INVX1_2/gnd DFFSR_51/S FILL
XFILL_30_DFFSR_156 INVX1_23/gnd DFFSR_91/S FILL
XFILL_15_DFFSR_84 BUFX2_43/A DFFSR_23/S FILL
XFILL_43_7 INVX1_4/gnd DFFSR_4/S FILL
XFILL_4_OR2X2_2 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_20_DFFSR_159 BUFX2_36/A DFFSR_6/S FILL
XFILL_10_DFFSR_162 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_5_NAND3X1_3 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_4_NAND2X1_235 INVX1_4/gnd DFFSR_51/S FILL
XINVX1_423 BUFX2_7/Y BUFX2_37/A DFFSR_185/R DFFSR_8/S INVX1
XFILL_0_INVX1_313 INVX1_8/gnd DFFSR_5/S FILL
XFILL_30_DFFSR_6 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_3_NAND3X1_133 INVX1_8/gnd DFFSR_5/S FILL
XFILL_5_NOR2X1_38 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_38_2_0 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_2_OAI21X1_217 INVX1_23/gnd DFFSR_91/S FILL
XFILL_5_NAND2X1_169 BUFX2_36/A DFFSR_8/S FILL
XFILL_4_INVX1_420 INVX1_2/gnd DFFSR_51/S FILL
XFILL_6_DFFSR_156 INVX1_23/gnd DFFSR_91/S FILL
XFILL_23_DFFSR_91 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_36_4_1 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_6_DFFSR_98 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_34_DFFSR_51 INVX1_2/gnd DFFSR_51/S FILL
XFILL_45_DFFSR_11 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_11_DFFPOSX1_2 INVX1_89/gnd DFFSR_36/S FILL
XFILL_47_DFFSR_187 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_5_BUFX2_36 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_37_DFFSR_190 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_10_DFFPOSX1_5 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_3_INVX1_240 BUFX2_35/A DFFSR_14/S FILL
XFILL_17_DFFPOSX1_26 BUFX2_37/A DFFSR_81/S FILL
XFILL_3_OAI21X1_151 BUFX2_37/A DFFSR_81/S FILL
XFILL_6_NAND2X1_103 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_9_DFFPOSX1_8 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_3_NAND2X1_265 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_3_INVX1_92 BUFX2_19/gnd DFFSR_54/S FILL
XNAND2X1_139 DFFSR_57/S NAND2X1_244/Y BUFX2_17/gnd NAND2X1_139/Y DFFSR_57/S NAND2X1
XFILL_31_DFFSR_98 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_42_DFFSR_58 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_8_AOI21X1_31 INVX1_23/gnd DFFSR_186/S FILL
XFILL_27_DFFPOSX1_15 BUFX2_35/A DFFSR_14/S FILL
XFILL_50_DFFSR_114 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_40_DFFSR_117 INVX1_23/gnd DFFSR_91/S FILL
XFILL_7_AOI21X1_34 INVX1_94/gnd DFFSR_25/S FILL
XFILL_9_DFFSR_15 INVX1_8/gnd DFFSR_7/S FILL
XFILL_15_DFFSR_48 INVX1_4/gnd DFFSR_4/S FILL
XFILL_6_AOI21X1_37 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_30_DFFSR_120 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_20_DFFSR_123 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_4_NAND2X1_199 BUFX2_36/A DFFSR_8/S FILL
XFILL_1_OAI21X1_247 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_5_AOI21X1_40 DFFSR_3/gnd DFFSR_4/S FILL
XAOI21X1_37 AOI21X1_37/A INVX1_261/A BUFX2_4/Y BUFX2_8/gnd AOI21X1_37/Y DFFSR_25/S
+ AOI21X1
XFILL_4_AOI21X1_43 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_10_DFFSR_126 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_0_AOI21X1_5 BUFX2_37/A DFFSR_81/S FILL
XINVX1_387 INVX1_387/A INVX1_94/gnd INVX1_387/Y DFFSR_25/S INVX1
XFILL_3_AOI21X1_46 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_0_INVX1_277 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_50_DFFSR_65 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_4_INVX1_384 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_5_NAND2X1_133 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_6_DFFSR_62 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_12_DFFSR_95 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_23_DFFSR_55 INVX1_89/gnd DFFSR_36/S FILL
XFILL_34_DFFSR_15 INVX1_8/gnd DFFSR_7/S FILL
XFILL_2_OAI21X1_181 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_6_DFFSR_120 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_47_DFFSR_151 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_37_DFFSR_154 BUFX2_36/A DFFSR_6/S FILL
XFILL_44_1_2 INVX1_2/gnd DFFSR_51/S FILL
XFILL_27_DFFSR_157 BUFX2_6/gnd DFFSR_91/S FILL
XBUFX2_40 BUFX2_35/A BUFX2_35/A BUFX2_40/Y DFFSR_14/S BUFX2
XFILL_3_OAI21X1_115 BUFX2_36/A DFFSR_6/S FILL
XFILL_3_INVX1_204 BUFX2_36/A DFFSR_8/S FILL
XFILL_17_DFFSR_160 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_2_NAND3X1_4 INVX1_94/gnd DFFSR_52/S FILL
XFILL_8_OAI21X1_79 INVX1_89/gnd DFFSR_36/S FILL
XFILL_31_DFFSR_62 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_42_DFFSR_22 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_7_OAI21X1_82 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_3_INVX1_56 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_3_NAND2X1_229 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_6_OAI21X1_85 DFFSR_79/gnd DFFSR_45/S FILL
XNAND2X1_103 BUFX2_22/Y DFFSR_95/Q DFFSR_5/gnd NAND2X1_103/Y DFFSR_2/S NAND2X1
XFILL_2_NOR2X1_39 INVX1_8/gnd DFFSR_5/S FILL
XFILL_12_0_0 BUFX2_36/A DFFSR_6/S FILL
XFILL_1_BUFX2_1 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_1_INVX1_421 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_5_OAI21X1_88 INVX1_4/gnd DFFSR_4/S FILL
XFILL_3_DFFSR_157 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_15_DFFSR_12 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_4_OAI21X1_91 BUFX2_43/A DFFSR_97/S FILL
XOAI21X1_85 BUFX2_23/Y INVX1_96/Y OAI21X1_85/C DFFSR_79/gnd DFFSR_85/D DFFSR_45/S
+ OAI21X1
XFILL_2_NAND3X1_127 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_10_2_1 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_1_OAI21X1_211 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_44_DFFSR_188 INVX1_2/gnd DFFSR_1/S FILL
XFILL_3_OAI21X1_94 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_34_DFFSR_191 INVX1_23/gnd DFFSR_91/S FILL
XFILL_2_OAI21X1_97 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_4_NAND2X1_163 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_0_INVX1_241 BUFX2_43/A DFFSR_23/S FILL
XFILL_39_DFFSR_69 BUFX2_43/A DFFSR_23/S FILL
XINVX1_351 DFFSR_83/Q BUFX2_19/gnd INVX1_351/Y DFFSR_54/S INVX1
XFILL_50_DFFSR_29 INVX1_4/gnd DFFSR_4/S FILL
XFILL_3_3 INVX1_23/gnd DFFSR_186/S FILL
XFILL_3_AOI21X1_10 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_2_OAI21X1_145 INVX1_23/gnd DFFSR_91/S FILL
XFILL_16_DFFPOSX1_20 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_2_AOI21X1_13 INVX1_8/gnd DFFSR_7/S FILL
XFILL_4_INVX1_348 INVX1_4/gnd DFFSR_4/S FILL
XFILL_1_AOI21X1_16 BUFX2_43/A DFFSR_23/S FILL
XFILL_23_DFFSR_19 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_6_DFFSR_26 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_12_DFFSR_59 INVX1_4/gnd DFFSR_51/S FILL
XFILL_47_DFFSR_115 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_0_AOI21X1_19 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_5_NOR2X1_7 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_37_DFFSR_118 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_3_INVX1_168 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_27_DFFSR_121 BUFX2_36/A DFFSR_6/S FILL
XFILL_47_DFFSR_76 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_9_OAI21X1_40 INVX1_8/gnd DFFSR_7/S FILL
XFILL_42_DFFSR_9 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_2_NAND2X1_259 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_8_OAI21X1_43 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_17_DFFSR_124 INVX1_89/gnd DFFSR_36/S FILL
XFILL_7_OAI21X1_46 BUFX2_37/A DFFSR_81/S FILL
XFILL_7_AOI21X1_3 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_6_NAND2X1_64 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_0_OAI21X1_241 BUFX2_35/A DFFSR_97/S FILL
XFILL_3_NAND2X1_193 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_3_INVX1_20 INVX1_8/gnd DFFSR_5/S FILL
XFILL_6_DFFPOSX1_31 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_31_DFFSR_26 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_5_NAND2X1_67 INVX1_2/gnd DFFSR_1/S FILL
XFILL_20_DFFSR_66 INVX1_2/gnd DFFSR_51/S FILL
XFILL_3_DFFSR_73 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_6_OAI21X1_49 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_5_OAI21X1_52 INVX1_94/gnd DFFSR_25/S FILL
XFILL_1_INVX1_385 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_4_NAND2X1_70 DFFSR_5/gnd DFFSR_2/S FILL
XNAND2X1_64 DFFSR_11/S DFFSR_56/Q BUFX2_16/gnd NAND2X1_64/Y DFFSR_65/S NAND2X1
XFILL_3_DFFSR_121 BUFX2_36/A DFFSR_6/S FILL
XFILL_25_4 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_4_OAI21X1_55 INVX1_89/gnd DFFSR_2/S FILL
XFILL_3_NAND2X1_73 DFFSR_73/gnd DFFSR_11/S FILL
XOAI21X1_49 DFFSR_13/S INVX1_56/Y NAND2X1_49/Y DFFSR_73/gnd DFFSR_49/D DFFSR_11/S
+ OAI21X1
XFILL_44_DFFSR_152 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_2_BUFX2_11 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_2_NAND2X1_76 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_7_XOR2X1_3 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_3_OAI21X1_58 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_1_OAI21X1_175 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_4_NAND2X1_127 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_34_DFFSR_155 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_24_DFFSR_158 BUFX2_43/A DFFSR_23/S FILL
XFILL_2_OAI21X1_61 BUFX2_36/A DFFSR_8/S FILL
XFILL_1_NAND2X1_79 INVX1_89/gnd DFFSR_36/S FILL
XFILL_14_DFFSR_161 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_39_DFFSR_33 INVX1_94/gnd DFFSR_52/S FILL
XFILL_0_INVX1_205 INVX1_94/gnd DFFSR_25/S FILL
XINVX1_315 DFFSR_55/Q BUFX2_8/gnd INVX1_315/Y DFFSR_25/S INVX1
XFILL_0_NAND2X1_82 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_0_INVX1_67 INVX1_4/gnd DFFSR_51/S FILL
XFILL_1_OAI21X1_64 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_28_DFFSR_73 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_4_INVX1_312 BUFX2_36/A DFFSR_6/S FILL
XFILL_0_OAI21X1_67 INVX1_2/gnd DFFSR_1/S FILL
XFILL_12_DFFSR_23 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_2_OAI21X1_109 BUFX2_5/gnd DFFSR_6/S FILL
XDFFSR_3 DFFSR_3/Q DFFSR_3/CLK DFFSR_6/R DFFSR_3/S DFFSR_3/D DFFSR_3/gnd DFFSR_4/S
+ DFFSR
XFILL_51_DFFSR_186 INVX1_23/gnd DFFSR_186/S FILL
XFILL_2_NAND2X1_223 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_0_DFFSR_158 BUFX2_43/A DFFSR_23/S FILL
XFILL_3_INVX1_132 BUFX2_35/A DFFSR_97/S FILL
XFILL_47_DFFSR_40 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_41_DFFSR_189 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_36_DFFSR_80 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_1_NAND3X1_121 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_45_2_0 INVX1_2/gnd DFFSR_1/S FILL
XFILL_0_OAI21X1_205 BUFX2_36/A DFFSR_8/S FILL
XFILL_6_NAND2X1_28 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_7_OAI21X1_10 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_20_DFFSR_30 INVX1_89/gnd DFFSR_36/S FILL
XFILL_3_DFFSR_37 INVX1_89/gnd DFFSR_2/S FILL
XFILL_3_NAND2X1_157 BUFX2_35/A DFFSR_97/S FILL
XFILL_5_NAND2X1_31 BUFX2_43/A DFFSR_97/S FILL
XNAND2X1_28 DFFSR_81/S DFFSR_20/Q BUFX2_7/gnd OAI21X1_28/C DFFSR_81/S NAND2X1
XFILL_6_OAI21X1_13 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_9_OAI21X1_260 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_5_OAI21X1_16 INVX1_89/gnd DFFSR_36/S FILL
XFILL_1_INVX1_349 INVX1_89/gnd DFFSR_2/S FILL
XFILL_4_NAND2X1_34 INVX1_2/gnd DFFSR_1/S FILL
XFILL_43_4_1 INVX1_4/gnd DFFSR_51/S FILL
XOAI21X1_13 DFFSR_13/S INVX1_15/Y NAND2X1_13/Y BUFX2_16/gnd DFFSR_13/D DFFSR_65/S
+ OAI21X1
XFILL_3_NAND2X1_37 INVX1_8/gnd DFFSR_5/S FILL
XDFFPOSX1_31 NOR2X1_2/A CLKBUF1_13/Y AOI21X1_48/Y BUFX2_17/gnd DFFSR_57/S DFFPOSX1
XFILL_4_OAI21X1_19 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_15_DFFPOSX1_14 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_3_OAI21X1_22 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_44_DFFSR_116 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_44_DFFSR_87 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_29_DFFSR_3 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_1_OAI21X1_139 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_2_NAND2X1_40 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_34_DFFSR_119 BUFX2_37/A DFFSR_81/S FILL
XFILL_2_OAI21X1_25 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_1_NAND2X1_43 INVX1_89/gnd DFFSR_2/S FILL
XFILL_0_INVX1_169 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_8_NAND3X1_99 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_0_DFFSR_84 BUFX2_43/A DFFSR_23/S FILL
XFILL_1_OAI21X1_28 BUFX2_7/gnd DFFSR_81/S FILL
XAOI21X1_7 AOI21X1_7/A AOI21X1_7/B AOI21X1_7/C BUFX2_19/gnd NOR3X1_1/C DFFSR_54/S
+ AOI21X1
XFILL_24_DFFSR_122 INVX1_94/gnd DFFSR_52/S FILL
XFILL_0_NAND2X1_46 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_28_DFFSR_37 INVX1_89/gnd DFFSR_2/S FILL
XFILL_0_INVX1_31 INVX1_2/gnd DFFSR_1/S FILL
XINVX1_279 INVX1_39/A INVX1_4/gnd INVX1_279/Y DFFSR_51/S INVX1
XFILL_14_DFFSR_125 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_0_OAI21X1_31 BUFX2_35/A DFFSR_97/S FILL
XFILL_17_DFFSR_77 INVX1_89/gnd DFFSR_2/S FILL
XFILL_4_AOI21X1_4 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_1_NAND2X1_253 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_4_INVX1_276 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_5_DFFPOSX1_25 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_0_DFFSR_122 INVX1_94/gnd DFFSR_52/S FILL
XFILL_8_DFFSR_91 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_41_DFFSR_153 BUFX2_36/A DFFSR_8/S FILL
XFILL_2_NAND2X1_187 BUFX2_37/A DFFSR_8/S FILL
XFILL_31_DFFSR_156 INVX1_23/gnd DFFSR_91/S FILL
XFILL_25_DFFSR_84 BUFX2_43/A DFFSR_23/S FILL
XFILL_36_DFFSR_44 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_4_AOI22X1_12 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_21_DFFSR_159 BUFX2_36/A DFFSR_6/S FILL
XFILL_11_DFFSR_162 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_9_OAI21X1_224 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_0_OAI21X1_169 BUFX2_36/A DFFSR_8/S FILL
XFILL_3_NAND2X1_121 BUFX2_36/A DFFSR_8/S FILL
XFILL_6_NAND3X1_3 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_1_INVX1_313 INVX1_8/gnd DFFSR_5/S FILL
XINVX1_5 DFFSR_4/Q INVX1_4/gnd INVX1_5/Y DFFSR_51/S INVX1
XFILL_6_NOR2X1_38 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_0_NAND2X1_283 INVX1_89/gnd DFFSR_36/S FILL
XFILL_10_OAI22X1_42 INVX1_8/gnd DFFSR_7/S FILL
XFILL_7_DFFSR_156 INVX1_23/gnd DFFSR_91/S FILL
XFILL_33_DFFSR_91 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_1_OAI21X1_103 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_44_DFFSR_51 INVX1_2/gnd DFFSR_51/S FILL
XFILL_8_NAND3X1_63 BUFX2_43/A DFFSR_23/S FILL
XFILL_9_OAI22X1_45 INVX1_89/gnd DFFSR_2/S FILL
XFILL_48_DFFSR_187 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_7_NAND3X1_66 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_8_OAI22X1_48 BUFX2_37/A DFFSR_81/S FILL
XINVX1_243 INVX1_243/A DFFSR_71/gnd INVX1_243/Y DFFSR_10/S INVX1
XFILL_0_NAND2X1_10 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_17_DFFSR_41 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_38_DFFSR_190 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_0_DFFSR_48 INVX1_4/gnd DFFSR_4/S FILL
XFILL_0_INVX1_133 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_6_NAND3X1_69 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_1_NAND2X1_217 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_7_OAI22X1_51 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_19_0_0 BUFX2_19/gnd DFFSR_52/S FILL
XNAND3X1_69 NAND3X1_66/Y NAND3X1_67/B NAND3X1_69/C BUFX2_6/gnd AOI22X1_13/C DFFSR_14/S
+ NAND3X1
XFILL_5_NAND3X1_72 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_0_NAND3X1_115 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_6_OAI22X1_54 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_4_NAND3X1_75 BUFX2_35/A DFFSR_97/S FILL
XFILL_17_2_1 BUFX2_7/gnd DFFSR_54/S FILL
XOAI22X1_54 INVX1_366/Y OAI22X1_38/B INVX1_367/Y OAI22X1_38/D BUFX2_8/gnd NOR2X1_36/A
+ DFFSR_10/S OAI22X1
XFILL_5_OAI22X1_57 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_41_DFFSR_98 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_8_OAI21X1_254 INVX1_23/gnd DFFSR_91/S FILL
XFILL_3_NAND3X1_78 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_2_NAND2X1_151 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_4_OAI22X1_60 INVX1_8/gnd DFFSR_5/S FILL
XFILL_41_DFFSR_117 INVX1_23/gnd DFFSR_91/S FILL
XFILL_2_AND2X2_7 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_2_NAND3X1_81 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_3_OAI22X1_63 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_8_DFFSR_55 INVX1_89/gnd DFFSR_36/S FILL
XFILL_25_DFFSR_48 INVX1_4/gnd DFFSR_4/S FILL
XFILL_14_DFFSR_88 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_15_4_2 BUFX2_37/A DFFSR_81/S FILL
XFILL_1_NAND3X1_84 INVX1_94/gnd DFFSR_25/S FILL
XFILL_2_OAI22X1_66 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_31_DFFSR_120 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_21_DFFSR_123 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_0_OAI21X1_133 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_0_NAND3X1_87 INVX1_94/gnd DFFSR_52/S FILL
XFILL_9_OAI21X1_188 INVX1_89/gnd DFFSR_2/S FILL
XFILL_11_DFFSR_126 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_1_AOI21X1_5 BUFX2_37/A DFFSR_81/S FILL
XFILL_1_INVX1_277 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_22_DFFSR_95 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_33_DFFSR_55 INVX1_89/gnd DFFSR_36/S FILL
XINVX1_89 DFFSR_79/Q INVX1_89/gnd INVX1_89/Y DFFSR_2/S INVX1
XFILL_0_NAND2X1_247 INVX1_8/gnd DFFSR_5/S FILL
XFILL_44_DFFSR_15 INVX1_8/gnd DFFSR_7/S FILL
XFILL_7_DFFSR_120 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_9_NAND3X1_24 BUFX2_37/A DFFSR_8/S FILL
XFILL_48_DFFSR_151 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_0_DFFSR_12 BUFX2_6/gnd DFFSR_14/S FILL
XINVX1_207 AND2X2_8/B BUFX2_36/A INVX1_207/Y DFFSR_6/S INVX1
XFILL_38_DFFSR_154 BUFX2_36/A DFFSR_6/S FILL
XFILL_8_NAND3X1_27 BUFX2_37/A DFFSR_81/S FILL
XFILL_28_DFFSR_157 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_4_BUFX2_40 BUFX2_35/A DFFSR_14/S FILL
XFILL_7_NAND3X1_30 INVX1_94/gnd DFFSR_52/S FILL
XFILL_8_OAI22X1_12 INVX1_4/gnd DFFSR_51/S FILL
XFILL_4_DFFPOSX1_19 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_1_NAND2X1_181 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_6_NAND3X1_33 INVX1_8/gnd DFFSR_7/S FILL
XFILL_18_DFFSR_160 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_7_OAI22X1_15 INVX1_4/gnd DFFSR_4/S FILL
XFILL_5_NAND3X1_36 BUFX2_35/A DFFSR_97/S FILL
XFILL_41_DFFSR_6 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_3_NAND3X1_4 INVX1_94/gnd DFFSR_52/S FILL
XFILL_6_OAI22X1_18 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_4_NAND3X1_39 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_41_DFFSR_62 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_2_INVX1_96 DFFSR_79/gnd DFFSR_36/S FILL
XNAND3X1_33 INVX1_237/A AOI21X1_17/A AOI21X1_17/B INVX1_8/gnd NAND3X1_33/Y DFFSR_7/S
+ NAND3X1
XFILL_5_OAI22X1_21 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_3_NAND3X1_42 BUFX2_43/A DFFSR_23/S FILL
XFILL_2_NAND2X1_115 BUFX2_36/A DFFSR_6/S FILL
XOAI22X1_18 INVX1_291/Y OAI22X1_6/B INVX1_292/Y OAI22X1_8/D BUFX2_8/gnd NOR2X1_18/A
+ DFFSR_10/S OAI22X1
XFILL_4_OAI22X1_24 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_3_NOR2X1_39 INVX1_8/gnd DFFSR_5/S FILL
XDFFSR_160 DFFSR_160/Q CLKBUF1_10/Y DFFSR_162/R DFFSR_57/S DFFSR_160/D BUFX2_17/gnd
+ DFFSR_57/S DFFSR
XFILL_8_OAI21X1_218 INVX1_23/gnd DFFSR_186/S FILL
XFILL_2_NAND3X1_45 BUFX2_35/A DFFSR_97/S FILL
XFILL_3_OAI22X1_27 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_2_INVX1_421 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_8_DFFSR_19 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_4_DFFSR_157 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_25_DFFSR_12 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_1_NAND3X1_48 BUFX2_43/A DFFSR_23/S FILL
XFILL_14_DFFSR_52 INVX1_94/gnd DFFSR_52/S FILL
XFILL_2_OAI22X1_30 INVX1_94/gnd DFFSR_25/S FILL
XFILL_0_NAND3X1_51 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_1_OAI22X1_33 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_45_DFFSR_188 INVX1_2/gnd DFFSR_1/S FILL
XFILL_35_DFFSR_191 INVX1_23/gnd DFFSR_91/S FILL
XFILL_5_0_2 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_23_DFFPOSX1_27 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_0_OAI22X1_36 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_1_INVX1_241 BUFX2_43/A DFFSR_23/S FILL
XFILL_49_DFFSR_69 BUFX2_43/A DFFSR_23/S FILL
XFILL_0_NAND2X1_211 BUFX2_6/gnd DFFSR_91/S FILL
XINVX1_53 INVX1_53/A INVX1_89/gnd INVX1_53/Y DFFSR_2/S INVX1
XFILL_11_DFFSR_99 BUFX2_35/A DFFSR_97/S FILL
XFILL_33_DFFSR_19 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_5_DFFSR_66 INVX1_2/gnd DFFSR_51/S FILL
XFILL_22_DFFSR_59 INVX1_4/gnd DFFSR_51/S FILL
XFILL_48_DFFSR_115 BUFX2_6/gnd DFFSR_14/S FILL
XINVX1_171 BUFX2_5/Y BUFX2_35/A DFFSR_148/R DFFSR_14/S INVX1
XFILL_38_DFFSR_118 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_4_INVX1_168 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_1_NAND2X1_145 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_28_DFFSR_121 BUFX2_36/A DFFSR_6/S FILL
XFILL_7_OAI21X1_248 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_18_DFFSR_124 INVX1_89/gnd DFFSR_36/S FILL
XFILL_8_AOI21X1_3 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_2_INVX1_60 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_41_DFFSR_26 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_30_DFFSR_66 INVX1_2/gnd DFFSR_51/S FILL
XDFFSR_124 INVX1_362/A CLKBUF1_1/Y DFFSR_123/R DFFSR_36/S DFFSR_124/D INVX1_89/gnd
+ DFFSR_36/S DFFSR
XFILL_8_OAI21X1_182 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_4_DFFSR_121 BUFX2_36/A DFFSR_6/S FILL
XFILL_2_INVX1_385 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_14_DFFSR_16 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_29_1 INVX1_89/gnd DFFSR_36/S FILL
XFILL_45_DFFSR_152 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_1_NAND3X1_12 INVX1_94/gnd DFFSR_52/S FILL
XFILL_35_DFFSR_155 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_0_NAND3X1_15 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_8_DFFSR_9 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_25_DFFSR_158 BUFX2_43/A DFFSR_23/S FILL
XFILL_15_DFFSR_161 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_16_5_0 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_49_DFFSR_33 INVX1_94/gnd DFFSR_52/S FILL
XFILL_1_INVX1_205 INVX1_94/gnd DFFSR_25/S FILL
XFILL_38_DFFSR_73 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_0_NAND3X1_5 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_3_DFFPOSX1_13 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_0_NAND2X1_175 BUFX2_35/A DFFSR_14/S FILL
XFILL_22_DFFSR_23 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_11_DFFSR_63 INVX1_94/gnd DFFSR_52/S FILL
XFILL_5_DFFSR_30 INVX1_89/gnd DFFSR_36/S FILL
XINVX1_17 DFFSR_15/Q BUFX2_17/gnd INVX1_17/Y DFFSR_7/S INVX1
XDFFSR_70 DFFSR_70/Q CLKBUF1_3/Y DFFSR_68/R DFFSR_57/S DFFSR_70/D BUFX2_17/gnd DFFSR_57/S
+ DFFSR
XFILL_0_NOR2X1_40 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_8_NAND3X1_128 DFFSR_5/gnd DFFSR_5/S FILL
XINVX1_135 INVX1_390/A BUFX2_16/gnd INVX1_135/Y DFFSR_11/S INVX1
XFILL_1_DFFSR_158 BUFX2_43/A DFFSR_23/S FILL
XFILL_4_INVX1_132 BUFX2_35/A DFFSR_97/S FILL
XFILL_7_OAI21X1_212 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_1_NAND2X1_109 INVX1_94/gnd DFFSR_25/S FILL
XFILL_42_DFFSR_189 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_46_DFFSR_80 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_30_DFFSR_30 INVX1_89/gnd DFFSR_36/S FILL
XFILL_2_DFFSR_77 INVX1_89/gnd DFFSR_2/S FILL
XFILL_19_DFFSR_70 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_2_INVX1_24 INVX1_2/gnd DFFSR_51/S FILL
XFILL_22_DFFPOSX1_21 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_8_OAI21X1_146 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_2_INVX1_349 INVX1_89/gnd DFFSR_2/S FILL
XFILL_1_BUFX2_15 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_6_XOR2X1_7 INVX1_23/gnd DFFSR_91/S FILL
XFILL_45_DFFSR_116 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_35_DFFSR_119 BUFX2_37/A DFFSR_81/S FILL
XNOR3X1_1 NOR3X1_1/A NOR3X1_1/B NOR3X1_1/C INVX1_94/gnd NOR3X1_1/Y DFFSR_52/S NOR3X1
XFILL_26_0_0 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_1_INVX1_169 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_25_DFFSR_122 INVX1_94/gnd DFFSR_52/S FILL
XFILL_38_DFFSR_37 INVX1_89/gnd DFFSR_2/S FILL
XFILL_15_DFFSR_125 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_27_DFFSR_77 INVX1_89/gnd DFFSR_2/S FILL
XFILL_5_AOI21X1_4 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_24_2_1 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_0_NAND2X1_139 BUFX2_17/gnd DFFSR_57/S FILL
XDFFSR_34 INVX1_39/A DFFSR_24/CLK DFFSR_33/R DFFSR_9/S DFFSR_34/D DFFSR_1/gnd DFFSR_9/S
+ DFFSR
XFILL_6_1_0 BUFX2_35/A DFFSR_14/S FILL
XFILL_6_OAI21X1_242 BUFX2_35/A DFFSR_97/S FILL
XFILL_11_DFFSR_27 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_22_4_2 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_4_3_1 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_1_DFFSR_122 INVX1_94/gnd DFFSR_52/S FILL
XFILL_42_DFFSR_153 BUFX2_36/A DFFSR_8/S FILL
XFILL_7_OAI21X1_176 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_34_6 INVX1_8/gnd DFFSR_7/S FILL
XFILL_32_DFFSR_156 INVX1_23/gnd DFFSR_91/S FILL
XFILL_35_DFFSR_84 BUFX2_43/A DFFSR_23/S FILL
XFILL_46_DFFSR_44 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_2_5_2 INVX1_23/gnd DFFSR_186/S FILL
XFILL_22_DFFSR_159 BUFX2_36/A DFFSR_6/S FILL
XFILL_12_DFFSR_162 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_7_NAND3X1_3 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_2_DFFSR_41 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_19_DFFSR_34 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_2_INVX1_313 INVX1_8/gnd DFFSR_5/S FILL
XFILL_8_OAI21X1_110 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_12_XOR2X1_4 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_20_CLKBUF1_24 INVX1_23/gnd DFFSR_186/S FILL
XFILL_19_DFFSR_7 INVX1_8/gnd DFFSR_7/S FILL
XFILL_8_DFFSR_156 INVX1_23/gnd DFFSR_91/S FILL
XFILL_43_DFFSR_91 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_49_DFFSR_187 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_16_DFFSR_81 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_7_NAND3X1_122 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_27_DFFSR_41 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_39_DFFSR_190 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_1_INVX1_133 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_11_DFFPOSX1_26 BUFX2_37/A DFFSR_81/S FILL
XFILL_3_BUFX2_8 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_6_OAI21X1_206 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_0_NAND2X1_103 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_40_DFFSR_3 DFFSR_3/gnd DFFSR_4/S FILL
XOAI21X1_242 INVX1_401/Y AOI21X1_41/B INVX1_400/Y BUFX2_35/A AOI21X1_41/C DFFSR_97/S
+ OAI21X1
XFILL_42_DFFSR_117 INVX1_23/gnd DFFSR_91/S FILL
XFILL_21_DFFPOSX1_15 BUFX2_35/A DFFSR_14/S FILL
XFILL_7_OAI21X1_140 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_7_DFFSR_95 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_35_DFFSR_48 INVX1_4/gnd DFFSR_4/S FILL
XFILL_24_DFFSR_88 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_32_DFFSR_120 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_22_DFFSR_123 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_6_BUFX2_33 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_12_DFFSR_126 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_2_AOI21X1_5 BUFX2_37/A DFFSR_81/S FILL
XFILL_2_INVX1_277 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_32_DFFSR_95 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_43_DFFSR_55 INVX1_89/gnd DFFSR_36/S FILL
XFILL_4_INVX1_89 INVX1_89/gnd DFFSR_2/S FILL
XFILL_8_DFFSR_120 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_5_OAI21X1_236 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_49_DFFSR_151 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_39_DFFSR_154 BUFX2_36/A DFFSR_6/S FILL
XFILL_29_DFFSR_157 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_16_DFFSR_45 DFFSR_79/gnd DFFSR_45/S FILL
XNAND3X1_7 AOI22X1_3/C AOI22X1_3/D NAND3X1_7/C BUFX2_7/gnd NAND3X1_7/Y DFFSR_54/S
+ NAND3X1
XFILL_19_DFFSR_160 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_4_NAND3X1_4 INVX1_94/gnd DFFSR_52/S FILL
XFILL_6_OAI21X1_170 INVX1_94/gnd DFFSR_25/S FILL
XNOR2X1_42 NOR2X1_42/A NOR2X1_42/B BUFX2_17/gnd NOR2X1_42/Y DFFSR_57/S NOR2X1
XOAI21X1_206 AOI21X1_16/Y AOI21X1_15/Y AOI21X1_26/C BUFX2_5/gnd AOI21X1_27/B DFFSR_23/S
+ OAI21X1
XFILL_4_NOR2X1_39 INVX1_8/gnd DFFSR_5/S FILL
XFILL_12_CLKBUF1_12 BUFX2_43/A DFFSR_23/S FILL
XFILL_6_NAND2X1_284 INVX1_8/gnd DFFSR_5/S FILL
XFILL_3_INVX1_421 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_7_OAI21X1_104 INVX1_4/gnd DFFSR_51/S FILL
XFILL_13_DFFSR_92 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_5_DFFSR_157 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_35_DFFSR_12 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_24_DFFSR_52 INVX1_94/gnd DFFSR_52/S FILL
XFILL_11_CLKBUF1_15 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_7_DFFSR_59 INVX1_4/gnd DFFSR_51/S FILL
XFILL_10_CLKBUF1_18 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_23_5_0 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_46_DFFSR_188 INVX1_2/gnd DFFSR_1/S FILL
XFILL_36_DFFSR_191 INVX1_23/gnd DFFSR_91/S FILL
XFILL_2_INVX1_241 BUFX2_43/A DFFSR_23/S FILL
XFILL_7_DFFSR_6 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_9_CLKBUF1_21 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_8_CLKBUF1_24 INVX1_23/gnd DFFSR_186/S FILL
XFILL_10_DFFPOSX1_20 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_6_NAND3X1_116 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_21_DFFSR_99 BUFX2_35/A DFFSR_97/S FILL
XFILL_5_OAI21X1_200 BUFX2_37/A DFFSR_8/S FILL
XFILL_4_INVX1_53 INVX1_89/gnd DFFSR_2/S FILL
XFILL_43_DFFSR_19 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_32_DFFSR_59 INVX1_4/gnd DFFSR_51/S FILL
XFILL_49_DFFSR_115 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_39_DFFSR_118 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_29_DFFSR_121 BUFX2_36/A DFFSR_6/S FILL
XFILL_6_OAI21X1_134 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_19_DFFSR_124 INVX1_89/gnd DFFSR_36/S FILL
XFILL_9_AOI21X1_3 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_51_DFFSR_26 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_40_DFFSR_66 INVX1_2/gnd DFFSR_51/S FILL
XFILL_16_3 BUFX2_37/A DFFSR_81/S FILL
XOAI21X1_170 DFFSR_25/S INVX1_205/Y OAI21X1_170/C INVX1_94/gnd DFFSR_170/D DFFSR_25/S
+ OAI21X1
XFILL_6_NAND2X1_248 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_0_DFFPOSX1_31 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_7_DFFSR_23 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_5_DFFSR_121 BUFX2_36/A DFFSR_6/S FILL
XFILL_3_INVX1_385 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_24_DFFSR_16 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_33_0_0 INVX1_8/gnd DFFSR_7/S FILL
XFILL_13_DFFSR_56 INVX1_2/gnd DFFSR_51/S FILL
XFILL_46_DFFSR_152 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_36_DFFSR_155 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_31_2_1 DFFSR_5/gnd DFFSR_5/S FILL
XNAND2X1_284 NAND3X1_133/Y OAI21X1_263/Y INVX1_8/gnd NAND2X1_284/Y DFFSR_5/S NAND2X1
XFILL_4_OAI21X1_230 INVX1_23/gnd DFFSR_186/S FILL
XFILL_26_DFFSR_158 BUFX2_43/A DFFSR_23/S FILL
XFILL_6_NOR2X1_4 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_16_DFFSR_161 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_2_INVX1_205 INVX1_94/gnd DFFSR_25/S FILL
XFILL_29_4_2 INVX1_89/gnd DFFSR_2/S FILL
XFILL_48_DFFSR_73 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_1_NAND3X1_5 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_32_DFFSR_23 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_21_DFFSR_63 INVX1_94/gnd DFFSR_52/S FILL
XFILL_4_DFFSR_70 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_1_NOR2X1_40 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_5_OAI21X1_164 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_0_INVX1_422 INVX1_23/gnd DFFSR_186/S FILL
XFILL_9_5_2 BUFX2_43/A DFFSR_23/S FILL
XNAND3X1_116 NOR2X1_2/A INVX1_266/Y INVX1_264/Y DFFSR_71/gnd OAI22X1_7/D DFFSR_45/S
+ NAND3X1
XFILL_2_DFFSR_158 BUFX2_43/A DFFSR_23/S FILL
XFILL_5_NAND2X1_278 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_43_DFFSR_189 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_1_INVX1_64 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_40_DFFSR_30 INVX1_89/gnd DFFSR_36/S FILL
XFILL_29_DFFSR_70 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_0_CLKBUF1_12 BUFX2_43/A DFFSR_23/S FILL
XOAI21X1_134 DFFSR_45/S INVX1_151/Y OAI21X1_134/C DFFSR_79/gnd DFFSR_134/D DFFSR_36/S
+ OAI21X1
XFILL_6_NAND2X1_212 INVX1_23/gnd DFFSR_186/S FILL
XFILL_3_INVX1_349 INVX1_89/gnd DFFSR_2/S FILL
XFILL_3_OAI21X1_260 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_13_DFFSR_20 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_5_NAND3X1_110 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_46_DFFSR_116 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_36_DFFSR_119 BUFX2_37/A DFFSR_81/S FILL
XFILL_4_OAI21X1_194 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_4_NOR3X1_1 INVX1_94/gnd DFFSR_52/S FILL
XNAND2X1_248 NOR2X1_41/Y NOR2X1_40/Y BUFX2_8/gnd NAND2X1_248/Y DFFSR_10/S NAND2X1
XFILL_2_INVX1_169 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_26_DFFSR_122 INVX1_94/gnd DFFSR_52/S FILL
XFILL_18_DFFSR_4 INVX1_4/gnd DFFSR_4/S FILL
XFILL_16_DFFSR_125 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_48_DFFSR_37 INVX1_89/gnd DFFSR_2/S FILL
XFILL_37_DFFSR_77 INVX1_89/gnd DFFSR_2/S FILL
XFILL_6_AOI21X1_4 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_2_BUFX2_5 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_5_OAI21X1_128 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_21_DFFSR_27 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_4_DFFSR_34 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_10_DFFSR_67 INVX1_2/gnd DFFSR_51/S FILL
XFILL_21_8 INVX1_94/gnd DFFSR_52/S FILL
XFILL_0_INVX1_386 INVX1_94/gnd DFFSR_52/S FILL
XFILL_2_DFFSR_122 INVX1_94/gnd DFFSR_52/S FILL
XFILL_43_DFFSR_153 BUFX2_36/A DFFSR_8/S FILL
XFILL_38_3 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_33_DFFSR_156 INVX1_23/gnd DFFSR_91/S FILL
XFILL_45_DFFSR_84 BUFX2_43/A DFFSR_23/S FILL
XFILL_5_NAND2X1_242 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_23_DFFSR_159 BUFX2_36/A DFFSR_6/S FILL
XFILL_13_DFFSR_162 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_1_DFFSR_81 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_8_NAND3X1_3 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_1_INVX1_28 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_29_DFFSR_34 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_18_DFFSR_74 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_3_OAI21X1_224 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_9_DFFPOSX1_14 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_6_NAND2X1_176 INVX1_94/gnd DFFSR_25/S FILL
XFILL_23_DFFPOSX1_3 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_3_INVX1_313 INVX1_8/gnd DFFSR_5/S FILL
XFILL_22_DFFPOSX1_6 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_21_DFFPOSX1_9 BUFX2_37/A DFFSR_8/S FILL
XFILL_0_BUFX2_19 BUFX2_19/gnd DFFSR_54/S FILL
XNAND2X1_212 NOR2X1_7/Y XOR2X1_4/Y INVX1_23/gnd AOI22X1_13/A DFFSR_186/S NAND2X1
XFILL_9_DFFSR_156 INVX1_23/gnd DFFSR_91/S FILL
XFILL_4_OAI21X1_158 BUFX2_43/A DFFSR_97/S FILL
XFILL_50_DFFSR_187 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_26_DFFSR_81 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_37_DFFSR_41 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_40_DFFSR_190 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_9_DFFSR_88 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_2_INVX1_133 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_10_DFFSR_31 BUFX2_35/A DFFSR_97/S FILL
XFILL_4_NAND2X1_272 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_0_INVX1_350 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_30_5_0 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_2_OAI21X1_254 INVX1_23/gnd DFFSR_91/S FILL
XFILL_43_DFFSR_117 INVX1_23/gnd DFFSR_91/S FILL
XFILL_5_NAND2X1_206 BUFX2_43/A DFFSR_97/S FILL
XFILL_45_DFFSR_48 INVX1_4/gnd DFFSR_4/S FILL
XFILL_34_DFFSR_88 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_33_DFFSR_120 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_23_DFFSR_123 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_4_NAND3X1_104 INVX1_23/gnd DFFSR_186/S FILL
XFILL_1_DFFSR_45 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_13_DFFSR_126 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_18_DFFSR_38 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_3_AOI21X1_5 BUFX2_37/A DFFSR_81/S FILL
XFILL_6_NAND2X1_140 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_3_OAI21X1_188 INVX1_89/gnd DFFSR_2/S FILL
XFILL_3_INVX1_277 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_6_DFFSR_3 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_11_XOR2X1_8 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_42_DFFSR_95 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_9_DFFSR_120 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_50_DFFSR_151 BUFX2_7/gnd DFFSR_81/S FILL
XNAND2X1_176 BUFX2_12/Y AND2X2_11/A INVX1_94/gnd NOR2X1_4/A DFFSR_25/S NAND2X1
XFILL_4_OAI21X1_122 INVX1_94/gnd DFFSR_25/S FILL
XFILL_40_DFFSR_154 BUFX2_36/A DFFSR_6/S FILL
XFILL_3_AND2X2_4 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_30_DFFSR_157 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_9_DFFSR_52 INVX1_94/gnd DFFSR_52/S FILL
XFILL_15_DFFSR_85 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_26_DFFSR_45 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_43_8 INVX1_4/gnd DFFSR_4/S FILL
XFILL_20_DFFSR_160 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_4_OR2X2_3 BUFX2_43/A DFFSR_23/S FILL
XFILL_5_NAND3X1_4 INVX1_94/gnd DFFSR_52/S FILL
XFILL_4_NAND2X1_236 INVX1_2/gnd DFFSR_1/S FILL
XFILL_40_0_0 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_10_DFFSR_163 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_3_NAND3X1_134 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_0_INVX1_314 INVX1_8/gnd DFFSR_5/S FILL
XFILL_5_NOR2X1_39 INVX1_8/gnd DFFSR_5/S FILL
XFILL_30_DFFSR_7 INVX1_8/gnd DFFSR_7/S FILL
XINVX1_424 INVX1_424/A BUFX2_16/gnd INVX1_424/Y DFFSR_65/S INVX1
XFILL_38_2_1 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_2_OAI21X1_218 INVX1_23/gnd DFFSR_186/S FILL
XFILL_4_INVX1_421 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_23_DFFSR_92 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_6_DFFSR_157 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_45_DFFSR_12 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_6_DFFSR_99 BUFX2_35/A DFFSR_97/S FILL
XFILL_34_DFFSR_52 INVX1_94/gnd DFFSR_52/S FILL
XFILL_36_4_2 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_5_NAND2X1_170 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_47_DFFSR_188 INVX1_2/gnd DFFSR_1/S FILL
XFILL_37_DFFSR_191 INVX1_23/gnd DFFSR_91/S FILL
XFILL_11_DFFPOSX1_3 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_3_INVX1_241 BUFX2_43/A DFFSR_23/S FILL
XFILL_3_OAI21X1_152 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_5_BUFX2_37 BUFX2_37/A DFFSR_81/S FILL
XFILL_17_DFFPOSX1_27 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_6_NAND2X1_104 INVX1_4/gnd DFFSR_51/S FILL
XFILL_10_DFFPOSX1_6 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_9_DFFPOSX1_9 BUFX2_37/A DFFSR_8/S FILL
XFILL_31_DFFSR_99 BUFX2_35/A DFFSR_97/S FILL
XNAND2X1_140 DFFSR_10/S NAND2X1_245/Y DFFSR_71/gnd NAND2X1_140/Y DFFSR_10/S NAND2X1
XFILL_3_INVX1_93 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_42_DFFSR_59 INVX1_4/gnd DFFSR_51/S FILL
XFILL_27_DFFPOSX1_16 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_50_DFFSR_115 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_8_AOI21X1_32 BUFX2_43/A DFFSR_23/S FILL
XFILL_3_NAND2X1_266 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_7_AOI21X1_35 INVX1_94/gnd DFFSR_25/S FILL
XFILL_9_DFFSR_16 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_40_DFFSR_118 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_15_DFFSR_49 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_30_DFFSR_121 BUFX2_36/A DFFSR_6/S FILL
XFILL_6_AOI21X1_38 BUFX2_36/A DFFSR_8/S FILL
XFILL_4_NAND2X1_200 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_5_AOI21X1_41 BUFX2_35/A DFFSR_14/S FILL
XFILL_20_DFFSR_124 INVX1_89/gnd DFFSR_36/S FILL
XFILL_1_OAI21X1_248 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_10_DFFSR_127 BUFX2_43/A DFFSR_97/S FILL
XAOI21X1_38 OR2X2_3/Y AOI21X1_38/B INVX1_251/Y BUFX2_36/A OAI22X1_4/A DFFSR_8/S AOI21X1
XFILL_4_AOI21X1_44 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_3_AOI21X1_47 BUFX2_43/A DFFSR_23/S FILL
XFILL_0_AOI21X1_6 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_50_DFFSR_66 INVX1_2/gnd DFFSR_51/S FILL
XFILL_0_INVX1_278 DFFSR_3/gnd DFFSR_4/S FILL
XINVX1_388 DFFSR_88/Q DFFSR_3/gnd INVX1_388/Y DFFSR_65/S INVX1
XFILL_6_DFFSR_121 BUFX2_36/A DFFSR_6/S FILL
XFILL_6_DFFSR_63 INVX1_94/gnd DFFSR_52/S FILL
XFILL_34_DFFSR_16 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_5_NAND2X1_134 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_2_OAI21X1_182 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_12_DFFSR_96 INVX1_2/gnd DFFSR_1/S FILL
XFILL_23_DFFSR_56 INVX1_2/gnd DFFSR_51/S FILL
XFILL_47_DFFSR_152 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_37_DFFSR_155 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_27_DFFSR_158 BUFX2_43/A DFFSR_23/S FILL
XBUFX2_41 BUFX2_36/A BUFX2_37/A BUFX2_41/Y DFFSR_81/S BUFX2
XFILL_17_DFFSR_161 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_3_INVX1_205 INVX1_94/gnd DFFSR_25/S FILL
XFILL_3_OAI21X1_116 INVX1_89/gnd DFFSR_2/S FILL
XFILL_2_NAND3X1_5 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_17_DFFSR_1 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_8_OAI21X1_80 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_42_DFFSR_23 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_31_DFFSR_63 INVX1_94/gnd DFFSR_52/S FILL
XFILL_7_OAI21X1_83 INVX1_94/gnd DFFSR_52/S FILL
XFILL_3_INVX1_57 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_3_NAND2X1_230 BUFX2_36/A DFFSR_6/S FILL
XFILL_2_NOR2X1_40 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_6_OAI21X1_86 INVX1_4/gnd DFFSR_51/S FILL
XNAND2X1_104 BUFX2_15/Y DFFSR_96/Q INVX1_4/gnd NAND2X1_104/Y DFFSR_51/S NAND2X1
XFILL_1_INVX1_422 INVX1_23/gnd DFFSR_186/S FILL
XFILL_5_OAI21X1_89 BUFX2_35/A DFFSR_14/S FILL
XFILL_1_BUFX2_2 BUFX2_43/A DFFSR_23/S FILL
XFILL_12_0_1 BUFX2_36/A DFFSR_6/S FILL
XFILL_3_DFFSR_158 BUFX2_43/A DFFSR_23/S FILL
XFILL_4_OAI21X1_92 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_2_NAND3X1_128 DFFSR_5/gnd DFFSR_5/S FILL
XOAI21X1_86 BUFX2_15/Y INVX1_97/Y NAND2X1_86/Y INVX1_4/gnd DFFSR_86/D DFFSR_51/S OAI21X1
XFILL_15_DFFSR_13 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_1_OAI21X1_212 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_10_2_2 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_3_OAI21X1_95 INVX1_89/gnd DFFSR_36/S FILL
XFILL_44_DFFSR_189 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_4_NAND2X1_164 INVX1_8/gnd DFFSR_5/S FILL
XFILL_2_OAI21X1_98 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_50_DFFSR_30 INVX1_89/gnd DFFSR_36/S FILL
XINVX1_352 DFFSR_99/Q BUFX2_5/gnd INVX1_352/Y DFFSR_6/S INVX1
XFILL_0_INVX1_242 BUFX2_36/A DFFSR_6/S FILL
XFILL_3_AOI21X1_11 INVX1_8/gnd DFFSR_5/S FILL
XFILL_39_DFFSR_70 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_2_OAI21X1_146 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_16_DFFPOSX1_21 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_2_AOI21X1_14 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_23_DFFSR_20 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_12_DFFSR_60 BUFX2_37/A DFFSR_8/S FILL
XFILL_1_AOI21X1_17 INVX1_8/gnd DFFSR_5/S FILL
XFILL_6_DFFSR_27 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_0_AOI21X1_20 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_47_DFFSR_116 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_5_NOR2X1_8 BUFX2_43/A DFFSR_23/S FILL
XFILL_37_DFFSR_119 BUFX2_37/A DFFSR_81/S FILL
XFILL_3_INVX1_169 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_2_NAND2X1_260 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_27_DFFSR_122 INVX1_94/gnd DFFSR_52/S FILL
XFILL_26_DFFPOSX1_10 INVX1_8/gnd DFFSR_5/S FILL
XFILL_17_DFFSR_125 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_8_OAI21X1_44 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_47_DFFSR_77 INVX1_89/gnd DFFSR_2/S FILL
XFILL_37_5_0 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_7_AOI21X1_4 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_7_OAI21X1_47 INVX1_89/gnd DFFSR_2/S FILL
XFILL_6_NAND2X1_65 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_0_OAI21X1_242 BUFX2_35/A DFFSR_97/S FILL
XFILL_3_NAND2X1_194 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_5_NAND2X1_68 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_6_OAI21X1_50 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_31_DFFSR_27 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_3_INVX1_21 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_3_DFFSR_74 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_20_DFFSR_67 INVX1_2/gnd DFFSR_51/S FILL
XFILL_4_NAND2X1_71 BUFX2_8/gnd DFFSR_10/S FILL
XNAND2X1_65 NAND2X1_65/A BUFX2_24/Y DFFSR_3/gnd OAI21X1_65/C DFFSR_4/S NAND2X1
XFILL_1_INVX1_386 INVX1_94/gnd DFFSR_52/S FILL
XFILL_3_DFFSR_122 INVX1_94/gnd DFFSR_52/S FILL
XFILL_25_5 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_5_OAI21X1_53 DFFSR_71/gnd DFFSR_45/S FILL
XOAI21X1_50 DFFSR_15/S INVX1_57/Y NAND2X1_50/Y BUFX2_17/gnd DFFSR_50/D DFFSR_7/S OAI21X1
XFILL_7_XOR2X1_4 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_44_DFFSR_153 BUFX2_36/A DFFSR_8/S FILL
XFILL_2_BUFX2_12 BUFX2_37/A DFFSR_81/S FILL
XFILL_3_NAND2X1_74 INVX1_2/gnd DFFSR_1/S FILL
XFILL_4_OAI21X1_56 INVX1_2/gnd DFFSR_51/S FILL
XFILL_34_DFFSR_156 INVX1_23/gnd DFFSR_91/S FILL
XFILL_1_OAI21X1_176 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_2_NAND2X1_77 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_4_NAND2X1_128 INVX1_89/gnd DFFSR_2/S FILL
XFILL_3_OAI21X1_59 INVX1_4/gnd DFFSR_51/S FILL
XFILL_24_DFFSR_159 BUFX2_36/A DFFSR_6/S FILL
XFILL_2_OAI21X1_62 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_1_NAND2X1_80 BUFX2_17/gnd DFFSR_57/S FILL
XINVX1_316 INVX1_26/A BUFX2_37/A INVX1_316/Y DFFSR_8/S INVX1
XFILL_0_INVX1_68 BUFX2_37/A DFFSR_81/S FILL
XFILL_0_INVX1_206 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_0_NAND2X1_83 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_39_DFFSR_34 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_28_DFFSR_74 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_1_OAI21X1_65 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_14_DFFSR_162 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_0_OAI21X1_68 BUFX2_37/A DFFSR_81/S FILL
XFILL_4_INVX1_313 INVX1_8/gnd DFFSR_5/S FILL
XFILL_12_DFFSR_24 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_2_OAI21X1_110 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_0_DFFSR_159 BUFX2_36/A DFFSR_6/S FILL
XFILL_2_NAND2X1_224 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_47_0_0 DFFSR_1/gnd DFFSR_9/S FILL
XDFFSR_4 DFFSR_4/Q DFFSR_3/CLK DFFSR_6/R DFFSR_4/S DFFSR_4/D INVX1_4/gnd DFFSR_4/S
+ DFFSR
XFILL_36_DFFSR_81 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_47_DFFSR_41 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_41_DFFSR_190 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_3_INVX1_133 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_1_NAND3X1_122 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_45_2_1 INVX1_2/gnd DFFSR_1/S FILL
XFILL_20_DFFSR_31 BUFX2_35/A DFFSR_97/S FILL
XFILL_3_DFFSR_38 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_6_NAND2X1_29 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_7_OAI21X1_11 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_3_NAND2X1_158 BUFX2_35/A DFFSR_97/S FILL
XFILL_6_OAI21X1_14 BUFX2_43/A DFFSR_23/S FILL
XFILL_0_OAI21X1_206 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_5_NAND2X1_32 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_1_INVX1_350 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_5_OAI21X1_17 INVX1_8/gnd DFFSR_5/S FILL
XFILL_4_NAND2X1_35 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_43_4_2 INVX1_4/gnd DFFSR_51/S FILL
XNAND2X1_29 DFFSR_4/S INVX1_24/A DFFSR_3/gnd OAI21X1_29/C DFFSR_4/S NAND2X1
XFILL_4_OAI21X1_20 DFFSR_89/gnd DFFSR_186/S FILL
XOAI21X1_14 DFFSR_23/S INVX1_16/Y OAI21X1_14/C BUFX2_43/A DFFSR_14/D DFFSR_23/S OAI21X1
XFILL_3_NAND2X1_38 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_44_DFFSR_117 INVX1_23/gnd DFFSR_91/S FILL
XFILL_15_DFFPOSX1_15 BUFX2_35/A DFFSR_14/S FILL
XFILL_3_OAI21X1_23 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_1_OAI21X1_140 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_13_XOR2X1_1 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_2_NAND2X1_41 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_29_DFFSR_4 INVX1_4/gnd DFFSR_4/S FILL
XFILL_44_DFFSR_88 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_9_NAND3X1_97 BUFX2_35/A DFFSR_97/S FILL
XFILL_1_NAND2X1_44 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_2_OAI21X1_26 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_34_DFFSR_120 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_24_DFFSR_123 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_0_INVX1_32 BUFX2_7/gnd DFFSR_54/S FILL
XAOI21X1_8 AOI21X1_8/A AOI21X1_8/B AOI21X1_2/Y INVX1_94/gnd AOI21X1_8/Y DFFSR_52/S
+ AOI21X1
XFILL_0_NAND2X1_47 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_1_OAI21X1_29 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_0_INVX1_170 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_0_DFFSR_85 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_14_DFFSR_126 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_28_DFFSR_38 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_17_DFFSR_78 DFFSR_1/gnd DFFSR_1/S FILL
XINVX1_280 INVX1_30/A INVX1_2/gnd INVX1_280/Y DFFSR_51/S INVX1
XFILL_0_OAI21X1_32 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_11_3_0 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_4_AOI21X1_5 BUFX2_37/A DFFSR_81/S FILL
XFILL_1_NAND2X1_254 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_5_DFFPOSX1_26 BUFX2_37/A DFFSR_81/S FILL
XFILL_0_DFFSR_123 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_41_DFFSR_154 BUFX2_36/A DFFSR_6/S FILL
XFILL_2_NAND2X1_188 INVX1_8/gnd DFFSR_7/S FILL
XFILL_8_DFFSR_92 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_5_AOI22X1_10 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_31_DFFSR_157 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_25_DFFSR_85 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_36_DFFSR_45 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_4_AOI22X1_13 INVX1_23/gnd DFFSR_186/S FILL
XFILL_21_DFFSR_160 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_6_NAND3X1_4 INVX1_94/gnd DFFSR_52/S FILL
XFILL_0_OAI21X1_170 INVX1_94/gnd DFFSR_25/S FILL
XFILL_3_NAND2X1_122 INVX1_94/gnd DFFSR_25/S FILL
XINVX1_6 DFFSR_5/Q INVX1_8/gnd INVX1_6/Y DFFSR_5/S INVX1
XFILL_11_DFFSR_163 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_11_OAI22X1_40 BUFX2_37/A DFFSR_8/S FILL
XFILL_1_INVX1_314 INVX1_8/gnd DFFSR_5/S FILL
XFILL_6_NOR2X1_39 INVX1_8/gnd DFFSR_5/S FILL
XFILL_10_OAI22X1_43 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_33_DFFSR_92 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_7_DFFSR_157 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_44_DFFSR_52 INVX1_94/gnd DFFSR_52/S FILL
XFILL_0_NAND2X1_284 INVX1_8/gnd DFFSR_5/S FILL
XFILL_1_OAI21X1_104 INVX1_4/gnd DFFSR_51/S FILL
XAND2X2_1 AND2X2_1/A AND2X2_1/B BUFX2_5/gnd AND2X2_1/Y DFFSR_23/S AND2X2
XFILL_48_DFFSR_188 INVX1_2/gnd DFFSR_1/S FILL
XFILL_38_DFFSR_191 INVX1_23/gnd DFFSR_91/S FILL
XFILL_8_NAND3X1_64 BUFX2_35/A DFFSR_14/S FILL
XFILL_0_INVX1_134 BUFX2_37/A DFFSR_8/S FILL
XFILL_9_OAI22X1_46 BUFX2_19/gnd DFFSR_52/S FILL
XINVX1_244 INVX1_244/A DFFSR_71/gnd INVX1_244/Y DFFSR_45/S INVX1
XFILL_17_DFFSR_42 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_0_NAND2X1_11 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_0_DFFSR_49 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_7_NAND3X1_67 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_8_OAI22X1_49 INVX1_94/gnd DFFSR_25/S FILL
XFILL_1_NAND2X1_218 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_6_NAND3X1_70 BUFX2_35/A DFFSR_14/S FILL
XFILL_19_0_1 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_7_OAI22X1_52 INVX1_94/gnd DFFSR_25/S FILL
XNAND3X1_70 NAND3X1_70/A INVX1_245/Y NAND3X1_70/C BUFX2_35/A NAND3X1_70/Y DFFSR_14/S
+ NAND3X1
XFILL_5_NAND3X1_73 BUFX2_43/A DFFSR_23/S FILL
XFILL_0_NAND3X1_116 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_6_OAI22X1_55 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_41_DFFSR_99 BUFX2_35/A DFFSR_97/S FILL
XFILL_4_NAND3X1_76 BUFX2_5/gnd DFFSR_6/S FILL
XOAI22X1_55 INVX1_369/Y OAI22X1_39/B INVX1_368/Y OAI22X1_39/D DFFSR_79/gnd NOR2X1_37/B
+ DFFSR_36/S OAI22X1
XFILL_5_OAI22X1_58 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_51_DFFSR_115 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_2_NAND2X1_152 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_3_NAND3X1_79 BUFX2_36/A DFFSR_6/S FILL
XFILL_17_2_2 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_4_OAI22X1_61 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_8_OAI21X1_255 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_14_DFFSR_89 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_2_AND2X2_8 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_2_NAND3X1_82 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_3_OAI22X1_64 INVX1_94/gnd DFFSR_25/S FILL
XFILL_8_DFFSR_56 INVX1_2/gnd DFFSR_51/S FILL
XFILL_41_DFFSR_118 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_25_DFFSR_49 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_31_DFFSR_121 BUFX2_36/A DFFSR_6/S FILL
XFILL_1_NAND3X1_85 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_2_OAI22X1_67 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_0_NAND3X1_88 INVX1_94/gnd DFFSR_52/S FILL
XFILL_21_DFFSR_124 INVX1_89/gnd DFFSR_36/S FILL
XFILL_11_DFFSR_127 BUFX2_43/A DFFSR_97/S FILL
XFILL_0_OAI21X1_134 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_9_OAI21X1_189 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_1_AOI21X1_6 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_1_INVX1_278 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_7_DFFSR_121 BUFX2_36/A DFFSR_6/S FILL
XFILL_0_NAND2X1_248 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_44_DFFSR_16 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_22_DFFSR_96 INVX1_2/gnd DFFSR_1/S FILL
XFILL_33_DFFSR_56 INVX1_2/gnd DFFSR_51/S FILL
XINVX1_90 INVX1_90/A DFFSR_73/gnd INVX1_90/Y DFFSR_11/S INVX1
XFILL_48_DFFSR_152 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_44_5_0 INVX1_2/gnd DFFSR_51/S FILL
XFILL_8_NAND3X1_28 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_38_DFFSR_155 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_9_OAI22X1_10 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_0_DFFSR_13 BUFX2_16/gnd DFFSR_65/S FILL
XINVX1_208 INVX1_246/A INVX1_23/gnd INVX1_208/Y DFFSR_186/S INVX1
XFILL_28_DFFSR_158 BUFX2_43/A DFFSR_23/S FILL
XFILL_4_BUFX2_41 BUFX2_37/A DFFSR_81/S FILL
XFILL_4_DFFPOSX1_20 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_7_NAND3X1_31 INVX1_94/gnd DFFSR_52/S FILL
XFILL_8_OAI22X1_13 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_1_NAND2X1_182 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_6_NAND3X1_34 INVX1_2/gnd DFFSR_1/S FILL
XFILL_7_OAI22X1_16 INVX1_4/gnd DFFSR_4/S FILL
XFILL_18_DFFSR_161 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_5_NAND3X1_37 BUFX2_43/A DFFSR_97/S FILL
XFILL_3_NAND3X1_5 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_6_OAI22X1_19 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_41_DFFSR_7 INVX1_8/gnd DFFSR_7/S FILL
XFILL_4_NAND3X1_40 BUFX2_43/A DFFSR_23/S FILL
XFILL_41_DFFSR_63 INVX1_94/gnd DFFSR_52/S FILL
XNAND3X1_34 NAND3X1_2/A NAND3X1_33/Y NAND3X1_34/C INVX1_2/gnd NAND3X1_34/Y DFFSR_1/S
+ NAND3X1
XFILL_2_INVX1_97 INVX1_4/gnd DFFSR_4/S FILL
XFILL_5_OAI22X1_22 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_3_NAND3X1_43 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_4_OAI22X1_25 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_3_NOR2X1_40 BUFX2_8/gnd DFFSR_10/S FILL
XOAI22X1_19 INVX1_294/Y OAI22X1_7/B INVX1_293/Y OAI22X1_7/D DFFSR_71/gnd NOR2X1_19/A
+ DFFSR_45/S OAI22X1
XDFFSR_161 DFFSR_161/Q CLKBUF1_14/Y DFFSR_162/R DFFSR_186/S DFFSR_161/D DFFSR_89/gnd
+ DFFSR_186/S DFFSR
XFILL_2_INVX1_422 INVX1_23/gnd DFFSR_186/S FILL
XFILL_2_NAND3X1_46 BUFX2_35/A DFFSR_97/S FILL
XFILL_8_OAI21X1_219 BUFX2_35/A DFFSR_97/S FILL
XFILL_3_OAI22X1_28 INVX1_94/gnd DFFSR_25/S FILL
XFILL_2_NAND2X1_116 INVX1_89/gnd DFFSR_36/S FILL
XFILL_8_DFFSR_20 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_4_DFFSR_158 BUFX2_43/A DFFSR_23/S FILL
XFILL_1_NAND3X1_49 BUFX2_37/A DFFSR_8/S FILL
XFILL_14_DFFSR_53 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_25_DFFSR_13 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_2_OAI22X1_31 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_45_DFFSR_189 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_0_NAND3X1_52 BUFX2_36/A DFFSR_8/S FILL
XFILL_23_DFFPOSX1_28 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_1_OAI22X1_34 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_0_OAI22X1_37 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_7_1 BUFX2_35/A DFFSR_14/S FILL
XFILL_1_INVX1_242 BUFX2_36/A DFFSR_6/S FILL
XFILL_49_DFFSR_70 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_33_DFFSR_20 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_0_NAND2X1_212 INVX1_23/gnd DFFSR_186/S FILL
XFILL_22_DFFSR_60 BUFX2_37/A DFFSR_8/S FILL
XFILL_5_DFFSR_67 INVX1_2/gnd DFFSR_51/S FILL
XINVX1_54 INVX1_54/A DFFSR_3/gnd INVX1_54/Y DFFSR_4/S INVX1
XFILL_48_DFFSR_116 DFFSR_5/gnd DFFSR_2/S FILL
XINVX1_172 INVX1_172/A DFFSR_89/gnd INVX1_172/Y DFFSR_186/S INVX1
XFILL_38_DFFSR_119 BUFX2_37/A DFFSR_81/S FILL
XFILL_1_NAND2X1_146 INVX1_23/gnd DFFSR_91/S FILL
XFILL_28_DFFSR_122 INVX1_94/gnd DFFSR_52/S FILL
XFILL_4_INVX1_169 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_7_OAI21X1_249 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_18_DFFSR_125 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_8_AOI21X1_4 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_2_INVX1_61 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_41_DFFSR_27 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_30_DFFSR_67 INVX1_2/gnd DFFSR_51/S FILL
XDFFSR_125 DFFSR_125/Q CLKBUF1_7/Y DFFSR_123/R DFFSR_91/S DFFSR_125/D BUFX2_6/gnd
+ DFFSR_91/S DFFSR
XFILL_8_OAI21X1_183 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_2_NAND3X1_10 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_2_INVX1_386 INVX1_94/gnd DFFSR_52/S FILL
XFILL_29_2 INVX1_89/gnd DFFSR_36/S FILL
XFILL_14_DFFSR_17 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_45_DFFSR_153 BUFX2_36/A DFFSR_8/S FILL
XFILL_4_DFFSR_122 INVX1_94/gnd DFFSR_52/S FILL
XFILL_1_NAND3X1_13 INVX1_94/gnd DFFSR_25/S FILL
XFILL_35_DFFSR_156 INVX1_23/gnd DFFSR_91/S FILL
XFILL_18_3_0 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_0_NAND3X1_16 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_25_DFFSR_159 BUFX2_36/A DFFSR_6/S FILL
XFILL_28_DFFSR_1 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_1_INVX1_206 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_49_DFFSR_34 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_38_DFFSR_74 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_15_DFFSR_162 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_16_5_1 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_0_NAND3X1_6 INVX1_8/gnd DFFSR_7/S FILL
XFILL_3_DFFPOSX1_14 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_5_DFFSR_31 BUFX2_35/A DFFSR_97/S FILL
XFILL_0_NAND2X1_176 INVX1_94/gnd DFFSR_25/S FILL
XDFFSR_71 INVX1_80/A CLKBUF1_1/Y DFFSR_68/R DFFSR_10/S DFFSR_71/D DFFSR_71/gnd DFFSR_10/S
+ DFFSR
XINVX1_18 DFFSR_16/Q INVX1_89/gnd INVX1_18/Y DFFSR_2/S INVX1
XFILL_22_DFFSR_24 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_11_DFFSR_64 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_0_NOR2X1_41 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_8_NAND3X1_129 BUFX2_35/A DFFSR_14/S FILL
XINVX1_136 BUFX2_5/Y BUFX2_43/A DFFSR_113/R DFFSR_97/S INVX1
XFILL_1_DFFSR_159 BUFX2_36/A DFFSR_6/S FILL
XFILL_7_OAI21X1_213 BUFX2_36/A DFFSR_6/S FILL
XFILL_46_DFFSR_81 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_42_DFFSR_190 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_4_INVX1_133 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_1_NAND2X1_110 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_2_INVX1_25 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_2_DFFSR_78 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_30_DFFSR_31 BUFX2_35/A DFFSR_97/S FILL
XFILL_19_DFFSR_71 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_8_OAI21X1_147 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_2_INVX1_350 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_22_DFFPOSX1_22 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_1_BUFX2_16 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_45_DFFSR_117 INVX1_23/gnd DFFSR_91/S FILL
XFILL_6_XOR2X1_8 BUFX2_5/gnd DFFSR_6/S FILL
XNOR3X1_2 NOR3X1_2/A NOR3X1_2/B NOR3X1_2/C INVX1_89/gnd NOR3X1_2/Y DFFSR_2/S NOR3X1
XFILL_35_DFFSR_120 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_25_DFFSR_123 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_26_0_1 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_1_INVX1_170 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_15_DFFSR_126 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_38_DFFSR_38 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_27_DFFSR_78 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_5_AOI21X1_5 BUFX2_37/A DFFSR_81/S FILL
XFILL_24_2_2 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_6_OAI21X1_243 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_6_1_1 BUFX2_35/A DFFSR_14/S FILL
XFILL_11_DFFSR_28 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_0_NAND2X1_140 DFFSR_71/gnd DFFSR_10/S FILL
XDFFSR_35 DFFSR_35/Q DFFSR_2/CLK DFFSR_33/R DFFSR_2/S DFFSR_35/D DFFSR_5/gnd DFFSR_2/S
+ DFFSR
XFILL_4_3_2 BUFX2_6/gnd DFFSR_91/S FILL
XINVX1_100 BUFX2_8/Y BUFX2_16/gnd DFFSR_84/R DFFSR_11/S INVX1
XFILL_1_DFFSR_123 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_42_DFFSR_154 BUFX2_36/A DFFSR_6/S FILL
XFILL_7_OAI21X1_177 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_34_7 INVX1_8/gnd DFFSR_7/S FILL
XFILL_32_DFFSR_157 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_35_DFFSR_85 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_46_DFFSR_45 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_7_NAND3X1_4 INVX1_94/gnd DFFSR_52/S FILL
XFILL_19_DFFSR_35 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_22_DFFSR_160 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_2_DFFSR_42 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_8_OAI21X1_111 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_12_DFFSR_163 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_21_CLKBUF1_22 INVX1_94/gnd DFFSR_25/S FILL
XFILL_2_INVX1_314 INVX1_8/gnd DFFSR_5/S FILL
XFILL_12_XOR2X1_5 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_43_DFFSR_92 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_8_DFFSR_157 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_19_DFFSR_8 BUFX2_36/A DFFSR_8/S FILL
XFILL_49_DFFSR_188 INVX1_2/gnd DFFSR_1/S FILL
XFILL_39_DFFSR_191 INVX1_23/gnd DFFSR_91/S FILL
XFILL_4_AND2X2_1 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_1_INVX1_134 BUFX2_37/A DFFSR_8/S FILL
XFILL_16_DFFSR_82 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_27_DFFSR_42 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_3_BUFX2_9 BUFX2_37/A DFFSR_8/S FILL
XFILL_11_DFFPOSX1_27 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_7_NAND3X1_123 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_6_OAI21X1_207 BUFX2_37/A DFFSR_8/S FILL
XFILL_0_NAND2X1_104 INVX1_4/gnd DFFSR_51/S FILL
XFILL_40_DFFSR_4 INVX1_4/gnd DFFSR_4/S FILL
XOAI21X1_243 INVX1_401/Y AOI21X1_41/B INVX1_402/A BUFX2_6/gnd AOI21X1_42/B DFFSR_14/S
+ OAI21X1
XFILL_24_DFFSR_89 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_21_DFFPOSX1_16 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_7_OAI21X1_141 INVX1_94/gnd DFFSR_52/S FILL
XFILL_7_DFFSR_96 INVX1_2/gnd DFFSR_1/S FILL
XFILL_42_DFFSR_118 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_35_DFFSR_49 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_32_DFFSR_121 BUFX2_36/A DFFSR_6/S FILL
XFILL_22_DFFSR_124 INVX1_89/gnd DFFSR_36/S FILL
XFILL_12_DFFSR_127 BUFX2_43/A DFFSR_97/S FILL
XFILL_6_BUFX2_34 BUFX2_37/A DFFSR_81/S FILL
XFILL_2_AOI21X1_6 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_2_INVX1_278 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_32_DFFSR_96 INVX1_2/gnd DFFSR_1/S FILL
XFILL_43_DFFSR_56 INVX1_2/gnd DFFSR_51/S FILL
XFILL_4_INVX1_90 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_49_DFFSR_152 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_8_DFFSR_121 BUFX2_36/A DFFSR_6/S FILL
XFILL_5_OAI21X1_237 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_39_DFFSR_155 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_29_DFFSR_158 BUFX2_43/A DFFSR_23/S FILL
XFILL_16_DFFSR_46 BUFX2_36/A DFFSR_6/S FILL
XNAND3X1_8 NAND3X1_8/A NAND3X1_8/B NAND3X1_8/C BUFX2_19/gnd NAND3X1_8/Y DFFSR_54/S
+ NAND3X1
XFILL_19_DFFSR_161 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_6_OAI21X1_171 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_4_NAND3X1_5 BUFX2_8/gnd DFFSR_10/S FILL
XNOR2X1_43 NOR2X1_43/A NOR2X1_43/B BUFX2_17/gnd NOR2X1_43/Y DFFSR_7/S NOR2X1
XFILL_51_DFFSR_63 INVX1_94/gnd DFFSR_52/S FILL
XOAI21X1_207 AOI22X1_7/Y AOI22X1_8/Y AOI21X1_26/C BUFX2_37/A NAND3X1_53/B DFFSR_8/S
+ OAI21X1
XFILL_4_NOR2X1_40 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_13_CLKBUF1_10 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_3_INVX1_422 INVX1_23/gnd DFFSR_186/S FILL
XFILL_7_OAI21X1_105 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_6_NAND2X1_285 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_25_3_0 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_12_CLKBUF1_13 INVX1_4/gnd DFFSR_51/S FILL
XFILL_5_DFFSR_158 BUFX2_43/A DFFSR_23/S FILL
XFILL_11_CLKBUF1_16 BUFX2_36/A DFFSR_6/S FILL
XFILL_7_DFFSR_60 BUFX2_37/A DFFSR_8/S FILL
XFILL_24_DFFSR_53 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_13_DFFSR_93 INVX1_2/gnd DFFSR_51/S FILL
XFILL_35_DFFSR_13 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_23_5_1 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_46_DFFSR_189 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_10_CLKBUF1_19 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_5_4_0 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_9_CLKBUF1_22 INVX1_94/gnd DFFSR_25/S FILL
XFILL_7_DFFSR_7 INVX1_8/gnd DFFSR_7/S FILL
XFILL_8_CLKBUF1_25 INVX1_23/gnd DFFSR_186/S FILL
XFILL_2_INVX1_242 BUFX2_36/A DFFSR_6/S FILL
XFILL_6_NAND3X1_117 INVX1_94/gnd DFFSR_25/S FILL
XFILL_43_DFFSR_20 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_5_OAI21X1_201 BUFX2_35/A DFFSR_97/S FILL
XFILL_10_DFFPOSX1_21 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_32_DFFSR_60 BUFX2_37/A DFFSR_8/S FILL
XFILL_4_INVX1_54 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_49_DFFSR_116 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_39_DFFSR_119 BUFX2_37/A DFFSR_81/S FILL
XFILL_16_DFFSR_10 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_29_DFFSR_122 INVX1_94/gnd DFFSR_52/S FILL
XFILL_19_DFFSR_125 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_6_OAI21X1_135 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_20_DFFPOSX1_10 INVX1_8/gnd DFFSR_5/S FILL
XFILL_9_AOI21X1_4 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_40_DFFSR_67 INVX1_2/gnd DFFSR_51/S FILL
XFILL_16_4 BUFX2_37/A DFFSR_81/S FILL
XOAI21X1_171 DFFSR_54/S INVX1_206/Y NAND2X1_171/Y BUFX2_19/gnd DFFSR_171/D DFFSR_54/S
+ OAI21X1
XFILL_3_INVX1_386 INVX1_94/gnd DFFSR_52/S FILL
XFILL_24_DFFSR_17 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_33_0_1 INVX1_8/gnd DFFSR_7/S FILL
XFILL_6_NAND2X1_249 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_13_DFFSR_57 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_7_DFFSR_24 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_46_DFFSR_153 BUFX2_36/A DFFSR_8/S FILL
XFILL_5_DFFSR_122 INVX1_94/gnd DFFSR_52/S FILL
XFILL_36_DFFSR_156 INVX1_23/gnd DFFSR_91/S FILL
XNAND2X1_285 NOR2X1_1/B NOR2X1_1/A DFFSR_71/gnd NAND2X1_285/Y DFFSR_10/S NAND2X1
XFILL_31_2_2 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_4_OAI21X1_231 BUFX2_36/A DFFSR_6/S FILL
XFILL_6_NOR2X1_5 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_26_DFFSR_159 BUFX2_36/A DFFSR_6/S FILL
XFILL_2_INVX1_206 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_48_DFFSR_74 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_16_DFFSR_162 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_1_NAND3X1_6 INVX1_8/gnd DFFSR_7/S FILL
XFILL_4_DFFSR_71 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_32_DFFSR_24 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_5_OAI21X1_165 BUFX2_35/A DFFSR_97/S FILL
XFILL_1_NOR2X1_41 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_21_DFFSR_64 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_0_INVX1_423 BUFX2_37/A DFFSR_8/S FILL
XNAND3X1_117 NOR2X1_1/B NOR2X1_1/A NOR2X1_2/A INVX1_94/gnd OAI22X1_8/B DFFSR_25/S
+ NAND3X1
XFILL_2_DFFSR_159 BUFX2_36/A DFFSR_6/S FILL
XFILL_8_XOR2X1_1 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_5_NAND2X1_279 INVX1_89/gnd DFFSR_2/S FILL
XFILL_43_DFFSR_190 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_1_CLKBUF1_10 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_40_DFFSR_31 BUFX2_35/A DFFSR_97/S FILL
XOAI21X1_135 DFFSR_97/S INVX1_152/Y OAI21X1_135/C BUFX2_5/gnd DFFSR_135/D DFFSR_23/S
+ OAI21X1
XFILL_29_DFFSR_71 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_0_CLKBUF1_13 INVX1_4/gnd DFFSR_51/S FILL
XFILL_1_INVX1_65 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_6_NAND2X1_213 BUFX2_35/A DFFSR_97/S FILL
XFILL_3_INVX1_350 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_3_OAI21X1_261 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_13_DFFSR_21 INVX1_2/gnd DFFSR_1/S FILL
XFILL_46_DFFSR_117 INVX1_23/gnd DFFSR_91/S FILL
XFILL_5_NAND3X1_111 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_4_NOR3X1_2 INVX1_89/gnd DFFSR_2/S FILL
XNAND2X1_249 NOR2X1_42/Y NOR2X1_43/Y BUFX2_17/gnd NAND2X1_144/B DFFSR_7/S NAND2X1
XFILL_36_DFFSR_120 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_26_DFFSR_123 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_4_OAI21X1_195 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_18_DFFSR_5 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_2_INVX1_170 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_16_DFFSR_126 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_48_DFFSR_38 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_37_DFFSR_78 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_6_AOI21X1_5 BUFX2_37/A DFFSR_81/S FILL
XFILL_2_BUFX2_6 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_10_DFFSR_68 BUFX2_35/A DFFSR_14/S FILL
XFILL_21_DFFSR_28 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_4_DFFSR_35 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_5_OAI21X1_129 INVX1_4/gnd DFFSR_4/S FILL
XFILL_0_INVX1_387 INVX1_94/gnd DFFSR_25/S FILL
XFILL_2_DFFSR_123 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_43_DFFSR_154 BUFX2_36/A DFFSR_6/S FILL
XFILL_38_4 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_33_DFFSR_157 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_45_DFFSR_85 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_39_DFFSR_1 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_5_NAND2X1_243 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_24_DFFPOSX1_1 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_8_NAND3X1_4 INVX1_94/gnd DFFSR_52/S FILL
XFILL_1_INVX1_29 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_29_DFFSR_35 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_23_DFFSR_160 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_1_DFFSR_82 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_18_DFFSR_75 INVX1_4/gnd DFFSR_51/S FILL
XFILL_3_OAI21X1_225 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_9_DFFPOSX1_15 BUFX2_35/A DFFSR_14/S FILL
XFILL_23_DFFPOSX1_4 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_13_DFFSR_163 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_22_DFFPOSX1_7 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_6_NAND2X1_177 INVX1_89/gnd DFFSR_36/S FILL
XFILL_3_INVX1_314 INVX1_8/gnd DFFSR_5/S FILL
XFILL_0_BUFX2_20 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_9_DFFSR_157 BUFX2_6/gnd DFFSR_91/S FILL
XNAND2X1_213 AND2X2_5/B AND2X2_8/B BUFX2_35/A XNOR2X1_3/A DFFSR_97/S NAND2X1
XFILL_4_OAI21X1_159 BUFX2_43/A DFFSR_97/S FILL
XFILL_50_DFFSR_188 INVX1_2/gnd DFFSR_1/S FILL
XFILL_9_DFFSR_89 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_40_DFFSR_191 INVX1_23/gnd DFFSR_91/S FILL
XFILL_2_INVX1_134 BUFX2_37/A DFFSR_8/S FILL
XFILL_26_DFFSR_82 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_37_DFFSR_42 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_32_3_0 INVX1_8/gnd DFFSR_5/S FILL
XFILL_10_DFFSR_32 INVX1_2/gnd DFFSR_1/S FILL
XFILL_4_NAND2X1_273 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_0_INVX1_351 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_30_5_1 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_34_DFFSR_89 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_5_NAND2X1_207 BUFX2_43/A DFFSR_97/S FILL
XFILL_2_OAI21X1_255 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_43_DFFSR_118 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_45_DFFSR_49 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_33_DFFSR_121 BUFX2_36/A DFFSR_6/S FILL
XFILL_4_NAND3X1_105 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_23_DFFSR_124 INVX1_89/gnd DFFSR_36/S FILL
XFILL_13_DFFSR_127 BUFX2_43/A DFFSR_97/S FILL
XFILL_1_DFFSR_46 BUFX2_36/A DFFSR_6/S FILL
XFILL_18_DFFSR_39 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_3_AOI21X1_6 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_6_NAND2X1_141 INVX1_94/gnd DFFSR_25/S FILL
XFILL_3_OAI21X1_189 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_3_INVX1_278 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_11_XOR2X1_9 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_6_DFFSR_4 INVX1_4/gnd DFFSR_4/S FILL
XFILL_4_OAI21X1_123 INVX1_23/gnd DFFSR_91/S FILL
XFILL_50_DFFSR_152 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_9_DFFSR_121 BUFX2_36/A DFFSR_6/S FILL
XNAND2X1_177 NAND3X1_1/C NAND3X1_2/A INVX1_89/gnd XOR2X1_1/A DFFSR_36/S NAND2X1
XFILL_42_DFFSR_96 INVX1_2/gnd DFFSR_1/S FILL
XFILL_3_AND2X2_5 BUFX2_37/A DFFSR_81/S FILL
XFILL_40_DFFSR_155 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_26_DFFSR_46 BUFX2_36/A DFFSR_6/S FILL
XFILL_9_DFFSR_53 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_15_DFFSR_86 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_30_DFFSR_158 BUFX2_43/A DFFSR_23/S FILL
XFILL_20_DFFSR_161 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_5_NAND3X1_5 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_4_NAND2X1_237 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_40_0_1 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_10_DFFSR_164 INVX1_89/gnd DFFSR_2/S FILL
XFILL_30_DFFSR_8 BUFX2_36/A DFFSR_8/S FILL
XFILL_0_INVX1_315 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_5_NOR2X1_40 BUFX2_8/gnd DFFSR_10/S FILL
XINVX1_425 XOR2X1_13/A BUFX2_17/gnd NOR2X1_47/A DFFSR_57/S INVX1
XFILL_38_2_2 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_4_INVX1_422 INVX1_23/gnd DFFSR_186/S FILL
XFILL_2_OAI21X1_219 BUFX2_35/A DFFSR_97/S FILL
XFILL_6_DFFSR_158 BUFX2_43/A DFFSR_23/S FILL
XFILL_5_NAND2X1_171 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_34_DFFSR_53 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_23_DFFSR_93 INVX1_2/gnd DFFSR_51/S FILL
XFILL_45_DFFSR_13 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_12_DFFPOSX1_1 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_47_DFFSR_189 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_1_DFFSR_10 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_11_DFFPOSX1_4 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_3_OAI21X1_153 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_5_BUFX2_38 BUFX2_37/A DFFSR_81/S FILL
XFILL_10_DFFPOSX1_7 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_17_DFFPOSX1_28 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_6_NAND2X1_105 BUFX2_35/A DFFSR_14/S FILL
XFILL_3_INVX1_242 BUFX2_36/A DFFSR_6/S FILL
XFILL_42_DFFSR_60 BUFX2_37/A DFFSR_8/S FILL
XFILL_3_INVX1_94 INVX1_94/gnd DFFSR_52/S FILL
XNAND2X1_141 DFFSR_25/S NAND2X1_246/Y INVX1_94/gnd OAI21X1_141/C DFFSR_25/S NAND2X1
XFILL_8_AOI21X1_33 BUFX2_35/A DFFSR_14/S FILL
XFILL_27_DFFPOSX1_17 BUFX2_37/A DFFSR_8/S FILL
XFILL_50_DFFSR_116 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_3_NAND2X1_267 INVX1_4/gnd DFFSR_4/S FILL
XFILL_40_DFFSR_119 BUFX2_37/A DFFSR_81/S FILL
XFILL_7_AOI21X1_36 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_26_DFFSR_10 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_9_DFFSR_17 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_15_DFFSR_50 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_6_AOI21X1_39 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_30_DFFSR_122 INVX1_94/gnd DFFSR_52/S FILL
XFILL_1_OAI21X1_249 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_5_AOI21X1_42 INVX1_23/gnd DFFSR_91/S FILL
XFILL_20_DFFSR_125 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_4_NAND2X1_201 BUFX2_35/A DFFSR_14/S FILL
XAOI21X1_39 AOI21X1_39/A AOI21X1_39/B INVX1_251/A BUFX2_7/gnd OAI22X1_4/B DFFSR_81/S
+ AOI21X1
XFILL_10_DFFSR_128 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_4_AOI21X1_45 INVX1_89/gnd DFFSR_36/S FILL
XFILL_0_AOI21X1_7 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_50_DFFSR_67 INVX1_2/gnd DFFSR_51/S FILL
XFILL_0_INVX1_279 INVX1_4/gnd DFFSR_51/S FILL
XINVX1_389 INVX1_90/A DFFSR_73/gnd INVX1_389/Y DFFSR_57/S INVX1
XFILL_20_1 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_3_AOI21X1_48 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_5_NAND2X1_135 BUFX2_36/A DFFSR_6/S FILL
XFILL_4_INVX1_386 INVX1_94/gnd DFFSR_52/S FILL
XFILL_34_DFFSR_17 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_2_OAI21X1_183 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_23_DFFSR_57 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_6_DFFSR_64 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_12_DFFSR_97 BUFX2_35/A DFFSR_97/S FILL
XFILL_47_DFFSR_153 BUFX2_36/A DFFSR_8/S FILL
XFILL_6_DFFSR_122 INVX1_94/gnd DFFSR_52/S FILL
XFILL_37_DFFSR_156 INVX1_23/gnd DFFSR_91/S FILL
XBUFX2_42 BUFX2_43/A BUFX2_5/gnd BUFX2_42/Y DFFSR_23/S BUFX2
XFILL_3_OAI21X1_117 BUFX2_35/A DFFSR_97/S FILL
XFILL_27_DFFSR_159 BUFX2_36/A DFFSR_6/S FILL
XFILL_3_INVX1_206 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_17_DFFSR_162 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_8_OAI21X1_81 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_17_DFFSR_2 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_2_NAND3X1_6 INVX1_8/gnd DFFSR_7/S FILL
XFILL_7_OAI21X1_84 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_42_DFFSR_24 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_3_INVX1_58 BUFX2_16/gnd DFFSR_65/S FILL
XNAND2X1_105 DFFSR_97/Q BUFX2_21/Y BUFX2_35/A OAI21X1_105/C DFFSR_14/S NAND2X1
XFILL_3_NAND2X1_231 BUFX2_37/A DFFSR_81/S FILL
XFILL_2_NOR2X1_41 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_6_OAI21X1_87 INVX1_4/gnd DFFSR_4/S FILL
XFILL_31_DFFSR_64 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_12_0_2 BUFX2_36/A DFFSR_6/S FILL
XFILL_1_INVX1_423 BUFX2_37/A DFFSR_8/S FILL
XFILL_1_BUFX2_3 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_5_OAI21X1_90 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_2_NAND3X1_129 BUFX2_35/A DFFSR_14/S FILL
XFILL_15_DFFSR_14 BUFX2_35/A DFFSR_14/S FILL
XFILL_3_DFFSR_159 BUFX2_36/A DFFSR_6/S FILL
XFILL_4_OAI21X1_93 INVX1_4/gnd DFFSR_51/S FILL
XOAI21X1_87 BUFX2_15/Y INVX1_98/Y NAND2X1_87/Y INVX1_4/gnd DFFSR_87/D DFFSR_4/S OAI21X1
XFILL_44_DFFSR_190 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_3_OAI21X1_96 INVX1_4/gnd DFFSR_51/S FILL
XFILL_2_OAI21X1_99 BUFX2_43/A DFFSR_97/S FILL
XFILL_1_OAI21X1_213 BUFX2_36/A DFFSR_6/S FILL
XFILL_4_NAND2X1_165 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_50_DFFSR_31 BUFX2_35/A DFFSR_97/S FILL
XINVX1_353 DFFSR_91/Q BUFX2_37/A INVX1_353/Y DFFSR_8/S INVX1
XFILL_0_INVX1_243 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_39_DFFSR_71 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_3_AOI21X1_12 INVX1_8/gnd DFFSR_7/S FILL
XFILL_2_OAI21X1_147 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_2_AOI21X1_15 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_4_INVX1_350 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_16_DFFPOSX1_22 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_0_DFFPOSX1_1 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_12_DFFSR_61 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_6_DFFSR_28 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_1_AOI21X1_18 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_23_DFFSR_21 INVX1_2/gnd DFFSR_1/S FILL
XFILL_47_DFFSR_117 INVX1_23/gnd DFFSR_91/S FILL
XFILL_0_AOI21X1_21 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_5_NOR2X1_9 BUFX2_43/A DFFSR_97/S FILL
XFILL_39_3_0 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_37_DFFSR_120 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_27_DFFSR_123 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_2_NAND2X1_261 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_26_DFFPOSX1_11 INVX1_4/gnd DFFSR_4/S FILL
XFILL_3_INVX1_170 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_8_OAI21X1_45 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_17_DFFSR_126 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_47_DFFSR_78 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_37_5_1 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_7_AOI21X1_5 BUFX2_37/A DFFSR_81/S FILL
XFILL_6_NAND2X1_66 INVX1_4/gnd DFFSR_51/S FILL
XFILL_0_OAI21X1_243 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_20_DFFSR_68 BUFX2_35/A DFFSR_14/S FILL
XFILL_31_DFFSR_28 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_3_INVX1_22 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_3_DFFSR_75 INVX1_4/gnd DFFSR_51/S FILL
XFILL_7_OAI21X1_48 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_3_NAND2X1_195 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_5_NAND2X1_69 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_6_OAI21X1_51 INVX1_2/gnd DFFSR_51/S FILL
XNAND2X1_66 BUFX2_24/Y NAND2X1_66/B INVX1_4/gnd OAI21X1_66/C DFFSR_51/S NAND2X1
XFILL_5_OAI21X1_54 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_1_INVX1_387 INVX1_94/gnd DFFSR_25/S FILL
XFILL_4_NAND2X1_72 DFFSR_5/gnd DFFSR_2/S FILL
XOAI21X1_51 DFFSR_1/S INVX1_58/Y OAI21X1_51/C INVX1_2/gnd DFFSR_51/D DFFSR_51/S OAI21X1
XFILL_7_XOR2X1_5 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_3_DFFSR_123 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_44_DFFSR_154 BUFX2_36/A DFFSR_6/S FILL
XFILL_2_BUFX2_13 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_3_NAND2X1_75 INVX1_4/gnd DFFSR_4/S FILL
XFILL_42_1 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_4_OAI21X1_57 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_3_OAI21X1_60 BUFX2_37/A DFFSR_81/S FILL
XFILL_10_AOI22X1_1 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_1_OAI21X1_177 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_4_NAND2X1_129 INVX1_4/gnd DFFSR_4/S FILL
XFILL_2_NAND2X1_78 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_34_DFFSR_157 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_2_OAI21X1_63 INVX1_94/gnd DFFSR_25/S FILL
XFILL_1_NAND2X1_81 INVX1_94/gnd DFFSR_25/S FILL
XFILL_0_INVX1_207 BUFX2_36/A DFFSR_6/S FILL
XFILL_0_NAND2X1_84 BUFX2_36/A DFFSR_6/S FILL
XFILL_0_INVX1_69 BUFX2_36/A DFFSR_8/S FILL
XFILL_9_NAND3X1_4 INVX1_94/gnd DFFSR_52/S FILL
XINVX1_317 DFFSR_39/Q DFFSR_79/gnd INVX1_317/Y DFFSR_45/S INVX1
XFILL_39_DFFSR_35 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_24_DFFSR_160 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_1_OAI21X1_66 INVX1_4/gnd DFFSR_51/S FILL
XFILL_28_DFFSR_75 INVX1_4/gnd DFFSR_51/S FILL
XFILL_0_OAI21X1_69 BUFX2_37/A DFFSR_8/S FILL
XFILL_14_DFFSR_163 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_2_OAI21X1_111 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_4_INVX1_314 INVX1_8/gnd DFFSR_5/S FILL
XFILL_12_DFFSR_25 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_2_NAND2X1_225 BUFX2_36/A DFFSR_8/S FILL
XDFFSR_5 DFFSR_5/Q DFFSR_2/CLK DFFSR_6/R DFFSR_5/S DFFSR_5/D DFFSR_5/gnd DFFSR_5/S
+ DFFSR
XFILL_0_DFFSR_160 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_5_DFFSR_1 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_47_0_1 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_41_DFFSR_191 INVX1_23/gnd DFFSR_91/S FILL
XFILL_3_INVX1_134 BUFX2_37/A DFFSR_8/S FILL
XFILL_36_DFFSR_82 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_47_DFFSR_42 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_1_NAND3X1_123 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_7_OAI21X1_12 BUFX2_35/A DFFSR_14/S FILL
XFILL_3_DFFSR_39 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_6_NAND2X1_30 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_45_2_2 INVX1_2/gnd DFFSR_1/S FILL
XFILL_3_NAND2X1_159 BUFX2_43/A DFFSR_97/S FILL
XFILL_0_OAI21X1_207 BUFX2_37/A DFFSR_8/S FILL
XFILL_5_NAND2X1_33 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_6_OAI21X1_15 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_20_DFFSR_32 INVX1_2/gnd DFFSR_1/S FILL
XFILL_1_INVX1_351 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_3_OR2X2_1 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_4_NAND2X1_36 DFFSR_71/gnd DFFSR_45/S FILL
XNAND2X1_30 DFFSR_2/S INVX1_25/A DFFSR_79/gnd NAND2X1_30/Y DFFSR_36/S NAND2X1
XFILL_5_OAI21X1_18 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_3_NAND2X1_39 DFFSR_71/gnd DFFSR_10/S FILL
XOAI21X1_15 DFFSR_15/S INVX1_17/Y NAND2X1_15/Y BUFX2_17/gnd DFFSR_15/D DFFSR_57/S
+ OAI21X1
XFILL_4_OAI21X1_21 INVX1_2/gnd DFFSR_51/S FILL
XFILL_44_DFFSR_89 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_15_DFFPOSX1_16 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_13_XOR2X1_2 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_29_DFFSR_5 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_2_NAND2X1_42 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_44_DFFSR_118 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_3_OAI21X1_24 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_34_DFFSR_121 BUFX2_36/A DFFSR_6/S FILL
XFILL_1_OAI21X1_141 INVX1_94/gnd DFFSR_52/S FILL
XFILL_1_NAND2X1_45 INVX1_89/gnd DFFSR_36/S FILL
XFILL_2_OAI21X1_27 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_13_1_0 BUFX2_36/A DFFSR_8/S FILL
XFILL_1_OAI21X1_30 INVX1_89/gnd DFFSR_36/S FILL
XFILL_24_DFFSR_124 INVX1_89/gnd DFFSR_36/S FILL
XFILL_0_NAND2X1_48 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_0_INVX1_171 BUFX2_35/A DFFSR_14/S FILL
XFILL_14_DFFSR_127 BUFX2_43/A DFFSR_97/S FILL
XFILL_0_OAI21X1_33 BUFX2_19/gnd DFFSR_52/S FILL
XAOI21X1_9 INVX1_224/Y AOI21X1_9/B AOI21X1_8/Y INVX1_94/gnd AOI21X1_9/Y DFFSR_52/S
+ AOI21X1
XFILL_28_DFFSR_39 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_17_DFFSR_79 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_0_DFFSR_86 DFFSR_1/gnd DFFSR_9/S FILL
XINVX1_281 DFFSR_3/Q DFFSR_3/gnd INVX1_281/Y DFFSR_65/S INVX1
XFILL_0_INVX1_33 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_11_3_1 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_4_AOI21X1_6 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_4_INVX1_278 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_1_NAND2X1_255 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_5_DFFPOSX1_27 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_50_DFFSR_1 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_2_NAND2X1_189 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_41_DFFSR_155 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_0_DFFSR_124 INVX1_89/gnd DFFSR_36/S FILL
XFILL_5_AOI22X1_11 INVX1_23/gnd DFFSR_91/S FILL
XFILL_36_DFFSR_46 BUFX2_36/A DFFSR_6/S FILL
XFILL_25_DFFSR_86 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_8_DFFSR_93 INVX1_2/gnd DFFSR_51/S FILL
XFILL_31_DFFSR_158 BUFX2_43/A DFFSR_23/S FILL
XFILL_4_AOI22X1_14 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_21_DFFSR_161 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_0_OAI21X1_171 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_6_NAND3X1_5 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_9_OAI21X1_226 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_3_NAND2X1_123 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_11_DFFSR_164 INVX1_89/gnd DFFSR_2/S FILL
XINVX1_7 DFFSR_6/Q BUFX2_36/A INVX1_7/Y DFFSR_8/S INVX1
XFILL_1_INVX1_315 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_6_NOR2X1_40 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_11_OAI22X1_41 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_10_OAI22X1_44 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_1_OAI21X1_105 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_7_DFFSR_158 BUFX2_43/A DFFSR_23/S FILL
XFILL_44_DFFSR_53 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_0_NAND2X1_285 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_33_DFFSR_93 INVX1_2/gnd DFFSR_51/S FILL
XFILL_48_DFFSR_189 DFFSR_1/gnd DFFSR_1/S FILL
XINVX1_245 XNOR2X1_1/Y BUFX2_35/A INVX1_245/Y DFFSR_14/S INVX1
XFILL_8_NAND3X1_65 BUFX2_35/A DFFSR_14/S FILL
XFILL_9_OAI22X1_47 BUFX2_37/A DFFSR_8/S FILL
XAND2X2_2 BUFX2_11/Y AND2X2_9/A BUFX2_7/gnd AND2X2_2/Y DFFSR_54/S AND2X2
XFILL_17_DFFSR_43 INVX1_94/gnd DFFSR_25/S FILL
XFILL_0_NAND2X1_12 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_0_INVX1_135 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_0_DFFSR_50 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_7_NAND3X1_68 BUFX2_35/A DFFSR_14/S FILL
XFILL_8_OAI22X1_50 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_6_NAND3X1_71 BUFX2_35/A DFFSR_14/S FILL
XFILL_1_NAND2X1_219 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_19_0_2 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_7_OAI22X1_53 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_5_NAND3X1_74 BUFX2_35/A DFFSR_14/S FILL
XFILL_6_OAI22X1_56 BUFX2_37/A DFFSR_8/S FILL
XFILL_0_NAND3X1_117 INVX1_94/gnd DFFSR_25/S FILL
XNAND3X1_71 XNOR2X1_1/Y NAND3X1_71/B NAND3X1_71/C BUFX2_35/A NAND3X1_71/Y DFFSR_14/S
+ NAND3X1
XFILL_4_NAND3X1_77 BUFX2_37/A DFFSR_81/S FILL
XFILL_5_OAI22X1_59 INVX1_8/gnd DFFSR_7/S FILL
XFILL_2_NAND2X1_153 BUFX2_5/gnd DFFSR_6/S FILL
XOAI22X1_56 INVX1_370/Y OAI22X1_40/B INVX1_371/Y OAI22X1_40/D BUFX2_37/A NOR2X1_37/A
+ DFFSR_8/S OAI22X1
XFILL_3_NAND3X1_80 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_4_OAI22X1_62 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_8_OAI21X1_256 INVX1_2/gnd DFFSR_51/S FILL
XFILL_2_AND2X2_9 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_2_NAND3X1_83 BUFX2_37/A DFFSR_81/S FILL
XFILL_41_DFFSR_119 BUFX2_37/A DFFSR_81/S FILL
XFILL_36_DFFSR_10 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_8_DFFSR_57 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_14_DFFSR_90 INVX1_2/gnd DFFSR_1/S FILL
XFILL_25_DFFSR_50 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_3_OAI22X1_65 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_10_XNOR2X1_1 BUFX2_35/A DFFSR_14/S FILL
XFILL_1_NAND3X1_86 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_31_DFFSR_122 INVX1_94/gnd DFFSR_52/S FILL
XFILL_2_OAI22X1_68 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_21_DFFSR_125 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_0_NAND3X1_89 BUFX2_43/A DFFSR_23/S FILL
XFILL_14_DFFPOSX1_10 INVX1_8/gnd DFFSR_5/S FILL
XFILL_0_OAI21X1_135 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_9_OAI21X1_190 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_11_DFFSR_128 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_1_AOI21X1_7 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_1_INVX1_279 INVX1_4/gnd DFFSR_51/S FILL
XFILL_46_3_0 DFFSR_1/gnd DFFSR_1/S FILL
XINVX1_91 BUFX2_9/Y BUFX2_19/gnd DFFSR_76/R DFFSR_52/S INVX1
XFILL_44_DFFSR_17 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_0_NAND2X1_249 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_22_DFFSR_97 BUFX2_35/A DFFSR_97/S FILL
XFILL_48_DFFSR_153 BUFX2_36/A DFFSR_8/S FILL
XFILL_7_DFFSR_122 INVX1_94/gnd DFFSR_52/S FILL
XFILL_33_DFFSR_57 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_8_NAND3X1_29 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_44_5_1 INVX1_2/gnd DFFSR_51/S FILL
XFILL_9_OAI22X1_11 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_38_DFFSR_156 INVX1_23/gnd DFFSR_91/S FILL
XFILL_0_DFFSR_14 BUFX2_35/A DFFSR_14/S FILL
XINVX1_209 AND2X2_11/B BUFX2_43/A INVX1_209/Y DFFSR_23/S INVX1
XFILL_4_BUFX2_42 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_7_NAND3X1_32 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_8_OAI22X1_14 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_6_NAND3X1_35 BUFX2_35/A DFFSR_97/S FILL
XFILL_4_DFFPOSX1_21 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_28_DFFSR_159 BUFX2_36/A DFFSR_6/S FILL
XFILL_7_OAI22X1_17 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_1_NAND2X1_183 INVX1_8/gnd DFFSR_7/S FILL
XFILL_18_DFFSR_162 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_5_NAND3X1_38 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_41_DFFSR_8 BUFX2_36/A DFFSR_8/S FILL
XFILL_6_OAI22X1_20 BUFX2_8/gnd DFFSR_25/S FILL
XNAND3X1_35 NAND3X1_35/A INVX1_239/Y NAND3X1_35/C BUFX2_35/A AOI22X1_7/A DFFSR_97/S
+ NAND3X1
XFILL_4_NAND3X1_41 BUFX2_43/A DFFSR_23/S FILL
XFILL_5_OAI22X1_23 INVX1_89/gnd DFFSR_2/S FILL
XFILL_3_NAND3X1_6 INVX1_8/gnd DFFSR_7/S FILL
XFILL_3_NAND3X1_44 BUFX2_5/gnd DFFSR_23/S FILL
XOAI22X1_20 INVX1_295/Y OAI22X1_8/B INVX1_296/Y OAI22X1_9/D BUFX2_8/gnd NOR2X1_19/B
+ DFFSR_25/S OAI22X1
XFILL_3_NOR2X1_41 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_2_INVX1_98 INVX1_4/gnd DFFSR_4/S FILL
XFILL_41_DFFSR_64 BUFX2_16/gnd DFFSR_11/S FILL
XDFFSR_162 DFFSR_162/Q CLKBUF1_14/Y DFFSR_162/R DFFSR_92/S DFFSR_162/D DFFSR_89/gnd
+ DFFSR_92/S DFFSR
XFILL_2_NAND2X1_117 BUFX2_35/A DFFSR_14/S FILL
XFILL_8_OAI21X1_220 BUFX2_43/A DFFSR_97/S FILL
XFILL_2_INVX1_423 BUFX2_37/A DFFSR_8/S FILL
XFILL_4_OAI22X1_26 INVX1_94/gnd DFFSR_52/S FILL
XFILL_25_DFFSR_14 BUFX2_35/A DFFSR_14/S FILL
XFILL_2_NAND3X1_47 BUFX2_43/A DFFSR_97/S FILL
XFILL_4_DFFSR_159 BUFX2_36/A DFFSR_6/S FILL
XFILL_14_DFFSR_54 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_3_OAI22X1_29 INVX1_8/gnd DFFSR_5/S FILL
XFILL_8_DFFSR_21 INVX1_2/gnd DFFSR_1/S FILL
XFILL_1_NAND3X1_50 BUFX2_37/A DFFSR_81/S FILL
XFILL_2_OAI22X1_32 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_45_DFFSR_190 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_0_NAND3X1_53 BUFX2_37/A DFFSR_81/S FILL
XFILL_1_OAI22X1_35 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_0_OAI22X1_38 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_23_DFFPOSX1_29 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_7_2 BUFX2_35/A DFFSR_14/S FILL
XFILL_1_INVX1_243 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_49_DFFSR_71 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_5_DFFSR_68 BUFX2_35/A DFFSR_14/S FILL
XFILL_0_NAND2X1_213 BUFX2_35/A DFFSR_97/S FILL
XFILL_22_DFFSR_61 BUFX2_5/gnd DFFSR_6/S FILL
XINVX1_55 BUFX2_7/Y BUFX2_36/A DFFSR_46/R DFFSR_8/S INVX1
XFILL_33_DFFSR_21 INVX1_2/gnd DFFSR_1/S FILL
XFILL_48_DFFSR_117 INVX1_23/gnd DFFSR_91/S FILL
XINVX1_173 BUFX2_5/Y BUFX2_35/A DFFSR_149/R DFFSR_14/S INVX1
XFILL_38_DFFSR_120 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_1_NAND2X1_147 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_28_DFFSR_123 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_4_INVX1_170 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_7_OAI21X1_250 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_18_DFFSR_126 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_8_AOI21X1_5 BUFX2_37/A DFFSR_81/S FILL
XFILL_30_DFFSR_68 BUFX2_35/A DFFSR_14/S FILL
XFILL_41_DFFSR_28 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_2_INVX1_62 INVX1_89/gnd DFFSR_2/S FILL
XFILL_8_OAI21X1_184 BUFX2_19/gnd DFFSR_52/S FILL
XDFFSR_126 INVX1_378/A CLKBUF1_4/Y DFFSR_123/R DFFSR_57/S DFFSR_126/D BUFX2_17/gnd
+ DFFSR_57/S DFFSR
XFILL_2_NAND3X1_11 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_20_1_0 INVX1_94/gnd DFFSR_52/S FILL
XFILL_2_INVX1_387 INVX1_94/gnd DFFSR_25/S FILL
XFILL_29_3 INVX1_89/gnd DFFSR_36/S FILL
XFILL_14_DFFSR_18 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_4_DFFSR_123 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_45_DFFSR_154 BUFX2_36/A DFFSR_6/S FILL
XFILL_1_NAND3X1_14 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_11_AOI22X1_1 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_18_3_1 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_0_NAND3X1_17 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_35_DFFSR_157 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_28_DFFSR_2 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_0_2_0 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_1_INVX1_207 BUFX2_36/A DFFSR_6/S FILL
XFILL_49_DFFSR_35 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_25_DFFSR_160 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_38_DFFSR_75 INVX1_4/gnd DFFSR_51/S FILL
XFILL_16_5_2 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_15_DFFSR_163 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_3_DFFPOSX1_15 BUFX2_35/A DFFSR_14/S FILL
XFILL_0_NAND3X1_7 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_0_NAND2X1_177 INVX1_89/gnd DFFSR_36/S FILL
XDFFSR_72 INVX1_81/A CLKBUF1_3/Y DFFSR_68/R DFFSR_7/S DFFSR_72/D BUFX2_17/gnd DFFSR_7/S
+ DFFSR
XFILL_5_DFFSR_32 INVX1_2/gnd DFFSR_1/S FILL
XINVX1_19 BUFX2_8/Y DFFSR_3/gnd DFFSR_9/R DFFSR_65/S INVX1
XFILL_22_DFFSR_25 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_0_NOR2X1_42 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_11_DFFSR_65 DFFSR_3/gnd DFFSR_65/S FILL
XINVX1_137 DFFSR_121/Q BUFX2_36/A INVX1_137/Y DFFSR_8/S INVX1
XFILL_8_NAND3X1_130 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_1_DFFSR_160 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_42_DFFSR_191 INVX1_23/gnd DFFSR_91/S FILL
XFILL_7_OAI21X1_214 BUFX2_35/A DFFSR_97/S FILL
XFILL_4_INVX1_134 BUFX2_37/A DFFSR_8/S FILL
XFILL_1_NAND2X1_111 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_46_DFFSR_82 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_2_INVX1_26 BUFX2_43/A DFFSR_23/S FILL
XFILL_2_DFFSR_79 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_19_DFFSR_72 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_30_DFFSR_32 INVX1_2/gnd DFFSR_1/S FILL
XFILL_8_OAI21X1_148 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_22_DFFPOSX1_23 INVX1_23/gnd DFFSR_91/S FILL
XFILL_2_INVX1_351 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_1_BUFX2_17 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_6_XOR2X1_9 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_45_DFFSR_118 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_35_DFFSR_121 BUFX2_36/A DFFSR_6/S FILL
XFILL_26_0_2 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_25_DFFSR_124 INVX1_89/gnd DFFSR_36/S FILL
XFILL_1_INVX1_171 BUFX2_35/A DFFSR_14/S FILL
XFILL_15_DFFSR_127 BUFX2_43/A DFFSR_97/S FILL
XFILL_38_DFFSR_39 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_27_DFFSR_79 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_5_AOI21X1_6 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_6_1_2 BUFX2_35/A DFFSR_14/S FILL
XFILL_0_NAND2X1_141 INVX1_94/gnd DFFSR_25/S FILL
XDFFSR_36 INVX1_41/A DFFSR_52/CLK DFFSR_33/R DFFSR_36/S DFFSR_36/D DFFSR_79/gnd DFFSR_36/S
+ DFFSR
XFILL_11_DFFSR_29 INVX1_4/gnd DFFSR_4/S FILL
XFILL_6_OAI21X1_244 DFFSR_3/gnd DFFSR_4/S FILL
XINVX1_101 DFFSR_89/Q BUFX2_35/A INVX1_101/Y DFFSR_14/S INVX1
XFILL_1_DFFSR_124 INVX1_89/gnd DFFSR_36/S FILL
XFILL_34_8 INVX1_8/gnd DFFSR_7/S FILL
XFILL_46_DFFSR_46 BUFX2_36/A DFFSR_6/S FILL
XFILL_42_DFFSR_155 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_7_OAI21X1_178 INVX1_94/gnd DFFSR_25/S FILL
XFILL_35_DFFSR_86 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_32_DFFSR_158 BUFX2_43/A DFFSR_23/S FILL
XFILL_22_DFFSR_161 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_2_DFFSR_43 INVX1_94/gnd DFFSR_25/S FILL
XFILL_19_DFFSR_36 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_7_NAND3X1_5 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_12_DFFSR_164 INVX1_89/gnd DFFSR_2/S FILL
XFILL_8_OAI21X1_112 INVX1_4/gnd DFFSR_4/S FILL
XFILL_2_INVX1_315 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_12_XOR2X1_6 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_8_DFFSR_158 BUFX2_43/A DFFSR_23/S FILL
XFILL_19_DFFSR_9 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_43_DFFSR_93 INVX1_2/gnd DFFSR_51/S FILL
XFILL_49_DFFSR_189 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_4_AND2X2_2 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_16_DFFSR_83 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_27_DFFSR_43 INVX1_94/gnd DFFSR_25/S FILL
XFILL_1_INVX1_135 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_7_NAND3X1_124 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_11_DFFPOSX1_28 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_0_NAND2X1_105 BUFX2_35/A DFFSR_14/S FILL
XFILL_6_OAI21X1_208 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_40_DFFSR_5 DFFSR_5/gnd DFFSR_5/S FILL
XOAI21X1_244 DFFSR_11/S INVX1_406/Y OAI21X1_244/C DFFSR_3/gnd DFFSR_176/D DFFSR_4/S
+ OAI21X1
XFILL_7_DFFSR_97 BUFX2_35/A DFFSR_97/S FILL
XFILL_21_DFFPOSX1_17 BUFX2_37/A DFFSR_8/S FILL
XFILL_42_DFFSR_119 BUFX2_37/A DFFSR_81/S FILL
XFILL_7_OAI21X1_142 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_46_DFFSR_10 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_35_DFFSR_50 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_11_XNOR2X1_1 BUFX2_35/A DFFSR_14/S FILL
XFILL_32_DFFSR_122 INVX1_94/gnd DFFSR_52/S FILL
XFILL_24_DFFSR_90 INVX1_2/gnd DFFSR_1/S FILL
XFILL_22_DFFSR_125 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_6_BUFX2_35 BUFX2_35/A DFFSR_14/S FILL
XFILL_12_DFFSR_128 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_2_AOI21X1_7 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_2_INVX1_279 INVX1_4/gnd DFFSR_51/S FILL
XFILL_32_DFFSR_97 BUFX2_35/A DFFSR_97/S FILL
XFILL_49_DFFSR_153 BUFX2_36/A DFFSR_8/S FILL
XFILL_5_OAI21X1_238 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_4_INVX1_91 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_8_DFFSR_122 INVX1_94/gnd DFFSR_52/S FILL
XFILL_43_DFFSR_57 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_39_DFFSR_156 INVX1_23/gnd DFFSR_91/S FILL
XFILL_16_DFFSR_47 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_29_DFFSR_159 BUFX2_36/A DFFSR_6/S FILL
XNAND3X1_9 NAND3X1_7/Y AOI21X1_6/C NAND3X1_8/Y BUFX2_19/gnd NAND3X1_9/Y DFFSR_52/S
+ NAND3X1
XFILL_19_DFFSR_162 DFFSR_89/gnd DFFSR_92/S FILL
XNOR2X1_44 NOR2X1_44/A BUFX2_6/Y BUFX2_6/gnd NOR2X1_44/Y DFFSR_91/S NOR2X1
XFILL_6_OAI21X1_172 BUFX2_36/A DFFSR_6/S FILL
XFILL_27_1_0 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_4_NAND3X1_6 INVX1_8/gnd DFFSR_7/S FILL
XFILL_13_CLKBUF1_11 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_4_NOR2X1_41 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_12_CLKBUF1_14 BUFX2_43/A DFFSR_23/S FILL
XOAI21X1_208 AOI21X1_16/Y AOI21X1_15/Y AOI21X1_23/C BUFX2_5/gnd NAND3X1_53/C DFFSR_6/S
+ OAI21X1
XFILL_3_INVX1_423 BUFX2_37/A DFFSR_8/S FILL
XFILL_25_3_1 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_6_NAND2X1_286 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_35_DFFSR_14 BUFX2_35/A DFFSR_14/S FILL
XFILL_7_2_0 BUFX2_35/A DFFSR_97/S FILL
XFILL_7_DFFSR_61 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_5_DFFSR_159 BUFX2_36/A DFFSR_6/S FILL
XFILL_24_DFFSR_54 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_11_CLKBUF1_17 INVX1_94/gnd DFFSR_25/S FILL
XFILL_7_OAI21X1_106 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_13_DFFSR_94 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_23_5_2 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_46_DFFSR_190 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_10_CLKBUF1_20 INVX1_4/gnd DFFSR_51/S FILL
XFILL_5_4_1 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_9_CLKBUF1_23 INVX1_89/gnd DFFSR_2/S FILL
XFILL_7_DFFSR_8 BUFX2_36/A DFFSR_8/S FILL
XFILL_2_INVX1_243 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_6_NAND3X1_118 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_5_OAI21X1_202 BUFX2_35/A DFFSR_14/S FILL
XFILL_32_DFFSR_61 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_4_INVX1_55 BUFX2_36/A DFFSR_8/S FILL
XFILL_43_DFFSR_21 INVX1_2/gnd DFFSR_1/S FILL
XFILL_10_DFFPOSX1_22 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_49_DFFSR_117 INVX1_23/gnd DFFSR_91/S FILL
XFILL_39_DFFSR_120 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_16_DFFSR_11 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_29_DFFSR_123 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_6_OAI21X1_136 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_19_DFFSR_126 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_20_DFFPOSX1_11 INVX1_4/gnd DFFSR_4/S FILL
XFILL_40_DFFSR_68 BUFX2_35/A DFFSR_14/S FILL
XOAI21X1_172 DFFSR_8/S INVX1_207/Y NAND2X1_172/Y BUFX2_36/A DFFSR_172/D DFFSR_6/S
+ OAI21X1
XFILL_3_INVX1_387 INVX1_94/gnd DFFSR_25/S FILL
XFILL_7_DFFSR_25 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_6_NAND2X1_250 INVX1_8/gnd DFFSR_5/S FILL
XFILL_33_0_2 INVX1_8/gnd DFFSR_7/S FILL
XFILL_5_DFFSR_123 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_24_DFFSR_18 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_13_DFFSR_58 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_46_DFFSR_154 BUFX2_36/A DFFSR_6/S FILL
XFILL_36_DFFSR_157 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_4_OAI21X1_232 BUFX2_35/A DFFSR_97/S FILL
XNAND2X1_286 NOR2X1_2/A NAND2X1_285/Y DFFSR_71/gnd AOI21X1_48/B DFFSR_45/S NAND2X1
XFILL_6_NOR2X1_6 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_2_INVX1_207 BUFX2_36/A DFFSR_6/S FILL
XFILL_26_DFFSR_160 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_48_DFFSR_75 INVX1_4/gnd DFFSR_51/S FILL
XFILL_16_DFFSR_163 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_1_NAND3X1_7 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_32_DFFSR_25 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_4_DFFSR_72 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_1_NOR2X1_42 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_5_OAI21X1_166 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_21_DFFSR_65 DFFSR_3/gnd DFFSR_65/S FILL
XNAND3X1_118 NOR2X1_1/B NOR2X1_2/A INVX1_264/Y DFFSR_79/gnd OAI22X1_8/D DFFSR_45/S
+ NAND3X1
XFILL_0_INVX1_424 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_3_BUFX2_10 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_2_DFFSR_160 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_43_DFFSR_191 INVX1_23/gnd DFFSR_91/S FILL
XFILL_8_XOR2X1_2 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_5_NAND2X1_280 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_6_OAI21X1_100 INVX1_23/gnd DFFSR_91/S FILL
XFILL_1_CLKBUF1_11 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_0_CLKBUF1_14 BUFX2_43/A DFFSR_23/S FILL
XFILL_29_DFFSR_72 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_40_DFFSR_32 INVX1_2/gnd DFFSR_1/S FILL
XFILL_1_INVX1_66 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_6_NAND2X1_214 BUFX2_35/A DFFSR_97/S FILL
XFILL_3_INVX1_351 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_3_OAI21X1_262 INVX1_89/gnd DFFSR_36/S FILL
XOAI21X1_136 DFFSR_5/S INVX1_153/Y NAND2X1_136/Y DFFSR_5/gnd DFFSR_136/D DFFSR_2/S
+ OAI21X1
XFILL_13_DFFSR_22 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_5_NAND3X1_112 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_46_DFFSR_118 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_36_DFFSR_121 BUFX2_36/A DFFSR_6/S FILL
XNAND2X1_250 INVX1_397/A INVX1_396/Y INVX1_8/gnd NAND2X1_250/Y DFFSR_5/S NAND2X1
XFILL_18_DFFSR_6 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_4_OAI21X1_196 INVX1_94/gnd DFFSR_25/S FILL
XFILL_26_DFFSR_124 INVX1_89/gnd DFFSR_36/S FILL
XFILL_2_INVX1_171 BUFX2_35/A DFFSR_14/S FILL
XFILL_16_DFFSR_127 BUFX2_43/A DFFSR_97/S FILL
XFILL_48_DFFSR_39 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_37_DFFSR_79 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_6_AOI21X1_6 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_10_DFFSR_69 BUFX2_43/A DFFSR_23/S FILL
XFILL_2_BUFX2_7 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_4_DFFSR_36 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_5_OAI21X1_130 INVX1_4/gnd DFFSR_4/S FILL
XFILL_21_DFFSR_29 INVX1_4/gnd DFFSR_4/S FILL
XFILL_0_INVX1_388 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_2_DFFSR_124 INVX1_89/gnd DFFSR_36/S FILL
XFILL_38_5 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_43_DFFSR_155 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_5_NAND2X1_244 INVX1_94/gnd DFFSR_52/S FILL
XFILL_39_DFFSR_2 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_45_DFFSR_86 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_33_DFFSR_158 BUFX2_43/A DFFSR_23/S FILL
XFILL_23_DFFSR_161 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_18_DFFSR_76 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_1_DFFSR_83 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_29_DFFSR_36 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_24_DFFPOSX1_2 INVX1_89/gnd DFFSR_36/S FILL
XFILL_1_INVX1_30 DFFSR_1/gnd DFFSR_9/S FILL
XOAI21X1_100 BUFX2_21/Y INVX1_113/Y OAI21X1_100/C INVX1_23/gnd DFFSR_100/D DFFSR_91/S
+ OAI21X1
XFILL_3_OAI21X1_226 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_9_DFFPOSX1_16 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_8_NAND3X1_5 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_13_DFFSR_164 INVX1_89/gnd DFFSR_2/S FILL
XFILL_6_NAND2X1_178 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_3_INVX1_315 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_23_DFFPOSX1_5 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_0_BUFX2_21 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_22_DFFPOSX1_8 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_9_DFFSR_158 BUFX2_43/A DFFSR_23/S FILL
XNAND2X1_214 INVX1_256/A AND2X2_6/B BUFX2_35/A INVX1_248/A DFFSR_97/S NAND2X1
XFILL_4_OAI21X1_160 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_50_DFFSR_189 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_26_DFFSR_83 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_37_DFFSR_43 INVX1_94/gnd DFFSR_25/S FILL
XFILL_34_1_0 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_9_DFFSR_90 INVX1_2/gnd DFFSR_1/S FILL
XFILL_2_INVX1_135 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_32_3_1 INVX1_8/gnd DFFSR_5/S FILL
XFILL_10_DFFSR_33 INVX1_94/gnd DFFSR_52/S FILL
XFILL_4_NAND2X1_274 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_0_INVX1_352 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_30_5_2 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_43_DFFSR_119 BUFX2_37/A DFFSR_81/S FILL
XFILL_5_NAND2X1_208 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_2_OAI21X1_256 INVX1_2/gnd DFFSR_51/S FILL
XFILL_45_DFFSR_50 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_12_XNOR2X1_1 BUFX2_35/A DFFSR_14/S FILL
XFILL_33_DFFSR_122 INVX1_94/gnd DFFSR_52/S FILL
XFILL_34_DFFSR_90 INVX1_2/gnd DFFSR_1/S FILL
XFILL_23_DFFSR_125 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_4_NAND3X1_106 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_13_DFFSR_128 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_1_DFFSR_47 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_18_DFFSR_40 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_3_OAI21X1_190 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_3_AOI21X1_7 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_6_NAND2X1_142 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_3_INVX1_279 INVX1_4/gnd DFFSR_51/S FILL
XFILL_6_DFFSR_5 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_42_DFFSR_97 BUFX2_35/A DFFSR_97/S FILL
XFILL_9_DFFSR_122 INVX1_94/gnd DFFSR_52/S FILL
XNAND2X1_178 AND2X2_8/A AND2X2_6/A BUFX2_8/gnd NOR2X1_3/A DFFSR_25/S NAND2X1
XFILL_3_AND2X2_6 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_50_DFFSR_153 BUFX2_36/A DFFSR_8/S FILL
XFILL_4_OAI21X1_124 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_40_DFFSR_156 INVX1_23/gnd DFFSR_91/S FILL
XFILL_9_DFFSR_54 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_26_DFFSR_47 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_15_DFFSR_87 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_30_DFFSR_159 BUFX2_36/A DFFSR_6/S FILL
XFILL_20_DFFSR_162 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_4_NAND2X1_238 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_40_0_2 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_10_DFFSR_165 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_5_NAND3X1_6 INVX1_8/gnd DFFSR_7/S FILL
XFILL_0_INVX1_316 BUFX2_37/A DFFSR_8/S FILL
XFILL_5_NOR2X1_41 BUFX2_8/gnd DFFSR_10/S FILL
XINVX1_426 DFFSR_140/Q BUFX2_17/gnd INVX1_426/Y DFFSR_57/S INVX1
XFILL_30_DFFSR_9 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_4_INVX1_423 BUFX2_37/A DFFSR_8/S FILL
XFILL_45_DFFSR_14 BUFX2_35/A DFFSR_14/S FILL
XFILL_2_OAI21X1_220 BUFX2_43/A DFFSR_97/S FILL
XFILL_6_DFFSR_159 BUFX2_36/A DFFSR_6/S FILL
XFILL_5_NAND2X1_172 BUFX2_36/A DFFSR_6/S FILL
XFILL_34_DFFSR_54 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_8_DFFPOSX1_10 INVX1_8/gnd DFFSR_5/S FILL
XFILL_23_DFFSR_94 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_12_DFFPOSX1_2 INVX1_89/gnd DFFSR_36/S FILL
XFILL_47_DFFSR_190 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_1_DFFSR_11 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_11_DFFPOSX1_5 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_5_BUFX2_39 BUFX2_43/A DFFSR_97/S FILL
XFILL_3_OAI21X1_154 BUFX2_37/A DFFSR_8/S FILL
XFILL_10_DFFPOSX1_8 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_17_DFFPOSX1_29 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_3_INVX1_243 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_6_NAND2X1_106 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_51_DFFSR_5 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_42_DFFSR_61 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_3_INVX1_95 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_50_DFFSR_117 INVX1_23/gnd DFFSR_91/S FILL
XFILL_3_NAND2X1_268 BUFX2_37/A DFFSR_8/S FILL
XFILL_27_DFFPOSX1_18 BUFX2_37/A DFFSR_8/S FILL
XFILL_8_AOI21X1_34 INVX1_94/gnd DFFSR_25/S FILL
XNAND2X1_142 DFFSR_36/S NAND2X1_142/B DFFSR_79/gnd OAI21X1_142/C DFFSR_36/S NAND2X1
XFILL_7_AOI21X1_37 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_9_DFFSR_18 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_40_DFFSR_120 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_26_DFFSR_11 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_30_DFFSR_123 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_15_DFFSR_51 INVX1_2/gnd DFFSR_51/S FILL
XFILL_6_AOI21X1_40 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_1_OAI21X1_250 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_20_DFFSR_126 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_4_NAND2X1_202 BUFX2_35/A DFFSR_97/S FILL
XFILL_5_AOI21X1_43 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_10_DFFSR_129 INVX1_2/gnd DFFSR_1/S FILL
XAOI21X1_40 INVX1_397/A INVX1_331/A BUFX2_8/Y DFFSR_3/gnd AOI21X1_40/Y DFFSR_4/S AOI21X1
XFILL_3_NAND3X1_100 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_50_DFFSR_68 BUFX2_35/A DFFSR_14/S FILL
XFILL_0_AOI21X1_8 INVX1_94/gnd DFFSR_52/S FILL
XFILL_4_AOI21X1_46 DFFSR_5/gnd DFFSR_5/S FILL
XINVX1_390 INVX1_390/A BUFX2_17/gnd INVX1_390/Y DFFSR_7/S INVX1
XFILL_0_INVX1_280 INVX1_2/gnd DFFSR_51/S FILL
XFILL_20_2 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_2_OAI21X1_184 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_5_NAND2X1_136 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_6_DFFSR_65 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_6_DFFSR_123 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_12_DFFSR_98 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_34_DFFSR_18 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_23_DFFSR_58 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_47_DFFSR_154 BUFX2_36/A DFFSR_6/S FILL
XFILL_37_DFFSR_157 BUFX2_6/gnd DFFSR_91/S FILL
XBUFX2_43 BUFX2_43/A BUFX2_35/A BUFX2_43/Y DFFSR_97/S BUFX2
XFILL_3_INVX1_207 BUFX2_36/A DFFSR_6/S FILL
XFILL_27_DFFSR_160 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_3_OAI21X1_118 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_8_OAI21X1_82 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_17_DFFSR_3 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_17_DFFSR_163 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_2_NAND3X1_7 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_7_OAI21X1_85 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_3_NAND2X1_232 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_3_INVX1_59 INVX1_94/gnd DFFSR_25/S FILL
XFILL_42_DFFSR_25 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_2_NOR2X1_42 BUFX2_17/gnd DFFSR_57/S FILL
XNAND2X1_106 BUFX2_24/Y DFFSR_98/Q DFFSR_1/gnd OAI21X1_106/C DFFSR_9/S NAND2X1
XFILL_6_OAI21X1_88 INVX1_4/gnd DFFSR_4/S FILL
XFILL_31_DFFSR_65 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_5_OAI21X1_91 BUFX2_43/A DFFSR_97/S FILL
XFILL_1_INVX1_424 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_2_NAND3X1_130 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_1_BUFX2_4 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_15_DFFSR_15 INVX1_8/gnd DFFSR_7/S FILL
XFILL_3_DFFSR_160 BUFX2_17/gnd DFFSR_57/S FILL
XOAI21X1_88 BUFX2_18/Y INVX1_99/Y NAND2X1_88/Y INVX1_4/gnd DFFSR_88/D DFFSR_4/S OAI21X1
XFILL_4_OAI21X1_94 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_44_DFFSR_191 INVX1_23/gnd DFFSR_91/S FILL
XFILL_3_OAI21X1_97 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_1_OAI21X1_214 BUFX2_35/A DFFSR_97/S FILL
XFILL_4_NAND2X1_166 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_4_AOI21X1_10 BUFX2_17/gnd DFFSR_57/S FILL
XINVX1_354 DFFSR_123/Q BUFX2_35/A INVX1_354/Y DFFSR_97/S INVX1
XFILL_0_INVX1_244 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_3_AOI21X1_13 INVX1_8/gnd DFFSR_7/S FILL
XFILL_39_DFFSR_72 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_50_DFFSR_32 INVX1_2/gnd DFFSR_1/S FILL
XFILL_16_DFFPOSX1_23 INVX1_23/gnd DFFSR_91/S FILL
XFILL_2_AOI21X1_16 BUFX2_43/A DFFSR_23/S FILL
XFILL_2_OAI21X1_148 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_5_NAND2X1_100 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_1_AOI21X1_19 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_12_DFFSR_62 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_23_DFFSR_22 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_0_DFFPOSX1_2 INVX1_89/gnd DFFSR_36/S FILL
XFILL_6_DFFSR_29 INVX1_4/gnd DFFSR_4/S FILL
XFILL_41_1_0 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_0_AOI21X1_22 BUFX2_43/A DFFSR_97/S FILL
XFILL_47_DFFSR_118 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_37_DFFSR_121 BUFX2_36/A DFFSR_6/S FILL
XFILL_39_3_1 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_2_NAND2X1_262 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_27_DFFSR_124 INVX1_89/gnd DFFSR_36/S FILL
XFILL_3_INVX1_171 BUFX2_35/A DFFSR_14/S FILL
XFILL_17_DFFSR_127 BUFX2_43/A DFFSR_97/S FILL
XFILL_47_DFFSR_79 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_26_DFFPOSX1_12 INVX1_8/gnd DFFSR_5/S FILL
XFILL_8_OAI21X1_46 BUFX2_37/A DFFSR_81/S FILL
XFILL_7_AOI21X1_6 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_37_5_2 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_3_INVX1_23 INVX1_23/gnd DFFSR_91/S FILL
XFILL_20_DFFSR_69 BUFX2_43/A DFFSR_23/S FILL
XFILL_3_DFFSR_76 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_6_NAND2X1_67 INVX1_2/gnd DFFSR_1/S FILL
XFILL_31_DFFSR_29 INVX1_4/gnd DFFSR_4/S FILL
XFILL_0_OAI21X1_244 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_7_OAI21X1_49 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_3_NAND2X1_196 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_6_OAI21X1_52 INVX1_94/gnd DFFSR_25/S FILL
XFILL_5_NAND2X1_70 DFFSR_5/gnd DFFSR_2/S FILL
XNAND2X1_67 BUFX2_24/Y NAND2X1_67/B INVX1_2/gnd NAND2X1_67/Y DFFSR_1/S NAND2X1
XOAI21X1_52 DFFSR_10/S INVX1_59/Y OAI21X1_52/C INVX1_94/gnd DFFSR_52/D DFFSR_25/S
+ OAI21X1
XFILL_5_OAI21X1_55 INVX1_89/gnd DFFSR_2/S FILL
XFILL_1_INVX1_388 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_4_NAND2X1_73 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_7_XOR2X1_6 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_2_BUFX2_14 BUFX2_37/A DFFSR_81/S FILL
XFILL_3_NAND2X1_76 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_3_DFFSR_124 INVX1_89/gnd DFFSR_36/S FILL
XFILL_42_2 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_4_OAI21X1_58 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_3_OAI21X1_61 BUFX2_36/A DFFSR_8/S FILL
XFILL_10_AOI22X1_2 BUFX2_37/A DFFSR_81/S FILL
XFILL_44_DFFSR_155 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_1_OAI21X1_178 INVX1_94/gnd DFFSR_25/S FILL
XFILL_2_NAND2X1_79 INVX1_89/gnd DFFSR_36/S FILL
XFILL_34_DFFSR_158 BUFX2_43/A DFFSR_23/S FILL
XFILL_1_NAND2X1_82 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_4_NAND2X1_130 INVX1_4/gnd DFFSR_4/S FILL
XFILL_2_OAI21X1_64 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_24_DFFSR_161 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_0_INVX1_208 INVX1_23/gnd DFFSR_186/S FILL
XFILL_28_DFFSR_76 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_0_INVX1_70 BUFX2_19/gnd DFFSR_54/S FILL
XINVX1_318 INVX1_35/A DFFSR_71/gnd INVX1_318/Y DFFSR_45/S INVX1
XFILL_0_NAND2X1_85 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_39_DFFSR_36 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_1_OAI21X1_67 INVX1_2/gnd DFFSR_1/S FILL
XFILL_9_NAND3X1_5 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_14_DFFSR_164 INVX1_89/gnd DFFSR_2/S FILL
XFILL_0_OAI21X1_70 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_4_INVX1_315 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_2_OAI21X1_112 INVX1_4/gnd DFFSR_4/S FILL
XFILL_12_DFFSR_26 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_0_DFFSR_161 DFFSR_89/gnd DFFSR_186/S FILL
XDFFSR_6 DFFSR_6/Q INVX1_1/A DFFSR_6/R DFFSR_6/S DFFSR_6/D BUFX2_5/gnd DFFSR_6/S DFFSR
XFILL_2_NAND2X1_226 BUFX2_36/A DFFSR_6/S FILL
XFILL_5_DFFSR_2 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_51_DFFSR_189 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_47_0_2 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_47_DFFSR_43 INVX1_94/gnd DFFSR_25/S FILL
XFILL_3_INVX1_135 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_36_DFFSR_83 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_8_OAI21X1_10 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_1_NAND3X1_124 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_6_NAND2X1_31 BUFX2_43/A DFFSR_97/S FILL
XFILL_7_OAI21X1_13 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_0_OAI21X1_208 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_20_DFFSR_33 INVX1_94/gnd DFFSR_52/S FILL
XFILL_6_OAI21X1_16 INVX1_89/gnd DFFSR_36/S FILL
XFILL_3_DFFSR_40 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_3_NAND2X1_160 INVX1_8/gnd DFFSR_5/S FILL
XFILL_5_NAND2X1_34 INVX1_2/gnd DFFSR_1/S FILL
XFILL_3_OR2X2_2 BUFX2_6/gnd DFFSR_91/S FILL
XNAND2X1_31 DFFSR_23/S INVX1_26/A BUFX2_43/A OAI21X1_31/C DFFSR_97/S NAND2X1
XFILL_1_INVX1_352 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_4_NAND2X1_37 INVX1_8/gnd DFFSR_5/S FILL
XFILL_5_OAI21X1_19 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_4_OAI21X1_22 BUFX2_8/gnd DFFSR_25/S FILL
XOAI21X1_16 DFFSR_45/S INVX1_18/Y NAND2X1_16/Y INVX1_89/gnd DFFSR_16/D DFFSR_36/S
+ OAI21X1
XFILL_3_NAND2X1_40 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_29_DFFSR_6 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_15_DFFPOSX1_17 BUFX2_37/A DFFSR_8/S FILL
XFILL_44_DFFSR_119 BUFX2_37/A DFFSR_81/S FILL
XFILL_3_OAI21X1_25 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_2_NAND2X1_43 INVX1_89/gnd DFFSR_2/S FILL
XFILL_13_XOR2X1_3 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_9_NAND3X1_99 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_13_XNOR2X1_1 BUFX2_35/A DFFSR_14/S FILL
XFILL_1_OAI21X1_142 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_34_DFFSR_122 INVX1_94/gnd DFFSR_52/S FILL
XFILL_1_NAND2X1_46 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_44_DFFSR_90 INVX1_2/gnd DFFSR_1/S FILL
XFILL_24_DFFSR_125 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_13_1_1 BUFX2_36/A DFFSR_8/S FILL
XFILL_2_OAI21X1_28 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_0_INVX1_172 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_1_OAI21X1_31 BUFX2_35/A DFFSR_97/S FILL
XFILL_14_DFFSR_128 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_0_INVX1_34 INVX1_89/gnd DFFSR_36/S FILL
XFILL_28_DFFSR_40 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_0_DFFSR_87 DFFSR_3/gnd DFFSR_4/S FILL
XINVX1_282 DFFSR_11/Q DFFSR_3/gnd INVX1_282/Y DFFSR_65/S INVX1
XFILL_17_DFFSR_80 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_0_NAND2X1_49 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_11_3_2 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_4_AOI21X1_7 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_1_NAND2X1_256 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_0_OAI21X1_34 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_50_DFFSR_2 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_0_DFFSR_125 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_2_NAND2X1_190 BUFX2_35/A DFFSR_97/S FILL
XFILL_5_DFFPOSX1_28 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_41_DFFSR_156 INVX1_23/gnd DFFSR_91/S FILL
XFILL_5_AOI22X1_12 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_36_DFFSR_47 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_25_DFFSR_87 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_8_DFFSR_94 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_31_DFFSR_159 BUFX2_36/A DFFSR_6/S FILL
XFILL_21_DFFSR_162 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_0_OAI21X1_172 BUFX2_36/A DFFSR_6/S FILL
XFILL_11_DFFSR_165 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_3_NAND2X1_124 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_6_NAND3X1_6 INVX1_8/gnd DFFSR_7/S FILL
XFILL_1_INVX1_316 BUFX2_37/A DFFSR_8/S FILL
XFILL_6_NOR2X1_41 BUFX2_8/gnd DFFSR_10/S FILL
XINVX1_8 INVX1_8/A INVX1_8/gnd INVX1_8/Y DFFSR_5/S INVX1
XFILL_11_OAI22X1_42 INVX1_8/gnd DFFSR_7/S FILL
XFILL_7_DFFSR_159 BUFX2_36/A DFFSR_6/S FILL
XFILL_44_DFFSR_54 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_0_NAND2X1_286 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_10_OAI22X1_45 INVX1_89/gnd DFFSR_2/S FILL
XFILL_1_OAI21X1_106 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_33_DFFSR_94 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_1_NAND2X1_10 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_48_DFFSR_190 DFFSR_9/gnd DFFSR_9/S FILL
XINVX1_246 INVX1_246/A DFFSR_89/gnd NOR2X1_7/B DFFSR_92/S INVX1
XFILL_8_NAND3X1_66 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_0_INVX1_136 BUFX2_43/A DFFSR_97/S FILL
XFILL_9_OAI22X1_48 BUFX2_37/A DFFSR_81/S FILL
XFILL_17_DFFSR_44 BUFX2_8/gnd DFFSR_10/S FILL
XAND2X2_3 AND2X2_3/A AND2X2_3/B BUFX2_17/gnd AND2X2_3/Y DFFSR_57/S AND2X2
XFILL_0_DFFSR_51 INVX1_2/gnd DFFSR_51/S FILL
XFILL_0_NAND2X1_13 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_7_NAND3X1_69 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_8_OAI22X1_51 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_1_NAND2X1_220 BUFX2_35/A DFFSR_14/S FILL
XFILL_6_NAND3X1_72 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_7_OAI22X1_54 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_4_INVX1_243 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_5_NAND3X1_75 BUFX2_35/A DFFSR_97/S FILL
XFILL_0_NAND3X1_118 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_6_OAI22X1_57 BUFX2_17/gnd DFFSR_57/S FILL
XNAND3X1_72 NAND3X1_71/Y NAND3X1_70/Y NAND3X1_72/C BUFX2_5/gnd XOR2X1_8/A DFFSR_23/S
+ NAND3X1
XFILL_4_NAND3X1_78 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_5_OAI22X1_60 INVX1_8/gnd DFFSR_5/S FILL
XFILL_2_NAND2X1_154 BUFX2_37/A DFFSR_8/S FILL
XFILL_3_NAND3X1_81 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_4_OAI22X1_63 BUFX2_8/gnd DFFSR_10/S FILL
XOAI22X1_57 INVX1_372/Y OAI22X1_38/D INVX1_373/Y OAI22X1_49/D BUFX2_17/gnd NOR2X1_38/B
+ DFFSR_57/S OAI22X1
XFILL_2_NAND3X1_84 INVX1_94/gnd DFFSR_25/S FILL
XFILL_3_OAI22X1_66 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_8_OAI21X1_257 INVX1_2/gnd DFFSR_51/S FILL
XFILL_8_DFFSR_58 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_41_DFFSR_120 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_36_DFFSR_11 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_31_DFFSR_123 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_14_DFFSR_91 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_10_XNOR2X1_2 BUFX2_36/A DFFSR_8/S FILL
XFILL_1_NAND3X1_87 INVX1_94/gnd DFFSR_52/S FILL
XFILL_25_DFFSR_51 INVX1_2/gnd DFFSR_51/S FILL
XFILL_0_NAND3X1_90 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_0_BUFX2_1 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_21_DFFSR_126 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_0_OAI21X1_136 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_48_1_0 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_11_DFFSR_129 INVX1_2/gnd DFFSR_1/S FILL
XFILL_14_DFFPOSX1_11 INVX1_4/gnd DFFSR_4/S FILL
XFILL_1_AOI21X1_8 INVX1_94/gnd DFFSR_52/S FILL
XFILL_1_INVX1_280 INVX1_2/gnd DFFSR_51/S FILL
XINVX1_92 DFFSR_81/Q BUFX2_19/gnd INVX1_92/Y DFFSR_54/S INVX1
XFILL_0_NAND2X1_250 INVX1_8/gnd DFFSR_5/S FILL
XFILL_46_3_1 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_7_DFFSR_123 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_9_NAND3X1_27 BUFX2_37/A DFFSR_81/S FILL
XFILL_22_DFFSR_98 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_44_DFFSR_18 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_33_DFFSR_58 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_48_DFFSR_154 BUFX2_36/A DFFSR_6/S FILL
XFILL_8_NAND3X1_30 INVX1_94/gnd DFFSR_52/S FILL
XFILL_44_5_2 INVX1_2/gnd DFFSR_51/S FILL
XFILL_9_OAI22X1_12 INVX1_4/gnd DFFSR_51/S FILL
XINVX1_210 DFFSR_175/Q BUFX2_6/gnd INVX1_210/Y DFFSR_91/S INVX1
XFILL_38_DFFSR_157 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_4_BUFX2_43 BUFX2_35/A DFFSR_97/S FILL
XFILL_7_NAND3X1_33 INVX1_8/gnd DFFSR_7/S FILL
XFILL_0_DFFSR_15 INVX1_8/gnd DFFSR_7/S FILL
XFILL_8_OAI22X1_15 INVX1_4/gnd DFFSR_4/S FILL
XFILL_0_INVX1_100 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_6_NAND3X1_36 BUFX2_35/A DFFSR_97/S FILL
XFILL_1_NAND2X1_184 BUFX2_37/A DFFSR_8/S FILL
XFILL_7_OAI22X1_18 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_28_DFFSR_160 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_4_DFFPOSX1_22 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_18_DFFSR_163 DFFSR_3/gnd DFFSR_65/S FILL
XNAND3X1_36 INVX1_239/A NAND3X1_36/B NAND3X1_36/C BUFX2_35/A AOI22X1_7/B DFFSR_97/S
+ NAND3X1
XFILL_5_NAND3X1_39 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_3_NAND3X1_7 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_41_DFFSR_9 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_6_OAI22X1_21 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_4_NAND3X1_42 BUFX2_43/A DFFSR_23/S FILL
XFILL_5_OAI22X1_24 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_3_NOR2X1_42 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_2_INVX1_99 INVX1_4/gnd DFFSR_4/S FILL
XFILL_41_DFFSR_65 DFFSR_3/gnd DFFSR_65/S FILL
XOAI22X1_21 INVX1_298/Y OAI22X1_9/B INVX1_297/Y OAI22X1_9/D DFFSR_73/gnd NOR2X1_20/B
+ DFFSR_11/S OAI22X1
XFILL_8_OAI21X1_221 BUFX2_35/A DFFSR_14/S FILL
XFILL_3_NAND3X1_45 BUFX2_35/A DFFSR_97/S FILL
XFILL_12_4_0 BUFX2_36/A DFFSR_6/S FILL
XFILL_4_OAI22X1_27 DFFSR_79/gnd DFFSR_36/S FILL
XDFFSR_163 DFFSR_163/Q CLKBUF1_10/Y DFFSR_162/R DFFSR_65/S DFFSR_163/D DFFSR_3/gnd
+ DFFSR_65/S DFFSR
XFILL_2_INVX1_424 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_2_NAND2X1_118 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_2_NAND3X1_48 BUFX2_43/A DFFSR_23/S FILL
XFILL_3_OAI22X1_30 INVX1_94/gnd DFFSR_25/S FILL
XFILL_8_DFFSR_22 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_14_DFFSR_55 INVX1_89/gnd DFFSR_36/S FILL
XFILL_25_DFFSR_15 INVX1_8/gnd DFFSR_7/S FILL
XFILL_4_DFFSR_160 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_45_DFFSR_191 INVX1_23/gnd DFFSR_91/S FILL
XFILL_1_NAND3X1_51 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_2_OAI22X1_33 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_0_OAI21X1_100 INVX1_23/gnd DFFSR_91/S FILL
XFILL_0_NAND3X1_54 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_1_OAI22X1_36 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_23_DFFPOSX1_30 BUFX2_43/A DFFSR_97/S FILL
XFILL_0_OAI22X1_39 BUFX2_37/A DFFSR_8/S FILL
XFILL_7_3 BUFX2_35/A DFFSR_14/S FILL
XFILL_1_INVX1_244 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_49_DFFSR_72 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_0_NAND2X1_214 BUFX2_35/A DFFSR_97/S FILL
XFILL_5_DFFSR_69 BUFX2_43/A DFFSR_23/S FILL
XFILL_22_DFFSR_62 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_33_DFFSR_22 BUFX2_8/gnd DFFSR_10/S FILL
XINVX1_56 DFFSR_49/Q DFFSR_73/gnd INVX1_56/Y DFFSR_11/S INVX1
XFILL_48_DFFSR_118 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_38_DFFSR_121 BUFX2_36/A DFFSR_6/S FILL
XINVX1_174 INVX1_174/A INVX1_94/gnd INVX1_174/Y DFFSR_25/S INVX1
XFILL_28_DFFSR_124 INVX1_89/gnd DFFSR_36/S FILL
XFILL_7_OAI21X1_251 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_1_NAND2X1_148 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_4_INVX1_171 BUFX2_35/A DFFSR_14/S FILL
XFILL_18_DFFSR_127 BUFX2_43/A DFFSR_97/S FILL
XFILL_8_AOI21X1_6 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_9_NAND3X1_101 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_30_DFFSR_69 BUFX2_43/A DFFSR_23/S FILL
XFILL_2_INVX1_63 INVX1_2/gnd DFFSR_51/S FILL
XFILL_41_DFFSR_29 INVX1_4/gnd DFFSR_4/S FILL
XDFFSR_127 DFFSR_127/Q CLKBUF1_6/Y DFFSR_123/R DFFSR_97/S DFFSR_127/D BUFX2_43/A DFFSR_97/S
+ DFFSR
XFILL_8_OAI21X1_185 BUFX2_36/A DFFSR_8/S FILL
XFILL_2_NAND3X1_12 INVX1_94/gnd DFFSR_52/S FILL
XFILL_20_1_1 INVX1_94/gnd DFFSR_52/S FILL
XFILL_29_4 INVX1_89/gnd DFFSR_36/S FILL
XFILL_2_INVX1_388 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_1_NAND3X1_15 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_4_DFFSR_124 INVX1_89/gnd DFFSR_36/S FILL
XFILL_14_DFFSR_19 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_2_0_0 INVX1_23/gnd DFFSR_186/S FILL
XFILL_11_AOI22X1_2 BUFX2_37/A DFFSR_81/S FILL
XFILL_45_DFFSR_155 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_0_NAND3X1_18 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_35_DFFSR_158 BUFX2_43/A DFFSR_23/S FILL
XFILL_18_3_2 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_28_DFFSR_3 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_0_2_1 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_25_DFFSR_161 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_1_INVX1_208 INVX1_23/gnd DFFSR_186/S FILL
XFILL_38_DFFSR_76 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_49_DFFSR_36 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_15_DFFSR_164 INVX1_89/gnd DFFSR_2/S FILL
XFILL_3_DFFPOSX1_16 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_0_NAND3X1_8 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_0_NAND2X1_178 BUFX2_8/gnd DFFSR_25/S FILL
XINVX1_20 DFFSR_17/Q INVX1_8/gnd INVX1_20/Y DFFSR_5/S INVX1
XDFFSR_73 DFFSR_73/Q CLKBUF1_4/Y DFFSR_76/R DFFSR_11/S DFFSR_73/D DFFSR_73/gnd DFFSR_11/S
+ DFFSR
XFILL_5_DFFSR_33 INVX1_94/gnd DFFSR_52/S FILL
XFILL_0_NOR2X1_43 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_22_DFFSR_26 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_11_DFFSR_66 INVX1_2/gnd DFFSR_51/S FILL
XFILL_1_DFFSR_161 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_8_NAND3X1_131 BUFX2_7/gnd DFFSR_54/S FILL
XINVX1_138 DFFSR_122/Q INVX1_94/gnd INVX1_138/Y DFFSR_25/S INVX1
XFILL_7_OAI21X1_215 BUFX2_43/A DFFSR_97/S FILL
XFILL_1_NAND2X1_112 INVX1_4/gnd DFFSR_4/S FILL
XFILL_4_INVX1_135 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_46_DFFSR_83 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_30_DFFSR_33 INVX1_94/gnd DFFSR_52/S FILL
XFILL_2_DFFSR_80 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_19_DFFSR_73 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_2_INVX1_27 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_8_OAI21X1_149 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_22_DFFPOSX1_24 BUFX2_43/A DFFSR_23/S FILL
XFILL_2_INVX1_352 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_45_DFFSR_119 BUFX2_37/A DFFSR_81/S FILL
XFILL_1_BUFX2_18 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_14_XNOR2X1_1 BUFX2_35/A DFFSR_14/S FILL
XFILL_35_DFFSR_122 INVX1_94/gnd DFFSR_52/S FILL
XFILL_25_DFFSR_125 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_1_INVX1_172 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_15_DFFSR_128 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_38_DFFSR_40 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_27_DFFSR_80 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_5_AOI21X1_7 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_0_NAND2X1_142 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_11_DFFSR_30 INVX1_89/gnd DFFSR_36/S FILL
XDFFSR_37 INVX1_42/A DFFSR_2/CLK DFFSR_33/R DFFSR_37/S DFFSR_37/D INVX1_89/gnd DFFSR_2/S
+ DFFSR
XFILL_6_OAI21X1_245 DFFSR_5/gnd DFFSR_2/S FILL
XINVX1_102 DFFSR_90/Q DFFSR_1/gnd INVX1_102/Y DFFSR_1/S INVX1
XFILL_1_DFFSR_125 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_34_9 INVX1_8/gnd DFFSR_7/S FILL
XFILL_42_DFFSR_156 INVX1_23/gnd DFFSR_91/S FILL
XFILL_7_OAI21X1_179 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_46_DFFSR_47 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_35_DFFSR_87 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_32_DFFSR_159 BUFX2_36/A DFFSR_6/S FILL
XFILL_22_DFFSR_162 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_2_DFFSR_44 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_19_DFFSR_37 INVX1_89/gnd DFFSR_2/S FILL
XFILL_12_DFFSR_165 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_7_NAND3X1_6 INVX1_8/gnd DFFSR_7/S FILL
XFILL_8_OAI21X1_113 INVX1_23/gnd DFFSR_91/S FILL
XFILL_2_INVX1_316 BUFX2_37/A DFFSR_8/S FILL
XFILL_12_XOR2X1_7 INVX1_23/gnd DFFSR_91/S FILL
XFILL_8_DFFSR_159 BUFX2_36/A DFFSR_6/S FILL
XFILL_2_DFFPOSX1_10 INVX1_8/gnd DFFSR_5/S FILL
XFILL_43_DFFSR_94 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_49_DFFSR_190 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_1_INVX1_136 BUFX2_43/A DFFSR_97/S FILL
XFILL_27_DFFSR_44 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_4_AND2X2_3 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_16_DFFSR_84 BUFX2_43/A DFFSR_23/S FILL
XFILL_7_NAND3X1_125 INVX1_8/gnd DFFSR_5/S FILL
XFILL_19_4_0 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_6_OAI21X1_209 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_11_DFFPOSX1_29 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_0_NAND2X1_106 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_40_DFFSR_6 BUFX2_5/gnd DFFSR_6/S FILL
XOAI21X1_245 DFFSR_7/S INVX1_407/Y OAI21X1_245/C DFFSR_5/gnd DFFSR_177/D DFFSR_2/S
+ OAI21X1
XFILL_21_DFFPOSX1_18 BUFX2_37/A DFFSR_8/S FILL
XFILL_7_OAI21X1_143 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_42_DFFSR_120 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_32_DFFSR_123 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_24_DFFSR_91 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_11_XNOR2X1_2 BUFX2_36/A DFFSR_8/S FILL
XFILL_7_DFFSR_98 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_35_DFFSR_51 INVX1_2/gnd DFFSR_51/S FILL
XFILL_46_DFFSR_11 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_22_DFFSR_126 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_6_BUFX2_36 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_12_DFFSR_129 INVX1_2/gnd DFFSR_1/S FILL
XFILL_11_1 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_2_AOI21X1_8 INVX1_94/gnd DFFSR_52/S FILL
XFILL_2_INVX1_280 INVX1_2/gnd DFFSR_51/S FILL
XFILL_8_DFFSR_123 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_32_DFFSR_98 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_5_OAI21X1_239 INVX1_4/gnd DFFSR_4/S FILL
XFILL_43_DFFSR_58 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_49_DFFSR_154 BUFX2_36/A DFFSR_6/S FILL
XFILL_39_DFFSR_157 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_16_DFFSR_48 INVX1_4/gnd DFFSR_4/S FILL
XFILL_1_INVX1_100 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_29_DFFSR_160 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_6_OAI21X1_173 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_19_DFFSR_163 DFFSR_3/gnd DFFSR_65/S FILL
XNOR2X1_45 NOR2X1_45/A NOR2X1_45/B BUFX2_35/A NOR2X1_45/Y DFFSR_14/S NOR2X1
XFILL_4_NAND3X1_7 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_27_1_1 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_13_CLKBUF1_12 BUFX2_43/A DFFSR_23/S FILL
XFILL_9_0_0 BUFX2_43/A DFFSR_23/S FILL
XFILL_4_NOR2X1_42 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_25_3_2 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_12_CLKBUF1_15 BUFX2_17/gnd DFFSR_7/S FILL
XOAI21X1_209 AOI21X1_13/Y AOI21X1_12/Y INVX1_237/A BUFX2_17/gnd NAND3X1_60/C DFFSR_57/S
+ OAI21X1
XFILL_7_2_1 BUFX2_35/A DFFSR_97/S FILL
XFILL_7_OAI21X1_107 BUFX2_36/A DFFSR_6/S FILL
XFILL_7_DFFSR_62 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_11_CLKBUF1_18 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_13_DFFSR_95 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_24_DFFSR_55 INVX1_89/gnd DFFSR_36/S FILL
XFILL_35_DFFSR_15 INVX1_8/gnd DFFSR_7/S FILL
XFILL_5_DFFSR_160 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_3_INVX1_424 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_46_DFFSR_191 INVX1_23/gnd DFFSR_91/S FILL
XFILL_10_CLKBUF1_21 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_5_4_2 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_9_CLKBUF1_24 INVX1_23/gnd DFFSR_186/S FILL
XFILL_2_INVX1_244 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_7_DFFSR_9 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_6_NAND3X1_119 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_10_DFFPOSX1_23 INVX1_23/gnd DFFSR_91/S FILL
XFILL_32_DFFSR_62 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_43_DFFSR_22 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_5_OAI21X1_203 BUFX2_35/A DFFSR_14/S FILL
XFILL_49_DFFSR_118 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_39_DFFSR_121 BUFX2_36/A DFFSR_6/S FILL
XFILL_16_DFFSR_12 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_29_DFFSR_124 INVX1_89/gnd DFFSR_36/S FILL
XFILL_19_DFFSR_127 BUFX2_43/A DFFSR_97/S FILL
XFILL_6_OAI21X1_137 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_20_DFFPOSX1_12 INVX1_8/gnd DFFSR_5/S FILL
XFILL_40_DFFSR_69 BUFX2_43/A DFFSR_23/S FILL
XFILL_51_DFFSR_29 INVX1_4/gnd DFFSR_4/S FILL
XOAI21X1_173 DFFSR_91/S INVX1_208/Y OAI21X1_173/C BUFX2_6/gnd DFFSR_173/D DFFSR_14/S
+ OAI21X1
XFILL_6_NAND2X1_251 BUFX2_35/A DFFSR_97/S FILL
XFILL_33_1 INVX1_8/gnd DFFSR_5/S FILL
XFILL_3_INVX1_388 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_5_DFFSR_124 INVX1_89/gnd DFFSR_36/S FILL
XFILL_24_DFFSR_19 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_7_DFFSR_26 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_13_DFFSR_59 INVX1_4/gnd DFFSR_51/S FILL
XFILL_46_DFFSR_155 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_6_NOR2X1_7 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_36_DFFSR_158 BUFX2_43/A DFFSR_23/S FILL
XFILL_4_OAI21X1_233 BUFX2_36/A DFFSR_8/S FILL
XFILL_26_DFFSR_161 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_2_INVX1_208 INVX1_23/gnd DFFSR_186/S FILL
XFILL_48_DFFSR_76 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_16_DFFSR_164 INVX1_89/gnd DFFSR_2/S FILL
XFILL_1_NAND3X1_8 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_5_OAI21X1_167 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_4_INVX1_20 INVX1_8/gnd DFFSR_5/S FILL
XFILL_1_NOR2X1_43 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_32_DFFSR_26 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_21_DFFSR_66 INVX1_2/gnd DFFSR_51/S FILL
XFILL_4_DFFSR_73 DFFSR_73/gnd DFFSR_11/S FILL
XNAND3X1_119 INVX1_397/A INVX1_331/Y INVX1_332/Y DFFSR_5/gnd OAI22X1_49/D DFFSR_2/S
+ NAND3X1
XFILL_2_DFFSR_161 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_0_INVX1_425 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_3_BUFX2_11 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_8_XOR2X1_3 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_5_NAND2X1_281 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_6_OAI21X1_101 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_1_CLKBUF1_12 BUFX2_43/A DFFSR_23/S FILL
XFILL_40_DFFSR_33 INVX1_94/gnd DFFSR_52/S FILL
XFILL_1_INVX1_67 INVX1_4/gnd DFFSR_51/S FILL
XFILL_29_DFFSR_73 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_6_NAND2X1_215 BUFX2_43/A DFFSR_23/S FILL
XFILL_3_INVX1_352 BUFX2_5/gnd DFFSR_6/S FILL
XOAI21X1_137 DFFSR_54/S INVX1_155/Y NAND2X1_137/Y BUFX2_19/gnd DFFSR_137/D DFFSR_52/S
+ OAI21X1
XFILL_3_OAI21X1_263 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_0_CLKBUF1_15 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_13_DFFSR_23 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_46_DFFSR_119 BUFX2_37/A DFFSR_81/S FILL
XFILL_5_NAND3X1_113 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_15_XNOR2X1_1 BUFX2_35/A DFFSR_14/S FILL
XNAND2X1_251 NOR2X1_44/A AND2X2_14/B BUFX2_35/A AOI21X1_41/B DFFSR_97/S NAND2X1
XFILL_36_DFFSR_122 INVX1_94/gnd DFFSR_52/S FILL
XFILL_26_DFFSR_125 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_26_4_0 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_4_OAI21X1_197 INVX1_8/gnd DFFSR_7/S FILL
XFILL_18_DFFSR_7 INVX1_8/gnd DFFSR_7/S FILL
XFILL_2_INVX1_172 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_16_DFFSR_128 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_48_DFFSR_40 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_37_DFFSR_80 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_6_AOI21X1_7 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_6_5_0 BUFX2_35/A DFFSR_14/S FILL
XFILL_21_DFFSR_30 INVX1_89/gnd DFFSR_36/S FILL
XFILL_4_DFFSR_37 INVX1_89/gnd DFFSR_2/S FILL
XFILL_10_DFFSR_70 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_2_BUFX2_8 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_5_OAI21X1_131 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_0_INVX1_389 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_2_DFFSR_125 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_38_6 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_43_DFFSR_156 INVX1_23/gnd DFFSR_91/S FILL
XFILL_5_NAND2X1_245 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_45_DFFSR_87 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_39_DFFSR_3 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_33_DFFSR_159 BUFX2_36/A DFFSR_6/S FILL
XFILL_23_DFFSR_162 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_1_DFFSR_84 BUFX2_43/A DFFSR_23/S FILL
XFILL_29_DFFSR_37 INVX1_89/gnd DFFSR_2/S FILL
XFILL_1_INVX1_31 INVX1_2/gnd DFFSR_1/S FILL
XFILL_13_DFFSR_165 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_24_DFFPOSX1_3 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_18_DFFSR_77 INVX1_89/gnd DFFSR_2/S FILL
XFILL_8_NAND3X1_6 INVX1_8/gnd DFFSR_7/S FILL
XOAI21X1_101 BUFX2_16/Y INVX1_114/Y NAND2X1_101/Y BUFX2_17/gnd DFFSR_101/D DFFSR_7/S
+ OAI21X1
XFILL_3_OAI21X1_227 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_9_DFFPOSX1_17 BUFX2_37/A DFFSR_8/S FILL
XFILL_3_INVX1_316 BUFX2_37/A DFFSR_8/S FILL
XFILL_6_NAND2X1_179 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_23_DFFPOSX1_6 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_22_DFFPOSX1_9 BUFX2_37/A DFFSR_8/S FILL
XFILL_0_BUFX2_22 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_9_DFFSR_159 BUFX2_36/A DFFSR_6/S FILL
XFILL_4_OAI21X1_161 INVX1_23/gnd DFFSR_186/S FILL
XNAND2X1_215 AND2X2_6/A AOI22X1_9/B BUFX2_43/A NOR2X1_9/B DFFSR_23/S NAND2X1
XFILL_10_NOR3X1_1 INVX1_94/gnd DFFSR_52/S FILL
XFILL_50_DFFSR_190 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_9_DFFSR_91 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_2_INVX1_136 BUFX2_43/A DFFSR_97/S FILL
XFILL_34_1_1 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_26_DFFSR_84 BUFX2_43/A DFFSR_23/S FILL
XFILL_37_DFFSR_44 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_32_3_2 INVX1_8/gnd DFFSR_5/S FILL
XFILL_4_NAND2X1_275 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_10_DFFSR_34 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_0_INVX1_353 BUFX2_37/A DFFSR_8/S FILL
XFILL_2_OAI21X1_257 INVX1_2/gnd DFFSR_51/S FILL
XFILL_43_DFFSR_120 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_33_DFFSR_123 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_34_DFFSR_91 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_12_XNOR2X1_2 BUFX2_36/A DFFSR_8/S FILL
XFILL_5_NAND2X1_209 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_45_DFFSR_51 INVX1_2/gnd DFFSR_51/S FILL
XFILL_4_NAND3X1_107 BUFX2_43/A DFFSR_97/S FILL
XFILL_23_DFFSR_126 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_18_DFFSR_41 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_13_DFFSR_129 INVX1_2/gnd DFFSR_1/S FILL
XFILL_1_DFFSR_48 INVX1_4/gnd DFFSR_4/S FILL
XFILL_3_OAI21X1_191 BUFX2_37/A DFFSR_8/S FILL
XFILL_3_AOI21X1_8 INVX1_94/gnd DFFSR_52/S FILL
XFILL_6_NAND2X1_143 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_3_INVX1_280 INVX1_2/gnd DFFSR_51/S FILL
XFILL_6_DFFSR_6 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_9_DFFSR_123 DFFSR_89/gnd DFFSR_186/S FILL
XNAND2X1_179 OR2X2_1/B OR2X2_1/A BUFX2_8/gnd NAND3X1_2/B DFFSR_25/S NAND2X1
XFILL_42_DFFSR_98 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_4_OAI21X1_125 BUFX2_35/A DFFSR_14/S FILL
XFILL_50_DFFSR_154 BUFX2_36/A DFFSR_6/S FILL
XFILL_40_DFFSR_157 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_3_AND2X2_7 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_9_DFFSR_55 INVX1_89/gnd DFFSR_36/S FILL
XFILL_26_DFFSR_48 INVX1_4/gnd DFFSR_4/S FILL
XFILL_15_DFFSR_88 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_2_INVX1_100 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_30_DFFSR_160 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_4_NAND2X1_239 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_20_DFFSR_163 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_5_NAND3X1_7 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_10_DFFSR_166 INVX1_4/gnd DFFSR_51/S FILL
XINVX1_427 DFFSR_133/Q DFFSR_71/gnd INVX1_427/Y DFFSR_10/S INVX1
XFILL_0_INVX1_317 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_5_NOR2X1_42 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_2_OAI21X1_221 BUFX2_35/A DFFSR_14/S FILL
XFILL_5_NAND2X1_173 BUFX2_35/A DFFSR_14/S FILL
XFILL_23_DFFSR_95 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_34_DFFSR_55 INVX1_89/gnd DFFSR_36/S FILL
XFILL_45_DFFSR_15 INVX1_8/gnd DFFSR_7/S FILL
XFILL_6_DFFSR_160 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_8_DFFPOSX1_11 INVX1_4/gnd DFFSR_4/S FILL
XFILL_4_INVX1_424 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_47_DFFSR_191 INVX1_23/gnd DFFSR_91/S FILL
XFILL_12_DFFPOSX1_3 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_1_DFFSR_12 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_11_DFFPOSX1_6 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_5_BUFX2_40 BUFX2_35/A DFFSR_14/S FILL
XFILL_17_DFFPOSX1_30 BUFX2_43/A DFFSR_97/S FILL
XFILL_10_DFFPOSX1_9 BUFX2_37/A DFFSR_8/S FILL
XFILL_3_OAI21X1_155 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_6_NAND2X1_107 BUFX2_36/A DFFSR_6/S FILL
XFILL_3_INVX1_244 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_9_AOI21X1_32 BUFX2_43/A DFFSR_23/S FILL
XFILL_42_DFFSR_62 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_3_INVX1_96 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_8_AOI21X1_35 INVX1_94/gnd DFFSR_25/S FILL
XNAND2X1_143 DFFSR_25/S NAND2X1_248/Y BUFX2_8/gnd NAND2X1_143/Y DFFSR_10/S NAND2X1
XFILL_3_NAND2X1_269 INVX1_4/gnd DFFSR_4/S FILL
XFILL_50_DFFSR_118 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_40_DFFSR_121 BUFX2_36/A DFFSR_6/S FILL
XFILL_9_DFFSR_19 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_27_DFFPOSX1_19 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_26_DFFSR_12 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_7_AOI21X1_38 BUFX2_36/A DFFSR_8/S FILL
XFILL_15_DFFSR_52 INVX1_94/gnd DFFSR_52/S FILL
XFILL_30_DFFSR_124 INVX1_89/gnd DFFSR_36/S FILL
XFILL_1_OAI21X1_251 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_6_AOI21X1_41 BUFX2_35/A DFFSR_14/S FILL
XFILL_20_DFFSR_127 BUFX2_43/A DFFSR_97/S FILL
XAOI21X1_41 INVX1_401/Y AOI21X1_41/B AOI21X1_41/C BUFX2_35/A AOI21X1_41/Y DFFSR_14/S
+ AOI21X1
XFILL_4_NAND2X1_203 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_5_AOI21X1_44 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_10_DFFSR_130 INVX1_4/gnd DFFSR_51/S FILL
XFILL_4_AOI21X1_47 BUFX2_43/A DFFSR_23/S FILL
XFILL_50_DFFSR_69 BUFX2_43/A DFFSR_23/S FILL
XFILL_0_AOI21X1_9 INVX1_94/gnd DFFSR_52/S FILL
XFILL_3_NAND3X1_101 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_20_3 BUFX2_19/gnd DFFSR_52/S FILL
XINVX1_391 INVX1_391/A BUFX2_17/gnd INVX1_391/Y DFFSR_7/S INVX1
XFILL_0_INVX1_281 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_2_OAI21X1_185 BUFX2_36/A DFFSR_8/S FILL
XFILL_33_4_0 INVX1_8/gnd DFFSR_7/S FILL
XFILL_4_INVX1_388 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_12_DFFSR_99 BUFX2_35/A DFFSR_97/S FILL
XFILL_5_NAND2X1_137 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_6_DFFSR_124 INVX1_89/gnd DFFSR_36/S FILL
XFILL_34_DFFSR_19 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_6_DFFSR_66 INVX1_2/gnd DFFSR_51/S FILL
XFILL_23_DFFSR_59 INVX1_4/gnd DFFSR_51/S FILL
XFILL_47_DFFSR_155 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_37_DFFSR_158 BUFX2_43/A DFFSR_23/S FILL
XFILL_27_DFFSR_161 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_3_INVX1_208 INVX1_23/gnd DFFSR_186/S FILL
XFILL_3_OAI21X1_119 BUFX2_37/A DFFSR_8/S FILL
XFILL_8_OAI21X1_83 INVX1_94/gnd DFFSR_52/S FILL
XFILL_17_DFFSR_164 INVX1_89/gnd DFFSR_2/S FILL
XFILL_17_DFFSR_4 INVX1_4/gnd DFFSR_4/S FILL
XFILL_2_NAND3X1_8 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_7_OAI21X1_86 INVX1_4/gnd DFFSR_51/S FILL
XFILL_6_OAI21X1_89 BUFX2_35/A DFFSR_14/S FILL
XNAND2X1_107 BUFX2_25/Y DFFSR_99/Q BUFX2_36/A OAI21X1_107/C DFFSR_6/S NAND2X1
XFILL_3_NAND2X1_233 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_3_INVX1_60 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_2_NOR2X1_43 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_42_DFFSR_26 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_31_DFFSR_66 INVX1_2/gnd DFFSR_51/S FILL
XFILL_5_OAI21X1_92 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_3_DFFSR_161 DFFSR_89/gnd DFFSR_186/S FILL
XOAI21X1_89 BUFX2_21/Y INVX1_101/Y OAI21X1_89/C BUFX2_35/A DFFSR_89/D DFFSR_14/S OAI21X1
XFILL_1_BUFX2_5 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_2_NAND3X1_131 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_15_DFFSR_16 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_1_INVX1_425 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_4_OAI21X1_95 INVX1_89/gnd DFFSR_36/S FILL
XFILL_1_OAI21X1_215 BUFX2_43/A DFFSR_97/S FILL
XFILL_3_OAI21X1_98 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_4_NAND2X1_167 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_4_AOI21X1_11 INVX1_8/gnd DFFSR_5/S FILL
XFILL_0_INVX1_245 BUFX2_35/A DFFSR_14/S FILL
XINVX1_355 INVX1_121/A BUFX2_37/A INVX1_355/Y DFFSR_8/S INVX1
XFILL_3_AOI21X1_14 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_50_DFFSR_33 INVX1_94/gnd DFFSR_52/S FILL
XFILL_39_DFFSR_73 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_16_DFFPOSX1_24 BUFX2_43/A DFFSR_23/S FILL
XFILL_2_AOI21X1_17 INVX1_8/gnd DFFSR_5/S FILL
XFILL_2_OAI21X1_149 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_23_DFFSR_23 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_4_INVX1_352 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_1_AOI21X1_20 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_12_DFFSR_63 INVX1_94/gnd DFFSR_52/S FILL
XFILL_0_DFFPOSX1_3 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_6_DFFSR_30 INVX1_89/gnd DFFSR_36/S FILL
XFILL_5_NAND2X1_101 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_41_1_1 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_47_DFFSR_119 BUFX2_37/A DFFSR_81/S FILL
XFILL_0_AOI21X1_23 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_37_DFFSR_122 INVX1_94/gnd DFFSR_52/S FILL
XFILL_39_3_2 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_27_DFFSR_125 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_2_NAND2X1_263 INVX1_2/gnd DFFSR_51/S FILL
XFILL_3_INVX1_172 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_26_DFFPOSX1_13 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_17_DFFSR_128 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_47_DFFSR_80 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_7_AOI21X1_7 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_8_OAI21X1_47 INVX1_89/gnd DFFSR_2/S FILL
XFILL_6_NAND2X1_68 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_31_DFFSR_30 INVX1_89/gnd DFFSR_36/S FILL
XFILL_3_DFFSR_77 INVX1_89/gnd DFFSR_2/S FILL
XFILL_7_OAI21X1_50 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_20_DFFSR_70 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_3_INVX1_24 INVX1_2/gnd DFFSR_51/S FILL
XFILL_5_NAND2X1_71 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_6_OAI21X1_53 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_0_OAI21X1_245 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_3_NAND2X1_197 INVX1_8/gnd DFFSR_5/S FILL
XNAND2X1_68 BUFX2_23/Y NAND2X1_68/B BUFX2_8/gnd OAI21X1_68/C DFFSR_10/S NAND2X1
XFILL_4_NAND2X1_74 INVX1_2/gnd DFFSR_1/S FILL
XFILL_5_OAI21X1_56 INVX1_2/gnd DFFSR_51/S FILL
XFILL_1_INVX1_389 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_3_DFFSR_125 BUFX2_6/gnd DFFSR_91/S FILL
XOAI21X1_53 DFFSR_10/S INVX1_60/Y OAI21X1_53/C DFFSR_71/gnd DFFSR_53/D DFFSR_45/S
+ OAI21X1
XFILL_3_NAND2X1_77 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_4_OAI21X1_59 INVX1_4/gnd DFFSR_51/S FILL
XFILL_42_3 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_2_BUFX2_15 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_7_XOR2X1_7 INVX1_23/gnd DFFSR_91/S FILL
XFILL_44_DFFSR_156 INVX1_23/gnd DFFSR_91/S FILL
XFILL_10_AOI22X1_3 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_3_OAI21X1_62 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_1_OAI21X1_179 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_2_NAND2X1_80 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_34_DFFSR_159 BUFX2_36/A DFFSR_6/S FILL
XFILL_1_NAND2X1_83 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_4_NAND2X1_131 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_2_OAI21X1_65 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_24_DFFSR_162 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_0_INVX1_209 BUFX2_43/A DFFSR_23/S FILL
XFILL_1_OAI21X1_68 BUFX2_37/A DFFSR_81/S FILL
XFILL_0_INVX1_71 INVX1_94/gnd DFFSR_25/S FILL
XFILL_39_DFFSR_37 INVX1_89/gnd DFFSR_2/S FILL
XFILL_0_NAND2X1_86 INVX1_4/gnd DFFSR_51/S FILL
XFILL_14_DFFSR_165 BUFX2_6/gnd DFFSR_14/S FILL
XINVX1_319 DFFSR_63/Q INVX1_94/gnd INVX1_319/Y DFFSR_25/S INVX1
XFILL_0_OAI21X1_71 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_28_DFFSR_77 INVX1_89/gnd DFFSR_2/S FILL
XFILL_2_OAI21X1_113 INVX1_23/gnd DFFSR_91/S FILL
XFILL_4_INVX1_316 BUFX2_37/A DFFSR_8/S FILL
XFILL_12_DFFSR_27 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_0_DFFSR_162 DFFSR_89/gnd DFFSR_92/S FILL
XDFFSR_7 INVX1_8/A DFFSR_2/CLK DFFSR_6/R DFFSR_7/S DFFSR_7/D INVX1_8/gnd DFFSR_7/S
+ DFFSR
XFILL_5_DFFSR_3 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_2_NAND2X1_227 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_3_INVX1_136 BUFX2_43/A DFFSR_97/S FILL
XFILL_36_DFFSR_84 BUFX2_43/A DFFSR_23/S FILL
XFILL_47_DFFSR_44 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_1_NAND3X1_125 INVX1_8/gnd DFFSR_5/S FILL
XFILL_8_OAI21X1_11 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_7_OAI21X1_14 BUFX2_43/A DFFSR_23/S FILL
XFILL_6_NAND2X1_32 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_3_NAND2X1_161 INVX1_23/gnd DFFSR_186/S FILL
XFILL_6_OAI21X1_17 INVX1_8/gnd DFFSR_5/S FILL
XFILL_5_NAND2X1_35 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_0_OAI21X1_209 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_3_DFFSR_41 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_20_DFFSR_34 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_5_OAI21X1_20 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_3_OR2X2_3 BUFX2_43/A DFFSR_23/S FILL
XFILL_4_NAND2X1_38 DFFSR_5/gnd DFFSR_5/S FILL
XNAND2X1_32 DFFSR_4/S INVX1_27/A DFFSR_3/gnd NAND2X1_32/Y DFFSR_65/S NAND2X1
XFILL_1_INVX1_353 BUFX2_37/A DFFSR_8/S FILL
XFILL_3_NAND2X1_41 DFFSR_5/gnd DFFSR_5/S FILL
XOAI21X1_17 DFFSR_17/S INVX1_20/Y OAI21X1_17/C INVX1_8/gnd DFFSR_17/D DFFSR_5/S OAI21X1
XFILL_13_XOR2X1_4 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_4_OAI21X1_23 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_29_DFFSR_7 INVX1_8/gnd DFFSR_7/S FILL
XFILL_44_DFFSR_120 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_34_DFFSR_123 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_44_DFFSR_91 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_13_XNOR2X1_2 BUFX2_36/A DFFSR_8/S FILL
XFILL_15_DFFPOSX1_18 BUFX2_37/A DFFSR_8/S FILL
XFILL_1_OAI21X1_143 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_2_NAND2X1_44 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_3_OAI21X1_26 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_13_1_2 BUFX2_36/A DFFSR_8/S FILL
XFILL_1_NAND2X1_47 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_24_DFFSR_126 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_2_OAI21X1_29 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_0_INVX1_173 BUFX2_35/A DFFSR_14/S FILL
XFILL_0_INVX1_35 BUFX2_35/A DFFSR_97/S FILL
XFILL_17_DFFSR_81 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_0_NAND2X1_50 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_28_DFFSR_41 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_14_DFFSR_129 INVX1_2/gnd DFFSR_1/S FILL
XINVX1_283 INVX1_58/A INVX1_4/gnd INVX1_283/Y DFFSR_4/S INVX1
XFILL_0_DFFSR_88 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_1_OAI21X1_32 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_4_AOI21X1_8 INVX1_94/gnd DFFSR_52/S FILL
XFILL_0_OAI21X1_35 INVX1_8/gnd DFFSR_5/S FILL
XFILL_1_NAND2X1_257 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_4_INVX1_280 INVX1_2/gnd DFFSR_51/S FILL
XFILL_50_DFFSR_3 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_6_AOI22X1_10 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_2_NAND2X1_191 BUFX2_37/A DFFSR_8/S FILL
XFILL_0_DFFSR_126 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_5_DFFPOSX1_29 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_5_AOI22X1_13 INVX1_23/gnd DFFSR_186/S FILL
XFILL_41_DFFSR_157 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_8_DFFSR_95 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_36_DFFSR_48 INVX1_4/gnd DFFSR_4/S FILL
XFILL_25_DFFSR_88 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_3_INVX1_100 BUFX2_16/gnd DFFSR_11/S FILL
XAOI22X1_10 AOI22X1_13/A AOI22X1_13/B AOI22X1_10/C AOI22X1_10/D BUFX2_6/gnd AOI22X1_10/Y
+ DFFSR_91/S AOI22X1
XFILL_31_DFFSR_160 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_40_4_0 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_21_DFFSR_163 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_0_OAI21X1_173 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_3_NAND2X1_125 BUFX2_35/A DFFSR_14/S FILL
XFILL_6_NAND3X1_7 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_9_OAI21X1_228 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_11_DFFSR_166 INVX1_4/gnd DFFSR_51/S FILL
XINVX1_9 INVX1_9/A BUFX2_36/A INVX1_9/Y DFFSR_6/S INVX1
XFILL_1_INVX1_317 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_6_NOR2X1_42 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_11_OAI22X1_43 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_1_OAI21X1_107 BUFX2_36/A DFFSR_6/S FILL
XFILL_10_OAI22X1_46 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_33_DFFSR_95 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_44_DFFSR_55 INVX1_89/gnd DFFSR_36/S FILL
XFILL_7_DFFSR_160 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_48_DFFSR_191 INVX1_23/gnd DFFSR_91/S FILL
XFILL_9_NAND3X1_64 BUFX2_35/A DFFSR_14/S FILL
XFILL_1_NAND2X1_11 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_8_NAND3X1_67 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_0_NAND2X1_14 BUFX2_43/A DFFSR_23/S FILL
XFILL_0_INVX1_137 BUFX2_36/A DFFSR_8/S FILL
XAND2X2_4 AND2X2_6/A AND2X2_9/A BUFX2_19/gnd AND2X2_4/Y DFFSR_54/S AND2X2
XFILL_0_DFFSR_52 INVX1_94/gnd DFFSR_52/S FILL
XFILL_9_OAI22X1_49 INVX1_94/gnd DFFSR_25/S FILL
XINVX1_247 AND2X2_9/Y BUFX2_6/gnd INVX1_247/Y DFFSR_91/S INVX1
XFILL_7_NAND3X1_70 BUFX2_35/A DFFSR_14/S FILL
XFILL_8_OAI22X1_52 INVX1_94/gnd DFFSR_25/S FILL
XFILL_17_DFFSR_45 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_1_NAND2X1_221 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_6_NAND3X1_73 BUFX2_43/A DFFSR_23/S FILL
XFILL_4_INVX1_244 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_7_OAI22X1_55 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_5_NAND3X1_76 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_6_OAI22X1_58 BUFX2_17/gnd DFFSR_7/S FILL
XNAND3X1_73 AOI22X1_8/C NAND3X1_73/B AOI22X1_8/D BUFX2_43/A NAND3X1_73/Y DFFSR_23/S
+ NAND3X1
XFILL_4_NAND3X1_79 BUFX2_36/A DFFSR_6/S FILL
XFILL_5_OAI22X1_61 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_0_NAND3X1_119 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_16_DFFSR_1 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_3_NAND3X1_82 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_4_OAI22X1_64 INVX1_94/gnd DFFSR_25/S FILL
XOAI22X1_58 INVX1_374/Y OAI22X1_38/B INVX1_375/Y OAI22X1_40/D BUFX2_17/gnd NOR2X1_38/A
+ DFFSR_7/S OAI22X1
XFILL_51_DFFSR_118 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_41_DFFSR_121 BUFX2_36/A DFFSR_6/S FILL
XFILL_2_NAND2X1_155 BUFX2_37/A DFFSR_81/S FILL
XFILL_2_NAND3X1_85 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_8_OAI21X1_258 INVX1_2/gnd DFFSR_51/S FILL
XFILL_3_OAI22X1_67 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_14_DFFSR_92 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_10_XNOR2X1_3 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_36_DFFSR_12 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_1_NAND3X1_88 INVX1_94/gnd DFFSR_52/S FILL
XFILL_25_DFFSR_52 INVX1_94/gnd DFFSR_52/S FILL
XFILL_31_DFFSR_124 INVX1_89/gnd DFFSR_36/S FILL
XFILL_8_DFFSR_59 INVX1_4/gnd DFFSR_51/S FILL
XFILL_21_DFFSR_127 BUFX2_43/A DFFSR_97/S FILL
XFILL_0_BUFX2_2 BUFX2_43/A DFFSR_23/S FILL
XFILL_0_NAND3X1_91 BUFX2_43/A DFFSR_97/S FILL
XFILL_0_OAI21X1_137 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_14_DFFPOSX1_12 INVX1_8/gnd DFFSR_5/S FILL
XFILL_48_1_1 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_11_DFFSR_130 INVX1_4/gnd DFFSR_51/S FILL
XFILL_1_AOI21X1_9 INVX1_94/gnd DFFSR_52/S FILL
XFILL_1_INVX1_281 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_46_3_2 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_10_OAI22X1_10 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_0_NAND2X1_251 BUFX2_35/A DFFSR_97/S FILL
XFILL_22_DFFSR_99 BUFX2_35/A DFFSR_97/S FILL
XFILL_7_DFFSR_124 INVX1_89/gnd DFFSR_36/S FILL
XFILL_44_DFFSR_19 DFFSR_1/gnd DFFSR_9/S FILL
XINVX1_93 DFFSR_82/Q DFFSR_9/gnd INVX1_93/Y DFFSR_9/S INVX1
XFILL_33_DFFSR_59 INVX1_4/gnd DFFSR_51/S FILL
XFILL_48_DFFSR_155 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_8_NAND3X1_31 INVX1_94/gnd DFFSR_52/S FILL
XFILL_9_OAI22X1_13 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_0_INVX1_101 BUFX2_35/A DFFSR_14/S FILL
XFILL_38_DFFSR_158 BUFX2_43/A DFFSR_23/S FILL
XINVX1_211 BUFX2_7/Y BUFX2_37/A DFFSR_175/R DFFSR_8/S INVX1
XFILL_0_DFFSR_16 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_28_DFFSR_161 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_4_DFFPOSX1_23 INVX1_23/gnd DFFSR_91/S FILL
XFILL_1_NAND2X1_185 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_7_NAND3X1_34 INVX1_2/gnd DFFSR_1/S FILL
XFILL_8_OAI22X1_16 INVX1_4/gnd DFFSR_4/S FILL
XFILL_6_NAND3X1_37 BUFX2_43/A DFFSR_97/S FILL
XFILL_7_OAI22X1_19 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_18_DFFSR_164 INVX1_89/gnd DFFSR_2/S FILL
XNAND3X1_37 INVX1_241/Y NAND3X1_37/B NAND3X1_37/C BUFX2_43/A NAND3X1_37/Y DFFSR_97/S
+ NAND3X1
XFILL_5_NAND3X1_40 BUFX2_43/A DFFSR_23/S FILL
XFILL_14_2_0 BUFX2_37/A DFFSR_8/S FILL
XFILL_3_NAND3X1_8 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_6_OAI22X1_22 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_4_NAND3X1_43 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_5_OAI22X1_25 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_3_NOR2X1_43 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_41_DFFSR_66 INVX1_2/gnd DFFSR_51/S FILL
XOAI22X1_22 INVX1_299/Y OAI22X1_6/B INVX1_300/Y OAI22X1_6/D BUFX2_16/gnd NOR2X1_20/A
+ DFFSR_11/S OAI22X1
XFILL_8_OAI21X1_222 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_3_NAND3X1_46 BUFX2_35/A DFFSR_97/S FILL
XFILL_12_4_1 BUFX2_36/A DFFSR_6/S FILL
XFILL_2_NAND2X1_119 BUFX2_37/A DFFSR_8/S FILL
XFILL_4_OAI22X1_28 INVX1_94/gnd DFFSR_25/S FILL
XDFFSR_164 DFFSR_164/Q CLKBUF1_10/Y DFFSR_162/R DFFSR_2/S DFFSR_164/D INVX1_89/gnd
+ DFFSR_2/S DFFSR
XFILL_4_DFFSR_161 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_8_DFFSR_23 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_2_NAND3X1_49 BUFX2_37/A DFFSR_8/S FILL
XFILL_3_OAI22X1_31 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_25_DFFSR_16 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_2_INVX1_425 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_14_DFFSR_56 INVX1_2/gnd DFFSR_51/S FILL
XFILL_1_NAND3X1_52 BUFX2_36/A DFFSR_8/S FILL
XFILL_2_OAI22X1_34 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_0_NAND3X1_55 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_1_OAI22X1_37 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_0_OAI21X1_101 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_0_OAI22X1_40 BUFX2_37/A DFFSR_8/S FILL
XFILL_23_DFFPOSX1_31 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_7_4 BUFX2_35/A DFFSR_14/S FILL
XFILL_1_INVX1_245 BUFX2_35/A DFFSR_14/S FILL
XFILL_49_DFFSR_73 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_0_NAND2X1_215 BUFX2_43/A DFFSR_23/S FILL
XFILL_33_DFFSR_23 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_22_DFFSR_63 INVX1_94/gnd DFFSR_52/S FILL
XINVX1_57 INVX1_57/A BUFX2_17/gnd INVX1_57/Y DFFSR_57/S INVX1
XFILL_5_DFFSR_70 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_48_DFFSR_119 BUFX2_37/A DFFSR_81/S FILL
XINVX1_175 BUFX2_9/Y INVX1_94/gnd INVX1_175/Y DFFSR_52/S INVX1
XFILL_38_DFFSR_122 INVX1_94/gnd DFFSR_52/S FILL
XFILL_28_DFFSR_125 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_1_NAND2X1_149 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_4_INVX1_172 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_18_DFFSR_128 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_7_OAI21X1_252 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_8_AOI21X1_7 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_2_INVX1_64 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_41_DFFSR_30 INVX1_89/gnd DFFSR_36/S FILL
XFILL_30_DFFSR_70 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_3_NAND3X1_10 BUFX2_7/gnd DFFSR_54/S FILL
XDFFSR_128 DFFSR_128/Q CLKBUF1_1/Y DFFSR_123/R DFFSR_52/S DFFSR_128/D BUFX2_19/gnd
+ DFFSR_52/S DFFSR
XFILL_8_OAI21X1_186 BUFX2_36/A DFFSR_8/S FILL
XFILL_20_1_2 INVX1_94/gnd DFFSR_52/S FILL
XFILL_2_NAND3X1_13 INVX1_94/gnd DFFSR_25/S FILL
XFILL_29_5 INVX1_89/gnd DFFSR_36/S FILL
XFILL_2_INVX1_389 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_14_DFFSR_20 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_4_DFFSR_125 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_1_NAND3X1_16 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_2_0_1 INVX1_23/gnd DFFSR_186/S FILL
XFILL_45_DFFSR_156 INVX1_23/gnd DFFSR_91/S FILL
XFILL_0_NAND3X1_19 INVX1_8/gnd DFFSR_5/S FILL
XFILL_35_DFFSR_159 BUFX2_36/A DFFSR_6/S FILL
XFILL_5_NOR3X1_1 INVX1_94/gnd DFFSR_52/S FILL
XFILL_25_DFFSR_162 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_0_2_2 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_28_DFFSR_4 INVX1_4/gnd DFFSR_4/S FILL
XFILL_15_DFFSR_165 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_1_INVX1_209 BUFX2_43/A DFFSR_23/S FILL
XFILL_49_DFFSR_37 INVX1_89/gnd DFFSR_2/S FILL
XFILL_38_DFFSR_77 INVX1_89/gnd DFFSR_2/S FILL
XFILL_3_DFFPOSX1_17 BUFX2_37/A DFFSR_8/S FILL
XFILL_0_NAND3X1_9 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_0_NAND2X1_179 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_0_NOR2X1_44 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_22_DFFSR_27 DFFSR_1/gnd DFFSR_1/S FILL
XINVX1_21 INVX1_21/A DFFSR_1/gnd INVX1_21/Y DFFSR_9/S INVX1
XFILL_5_DFFSR_34 DFFSR_1/gnd DFFSR_9/S FILL
XDFFSR_74 DFFSR_74/Q CLKBUF1_5/Y DFFSR_76/R DFFSR_9/S DFFSR_74/D DFFSR_9/gnd DFFSR_9/S
+ DFFSR
XFILL_11_DFFSR_67 INVX1_2/gnd DFFSR_51/S FILL
XINVX1_139 DFFSR_123/Q BUFX2_6/gnd INVX1_139/Y DFFSR_91/S INVX1
XFILL_8_NAND3X1_132 INVX1_8/gnd DFFSR_7/S FILL
XFILL_47_4_0 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_1_DFFSR_162 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_1_NAND2X1_113 INVX1_23/gnd DFFSR_91/S FILL
XFILL_7_OAI21X1_216 BUFX2_35/A DFFSR_14/S FILL
XFILL_4_INVX1_136 BUFX2_43/A DFFSR_97/S FILL
XFILL_46_DFFSR_84 BUFX2_43/A DFFSR_23/S FILL
XFILL_2_DFFSR_81 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_2_INVX1_28 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_30_DFFSR_34 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_19_DFFSR_74 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_22_DFFPOSX1_25 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_8_OAI21X1_150 INVX1_94/gnd DFFSR_52/S FILL
XFILL_2_INVX1_353 BUFX2_37/A DFFSR_8/S FILL
XFILL_1_BUFX2_19 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_4_INVX1_2 INVX1_2/gnd DFFSR_51/S FILL
XFILL_45_DFFSR_120 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_35_DFFSR_123 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_14_XNOR2X1_2 BUFX2_36/A DFFSR_8/S FILL
XFILL_25_DFFSR_126 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_1_INVX1_173 BUFX2_35/A DFFSR_14/S FILL
XFILL_27_DFFSR_81 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_38_DFFSR_41 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_15_DFFSR_129 INVX1_2/gnd DFFSR_1/S FILL
XFILL_5_AOI21X1_8 INVX1_94/gnd DFFSR_52/S FILL
XFILL_11_DFFSR_31 BUFX2_35/A DFFSR_97/S FILL
XFILL_0_NAND2X1_143 BUFX2_8/gnd DFFSR_10/S FILL
XDFFSR_38 INVX1_43/A DFFSR_15/CLK DFFSR_33/R DFFSR_57/S DFFSR_38/D DFFSR_73/gnd DFFSR_57/S
+ DFFSR
XFILL_6_OAI21X1_246 DFFSR_9/gnd DFFSR_9/S FILL
XINVX1_103 DFFSR_91/Q BUFX2_43/A INVX1_103/Y DFFSR_97/S INVX1
XFILL_1_DFFSR_126 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_42_DFFSR_157 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_7_OAI21X1_180 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_46_DFFSR_48 INVX1_4/gnd DFFSR_4/S FILL
XFILL_35_DFFSR_88 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_32_DFFSR_160 BUFX2_17/gnd DFFSR_57/S FILL
XAOI22X1_1 BUFX2_12/Y AND2X2_9/A AND2X2_8/A AND2X2_6/A BUFX2_19/gnd AOI22X1_1/Y DFFSR_54/S
+ AOI22X1
XFILL_2_DFFSR_45 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_22_DFFSR_163 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_7_NAND3X1_7 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_19_DFFSR_38 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_12_DFFSR_166 INVX1_4/gnd DFFSR_51/S FILL
XFILL_2_INVX1_317 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_8_OAI21X1_114 INVX1_89/gnd DFFSR_36/S FILL
XFILL_12_XOR2X1_8 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_43_DFFSR_95 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_8_DFFSR_160 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_2_DFFPOSX1_11 INVX1_4/gnd DFFSR_4/S FILL
XFILL_49_DFFSR_191 INVX1_23/gnd DFFSR_91/S FILL
XFILL_1_INVX1_137 BUFX2_36/A DFFSR_8/S FILL
XFILL_4_AND2X2_4 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_21_2_0 INVX1_94/gnd DFFSR_25/S FILL
XFILL_16_DFFSR_85 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_27_DFFSR_45 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_7_NAND3X1_126 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_11_DFFPOSX1_30 BUFX2_43/A DFFSR_97/S FILL
XFILL_0_NAND2X1_107 BUFX2_36/A DFFSR_6/S FILL
XFILL_19_4_1 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_6_OAI21X1_210 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_1_3_0 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_40_DFFSR_7 INVX1_8/gnd DFFSR_7/S FILL
XOAI21X1_246 DFFSR_9/S INVX1_408/Y NAND2X1_257/Y DFFSR_9/gnd DFFSR_178/D DFFSR_9/S
+ OAI21X1
XFILL_42_DFFSR_121 BUFX2_36/A DFFSR_6/S FILL
XFILL_7_OAI21X1_144 INVX1_8/gnd DFFSR_7/S FILL
XFILL_21_DFFPOSX1_19 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_24_DFFSR_92 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_11_XNOR2X1_3 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_46_DFFSR_12 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_7_DFFSR_99 BUFX2_35/A DFFSR_97/S FILL
XFILL_35_DFFSR_52 INVX1_94/gnd DFFSR_52/S FILL
XFILL_32_DFFSR_124 INVX1_89/gnd DFFSR_36/S FILL
XFILL_22_DFFSR_127 BUFX2_43/A DFFSR_97/S FILL
XFILL_11_2 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_6_BUFX2_37 BUFX2_37/A DFFSR_81/S FILL
XFILL_2_AOI21X1_9 INVX1_94/gnd DFFSR_52/S FILL
XFILL_12_DFFSR_130 INVX1_4/gnd DFFSR_51/S FILL
XFILL_2_INVX1_281 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_32_DFFSR_99 BUFX2_35/A DFFSR_97/S FILL
XFILL_8_DFFSR_124 INVX1_89/gnd DFFSR_36/S FILL
XFILL_5_OAI21X1_240 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_43_DFFSR_59 INVX1_4/gnd DFFSR_51/S FILL
XFILL_49_DFFSR_155 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_1_INVX1_101 BUFX2_35/A DFFSR_14/S FILL
XFILL_39_DFFSR_158 BUFX2_43/A DFFSR_23/S FILL
XFILL_16_DFFSR_49 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_29_DFFSR_161 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_6_OAI21X1_174 BUFX2_43/A DFFSR_23/S FILL
XFILL_19_DFFSR_164 INVX1_89/gnd DFFSR_2/S FILL
XFILL_4_NAND3X1_8 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_27_1_2 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_14_CLKBUF1_10 DFFSR_73/gnd DFFSR_57/S FILL
XNOR2X1_46 NOR2X1_46/A INVX1_156/A BUFX2_16/gnd INVX1_424/A DFFSR_65/S NOR2X1
XFILL_9_0_1 BUFX2_43/A DFFSR_23/S FILL
XFILL_4_NOR2X1_43 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_13_CLKBUF1_13 INVX1_4/gnd DFFSR_51/S FILL
XFILL_12_CLKBUF1_16 BUFX2_36/A DFFSR_6/S FILL
XOAI21X1_210 AOI21X1_18/Y INVX1_244/Y AOI21X1_17/Y DFFSR_71/gnd NAND3X1_61/C DFFSR_45/S
+ OAI21X1
XFILL_7_2_2 BUFX2_35/A DFFSR_97/S FILL
XFILL_7_DFFSR_63 INVX1_94/gnd DFFSR_52/S FILL
XFILL_7_OAI21X1_108 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_35_DFFSR_16 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_3_INVX1_425 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_13_DFFSR_96 INVX1_2/gnd DFFSR_1/S FILL
XFILL_11_CLKBUF1_19 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_24_DFFSR_56 INVX1_2/gnd DFFSR_51/S FILL
XFILL_5_DFFSR_161 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_10_CLKBUF1_22 INVX1_94/gnd DFFSR_25/S FILL
XFILL_9_CLKBUF1_25 INVX1_23/gnd DFFSR_186/S FILL
XFILL_2_INVX1_245 BUFX2_35/A DFFSR_14/S FILL
XFILL_6_NAND3X1_120 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_27_DFFSR_1 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_10_DFFPOSX1_24 BUFX2_43/A DFFSR_23/S FILL
XFILL_43_DFFSR_23 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_32_DFFSR_63 INVX1_94/gnd DFFSR_52/S FILL
XFILL_5_OAI21X1_204 BUFX2_36/A DFFSR_6/S FILL
XFILL_49_DFFSR_119 BUFX2_37/A DFFSR_81/S FILL
XFILL_39_DFFSR_122 INVX1_94/gnd DFFSR_52/S FILL
XFILL_29_DFFSR_125 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_16_DFFSR_13 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_20_DFFPOSX1_13 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_19_DFFSR_128 BUFX2_19/gnd DFFSR_52/S FILL
XXNOR2X1_1 XNOR2X1_1/A AND2X2_11/Y BUFX2_35/A XNOR2X1_1/Y DFFSR_14/S XNOR2X1
XNOR2X1_10 NOR2X1_10/A NOR2X1_10/B BUFX2_36/A NOR2X1_10/Y DFFSR_6/S NOR2X1
XFILL_9_AOI21X1_7 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_6_OAI21X1_138 DFFSR_73/gnd DFFSR_57/S FILL
XOAI21X1_174 DFFSR_6/S INVX1_209/Y NAND2X1_174/Y BUFX2_43/A DFFSR_174/D DFFSR_23/S
+ OAI21X1
XFILL_40_DFFSR_70 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_6_NAND2X1_252 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_33_2 INVX1_8/gnd DFFSR_5/S FILL
XFILL_3_INVX1_389 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_24_DFFSR_20 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_5_DFFSR_125 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_13_DFFSR_60 BUFX2_37/A DFFSR_8/S FILL
XFILL_7_DFFSR_27 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_46_DFFSR_156 INVX1_23/gnd DFFSR_91/S FILL
XFILL_4_OAI21X1_234 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_6_NOR2X1_8 BUFX2_43/A DFFSR_23/S FILL
XFILL_36_DFFSR_159 BUFX2_36/A DFFSR_6/S FILL
XFILL_26_DFFSR_162 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_16_DFFSR_165 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_2_INVX1_209 BUFX2_43/A DFFSR_23/S FILL
XFILL_48_DFFSR_77 INVX1_89/gnd DFFSR_2/S FILL
XFILL_1_NAND3X1_9 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_1_NOR2X1_44 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_5_OAI21X1_168 BUFX2_36/A DFFSR_6/S FILL
XFILL_32_DFFSR_27 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_4_INVX1_21 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_4_DFFSR_74 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_21_DFFSR_67 INVX1_2/gnd DFFSR_51/S FILL
XNAND3X1_120 INVX1_333/Y INVX1_331/Y INVX1_332/Y DFFSR_5/gnd OAI22X1_52/D DFFSR_5/S
+ NAND3X1
XFILL_0_INVX1_426 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_2_DFFSR_162 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_8_XOR2X1_4 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_3_BUFX2_12 BUFX2_37/A DFFSR_81/S FILL
XFILL_5_NAND2X1_282 INVX1_89/gnd DFFSR_2/S FILL
XFILL_6_OAI21X1_102 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_2_CLKBUF1_10 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_1_INVX1_68 BUFX2_37/A DFFSR_81/S FILL
XFILL_40_DFFSR_34 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_29_DFFSR_74 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_1_CLKBUF1_13 INVX1_4/gnd DFFSR_51/S FILL
XFILL_0_CLKBUF1_16 BUFX2_36/A DFFSR_6/S FILL
XFILL_3_OAI21X1_264 DFFSR_5/gnd DFFSR_5/S FILL
XOAI21X1_138 DFFSR_11/S INVX1_156/Y NAND2X1_138/Y DFFSR_73/gnd DFFSR_138/D DFFSR_57/S
+ OAI21X1
XFILL_6_NAND2X1_216 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_3_INVX1_353 BUFX2_37/A DFFSR_8/S FILL
XFILL_28_2_0 INVX1_89/gnd DFFSR_36/S FILL
XFILL_13_DFFSR_24 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_5_NAND3X1_114 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_46_DFFSR_120 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_36_DFFSR_123 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_15_XNOR2X1_2 BUFX2_36/A DFFSR_8/S FILL
XNAND2X1_252 NOR2X1_1/B NOR2X1_1/A BUFX2_7/gnd NAND2X1_252/Y DFFSR_54/S NAND2X1
XFILL_18_DFFSR_8 BUFX2_36/A DFFSR_8/S FILL
XFILL_26_4_1 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_4_OAI21X1_198 INVX1_8/gnd DFFSR_7/S FILL
XFILL_26_DFFSR_126 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_2_INVX1_173 BUFX2_35/A DFFSR_14/S FILL
XFILL_8_3_0 BUFX2_43/A DFFSR_97/S FILL
XFILL_37_DFFSR_81 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_48_DFFSR_41 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_6_AOI21X1_8 INVX1_94/gnd DFFSR_52/S FILL
XFILL_16_DFFSR_129 INVX1_2/gnd DFFSR_1/S FILL
XFILL_6_5_1 BUFX2_35/A DFFSR_14/S FILL
XFILL_21_DFFSR_31 BUFX2_35/A DFFSR_97/S FILL
XFILL_4_DFFSR_38 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_2_BUFX2_9 BUFX2_37/A DFFSR_8/S FILL
XFILL_10_DFFSR_71 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_5_OAI21X1_132 INVX1_4/gnd DFFSR_4/S FILL
XFILL_0_INVX1_390 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_2_DFFSR_126 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_38_7 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_43_DFFSR_157 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_5_NAND2X1_246 INVX1_94/gnd DFFSR_25/S FILL
XFILL_14_XOR2X1_1 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_39_DFFSR_4 INVX1_4/gnd DFFSR_4/S FILL
XFILL_45_DFFSR_88 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_33_DFFSR_160 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_25_DFFPOSX1_1 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_1_INVX1_32 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_23_DFFSR_163 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_8_NAND3X1_7 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_1_DFFSR_85 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_24_DFFPOSX1_4 BUFX2_17/gnd DFFSR_7/S FILL
XOAI21X1_102 BUFX2_17/Y INVX1_115/Y NAND2X1_102/Y BUFX2_17/gnd DFFSR_102/D DFFSR_57/S
+ OAI21X1
XFILL_29_DFFSR_38 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_18_DFFSR_78 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_13_DFFSR_166 INVX1_4/gnd DFFSR_51/S FILL
XFILL_9_DFFPOSX1_18 BUFX2_37/A DFFSR_8/S FILL
XFILL_6_NAND2X1_180 INVX1_94/gnd DFFSR_52/S FILL
XFILL_3_OAI21X1_228 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_23_DFFPOSX1_7 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_3_INVX1_317 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_0_BUFX2_23 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_50_DFFSR_191 INVX1_23/gnd DFFSR_91/S FILL
XFILL_4_OAI21X1_162 INVX1_23/gnd DFFSR_91/S FILL
XNAND2X1_216 NOR2X1_7/Y OAI21X1_218/C BUFX2_5/gnd AOI22X1_11/B DFFSR_6/S NAND2X1
XFILL_10_NOR3X1_2 INVX1_89/gnd DFFSR_2/S FILL
XFILL_9_DFFSR_160 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_34_1_2 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_9_DFFSR_92 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_2_INVX1_137 BUFX2_36/A DFFSR_8/S FILL
XFILL_26_DFFSR_85 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_37_DFFSR_45 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_4_NAND2X1_276 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_10_DFFSR_35 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_0_INVX1_354 BUFX2_35/A DFFSR_97/S FILL
XFILL_43_DFFSR_121 BUFX2_36/A DFFSR_6/S FILL
XFILL_2_OAI21X1_258 INVX1_2/gnd DFFSR_51/S FILL
XFILL_34_DFFSR_92 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_12_XNOR2X1_3 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_5_NAND2X1_210 BUFX2_35/A DFFSR_97/S FILL
XFILL_45_DFFSR_52 INVX1_94/gnd DFFSR_52/S FILL
XFILL_33_DFFSR_124 INVX1_89/gnd DFFSR_36/S FILL
XFILL_23_DFFSR_127 BUFX2_43/A DFFSR_97/S FILL
XFILL_4_NAND3X1_108 BUFX2_37/A DFFSR_81/S FILL
XFILL_18_DFFSR_42 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_1_DFFSR_49 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_3_OAI21X1_192 BUFX2_37/A DFFSR_81/S FILL
XFILL_3_AOI21X1_9 INVX1_94/gnd DFFSR_52/S FILL
XFILL_13_DFFSR_130 INVX1_4/gnd DFFSR_51/S FILL
XFILL_6_NAND2X1_144 INVX1_8/gnd DFFSR_7/S FILL
XFILL_3_INVX1_281 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_6_DFFSR_7 INVX1_8/gnd DFFSR_7/S FILL
XFILL_42_DFFSR_99 BUFX2_35/A DFFSR_97/S FILL
XNAND2X1_180 AND2X2_11/A INVX1_256/A INVX1_94/gnd INVX1_219/A DFFSR_52/S NAND2X1
XFILL_9_DFFSR_124 INVX1_89/gnd DFFSR_36/S FILL
XFILL_50_DFFSR_155 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_4_OAI21X1_126 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_15_DFFSR_89 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_2_INVX1_101 BUFX2_35/A DFFSR_14/S FILL
XFILL_40_DFFSR_158 BUFX2_43/A DFFSR_23/S FILL
XFILL_3_AND2X2_8 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_9_DFFSR_56 INVX1_2/gnd DFFSR_51/S FILL
XFILL_26_DFFSR_49 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_30_DFFSR_161 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_4_NAND2X1_240 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_20_DFFSR_164 INVX1_89/gnd DFFSR_2/S FILL
XFILL_5_NAND3X1_8 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_10_DFFSR_167 DFFSR_79/gnd DFFSR_36/S FILL
XINVX1_428 INVX1_159/A DFFSR_71/gnd INVX1_428/Y DFFSR_10/S INVX1
XFILL_0_INVX1_318 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_5_NOR2X1_43 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_2_OAI21X1_222 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_13_DFFPOSX1_1 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_5_NAND2X1_174 BUFX2_43/A DFFSR_97/S FILL
XFILL_45_DFFSR_16 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_8_DFFPOSX1_12 INVX1_8/gnd DFFSR_5/S FILL
XFILL_4_INVX1_425 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_23_DFFSR_96 INVX1_2/gnd DFFSR_1/S FILL
XFILL_34_DFFSR_56 INVX1_2/gnd DFFSR_51/S FILL
XFILL_6_DFFSR_161 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_12_DFFPOSX1_4 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_11_DFFPOSX1_7 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_1_DFFSR_13 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_5_BUFX2_41 BUFX2_37/A DFFSR_81/S FILL
XFILL_17_DFFPOSX1_31 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_3_OAI21X1_156 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_3_INVX1_245 BUFX2_35/A DFFSR_14/S FILL
XFILL_6_NAND2X1_108 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_42_DFFSR_63 INVX1_94/gnd DFFSR_52/S FILL
XFILL_3_INVX1_97 INVX1_4/gnd DFFSR_4/S FILL
XFILL_9_AOI21X1_33 BUFX2_35/A DFFSR_14/S FILL
XFILL_50_DFFSR_119 BUFX2_37/A DFFSR_81/S FILL
XFILL_3_NAND2X1_270 BUFX2_19/gnd DFFSR_52/S FILL
XNAND2X1_144 DFFSR_5/S NAND2X1_144/B INVX1_8/gnd NAND2X1_144/Y DFFSR_7/S NAND2X1
XFILL_27_DFFPOSX1_20 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_40_DFFSR_122 INVX1_94/gnd DFFSR_52/S FILL
XFILL_8_AOI21X1_36 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_9_DFFSR_20 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_30_DFFSR_125 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_7_AOI21X1_39 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_15_DFFSR_53 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_26_DFFSR_13 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_6_AOI21X1_42 INVX1_23/gnd DFFSR_91/S FILL
XAOI21X1_42 AOI21X1_42/A AOI21X1_42/B BUFX2_6/Y INVX1_23/gnd AOI21X1_42/Y DFFSR_91/S
+ AOI21X1
XFILL_4_NAND2X1_204 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_20_DFFSR_128 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_5_AOI21X1_45 INVX1_89/gnd DFFSR_36/S FILL
XFILL_1_OAI21X1_252 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_4_AOI21X1_48 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_35_2_0 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_10_DFFSR_131 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_3_NAND3X1_102 INVX1_23/gnd DFFSR_186/S FILL
XFILL_20_4 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_50_DFFSR_70 BUFX2_17/gnd DFFSR_57/S FILL
XINVX1_392 INVX1_392/A DFFSR_3/gnd INVX1_392/Y DFFSR_65/S INVX1
XFILL_0_INVX1_282 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_2_OAI21X1_186 BUFX2_36/A DFFSR_8/S FILL
XFILL_33_4_1 INVX1_8/gnd DFFSR_7/S FILL
XFILL_34_DFFSR_20 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_6_DFFSR_125 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_23_DFFSR_60 BUFX2_37/A DFFSR_8/S FILL
XFILL_6_DFFSR_67 INVX1_2/gnd DFFSR_51/S FILL
XFILL_5_NAND2X1_138 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_47_DFFSR_156 INVX1_23/gnd DFFSR_91/S FILL
XFILL_37_DFFSR_159 BUFX2_36/A DFFSR_6/S FILL
XFILL_27_DFFSR_162 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_9_OAI21X1_81 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_3_OAI21X1_120 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_17_DFFSR_165 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_3_INVX1_209 BUFX2_43/A DFFSR_23/S FILL
XFILL_8_OAI21X1_84 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_17_DFFSR_5 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_2_NAND3X1_9 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_7_OAI21X1_87 INVX1_4/gnd DFFSR_4/S FILL
XFILL_2_NOR2X1_44 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_3_INVX1_61 BUFX2_7/gnd DFFSR_54/S FILL
XNAND2X1_108 BUFX2_23/Y DFFSR_100/Q BUFX2_7/gnd NAND2X1_108/Y DFFSR_54/S NAND2X1
XFILL_42_DFFSR_27 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_31_DFFSR_67 INVX1_2/gnd DFFSR_51/S FILL
XFILL_6_OAI21X1_90 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_3_NAND2X1_234 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_1_BUFX2_6 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_15_DFFSR_17 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_2_NAND3X1_132 INVX1_8/gnd DFFSR_7/S FILL
XFILL_1_INVX1_426 BUFX2_17/gnd DFFSR_57/S FILL
XOAI21X1_90 BUFX2_18/Y INVX1_102/Y NAND2X1_90/Y DFFSR_1/gnd DFFSR_90/D DFFSR_1/S OAI21X1
XFILL_5_OAI21X1_93 INVX1_4/gnd DFFSR_51/S FILL
XFILL_3_DFFSR_162 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_4_OAI21X1_96 INVX1_4/gnd DFFSR_51/S FILL
XFILL_1_OAI21X1_216 BUFX2_35/A DFFSR_14/S FILL
XFILL_3_OAI21X1_99 BUFX2_43/A DFFSR_97/S FILL
XFILL_4_NAND2X1_168 BUFX2_36/A DFFSR_6/S FILL
XFILL_4_AOI21X1_12 INVX1_8/gnd DFFSR_7/S FILL
XFILL_38_DFFSR_1 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_0_INVX1_246 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_3_AOI21X1_15 BUFX2_5/gnd DFFSR_23/S FILL
XINVX1_356 DFFSR_84/Q BUFX2_5/gnd INVX1_356/Y DFFSR_6/S INVX1
XFILL_50_DFFSR_34 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_39_DFFSR_74 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_1_DFFPOSX1_1 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_6_DFFSR_31 BUFX2_35/A DFFSR_97/S FILL
XFILL_16_DFFPOSX1_25 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_2_OAI21X1_150 INVX1_94/gnd DFFSR_52/S FILL
XFILL_2_AOI21X1_18 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_5_NAND2X1_102 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_41_1_2 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_23_DFFSR_24 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_12_DFFSR_64 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_1_AOI21X1_21 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_0_DFFPOSX1_4 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_47_DFFSR_120 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_37_DFFSR_123 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_0_AOI21X1_24 BUFX2_43/A DFFSR_97/S FILL
XFILL_2_NAND2X1_264 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_26_DFFPOSX1_14 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_3_INVX1_173 BUFX2_35/A DFFSR_14/S FILL
XFILL_47_DFFSR_81 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_27_DFFSR_126 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_7_AOI21X1_8 INVX1_94/gnd DFFSR_52/S FILL
XFILL_17_DFFSR_129 INVX1_2/gnd DFFSR_1/S FILL
XFILL_8_OAI21X1_48 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_6_NAND2X1_69 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_3_INVX1_25 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_3_DFFSR_78 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_7_OAI21X1_51 INVX1_2/gnd DFFSR_51/S FILL
XFILL_31_DFFSR_31 BUFX2_35/A DFFSR_97/S FILL
XFILL_6_OAI21X1_54 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_20_DFFSR_71 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_5_NAND2X1_72 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_3_NAND2X1_198 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_0_OAI21X1_246 DFFSR_9/gnd DFFSR_9/S FILL
XNAND2X1_69 BUFX2_23/Y NAND2X1_69/B BUFX2_19/gnd OAI21X1_69/C DFFSR_54/S NAND2X1
XFILL_1_INVX1_390 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_4_NAND2X1_75 INVX1_4/gnd DFFSR_4/S FILL
XFILL_5_OAI21X1_57 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_4_OAI21X1_60 BUFX2_37/A DFFSR_81/S FILL
XOAI21X1_54 DFFSR_54/S INVX1_61/Y OAI21X1_54/C BUFX2_7/gnd DFFSR_54/D DFFSR_54/S OAI21X1
XFILL_3_DFFSR_126 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_42_4 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_2_BUFX2_16 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_3_NAND2X1_78 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_44_DFFSR_157 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_7_XOR2X1_8 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_10_AOI22X1_4 INVX1_94/gnd DFFSR_25/S FILL
XFILL_3_OAI21X1_63 INVX1_94/gnd DFFSR_25/S FILL
XFILL_2_NAND2X1_81 INVX1_94/gnd DFFSR_25/S FILL
XFILL_1_NAND2X1_84 BUFX2_36/A DFFSR_6/S FILL
XFILL_1_OAI21X1_180 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_4_NAND2X1_132 INVX1_8/gnd DFFSR_5/S FILL
XFILL_34_DFFSR_160 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_2_OAI21X1_66 INVX1_4/gnd DFFSR_51/S FILL
XFILL_1_OAI21X1_69 BUFX2_37/A DFFSR_8/S FILL
XFILL_0_NAND2X1_87 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_24_DFFSR_163 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_0_INVX1_210 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_9_NAND3X1_7 BUFX2_7/gnd DFFSR_54/S FILL
XINVX1_320 INVX1_53/A INVX1_89/gnd INVX1_320/Y DFFSR_2/S INVX1
XFILL_0_OAI21X1_72 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_39_DFFSR_38 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_28_DFFSR_78 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_14_DFFSR_166 INVX1_4/gnd DFFSR_51/S FILL
XFILL_0_INVX1_72 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_4_INVX1_317 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_2_OAI21X1_114 INVX1_89/gnd DFFSR_36/S FILL
XFILL_12_DFFSR_28 BUFX2_19/gnd DFFSR_54/S FILL
XDFFSR_8 INVX1_9/A INVX1_1/A DFFSR_6/R DFFSR_8/S DFFSR_8/D BUFX2_36/A DFFSR_8/S DFFSR
XFILL_5_DFFSR_4 INVX1_4/gnd DFFSR_4/S FILL
XFILL_2_NAND2X1_228 INVX1_23/gnd DFFSR_91/S FILL
XFILL_0_DFFSR_163 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_8_OAI21X1_12 BUFX2_35/A DFFSR_14/S FILL
XFILL_3_INVX1_137 BUFX2_36/A DFFSR_8/S FILL
XFILL_36_DFFSR_85 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_47_DFFSR_45 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_6_NAND2X1_33 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_1_NAND3X1_126 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_7_OAI21X1_15 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_0_OAI21X1_210 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_20_DFFSR_35 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_3_DFFSR_42 DFFSR_3/gnd DFFSR_65/S FILL
XNAND2X1_33 DFFSR_25/Q DFFSR_25/S BUFX2_19/gnd OAI21X1_33/C DFFSR_52/S NAND2X1
XFILL_3_NAND2X1_162 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_5_NAND2X1_36 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_6_OAI21X1_18 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_1_INVX1_354 BUFX2_35/A DFFSR_97/S FILL
XFILL_4_NAND2X1_39 DFFSR_71/gnd DFFSR_10/S FILL
XOAI21X1_18 DFFSR_9/S INVX1_21/Y NAND2X1_18/Y DFFSR_9/gnd DFFSR_18/D DFFSR_9/S OAI21X1
XFILL_5_OAI21X1_21 INVX1_2/gnd DFFSR_51/S FILL
XFILL_13_XOR2X1_5 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_44_DFFSR_121 BUFX2_36/A DFFSR_6/S FILL
XFILL_3_NAND2X1_42 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_4_OAI21X1_24 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_44_DFFSR_92 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_13_XNOR2X1_3 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_29_DFFSR_8 BUFX2_36/A DFFSR_8/S FILL
XFILL_2_NAND2X1_45 INVX1_89/gnd DFFSR_36/S FILL
XFILL_34_DFFSR_124 INVX1_89/gnd DFFSR_36/S FILL
XFILL_1_OAI21X1_144 INVX1_8/gnd DFFSR_7/S FILL
XFILL_3_OAI21X1_27 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_15_DFFPOSX1_19 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_2_OAI21X1_30 INVX1_89/gnd DFFSR_36/S FILL
XFILL_1_NAND2X1_48 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_0_DFFSR_89 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_24_DFFSR_127 BUFX2_43/A DFFSR_97/S FILL
XFILL_5_AND2X2_1 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_1_OAI21X1_33 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_0_INVX1_174 INVX1_94/gnd DFFSR_25/S FILL
XINVX1_284 INVX1_22/A DFFSR_1/gnd INVX1_284/Y DFFSR_1/S INVX1
XFILL_17_DFFSR_82 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_0_NAND2X1_51 INVX1_2/gnd DFFSR_51/S FILL
XFILL_0_INVX1_36 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_28_DFFSR_42 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_4_AOI21X1_9 INVX1_94/gnd DFFSR_52/S FILL
XFILL_0_OAI21X1_36 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_1_NAND2X1_258 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_14_DFFSR_130 INVX1_4/gnd DFFSR_51/S FILL
XFILL_50_DFFSR_4 INVX1_4/gnd DFFSR_4/S FILL
XFILL_5_DFFPOSX1_30 BUFX2_43/A DFFSR_97/S FILL
XFILL_0_DFFSR_127 BUFX2_43/A DFFSR_97/S FILL
XFILL_2_NAND2X1_192 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_25_DFFSR_89 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_6_AOI22X1_11 INVX1_23/gnd DFFSR_91/S FILL
XFILL_3_INVX1_101 BUFX2_35/A DFFSR_14/S FILL
XFILL_41_DFFSR_158 BUFX2_43/A DFFSR_23/S FILL
XFILL_8_DFFSR_96 INVX1_2/gnd DFFSR_1/S FILL
XFILL_42_2_0 INVX1_4/gnd DFFSR_4/S FILL
XFILL_36_DFFSR_49 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_31_DFFSR_161 DFFSR_89/gnd DFFSR_186/S FILL
XAOI22X1_11 AOI22X1_11/A AOI22X1_11/B AOI22X1_13/C INVX1_255/A INVX1_23/gnd AOI22X1_11/Y
+ DFFSR_91/S AOI22X1
XFILL_5_AOI22X1_14 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_21_DFFSR_164 INVX1_89/gnd DFFSR_2/S FILL
XFILL_40_4_1 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_0_OAI21X1_174 BUFX2_43/A DFFSR_23/S FILL
XFILL_6_NAND3X1_8 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_9_OAI21X1_229 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_11_DFFSR_167 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_3_NAND2X1_126 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_1_INVX1_318 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_6_NOR2X1_43 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_11_OAI22X1_44 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_10_OAI22X1_47 BUFX2_37/A DFFSR_8/S FILL
XFILL_1_OAI21X1_108 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_33_DFFSR_96 INVX1_2/gnd DFFSR_1/S FILL
XFILL_44_DFFSR_56 INVX1_2/gnd DFFSR_51/S FILL
XFILL_7_DFFSR_161 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_1_NAND2X1_12 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_8_NAND3X1_68 BUFX2_35/A DFFSR_14/S FILL
XAND2X2_5 BUFX2_14/Y AND2X2_5/B BUFX2_37/A AND2X2_5/Y DFFSR_81/S AND2X2
XFILL_9_OAI22X1_50 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_0_NAND2X1_15 BUFX2_17/gnd DFFSR_7/S FILL
XINVX1_248 INVX1_248/A BUFX2_6/gnd INVX1_248/Y DFFSR_14/S INVX1
XFILL_7_NAND3X1_71 BUFX2_35/A DFFSR_14/S FILL
XFILL_17_DFFSR_46 BUFX2_36/A DFFSR_6/S FILL
XFILL_0_INVX1_138 INVX1_94/gnd DFFSR_25/S FILL
XFILL_0_DFFSR_53 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_8_OAI22X1_53 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_1_NAND2X1_222 INVX1_23/gnd DFFSR_186/S FILL
XFILL_6_NAND3X1_74 BUFX2_35/A DFFSR_14/S FILL
XFILL_4_INVX1_245 BUFX2_35/A DFFSR_14/S FILL
XFILL_7_OAI22X1_56 BUFX2_37/A DFFSR_8/S FILL
XFILL_5_NAND3X1_77 BUFX2_37/A DFFSR_81/S FILL
XFILL_6_OAI22X1_59 INVX1_8/gnd DFFSR_7/S FILL
XNAND3X1_74 XNOR2X1_1/Y NAND3X1_70/A NAND3X1_70/C BUFX2_35/A NAND3X1_74/Y DFFSR_14/S
+ NAND3X1
XFILL_4_NAND3X1_80 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_5_OAI22X1_62 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_0_NAND3X1_120 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_3_NAND3X1_83 BUFX2_37/A DFFSR_81/S FILL
XFILL_16_DFFSR_2 DFFSR_5/gnd DFFSR_2/S FILL
XOAI22X1_59 INVX1_377/Y OAI22X1_39/B INVX1_376/Y OAI22X1_39/D INVX1_8/gnd NOR2X1_39/A
+ DFFSR_7/S OAI22X1
XFILL_4_OAI22X1_65 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_8_OAI21X1_259 INVX1_23/gnd DFFSR_186/S FILL
XFILL_2_NAND2X1_156 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_41_DFFSR_122 INVX1_94/gnd DFFSR_52/S FILL
XFILL_8_DFFSR_60 BUFX2_37/A DFFSR_8/S FILL
XFILL_2_NAND3X1_86 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_25_DFFSR_53 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_3_OAI22X1_68 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_10_XNOR2X1_4 INVX1_8/gnd DFFSR_7/S FILL
XFILL_14_DFFSR_93 INVX1_2/gnd DFFSR_51/S FILL
XFILL_36_DFFSR_13 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_31_DFFSR_125 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_1_NAND3X1_89 BUFX2_43/A DFFSR_23/S FILL
XFILL_0_BUFX2_3 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_14_DFFPOSX1_13 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_0_NAND3X1_92 BUFX2_43/A DFFSR_23/S FILL
XFILL_21_DFFSR_128 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_0_OAI21X1_138 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_11_DFFSR_131 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_48_1_2 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_1_INVX1_282 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_10_OAI22X1_11 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_44_DFFSR_20 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_7_DFFSR_125 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_33_DFFSR_60 BUFX2_37/A DFFSR_8/S FILL
XFILL_0_NAND2X1_252 BUFX2_7/gnd DFFSR_54/S FILL
XINVX1_94 DFFSR_83/Q INVX1_94/gnd INVX1_94/Y DFFSR_52/S INVX1
XFILL_48_DFFSR_156 INVX1_23/gnd DFFSR_91/S FILL
XFILL_38_DFFSR_159 BUFX2_36/A DFFSR_6/S FILL
XFILL_17_DFFSR_10 DFFSR_71/gnd DFFSR_10/S FILL
XINVX1_212 BUFX2_3/Y DFFSR_5/gnd NAND3X1_2/A DFFSR_2/S INVX1
XFILL_0_DFFSR_17 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_8_NAND3X1_32 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_0_INVX1_102 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_9_OAI22X1_14 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_28_DFFSR_162 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_7_NAND3X1_35 BUFX2_35/A DFFSR_97/S FILL
XFILL_4_DFFPOSX1_24 BUFX2_43/A DFFSR_23/S FILL
XFILL_1_NAND2X1_186 BUFX2_37/A DFFSR_81/S FILL
XFILL_16_0_0 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_8_OAI22X1_17 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_18_DFFSR_165 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_6_NAND3X1_38 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_7_OAI22X1_20 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_5_NAND3X1_41 BUFX2_43/A DFFSR_23/S FILL
XNAND3X1_38 BUFX2_12/Y AND2X2_10/B NOR2X1_8/A BUFX2_5/gnd NAND3X1_40/B DFFSR_6/S NAND3X1
XFILL_14_2_1 BUFX2_37/A DFFSR_8/S FILL
XFILL_3_NAND3X1_9 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_6_OAI22X1_23 INVX1_89/gnd DFFSR_2/S FILL
XFILL_3_NOR2X1_44 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_4_NAND3X1_44 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_5_OAI22X1_26 INVX1_94/gnd DFFSR_52/S FILL
XFILL_41_DFFSR_67 INVX1_2/gnd DFFSR_51/S FILL
XFILL_8_OAI21X1_223 BUFX2_6/gnd DFFSR_91/S FILL
XDFFSR_165 DFFSR_165/Q CLKBUF1_14/Y DFFSR_162/R DFFSR_14/S DFFSR_165/D BUFX2_6/gnd
+ DFFSR_14/S DFFSR
XFILL_3_NAND3X1_47 BUFX2_43/A DFFSR_97/S FILL
XFILL_12_4_2 BUFX2_36/A DFFSR_6/S FILL
XOAI22X1_23 INVX1_302/Y OAI22X1_7/B INVX1_301/Y OAI22X1_7/D INVX1_89/gnd NOR2X1_21/B
+ DFFSR_2/S OAI22X1
XFILL_4_OAI22X1_29 INVX1_8/gnd DFFSR_5/S FILL
XFILL_2_NAND2X1_120 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_2_NAND3X1_50 BUFX2_37/A DFFSR_81/S FILL
XFILL_3_OAI22X1_32 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_25_DFFSR_17 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_2_INVX1_426 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_14_DFFSR_57 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_8_DFFSR_24 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_4_DFFSR_162 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_1_NAND3X1_53 BUFX2_37/A DFFSR_81/S FILL
XFILL_2_OAI22X1_35 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_0_NAND3X1_56 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_1_OAI22X1_38 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_0_OAI21X1_102 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_0_OAI22X1_41 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_1_INVX1_246 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_49_DFFSR_74 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_7_5 BUFX2_35/A DFFSR_14/S FILL
XFILL_0_NAND2X1_216 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_5_DFFSR_71 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_33_DFFSR_24 BUFX2_16/gnd DFFSR_65/S FILL
XINVX1_58 INVX1_58/A BUFX2_16/gnd INVX1_58/Y DFFSR_65/S INVX1
XFILL_48_DFFSR_120 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_22_DFFSR_64 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_38_DFFSR_123 DFFSR_89/gnd DFFSR_186/S FILL
XINVX1_176 INVX1_176/A BUFX2_37/A INVX1_176/Y DFFSR_81/S INVX1
XFILL_7_OAI21X1_253 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_4_INVX1_173 BUFX2_35/A DFFSR_14/S FILL
XFILL_1_NAND2X1_150 BUFX2_37/A DFFSR_81/S FILL
XFILL_9_XOR2X1_1 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_28_DFFSR_126 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_4_DFFSR_1 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_8_AOI21X1_8 INVX1_94/gnd DFFSR_52/S FILL
XFILL_18_DFFSR_129 INVX1_2/gnd DFFSR_1/S FILL
XFILL_41_DFFSR_31 BUFX2_35/A DFFSR_97/S FILL
XFILL_3_NAND3X1_11 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_30_DFFSR_71 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_2_INVX1_65 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_8_OAI21X1_187 BUFX2_37/A DFFSR_8/S FILL
XFILL_2_INVX1_390 BUFX2_17/gnd DFFSR_7/S FILL
XDFFSR_129 XOR2X1_17/A CLKBUF1_13/Y DFFSR_135/R DFFSR_1/S DFFSR_129/D INVX1_2/gnd
+ DFFSR_1/S DFFSR
XFILL_2_NAND3X1_14 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_4_DFFSR_126 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_14_DFFSR_21 INVX1_2/gnd DFFSR_1/S FILL
XFILL_46_1 INVX1_2/gnd DFFSR_1/S FILL
XFILL_2_0_2 INVX1_23/gnd DFFSR_186/S FILL
XFILL_45_DFFSR_157 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_11_AOI22X1_4 INVX1_94/gnd DFFSR_25/S FILL
XFILL_2_OR2X2_1 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_1_NAND3X1_17 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_0_NAND3X1_20 BUFX2_37/A DFFSR_8/S FILL
XFILL_5_NOR3X1_2 INVX1_89/gnd DFFSR_2/S FILL
XFILL_35_DFFSR_160 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_28_DFFSR_5 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_25_DFFSR_163 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_1_INVX1_210 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_49_DFFSR_38 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_38_DFFSR_78 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_15_DFFSR_166 INVX1_4/gnd DFFSR_51/S FILL
XFILL_3_DFFPOSX1_18 BUFX2_37/A DFFSR_8/S FILL
XFILL_0_NOR2X1_45 BUFX2_35/A DFFSR_14/S FILL
XFILL_11_DFFSR_68 BUFX2_35/A DFFSR_14/S FILL
XFILL_22_DFFSR_28 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_0_NAND2X1_180 INVX1_94/gnd DFFSR_52/S FILL
XFILL_5_DFFSR_35 DFFSR_5/gnd DFFSR_2/S FILL
XINVX1_22 INVX1_22/A DFFSR_1/gnd INVX1_22/Y DFFSR_1/S INVX1
XDFFSR_75 INVX1_85/A CLKBUF1_2/Y DFFSR_76/R DFFSR_51/S DFFSR_75/D INVX1_4/gnd DFFSR_51/S
+ DFFSR
XINVX1_140 INVX1_362/A DFFSR_79/gnd INVX1_140/Y DFFSR_45/S INVX1
XFILL_8_NAND3X1_133 INVX1_8/gnd DFFSR_5/S FILL
XFILL_1_NAND2X1_114 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_47_4_1 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_1_DFFSR_163 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_7_OAI21X1_217 INVX1_23/gnd DFFSR_91/S FILL
XFILL_4_INVX1_137 BUFX2_36/A DFFSR_8/S FILL
XFILL_46_DFFSR_85 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_49_DFFSR_1 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_2_INVX1_29 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_30_DFFSR_35 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_2_DFFSR_82 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_19_DFFSR_75 INVX1_4/gnd DFFSR_51/S FILL
XFILL_22_DFFPOSX1_26 BUFX2_37/A DFFSR_81/S FILL
XFILL_8_OAI21X1_151 BUFX2_37/A DFFSR_81/S FILL
XFILL_2_INVX1_354 BUFX2_35/A DFFSR_97/S FILL
XFILL_1_BUFX2_20 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_45_DFFSR_121 BUFX2_36/A DFFSR_6/S FILL
XFILL_4_INVX1_3 INVX1_8/gnd DFFSR_5/S FILL
XFILL_14_XNOR2X1_3 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_13_5_0 BUFX2_36/A DFFSR_8/S FILL
XFILL_35_DFFSR_124 INVX1_89/gnd DFFSR_36/S FILL
XFILL_25_DFFSR_127 BUFX2_43/A DFFSR_97/S FILL
XFILL_1_INVX1_174 INVX1_94/gnd DFFSR_25/S FILL
XFILL_27_DFFSR_82 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_38_DFFSR_42 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_15_DFFSR_130 INVX1_4/gnd DFFSR_51/S FILL
XFILL_5_AOI21X1_9 INVX1_94/gnd DFFSR_52/S FILL
XDFFSR_39 DFFSR_39/Q DFFSR_52/CLK DFFSR_33/R DFFSR_45/S DFFSR_39/D DFFSR_79/gnd DFFSR_45/S
+ DFFSR
XFILL_0_NAND2X1_144 INVX1_8/gnd DFFSR_7/S FILL
XFILL_6_OAI21X1_247 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_11_DFFSR_32 INVX1_2/gnd DFFSR_1/S FILL
XFILL_1_DFFSR_127 BUFX2_43/A DFFSR_97/S FILL
XINVX1_104 DFFSR_92/Q BUFX2_5/gnd INVX1_104/Y DFFSR_23/S INVX1
XFILL_35_DFFSR_89 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_4_INVX1_101 BUFX2_35/A DFFSR_14/S FILL
XFILL_42_DFFSR_158 BUFX2_43/A DFFSR_23/S FILL
XFILL_7_OAI21X1_181 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_46_DFFSR_49 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_32_DFFSR_161 DFFSR_89/gnd DFFSR_186/S FILL
XAOI22X1_2 BUFX2_12/Y AND2X2_5/B AND2X2_6/A AND2X2_9/A BUFX2_37/A AOI22X1_2/Y DFFSR_81/S
+ AOI22X1
XFILL_22_DFFSR_164 INVX1_89/gnd DFFSR_2/S FILL
XFILL_2_DFFSR_46 BUFX2_36/A DFFSR_6/S FILL
XFILL_7_NAND3X1_8 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_19_DFFSR_39 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_12_DFFSR_167 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_8_OAI21X1_115 BUFX2_36/A DFFSR_6/S FILL
XFILL_2_INVX1_318 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_12_XOR2X1_9 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_23_0_0 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_2_DFFPOSX1_12 INVX1_8/gnd DFFSR_5/S FILL
XFILL_8_DFFSR_161 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_43_DFFSR_96 INVX1_2/gnd DFFSR_1/S FILL
XFILL_4_AND2X2_5 BUFX2_37/A DFFSR_81/S FILL
XFILL_21_2_1 INVX1_94/gnd DFFSR_25/S FILL
XFILL_27_DFFSR_46 BUFX2_36/A DFFSR_6/S FILL
XFILL_1_INVX1_138 INVX1_94/gnd DFFSR_25/S FILL
XFILL_7_NAND3X1_127 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_16_DFFSR_86 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_3_1_0 INVX1_23/gnd DFFSR_91/S FILL
XFILL_11_DFFPOSX1_31 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_0_NAND2X1_108 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_19_4_2 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_6_OAI21X1_211 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_1_3_1 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_40_DFFSR_8 BUFX2_36/A DFFSR_8/S FILL
XFILL_21_DFFPOSX1_20 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_42_DFFSR_122 INVX1_94/gnd DFFSR_52/S FILL
XOAI21X1_247 DFFSR_1/S INVX1_409/Y OAI21X1_247/C DFFSR_1/gnd DFFSR_179/D DFFSR_1/S
+ OAI21X1
XFILL_7_OAI21X1_145 INVX1_23/gnd DFFSR_91/S FILL
XFILL_35_DFFSR_53 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_11_XNOR2X1_4 INVX1_8/gnd DFFSR_7/S FILL
XFILL_24_DFFSR_93 INVX1_2/gnd DFFSR_51/S FILL
XFILL_46_DFFSR_13 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_32_DFFSR_125 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_22_DFFSR_128 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_2_DFFSR_10 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_11_3 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_6_BUFX2_38 BUFX2_37/A DFFSR_81/S FILL
XFILL_12_DFFSR_131 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_2_INVX1_282 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_8_DFFSR_125 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_5_OAI21X1_241 BUFX2_35/A DFFSR_97/S FILL
XFILL_43_DFFSR_60 BUFX2_37/A DFFSR_8/S FILL
XFILL_49_DFFSR_156 INVX1_23/gnd DFFSR_91/S FILL
XFILL_39_DFFSR_159 BUFX2_36/A DFFSR_6/S FILL
XFILL_27_DFFSR_10 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_1_INVX1_102 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_16_DFFSR_50 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_29_DFFSR_162 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_6_OAI21X1_175 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_19_DFFSR_165 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_14_CLKBUF1_11 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_4_NAND3X1_9 BUFX2_19/gnd DFFSR_52/S FILL
XNOR2X1_47 NOR2X1_47/A INVX1_426/Y BUFX2_17/gnd NOR2X1_47/Y DFFSR_57/S NOR2X1
XFILL_4_NOR2X1_44 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_13_CLKBUF1_14 BUFX2_43/A DFFSR_23/S FILL
XFILL_9_0_2 BUFX2_43/A DFFSR_23/S FILL
XFILL_51_DFFSR_67 INVX1_2/gnd DFFSR_51/S FILL
XFILL_12_CLKBUF1_17 INVX1_94/gnd DFFSR_25/S FILL
XOAI21X1_211 NAND3X1_2/A NAND2X1_208/Y NAND3X1_61/Y DFFSR_71/gnd DFFPOSX1_7/D DFFSR_10/S
+ OAI21X1
XFILL_7_OAI21X1_109 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_35_DFFSR_17 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_3_INVX1_426 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_24_DFFSR_57 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_11_CLKBUF1_20 INVX1_4/gnd DFFSR_51/S FILL
XFILL_7_DFFSR_64 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_5_DFFSR_162 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_13_DFFSR_97 BUFX2_35/A DFFSR_97/S FILL
XFILL_10_CLKBUF1_23 INVX1_89/gnd DFFSR_2/S FILL
XFILL_2_INVX1_246 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_27_DFFSR_2 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_6_NAND3X1_121 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_10_DFFPOSX1_25 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_43_DFFSR_24 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_5_OAI21X1_205 BUFX2_36/A DFFSR_8/S FILL
XFILL_49_DFFSR_120 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_32_DFFSR_64 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_39_DFFSR_123 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_16_DFFSR_14 BUFX2_35/A DFFSR_14/S FILL
XFILL_29_DFFSR_126 BUFX2_17/gnd DFFSR_57/S FILL
XNOR2X1_11 OR2X2_2/B OR2X2_2/A BUFX2_6/gnd NOR2X1_11/Y DFFSR_14/S NOR2X1
XFILL_20_DFFPOSX1_14 BUFX2_6/gnd DFFSR_14/S FILL
XXNOR2X1_2 NOR2X1_9/B XNOR2X1_2/B BUFX2_36/A XNOR2X1_2/Y DFFSR_8/S XNOR2X1
XFILL_19_DFFSR_129 INVX1_2/gnd DFFSR_1/S FILL
XFILL_6_OAI21X1_139 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_9_AOI21X1_8 INVX1_94/gnd DFFSR_52/S FILL
XFILL_40_DFFSR_71 DFFSR_71/gnd DFFSR_10/S FILL
XOAI21X1_175 DFFSR_14/S INVX1_210/Y OAI21X1_175/C BUFX2_6/gnd DFFSR_175/D DFFSR_91/S
+ OAI21X1
XFILL_6_NAND2X1_253 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_20_5_0 INVX1_94/gnd DFFSR_52/S FILL
XFILL_33_3 INVX1_8/gnd DFFSR_5/S FILL
XFILL_3_INVX1_390 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_13_DFFSR_61 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_7_DFFSR_28 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_5_DFFSR_126 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_24_DFFSR_21 INVX1_2/gnd DFFSR_1/S FILL
XFILL_46_DFFSR_157 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_6_NOR2X1_9 BUFX2_43/A DFFSR_97/S FILL
XFILL_36_DFFSR_160 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_4_OAI21X1_235 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_26_DFFSR_163 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_2_INVX1_210 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_48_DFFSR_78 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_16_DFFSR_166 INVX1_4/gnd DFFSR_51/S FILL
XFILL_1_NOR2X1_45 BUFX2_35/A DFFSR_14/S FILL
XFILL_21_DFFSR_68 BUFX2_35/A DFFSR_14/S FILL
XFILL_5_OAI21X1_169 BUFX2_36/A DFFSR_8/S FILL
XFILL_32_DFFSR_28 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_4_INVX1_22 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_4_DFFSR_75 INVX1_4/gnd DFFSR_51/S FILL
XFILL_0_INVX1_427 DFFSR_71/gnd DFFSR_10/S FILL
XNAND3X1_121 INVX1_331/A INVX1_333/Y INVX1_332/Y DFFSR_5/gnd OAI22X1_38/D DFFSR_5/S
+ NAND3X1
XFILL_8_XOR2X1_5 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_3_BUFX2_13 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_2_DFFSR_163 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_5_NAND2X1_283 INVX1_89/gnd DFFSR_36/S FILL
XFILL_6_OAI21X1_103 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_2_CLKBUF1_11 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_1_CLKBUF1_14 BUFX2_43/A DFFSR_23/S FILL
XFILL_1_INVX1_69 BUFX2_36/A DFFSR_8/S FILL
XFILL_40_DFFSR_35 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_30_0_0 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_29_DFFSR_75 INVX1_4/gnd DFFSR_51/S FILL
XFILL_3_OAI21X1_265 BUFX2_43/A DFFSR_97/S FILL
XFILL_0_CLKBUF1_17 INVX1_94/gnd DFFSR_25/S FILL
XOAI21X1_139 DFFSR_65/S INVX1_157/Y NAND2X1_139/Y DFFSR_3/gnd DFFSR_139/D DFFSR_65/S
+ OAI21X1
XFILL_3_INVX1_354 BUFX2_35/A DFFSR_97/S FILL
XFILL_6_NAND2X1_217 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_46_DFFSR_121 BUFX2_36/A DFFSR_6/S FILL
XFILL_13_DFFSR_25 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_28_2_1 INVX1_89/gnd DFFSR_36/S FILL
XFILL_15_XNOR2X1_3 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_5_NAND3X1_115 BUFX2_8/gnd DFFSR_10/S FILL
XNAND2X1_253 NOR2X1_2/A NAND2X1_252/Y BUFX2_7/gnd NAND2X1_253/Y DFFSR_54/S NAND2X1
XFILL_26_4_2 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_36_DFFSR_124 INVX1_89/gnd DFFSR_36/S FILL
XFILL_4_OAI21X1_199 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_18_DFFSR_9 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_8_3_1 BUFX2_43/A DFFSR_97/S FILL
XFILL_26_DFFSR_127 BUFX2_43/A DFFSR_97/S FILL
XFILL_2_INVX1_174 INVX1_94/gnd DFFSR_25/S FILL
XFILL_37_DFFSR_82 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_48_DFFSR_42 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_16_DFFSR_130 INVX1_4/gnd DFFSR_51/S FILL
XFILL_6_AOI21X1_9 INVX1_94/gnd DFFSR_52/S FILL
XFILL_4_DFFSR_39 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_6_5_2 BUFX2_35/A DFFSR_14/S FILL
XFILL_5_OAI21X1_133 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_10_DFFSR_72 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_21_DFFSR_32 INVX1_2/gnd DFFSR_1/S FILL
XFILL_0_INVX1_391 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_2_DFFSR_127 BUFX2_43/A DFFSR_97/S FILL
XFILL_45_DFFSR_89 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_43_DFFSR_158 BUFX2_43/A DFFSR_23/S FILL
XFILL_14_XOR2X1_2 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_39_DFFSR_5 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_5_NAND2X1_247 INVX1_8/gnd DFFSR_5/S FILL
XFILL_38_8 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_33_DFFSR_161 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_25_DFFPOSX1_2 INVX1_89/gnd DFFSR_36/S FILL
XFILL_23_DFFSR_164 INVX1_89/gnd DFFSR_2/S FILL
XFILL_8_NAND3X1_8 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_29_DFFSR_39 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_13_DFFSR_167 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_18_DFFSR_79 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_1_DFFSR_86 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_1_INVX1_33 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_24_DFFPOSX1_5 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_6_NAND2X1_181 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_3_OAI21X1_229 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_3_INVX1_318 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_23_DFFPOSX1_8 DFFSR_79/gnd DFFSR_36/S FILL
XOAI21X1_103 BUFX2_22/Y INVX1_116/Y NAND2X1_103/Y DFFSR_5/gnd DFFSR_103/D DFFSR_5/S
+ OAI21X1
XFILL_9_DFFPOSX1_19 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_0_BUFX2_24 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_9_DFFSR_161 DFFSR_89/gnd DFFSR_186/S FILL
XNAND2X1_217 NAND3X1_81/Y NAND3X1_84/Y BUFX2_8/gnd OAI22X1_3/B DFFSR_10/S NAND2X1
XFILL_4_OAI21X1_163 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_37_DFFSR_46 BUFX2_36/A DFFSR_6/S FILL
XFILL_2_INVX1_138 INVX1_94/gnd DFFSR_25/S FILL
XFILL_26_DFFSR_86 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_9_DFFSR_93 INVX1_2/gnd DFFSR_51/S FILL
XFILL_4_NAND2X1_277 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_10_DFFSR_36 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_0_INVX1_355 BUFX2_37/A DFFSR_8/S FILL
XFILL_2_OAI21X1_259 INVX1_23/gnd DFFSR_186/S FILL
XFILL_5_NAND2X1_211 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_43_DFFSR_122 INVX1_94/gnd DFFSR_52/S FILL
XFILL_45_DFFSR_53 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_12_XNOR2X1_4 INVX1_8/gnd DFFSR_7/S FILL
XFILL_34_DFFSR_93 INVX1_2/gnd DFFSR_51/S FILL
XFILL_33_DFFSR_125 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_4_NAND3X1_109 BUFX2_36/A DFFSR_8/S FILL
XFILL_23_DFFSR_128 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_18_DFFSR_43 INVX1_94/gnd DFFSR_25/S FILL
XFILL_1_DFFSR_50 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_3_OAI21X1_193 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_13_DFFSR_131 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_6_NAND2X1_145 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_3_INVX1_282 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_6_DFFSR_8 BUFX2_36/A DFFSR_8/S FILL
XFILL_9_DFFSR_125 BUFX2_6/gnd DFFSR_91/S FILL
XNAND2X1_181 BUFX2_13/Y AND2X2_9/A BUFX2_19/gnd NOR2X1_3/B DFFSR_52/S NAND2X1
XFILL_50_DFFSR_156 INVX1_23/gnd DFFSR_91/S FILL
XFILL_4_OAI21X1_127 BUFX2_43/A DFFSR_23/S FILL
XFILL_3_AND2X2_9 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_40_DFFSR_159 BUFX2_36/A DFFSR_6/S FILL
XFILL_37_DFFSR_10 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_9_DFFSR_57 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_2_INVX1_102 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_15_DFFSR_90 INVX1_2/gnd DFFSR_1/S FILL
XFILL_26_DFFSR_50 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_30_DFFSR_162 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_10_XOR2X1_10 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_20_DFFSR_165 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_10_DFFSR_168 BUFX2_36/A DFFSR_8/S FILL
XFILL_5_NAND3X1_9 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_27_5_0 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_4_NAND2X1_241 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_5_NOR2X1_44 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_0_INVX1_319 INVX1_94/gnd DFFSR_25/S FILL
XINVX1_429 DFFSR_134/Q INVX1_89/gnd NOR2X1_48/A DFFSR_2/S INVX1
XFILL_2_OAI21X1_223 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_8_DFFPOSX1_13 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_5_NAND2X1_175 BUFX2_35/A DFFSR_14/S FILL
XFILL_13_DFFPOSX1_2 INVX1_89/gnd DFFSR_36/S FILL
XFILL_45_DFFSR_17 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_6_DFFSR_162 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_23_DFFSR_97 BUFX2_35/A DFFSR_97/S FILL
XFILL_34_DFFSR_57 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_12_DFFPOSX1_5 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_11_DFFPOSX1_8 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_1_DFFSR_14 BUFX2_35/A DFFSR_14/S FILL
XFILL_5_BUFX2_42 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_3_INVX1_246 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_3_OAI21X1_157 BUFX2_35/A DFFSR_97/S FILL
XFILL_6_NAND2X1_109 INVX1_94/gnd DFFSR_25/S FILL
XFILL_51_DFFSR_8 BUFX2_36/A DFFSR_8/S FILL
XNAND2X1_145 DFFPOSX1_1/Q DFFSR_14/S BUFX2_6/gnd OAI21X1_145/C DFFSR_91/S NAND2X1
XFILL_3_NAND2X1_271 INVX1_89/gnd DFFSR_2/S FILL
XFILL_3_INVX1_98 INVX1_4/gnd DFFSR_4/S FILL
XFILL_50_DFFSR_120 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_42_DFFSR_64 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_27_DFFPOSX1_21 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_8_AOI21X1_37 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_40_DFFSR_123 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_26_DFFSR_14 BUFX2_35/A DFFSR_14/S FILL
XFILL_15_DFFSR_54 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_9_DFFSR_21 INVX1_2/gnd DFFSR_1/S FILL
XFILL_7_AOI21X1_40 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_6_AOI21X1_43 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_30_DFFSR_126 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_37_0_0 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_1_OAI21X1_253 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_4_NAND2X1_205 BUFX2_36/A DFFSR_6/S FILL
XFILL_5_AOI21X1_46 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_20_DFFSR_129 INVX1_2/gnd DFFSR_1/S FILL
XAOI21X1_43 XOR2X1_12/A XOR2X1_12/B AND2X2_15/Y BUFX2_17/gnd XNOR2X1_4/A DFFSR_7/S
+ AOI21X1
XFILL_35_2_1 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_10_DFFSR_132 INVX1_2/gnd DFFSR_51/S FILL
XFILL_3_NAND3X1_103 INVX1_23/gnd DFFSR_186/S FILL
XFILL_20_5 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_50_DFFSR_71 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_0_INVX1_283 INVX1_4/gnd DFFSR_4/S FILL
XINVX1_393 DFFSR_96/Q DFFSR_3/gnd INVX1_393/Y DFFSR_4/S INVX1
XFILL_2_OAI21X1_187 BUFX2_37/A DFFSR_8/S FILL
XFILL_33_4_2 INVX1_8/gnd DFFSR_7/S FILL
XFILL_4_INVX1_390 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_6_DFFSR_68 BUFX2_35/A DFFSR_14/S FILL
XFILL_23_DFFSR_61 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_5_NAND2X1_139 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_6_DFFSR_126 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_34_DFFSR_21 INVX1_2/gnd DFFSR_1/S FILL
XFILL_47_DFFSR_157 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_37_DFFSR_160 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_3_OAI21X1_121 BUFX2_36/A DFFSR_8/S FILL
XFILL_27_DFFSR_163 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_3_INVX1_210 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_9_OAI21X1_82 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_17_DFFSR_166 INVX1_4/gnd DFFSR_51/S FILL
XFILL_17_DFFSR_6 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_8_OAI21X1_85 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_2_NOR2X1_45 BUFX2_35/A DFFSR_14/S FILL
XFILL_31_DFFSR_68 BUFX2_35/A DFFSR_14/S FILL
XFILL_42_DFFSR_28 BUFX2_19/gnd DFFSR_54/S FILL
XNAND2X1_109 BUFX2_19/Y INVX1_368/A INVX1_94/gnd OAI21X1_109/C DFFSR_25/S NAND2X1
XFILL_3_INVX1_62 INVX1_89/gnd DFFSR_2/S FILL
XFILL_7_OAI21X1_88 INVX1_4/gnd DFFSR_4/S FILL
XFILL_6_OAI21X1_91 BUFX2_43/A DFFSR_97/S FILL
XFILL_3_NAND2X1_235 INVX1_4/gnd DFFSR_51/S FILL
XOAI21X1_91 BUFX2_25/Y INVX1_103/Y OAI21X1_91/C BUFX2_43/A DFFSR_91/D DFFSR_97/S OAI21X1
XFILL_1_BUFX2_7 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_1_INVX1_427 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_15_DFFSR_18 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_5_OAI21X1_94 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_4_OAI21X1_97 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_2_NAND3X1_133 INVX1_8/gnd DFFSR_5/S FILL
XFILL_3_DFFSR_163 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_1_OAI21X1_217 INVX1_23/gnd DFFSR_91/S FILL
XFILL_5_AOI21X1_10 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_4_NAND2X1_169 BUFX2_36/A DFFSR_8/S FILL
XFILL_38_DFFSR_2 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_0_INVX1_247 BUFX2_6/gnd DFFSR_91/S FILL
XINVX1_357 DFFSR_76/Q BUFX2_19/gnd INVX1_357/Y DFFSR_52/S INVX1
XFILL_50_DFFSR_35 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_4_AOI21X1_13 INVX1_8/gnd DFFSR_7/S FILL
XFILL_39_DFFSR_75 INVX1_4/gnd DFFSR_51/S FILL
XFILL_3_AOI21X1_16 BUFX2_43/A DFFSR_23/S FILL
XFILL_4_INVX1_354 BUFX2_35/A DFFSR_97/S FILL
XFILL_16_DFFPOSX1_26 BUFX2_37/A DFFSR_81/S FILL
XFILL_2_OAI21X1_151 BUFX2_37/A DFFSR_81/S FILL
XFILL_2_AOI21X1_19 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_1_DFFPOSX1_2 INVX1_89/gnd DFFSR_36/S FILL
XFILL_5_NAND2X1_103 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_6_DFFSR_32 INVX1_2/gnd DFFSR_1/S FILL
XFILL_1_AOI21X1_22 BUFX2_43/A DFFSR_97/S FILL
XFILL_23_DFFSR_25 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_12_DFFSR_65 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_0_DFFPOSX1_5 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_0_AOI21X1_25 BUFX2_43/A DFFSR_97/S FILL
XFILL_47_DFFSR_121 BUFX2_36/A DFFSR_6/S FILL
XFILL_2_NAND2X1_265 DFFSR_89/gnd DFFSR_186/S FILL
XBUFX2_10 rst BUFX2_7/gnd BUFX2_10/Y DFFSR_81/S BUFX2
XFILL_37_DFFSR_124 INVX1_89/gnd DFFSR_36/S FILL
XFILL_26_DFFPOSX1_15 BUFX2_35/A DFFSR_14/S FILL
XFILL_27_DFFSR_127 BUFX2_43/A DFFSR_97/S FILL
XFILL_3_INVX1_174 INVX1_94/gnd DFFSR_25/S FILL
XFILL_47_DFFSR_82 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_17_DFFSR_130 INVX1_4/gnd DFFSR_51/S FILL
XFILL_8_OAI21X1_49 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_7_AOI21X1_9 INVX1_94/gnd DFFSR_52/S FILL
XFILL_7_OAI21X1_52 INVX1_94/gnd DFFSR_25/S FILL
XFILL_6_NAND2X1_70 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_3_INVX1_26 BUFX2_43/A DFFSR_23/S FILL
XFILL_3_NAND2X1_199 BUFX2_36/A DFFSR_8/S FILL
XFILL_3_DFFSR_79 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_6_OAI21X1_55 INVX1_89/gnd DFFSR_2/S FILL
XFILL_20_DFFSR_72 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_0_OAI21X1_247 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_31_DFFSR_32 INVX1_2/gnd DFFSR_1/S FILL
XFILL_5_NAND2X1_73 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_4_NAND2X1_76 BUFX2_19/gnd DFFSR_52/S FILL
XNAND2X1_70 BUFX2_17/Y NAND2X1_70/B DFFSR_5/gnd NAND2X1_70/Y DFFSR_2/S NAND2X1
XFILL_1_INVX1_391 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_5_OAI21X1_58 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_3_DFFSR_127 BUFX2_43/A DFFSR_97/S FILL
XFILL_4_OAI21X1_61 BUFX2_36/A DFFSR_8/S FILL
XFILL_3_NAND2X1_79 INVX1_89/gnd DFFSR_36/S FILL
XOAI21X1_55 DFFSR_5/S INVX1_62/Y OAI21X1_55/C INVX1_89/gnd DFFSR_55/D DFFSR_2/S OAI21X1
XFILL_2_BUFX2_17 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_42_5 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_44_DFFSR_158 BUFX2_43/A DFFSR_23/S FILL
XFILL_10_AOI22X1_5 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_7_XOR2X1_9 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_2_NAND2X1_82 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_3_OAI21X1_64 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_34_DFFSR_161 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_4_NAND2X1_133 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_1_NAND2X1_85 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_1_OAI21X1_181 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_2_OAI21X1_67 INVX1_2/gnd DFFSR_1/S FILL
XFILL_24_DFFSR_164 INVX1_89/gnd DFFSR_2/S FILL
XFILL_0_INVX1_211 BUFX2_37/A DFFSR_8/S FILL
XFILL_0_INVX1_73 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_39_DFFSR_39 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_14_DFFSR_167 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_28_DFFSR_79 DFFSR_79/gnd DFFSR_36/S FILL
XINVX1_321 INVX1_27/A DFFSR_73/gnd INVX1_321/Y DFFSR_57/S INVX1
XFILL_0_NAND2X1_88 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_1_OAI21X1_70 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_2_OAI21X1_115 BUFX2_36/A DFFSR_6/S FILL
XFILL_4_INVX1_318 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_0_OAI21X1_73 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_12_DFFSR_29 INVX1_4/gnd DFFSR_4/S FILL
XFILL_5_DFFSR_5 DFFSR_5/gnd DFFSR_5/S FILL
XDFFSR_9 DFFSR_9/Q DFFSR_1/CLK DFFSR_9/R DFFSR_9/S DFFSR_9/D DFFSR_9/gnd DFFSR_9/S
+ DFFSR
XFILL_2_NAND2X1_229 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_9_OAI21X1_10 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_0_DFFSR_164 INVX1_89/gnd DFFSR_2/S FILL
XFILL_34_5_0 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_47_DFFSR_46 BUFX2_36/A DFFSR_6/S FILL
XFILL_3_INVX1_138 INVX1_94/gnd DFFSR_25/S FILL
XFILL_36_DFFSR_86 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_1_NAND3X1_127 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_8_OAI21X1_13 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_3_DFFSR_43 INVX1_94/gnd DFFSR_25/S FILL
XFILL_0_OAI21X1_211 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_20_DFFSR_36 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_7_OAI21X1_16 INVX1_89/gnd DFFSR_36/S FILL
XFILL_6_NAND2X1_34 INVX1_2/gnd DFFSR_1/S FILL
XFILL_5_NAND2X1_37 INVX1_8/gnd DFFSR_5/S FILL
XFILL_3_NAND2X1_163 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_6_OAI21X1_19 DFFSR_1/gnd DFFSR_1/S FILL
XNAND2X1_34 DFFSR_51/S INVX1_30/A INVX1_2/gnd NAND2X1_34/Y DFFSR_1/S NAND2X1
XFILL_1_INVX1_355 BUFX2_37/A DFFSR_8/S FILL
XFILL_5_OAI21X1_22 BUFX2_8/gnd DFFSR_25/S FILL
XOAI21X1_19 DFFSR_9/S INVX1_22/Y OAI21X1_19/C DFFSR_1/gnd DFFSR_19/D DFFSR_1/S OAI21X1
XFILL_4_NAND2X1_40 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_4_OAI21X1_25 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_3_NAND2X1_43 INVX1_89/gnd DFFSR_2/S FILL
XFILL_13_XOR2X1_6 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_1_OAI21X1_145 INVX1_23/gnd DFFSR_91/S FILL
XFILL_3_OAI21X1_28 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_15_DFFPOSX1_20 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_44_DFFSR_122 INVX1_94/gnd DFFSR_52/S FILL
XFILL_2_NAND2X1_46 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_13_XNOR2X1_4 INVX1_8/gnd DFFSR_7/S FILL
XFILL_29_DFFSR_9 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_44_DFFSR_93 INVX1_2/gnd DFFSR_51/S FILL
XFILL_34_DFFSR_125 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_2_OAI21X1_31 BUFX2_35/A DFFSR_97/S FILL
XFILL_1_NAND2X1_49 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_5_AND2X2_2 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_17_DFFSR_83 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_24_DFFSR_128 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_0_INVX1_37 INVX1_94/gnd DFFSR_52/S FILL
XFILL_0_INVX1_175 INVX1_94/gnd DFFSR_52/S FILL
XFILL_28_DFFSR_43 INVX1_94/gnd DFFSR_25/S FILL
XFILL_0_NAND2X1_52 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_0_DFFSR_90 INVX1_2/gnd DFFSR_1/S FILL
XFILL_1_OAI21X1_34 DFFSR_1/gnd DFFSR_1/S FILL
XINVX1_285 DFFSR_35/Q BUFX2_16/gnd INVX1_285/Y DFFSR_65/S INVX1
XFILL_0_OAI21X1_37 INVX1_89/gnd DFFSR_2/S FILL
XFILL_14_DFFSR_131 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_4_INVX1_282 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_1_NAND2X1_259 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_44_0_0 INVX1_2/gnd DFFSR_51/S FILL
XFILL_2_NAND2X1_193 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_0_DFFSR_128 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_50_DFFSR_5 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_5_DFFPOSX1_31 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_6_AOI22X1_12 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_8_DFFSR_97 BUFX2_35/A DFFSR_97/S FILL
XFILL_41_DFFSR_159 BUFX2_36/A DFFSR_6/S FILL
XFILL_47_DFFSR_10 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_3_INVX1_102 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_42_2_1 INVX1_4/gnd DFFSR_4/S FILL
XFILL_36_DFFSR_50 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_31_DFFSR_162 DFFSR_89/gnd DFFSR_92/S FILL
XAOI22X1_12 AOI22X1_11/A AOI22X1_11/B AOI22X1_10/C AOI22X1_10/D BUFX2_6/gnd OR2X2_2/A
+ DFFSR_91/S AOI22X1
XFILL_25_DFFSR_90 INVX1_2/gnd DFFSR_1/S FILL
XFILL_11_XOR2X1_10 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_21_DFFSR_165 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_40_4_2 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_9_OAI21X1_230 INVX1_23/gnd DFFSR_186/S FILL
XFILL_0_OAI21X1_175 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_3_NAND2X1_127 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_11_DFFSR_168 BUFX2_36/A DFFSR_8/S FILL
XFILL_6_NAND3X1_9 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_6_NOR2X1_44 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_1_INVX1_319 INVX1_94/gnd DFFSR_25/S FILL
XFILL_11_OAI22X1_45 INVX1_89/gnd DFFSR_2/S FILL
XFILL_10_OAI22X1_48 BUFX2_37/A DFFSR_81/S FILL
XFILL_2_NAND2X1_10 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_7_DFFSR_162 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_33_DFFSR_97 BUFX2_35/A DFFSR_97/S FILL
XFILL_1_OAI21X1_109 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_44_DFFSR_57 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_1_NAND2X1_13 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_8_NAND3X1_69 BUFX2_6/gnd DFFSR_14/S FILL
XAND2X2_6 AND2X2_6/A AND2X2_6/B BUFX2_5/gnd AND2X2_6/Y DFFSR_6/S AND2X2
XFILL_9_OAI22X1_51 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_0_NAND2X1_16 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_2_1 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_0_INVX1_139 BUFX2_6/gnd DFFSR_91/S FILL
XINVX1_249 INVX1_249/A BUFX2_35/A INVX1_249/Y DFFSR_14/S INVX1
XFILL_7_NAND3X1_72 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_0_DFFSR_54 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_8_OAI22X1_54 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_17_DFFSR_47 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_4_INVX1_246 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_1_NAND2X1_223 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_6_NAND3X1_75 BUFX2_35/A DFFSR_97/S FILL
XFILL_7_OAI22X1_57 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_5_NAND3X1_78 BUFX2_19/gnd DFFSR_54/S FILL
XNAND3X1_75 NAND3X1_71/B INVX1_245/Y NAND3X1_71/C BUFX2_35/A NAND3X1_75/Y DFFSR_97/S
+ NAND3X1
XFILL_0_NAND3X1_121 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_6_OAI22X1_60 INVX1_8/gnd DFFSR_5/S FILL
XFILL_4_NAND3X1_81 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_5_OAI22X1_63 BUFX2_8/gnd DFFSR_10/S FILL
XOAI22X1_60 INVX1_378/Y OAI22X1_40/B INVX1_379/Y OAI22X1_52/D INVX1_8/gnd NOR2X1_39/B
+ DFFSR_5/S OAI22X1
XFILL_16_DFFSR_3 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_2_NAND2X1_157 BUFX2_35/A DFFSR_97/S FILL
XFILL_3_NAND3X1_84 INVX1_94/gnd DFFSR_25/S FILL
XFILL_4_OAI22X1_66 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_8_OAI21X1_260 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_41_DFFSR_123 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_36_DFFSR_14 BUFX2_35/A DFFSR_14/S FILL
XFILL_8_DFFSR_61 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_25_DFFSR_54 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_2_NAND3X1_87 INVX1_94/gnd DFFSR_52/S FILL
XFILL_14_DFFSR_94 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_1_NAND3X1_90 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_0_BUFX2_4 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_31_DFFSR_126 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_14_DFFPOSX1_14 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_0_NAND3X1_93 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_21_DFFSR_129 INVX1_2/gnd DFFSR_1/S FILL
XFILL_0_OAI21X1_139 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_9_OAI21X1_194 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_11_DFFSR_132 INVX1_2/gnd DFFSR_51/S FILL
XFILL_1_INVX1_283 INVX1_4/gnd DFFSR_4/S FILL
XFILL_33_DFFSR_61 BUFX2_5/gnd DFFSR_6/S FILL
XINVX1_95 DFFSR_84/Q BUFX2_5/gnd INVX1_95/Y DFFSR_6/S INVX1
XFILL_0_NAND2X1_253 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_7_DFFSR_126 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_44_DFFSR_21 INVX1_2/gnd DFFSR_1/S FILL
XFILL_10_OAI22X1_12 INVX1_4/gnd DFFSR_51/S FILL
XFILL_48_DFFSR_157 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_0_INVX1_103 BUFX2_43/A DFFSR_97/S FILL
XINVX1_213 BUFX2_13/Y BUFX2_36/A INVX1_213/Y DFFSR_8/S INVX1
XFILL_8_NAND3X1_33 INVX1_8/gnd DFFSR_7/S FILL
XFILL_38_DFFSR_160 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_0_DFFSR_18 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_9_OAI22X1_15 INVX1_4/gnd DFFSR_4/S FILL
XFILL_17_DFFSR_11 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_7_NAND3X1_36 BUFX2_35/A DFFSR_97/S FILL
XFILL_16_0_1 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_4_DFFPOSX1_25 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_8_OAI22X1_18 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_28_DFFSR_163 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_6_NAND3X1_39 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_1_NAND2X1_187 BUFX2_37/A DFFSR_8/S FILL
XFILL_18_DFFSR_166 INVX1_4/gnd DFFSR_51/S FILL
XFILL_7_OAI22X1_21 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_5_NAND3X1_42 BUFX2_43/A DFFSR_23/S FILL
XFILL_14_2_2 BUFX2_37/A DFFSR_8/S FILL
XFILL_6_OAI22X1_24 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_3_NOR2X1_45 BUFX2_35/A DFFSR_14/S FILL
XFILL_41_DFFSR_68 BUFX2_35/A DFFSR_14/S FILL
XFILL_4_NAND3X1_45 BUFX2_35/A DFFSR_97/S FILL
XNAND3X1_39 AND2X2_6/A AND2X2_6/B NOR2X1_9/A BUFX2_5/gnd NAND3X1_40/C DFFSR_23/S NAND3X1
XFILL_0_AOI22X1_1 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_5_OAI22X1_27 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_3_NAND3X1_48 BUFX2_43/A DFFSR_23/S FILL
XFILL_2_NAND2X1_121 BUFX2_36/A DFFSR_8/S FILL
XFILL_4_OAI22X1_30 INVX1_94/gnd DFFSR_25/S FILL
XOAI22X1_24 INVX1_303/Y OAI22X1_8/B INVX1_304/Y OAI22X1_8/D DFFSR_79/gnd NOR2X1_21/A
+ DFFSR_36/S OAI22X1
XDFFSR_166 INVX1_200/A CLKBUF1_10/Y DFFSR_162/R DFFSR_166/S DFFSR_166/D INVX1_4/gnd
+ DFFSR_51/S DFFSR
XFILL_8_OAI21X1_224 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_2_NAND3X1_51 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_8_DFFSR_25 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_2_INVX1_427 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_3_OAI22X1_33 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_1_NAND3X1_54 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_2_OAI22X1_36 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_25_DFFSR_18 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_14_DFFSR_58 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_4_DFFSR_163 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_1_OAI22X1_39 BUFX2_37/A DFFSR_8/S FILL
XFILL_0_NAND3X1_57 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_0_OAI21X1_103 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_0_OAI22X1_42 INVX1_8/gnd DFFSR_7/S FILL
XFILL_1_INVX1_247 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_49_DFFSR_75 INVX1_4/gnd DFFSR_51/S FILL
XFILL_7_6 BUFX2_35/A DFFSR_14/S FILL
XINVX1_59 DFFSR_52/Q INVX1_94/gnd INVX1_59/Y DFFSR_25/S INVX1
XFILL_0_NAND2X1_217 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_41_5_0 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_33_DFFSR_25 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_5_DFFSR_72 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_22_DFFSR_65 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_48_DFFSR_121 BUFX2_36/A DFFSR_6/S FILL
XINVX1_177 BUFX2_9/Y BUFX2_37/A INVX1_177/Y DFFSR_81/S INVX1
XFILL_4_BUFX2_10 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_38_DFFSR_124 INVX1_89/gnd DFFSR_36/S FILL
XFILL_7_OAI21X1_254 INVX1_23/gnd DFFSR_91/S FILL
XFILL_28_DFFSR_127 BUFX2_43/A DFFSR_97/S FILL
XFILL_1_NAND2X1_151 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_4_INVX1_174 INVX1_94/gnd DFFSR_25/S FILL
XFILL_9_XOR2X1_2 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_4_DFFSR_2 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_18_DFFSR_130 INVX1_4/gnd DFFSR_51/S FILL
XFILL_8_AOI21X1_9 INVX1_94/gnd DFFSR_52/S FILL
XFILL_30_DFFSR_72 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_41_DFFSR_32 INVX1_2/gnd DFFSR_1/S FILL
XFILL_2_INVX1_66 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_3_NAND3X1_12 INVX1_94/gnd DFFSR_52/S FILL
XFILL_8_OAI21X1_188 INVX1_89/gnd DFFSR_2/S FILL
XFILL_2_INVX1_391 BUFX2_17/gnd DFFSR_7/S FILL
XDFFSR_130 NOR2X1_46/A CLKBUF1_13/Y DFFSR_135/R DFFSR_51/S DFFSR_130/D INVX1_4/gnd
+ DFFSR_51/S DFFSR
XFILL_4_DFFSR_127 BUFX2_43/A DFFSR_97/S FILL
XFILL_2_NAND3X1_15 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_14_DFFSR_22 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_46_2 INVX1_2/gnd DFFSR_1/S FILL
XFILL_2_OR2X2_2 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_45_DFFSR_158 BUFX2_43/A DFFSR_23/S FILL
XFILL_11_AOI22X1_5 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_1_NAND3X1_18 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_35_DFFSR_161 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_0_NAND3X1_21 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_28_DFFSR_6 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_25_DFFSR_164 INVX1_89/gnd DFFSR_2/S FILL
XFILL_1_INVX1_211 BUFX2_37/A DFFSR_8/S FILL
XFILL_49_DFFSR_39 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_15_DFFSR_167 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_38_DFFSR_79 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_3_DFFPOSX1_19 BUFX2_16/gnd DFFSR_65/S FILL
XINVX1_23 DFFSR_20/Q INVX1_23/gnd INVX1_23/Y DFFSR_91/S INVX1
XFILL_11_DFFSR_69 BUFX2_43/A DFFSR_23/S FILL
XDFFSR_76 DFFSR_76/Q CLKBUF1_6/Y DFFSR_76/R DFFSR_54/S DFFSR_76/D BUFX2_7/gnd DFFSR_54/S
+ DFFSR
XFILL_0_NAND2X1_181 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_5_DFFSR_36 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_22_DFFSR_29 INVX1_4/gnd DFFSR_4/S FILL
XFILL_0_NOR2X1_46 BUFX2_16/gnd DFFSR_65/S FILL
XINVX1_141 DFFSR_125/Q BUFX2_35/A INVX1_141/Y DFFSR_14/S INVX1
XFILL_8_NAND3X1_134 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_1_DFFSR_164 INVX1_89/gnd DFFSR_2/S FILL
XFILL_47_4_2 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_7_OAI21X1_218 INVX1_23/gnd DFFSR_186/S FILL
XFILL_1_NAND2X1_115 BUFX2_36/A DFFSR_6/S FILL
XFILL_4_INVX1_138 INVX1_94/gnd DFFSR_25/S FILL
XFILL_49_DFFSR_2 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_46_DFFSR_86 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_19_DFFSR_76 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_2_DFFSR_83 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_30_DFFSR_36 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_2_INVX1_30 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_22_DFFPOSX1_27 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_8_OAI21X1_152 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_2_INVX1_355 BUFX2_37/A DFFSR_8/S FILL
XFILL_1_BUFX2_21 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_15_3_0 BUFX2_37/A DFFSR_81/S FILL
XFILL_4_INVX1_4 INVX1_4/gnd DFFSR_4/S FILL
XFILL_45_DFFSR_122 INVX1_94/gnd DFFSR_52/S FILL
XFILL_14_XNOR2X1_4 INVX1_8/gnd DFFSR_7/S FILL
XFILL_35_DFFSR_125 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_13_5_1 BUFX2_36/A DFFSR_8/S FILL
XFILL_27_DFFSR_83 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_25_DFFSR_128 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_1_INVX1_175 INVX1_94/gnd DFFSR_52/S FILL
XFILL_38_DFFSR_43 INVX1_94/gnd DFFSR_25/S FILL
XFILL_15_DFFSR_131 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_0_NAND2X1_145 BUFX2_6/gnd DFFSR_91/S FILL
XDFFSR_40 DFFSR_40/Q DFFSR_28/CLK DFFSR_33/R DFFSR_2/S DFFSR_40/D DFFSR_5/gnd DFFSR_2/S
+ DFFSR
XFILL_6_OAI21X1_248 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_0_XNOR2X1_1 BUFX2_35/A DFFSR_14/S FILL
XFILL_0_NOR2X1_10 BUFX2_36/A DFFSR_6/S FILL
XFILL_11_DFFSR_33 INVX1_94/gnd DFFSR_52/S FILL
XFILL_1_DFFSR_128 BUFX2_19/gnd DFFSR_52/S FILL
XINVX1_105 DFFSR_93/Q INVX1_4/gnd INVX1_105/Y DFFSR_51/S INVX1
XFILL_42_DFFSR_159 BUFX2_36/A DFFSR_6/S FILL
XFILL_7_OAI21X1_182 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_4_INVX1_102 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_46_DFFSR_50 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_32_DFFSR_162 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_35_DFFSR_90 INVX1_2/gnd DFFSR_1/S FILL
XFILL_12_XOR2X1_10 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_22_DFFSR_165 BUFX2_6/gnd DFFSR_14/S FILL
XAOI22X1_3 AND2X2_2/Y AND2X2_7/Y AOI22X1_3/C AOI22X1_3/D BUFX2_7/gnd AOI21X1_4/C DFFSR_54/S
+ AOI22X1
XFILL_12_DFFSR_168 BUFX2_36/A DFFSR_8/S FILL
XFILL_7_NAND3X1_9 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_2_DFFSR_47 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_19_DFFSR_40 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_2_INVX1_319 INVX1_94/gnd DFFSR_25/S FILL
XFILL_8_OAI21X1_116 INVX1_89/gnd DFFSR_2/S FILL
XFILL_23_0_1 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_8_DFFSR_162 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_2_DFFPOSX1_13 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_43_DFFSR_97 BUFX2_35/A DFFSR_97/S FILL
XFILL_4_AND2X2_6 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_1_INVX1_139 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_21_2_2 INVX1_94/gnd DFFSR_25/S FILL
XFILL_27_DFFSR_47 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_7_NAND3X1_128 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_16_DFFSR_87 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_3_1_1 INVX1_23/gnd DFFSR_91/S FILL
XFILL_6_OAI21X1_212 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_0_NAND2X1_109 INVX1_94/gnd DFFSR_25/S FILL
XFILL_1_3_2 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_40_DFFSR_9 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_21_DFFPOSX1_21 BUFX2_5/gnd DFFSR_23/S FILL
XOAI21X1_248 DFFSR_11/S INVX1_410/Y OAI21X1_248/C DFFSR_73/gnd DFFSR_180/D DFFSR_57/S
+ OAI21X1
XFILL_7_OAI21X1_146 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_42_DFFSR_123 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_46_DFFSR_14 BUFX2_35/A DFFSR_14/S FILL
XFILL_35_DFFSR_54 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_24_DFFSR_94 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_32_DFFSR_126 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_22_DFFSR_129 INVX1_2/gnd DFFSR_1/S FILL
XFILL_2_DFFSR_11 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_6_BUFX2_39 BUFX2_43/A DFFSR_97/S FILL
XFILL_11_4 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_48_5_0 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_12_DFFSR_132 INVX1_2/gnd DFFSR_51/S FILL
XFILL_2_INVX1_283 INVX1_4/gnd DFFSR_4/S FILL
XFILL_43_DFFSR_61 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_8_DFFSR_126 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_49_DFFSR_157 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_5_OAI21X1_242 BUFX2_35/A DFFSR_97/S FILL
XFILL_1_INVX1_103 BUFX2_43/A DFFSR_97/S FILL
XFILL_39_DFFSR_160 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_27_DFFSR_11 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_16_DFFSR_51 INVX1_2/gnd DFFSR_51/S FILL
XFILL_29_DFFSR_163 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_6_OAI21X1_176 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_19_DFFSR_166 INVX1_4/gnd DFFSR_51/S FILL
XFILL_14_CLKBUF1_12 BUFX2_43/A DFFSR_23/S FILL
XNOR2X1_48 NOR2X1_48/A NOR2X1_48/B INVX1_89/gnd NOR3X1_2/A DFFSR_36/S NOR2X1
XFILL_1_AOI22X1_1 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_13_CLKBUF1_15 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_4_NOR2X1_45 BUFX2_35/A DFFSR_14/S FILL
XOAI21X1_212 AOI21X1_25/C AOI21X1_22/Y NAND3X1_73/B BUFX2_5/gnd AOI21X1_23/A DFFSR_23/S
+ OAI21X1
XFILL_12_CLKBUF1_18 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_3_INVX1_427 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_7_DFFSR_65 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_7_OAI21X1_110 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_11_CLKBUF1_21 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_13_DFFSR_98 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_35_DFFSR_18 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_24_DFFSR_58 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_5_DFFSR_163 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_10_CLKBUF1_24 INVX1_23/gnd DFFSR_186/S FILL
XFILL_2_INVX1_247 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_27_DFFSR_3 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_10_DFFPOSX1_26 BUFX2_37/A DFFSR_81/S FILL
XFILL_6_NAND3X1_122 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_5_OAI21X1_206 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_4_INVX1_59 INVX1_94/gnd DFFSR_25/S FILL
XFILL_43_DFFSR_25 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_32_DFFSR_65 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_49_DFFSR_121 BUFX2_36/A DFFSR_6/S FILL
XFILL_39_DFFSR_124 INVX1_89/gnd DFFSR_36/S FILL
XFILL_16_DFFSR_15 INVX1_8/gnd DFFSR_7/S FILL
XFILL_29_DFFSR_127 BUFX2_43/A DFFSR_97/S FILL
XXNOR2X1_3 XNOR2X1_3/A XNOR2X1_3/B BUFX2_6/gnd XOR2X1_7/A DFFSR_91/S XNOR2X1
XFILL_20_DFFPOSX1_15 BUFX2_35/A DFFSR_14/S FILL
XFILL_6_OAI21X1_140 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_19_DFFSR_130 INVX1_4/gnd DFFSR_51/S FILL
XFILL_22_3_0 BUFX2_8/gnd DFFSR_25/S FILL
XNOR2X1_12 OAI22X1_6/Y NOR2X1_12/B BUFX2_16/gnd NOR2X1_12/Y DFFSR_65/S NOR2X1
XFILL_40_DFFSR_72 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_51_DFFSR_32 INVX1_2/gnd DFFSR_1/S FILL
XFILL_6_NAND2X1_254 BUFX2_19/gnd DFFSR_52/S FILL
XOAI21X1_176 NOR2X1_4/A NOR2X1_3/A OAI22X1_1/Y BUFX2_8/gnd XOR2X1_2/A DFFSR_25/S OAI21X1
XFILL_33_4 INVX1_8/gnd DFFSR_5/S FILL
XFILL_3_INVX1_391 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_5_DFFSR_127 BUFX2_43/A DFFSR_97/S FILL
XFILL_13_DFFSR_62 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_20_5_1 INVX1_94/gnd DFFSR_52/S FILL
XFILL_24_DFFSR_22 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_7_DFFSR_29 INVX1_4/gnd DFFSR_4/S FILL
XFILL_2_4_0 INVX1_23/gnd DFFSR_186/S FILL
XFILL_46_DFFSR_158 BUFX2_43/A DFFSR_23/S FILL
XFILL_36_DFFSR_161 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_3_INVX1_1 BUFX2_37/A DFFSR_81/S FILL
XFILL_4_OAI21X1_236 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_26_DFFSR_164 INVX1_89/gnd DFFSR_2/S FILL
XFILL_2_INVX1_211 BUFX2_37/A DFFSR_8/S FILL
XFILL_16_DFFSR_167 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_48_DFFSR_79 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_4_INVX1_23 INVX1_23/gnd DFFSR_91/S FILL
XFILL_21_DFFSR_69 BUFX2_43/A DFFSR_23/S FILL
XFILL_4_DFFSR_76 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_32_DFFSR_29 INVX1_4/gnd DFFSR_4/S FILL
XFILL_5_OAI21X1_170 INVX1_94/gnd DFFSR_25/S FILL
XFILL_1_NOR2X1_46 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_0_INVX1_428 DFFSR_71/gnd DFFSR_10/S FILL
XNAND3X1_122 INVX1_331/A INVX1_332/A INVX1_333/Y DFFSR_5/gnd OAI22X1_38/B DFFSR_5/S
+ NAND3X1
XFILL_8_XOR2X1_6 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_3_BUFX2_14 BUFX2_37/A DFFSR_81/S FILL
XFILL_2_DFFSR_164 INVX1_89/gnd DFFSR_2/S FILL
XFILL_5_NAND2X1_284 INVX1_8/gnd DFFSR_5/S FILL
XFILL_6_OAI21X1_104 INVX1_4/gnd DFFSR_51/S FILL
XFILL_2_CLKBUF1_12 BUFX2_43/A DFFSR_23/S FILL
XFILL_29_DFFSR_76 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_1_INVX1_70 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_40_DFFSR_36 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_1_CLKBUF1_15 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_0_CLKBUF1_18 BUFX2_8/gnd DFFSR_25/S FILL
XOAI21X1_140 DFFSR_10/S INVX1_158/Y NAND2X1_140/Y DFFSR_71/gnd DFFSR_140/D DFFSR_45/S
+ OAI21X1
XFILL_30_0_1 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_3_INVX1_355 BUFX2_37/A DFFSR_8/S FILL
XFILL_6_NAND2X1_218 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_28_2_2 INVX1_89/gnd DFFSR_36/S FILL
XFILL_13_DFFSR_26 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_46_DFFSR_122 INVX1_94/gnd DFFSR_52/S FILL
XFILL_5_NAND3X1_116 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_15_XNOR2X1_4 INVX1_8/gnd DFFSR_7/S FILL
XFILL_36_DFFSR_125 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_4_OAI21X1_200 BUFX2_37/A DFFSR_8/S FILL
XNAND2X1_254 NAND2X1_253/Y NAND3X1_130/Y BUFX2_19/gnd NAND2X1_254/Y DFFSR_52/S NAND2X1
XFILL_8_3_2 BUFX2_43/A DFFSR_97/S FILL
XFILL_26_DFFSR_128 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_2_INVX1_175 INVX1_94/gnd DFFSR_52/S FILL
XFILL_48_DFFSR_43 INVX1_94/gnd DFFSR_25/S FILL
XFILL_37_DFFSR_83 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_16_DFFSR_131 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_1_XNOR2X1_1 BUFX2_35/A DFFSR_14/S FILL
XFILL_1_NOR2X1_10 BUFX2_36/A DFFSR_6/S FILL
XFILL_21_DFFSR_33 INVX1_94/gnd DFFSR_52/S FILL
XFILL_5_OAI21X1_134 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_4_DFFSR_40 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_10_DFFSR_73 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_2_DFFSR_128 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_0_INVX1_392 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_39_DFFSR_6 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_43_DFFSR_159 BUFX2_36/A DFFSR_6/S FILL
XFILL_14_XOR2X1_3 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_33_DFFSR_162 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_5_NAND2X1_248 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_45_DFFSR_90 INVX1_2/gnd DFFSR_1/S FILL
XFILL_13_XOR2X1_10 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_23_DFFSR_165 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_25_DFFPOSX1_3 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_13_DFFSR_168 BUFX2_36/A DFFSR_8/S FILL
XFILL_8_NAND3X1_9 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_1_INVX1_34 INVX1_89/gnd DFFSR_36/S FILL
XFILL_29_DFFSR_40 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_1_DFFSR_87 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_24_DFFPOSX1_6 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_18_DFFSR_80 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_3_OAI21X1_230 INVX1_23/gnd DFFSR_186/S FILL
XFILL_23_DFFPOSX1_9 BUFX2_37/A DFFSR_8/S FILL
XFILL_9_DFFPOSX1_20 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_3_INVX1_319 INVX1_94/gnd DFFSR_25/S FILL
XFILL_6_NAND2X1_182 BUFX2_8/gnd DFFSR_25/S FILL
XOAI21X1_104 BUFX2_15/Y INVX1_117/Y NAND2X1_104/Y INVX1_4/gnd DFFSR_104/D DFFSR_51/S
+ OAI21X1
XFILL_0_BUFX2_25 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_9_DFFSR_162 DFFSR_89/gnd DFFSR_92/S FILL
XNAND2X1_218 NAND3X1_85/Y NAND3X1_88/Y DFFSR_73/gnd OAI21X1_229/B DFFSR_57/S NAND2X1
XFILL_4_OAI21X1_164 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_2_INVX1_139 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_37_DFFSR_47 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_26_DFFSR_87 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_9_DFFSR_94 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_4_NAND2X1_278 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_10_DFFSR_37 INVX1_89/gnd DFFSR_2/S FILL
XFILL_0_INVX1_356 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_43_DFFSR_123 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_5_NAND2X1_212 INVX1_23/gnd DFFSR_186/S FILL
XFILL_45_DFFSR_54 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_34_DFFSR_94 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_2_OAI21X1_260 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_33_DFFSR_126 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_4_NAND3X1_110 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_18_DFFSR_44 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_23_DFFSR_129 INVX1_2/gnd DFFSR_1/S FILL
XFILL_1_DFFSR_51 INVX1_2/gnd DFFSR_51/S FILL
XFILL_15_1 BUFX2_37/A DFFSR_8/S FILL
XFILL_3_OAI21X1_194 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_13_DFFSR_132 INVX1_2/gnd DFFSR_51/S FILL
XFILL_6_NAND2X1_146 INVX1_23/gnd DFFSR_91/S FILL
XFILL_3_INVX1_283 INVX1_4/gnd DFFSR_4/S FILL
XFILL_6_DFFSR_9 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_9_DFFSR_126 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_50_DFFSR_157 BUFX2_6/gnd DFFSR_91/S FILL
XNAND2X1_182 NAND3X1_4/Y NAND3X1_5/C BUFX2_8/gnd NAND2X1_182/Y DFFSR_25/S NAND2X1
XFILL_4_OAI21X1_128 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_2_INVX1_103 BUFX2_43/A DFFSR_97/S FILL
XFILL_40_DFFSR_160 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_9_DFFSR_58 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_37_DFFSR_11 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_15_DFFSR_91 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_29_3_0 INVX1_89/gnd DFFSR_2/S FILL
XFILL_26_DFFSR_51 INVX1_2/gnd DFFSR_51/S FILL
XFILL_30_DFFSR_163 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_10_XOR2X1_11 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_20_DFFSR_166 INVX1_4/gnd DFFSR_51/S FILL
XFILL_10_DFFSR_169 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_4_NAND2X1_242 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_27_5_1 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_9_4_0 BUFX2_43/A DFFSR_23/S FILL
XFILL_2_AOI22X1_1 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_0_INVX1_320 INVX1_89/gnd DFFSR_2/S FILL
XFILL_5_NOR2X1_45 BUFX2_35/A DFFSR_14/S FILL
XINVX1_430 DFFSR_142/Q INVX1_89/gnd NOR2X1_48/B DFFSR_36/S INVX1
XFILL_2_OAI21X1_224 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_8_DFFPOSX1_14 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_13_DFFPOSX1_3 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_5_NAND2X1_176 INVX1_94/gnd DFFSR_25/S FILL
XFILL_23_DFFSR_98 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_45_DFFSR_18 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_34_DFFSR_58 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_6_DFFSR_163 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_12_DFFPOSX1_6 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_11_DFFPOSX1_9 BUFX2_37/A DFFSR_8/S FILL
XFILL_5_BUFX2_43 BUFX2_35/A DFFSR_97/S FILL
XFILL_1_DFFSR_15 INVX1_8/gnd DFFSR_7/S FILL
XFILL_3_INVX1_247 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_3_OAI21X1_158 BUFX2_43/A DFFSR_97/S FILL
XFILL_6_NAND2X1_110 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_51_DFFSR_9 DFFSR_9/gnd DFFSR_9/S FILL
XNAND2X1_146 DFFSR_145/Q DFFSR_91/S INVX1_23/gnd OAI21X1_146/C DFFSR_91/S NAND2X1
XFILL_9_AOI21X1_35 INVX1_94/gnd DFFSR_25/S FILL
XFILL_10_CLKBUF1_1 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_3_INVX1_99 INVX1_4/gnd DFFSR_4/S FILL
XFILL_42_DFFSR_65 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_3_NAND2X1_272 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_50_DFFSR_121 BUFX2_36/A DFFSR_6/S FILL
XFILL_8_AOI21X1_38 BUFX2_36/A DFFSR_8/S FILL
XFILL_27_DFFPOSX1_22 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_7_AOI21X1_41 BUFX2_35/A DFFSR_14/S FILL
XFILL_9_DFFSR_22 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_15_DFFSR_55 INVX1_89/gnd DFFSR_36/S FILL
XFILL_40_DFFSR_124 INVX1_89/gnd DFFSR_36/S FILL
XFILL_26_DFFSR_15 INVX1_8/gnd DFFSR_7/S FILL
XFILL_30_DFFSR_127 BUFX2_43/A DFFSR_97/S FILL
XFILL_6_AOI21X1_44 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_37_0_1 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_1_OAI21X1_254 INVX1_23/gnd DFFSR_91/S FILL
XFILL_4_NAND2X1_206 BUFX2_43/A DFFSR_97/S FILL
XFILL_5_AOI21X1_47 BUFX2_43/A DFFSR_23/S FILL
XFILL_20_DFFSR_130 INVX1_4/gnd DFFSR_51/S FILL
XFILL_10_DFFSR_133 BUFX2_37/A DFFSR_81/S FILL
XAOI21X1_44 AND2X2_15/Y AOI21X1_44/B NOR2X1_47/Y BUFX2_17/gnd AND2X2_17/B DFFSR_7/S
+ AOI21X1
XFILL_35_2_2 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_3_NAND3X1_104 INVX1_23/gnd DFFSR_186/S FILL
XFILL_20_6 BUFX2_19/gnd DFFSR_52/S FILL
XINVX1_394 DFFSR_128/Q INVX1_89/gnd INVX1_394/Y DFFSR_2/S INVX1
XFILL_50_DFFSR_72 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_0_INVX1_284 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_6_DFFSR_127 BUFX2_43/A DFFSR_97/S FILL
XFILL_6_DFFSR_69 BUFX2_43/A DFFSR_23/S FILL
XFILL_23_DFFSR_62 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_34_DFFSR_22 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_5_NAND2X1_140 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_2_OAI21X1_188 INVX1_89/gnd DFFSR_2/S FILL
XFILL_47_DFFSR_158 BUFX2_43/A DFFSR_23/S FILL
XFILL_37_DFFSR_161 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_3_OAI21X1_122 INVX1_94/gnd DFFSR_25/S FILL
XFILL_27_DFFSR_164 INVX1_89/gnd DFFSR_2/S FILL
XFILL_3_INVX1_211 BUFX2_37/A DFFSR_8/S FILL
XFILL_9_OAI21X1_83 INVX1_94/gnd DFFSR_52/S FILL
XFILL_17_DFFSR_167 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_17_DFFSR_7 INVX1_8/gnd DFFSR_7/S FILL
XFILL_8_OAI21X1_86 INVX1_4/gnd DFFSR_51/S FILL
XFILL_7_OAI21X1_89 BUFX2_35/A DFFSR_14/S FILL
XFILL_31_DFFSR_69 BUFX2_43/A DFFSR_23/S FILL
XFILL_3_INVX1_63 INVX1_2/gnd DFFSR_51/S FILL
XFILL_42_DFFSR_29 INVX1_4/gnd DFFSR_4/S FILL
XFILL_6_OAI21X1_92 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_3_NAND2X1_236 INVX1_2/gnd DFFSR_1/S FILL
XFILL_2_NOR2X1_46 BUFX2_16/gnd DFFSR_65/S FILL
XNAND2X1_110 BUFX2_17/Y INVX1_376/A DFFSR_73/gnd NAND2X1_110/Y DFFSR_11/S NAND2X1
XFILL_1_BUFX2_8 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_1_INVX1_428 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_5_OAI21X1_95 INVX1_89/gnd DFFSR_36/S FILL
XOAI21X1_92 BUFX2_25/Y INVX1_104/Y NAND2X1_92/Y BUFX2_5/gnd DFFSR_92/D DFFSR_23/S
+ OAI21X1
XFILL_2_NAND3X1_134 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_3_DFFSR_164 INVX1_89/gnd DFFSR_2/S FILL
XFILL_15_DFFSR_19 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_4_OAI21X1_98 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_1_OAI21X1_218 INVX1_23/gnd DFFSR_186/S FILL
XFILL_5_AOI21X1_11 INVX1_8/gnd DFFSR_5/S FILL
XFILL_38_DFFSR_3 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_4_NAND2X1_170 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_0_INVX1_248 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_4_AOI21X1_14 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_39_DFFSR_76 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_50_DFFSR_36 DFFSR_79/gnd DFFSR_36/S FILL
XINVX1_358 INVX1_131/A INVX1_89/gnd INVX1_358/Y DFFSR_36/S INVX1
XFILL_3_AOI21X1_17 INVX1_8/gnd DFFSR_5/S FILL
XFILL_2_OAI21X1_152 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_2_AOI21X1_20 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_1_DFFPOSX1_3 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_16_DFFPOSX1_27 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_1_AOI21X1_23 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_6_DFFSR_33 INVX1_94/gnd DFFSR_52/S FILL
XFILL_23_DFFSR_26 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_12_DFFSR_66 INVX1_2/gnd DFFSR_51/S FILL
XFILL_5_NAND2X1_104 INVX1_4/gnd DFFSR_51/S FILL
XFILL_0_DFFPOSX1_6 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_0_AOI21X1_26 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_47_DFFSR_122 INVX1_94/gnd DFFSR_52/S FILL
XFILL_16_XNOR2X1_4 INVX1_8/gnd DFFSR_7/S FILL
XFILL_37_DFFSR_125 BUFX2_6/gnd DFFSR_91/S FILL
XBUFX2_11 BUFX2_14/A BUFX2_7/gnd BUFX2_11/Y DFFSR_54/S BUFX2
XFILL_26_DFFPOSX1_16 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_27_DFFSR_128 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_3_INVX1_175 INVX1_94/gnd DFFSR_52/S FILL
XFILL_2_NAND2X1_266 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_47_DFFSR_83 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_8_OAI21X1_50 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_17_DFFSR_131 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_6_NAND2X1_71 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_7_OAI21X1_53 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_3_NAND2X1_200 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_2_XNOR2X1_1 BUFX2_35/A DFFSR_14/S FILL
XFILL_2_NOR2X1_10 BUFX2_36/A DFFSR_6/S FILL
XFILL_31_DFFSR_33 INVX1_94/gnd DFFSR_52/S FILL
XFILL_0_OAI21X1_248 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_5_NAND2X1_74 INVX1_2/gnd DFFSR_1/S FILL
XFILL_6_OAI21X1_56 INVX1_2/gnd DFFSR_51/S FILL
XFILL_3_DFFSR_80 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_20_DFFSR_73 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_3_INVX1_27 DFFSR_73/gnd DFFSR_11/S FILL
XNAND2X1_71 BUFX2_23/Y NAND2X1_71/B BUFX2_8/gnd OAI21X1_71/C DFFSR_10/S NAND2X1
XFILL_4_NAND2X1_77 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_5_OAI21X1_59 INVX1_4/gnd DFFSR_51/S FILL
XFILL_4_OAI21X1_62 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_3_DFFSR_128 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_3_NAND2X1_80 BUFX2_17/gnd DFFSR_57/S FILL
XOAI21X1_56 DFFSR_1/S INVX1_63/Y NAND2X1_56/Y INVX1_2/gnd DFFSR_56/D DFFSR_51/S OAI21X1
XFILL_1_INVX1_392 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_44_DFFSR_159 BUFX2_36/A DFFSR_6/S FILL
XFILL_10_AOI22X1_6 BUFX2_37/A DFFSR_81/S FILL
XFILL_2_BUFX2_18 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_34_DFFSR_162 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_2_NAND2X1_83 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_4_NAND2X1_134 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_1_OAI21X1_182 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_3_OAI21X1_65 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_14_XOR2X1_10 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_24_DFFSR_165 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_2_OAI21X1_68 BUFX2_37/A DFFSR_81/S FILL
XFILL_1_NAND2X1_86 INVX1_4/gnd DFFSR_51/S FILL
XFILL_14_DFFSR_168 BUFX2_36/A DFFSR_8/S FILL
XFILL_0_NAND2X1_89 BUFX2_37/A DFFSR_8/S FILL
XFILL_9_NAND3X1_9 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_1_OAI21X1_71 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_0_INVX1_212 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_39_DFFSR_40 DFFSR_5/gnd DFFSR_2/S FILL
XINVX1_322 DFFSR_16/Q BUFX2_17/gnd INVX1_322/Y DFFSR_7/S INVX1
XFILL_0_INVX1_74 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_28_DFFSR_80 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_4_INVX1_319 INVX1_94/gnd DFFSR_25/S FILL
XFILL_0_OAI21X1_74 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_12_DFFSR_30 INVX1_89/gnd DFFSR_36/S FILL
XFILL_2_OAI21X1_116 INVX1_89/gnd DFFSR_2/S FILL
XFILL_36_3_0 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_0_DFFSR_165 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_5_DFFSR_6 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_2_NAND2X1_230 BUFX2_36/A DFFSR_6/S FILL
XFILL_34_5_1 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_3_INVX1_139 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_47_DFFSR_47 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_36_DFFSR_87 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_9_OAI21X1_11 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_8_OAI21X1_14 BUFX2_43/A DFFSR_23/S FILL
XFILL_1_NAND3X1_128 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_0_OAI21X1_212 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_3_DFFSR_44 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_20_DFFSR_37 INVX1_89/gnd DFFSR_2/S FILL
XFILL_7_OAI21X1_17 INVX1_8/gnd DFFSR_5/S FILL
XFILL_6_NAND2X1_35 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_6_OAI21X1_20 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_5_NAND2X1_38 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_3_NAND2X1_164 INVX1_8/gnd DFFSR_5/S FILL
XNAND2X1_35 DFFSR_57/S INVX1_31/A BUFX2_17/gnd OAI21X1_35/C DFFSR_7/S NAND2X1
XFILL_5_OAI21X1_23 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_1_INVX1_356 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_4_NAND2X1_41 DFFSR_5/gnd DFFSR_5/S FILL
XOAI21X1_20 DFFSR_92/S INVX1_23/Y OAI21X1_20/C DFFSR_89/gnd DFFSR_20/D DFFSR_186/S
+ OAI21X1
XFILL_3_NAND2X1_44 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_4_OAI21X1_26 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_1_OAI21X1_146 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_44_DFFSR_123 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_13_XOR2X1_7 INVX1_23/gnd DFFSR_91/S FILL
XFILL_15_DFFPOSX1_21 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_2_NAND2X1_47 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_3_OAI21X1_29 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_44_DFFSR_94 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_1_NAND2X1_50 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_34_DFFSR_126 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_2_OAI21X1_32 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_0_DFFSR_91 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_0_INVX1_176 BUFX2_37/A DFFSR_81/S FILL
XFILL_0_INVX1_38 INVX1_94/gnd DFFSR_52/S FILL
XFILL_28_DFFSR_44 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_0_NAND2X1_53 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_1_OAI21X1_35 INVX1_8/gnd DFFSR_5/S FILL
XFILL_5_AND2X2_3 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_24_DFFSR_129 INVX1_2/gnd DFFSR_1/S FILL
XINVX1_286 INVX1_31/A INVX1_4/gnd INVX1_286/Y DFFSR_51/S INVX1
XFILL_17_DFFSR_84 BUFX2_43/A DFFSR_23/S FILL
XFILL_0_OAI21X1_38 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_14_DFFSR_132 INVX1_2/gnd DFFSR_51/S FILL
XFILL_1_NAND2X1_260 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_25_DFFPOSX1_10 INVX1_8/gnd DFFSR_5/S FILL
XFILL_44_0_1 INVX1_2/gnd DFFSR_51/S FILL
XFILL_7_AOI22X1_10 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_50_DFFSR_6 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_0_DFFSR_129 INVX1_2/gnd DFFSR_1/S FILL
XFILL_6_AOI22X1_13 INVX1_23/gnd DFFSR_186/S FILL
XFILL_3_INVX1_103 BUFX2_43/A DFFSR_97/S FILL
XFILL_2_NAND2X1_194 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_41_DFFSR_160 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_42_2_2 INVX1_4/gnd DFFSR_4/S FILL
XFILL_25_DFFSR_91 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_8_DFFSR_98 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_36_DFFSR_51 INVX1_2/gnd DFFSR_51/S FILL
XFILL_31_DFFSR_163 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_47_DFFSR_11 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_11_XOR2X1_11 DFFSR_73/gnd DFFSR_57/S FILL
XAOI22X1_13 AOI22X1_13/A AOI22X1_13/B AOI22X1_13/C INVX1_255/A INVX1_23/gnd AOI22X1_13/Y
+ DFFSR_186/S AOI22X1
XFILL_21_DFFSR_166 INVX1_4/gnd DFFSR_51/S FILL
XFILL_11_DFFSR_169 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_0_OAI21X1_176 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_3_NAND2X1_128 INVX1_89/gnd DFFSR_2/S FILL
XFILL_3_AOI22X1_1 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_6_NOR2X1_45 BUFX2_35/A DFFSR_14/S FILL
XFILL_11_OAI22X1_46 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_1_INVX1_320 INVX1_89/gnd DFFSR_2/S FILL
XFILL_10_OAI22X1_49 INVX1_94/gnd DFFSR_25/S FILL
XFILL_10_1_0 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_33_DFFSR_98 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_44_DFFSR_58 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_7_DFFSR_163 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_2_NAND2X1_11 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_1_OAI21X1_110 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_8_NAND3X1_70 BUFX2_35/A DFFSR_14/S FILL
XFILL_1_NAND2X1_14 BUFX2_43/A DFFSR_23/S FILL
XAND2X2_7 AND2X2_6/A AND2X2_5/B BUFX2_7/gnd AND2X2_7/Y DFFSR_54/S AND2X2
XFILL_9_OAI22X1_52 INVX1_94/gnd DFFSR_25/S FILL
XFILL_7_NAND3X1_73 BUFX2_43/A DFFSR_23/S FILL
XINVX1_250 INVX1_250/A INVX1_94/gnd INVX1_250/Y DFFSR_25/S INVX1
XFILL_0_INVX1_140 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_0_DFFSR_55 INVX1_89/gnd DFFSR_36/S FILL
XFILL_0_NAND2X1_17 INVX1_8/gnd DFFSR_7/S FILL
XFILL_17_DFFSR_48 INVX1_4/gnd DFFSR_4/S FILL
XFILL_2_2 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_4_INVX1_247 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_1_NAND2X1_224 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_8_OAI22X1_55 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_6_NAND3X1_76 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_7_OAI22X1_58 BUFX2_17/gnd DFFSR_7/S FILL
XNAND3X1_76 NAND3X1_74/Y NAND3X1_75/Y AOI21X1_27/Y BUFX2_5/gnd NAND3X1_76/Y DFFSR_6/S
+ NAND3X1
XFILL_5_NAND3X1_79 BUFX2_36/A DFFSR_6/S FILL
XFILL_6_OAI22X1_61 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_0_NAND3X1_122 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_4_NAND3X1_82 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_5_OAI22X1_64 INVX1_94/gnd DFFSR_25/S FILL
XFILL_11_CLKBUF1_1 BUFX2_8/gnd DFFSR_25/S FILL
XOAI22X1_61 INVX1_381/Y OAI22X1_49/D INVX1_380/Y OAI22X1_52/D DFFSR_79/gnd NOR2X1_40/B
+ DFFSR_45/S OAI22X1
XFILL_16_DFFSR_4 INVX1_4/gnd DFFSR_4/S FILL
XFILL_2_NAND2X1_158 BUFX2_35/A DFFSR_97/S FILL
XFILL_3_NAND3X1_85 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_8_OAI21X1_261 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_4_OAI22X1_67 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_8_DFFSR_62 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_2_NAND3X1_88 INVX1_94/gnd DFFSR_52/S FILL
XFILL_14_DFFSR_95 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_25_DFFSR_55 INVX1_89/gnd DFFSR_36/S FILL
XFILL_41_DFFSR_124 INVX1_89/gnd DFFSR_36/S FILL
XFILL_36_DFFSR_15 INVX1_8/gnd DFFSR_7/S FILL
XFILL_1_NAND3X1_91 BUFX2_43/A DFFSR_97/S FILL
XFILL_31_DFFSR_127 BUFX2_43/A DFFSR_97/S FILL
XFILL_0_BUFX2_5 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_14_DFFPOSX1_15 BUFX2_35/A DFFSR_14/S FILL
XFILL_0_NAND3X1_94 BUFX2_35/A DFFSR_97/S FILL
XFILL_0_OAI21X1_140 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_21_DFFSR_130 INVX1_4/gnd DFFSR_51/S FILL
XFILL_11_DFFSR_133 BUFX2_37/A DFFSR_81/S FILL
XFILL_1_INVX1_284 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_11_OAI22X1_10 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_7_DFFSR_127 BUFX2_43/A DFFSR_97/S FILL
XFILL_0_NAND2X1_254 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_33_DFFSR_62 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_44_DFFSR_22 BUFX2_8/gnd DFFSR_10/S FILL
XINVX1_96 DFFSR_85/Q DFFSR_79/gnd INVX1_96/Y DFFSR_36/S INVX1
XFILL_10_OAI22X1_13 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_48_DFFSR_158 BUFX2_43/A DFFSR_23/S FILL
XFILL_9_NAND3X1_31 INVX1_94/gnd DFFSR_52/S FILL
XFILL_38_DFFSR_161 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_0_INVX1_104 BUFX2_5/gnd DFFSR_23/S FILL
XINVX1_214 AND2X2_11/A BUFX2_5/gnd INVX1_214/Y DFFSR_6/S INVX1
XFILL_0_DFFSR_19 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_8_NAND3X1_34 INVX1_2/gnd DFFSR_1/S FILL
XFILL_9_OAI22X1_16 INVX1_4/gnd DFFSR_4/S FILL
XFILL_17_DFFSR_12 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_7_NAND3X1_37 BUFX2_43/A DFFSR_97/S FILL
XFILL_4_DFFPOSX1_26 BUFX2_37/A DFFSR_81/S FILL
XFILL_16_0_2 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_8_OAI22X1_19 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_28_DFFSR_164 INVX1_89/gnd DFFSR_2/S FILL
XFILL_6_NAND3X1_40 BUFX2_43/A DFFSR_23/S FILL
XFILL_18_DFFSR_167 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_1_NAND2X1_188 INVX1_8/gnd DFFSR_7/S FILL
XFILL_7_OAI22X1_22 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_5_NAND3X1_43 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_6_OAI22X1_25 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_4_NAND3X1_46 BUFX2_35/A DFFSR_97/S FILL
XNAND3X1_40 INVX1_241/A NAND3X1_40/B NAND3X1_40/C BUFX2_43/A NAND3X1_47/B DFFSR_23/S
+ NAND3X1
XFILL_41_DFFSR_69 BUFX2_43/A DFFSR_23/S FILL
XFILL_0_AOI22X1_2 BUFX2_37/A DFFSR_81/S FILL
XFILL_5_OAI22X1_28 INVX1_94/gnd DFFSR_25/S FILL
XFILL_3_NAND3X1_49 BUFX2_37/A DFFSR_8/S FILL
XOAI22X1_25 INVX1_305/Y OAI22X1_6/D INVX1_306/Y OAI22X1_9/B BUFX2_8/gnd NOR2X1_22/B
+ DFFSR_25/S OAI22X1
XFILL_4_OAI22X1_31 DFFSR_71/gnd DFFSR_45/S FILL
XDFFSR_167 INVX1_201/A CLKBUF1_15/Y DFFSR_162/R DFFSR_36/S DFFSR_167/D DFFSR_79/gnd
+ DFFSR_36/S DFFSR
XFILL_3_NOR2X1_46 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_8_OAI21X1_225 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_2_NAND3X1_52 BUFX2_36/A DFFSR_8/S FILL
XFILL_2_NAND2X1_122 INVX1_94/gnd DFFSR_25/S FILL
XFILL_2_INVX1_428 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_3_OAI22X1_34 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_1_NAND3X1_55 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_2_OAI22X1_37 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_4_DFFSR_164 INVX1_89/gnd DFFSR_2/S FILL
XFILL_25_DFFSR_19 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_8_DFFSR_26 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_14_DFFSR_59 INVX1_4/gnd DFFSR_51/S FILL
XFILL_1_OAI22X1_40 BUFX2_37/A DFFSR_8/S FILL
XFILL_0_NAND3X1_58 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_0_OAI21X1_104 INVX1_4/gnd DFFSR_51/S FILL
XFILL_1_INVX1_248 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_49_DFFSR_76 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_0_OAI22X1_43 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_43_3_0 INVX1_4/gnd DFFSR_51/S FILL
XFILL_7_7 BUFX2_35/A DFFSR_14/S FILL
XINVX1_60 DFFSR_53/Q DFFSR_71/gnd INVX1_60/Y DFFSR_45/S INVX1
XFILL_0_NAND2X1_218 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_41_5_1 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_33_DFFSR_26 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_22_DFFSR_66 INVX1_2/gnd DFFSR_51/S FILL
XFILL_5_DFFSR_73 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_48_DFFSR_122 INVX1_94/gnd DFFSR_52/S FILL
XFILL_38_DFFSR_125 BUFX2_6/gnd DFFSR_91/S FILL
XINVX1_178 DFFSR_152/Q BUFX2_5/gnd INVX1_178/Y DFFSR_6/S INVX1
XFILL_1_NAND2X1_152 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_4_BUFX2_11 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_28_DFFSR_128 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_4_INVX1_175 INVX1_94/gnd DFFSR_52/S FILL
XFILL_9_XOR2X1_3 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_7_OAI21X1_255 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_18_DFFSR_131 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_4_DFFSR_3 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_3_XNOR2X1_1 BUFX2_35/A DFFSR_14/S FILL
XFILL_3_NOR2X1_10 BUFX2_36/A DFFSR_6/S FILL
XFILL_4_NAND3X1_10 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_41_DFFSR_33 INVX1_94/gnd DFFSR_52/S FILL
XFILL_2_INVX1_67 INVX1_4/gnd DFFSR_51/S FILL
XFILL_30_DFFSR_73 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_3_NAND3X1_13 INVX1_94/gnd DFFSR_25/S FILL
XFILL_8_OAI21X1_189 DFFSR_73/gnd DFFSR_57/S FILL
XDFFSR_131 XOR2X1_11/A CLKBUF1_13/Y DFFSR_135/R DFFSR_51/S DFFSR_131/D DFFSR_1/gnd
+ DFFSR_1/S DFFSR
XFILL_14_DFFSR_23 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_2_NAND3X1_16 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_4_DFFSR_128 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_46_3 INVX1_2/gnd DFFSR_1/S FILL
XFILL_2_INVX1_392 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_2_OR2X2_3 BUFX2_43/A DFFSR_23/S FILL
XFILL_45_DFFSR_159 BUFX2_36/A DFFSR_6/S FILL
XFILL_1_NAND3X1_19 INVX1_8/gnd DFFSR_5/S FILL
XFILL_35_DFFSR_162 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_0_NAND3X1_22 BUFX2_37/A DFFSR_81/S FILL
XFILL_11_AOI22X1_6 BUFX2_37/A DFFSR_81/S FILL
XFILL_15_XOR2X1_10 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_25_DFFSR_165 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_28_DFFSR_7 INVX1_8/gnd DFFSR_7/S FILL
XFILL_15_DFFSR_168 BUFX2_36/A DFFSR_8/S FILL
XFILL_1_INVX1_212 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_49_DFFSR_40 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_38_DFFSR_80 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_3_DFFPOSX1_20 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_0_NAND2X1_182 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_22_DFFSR_30 INVX1_89/gnd DFFSR_36/S FILL
XFILL_5_DFFSR_37 INVX1_89/gnd DFFSR_2/S FILL
XDFFSR_77 INVX1_87/A CLKBUF1_3/Y DFFSR_76/R DFFSR_2/S DFFSR_77/D INVX1_89/gnd DFFSR_2/S
+ DFFSR
XFILL_11_DFFSR_70 BUFX2_17/gnd DFFSR_57/S FILL
XINVX1_24 INVX1_24/A INVX1_2/gnd INVX1_24/Y DFFSR_51/S INVX1
XFILL_0_NOR2X1_47 BUFX2_17/gnd DFFSR_57/S FILL
XINVX1_142 INVX1_378/A BUFX2_17/gnd INVX1_142/Y DFFSR_7/S INVX1
XFILL_1_DFFSR_165 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_4_INVX1_139 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_7_OAI21X1_219 BUFX2_35/A DFFSR_97/S FILL
XFILL_1_NAND2X1_116 INVX1_89/gnd DFFSR_36/S FILL
XFILL_46_DFFSR_87 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_49_DFFSR_3 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_2_DFFSR_84 BUFX2_43/A DFFSR_23/S FILL
XFILL_30_DFFSR_37 INVX1_89/gnd DFFSR_2/S FILL
XFILL_2_INVX1_31 INVX1_2/gnd DFFSR_1/S FILL
XFILL_17_1_0 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_19_DFFSR_77 INVX1_89/gnd DFFSR_2/S FILL
XFILL_22_DFFPOSX1_28 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_8_OAI21X1_153 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_2_INVX1_356 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_15_3_1 BUFX2_37/A DFFSR_81/S FILL
XFILL_1_BUFX2_22 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_4_INVX1_5 INVX1_4/gnd DFFSR_51/S FILL
XFILL_45_DFFSR_123 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_13_5_2 BUFX2_36/A DFFSR_8/S FILL
XFILL_11_NOR3X1_1 INVX1_94/gnd DFFSR_52/S FILL
XFILL_35_DFFSR_126 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_1_INVX1_176 BUFX2_37/A DFFSR_81/S FILL
XFILL_25_DFFSR_129 INVX1_2/gnd DFFSR_1/S FILL
XFILL_27_DFFSR_84 BUFX2_43/A DFFSR_23/S FILL
XFILL_38_DFFSR_44 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_15_DFFSR_132 INVX1_2/gnd DFFSR_51/S FILL
XFILL_0_NAND2X1_146 INVX1_23/gnd DFFSR_91/S FILL
XFILL_6_OAI21X1_249 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_0_NOR2X1_11 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_0_XNOR2X1_2 BUFX2_36/A DFFSR_8/S FILL
XDFFSR_41 INVX1_47/A DFFSR_2/CLK DFFSR_46/R DFFSR_57/S DFFSR_41/D BUFX2_17/gnd DFFSR_57/S
+ DFFSR
XFILL_11_DFFSR_34 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_1_DFFSR_129 INVX1_2/gnd DFFSR_1/S FILL
XINVX1_106 DFFSR_94/Q BUFX2_16/gnd INVX1_106/Y DFFSR_11/S INVX1
XFILL_4_INVX1_103 BUFX2_43/A DFFSR_97/S FILL
XFILL_7_OAI21X1_183 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_42_DFFSR_160 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_15_DFFSR_1 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_35_DFFSR_91 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_46_DFFSR_51 INVX1_2/gnd DFFSR_51/S FILL
XFILL_32_DFFSR_163 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_12_XOR2X1_11 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_22_DFFSR_166 INVX1_4/gnd DFFSR_51/S FILL
XAOI22X1_4 NAND3X1_9/Y AOI22X1_4/B AOI22X1_4/C AOI22X1_4/D INVX1_94/gnd NOR3X1_1/B
+ DFFSR_25/S AOI22X1
XFILL_19_DFFSR_41 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_2_DFFSR_48 INVX1_4/gnd DFFSR_4/S FILL
XFILL_8_OAI21X1_117 BUFX2_35/A DFFSR_97/S FILL
XFILL_12_DFFSR_169 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_4_AOI22X1_1 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_2_INVX1_320 INVX1_89/gnd DFFSR_2/S FILL
XFILL_23_0_2 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_2_DFFPOSX1_14 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_43_DFFSR_98 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_8_DFFSR_163 DFFSR_3/gnd DFFSR_65/S FILL
XAND2X2_10 BUFX2_11/Y AND2X2_10/B BUFX2_5/gnd AND2X2_10/Y DFFSR_23/S AND2X2
XFILL_4_AND2X2_7 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_1_INVX1_140 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_27_DFFSR_48 INVX1_4/gnd DFFSR_4/S FILL
XFILL_16_DFFSR_88 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_3_1_2 INVX1_23/gnd DFFSR_91/S FILL
XFILL_7_NAND3X1_129 BUFX2_35/A DFFSR_14/S FILL
XFILL_6_OAI21X1_213 BUFX2_36/A DFFSR_6/S FILL
XFILL_0_NAND2X1_110 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_12_CLKBUF1_1 BUFX2_8/gnd DFFSR_25/S FILL
XOAI21X1_249 DFFSR_186/S INVX1_411/Y OAI21X1_249/C DFFSR_89/gnd DFFSR_181/D DFFSR_186/S
+ OAI21X1
XFILL_7_OAI21X1_147 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_24_DFFSR_95 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_35_DFFSR_55 INVX1_89/gnd DFFSR_36/S FILL
XFILL_42_DFFSR_124 INVX1_89/gnd DFFSR_36/S FILL
XFILL_46_DFFSR_15 INVX1_8/gnd DFFSR_7/S FILL
XFILL_21_DFFPOSX1_22 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_32_DFFSR_127 BUFX2_43/A DFFSR_97/S FILL
XFILL_2_DFFSR_12 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_22_DFFSR_130 INVX1_4/gnd DFFSR_51/S FILL
XFILL_6_BUFX2_40 BUFX2_35/A DFFSR_14/S FILL
XFILL_11_5 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_12_DFFSR_133 BUFX2_37/A DFFSR_81/S FILL
XFILL_48_5_1 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_2_INVX1_284 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_8_DFFSR_127 BUFX2_43/A DFFSR_97/S FILL
XFILL_43_DFFSR_62 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_5_OAI21X1_243 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_49_DFFSR_158 BUFX2_43/A DFFSR_23/S FILL
XFILL_39_DFFSR_161 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_1_INVX1_104 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_27_DFFSR_12 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_16_DFFSR_52 INVX1_94/gnd DFFSR_52/S FILL
XFILL_29_DFFSR_164 INVX1_89/gnd DFFSR_2/S FILL
XFILL_19_DFFSR_167 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_15_CLKBUF1_10 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_6_OAI21X1_177 DFFSR_71/gnd DFFSR_10/S FILL
XNOR2X1_49 DFFSR_134/Q DFFSR_142/Q INVX1_89/gnd NOR3X1_2/B DFFSR_36/S NOR2X1
XFILL_1_AOI22X1_2 BUFX2_37/A DFFSR_81/S FILL
XFILL_14_CLKBUF1_13 INVX1_4/gnd DFFSR_51/S FILL
XOAI21X1_213 INVX1_238/A AOI21X1_23/Y NAND3X1_52/B BUFX2_36/A NAND3X1_72/C DFFSR_6/S
+ OAI21X1
XFILL_13_CLKBUF1_16 BUFX2_36/A DFFSR_6/S FILL
XFILL_4_NOR2X1_46 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_3_INVX1_428 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_7_OAI21X1_111 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_12_CLKBUF1_19 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_13_DFFSR_99 BUFX2_35/A DFFSR_97/S FILL
XFILL_11_CLKBUF1_22 INVX1_94/gnd DFFSR_25/S FILL
XFILL_5_DFFSR_164 INVX1_89/gnd DFFSR_2/S FILL
XFILL_35_DFFSR_19 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_7_DFFSR_66 INVX1_2/gnd DFFSR_51/S FILL
XFILL_24_DFFSR_59 INVX1_4/gnd DFFSR_51/S FILL
XFILL_10_CLKBUF1_25 INVX1_23/gnd DFFSR_186/S FILL
XFILL_2_INVX1_248 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_27_DFFSR_4 INVX1_4/gnd DFFSR_4/S FILL
XFILL_10_DFFPOSX1_27 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_6_NAND3X1_123 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_5_OAI21X1_207 BUFX2_37/A DFFSR_8/S FILL
XFILL_4_INVX1_60 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_43_DFFSR_26 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_32_DFFSR_66 INVX1_2/gnd DFFSR_51/S FILL
XFILL_49_DFFSR_122 INVX1_94/gnd DFFSR_52/S FILL
XFILL_39_DFFSR_125 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_16_DFFSR_16 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_29_DFFSR_128 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_24_1_0 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_20_DFFPOSX1_16 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_6_OAI21X1_141 INVX1_94/gnd DFFSR_52/S FILL
XXNOR2X1_4 XNOR2X1_4/A XOR2X1_13/Y INVX1_8/gnd XNOR2X1_4/Y DFFSR_7/S XNOR2X1
XFILL_19_DFFSR_131 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_22_3_1 BUFX2_8/gnd DFFSR_25/S FILL
XNOR2X1_13 NOR2X1_13/A OAI22X1_7/Y BUFX2_17/gnd NOR2X1_13/Y DFFSR_57/S NOR2X1
XFILL_4_XNOR2X1_1 BUFX2_35/A DFFSR_14/S FILL
XFILL_4_NOR2X1_10 BUFX2_36/A DFFSR_6/S FILL
XFILL_51_DFFSR_33 INVX1_94/gnd DFFSR_52/S FILL
XFILL_40_DFFSR_73 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_4_2_0 BUFX2_6/gnd DFFSR_91/S FILL
XOAI21X1_177 NAND3X1_2/A XOR2X1_2/A NAND3X1_2/Y DFFSR_71/gnd DFFPOSX1_3/D DFFSR_10/S
+ OAI21X1
XFILL_33_5 INVX1_8/gnd DFFSR_5/S FILL
XFILL_24_DFFSR_23 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_5_DFFSR_128 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_20_5_2 INVX1_94/gnd DFFSR_52/S FILL
XFILL_13_DFFSR_63 INVX1_94/gnd DFFSR_52/S FILL
XFILL_7_DFFSR_30 INVX1_89/gnd DFFSR_36/S FILL
XFILL_6_NAND2X1_255 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_3_INVX1_392 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_2_4_1 INVX1_23/gnd DFFSR_186/S FILL
XFILL_46_DFFSR_159 BUFX2_36/A DFFSR_6/S FILL
XFILL_36_DFFSR_162 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_26_DFFSR_165 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_4_OAI21X1_237 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_3_INVX1_2 INVX1_2/gnd DFFSR_51/S FILL
XFILL_2_INVX1_212 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_48_DFFSR_80 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_16_DFFSR_168 BUFX2_36/A DFFSR_8/S FILL
XFILL_32_DFFSR_30 INVX1_89/gnd DFFSR_36/S FILL
XFILL_4_DFFSR_77 INVX1_89/gnd DFFSR_2/S FILL
XFILL_21_DFFSR_70 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_4_INVX1_24 INVX1_2/gnd DFFSR_51/S FILL
XFILL_5_OAI21X1_171 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_1_NOR2X1_47 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_0_INVX1_429 INVX1_89/gnd DFFSR_2/S FILL
XNAND3X1_123 INVX1_397/A INVX1_331/A INVX1_332/Y DFFSR_5/gnd OAI22X1_39/B DFFSR_2/S
+ NAND3X1
XFILL_2_DFFSR_165 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_3_BUFX2_15 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_8_XOR2X1_7 INVX1_23/gnd DFFSR_91/S FILL
XFILL_5_NAND2X1_285 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_3_CLKBUF1_10 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_6_OAI21X1_105 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_2_CLKBUF1_13 INVX1_4/gnd DFFSR_51/S FILL
XFILL_1_CLKBUF1_16 BUFX2_36/A DFFSR_6/S FILL
XFILL_1_INVX1_71 INVX1_94/gnd DFFSR_25/S FILL
XFILL_40_DFFSR_37 INVX1_89/gnd DFFSR_2/S FILL
XOAI21X1_141 DFFSR_25/S INVX1_159/Y OAI21X1_141/C INVX1_94/gnd DFFSR_141/D DFFSR_52/S
+ OAI21X1
XFILL_29_DFFSR_77 INVX1_89/gnd DFFSR_2/S FILL
XFILL_30_0_2 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_0_CLKBUF1_19 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_3_INVX1_356 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_6_NAND2X1_219 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_13_DFFSR_27 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_46_DFFSR_123 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_5_NAND3X1_117 INVX1_94/gnd DFFSR_25/S FILL
XFILL_4_OAI21X1_201 BUFX2_35/A DFFSR_97/S FILL
XFILL_36_DFFSR_126 BUFX2_17/gnd DFFSR_57/S FILL
XNAND2X1_255 din[0] DFFSR_4/S DFFSR_3/gnd OAI21X1_244/C DFFSR_4/S NAND2X1
XFILL_2_INVX1_176 BUFX2_37/A DFFSR_81/S FILL
XFILL_26_DFFSR_129 INVX1_2/gnd DFFSR_1/S FILL
XFILL_37_DFFSR_84 BUFX2_43/A DFFSR_23/S FILL
XFILL_48_DFFSR_44 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_16_DFFSR_132 INVX1_2/gnd DFFSR_51/S FILL
XFILL_1_NOR2X1_11 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_5_OAI21X1_135 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_1_XNOR2X1_2 BUFX2_36/A DFFSR_8/S FILL
XFILL_19_DFFPOSX1_10 INVX1_8/gnd DFFSR_5/S FILL
XFILL_4_DFFSR_41 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_21_DFFSR_34 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_10_DFFSR_74 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_0_INVX1_393 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_14_XOR2X1_4 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_39_DFFSR_7 INVX1_8/gnd DFFSR_7/S FILL
XFILL_43_DFFSR_160 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_2_DFFSR_129 INVX1_2/gnd DFFSR_1/S FILL
XFILL_45_DFFSR_91 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_26_DFFPOSX1_1 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_5_NAND2X1_249 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_33_DFFSR_163 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_13_XOR2X1_11 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_25_DFFPOSX1_4 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_23_DFFSR_166 INVX1_4/gnd DFFSR_51/S FILL
XFILL_1_INVX1_35 BUFX2_35/A DFFSR_97/S FILL
XFILL_18_DFFSR_81 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_24_DFFPOSX1_7 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_29_DFFSR_41 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_1_DFFSR_88 DFFSR_3/gnd DFFSR_4/S FILL
XOAI21X1_105 BUFX2_21/Y INVX1_119/Y OAI21X1_105/C BUFX2_6/gnd DFFSR_105/D DFFSR_14/S
+ OAI21X1
XFILL_9_DFFPOSX1_21 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_13_DFFSR_169 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_3_OAI21X1_231 BUFX2_36/A DFFSR_6/S FILL
XFILL_5_AOI22X1_1 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_3_INVX1_320 INVX1_89/gnd DFFSR_2/S FILL
XFILL_6_NAND2X1_183 INVX1_8/gnd DFFSR_7/S FILL
XFILL_0_BUFX2_26 DFFSR_9/gnd DFFSR_9/S FILL
XNAND2X1_219 NAND3X1_77/Y NAND3X1_81/Y BUFX2_19/gnd INVX1_251/A DFFSR_54/S NAND2X1
XFILL_9_DFFSR_163 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_4_OAI21X1_165 BUFX2_35/A DFFSR_97/S FILL
XFILL_2_INVX1_140 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_9_DFFSR_95 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_37_DFFSR_48 INVX1_4/gnd DFFSR_4/S FILL
XFILL_26_DFFSR_88 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_4_NAND2X1_279 INVX1_89/gnd DFFSR_2/S FILL
XFILL_10_DFFSR_38 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_0_INVX1_357 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_13_CLKBUF1_1 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_5_NAND2X1_213 BUFX2_35/A DFFSR_97/S FILL
XFILL_34_DFFSR_95 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_2_OAI21X1_261 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_45_DFFSR_55 INVX1_89/gnd DFFSR_36/S FILL
XFILL_43_DFFSR_124 INVX1_89/gnd DFFSR_36/S FILL
XFILL_33_DFFSR_127 BUFX2_43/A DFFSR_97/S FILL
XFILL_1_DFFSR_52 INVX1_94/gnd DFFSR_52/S FILL
XFILL_4_NAND3X1_111 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_23_DFFSR_130 INVX1_4/gnd DFFSR_51/S FILL
XFILL_15_2 BUFX2_37/A DFFSR_8/S FILL
XFILL_13_DFFSR_133 BUFX2_37/A DFFSR_81/S FILL
XFILL_18_DFFSR_45 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_6_NAND2X1_147 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_3_OAI21X1_195 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_3_INVX1_284 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_9_DFFSR_127 BUFX2_43/A DFFSR_97/S FILL
XFILL_31_1_0 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_26_DFFSR_1 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_50_DFFSR_158 BUFX2_43/A DFFSR_23/S FILL
XNAND2X1_183 INVX1_223/A AOI21X1_1/A INVX1_8/gnd NAND2X1_183/Y DFFSR_7/S NAND2X1
XFILL_4_OAI21X1_129 INVX1_4/gnd DFFSR_4/S FILL
XFILL_40_DFFSR_161 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_2_INVX1_104 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_15_DFFSR_92 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_37_DFFSR_12 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_26_DFFSR_52 INVX1_94/gnd DFFSR_52/S FILL
XFILL_30_DFFSR_164 INVX1_89/gnd DFFSR_2/S FILL
XFILL_29_3_1 INVX1_89/gnd DFFSR_2/S FILL
XFILL_10_XOR2X1_12 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_9_DFFSR_59 INVX1_4/gnd DFFSR_51/S FILL
XFILL_27_5_2 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_20_DFFSR_167 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_4_NAND2X1_243 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_9_4_1 BUFX2_43/A DFFSR_23/S FILL
XFILL_2_AOI22X1_2 BUFX2_37/A DFFSR_81/S FILL
XFILL_10_DFFSR_170 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_14_DFFPOSX1_1 BUFX2_6/gnd DFFSR_14/S FILL
XINVX1_431 AND2X2_16/B INVX1_89/gnd INVX1_431/Y DFFSR_36/S INVX1
XFILL_0_INVX1_321 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_5_NOR2X1_46 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_2_OAI21X1_225 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_8_DFFPOSX1_15 BUFX2_35/A DFFSR_14/S FILL
XFILL_4_INVX1_428 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_13_DFFPOSX1_4 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_23_DFFSR_99 BUFX2_35/A DFFSR_97/S FILL
XFILL_5_NAND2X1_177 INVX1_89/gnd DFFSR_36/S FILL
XFILL_6_DFFSR_164 INVX1_89/gnd DFFSR_2/S FILL
XFILL_45_DFFSR_19 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_34_DFFSR_59 INVX1_4/gnd DFFSR_51/S FILL
XFILL_12_DFFPOSX1_7 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_1_DFFSR_16 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_3_OAI21X1_159 BUFX2_43/A DFFSR_97/S FILL
XFILL_3_INVX1_248 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_6_NAND2X1_111 DFFSR_5/gnd DFFSR_5/S FILL
XNAND2X1_147 DFFSR_146/Q DFFSR_92/S DFFSR_89/gnd NAND2X1_147/Y DFFSR_92/S NAND2X1
XFILL_42_DFFSR_66 INVX1_2/gnd DFFSR_51/S FILL
XFILL_27_DFFPOSX1_23 INVX1_23/gnd DFFSR_91/S FILL
XFILL_8_AOI21X1_39 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_50_DFFSR_122 INVX1_94/gnd DFFSR_52/S FILL
XFILL_10_CLKBUF1_2 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_3_NAND2X1_273 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_7_AOI21X1_42 INVX1_23/gnd DFFSR_91/S FILL
XFILL_40_DFFSR_125 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_9_DFFSR_23 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_26_DFFSR_16 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_15_DFFSR_56 INVX1_2/gnd DFFSR_51/S FILL
XFILL_30_DFFSR_128 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_6_AOI21X1_45 INVX1_89/gnd DFFSR_36/S FILL
XFILL_37_0_2 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_4_NAND2X1_207 BUFX2_43/A DFFSR_97/S FILL
XFILL_5_AOI21X1_48 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_20_DFFSR_131 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_1_OAI21X1_255 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_10_DFFSR_134 DFFSR_79/gnd DFFSR_45/S FILL
XAOI21X1_45 XOR2X1_15/B INVX1_431/Y NOR3X1_2/A INVX1_89/gnd INVX1_436/A DFFSR_36/S
+ AOI21X1
XFILL_3_NAND3X1_105 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_5_XNOR2X1_1 BUFX2_35/A DFFSR_14/S FILL
XFILL_5_NOR2X1_10 BUFX2_36/A DFFSR_6/S FILL
XINVX1_395 INVX1_81/A DFFSR_5/gnd INVX1_395/Y DFFSR_5/S INVX1
XFILL_0_INVX1_285 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_50_DFFSR_73 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_20_7 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_34_DFFSR_23 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_23_DFFSR_63 INVX1_94/gnd DFFSR_52/S FILL
XFILL_5_NAND2X1_141 INVX1_94/gnd DFFSR_25/S FILL
XFILL_6_DFFSR_70 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_2_OAI21X1_189 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_4_INVX1_392 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_47_DFFSR_159 BUFX2_36/A DFFSR_6/S FILL
XFILL_6_DFFSR_128 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_37_DFFSR_162 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_27_DFFSR_165 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_3_OAI21X1_123 INVX1_23/gnd DFFSR_91/S FILL
XFILL_9_OAI21X1_84 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_3_INVX1_212 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_17_DFFSR_168 BUFX2_36/A DFFSR_8/S FILL
XFILL_17_DFFSR_8 BUFX2_36/A DFFSR_8/S FILL
XFILL_8_OAI21X1_87 INVX1_4/gnd DFFSR_4/S FILL
XFILL_3_INVX1_64 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_42_DFFSR_30 INVX1_89/gnd DFFSR_36/S FILL
XFILL_31_DFFSR_70 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_7_OAI21X1_90 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_3_NAND2X1_237 BUFX2_8/gnd DFFSR_10/S FILL
XNAND2X1_111 BUFX2_22/Y INVX1_116/A DFFSR_5/gnd NAND2X1_111/Y DFFSR_5/S NAND2X1
XFILL_2_NOR2X1_47 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_6_OAI21X1_93 INVX1_4/gnd DFFSR_51/S FILL
XFILL_1_BUFX2_9 BUFX2_37/A DFFSR_8/S FILL
XFILL_1_INVX1_429 INVX1_89/gnd DFFSR_2/S FILL
XFILL_5_OAI21X1_96 INVX1_4/gnd DFFSR_51/S FILL
XFILL_15_DFFSR_20 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_3_DFFSR_165 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_4_OAI21X1_99 BUFX2_43/A DFFSR_97/S FILL
XOAI21X1_93 BUFX2_15/Y INVX1_105/Y NAND2X1_93/Y INVX1_4/gnd DFFSR_93/D DFFSR_51/S
+ OAI21X1
XFILL_1_OAI21X1_219 BUFX2_35/A DFFSR_97/S FILL
XFILL_4_NAND2X1_171 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_6_NOR3X1_1 INVX1_94/gnd DFFSR_52/S FILL
XFILL_5_AOI21X1_12 INVX1_8/gnd DFFSR_7/S FILL
XFILL_4_AOI21X1_15 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_38_DFFSR_4 INVX1_4/gnd DFFSR_4/S FILL
XFILL_2_DFFPOSX1_1 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_0_INVX1_249 BUFX2_35/A DFFSR_14/S FILL
XFILL_3_AOI21X1_18 BUFX2_8/gnd DFFSR_10/S FILL
XINVX1_359 INVX1_122/A DFFSR_79/gnd INVX1_359/Y DFFSR_36/S INVX1
XFILL_50_DFFSR_37 INVX1_89/gnd DFFSR_2/S FILL
XFILL_39_DFFSR_77 INVX1_89/gnd DFFSR_2/S FILL
XFILL_2_AOI21X1_21 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_2_OAI21X1_153 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_4_INVX1_356 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_1_DFFPOSX1_4 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_16_DFFPOSX1_28 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_5_NAND2X1_105 BUFX2_35/A DFFSR_14/S FILL
XFILL_1_AOI21X1_24 BUFX2_43/A DFFSR_97/S FILL
XFILL_0_DFFPOSX1_7 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_23_DFFSR_27 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_6_DFFSR_34 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_12_DFFSR_67 INVX1_2/gnd DFFSR_51/S FILL
XFILL_47_DFFSR_123 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_0_AOI21X1_27 BUFX2_5/gnd DFFSR_6/S FILL
XBUFX2_12 BUFX2_14/A BUFX2_37/A BUFX2_12/Y DFFSR_81/S BUFX2
XFILL_37_DFFSR_126 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_26_DFFPOSX1_17 BUFX2_37/A DFFSR_8/S FILL
XFILL_27_DFFSR_129 INVX1_2/gnd DFFSR_1/S FILL
XFILL_2_NAND2X1_267 INVX1_4/gnd DFFSR_4/S FILL
XFILL_47_DFFSR_84 BUFX2_43/A DFFSR_23/S FILL
XFILL_3_INVX1_176 BUFX2_37/A DFFSR_81/S FILL
XFILL_17_DFFSR_132 INVX1_2/gnd DFFSR_51/S FILL
XFILL_8_OAI21X1_51 INVX1_2/gnd DFFSR_51/S FILL
XFILL_7_OAI21X1_54 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_6_NAND2X1_72 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_0_OAI21X1_249 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_2_NOR2X1_11 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_2_XNOR2X1_2 BUFX2_36/A DFFSR_8/S FILL
XFILL_3_DFFSR_81 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_3_INVX1_28 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_31_DFFSR_34 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_20_DFFSR_74 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_5_NAND2X1_75 INVX1_4/gnd DFFSR_4/S FILL
XFILL_3_NAND2X1_201 BUFX2_35/A DFFSR_14/S FILL
XNAND2X1_72 BUFX2_17/Y NAND2X1_72/B DFFSR_5/gnd OAI21X1_72/C DFFSR_2/S NAND2X1
XFILL_6_OAI21X1_57 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_5_OAI21X1_60 BUFX2_37/A DFFSR_81/S FILL
XFILL_1_INVX1_393 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_4_NAND2X1_78 DFFSR_73/gnd DFFSR_11/S FILL
XOAI21X1_57 DFFSR_11/S INVX1_65/Y NAND2X1_57/Y DFFSR_73/gnd DFFSR_57/D DFFSR_11/S
+ OAI21X1
XFILL_2_BUFX2_19 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_4_OAI21X1_63 INVX1_94/gnd DFFSR_25/S FILL
XFILL_3_NAND2X1_81 INVX1_94/gnd DFFSR_25/S FILL
XFILL_44_DFFSR_160 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_3_DFFSR_129 INVX1_2/gnd DFFSR_1/S FILL
XFILL_10_AOI22X1_7 BUFX2_43/A DFFSR_23/S FILL
XFILL_4_NAND2X1_135 BUFX2_36/A DFFSR_6/S FILL
XFILL_2_NAND2X1_84 BUFX2_36/A DFFSR_6/S FILL
XFILL_1_OAI21X1_183 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_3_OAI21X1_66 INVX1_4/gnd DFFSR_51/S FILL
XFILL_34_DFFSR_163 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_14_XOR2X1_11 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_2_OAI21X1_69 BUFX2_37/A DFFSR_8/S FILL
XFILL_1_NAND2X1_87 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_0_INVX1_213 BUFX2_36/A DFFSR_8/S FILL
XFILL_28_DFFSR_81 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_1_OAI21X1_72 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_39_DFFSR_41 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_0_NAND2X1_90 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_0_INVX1_75 INVX1_4/gnd DFFSR_51/S FILL
XFILL_24_DFFSR_166 INVX1_4/gnd DFFSR_51/S FILL
XINVX1_323 DFFSR_56/Q BUFX2_16/gnd INVX1_323/Y DFFSR_65/S INVX1
XFILL_14_DFFSR_169 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_6_AOI22X1_1 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_0_OAI21X1_75 INVX1_4/gnd DFFSR_4/S FILL
XFILL_38_1_0 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_12_DFFSR_31 BUFX2_35/A DFFSR_97/S FILL
XFILL_2_OAI21X1_117 BUFX2_35/A DFFSR_97/S FILL
XFILL_4_INVX1_320 INVX1_89/gnd DFFSR_2/S FILL
XFILL_36_3_1 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_2_NAND2X1_231 BUFX2_37/A DFFSR_81/S FILL
XFILL_5_DFFSR_7 INVX1_8/gnd DFFSR_7/S FILL
XFILL_34_5_2 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_0_DFFSR_166 INVX1_4/gnd DFFSR_51/S FILL
XFILL_9_OAI21X1_12 BUFX2_35/A DFFSR_14/S FILL
XFILL_3_INVX1_140 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_47_DFFSR_48 INVX1_4/gnd DFFSR_4/S FILL
XFILL_36_DFFSR_88 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_1_NAND3X1_129 BUFX2_35/A DFFSR_14/S FILL
XFILL_8_OAI21X1_15 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_6_NAND2X1_36 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_3_DFFSR_45 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_7_OAI21X1_18 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_0_OAI21X1_213 BUFX2_36/A DFFSR_6/S FILL
XFILL_3_NAND2X1_165 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_5_NAND2X1_39 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_20_DFFSR_38 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_6_OAI21X1_21 INVX1_2/gnd DFFSR_51/S FILL
XFILL_1_INVX1_357 BUFX2_19/gnd DFFSR_52/S FILL
XNAND2X1_36 DFFSR_45/S INVX1_32/A DFFSR_71/gnd NAND2X1_36/Y DFFSR_45/S NAND2X1
XFILL_4_NAND2X1_42 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_5_OAI21X1_24 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_14_CLKBUF1_1 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_3_NAND2X1_45 INVX1_89/gnd DFFSR_36/S FILL
XFILL_4_OAI21X1_27 DFFSR_1/gnd DFFSR_1/S FILL
XOAI21X1_21 DFFSR_51/S INVX1_24/Y NAND2X1_21/Y INVX1_2/gnd DFFSR_21/D DFFSR_51/S OAI21X1
XFILL_1_OAI21X1_147 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_13_XOR2X1_8 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_44_DFFSR_95 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_3_OAI21X1_30 INVX1_89/gnd DFFSR_36/S FILL
XFILL_44_DFFSR_124 INVX1_89/gnd DFFSR_36/S FILL
XFILL_15_DFFPOSX1_22 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_2_NAND2X1_48 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_34_DFFSR_127 BUFX2_43/A DFFSR_97/S FILL
XFILL_2_OAI21X1_33 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_1_NAND2X1_51 INVX1_2/gnd DFFSR_51/S FILL
XFILL_0_NAND2X1_54 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_5_AND2X2_4 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_1_OAI21X1_36 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_24_DFFSR_130 INVX1_4/gnd DFFSR_51/S FILL
XFILL_0_DFFSR_92 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_14_DFFSR_133 BUFX2_37/A DFFSR_81/S FILL
XFILL_0_INVX1_177 BUFX2_37/A DFFSR_81/S FILL
XFILL_0_OAI21X1_39 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_17_DFFSR_85 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_28_DFFSR_45 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_0_INVX1_39 DFFSR_1/gnd DFFSR_1/S FILL
XINVX1_287 INVX1_67/A INVX1_4/gnd INVX1_287/Y DFFSR_51/S INVX1
XFILL_1_NAND2X1_261 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_4_INVX1_284 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_25_DFFPOSX1_11 INVX1_4/gnd DFFSR_4/S FILL
XFILL_44_0_2 INVX1_2/gnd DFFSR_51/S FILL
XFILL_7_AOI22X1_11 INVX1_23/gnd DFFSR_91/S FILL
XFILL_50_DFFSR_7 INVX1_8/gnd DFFSR_7/S FILL
XFILL_41_DFFSR_161 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_2_NAND2X1_195 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_6_AOI22X1_14 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_0_DFFSR_130 INVX1_4/gnd DFFSR_51/S FILL
XFILL_25_DFFSR_92 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_47_DFFSR_12 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_8_DFFSR_99 BUFX2_35/A DFFSR_97/S FILL
XFILL_3_INVX1_104 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_36_DFFSR_52 INVX1_94/gnd DFFSR_52/S FILL
XFILL_31_DFFSR_164 INVX1_89/gnd DFFSR_2/S FILL
XFILL_11_XOR2X1_12 BUFX2_17/gnd DFFSR_7/S FILL
XAOI22X1_14 AOI22X1_14/A AOI22X1_14/B AOI22X1_14/C INVX1_436/A DFFSR_79/gnd NOR2X1_52/A
+ DFFSR_36/S AOI22X1
XFILL_0_OAI21X1_177 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_21_DFFSR_167 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_3_AOI22X1_2 BUFX2_37/A DFFSR_81/S FILL
XFILL_11_DFFSR_170 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_3_NAND2X1_129 INVX1_4/gnd DFFSR_4/S FILL
XFILL_11_OAI22X1_47 BUFX2_37/A DFFSR_8/S FILL
XFILL_1_INVX1_321 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_6_NOR2X1_46 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_10_OAI22X1_50 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_33_DFFSR_99 BUFX2_35/A DFFSR_97/S FILL
XFILL_10_1_1 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_2_NAND2X1_12 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_7_DFFSR_164 INVX1_89/gnd DFFSR_2/S FILL
XFILL_1_OAI21X1_111 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_44_DFFSR_59 INVX1_4/gnd DFFSR_51/S FILL
XAND2X2_8 AND2X2_8/A AND2X2_8/B BUFX2_5/gnd AND2X2_8/Y DFFSR_23/S AND2X2
XFILL_1_NAND2X1_15 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_8_NAND3X1_71 BUFX2_35/A DFFSR_14/S FILL
XFILL_0_INVX1_141 BUFX2_35/A DFFSR_14/S FILL
XINVX1_251 INVX1_251/A BUFX2_36/A INVX1_251/Y DFFSR_8/S INVX1
XFILL_9_OAI22X1_53 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_0_NAND2X1_18 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_0_DFFSR_56 INVX1_2/gnd DFFSR_51/S FILL
XFILL_17_DFFSR_49 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_2_3 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_7_NAND3X1_74 BUFX2_35/A DFFSR_14/S FILL
XFILL_1_NAND2X1_225 BUFX2_36/A DFFSR_8/S FILL
XFILL_8_OAI22X1_56 BUFX2_37/A DFFSR_8/S FILL
XFILL_4_INVX1_248 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_6_NAND3X1_77 BUFX2_37/A DFFSR_81/S FILL
XFILL_7_OAI22X1_59 INVX1_8/gnd DFFSR_7/S FILL
XNAND3X1_77 NAND3X1_83/A NAND3X1_76/Y XOR2X1_8/A BUFX2_37/A NAND3X1_77/Y DFFSR_81/S
+ NAND3X1
XFILL_5_NAND3X1_80 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_6_OAI22X1_62 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_0_NAND3X1_123 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_4_NAND3X1_83 BUFX2_37/A DFFSR_81/S FILL
XFILL_16_DFFSR_5 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_5_OAI22X1_65 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_2_NAND2X1_159 BUFX2_43/A DFFSR_97/S FILL
XFILL_3_NAND3X1_86 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_51_DFFSR_122 INVX1_94/gnd DFFSR_52/S FILL
XOAI22X1_62 INVX1_382/Y OAI22X1_38/B INVX1_383/Y OAI22X1_38/D BUFX2_8/gnd NOR2X1_40/A
+ DFFSR_25/S OAI22X1
XFILL_11_CLKBUF1_2 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_8_OAI21X1_262 INVX1_89/gnd DFFSR_36/S FILL
XFILL_4_OAI22X1_68 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_41_DFFSR_125 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_2_NAND3X1_89 BUFX2_43/A DFFSR_23/S FILL
XFILL_8_DFFSR_63 INVX1_94/gnd DFFSR_52/S FILL
XFILL_36_DFFSR_16 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_14_DFFSR_96 INVX1_2/gnd DFFSR_1/S FILL
XFILL_25_DFFSR_56 INVX1_2/gnd DFFSR_51/S FILL
XFILL_1_NAND3X1_92 BUFX2_43/A DFFSR_23/S FILL
XFILL_31_DFFSR_128 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_0_NAND3X1_95 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_14_DFFPOSX1_16 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_0_BUFX2_6 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_21_DFFSR_131 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_0_OAI21X1_141 INVX1_94/gnd DFFSR_52/S FILL
XFILL_11_DFFSR_134 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_6_XNOR2X1_1 BUFX2_35/A DFFSR_14/S FILL
XFILL_6_NOR2X1_10 BUFX2_36/A DFFSR_6/S FILL
XFILL_1_INVX1_285 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_37_DFFSR_1 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_11_OAI22X1_11 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_44_DFFSR_23 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_33_DFFSR_63 INVX1_94/gnd DFFSR_52/S FILL
XINVX1_97 INVX1_97/A INVX1_4/gnd INVX1_97/Y DFFSR_4/S INVX1
XFILL_10_OAI22X1_14 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_0_NAND2X1_255 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_48_DFFSR_159 BUFX2_36/A DFFSR_6/S FILL
XFILL_7_DFFSR_128 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_9_NAND3X1_32 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_38_DFFSR_162 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_8_NAND3X1_35 BUFX2_35/A DFFSR_97/S FILL
XFILL_9_OAI22X1_17 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_0_DFFSR_20 DFFSR_89/gnd DFFSR_92/S FILL
XINVX1_215 AND2X2_8/A BUFX2_6/gnd NOR2X1_7/A DFFSR_14/S INVX1
XFILL_7_NAND3X1_38 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_8_OAI22X1_20 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_0_INVX1_105 INVX1_4/gnd DFFSR_51/S FILL
XFILL_17_DFFSR_13 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_28_DFFSR_165 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_6_NAND3X1_41 BUFX2_43/A DFFSR_23/S FILL
XFILL_1_NAND2X1_189 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_4_DFFPOSX1_27 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_7_OAI22X1_23 INVX1_89/gnd DFFSR_2/S FILL
XFILL_4_INVX1_212 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_5_NAND3X1_44 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_18_DFFSR_168 BUFX2_36/A DFFSR_8/S FILL
XFILL_6_OAI22X1_26 INVX1_94/gnd DFFSR_52/S FILL
XXOR2X1_10 XOR2X1_10/A XOR2X1_10/B BUFX2_16/gnd XOR2X1_10/Y DFFSR_11/S XOR2X1
XFILL_4_NAND3X1_47 BUFX2_43/A DFFSR_97/S FILL
XNAND3X1_41 AOI22X1_5/Y NAND3X1_47/B NAND3X1_37/Y BUFX2_43/A AOI22X1_7/C DFFSR_23/S
+ NAND3X1
XFILL_0_AOI22X1_3 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_5_OAI22X1_29 INVX1_8/gnd DFFSR_5/S FILL
XFILL_3_NAND3X1_50 BUFX2_37/A DFFSR_81/S FILL
XOAI22X1_26 INVX1_307/Y OAI22X1_6/B INVX1_308/Y OAI22X1_8/D INVX1_94/gnd NOR2X1_22/A
+ DFFSR_52/S OAI22X1
XFILL_4_OAI22X1_32 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_3_NOR2X1_47 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_41_DFFSR_70 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_8_OAI21X1_226 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_2_NAND2X1_123 BUFX2_6/gnd DFFSR_14/S FILL
XDFFSR_168 BUFX2_14/A CLKBUF1_16/Y DFFSR_175/R DFFSR_8/S DFFSR_168/D BUFX2_36/A DFFSR_8/S
+ DFFSR
XFILL_2_NAND3X1_53 BUFX2_37/A DFFSR_81/S FILL
XFILL_2_INVX1_429 INVX1_89/gnd DFFSR_2/S FILL
XFILL_25_DFFSR_20 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_4_DFFSR_165 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_14_DFFSR_60 BUFX2_37/A DFFSR_8/S FILL
XFILL_3_OAI22X1_35 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_8_DFFSR_27 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_1_NAND3X1_56 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_2_OAI22X1_38 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_45_1_0 INVX1_2/gnd DFFSR_1/S FILL
XFILL_0_OAI21X1_105 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_0_NAND3X1_59 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_1_OAI22X1_41 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_43_3_1 INVX1_4/gnd DFFSR_51/S FILL
XFILL_0_OAI22X1_44 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_1_INVX1_249 BUFX2_35/A DFFSR_14/S FILL
XFILL_49_DFFSR_77 INVX1_89/gnd DFFSR_2/S FILL
XINVX1_61 DFFSR_54/Q BUFX2_7/gnd INVX1_61/Y DFFSR_54/S INVX1
XFILL_0_NAND2X1_219 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_33_DFFSR_27 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_5_DFFSR_74 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_22_DFFSR_67 INVX1_2/gnd DFFSR_51/S FILL
XFILL_41_5_2 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_48_DFFSR_123 DFFSR_89/gnd DFFSR_186/S FILL
XINVX1_179 BUFX2_5/Y BUFX2_5/gnd DFFSR_152/R DFFSR_23/S INVX1
XFILL_38_DFFSR_126 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_9_XOR2X1_4 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_1_NAND2X1_153 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_4_BUFX2_12 BUFX2_37/A DFFSR_81/S FILL
XFILL_28_DFFSR_129 INVX1_2/gnd DFFSR_1/S FILL
XFILL_4_INVX1_176 BUFX2_37/A DFFSR_81/S FILL
XFILL_18_DFFSR_132 INVX1_2/gnd DFFSR_51/S FILL
XFILL_7_OAI21X1_256 INVX1_2/gnd DFFSR_51/S FILL
XFILL_4_DFFSR_4 INVX1_4/gnd DFFSR_4/S FILL
XFILL_3_NOR2X1_11 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_9_NAND3X1_106 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_3_XNOR2X1_2 BUFX2_36/A DFFSR_8/S FILL
XFILL_2_INVX1_68 BUFX2_37/A DFFSR_81/S FILL
XFILL_4_NAND3X1_11 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_41_DFFSR_34 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_30_DFFSR_74 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_8_OAI21X1_190 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_3_NAND3X1_14 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_13_DFFPOSX1_10 INVX1_8/gnd DFFSR_5/S FILL
XDFFSR_132 XOR2X1_13/A CLKBUF1_13/Y DFFSR_135/R DFFSR_51/S DFFSR_132/D INVX1_2/gnd
+ DFFSR_51/S DFFSR
XFILL_2_NAND3X1_17 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_46_4 INVX1_2/gnd DFFSR_1/S FILL
XFILL_2_INVX1_393 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_14_DFFSR_24 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_1_NAND3X1_20 BUFX2_37/A DFFSR_8/S FILL
XFILL_45_DFFSR_160 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_4_DFFSR_129 INVX1_2/gnd DFFSR_1/S FILL
XFILL_0_NAND3X1_23 BUFX2_37/A DFFSR_81/S FILL
XFILL_35_DFFSR_163 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_15_XOR2X1_11 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_28_DFFSR_8 BUFX2_36/A DFFSR_8/S FILL
XFILL_1_INVX1_213 BUFX2_36/A DFFSR_8/S FILL
XFILL_38_DFFSR_81 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_49_DFFSR_41 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_25_DFFSR_166 INVX1_4/gnd DFFSR_51/S FILL
XFILL_15_DFFSR_169 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_7_AOI22X1_1 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_22_DFFSR_31 BUFX2_35/A DFFSR_97/S FILL
XFILL_3_DFFPOSX1_21 BUFX2_5/gnd DFFSR_23/S FILL
XINVX1_25 INVX1_25/A BUFX2_8/gnd INVX1_25/Y DFFSR_25/S INVX1
XFILL_0_NAND2X1_183 INVX1_8/gnd DFFSR_7/S FILL
XFILL_5_DFFSR_38 DFFSR_73/gnd DFFSR_57/S FILL
XDFFSR_78 INVX1_88/A CLKBUF1_5/Y DFFSR_76/R DFFSR_51/S DFFSR_78/D DFFSR_1/gnd DFFSR_1/S
+ DFFSR
XFILL_11_DFFSR_71 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_0_NOR2X1_48 INVX1_89/gnd DFFSR_36/S FILL
XINVX1_143 DFFSR_127/Q BUFX2_5/gnd INVX1_143/Y DFFSR_23/S INVX1
XFILL_1_DFFSR_166 INVX1_4/gnd DFFSR_51/S FILL
XFILL_1_NAND2X1_117 BUFX2_35/A DFFSR_14/S FILL
XFILL_7_OAI21X1_220 BUFX2_43/A DFFSR_97/S FILL
XFILL_15_XOR2X1_1 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_4_INVX1_140 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_49_DFFSR_4 INVX1_4/gnd DFFSR_4/S FILL
XFILL_46_DFFSR_88 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_2_INVX1_32 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_17_1_1 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_2_DFFSR_85 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_30_DFFSR_38 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_19_DFFSR_78 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_8_OAI21X1_154 BUFX2_37/A DFFSR_8/S FILL
XFILL_2_INVX1_357 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_22_DFFPOSX1_29 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_15_3_2 BUFX2_37/A DFFSR_81/S FILL
XFILL_1_BUFX2_23 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_15_CLKBUF1_1 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_45_DFFSR_124 INVX1_89/gnd DFFSR_36/S FILL
XFILL_4_INVX1_6 INVX1_8/gnd DFFSR_5/S FILL
XFILL_35_DFFSR_127 BUFX2_43/A DFFSR_97/S FILL
XFILL_11_NOR3X1_2 INVX1_89/gnd DFFSR_2/S FILL
XFILL_25_DFFSR_130 INVX1_4/gnd DFFSR_51/S FILL
XFILL_15_DFFSR_133 BUFX2_37/A DFFSR_81/S FILL
XFILL_1_INVX1_177 BUFX2_37/A DFFSR_81/S FILL
XFILL_27_DFFSR_85 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_38_DFFSR_45 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_0_NAND2X1_147 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_0_XNOR2X1_3 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_6_OAI21X1_250 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_11_DFFSR_35 DFFSR_5/gnd DFFSR_2/S FILL
XDFFSR_42 INVX1_48/A DFFSR_24/CLK DFFSR_46/R DFFSR_65/S DFFSR_42/D DFFSR_3/gnd DFFSR_65/S
+ DFFSR
XFILL_0_NOR2X1_12 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_8_NAND3X1_100 BUFX2_6/gnd DFFSR_14/S FILL
XINVX1_107 DFFSR_95/Q INVX1_89/gnd INVX1_107/Y DFFSR_36/S INVX1
XFILL_42_DFFSR_161 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_15_DFFSR_2 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_1_DFFSR_130 INVX1_4/gnd DFFSR_51/S FILL
XFILL_35_DFFSR_92 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_4_INVX1_104 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_7_OAI21X1_184 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_46_DFFSR_52 INVX1_94/gnd DFFSR_52/S FILL
XFILL_12_XOR2X1_12 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_32_DFFSR_164 INVX1_89/gnd DFFSR_2/S FILL
XAOI22X1_5 AND2X2_5/Y AND2X2_6/Y AOI22X1_5/C AOI22X1_5/D BUFX2_5/gnd AOI22X1_5/Y DFFSR_6/S
+ AOI22X1
XFILL_22_DFFSR_167 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_19_DFFSR_42 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_2_DFFSR_49 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_4_AOI22X1_2 BUFX2_37/A DFFSR_81/S FILL
XFILL_12_DFFSR_170 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_8_OAI21X1_118 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_2_INVX1_321 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_2_DFFPOSX1_15 BUFX2_35/A DFFSR_14/S FILL
XFILL_43_DFFSR_99 BUFX2_35/A DFFSR_97/S FILL
XFILL_8_DFFSR_164 INVX1_89/gnd DFFSR_2/S FILL
XAND2X2_11 AND2X2_11/A AND2X2_11/B BUFX2_35/A AND2X2_11/Y DFFSR_14/S AND2X2
XFILL_16_DFFSR_89 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_1_INVX1_141 BUFX2_35/A DFFSR_14/S FILL
XFILL_4_AND2X2_8 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_27_DFFSR_49 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_7_NAND3X1_130 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_6_OAI21X1_214 BUFX2_35/A DFFSR_97/S FILL
XFILL_0_NAND2X1_111 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_12_CLKBUF1_2 DFFSR_79/gnd DFFSR_45/S FILL
XOAI21X1_250 DFFSR_45/S INVX1_412/Y NAND2X1_261/Y DFFSR_79/gnd DFFSR_182/D DFFSR_36/S
+ OAI21X1
XFILL_7_OAI21X1_148 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_21_DFFPOSX1_23 INVX1_23/gnd DFFSR_91/S FILL
XFILL_42_DFFSR_125 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_46_DFFSR_16 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_24_DFFSR_96 INVX1_2/gnd DFFSR_1/S FILL
XFILL_35_DFFSR_56 INVX1_2/gnd DFFSR_51/S FILL
XFILL_32_DFFSR_128 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_22_DFFSR_131 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_6_BUFX2_41 BUFX2_37/A DFFSR_81/S FILL
XFILL_12_DFFSR_134 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_48_5_2 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_2_DFFSR_13 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_7_XNOR2X1_1 BUFX2_35/A DFFSR_14/S FILL
XFILL_11_6 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_28_1 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_2_INVX1_285 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_43_DFFSR_63 INVX1_94/gnd DFFSR_52/S FILL
XFILL_49_DFFSR_159 BUFX2_36/A DFFSR_6/S FILL
XFILL_8_DFFSR_128 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_5_OAI21X1_244 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_39_DFFSR_162 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_16_4_0 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_16_DFFSR_53 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_1_INVX1_105 INVX1_4/gnd DFFSR_51/S FILL
XFILL_27_DFFSR_13 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_29_DFFSR_165 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_19_DFFSR_168 BUFX2_36/A DFFSR_8/S FILL
XFILL_15_CLKBUF1_11 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_6_OAI21X1_178 INVX1_94/gnd DFFSR_25/S FILL
XNOR2X1_50 NOR3X1_2/B NOR3X1_2/A INVX1_89/gnd XOR2X1_15/B DFFSR_36/S NOR2X1
XFILL_14_CLKBUF1_14 BUFX2_43/A DFFSR_23/S FILL
XFILL_1_AOI22X1_3 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_3_DFFSR_1 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_13_CLKBUF1_17 INVX1_94/gnd DFFSR_25/S FILL
XFILL_4_NOR2X1_47 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_51_DFFSR_70 BUFX2_17/gnd DFFSR_57/S FILL
XOAI21X1_214 NAND2X1_190/Y XOR2X1_4/A AOI22X1_7/A BUFX2_35/A XNOR2X1_1/A DFFSR_97/S
+ OAI21X1
XFILL_3_INVX1_429 INVX1_89/gnd DFFSR_2/S FILL
XFILL_12_CLKBUF1_20 INVX1_4/gnd DFFSR_51/S FILL
XFILL_35_DFFSR_20 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_5_DFFSR_165 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_24_DFFSR_60 BUFX2_37/A DFFSR_8/S FILL
XFILL_11_CLKBUF1_23 INVX1_89/gnd DFFSR_2/S FILL
XFILL_7_DFFSR_67 INVX1_2/gnd DFFSR_51/S FILL
XFILL_7_OAI21X1_112 INVX1_4/gnd DFFSR_4/S FILL
XFILL_1_OR2X2_1 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_2_INVX1_249 BUFX2_35/A DFFSR_14/S FILL
XFILL_27_DFFSR_5 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_6_NAND3X1_124 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_5_OAI21X1_208 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_4_INVX1_61 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_43_DFFSR_27 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_32_DFFSR_67 INVX1_2/gnd DFFSR_51/S FILL
XFILL_10_DFFPOSX1_28 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_49_DFFSR_123 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_16_DFFSR_17 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_39_DFFSR_126 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_24_1_1 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_29_DFFSR_129 INVX1_2/gnd DFFSR_1/S FILL
XFILL_20_DFFPOSX1_17 BUFX2_37/A DFFSR_8/S FILL
XFILL_6_OAI21X1_142 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_19_DFFSR_132 INVX1_2/gnd DFFSR_51/S FILL
XFILL_6_0_0 BUFX2_35/A DFFSR_14/S FILL
XFILL_48_DFFSR_1 DFFSR_1/gnd DFFSR_1/S FILL
XNOR2X1_14 NOR2X1_14/A OAI22X1_9/Y DFFSR_3/gnd NOR2X1_14/Y DFFSR_4/S NOR2X1
XFILL_4_NOR2X1_11 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_4_XNOR2X1_2 BUFX2_36/A DFFSR_8/S FILL
XFILL_22_3_2 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_40_DFFSR_74 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_4_2_1 BUFX2_6/gnd DFFSR_91/S FILL
XOAI21X1_178 AOI22X1_1/Y NOR2X1_3/Y INVX1_219/A INVX1_94/gnd NAND3X1_5/C DFFSR_25/S
+ OAI21X1
XFILL_7_DFFSR_31 BUFX2_35/A DFFSR_97/S FILL
XFILL_6_NAND2X1_256 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_33_6 INVX1_8/gnd DFFSR_5/S FILL
XFILL_3_INVX1_393 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_24_DFFSR_24 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_2_4_2 INVX1_23/gnd DFFSR_186/S FILL
XFILL_46_DFFSR_160 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_5_DFFSR_129 INVX1_2/gnd DFFSR_1/S FILL
XFILL_13_DFFSR_64 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_4_OAI21X1_238 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_3_INVX1_3 INVX1_8/gnd DFFSR_5/S FILL
XFILL_36_DFFSR_163 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_2_INVX1_213 BUFX2_36/A DFFSR_8/S FILL
XFILL_48_DFFSR_81 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_0_XOR2X1_1 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_26_DFFSR_166 INVX1_4/gnd DFFSR_51/S FILL
XFILL_16_DFFSR_169 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_8_AOI22X1_1 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_4_INVX1_25 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_4_DFFSR_78 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_32_DFFSR_31 BUFX2_35/A DFFSR_97/S FILL
XFILL_5_OAI21X1_172 BUFX2_36/A DFFSR_6/S FILL
XFILL_21_DFFSR_71 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_1_NOR2X1_48 INVX1_89/gnd DFFSR_36/S FILL
XFILL_0_INVX1_430 INVX1_89/gnd DFFSR_36/S FILL
XNAND3X1_124 INVX1_332/A INVX1_333/Y INVX1_331/Y DFFSR_5/gnd OAI22X1_39/D DFFSR_5/S
+ NAND3X1
XFILL_2_DFFSR_166 INVX1_4/gnd DFFSR_51/S FILL
XFILL_3_BUFX2_16 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_8_XOR2X1_8 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_3_CLKBUF1_11 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_5_NAND2X1_286 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_2_CLKBUF1_14 BUFX2_43/A DFFSR_23/S FILL
XFILL_6_OAI21X1_106 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_1_CLKBUF1_17 INVX1_94/gnd DFFSR_25/S FILL
XOAI21X1_142 DFFSR_54/S INVX1_160/Y OAI21X1_142/C BUFX2_19/gnd DFFSR_142/D DFFSR_52/S
+ OAI21X1
XFILL_40_DFFSR_38 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_29_DFFSR_78 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_0_CLKBUF1_20 INVX1_4/gnd DFFSR_51/S FILL
XFILL_1_INVX1_72 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_6_NAND2X1_220 BUFX2_35/A DFFSR_14/S FILL
XFILL_3_INVX1_357 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_13_DFFSR_28 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_16_CLKBUF1_1 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_5_NAND3X1_118 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_46_DFFSR_124 INVX1_89/gnd DFFSR_36/S FILL
XFILL_36_DFFSR_127 BUFX2_43/A DFFSR_97/S FILL
XNAND2X1_256 DFFSR_5/S din[1] DFFSR_5/gnd OAI21X1_245/C DFFSR_2/S NAND2X1
XFILL_4_OAI21X1_202 BUFX2_35/A DFFSR_14/S FILL
XFILL_26_DFFSR_130 INVX1_4/gnd DFFSR_51/S FILL
XFILL_16_DFFSR_133 BUFX2_37/A DFFSR_81/S FILL
XFILL_2_INVX1_177 BUFX2_37/A DFFSR_81/S FILL
XFILL_37_DFFSR_85 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_48_DFFSR_45 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_1_XNOR2X1_3 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_21_DFFSR_35 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_5_OAI21X1_136 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_10_DFFSR_75 INVX1_4/gnd DFFSR_51/S FILL
XFILL_19_DFFPOSX1_11 INVX1_4/gnd DFFSR_4/S FILL
XFILL_4_DFFSR_42 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_1_NOR2X1_12 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_0_INVX1_394 INVX1_89/gnd DFFSR_2/S FILL
XFILL_43_DFFSR_161 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_14_XOR2X1_5 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_2_DFFSR_130 INVX1_4/gnd DFFSR_51/S FILL
XFILL_45_DFFSR_92 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_39_DFFSR_8 BUFX2_36/A DFFSR_8/S FILL
XFILL_26_DFFPOSX1_2 INVX1_89/gnd DFFSR_36/S FILL
XFILL_5_NAND2X1_250 INVX1_8/gnd DFFSR_5/S FILL
XFILL_13_XOR2X1_12 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_33_DFFSR_164 INVX1_89/gnd DFFSR_2/S FILL
XFILL_25_DFFPOSX1_5 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_1_DFFSR_89 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_6_AND2X2_1 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_24_DFFPOSX1_8 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_23_DFFSR_167 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_18_DFFSR_82 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_1_INVX1_36 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_29_DFFSR_42 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_3_OAI21X1_232 BUFX2_35/A DFFSR_97/S FILL
XFILL_5_AOI22X1_2 BUFX2_37/A DFFSR_81/S FILL
XFILL_13_DFFSR_170 BUFX2_7/gnd DFFSR_81/S FILL
XOAI21X1_106 BUFX2_24/Y INVX1_120/Y OAI21X1_106/C DFFSR_1/gnd DFFSR_106/D DFFSR_9/S
+ OAI21X1
XFILL_9_DFFPOSX1_22 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_6_NAND2X1_184 BUFX2_37/A DFFSR_8/S FILL
XFILL_3_INVX1_321 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_0_BUFX2_27 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_23_4_0 BUFX2_8/gnd DFFSR_10/S FILL
XNAND2X1_220 AND2X2_11/Y XNOR2X1_1/A BUFX2_35/A INVX1_253/A DFFSR_14/S NAND2X1
XFILL_9_DFFSR_164 INVX1_89/gnd DFFSR_2/S FILL
XFILL_4_OAI21X1_166 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_26_DFFSR_89 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_2_INVX1_141 BUFX2_35/A DFFSR_14/S FILL
XFILL_9_DFFSR_96 INVX1_2/gnd DFFSR_1/S FILL
XFILL_37_DFFSR_49 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_3_5_0 INVX1_23/gnd DFFSR_91/S FILL
XFILL_5_OAI21X1_100 INVX1_23/gnd DFFSR_91/S FILL
XFILL_10_DFFSR_39 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_4_NAND2X1_280 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_0_INVX1_358 INVX1_89/gnd DFFSR_36/S FILL
XFILL_13_CLKBUF1_2 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_43_DFFSR_125 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_5_NAND2X1_214 BUFX2_35/A DFFSR_97/S FILL
XFILL_2_OAI21X1_262 INVX1_89/gnd DFFSR_36/S FILL
XFILL_34_DFFSR_96 INVX1_2/gnd DFFSR_1/S FILL
XFILL_45_DFFSR_56 INVX1_2/gnd DFFSR_51/S FILL
XFILL_33_DFFSR_128 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_4_NAND3X1_112 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_23_DFFSR_131 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_18_DFFSR_46 BUFX2_36/A DFFSR_6/S FILL
XFILL_1_DFFSR_53 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_13_DFFSR_134 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_6_NAND2X1_148 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_8_XNOR2X1_1 BUFX2_35/A DFFSR_14/S FILL
XFILL_3_OAI21X1_196 INVX1_94/gnd DFFSR_25/S FILL
XFILL_3_INVX1_285 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_50_DFFSR_159 BUFX2_36/A DFFSR_6/S FILL
XNAND2X1_184 AND2X2_11/A AND2X2_9/B BUFX2_37/A INVX1_224/A DFFSR_8/S NAND2X1
XFILL_9_DFFSR_128 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_26_DFFSR_2 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_31_1_1 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_4_OAI21X1_130 INVX1_4/gnd DFFSR_4/S FILL
XFILL_40_DFFSR_162 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_9_DFFSR_60 BUFX2_37/A DFFSR_8/S FILL
XFILL_26_DFFSR_53 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_29_3_2 INVX1_89/gnd DFFSR_2/S FILL
XFILL_10_XOR2X1_13 INVX1_8/gnd DFFSR_7/S FILL
XFILL_15_DFFSR_93 INVX1_2/gnd DFFSR_51/S FILL
XFILL_2_INVX1_105 INVX1_4/gnd DFFSR_51/S FILL
XFILL_37_DFFSR_13 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_30_DFFSR_165 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_20_DFFSR_168 BUFX2_36/A DFFSR_8/S FILL
XFILL_4_NAND2X1_244 INVX1_94/gnd DFFSR_52/S FILL
XFILL_9_4_2 BUFX2_43/A DFFSR_23/S FILL
XFILL_2_AOI22X1_3 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_10_DFFSR_171 BUFX2_19/gnd DFFSR_52/S FILL
XINVX1_432 DFFSR_135/Q DFFSR_71/gnd INVX1_432/Y DFFSR_45/S INVX1
XFILL_0_INVX1_322 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_5_NOR2X1_47 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_2_OAI21X1_226 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_14_DFFPOSX1_2 INVX1_89/gnd DFFSR_36/S FILL
XFILL_4_INVX1_429 INVX1_89/gnd DFFSR_2/S FILL
XFILL_45_DFFSR_20 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_8_DFFPOSX1_16 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_6_DFFSR_165 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_34_DFFSR_60 BUFX2_37/A DFFSR_8/S FILL
XFILL_5_NAND2X1_178 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_13_DFFPOSX1_5 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_12_DFFPOSX1_8 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_18_DFFSR_10 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_1_DFFSR_17 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_3_OAI21X1_160 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_3_INVX1_249 BUFX2_35/A DFFSR_14/S FILL
XFILL_6_NAND2X1_112 INVX1_4/gnd DFFSR_4/S FILL
XNAND2X1_148 INVX1_168/A DFFSR_186/S DFFSR_89/gnd NAND2X1_148/Y DFFSR_92/S NAND2X1
XFILL_9_AOI21X1_37 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_42_DFFSR_67 INVX1_2/gnd DFFSR_51/S FILL
XFILL_50_DFFSR_123 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_27_DFFPOSX1_24 BUFX2_43/A DFFSR_23/S FILL
XFILL_10_CLKBUF1_3 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_3_NAND2X1_274 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_8_AOI21X1_40 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_26_DFFSR_17 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_7_AOI21X1_43 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_40_DFFSR_126 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_15_DFFSR_57 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_9_DFFSR_24 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_6_AOI21X1_46 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_30_DFFSR_129 INVX1_2/gnd DFFSR_1/S FILL
XFILL_20_DFFSR_132 INVX1_2/gnd DFFSR_51/S FILL
XFILL_1_OAI21X1_256 INVX1_2/gnd DFFSR_51/S FILL
XFILL_10_DFFSR_135 BUFX2_43/A DFFSR_97/S FILL
XFILL_4_NAND2X1_208 BUFX2_8/gnd DFFSR_10/S FILL
XAOI21X1_46 AND2X2_17/A AND2X2_17/B AOI21X1_46/C DFFSR_5/gnd AOI21X1_46/Y DFFSR_5/S
+ AOI21X1
XFILL_5_NOR2X1_11 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_3_NAND3X1_106 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_5_XNOR2X1_2 BUFX2_36/A DFFSR_8/S FILL
XINVX1_396 BUFX2_8/Y DFFSR_5/gnd INVX1_396/Y DFFSR_5/S INVX1
XFILL_50_DFFSR_74 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_0_INVX1_286 INVX1_4/gnd DFFSR_51/S FILL
XFILL_20_8 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_2_OAI21X1_190 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_6_DFFSR_71 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_5_NAND2X1_142 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_34_DFFSR_24 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_47_DFFSR_160 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_6_DFFSR_129 INVX1_2/gnd DFFSR_1/S FILL
XFILL_23_DFFSR_64 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_37_DFFSR_163 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_3_INVX1_213 BUFX2_36/A DFFSR_8/S FILL
XFILL_9_OAI21X1_85 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_3_OAI21X1_124 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_27_DFFSR_166 INVX1_4/gnd DFFSR_51/S FILL
XFILL_17_DFFSR_169 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_9_AOI22X1_1 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_17_DFFSR_9 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_8_OAI21X1_88 INVX1_4/gnd DFFSR_4/S FILL
XFILL_7_OAI21X1_91 BUFX2_43/A DFFSR_97/S FILL
XFILL_42_DFFSR_31 BUFX2_35/A DFFSR_97/S FILL
XFILL_31_DFFSR_71 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_3_NAND2X1_238 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_2_NOR2X1_48 INVX1_89/gnd DFFSR_36/S FILL
XNAND2X1_112 BUFX2_15/Y INVX1_392/A INVX1_4/gnd OAI21X1_112/C DFFSR_4/S NAND2X1
XFILL_6_OAI21X1_94 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_3_INVX1_65 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_5_OAI21X1_97 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_1_INVX1_430 INVX1_89/gnd DFFSR_36/S FILL
XFILL_15_DFFSR_21 INVX1_2/gnd DFFSR_1/S FILL
XFILL_3_DFFSR_166 INVX1_4/gnd DFFSR_51/S FILL
XOAI21X1_94 BUFX2_16/Y INVX1_106/Y NAND2X1_94/Y BUFX2_16/gnd DFFSR_94/D DFFSR_11/S
+ OAI21X1
XFILL_6_AOI21X1_10 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_1_OAI21X1_220 BUFX2_43/A DFFSR_97/S FILL
XFILL_4_NAND2X1_172 BUFX2_36/A DFFSR_6/S FILL
XFILL_6_NOR3X1_2 INVX1_89/gnd DFFSR_2/S FILL
XFILL_7_DFFPOSX1_10 INVX1_8/gnd DFFSR_5/S FILL
XFILL_5_AOI21X1_13 INVX1_8/gnd DFFSR_7/S FILL
XFILL_4_AOI21X1_16 BUFX2_43/A DFFSR_23/S FILL
XFILL_38_DFFSR_5 DFFSR_5/gnd DFFSR_5/S FILL
XAOI21X1_10 INVX1_234/Y INVX1_221/A NOR2X1_5/B BUFX2_17/gnd AOI21X1_10/Y DFFSR_57/S
+ AOI21X1
XINVX1_360 DFFSR_100/Q BUFX2_7/gnd INVX1_360/Y DFFSR_81/S INVX1
XFILL_3_AOI21X1_19 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_0_INVX1_250 INVX1_94/gnd DFFSR_25/S FILL
XFILL_2_DFFPOSX1_2 INVX1_89/gnd DFFSR_36/S FILL
XFILL_30_4_0 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_50_DFFSR_38 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_39_DFFSR_78 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_2_AOI21X1_22 BUFX2_43/A DFFSR_97/S FILL
XFILL_2_OAI21X1_154 BUFX2_37/A DFFSR_8/S FILL
XFILL_16_DFFPOSX1_29 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_1_DFFPOSX1_5 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_12_DFFSR_68 BUFX2_35/A DFFSR_14/S FILL
XFILL_1_AOI21X1_25 BUFX2_43/A DFFSR_97/S FILL
XFILL_23_DFFSR_28 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_17_CLKBUF1_1 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_0_DFFPOSX1_8 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_6_DFFSR_35 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_5_NAND2X1_106 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_0_AOI21X1_28 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_47_DFFSR_124 INVX1_89/gnd DFFSR_36/S FILL
XFILL_37_DFFSR_127 BUFX2_43/A DFFSR_97/S FILL
XFILL_2_NAND2X1_268 BUFX2_37/A DFFSR_8/S FILL
XBUFX2_13 BUFX2_14/A BUFX2_7/gnd BUFX2_13/Y DFFSR_54/S BUFX2
XFILL_27_DFFSR_130 INVX1_4/gnd DFFSR_51/S FILL
XFILL_9_OAI21X1_49 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_26_DFFPOSX1_18 BUFX2_37/A DFFSR_8/S FILL
XFILL_17_DFFSR_133 BUFX2_37/A DFFSR_81/S FILL
XFILL_3_INVX1_177 BUFX2_37/A DFFSR_81/S FILL
XFILL_47_DFFSR_85 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_8_OAI21X1_52 INVX1_94/gnd DFFSR_25/S FILL
XFILL_2_XNOR2X1_3 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_3_INVX1_29 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_0_OAI21X1_250 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_7_OAI21X1_55 INVX1_89/gnd DFFSR_2/S FILL
XFILL_31_DFFSR_35 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_3_DFFSR_82 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_20_DFFSR_75 INVX1_4/gnd DFFSR_51/S FILL
XFILL_2_NOR2X1_12 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_6_NAND2X1_73 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_3_NAND2X1_202 BUFX2_35/A DFFSR_97/S FILL
XFILL_5_NAND2X1_76 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_6_OAI21X1_58 DFFSR_3/gnd DFFSR_65/S FILL
XNAND2X1_73 DFFSR_65/Q BUFX2_16/Y DFFSR_73/gnd OAI21X1_73/C DFFSR_11/S NAND2X1
XFILL_5_OAI21X1_61 BUFX2_36/A DFFSR_8/S FILL
XFILL_4_NAND2X1_79 INVX1_89/gnd DFFSR_36/S FILL
XFILL_1_INVX1_394 INVX1_89/gnd DFFSR_2/S FILL
XOAI21X1_58 DFFSR_4/S INVX1_66/Y NAND2X1_58/Y DFFSR_3/gnd DFFSR_58/D DFFSR_65/S OAI21X1
XFILL_2_NAND3X1_100 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_2_BUFX2_20 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_3_NAND2X1_82 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_3_DFFSR_130 INVX1_4/gnd DFFSR_51/S FILL
XFILL_4_OAI21X1_64 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_44_DFFSR_161 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_10_AOI22X1_8 BUFX2_43/A DFFSR_97/S FILL
XFILL_1_OAI21X1_184 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_2_NAND2X1_85 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_14_XOR2X1_12 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_3_OAI21X1_67 INVX1_2/gnd DFFSR_1/S FILL
XFILL_34_DFFSR_164 INVX1_89/gnd DFFSR_2/S FILL
XFILL_4_NAND2X1_136 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_1_NAND2X1_88 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_2_OAI21X1_70 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_0_NAND2X1_91 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_0_INVX1_214 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_24_DFFSR_167 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_28_DFFSR_82 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_0_INVX1_76 INVX1_2/gnd DFFSR_1/S FILL
XFILL_39_DFFSR_42 DFFSR_3/gnd DFFSR_65/S FILL
XINVX1_324 INVX1_54/A BUFX2_16/gnd INVX1_324/Y DFFSR_11/S INVX1
XFILL_1_OAI21X1_73 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_6_AOI22X1_2 BUFX2_37/A DFFSR_81/S FILL
XFILL_14_DFFSR_170 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_0_OAI21X1_76 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_38_1_1 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_4_INVX1_321 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_2_OAI21X1_118 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_36_3_2 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_12_DFFSR_32 INVX1_2/gnd DFFSR_1/S FILL
XFILL_5_DFFSR_8 BUFX2_36/A DFFSR_8/S FILL
XFILL_2_NAND2X1_232 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_0_DFFSR_167 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_36_DFFSR_89 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_3_INVX1_141 BUFX2_35/A DFFSR_14/S FILL
XFILL_9_OAI21X1_13 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_47_DFFSR_49 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_1_NAND3X1_130 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_8_OAI21X1_16 INVX1_89/gnd DFFSR_36/S FILL
XFILL_6_NAND2X1_37 INVX1_8/gnd DFFSR_5/S FILL
XFILL_7_OAI21X1_19 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_0_OAI21X1_214 BUFX2_35/A DFFSR_97/S FILL
XFILL_3_DFFSR_46 BUFX2_36/A DFFSR_6/S FILL
XFILL_6_OAI21X1_22 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_20_DFFSR_39 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_3_NAND2X1_166 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_5_NAND2X1_40 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_5_OAI21X1_25 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_1_INVX1_358 INVX1_89/gnd DFFSR_36/S FILL
XFILL_4_NAND2X1_43 INVX1_89/gnd DFFSR_2/S FILL
XNAND2X1_37 DFFSR_7/S INVX1_33/A INVX1_8/gnd OAI21X1_37/C DFFSR_5/S NAND2X1
XFILL_4_OAI21X1_28 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_3_NAND2X1_46 BUFX2_8/gnd DFFSR_25/S FILL
XOAI21X1_22 DFFSR_25/S INVX1_25/Y NAND2X1_22/Y BUFX2_8/gnd DFFSR_22/D DFFSR_25/S OAI21X1
XFILL_14_CLKBUF1_2 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_15_DFFPOSX1_23 INVX1_23/gnd DFFSR_91/S FILL
XFILL_44_DFFSR_125 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_3_OAI21X1_31 BUFX2_35/A DFFSR_97/S FILL
XFILL_13_XOR2X1_9 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_2_NAND2X1_49 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_1_OAI21X1_148 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_4_NAND2X1_100 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_34_DFFSR_128 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_1_NAND2X1_52 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_44_DFFSR_96 INVX1_2/gnd DFFSR_1/S FILL
XFILL_2_OAI21X1_34 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_5_AND2X2_5 BUFX2_37/A DFFSR_81/S FILL
XFILL_1_OAI21X1_37 INVX1_89/gnd DFFSR_2/S FILL
XFILL_0_NAND2X1_55 INVX1_89/gnd DFFSR_2/S FILL
XFILL_24_DFFSR_131 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_0_INVX1_178 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_28_DFFSR_46 BUFX2_36/A DFFSR_6/S FILL
XFILL_14_DFFSR_134 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_0_INVX1_40 INVX1_8/gnd DFFSR_5/S FILL
XFILL_17_DFFSR_86 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_0_DFFSR_93 INVX1_2/gnd DFFSR_51/S FILL
XINVX1_288 DFFSR_43/Q INVX1_4/gnd INVX1_288/Y DFFSR_4/S INVX1
XFILL_1_NAND2X1_262 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_9_XNOR2X1_1 BUFX2_35/A DFFSR_14/S FILL
XFILL_0_OAI21X1_40 INVX1_8/gnd DFFSR_7/S FILL
XFILL_25_DFFPOSX1_12 INVX1_8/gnd DFFSR_5/S FILL
XFILL_7_AOI22X1_12 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_50_DFFSR_8 BUFX2_36/A DFFSR_8/S FILL
XFILL_2_NAND2X1_196 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_0_DFFSR_131 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_41_DFFSR_162 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_36_DFFSR_53 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_11_XOR2X1_13 INVX1_8/gnd DFFSR_7/S FILL
XFILL_25_DFFSR_93 INVX1_2/gnd DFFSR_51/S FILL
XFILL_3_INVX1_105 INVX1_4/gnd DFFSR_51/S FILL
XFILL_47_DFFSR_13 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_31_DFFSR_165 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_21_DFFSR_168 BUFX2_36/A DFFSR_8/S FILL
XFILL_0_OAI21X1_178 INVX1_94/gnd DFFSR_25/S FILL
XFILL_3_DFFSR_10 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_9_OAI21X1_233 BUFX2_36/A DFFSR_8/S FILL
XFILL_3_AOI22X1_3 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_11_DFFSR_171 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_3_NAND2X1_130 INVX1_4/gnd DFFSR_4/S FILL
XFILL_11_OAI22X1_48 BUFX2_37/A DFFSR_81/S FILL
XFILL_1_INVX1_322 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_6_NOR2X1_47 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_3_NAND2X1_10 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_7_DFFSR_165 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_10_1_2 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_44_DFFSR_60 BUFX2_37/A DFFSR_8/S FILL
XFILL_10_OAI22X1_51 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_1_OAI21X1_112 INVX1_4/gnd DFFSR_4/S FILL
XFILL_2_NAND2X1_13 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_9_NAND3X1_69 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_1_NAND2X1_16 DFFSR_79/gnd DFFSR_36/S FILL
XAND2X2_9 AND2X2_9/A AND2X2_9/B BUFX2_6/gnd AND2X2_9/Y DFFSR_14/S AND2X2
XFILL_8_NAND3X1_72 BUFX2_5/gnd DFFSR_23/S FILL
XINVX1_252 XOR2X1_8/A BUFX2_36/A INVX1_252/Y DFFSR_6/S INVX1
XFILL_9_OAI22X1_54 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_28_DFFSR_10 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_0_INVX1_142 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_0_DFFSR_57 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_0_NAND2X1_19 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_17_DFFSR_50 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_2_4 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_7_NAND3X1_75 BUFX2_35/A DFFSR_97/S FILL
XFILL_8_OAI22X1_57 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_1_NAND2X1_226 BUFX2_36/A DFFSR_6/S FILL
XFILL_6_NAND3X1_78 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_7_OAI22X1_60 INVX1_8/gnd DFFSR_5/S FILL
XFILL_5_NAND3X1_81 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_6_OAI22X1_63 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_0_NAND3X1_124 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_16_DFFSR_6 BUFX2_5/gnd DFFSR_6/S FILL
XNAND3X1_78 NAND3X1_71/Y NAND3X1_70/Y AOI21X1_27/Y BUFX2_19/gnd NAND3X1_83/B DFFSR_54/S
+ NAND3X1
XFILL_4_NAND3X1_84 INVX1_94/gnd DFFSR_25/S FILL
XFILL_5_OAI22X1_66 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_3_NAND3X1_87 INVX1_94/gnd DFFSR_52/S FILL
XOAI22X1_63 INVX1_385/Y OAI22X1_39/B INVX1_384/Y OAI22X1_39/D BUFX2_8/gnd NOR2X1_41/B
+ DFFSR_10/S OAI22X1
XFILL_11_CLKBUF1_3 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_2_NAND2X1_160 INVX1_8/gnd DFFSR_5/S FILL
XFILL_2_NAND3X1_90 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_36_DFFSR_17 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_8_OAI21X1_263 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_41_DFFSR_126 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_25_DFFSR_57 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_8_DFFSR_64 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_14_DFFSR_97 BUFX2_35/A DFFSR_97/S FILL
XFILL_1_NAND3X1_93 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_31_DFFSR_129 INVX1_2/gnd DFFSR_1/S FILL
XFILL_37_4_0 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_0_NAND3X1_96 BUFX2_43/A DFFSR_97/S FILL
XFILL_0_BUFX2_7 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_21_DFFSR_132 INVX1_2/gnd DFFSR_51/S FILL
XFILL_11_DFFSR_135 BUFX2_43/A DFFSR_97/S FILL
XFILL_14_DFFPOSX1_17 BUFX2_37/A DFFSR_8/S FILL
XFILL_0_OAI21X1_142 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_6_NOR2X1_11 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_6_XNOR2X1_2 BUFX2_36/A DFFSR_8/S FILL
XFILL_1_INVX1_286 INVX1_4/gnd DFFSR_51/S FILL
XFILL_37_DFFSR_2 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_11_OAI22X1_12 INVX1_4/gnd DFFSR_51/S FILL
XFILL_0_NAND2X1_256 DFFSR_5/gnd DFFSR_2/S FILL
XINVX1_98 DFFSR_87/Q INVX1_4/gnd INVX1_98/Y DFFSR_4/S INVX1
XFILL_10_OAI22X1_15 INVX1_4/gnd DFFSR_4/S FILL
XFILL_44_DFFSR_24 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_9_NAND3X1_33 INVX1_8/gnd DFFSR_7/S FILL
XFILL_7_DFFSR_129 INVX1_2/gnd DFFSR_1/S FILL
XFILL_33_DFFSR_64 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_8_NAND3X1_36 BUFX2_35/A DFFSR_97/S FILL
XFILL_9_OAI22X1_18 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_48_DFFSR_160 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_17_DFFSR_14 BUFX2_35/A DFFSR_14/S FILL
XFILL_7_NAND3X1_39 BUFX2_5/gnd DFFSR_23/S FILL
XINVX1_216 AND2X2_6/A BUFX2_36/A INVX1_216/Y DFFSR_6/S INVX1
XFILL_0_DFFSR_21 INVX1_2/gnd DFFSR_1/S FILL
XFILL_38_DFFSR_163 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_0_INVX1_106 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_8_OAI22X1_21 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_1_NAND2X1_190 BUFX2_35/A DFFSR_97/S FILL
XFILL_6_NAND3X1_42 BUFX2_43/A DFFSR_23/S FILL
XFILL_4_INVX1_213 BUFX2_36/A DFFSR_8/S FILL
XFILL_7_OAI22X1_24 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_28_DFFSR_166 INVX1_4/gnd DFFSR_51/S FILL
XFILL_4_DFFPOSX1_28 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_5_NAND3X1_45 BUFX2_35/A DFFSR_97/S FILL
XFILL_18_DFFSR_169 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_6_OAI22X1_27 DFFSR_79/gnd DFFSR_36/S FILL
XXOR2X1_11 XOR2X1_11/A XOR2X1_11/B DFFSR_73/gnd XOR2X1_12/B DFFSR_57/S XOR2X1
XFILL_4_NAND3X1_48 BUFX2_43/A DFFSR_23/S FILL
XNAND3X1_42 INVX1_241/A NAND3X1_37/B NAND3X1_37/C BUFX2_43/A NAND3X1_42/Y DFFSR_23/S
+ NAND3X1
XFILL_0_AOI22X1_4 INVX1_94/gnd DFFSR_25/S FILL
XFILL_5_OAI22X1_30 INVX1_94/gnd DFFSR_25/S FILL
XFILL_41_DFFSR_71 DFFSR_71/gnd DFFSR_10/S FILL
XOAI22X1_27 INVX1_310/Y OAI22X1_7/B INVX1_309/Y OAI22X1_7/D DFFSR_79/gnd NOR2X1_23/A
+ DFFSR_36/S OAI22X1
XFILL_3_NOR2X1_48 INVX1_89/gnd DFFSR_36/S FILL
XFILL_8_OAI21X1_227 BUFX2_5/gnd DFFSR_23/S FILL
XDFFSR_169 AND2X2_6/A CLKBUF1_16/Y DFFSR_175/R DFFSR_6/S DFFSR_169/D BUFX2_5/gnd DFFSR_6/S
+ DFFSR
XFILL_3_NAND3X1_51 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_2_NAND2X1_124 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_2_INVX1_430 INVX1_89/gnd DFFSR_36/S FILL
XFILL_4_OAI22X1_33 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_14_DFFSR_61 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_2_NAND3X1_54 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_8_DFFSR_28 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_3_OAI22X1_36 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_25_DFFSR_21 INVX1_2/gnd DFFSR_1/S FILL
XFILL_4_DFFSR_166 INVX1_4/gnd DFFSR_51/S FILL
XFILL_2_OAI22X1_39 BUFX2_37/A DFFSR_8/S FILL
XFILL_1_NAND3X1_57 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_45_1_1 INVX1_2/gnd DFFSR_1/S FILL
XFILL_0_AND2X2_10 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_0_NAND3X1_60 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_1_OAI22X1_42 INVX1_8/gnd DFFSR_7/S FILL
XFILL_0_OAI21X1_106 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_0_OAI22X1_45 INVX1_89/gnd DFFSR_2/S FILL
XFILL_43_3_2 INVX1_4/gnd DFFSR_51/S FILL
XFILL_1_INVX1_250 INVX1_94/gnd DFFSR_25/S FILL
XFILL_49_DFFSR_78 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_0_NAND2X1_220 BUFX2_35/A DFFSR_14/S FILL
XFILL_22_DFFSR_68 BUFX2_35/A DFFSR_14/S FILL
XFILL_33_DFFSR_28 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_18_CLKBUF1_1 BUFX2_8/gnd DFFSR_25/S FILL
XINVX1_62 DFFSR_55/Q INVX1_89/gnd INVX1_62/Y DFFSR_2/S INVX1
XFILL_5_DFFSR_75 INVX1_4/gnd DFFSR_51/S FILL
XFILL_48_DFFSR_124 INVX1_89/gnd DFFSR_36/S FILL
XFILL_38_DFFSR_127 BUFX2_43/A DFFSR_97/S FILL
XINVX1_180 DFFSR_153/Q BUFX2_37/A INVX1_180/Y DFFSR_8/S INVX1
XFILL_9_XOR2X1_5 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_4_BUFX2_13 BUFX2_7/gnd DFFSR_54/S FILL
XCLKBUF1_1 DFFSR_149/Q BUFX2_8/gnd CLKBUF1_1/Y DFFSR_25/S CLKBUF1
XFILL_28_DFFSR_130 INVX1_4/gnd DFFSR_51/S FILL
XFILL_11_2_0 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_1_NAND2X1_154 BUFX2_37/A DFFSR_8/S FILL
XFILL_18_DFFSR_133 BUFX2_37/A DFFSR_81/S FILL
XFILL_4_INVX1_177 BUFX2_37/A DFFSR_81/S FILL
XFILL_4_DFFSR_5 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_7_OAI21X1_257 INVX1_2/gnd DFFSR_51/S FILL
XFILL_3_XNOR2X1_3 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_2_INVX1_69 BUFX2_36/A DFFSR_8/S FILL
XFILL_4_NAND3X1_12 INVX1_94/gnd DFFSR_52/S FILL
XFILL_41_DFFSR_35 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_30_DFFSR_75 INVX1_4/gnd DFFSR_51/S FILL
XFILL_3_NOR2X1_12 BUFX2_16/gnd DFFSR_65/S FILL
XDFFSR_133 DFFSR_133/Q CLKBUF1_11/Y DFFSR_135/R DFFSR_8/S DFFSR_133/D BUFX2_37/A DFFSR_81/S
+ DFFSR
XFILL_3_NAND3X1_15 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_13_DFFPOSX1_11 INVX1_4/gnd DFFSR_4/S FILL
XFILL_8_OAI21X1_191 BUFX2_37/A DFFSR_8/S FILL
XFILL_2_INVX1_394 INVX1_89/gnd DFFSR_2/S FILL
XFILL_2_NAND3X1_18 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_1_NAND3X1_21 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_14_DFFSR_25 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_4_DFFSR_130 INVX1_4/gnd DFFSR_51/S FILL
XFILL_45_DFFSR_161 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_0_NAND3X1_24 BUFX2_37/A DFFSR_8/S FILL
XFILL_15_XOR2X1_12 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_35_DFFSR_164 INVX1_89/gnd DFFSR_2/S FILL
XFILL_28_DFFSR_9 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_1_INVX1_214 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_25_DFFSR_167 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_38_DFFSR_82 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_49_DFFSR_42 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_7_AOI22X1_2 BUFX2_37/A DFFSR_81/S FILL
XFILL_15_DFFSR_170 BUFX2_7/gnd DFFSR_81/S FILL
XINVX1_26 INVX1_26/A BUFX2_43/A INVX1_26/Y DFFSR_23/S INVX1
XFILL_0_NAND2X1_184 BUFX2_37/A DFFSR_8/S FILL
XFILL_5_DFFSR_39 DFFSR_79/gnd DFFSR_45/S FILL
XDFFSR_79 DFFSR_79/Q CLKBUF1_1/Y DFFSR_76/R DFFSR_36/S DFFSR_79/D DFFSR_79/gnd DFFSR_36/S
+ DFFSR
XFILL_3_DFFPOSX1_22 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_0_NOR2X1_49 INVX1_89/gnd DFFSR_36/S FILL
XFILL_11_DFFSR_72 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_22_DFFSR_32 INVX1_2/gnd DFFSR_1/S FILL
XINVX1_144 DFFSR_128/Q BUFX2_8/gnd INVX1_144/Y DFFSR_25/S INVX1
XFILL_1_DFFSR_167 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_46_DFFSR_89 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_7_OAI21X1_221 BUFX2_35/A DFFSR_14/S FILL
XFILL_4_INVX1_141 BUFX2_35/A DFFSR_14/S FILL
XFILL_15_XOR2X1_2 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_49_DFFSR_5 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_1_NAND2X1_118 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_17_1_2 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_30_DFFSR_39 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_19_DFFSR_79 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_2_DFFSR_86 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_2_INVX1_33 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_22_DFFPOSX1_30 BUFX2_43/A DFFSR_97/S FILL
XFILL_8_OAI21X1_155 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_2_INVX1_358 INVX1_89/gnd DFFSR_36/S FILL
XFILL_15_CLKBUF1_2 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_45_DFFSR_125 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_4_INVX1_7 BUFX2_36/A DFFSR_8/S FILL
XFILL_1_BUFX2_24 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_35_DFFSR_128 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_25_DFFSR_131 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_1_INVX1_178 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_38_DFFSR_46 BUFX2_36/A DFFSR_6/S FILL
XFILL_15_DFFSR_134 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_27_DFFSR_86 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_6_OAI21X1_251 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_0_NAND2X1_148 DFFSR_89/gnd DFFSR_92/S FILL
XDFFSR_43 DFFSR_43/Q DFFSR_52/CLK DFFSR_46/R DFFSR_25/S DFFSR_43/D INVX1_94/gnd DFFSR_25/S
+ DFFSR
XFILL_11_DFFSR_36 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_0_XNOR2X1_4 INVX1_8/gnd DFFSR_7/S FILL
XFILL_0_NOR2X1_13 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_44_4_0 INVX1_2/gnd DFFSR_51/S FILL
XFILL_8_NAND3X1_101 DFFSR_89/gnd DFFSR_186/S FILL
XINVX1_108 DFFSR_96/Q INVX1_2/gnd INVX1_108/Y DFFSR_51/S INVX1
XFILL_1_DFFSR_131 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_15_DFFSR_3 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_42_DFFSR_162 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_7_OAI21X1_185 BUFX2_36/A DFFSR_8/S FILL
XFILL_46_DFFSR_53 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_12_XOR2X1_13 INVX1_8/gnd DFFSR_7/S FILL
XFILL_35_DFFSR_93 INVX1_2/gnd DFFSR_51/S FILL
XFILL_4_INVX1_105 INVX1_4/gnd DFFSR_51/S FILL
XFILL_32_DFFSR_165 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_22_DFFSR_168 BUFX2_36/A DFFSR_8/S FILL
XAOI22X1_6 BUFX2_14/Y AND2X2_6/B AND2X2_6/A AND2X2_5/B BUFX2_37/A OAI22X1_2/D DFFSR_81/S
+ AOI22X1
XFILL_19_DFFSR_43 INVX1_94/gnd DFFSR_25/S FILL
XFILL_2_DFFSR_50 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_4_AOI22X1_3 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_12_DFFSR_171 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_8_OAI21X1_119 BUFX2_37/A DFFSR_8/S FILL
XFILL_2_INVX1_322 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_2_DFFPOSX1_16 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_8_DFFSR_165 BUFX2_6/gnd DFFSR_14/S FILL
XAND2X2_12 NOR2X1_8/A NOR2X1_9/A BUFX2_43/A AND2X2_12/Y DFFSR_97/S AND2X2
XFILL_4_AND2X2_9 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_38_DFFSR_10 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_1_INVX1_142 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_16_DFFSR_90 INVX1_2/gnd DFFSR_1/S FILL
XFILL_27_DFFSR_50 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_6_1 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_7_NAND3X1_131 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_6_OAI21X1_215 BUFX2_43/A DFFSR_97/S FILL
XFILL_0_NAND2X1_112 INVX1_4/gnd DFFSR_4/S FILL
XOAI21X1_251 DFFSR_186/S INVX1_413/Y NAND2X1_262/Y DFFSR_89/gnd DFFSR_183/D DFFSR_92/S
+ OAI21X1
XFILL_12_CLKBUF1_3 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_7_OAI21X1_149 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_21_DFFPOSX1_24 BUFX2_43/A DFFSR_23/S FILL
XFILL_46_DFFSR_17 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_42_DFFSR_126 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_24_DFFSR_97 BUFX2_35/A DFFSR_97/S FILL
XFILL_35_DFFSR_57 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_32_DFFSR_129 INVX1_2/gnd DFFSR_1/S FILL
XFILL_22_DFFSR_132 INVX1_2/gnd DFFSR_51/S FILL
XFILL_2_DFFSR_14 BUFX2_35/A DFFSR_14/S FILL
XFILL_12_DFFSR_135 BUFX2_43/A DFFSR_97/S FILL
XFILL_6_BUFX2_42 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_11_7 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_7_XNOR2X1_2 BUFX2_36/A DFFSR_8/S FILL
XFILL_2_INVX1_286 INVX1_4/gnd DFFSR_51/S FILL
XFILL_18_2_0 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_5_OAI21X1_245 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_8_DFFSR_129 INVX1_2/gnd DFFSR_1/S FILL
XFILL_43_DFFSR_64 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_49_DFFSR_160 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_27_DFFSR_14 BUFX2_35/A DFFSR_14/S FILL
XFILL_16_4_1 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_16_DFFSR_54 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_39_DFFSR_163 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_1_INVX1_106 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_29_DFFSR_166 INVX1_4/gnd DFFSR_51/S FILL
XFILL_15_CLKBUF1_12 BUFX2_43/A DFFSR_23/S FILL
XFILL_19_DFFSR_169 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_6_OAI21X1_179 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_1_AOI22X1_4 INVX1_94/gnd DFFSR_25/S FILL
XNOR2X1_51 NOR2X1_51/A NOR2X1_51/B INVX1_89/gnd NOR2X1_52/B DFFSR_36/S NOR2X1
XFILL_3_DFFSR_2 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_14_CLKBUF1_15 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_13_CLKBUF1_18 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_4_NOR2X1_48 INVX1_89/gnd DFFSR_36/S FILL
XOAI21X1_215 NAND3X1_73/B AOI21X1_22/Y AOI22X1_8/C BUFX2_43/A OAI21X1_223/C DFFSR_97/S
+ OAI21X1
XFILL_3_INVX1_430 INVX1_89/gnd DFFSR_36/S FILL
XFILL_12_CLKBUF1_21 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_11_CLKBUF1_24 INVX1_23/gnd DFFSR_186/S FILL
XFILL_7_OAI21X1_113 INVX1_23/gnd DFFSR_91/S FILL
XFILL_7_DFFSR_68 BUFX2_35/A DFFSR_14/S FILL
XFILL_24_DFFSR_61 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_35_DFFSR_21 INVX1_2/gnd DFFSR_1/S FILL
XFILL_5_DFFSR_166 INVX1_4/gnd DFFSR_51/S FILL
XFILL_1_OR2X2_2 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_1_DFFPOSX1_10 INVX1_8/gnd DFFSR_5/S FILL
XFILL_1_AND2X2_10 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_2_INVX1_250 INVX1_94/gnd DFFSR_25/S FILL
XFILL_27_DFFSR_6 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_6_NAND3X1_125 INVX1_8/gnd DFFSR_5/S FILL
XFILL_32_DFFSR_68 BUFX2_35/A DFFSR_14/S FILL
XFILL_43_DFFSR_28 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_19_CLKBUF1_1 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_4_INVX1_62 INVX1_89/gnd DFFSR_2/S FILL
XFILL_10_DFFPOSX1_29 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_49_DFFSR_124 INVX1_89/gnd DFFSR_36/S FILL
XFILL_5_OAI21X1_209 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_39_DFFSR_127 BUFX2_43/A DFFSR_97/S FILL
XFILL_16_DFFSR_18 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_24_1_2 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_29_DFFSR_130 INVX1_4/gnd DFFSR_51/S FILL
XFILL_20_DFFPOSX1_18 BUFX2_37/A DFFSR_8/S FILL
XFILL_19_DFFSR_133 BUFX2_37/A DFFSR_81/S FILL
XFILL_6_OAI21X1_143 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_6_0_1 BUFX2_35/A DFFSR_14/S FILL
XFILL_48_DFFSR_2 DFFSR_5/gnd DFFSR_2/S FILL
XNOR2X1_15 NOR2X1_15/A NOR2X1_15/B INVX1_4/gnd NOR2X1_15/Y DFFSR_51/S NOR2X1
XFILL_4_XNOR2X1_3 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_40_DFFSR_75 INVX1_4/gnd DFFSR_51/S FILL
XFILL_4_NOR2X1_12 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_4_2_2 BUFX2_6/gnd DFFSR_91/S FILL
XOAI21X1_179 NOR2X1_4/A NOR2X1_3/A NAND2X1_182/Y DFFSR_71/gnd AOI21X1_1/A DFFSR_10/S
+ OAI21X1
XFILL_3_INVX1_394 INVX1_89/gnd DFFSR_2/S FILL
XFILL_33_7 INVX1_8/gnd DFFSR_5/S FILL
XFILL_6_NAND2X1_257 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_7_DFFSR_32 INVX1_2/gnd DFFSR_1/S FILL
XFILL_24_DFFSR_25 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_5_DFFSR_130 INVX1_4/gnd DFFSR_51/S FILL
XFILL_13_DFFSR_65 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_46_DFFSR_161 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_36_DFFSR_164 INVX1_89/gnd DFFSR_2/S FILL
XFILL_4_OAI21X1_239 INVX1_4/gnd DFFSR_4/S FILL
XFILL_3_INVX1_4 INVX1_4/gnd DFFSR_4/S FILL
XFILL_2_INVX1_214 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_0_XOR2X1_2 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_26_DFFSR_167 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_48_DFFSR_82 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_8_AOI22X1_2 BUFX2_37/A DFFSR_81/S FILL
XFILL_16_DFFSR_170 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_5_OAI21X1_173 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_4_INVX1_26 BUFX2_43/A DFFSR_23/S FILL
XFILL_4_DFFSR_79 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_1_NOR2X1_49 INVX1_89/gnd DFFSR_36/S FILL
XFILL_21_DFFSR_72 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_32_DFFSR_32 INVX1_2/gnd DFFSR_1/S FILL
XFILL_0_INVX1_431 INVX1_89/gnd DFFSR_36/S FILL
XNAND3X1_125 INVX1_397/A INVX1_331/A INVX1_332/A INVX1_8/gnd OAI22X1_40/B DFFSR_5/S
+ NAND3X1
XFILL_2_DFFSR_167 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_3_CLKBUF1_12 BUFX2_43/A DFFSR_23/S FILL
XFILL_8_XOR2X1_9 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_3_BUFX2_17 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_6_OAI21X1_107 BUFX2_36/A DFFSR_6/S FILL
XFILL_2_CLKBUF1_15 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_1_CLKBUF1_18 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_1_INVX1_73 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_40_DFFSR_39 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_29_DFFSR_79 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_0_CLKBUF1_21 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_6_NAND2X1_221 BUFX2_6/gnd DFFSR_14/S FILL
XOAI21X1_143 DFFSR_25/S INVX1_161/Y NAND2X1_143/Y BUFX2_8/gnd DFFSR_143/D DFFSR_10/S
+ OAI21X1
XFILL_3_INVX1_358 INVX1_89/gnd DFFSR_36/S FILL
XFILL_16_CLKBUF1_2 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_13_DFFSR_29 INVX1_4/gnd DFFSR_4/S FILL
XFILL_46_DFFSR_125 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_5_NAND3X1_119 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_36_DFFSR_128 BUFX2_19/gnd DFFSR_52/S FILL
XNAND2X1_257 DFFSR_9/S din[2] DFFSR_9/gnd NAND2X1_257/Y DFFSR_9/S NAND2X1
XFILL_4_OAI21X1_203 BUFX2_35/A DFFSR_14/S FILL
XFILL_26_DFFSR_131 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_2_INVX1_178 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_48_DFFSR_46 BUFX2_36/A DFFSR_6/S FILL
XFILL_16_DFFSR_134 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_37_DFFSR_86 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_10_DFFSR_76 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_4_DFFSR_43 INVX1_94/gnd DFFSR_25/S FILL
XFILL_21_DFFSR_36 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_19_DFFPOSX1_12 INVX1_8/gnd DFFSR_5/S FILL
XFILL_1_XNOR2X1_4 INVX1_8/gnd DFFSR_7/S FILL
XFILL_5_OAI21X1_137 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_1_NOR2X1_13 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_0_INVX1_395 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_2_DFFSR_131 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_43_DFFSR_162 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_14_XOR2X1_6 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_5_NAND2X1_251 BUFX2_35/A DFFSR_97/S FILL
XFILL_26_DFFPOSX1_3 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_13_XOR2X1_13 INVX1_8/gnd DFFSR_7/S FILL
XFILL_39_DFFSR_9 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_45_DFFSR_93 INVX1_2/gnd DFFSR_51/S FILL
XFILL_33_DFFSR_165 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_25_DFFPOSX1_6 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_23_DFFSR_168 BUFX2_36/A DFFSR_8/S FILL
XFILL_6_AND2X2_2 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_18_DFFSR_83 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_1_INVX1_37 INVX1_94/gnd DFFSR_52/S FILL
XFILL_29_DFFSR_43 INVX1_94/gnd DFFSR_25/S FILL
XFILL_1_DFFSR_90 INVX1_2/gnd DFFSR_1/S FILL
XFILL_9_DFFPOSX1_23 INVX1_23/gnd DFFSR_91/S FILL
XOAI21X1_107 BUFX2_25/Y INVX1_121/Y OAI21X1_107/C BUFX2_36/A DFFSR_107/D DFFSR_6/S
+ OAI21X1
XFILL_3_OAI21X1_233 BUFX2_36/A DFFSR_8/S FILL
XFILL_24_DFFPOSX1_9 BUFX2_37/A DFFSR_8/S FILL
XFILL_5_AOI22X1_3 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_13_DFFSR_171 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_25_2_0 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_6_NAND2X1_185 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_3_INVX1_322 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_0_BUFX2_28 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_9_DFFSR_165 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_23_4_1 BUFX2_8/gnd DFFSR_10/S FILL
XNAND2X1_221 NAND3X1_70/A NAND3X1_70/Y BUFX2_6/gnd INVX1_260/A DFFSR_14/S NAND2X1
XFILL_5_3_0 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_4_OAI21X1_167 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_9_DFFSR_97 BUFX2_35/A DFFSR_97/S FILL
XFILL_48_DFFSR_10 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_2_INVX1_142 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_37_DFFSR_50 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_3_5_1 INVX1_23/gnd DFFSR_91/S FILL
XFILL_26_DFFSR_90 INVX1_2/gnd DFFSR_1/S FILL
XFILL_4_NAND2X1_281 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_10_DFFSR_40 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_5_OAI21X1_101 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_0_INVX1_359 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_13_CLKBUF1_3 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_2_OAI21X1_263 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_43_DFFSR_126 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_34_DFFSR_97 BUFX2_35/A DFFSR_97/S FILL
XFILL_5_NAND2X1_215 BUFX2_43/A DFFSR_23/S FILL
XFILL_45_DFFSR_57 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_33_DFFSR_129 INVX1_2/gnd DFFSR_1/S FILL
XFILL_4_NAND3X1_113 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_23_DFFSR_132 INVX1_2/gnd DFFSR_51/S FILL
XFILL_13_DFFSR_135 BUFX2_43/A DFFSR_97/S FILL
XFILL_1_DFFSR_54 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_18_DFFSR_47 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_6_NAND2X1_149 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_8_XNOR2X1_2 BUFX2_36/A DFFSR_8/S FILL
XFILL_3_OAI21X1_197 INVX1_8/gnd DFFSR_7/S FILL
XFILL_3_INVX1_286 INVX1_4/gnd DFFSR_51/S FILL
XNAND2X1_185 AND2X2_8/A INVX1_256/A BUFX2_19/gnd NAND3X1_8/A DFFSR_52/S NAND2X1
XFILL_31_1_2 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_9_DFFSR_129 INVX1_2/gnd DFFSR_1/S FILL
XFILL_26_DFFSR_3 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_50_DFFSR_160 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_4_OAI21X1_131 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_37_DFFSR_14 BUFX2_35/A DFFSR_14/S FILL
XFILL_9_DFFSR_61 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_26_DFFSR_54 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_40_DFFSR_163 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_15_DFFSR_94 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_2_INVX1_106 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_10_XOR2X1_14 INVX1_89/gnd DFFSR_2/S FILL
XFILL_30_DFFSR_166 INVX1_4/gnd DFFSR_51/S FILL
XFILL_20_DFFSR_169 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_4_NAND2X1_245 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_10_DFFSR_172 BUFX2_37/A DFFSR_8/S FILL
XFILL_2_AOI22X1_4 INVX1_94/gnd DFFSR_25/S FILL
XINVX1_433 DFFSR_143/Q DFFSR_79/gnd NOR2X1_53/B DFFSR_45/S INVX1
XFILL_5_NOR2X1_48 INVX1_89/gnd DFFSR_36/S FILL
XFILL_0_INVX1_323 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_14_DFFPOSX1_3 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_4_INVX1_430 INVX1_89/gnd DFFSR_36/S FILL
XFILL_2_OAI21X1_227 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_34_DFFSR_61 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_8_DFFPOSX1_17 BUFX2_37/A DFFSR_8/S FILL
XFILL_5_NAND2X1_179 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_45_DFFSR_21 INVX1_2/gnd DFFSR_1/S FILL
XFILL_6_DFFSR_166 INVX1_4/gnd DFFSR_51/S FILL
XFILL_13_DFFPOSX1_6 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_12_DFFPOSX1_9 BUFX2_37/A DFFSR_8/S FILL
XFILL_1_DFFSR_18 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_18_DFFSR_11 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_3_OAI21X1_161 INVX1_23/gnd DFFSR_186/S FILL
XFILL_2_AND2X2_10 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_6_NAND2X1_113 INVX1_23/gnd DFFSR_91/S FILL
XFILL_2_INVX1_1 BUFX2_37/A DFFSR_81/S FILL
XFILL_3_INVX1_250 INVX1_94/gnd DFFSR_25/S FILL
XFILL_42_DFFSR_68 BUFX2_35/A DFFSR_14/S FILL
XFILL_20_CLKBUF1_1 BUFX2_8/gnd DFFSR_25/S FILL
XNAND2X1_149 DFFSR_148/Q DFFSR_91/S DFFSR_89/gnd OAI21X1_149/C DFFSR_186/S NAND2X1
XFILL_8_AOI21X1_41 BUFX2_35/A DFFSR_14/S FILL
XFILL_10_CLKBUF1_4 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_50_DFFSR_124 INVX1_89/gnd DFFSR_36/S FILL
XFILL_3_NAND2X1_275 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_40_DFFSR_127 BUFX2_43/A DFFSR_97/S FILL
XFILL_27_DFFPOSX1_25 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_9_DFFSR_25 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_7_AOI21X1_44 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_26_DFFSR_18 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_30_DFFSR_130 INVX1_4/gnd DFFSR_51/S FILL
XFILL_15_DFFSR_58 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_6_AOI21X1_47 BUFX2_43/A DFFSR_23/S FILL
XFILL_20_DFFSR_133 BUFX2_37/A DFFSR_81/S FILL
XFILL_1_OAI21X1_257 INVX1_2/gnd DFFSR_51/S FILL
XAOI21X1_47 NOR2X1_1/B NOR2X1_1/A AOI21X1_47/C BUFX2_43/A AOI21X1_47/Y DFFSR_23/S
+ AOI21X1
XFILL_4_NAND2X1_209 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_10_DFFSR_136 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_5_XNOR2X1_3 BUFX2_6/gnd DFFSR_91/S FILL
XINVX1_397 INVX1_397/A INVX1_89/gnd INVX1_397/Y DFFSR_36/S INVX1
XFILL_50_DFFSR_75 INVX1_4/gnd DFFSR_51/S FILL
XFILL_0_INVX1_287 INVX1_4/gnd DFFSR_51/S FILL
XFILL_3_NAND3X1_107 BUFX2_43/A DFFSR_97/S FILL
XFILL_20_9 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_5_NOR2X1_12 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_2_OAI21X1_191 BUFX2_37/A DFFSR_8/S FILL
XFILL_5_NAND2X1_143 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_4_INVX1_394 INVX1_89/gnd DFFSR_2/S FILL
XFILL_34_DFFSR_25 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_6_DFFSR_72 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_6_DFFSR_130 INVX1_4/gnd DFFSR_51/S FILL
XFILL_23_DFFSR_65 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_47_DFFSR_161 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_5_BUFX2_10 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_37_DFFSR_164 INVX1_89/gnd DFFSR_2/S FILL
XFILL_3_OAI21X1_125 BUFX2_35/A DFFSR_14/S FILL
XFILL_3_INVX1_214 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_27_DFFSR_167 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_9_OAI21X1_86 INVX1_4/gnd DFFSR_51/S FILL
XFILL_8_OAI21X1_89 BUFX2_35/A DFFSR_14/S FILL
XFILL_9_AOI22X1_2 BUFX2_37/A DFFSR_81/S FILL
XFILL_17_DFFSR_170 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_7_OAI21X1_92 BUFX2_5/gnd DFFSR_23/S FILL
XNAND2X1_113 DFFSR_105/Q BUFX2_21/Y INVX1_23/gnd NAND2X1_113/Y DFFSR_91/S NAND2X1
XFILL_3_NAND2X1_239 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_2_NOR2X1_49 INVX1_89/gnd DFFSR_36/S FILL
XFILL_6_OAI21X1_95 INVX1_89/gnd DFFSR_36/S FILL
XFILL_31_DFFSR_72 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_42_DFFSR_32 INVX1_2/gnd DFFSR_1/S FILL
XFILL_3_INVX1_66 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_5_OAI21X1_98 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_15_DFFSR_22 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_3_DFFSR_167 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_1_INVX1_431 INVX1_89/gnd DFFSR_36/S FILL
XOAI21X1_95 BUFX2_22/Y INVX1_107/Y NAND2X1_95/Y INVX1_89/gnd DFFSR_95/D DFFSR_36/S
+ OAI21X1
XFILL_6_AOI21X1_11 INVX1_8/gnd DFFSR_5/S FILL
XFILL_1_OAI21X1_221 BUFX2_35/A DFFSR_14/S FILL
XFILL_4_NAND2X1_173 BUFX2_35/A DFFSR_14/S FILL
XFILL_5_AOI21X1_14 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_32_2_0 INVX1_8/gnd DFFSR_5/S FILL
XFILL_7_DFFPOSX1_11 INVX1_4/gnd DFFSR_4/S FILL
XFILL_10_DFFSR_100 INVX1_23/gnd DFFSR_186/S FILL
XFILL_38_DFFSR_6 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_4_AOI21X1_17 INVX1_8/gnd DFFSR_5/S FILL
XAOI21X1_11 INVX1_228/Y NOR3X1_1/A INVX1_229/A INVX1_8/gnd AOI21X1_11/Y DFFSR_5/S
+ AOI21X1
XFILL_0_INVX1_251 BUFX2_36/A DFFSR_8/S FILL
XFILL_3_AOI21X1_20 BUFX2_7/gnd DFFSR_81/S FILL
XINVX1_361 DFFSR_92/Q BUFX2_7/gnd INVX1_361/Y DFFSR_81/S INVX1
XFILL_2_DFFPOSX1_3 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_50_DFFSR_39 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_39_DFFSR_79 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_30_4_1 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_16_DFFPOSX1_30 BUFX2_43/A DFFSR_97/S FILL
XFILL_2_AOI21X1_23 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_4_INVX1_358 INVX1_89/gnd DFFSR_36/S FILL
XFILL_1_DFFPOSX1_6 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_12_DFFSR_69 BUFX2_43/A DFFSR_23/S FILL
XFILL_1_AOI21X1_26 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_5_NAND2X1_107 BUFX2_36/A DFFSR_6/S FILL
XFILL_0_DFFPOSX1_9 BUFX2_37/A DFFSR_8/S FILL
XFILL_2_OAI21X1_155 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_17_CLKBUF1_2 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_6_DFFSR_36 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_23_DFFSR_29 INVX1_4/gnd DFFSR_4/S FILL
XFILL_47_DFFSR_125 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_0_AOI21X1_29 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_37_DFFSR_128 BUFX2_19/gnd DFFSR_52/S FILL
XBUFX2_14 BUFX2_14/A BUFX2_37/A BUFX2_14/Y DFFSR_81/S BUFX2
XFILL_27_DFFSR_131 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_2_NAND2X1_269 INVX1_4/gnd DFFSR_4/S FILL
XFILL_3_INVX1_178 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_17_DFFSR_134 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_9_OAI21X1_50 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_47_DFFSR_86 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_26_DFFPOSX1_19 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_8_OAI21X1_53 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_0_OAI21X1_251 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_20_DFFSR_76 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_3_DFFSR_83 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_31_DFFSR_36 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_2_XNOR2X1_4 INVX1_8/gnd DFFSR_7/S FILL
XFILL_6_NAND2X1_74 INVX1_2/gnd DFFSR_1/S FILL
XFILL_3_INVX1_30 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_7_OAI21X1_56 INVX1_2/gnd DFFSR_51/S FILL
XFILL_3_NAND2X1_203 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_5_NAND2X1_77 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_2_NOR2X1_13 BUFX2_17/gnd DFFSR_57/S FILL
XNAND2X1_74 BUFX2_18/Y INVX1_75/A INVX1_2/gnd NAND2X1_74/Y DFFSR_1/S NAND2X1
XFILL_6_OAI21X1_59 INVX1_4/gnd DFFSR_51/S FILL
XFILL_5_OAI21X1_62 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_1_INVX1_395 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_4_NAND2X1_80 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_2_NAND3X1_101 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_2_BUFX2_21 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_3_NAND2X1_83 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_3_DFFSR_131 DFFSR_1/gnd DFFSR_1/S FILL
XOAI21X1_59 DFFSR_51/S INVX1_67/Y OAI21X1_59/C INVX1_4/gnd DFFSR_59/D DFFSR_51/S OAI21X1
XFILL_4_OAI21X1_65 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_44_DFFSR_162 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_10_AOI22X1_9 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_1_OAI21X1_185 BUFX2_36/A DFFSR_8/S FILL
XFILL_3_OAI21X1_68 BUFX2_37/A DFFSR_81/S FILL
XFILL_2_NAND2X1_86 INVX1_4/gnd DFFSR_51/S FILL
XFILL_34_DFFSR_165 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_1_NAND2X1_89 BUFX2_37/A DFFSR_8/S FILL
XFILL_4_NAND2X1_137 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_2_OAI21X1_71 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_14_XOR2X1_13 INVX1_8/gnd DFFSR_7/S FILL
XFILL_0_INVX1_215 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_0_NAND2X1_92 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_24_DFFSR_168 BUFX2_36/A DFFSR_8/S FILL
XFILL_0_INVX1_77 BUFX2_37/A DFFSR_81/S FILL
XFILL_28_DFFSR_83 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_39_DFFSR_43 INVX1_94/gnd DFFSR_25/S FILL
XINVX1_325 DFFSR_40/Q BUFX2_17/gnd INVX1_325/Y DFFSR_7/S INVX1
XFILL_1_OAI21X1_74 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_6_AOI22X1_3 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_14_DFFSR_171 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_0_OAI21X1_77 INVX1_89/gnd DFFSR_36/S FILL
XFILL_38_1_2 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_2_OAI21X1_119 BUFX2_37/A DFFSR_8/S FILL
XFILL_4_INVX1_322 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_12_DFFSR_33 INVX1_94/gnd DFFSR_52/S FILL
XFILL_0_XOR2X1_10 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_0_DFFSR_168 BUFX2_36/A DFFSR_8/S FILL
XFILL_5_DFFSR_9 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_9_OAI21X1_14 BUFX2_43/A DFFSR_23/S FILL
XFILL_2_NAND2X1_233 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_3_INVX1_142 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_47_DFFSR_50 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_1_NAND3X1_131 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_8_OAI21X1_17 INVX1_8/gnd DFFSR_5/S FILL
XFILL_36_DFFSR_90 INVX1_2/gnd DFFSR_1/S FILL
XFILL_7_OAI21X1_20 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_6_NAND2X1_38 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_0_OAI21X1_215 BUFX2_43/A DFFSR_97/S FILL
XFILL_6_OAI21X1_23 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_3_DFFSR_47 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_20_DFFSR_40 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_5_NAND2X1_41 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_3_NAND2X1_167 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_4_NAND2X1_44 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_1_INVX1_359 DFFSR_79/gnd DFFSR_36/S FILL
XNAND2X1_38 DFFSR_5/S DFFSR_30/Q DFFSR_5/gnd OAI21X1_38/C DFFSR_5/S NAND2X1
XFILL_5_OAI21X1_26 DFFSR_1/gnd DFFSR_9/S FILL
XOAI21X1_23 DFFSR_158/S INVX1_26/Y OAI21X1_23/C BUFX2_5/gnd DFFSR_23/D DFFSR_23/S
+ OAI21X1
XFILL_3_NAND2X1_47 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_14_CLKBUF1_3 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_4_OAI21X1_29 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_2_NAND2X1_50 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_44_DFFSR_126 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_1_OAI21X1_149 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_44_DFFSR_97 BUFX2_35/A DFFSR_97/S FILL
XFILL_15_DFFPOSX1_24 BUFX2_43/A DFFSR_23/S FILL
XFILL_4_NAND2X1_101 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_34_DFFSR_129 INVX1_2/gnd DFFSR_1/S FILL
XFILL_3_OAI21X1_32 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_5_AND2X2_6 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_1_NAND2X1_53 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_2_OAI21X1_35 INVX1_8/gnd DFFSR_5/S FILL
XFILL_24_DFFSR_132 INVX1_2/gnd DFFSR_51/S FILL
XFILL_14_DFFSR_135 BUFX2_43/A DFFSR_97/S FILL
XFILL_0_INVX1_179 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_19_1 BUFX2_19/gnd DFFSR_54/S FILL
XINVX1_289 DFFSR_20/Q BUFX2_19/gnd INVX1_289/Y DFFSR_52/S INVX1
XFILL_0_INVX1_41 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_28_DFFSR_47 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_1_OAI21X1_38 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_0_NAND2X1_56 INVX1_4/gnd DFFSR_51/S FILL
XFILL_17_DFFSR_87 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_0_DFFSR_94 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_9_XNOR2X1_2 BUFX2_36/A DFFSR_8/S FILL
XFILL_0_OAI21X1_41 INVX1_8/gnd DFFSR_7/S FILL
XFILL_1_NAND2X1_263 INVX1_2/gnd DFFSR_51/S FILL
XFILL_4_INVX1_286 INVX1_4/gnd DFFSR_51/S FILL
XFILL_25_DFFPOSX1_13 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_8_AOI22X1_10 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_7_AOI22X1_13 INVX1_23/gnd DFFSR_186/S FILL
XFILL_50_DFFSR_9 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_2_NAND2X1_197 INVX1_8/gnd DFFSR_5/S FILL
XFILL_0_DFFSR_132 INVX1_2/gnd DFFSR_51/S FILL
XFILL_47_DFFSR_14 BUFX2_35/A DFFSR_14/S FILL
XFILL_36_DFFSR_54 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_41_DFFSR_163 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_25_DFFSR_94 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_3_INVX1_106 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_11_XOR2X1_14 INVX1_89/gnd DFFSR_2/S FILL
XFILL_31_DFFSR_166 INVX1_4/gnd DFFSR_51/S FILL
XFILL_21_DFFSR_169 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_0_OAI21X1_179 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_3_DFFSR_11 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_9_OAI21X1_234 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_11_DFFSR_172 BUFX2_37/A DFFSR_8/S FILL
XFILL_3_AOI22X1_4 INVX1_94/gnd DFFSR_25/S FILL
XFILL_3_NAND2X1_131 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_6_NOR2X1_48 INVX1_89/gnd DFFSR_36/S FILL
XFILL_1_INVX1_323 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_11_OAI22X1_49 INVX1_94/gnd DFFSR_25/S FILL
XFILL_3_NAND2X1_11 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_1_OAI21X1_113 INVX1_23/gnd DFFSR_91/S FILL
XFILL_2_NAND2X1_14 BUFX2_43/A DFFSR_23/S FILL
XFILL_44_DFFSR_61 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_10_OAI22X1_52 INVX1_94/gnd DFFSR_25/S FILL
XFILL_7_DFFSR_166 INVX1_4/gnd DFFSR_51/S FILL
XFILL_1_NAND2X1_17 INVX1_8/gnd DFFSR_7/S FILL
XFILL_0_NAND2X1_20 INVX1_23/gnd DFFSR_186/S FILL
XINVX1_253 INVX1_253/A BUFX2_35/A XOR2X1_8/B DFFSR_97/S INVX1
XFILL_8_NAND3X1_73 BUFX2_43/A DFFSR_23/S FILL
XFILL_0_INVX1_143 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_9_OAI22X1_55 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_0_DFFSR_58 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_28_DFFSR_11 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_3_AND2X2_10 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_7_NAND3X1_76 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_8_OAI22X1_58 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_17_DFFSR_51 INVX1_2/gnd DFFSR_51/S FILL
XFILL_1_NAND2X1_227 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_6_NAND3X1_79 BUFX2_36/A DFFSR_6/S FILL
XFILL_4_INVX1_250 INVX1_94/gnd DFFSR_25/S FILL
XFILL_7_OAI22X1_61 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_5_NAND3X1_82 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_6_OAI22X1_64 INVX1_94/gnd DFFSR_25/S FILL
XNAND3X1_79 NAND3X1_74/Y NAND3X1_75/Y NAND3X1_72/C BUFX2_36/A NAND3X1_79/Y DFFSR_6/S
+ NAND3X1
XFILL_4_NAND3X1_85 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_0_NAND3X1_125 INVX1_8/gnd DFFSR_5/S FILL
XFILL_16_DFFSR_7 INVX1_8/gnd DFFSR_7/S FILL
XFILL_5_OAI22X1_67 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_3_NAND3X1_88 INVX1_94/gnd DFFSR_52/S FILL
XOAI22X1_64 INVX1_386/Y OAI22X1_40/B INVX1_387/Y OAI22X1_40/D INVX1_94/gnd NOR2X1_41/A
+ DFFSR_25/S OAI22X1
XFILL_11_CLKBUF1_4 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_39_2_0 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_2_NAND2X1_161 INVX1_23/gnd DFFSR_186/S FILL
XFILL_2_NAND3X1_91 BUFX2_43/A DFFSR_97/S FILL
XFILL_41_DFFSR_127 BUFX2_43/A DFFSR_97/S FILL
XFILL_8_OAI21X1_264 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_8_DFFSR_65 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_1_NAND3X1_94 BUFX2_35/A DFFSR_97/S FILL
XFILL_14_DFFSR_98 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_36_DFFSR_18 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_31_DFFSR_130 INVX1_4/gnd DFFSR_51/S FILL
XFILL_25_DFFSR_58 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_37_4_1 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_0_NAND3X1_97 BUFX2_35/A DFFSR_97/S FILL
XFILL_21_DFFSR_133 BUFX2_37/A DFFSR_81/S FILL
XFILL_0_BUFX2_8 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_14_DFFPOSX1_18 BUFX2_37/A DFFSR_8/S FILL
XFILL_0_OAI21X1_143 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_11_DFFSR_136 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_6_XNOR2X1_3 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_1_INVX1_287 INVX1_4/gnd DFFSR_51/S FILL
XFILL_37_DFFSR_3 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_11_OAI22X1_13 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_41_1 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_6_NOR2X1_12 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_0_NAND2X1_257 DFFSR_9/gnd DFFSR_9/S FILL
XINVX1_99 DFFSR_88/Q INVX1_4/gnd INVX1_99/Y DFFSR_4/S INVX1
XFILL_10_OAI22X1_16 INVX1_4/gnd DFFSR_4/S FILL
XFILL_44_DFFSR_25 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_7_DFFSR_130 INVX1_4/gnd DFFSR_51/S FILL
XFILL_33_DFFSR_65 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_48_DFFSR_161 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_8_NAND3X1_37 BUFX2_43/A DFFSR_97/S FILL
XFILL_9_OAI22X1_19 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_7_NAND3X1_40 BUFX2_43/A DFFSR_23/S FILL
XINVX1_217 NAND3X1_1/Y INVX1_94/gnd OR2X2_1/B DFFSR_25/S INVX1
XFILL_0_DFFSR_22 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_0_INVX1_107 INVX1_89/gnd DFFSR_36/S FILL
XFILL_38_DFFSR_164 INVX1_89/gnd DFFSR_2/S FILL
XFILL_17_DFFSR_15 INVX1_8/gnd DFFSR_7/S FILL
XFILL_8_OAI22X1_22 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_1_NAND2X1_191 BUFX2_37/A DFFSR_8/S FILL
XFILL_28_DFFSR_167 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_4_DFFPOSX1_29 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_6_NAND3X1_43 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_18_DFFSR_170 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_7_OAI22X1_25 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_5_NAND3X1_46 BUFX2_35/A DFFSR_97/S FILL
XNAND3X1_43 INVX1_241/Y NAND3X1_40/B NAND3X1_40/C BUFX2_5/gnd NAND3X1_48/B DFFSR_23/S
+ NAND3X1
XFILL_0_AOI22X1_5 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_6_OAI22X1_28 INVX1_94/gnd DFFSR_25/S FILL
XXOR2X1_12 XOR2X1_12/A XOR2X1_12/B BUFX2_17/gnd XOR2X1_12/Y DFFSR_7/S XOR2X1
XFILL_4_NAND3X1_49 BUFX2_37/A DFFSR_8/S FILL
XOAI22X1_28 INVX1_311/Y OAI22X1_8/B INVX1_312/Y OAI22X1_9/D INVX1_94/gnd NOR2X1_23/B
+ DFFSR_25/S OAI22X1
XFILL_5_OAI22X1_31 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_3_NOR2X1_49 INVX1_89/gnd DFFSR_36/S FILL
XFILL_41_DFFSR_72 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_2_NAND2X1_125 BUFX2_35/A DFFSR_14/S FILL
XFILL_3_NAND3X1_52 BUFX2_36/A DFFSR_8/S FILL
XDFFSR_170 INVX1_256/A CLKBUF1_16/Y DFFSR_175/R DFFSR_81/S DFFSR_170/D BUFX2_7/gnd
+ DFFSR_81/S DFFSR
XFILL_8_OAI21X1_228 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_4_OAI22X1_34 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_2_NAND3X1_55 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_14_DFFSR_62 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_25_DFFSR_22 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_3_OAI22X1_37 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_4_DFFSR_167 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_2_INVX1_431 INVX1_89/gnd DFFSR_36/S FILL
XFILL_8_DFFSR_29 INVX1_4/gnd DFFSR_4/S FILL
XFILL_2_OAI22X1_40 BUFX2_37/A DFFSR_8/S FILL
XFILL_1_NAND3X1_58 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_45_1_2 INVX1_2/gnd DFFSR_1/S FILL
XFILL_0_OAI21X1_107 BUFX2_36/A DFFSR_6/S FILL
XFILL_1_OAI22X1_43 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_0_NAND3X1_61 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_11_DFFSR_100 INVX1_23/gnd DFFSR_186/S FILL
XFILL_0_AND2X2_11 BUFX2_35/A DFFSR_14/S FILL
XFILL_0_OAI22X1_46 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_1_INVX1_251 BUFX2_36/A DFFSR_8/S FILL
XFILL_49_DFFSR_79 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_0_NAND2X1_221 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_22_DFFSR_69 BUFX2_43/A DFFSR_23/S FILL
XFILL_5_DFFSR_76 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_18_CLKBUF1_2 DFFSR_79/gnd DFFSR_45/S FILL
XINVX1_63 DFFSR_56/Q INVX1_2/gnd INVX1_63/Y DFFSR_51/S INVX1
XFILL_33_DFFSR_29 INVX1_4/gnd DFFSR_4/S FILL
XFILL_48_DFFSR_125 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_13_0_0 BUFX2_36/A DFFSR_8/S FILL
XINVX1_181 BUFX2_9/Y BUFX2_37/A DFFSR_153/R DFFSR_8/S INVX1
XFILL_38_DFFSR_128 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_9_XOR2X1_6 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_4_BUFX2_14 BUFX2_37/A DFFSR_81/S FILL
XCLKBUF1_2 DFFSR_149/Q DFFSR_79/gnd CLKBUF1_2/Y DFFSR_45/S CLKBUF1
XFILL_28_DFFSR_131 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_11_2_1 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_4_DFFSR_6 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_4_INVX1_178 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_1_NAND2X1_155 BUFX2_37/A DFFSR_81/S FILL
XFILL_18_DFFSR_134 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_7_OAI21X1_258 INVX1_2/gnd DFFSR_51/S FILL
XFILL_5_NAND3X1_10 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_30_DFFSR_76 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_2_INVX1_70 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_4_NAND3X1_13 INVX1_94/gnd DFFSR_25/S FILL
XFILL_41_DFFSR_36 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_3_XNOR2X1_4 INVX1_8/gnd DFFSR_7/S FILL
XFILL_3_NAND3X1_16 BUFX2_19/gnd DFFSR_52/S FILL
XDFFSR_134 DFFSR_134/Q CLKBUF1_9/Y DFFSR_135/R DFFSR_45/S DFFSR_134/D DFFSR_79/gnd
+ DFFSR_45/S DFFSR
XFILL_13_DFFPOSX1_12 INVX1_8/gnd DFFSR_5/S FILL
XFILL_3_NOR2X1_13 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_8_OAI21X1_192 BUFX2_37/A DFFSR_81/S FILL
XFILL_2_INVX1_395 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_2_NAND3X1_19 INVX1_8/gnd DFFSR_5/S FILL
XFILL_1_NAND3X1_22 BUFX2_37/A DFFSR_81/S FILL
XFILL_4_DFFSR_131 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_14_DFFSR_26 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_45_DFFSR_162 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_11_AOI22X1_9 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_0_NAND3X1_25 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_35_DFFSR_165 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_15_XOR2X1_13 INVX1_8/gnd DFFSR_7/S FILL
XFILL_1_INVX1_215 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_25_DFFSR_168 BUFX2_36/A DFFSR_8/S FILL
XFILL_49_DFFSR_43 INVX1_94/gnd DFFSR_25/S FILL
XFILL_0_OAI22X1_10 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_7_AOI22X1_3 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_38_DFFSR_83 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_15_DFFSR_171 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_3_DFFPOSX1_23 INVX1_23/gnd DFFSR_91/S FILL
XFILL_0_NAND2X1_185 BUFX2_19/gnd DFFSR_52/S FILL
XDFFSR_80 INVX1_90/A CLKBUF1_3/Y DFFSR_76/R DFFSR_65/S DFFSR_80/D BUFX2_16/gnd DFFSR_65/S
+ DFFSR
XINVX1_27 INVX1_27/A DFFSR_73/gnd INVX1_27/Y DFFSR_11/S INVX1
XFILL_22_DFFSR_33 INVX1_94/gnd DFFSR_52/S FILL
XFILL_0_NOR2X1_50 INVX1_89/gnd DFFSR_36/S FILL
XFILL_5_DFFSR_40 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_1_XOR2X1_10 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_11_DFFSR_73 DFFSR_73/gnd DFFSR_11/S FILL
XINVX1_145 BUFX2_5/Y BUFX2_43/A DFFSR_123/R DFFSR_97/S INVX1
XFILL_1_DFFSR_168 BUFX2_36/A DFFSR_8/S FILL
XFILL_7_OAI21X1_222 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_49_DFFSR_6 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_1_NAND2X1_119 BUFX2_37/A DFFSR_8/S FILL
XFILL_15_XOR2X1_3 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_4_INVX1_142 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_46_DFFSR_90 INVX1_2/gnd DFFSR_1/S FILL
XFILL_2_INVX1_34 INVX1_89/gnd DFFSR_36/S FILL
XFILL_30_DFFSR_40 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_2_DFFSR_87 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_19_DFFSR_80 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_8_OAI21X1_156 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_22_DFFPOSX1_31 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_15_CLKBUF1_3 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_2_INVX1_359 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_1_BUFX2_25 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_4_INVX1_8 INVX1_8/gnd DFFSR_5/S FILL
XFILL_45_DFFSR_126 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_35_DFFSR_129 INVX1_2/gnd DFFSR_1/S FILL
XFILL_25_DFFSR_132 INVX1_2/gnd DFFSR_51/S FILL
XFILL_15_DFFSR_135 BUFX2_43/A DFFSR_97/S FILL
XFILL_1_INVX1_179 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_38_DFFSR_47 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_27_DFFSR_87 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_46_2_0 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_0_NAND2X1_149 DFFSR_89/gnd DFFSR_186/S FILL
XDFFSR_44 INVX1_50/A DFFSR_52/CLK DFFSR_46/R DFFSR_44/S DFFSR_44/D BUFX2_8/gnd DFFSR_10/S
+ DFFSR
XFILL_11_DFFSR_37 INVX1_89/gnd DFFSR_2/S FILL
XFILL_6_OAI21X1_252 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_44_4_1 INVX1_2/gnd DFFSR_51/S FILL
XFILL_0_NOR2X1_14 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_8_NAND3X1_102 INVX1_23/gnd DFFSR_186/S FILL
XINVX1_109 BUFX2_5/Y BUFX2_35/A DFFSR_89/R DFFSR_97/S INVX1
XFILL_1_DFFSR_132 INVX1_2/gnd DFFSR_51/S FILL
XFILL_15_DFFSR_4 INVX1_4/gnd DFFSR_4/S FILL
XFILL_7_OAI21X1_186 BUFX2_36/A DFFSR_8/S FILL
XFILL_46_DFFSR_54 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_42_DFFSR_163 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_35_DFFSR_94 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_4_INVX1_106 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_12_XOR2X1_14 INVX1_89/gnd DFFSR_2/S FILL
XFILL_32_DFFSR_166 INVX1_4/gnd DFFSR_51/S FILL
XAOI22X1_7 AOI22X1_7/A AOI22X1_7/B AOI22X1_7/C AOI22X1_7/D BUFX2_43/A AOI22X1_7/Y
+ DFFSR_23/S AOI22X1
XFILL_22_DFFSR_169 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_19_DFFSR_44 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_2_DFFSR_51 INVX1_2/gnd DFFSR_51/S FILL
XFILL_12_DFFSR_172 BUFX2_37/A DFFSR_8/S FILL
XFILL_4_AOI22X1_4 INVX1_94/gnd DFFSR_25/S FILL
XFILL_8_OAI21X1_120 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_2_INVX1_323 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_10_5_0 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_2_DFFPOSX1_17 BUFX2_37/A DFFSR_8/S FILL
XFILL_8_DFFSR_166 INVX1_4/gnd DFFSR_51/S FILL
XAND2X2_13 AND2X2_13/A AND2X2_13/B BUFX2_19/gnd OAI22X1_4/D DFFSR_54/S AND2X2
XFILL_1_INVX1_143 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_38_DFFSR_11 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_16_DFFSR_91 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_6_2 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_4_AND2X2_10 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_7_NAND3X1_132 INVX1_8/gnd DFFSR_7/S FILL
XFILL_27_DFFSR_51 INVX1_2/gnd DFFSR_51/S FILL
XFILL_0_NAND2X1_113 INVX1_23/gnd DFFSR_91/S FILL
XFILL_6_OAI21X1_216 BUFX2_35/A DFFSR_14/S FILL
XFILL_12_CLKBUF1_4 BUFX2_8/gnd DFFSR_10/S FILL
XOAI21X1_252 DFFSR_1/S INVX1_415/Y NAND2X1_263/Y DFFSR_1/gnd DFFSR_184/D DFFSR_1/S
+ OAI21X1
XFILL_42_DFFSR_127 BUFX2_43/A DFFSR_97/S FILL
XFILL_21_DFFPOSX1_25 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_7_OAI21X1_150 INVX1_94/gnd DFFSR_52/S FILL
XFILL_24_DFFSR_98 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_46_DFFSR_18 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_32_DFFSR_130 INVX1_4/gnd DFFSR_51/S FILL
XFILL_35_DFFSR_58 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_22_DFFSR_133 BUFX2_37/A DFFSR_81/S FILL
XFILL_6_BUFX2_43 BUFX2_35/A DFFSR_97/S FILL
XFILL_12_DFFSR_136 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_2_DFFSR_15 INVX1_8/gnd DFFSR_7/S FILL
XFILL_7_XNOR2X1_3 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_20_0_0 INVX1_94/gnd DFFSR_52/S FILL
XFILL_2_INVX1_287 INVX1_4/gnd DFFSR_51/S FILL
XFILL_18_2_1 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_5_OAI21X1_246 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_8_DFFSR_130 INVX1_4/gnd DFFSR_51/S FILL
XFILL_43_DFFSR_65 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_0_1_0 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_49_DFFSR_161 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_16_4_2 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_16_DFFSR_55 INVX1_89/gnd DFFSR_36/S FILL
XFILL_1_INVX1_107 INVX1_89/gnd DFFSR_36/S FILL
XFILL_39_DFFSR_164 INVX1_89/gnd DFFSR_2/S FILL
XFILL_27_DFFSR_15 INVX1_8/gnd DFFSR_7/S FILL
XFILL_29_DFFSR_167 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_16_CLKBUF1_10 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_19_DFFSR_170 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_6_OAI21X1_180 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_15_CLKBUF1_13 INVX1_4/gnd DFFSR_51/S FILL
XFILL_1_AOI22X1_5 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_14_CLKBUF1_16 BUFX2_36/A DFFSR_6/S FILL
XNOR2X1_52 NOR2X1_52/A NOR2X1_52/B DFFSR_79/gnd NOR2X1_52/Y DFFSR_36/S NOR2X1
XFILL_3_DFFSR_3 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_4_NOR2X1_49 INVX1_89/gnd DFFSR_36/S FILL
XFILL_13_CLKBUF1_19 DFFSR_9/gnd DFFSR_9/S FILL
XOAI21X1_216 INVX1_227/Y INVX1_240/Y XOR2X1_4/A BUFX2_35/A OAI21X1_217/C DFFSR_14/S
+ OAI21X1
XFILL_12_CLKBUF1_22 INVX1_94/gnd DFFSR_25/S FILL
XFILL_11_CLKBUF1_25 INVX1_23/gnd DFFSR_186/S FILL
XFILL_7_DFFSR_69 BUFX2_43/A DFFSR_23/S FILL
XFILL_24_DFFSR_62 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_35_DFFSR_22 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_5_DFFSR_167 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_3_INVX1_431 INVX1_89/gnd DFFSR_36/S FILL
XFILL_7_OAI21X1_114 INVX1_89/gnd DFFSR_36/S FILL
XFILL_1_OR2X2_3 BUFX2_43/A DFFSR_23/S FILL
XFILL_1_DFFPOSX1_11 INVX1_4/gnd DFFSR_4/S FILL
XFILL_12_DFFSR_100 INVX1_23/gnd DFFSR_186/S FILL
XFILL_1_AND2X2_11 BUFX2_35/A DFFSR_14/S FILL
XFILL_2_INVX1_251 BUFX2_36/A DFFSR_8/S FILL
XFILL_6_NAND3X1_126 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_27_DFFSR_7 INVX1_8/gnd DFFSR_7/S FILL
XFILL_10_DFFPOSX1_30 BUFX2_43/A DFFSR_97/S FILL
XFILL_32_DFFSR_69 BUFX2_43/A DFFSR_23/S FILL
XFILL_19_CLKBUF1_2 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_4_INVX1_63 INVX1_2/gnd DFFSR_51/S FILL
XFILL_43_DFFSR_29 INVX1_4/gnd DFFSR_4/S FILL
XFILL_49_DFFSR_125 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_5_OAI21X1_210 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_39_DFFSR_128 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_29_DFFSR_131 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_16_DFFSR_19 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_19_DFFSR_134 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_20_DFFPOSX1_19 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_6_0_2 BUFX2_35/A DFFSR_14/S FILL
XFILL_6_OAI21X1_144 INVX1_8/gnd DFFSR_7/S FILL
XFILL_48_DFFSR_3 DFFSR_3/gnd DFFSR_4/S FILL
XNOR2X1_16 NOR2X1_16/A NOR2X1_16/B DFFSR_3/gnd NOR2X1_16/Y DFFSR_65/S NOR2X1
XFILL_40_DFFSR_76 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_51_DFFSR_36 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_4_XNOR2X1_4 INVX1_8/gnd DFFSR_7/S FILL
XOAI21X1_180 XOR2X1_2/B XOR2X1_2/A NAND3X1_2/B DFFSR_71/gnd INVX1_221/A DFFSR_10/S
+ OAI21X1
XFILL_4_NOR2X1_13 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_3_INVX1_395 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_33_8 INVX1_8/gnd DFFSR_5/S FILL
XFILL_6_NAND2X1_258 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_7_DFFSR_33 INVX1_94/gnd DFFSR_52/S FILL
XFILL_5_DFFSR_131 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_24_DFFSR_26 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_13_DFFSR_66 INVX1_2/gnd DFFSR_51/S FILL
XFILL_46_DFFSR_162 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_36_DFFSR_165 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_4_OAI21X1_240 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_3_INVX1_5 INVX1_4/gnd DFFSR_51/S FILL
XFILL_2_INVX1_215 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_26_DFFSR_168 BUFX2_36/A DFFSR_8/S FILL
XFILL_0_XOR2X1_3 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_8_AOI22X1_3 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_48_DFFSR_83 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_16_DFFSR_171 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_5_OAI21X1_174 BUFX2_43/A DFFSR_23/S FILL
XFILL_32_DFFSR_33 INVX1_94/gnd DFFSR_52/S FILL
XFILL_1_NOR2X1_50 INVX1_89/gnd DFFSR_36/S FILL
XFILL_4_DFFSR_80 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_2_XOR2X1_10 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_21_DFFSR_73 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_4_INVX1_27 DFFSR_73/gnd DFFSR_11/S FILL
XNAND3X1_126 INVX1_397/A INVX1_332/A INVX1_331/Y DFFSR_5/gnd OAI22X1_40/D DFFSR_5/S
+ NAND3X1
XFILL_2_DFFSR_168 BUFX2_36/A DFFSR_8/S FILL
XFILL_0_INVX1_432 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_4_CLKBUF1_10 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_3_CLKBUF1_13 INVX1_4/gnd DFFSR_51/S FILL
XFILL_3_BUFX2_18 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_2_CLKBUF1_16 BUFX2_36/A DFFSR_6/S FILL
XFILL_6_OAI21X1_108 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_14_DFFSR_1 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_17_5_0 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_40_DFFSR_40 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_1_CLKBUF1_19 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_1_INVX1_74 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_29_DFFSR_80 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_0_CLKBUF1_22 INVX1_94/gnd DFFSR_25/S FILL
XOAI21X1_144 DFFSR_5/S INVX1_162/Y NAND2X1_144/Y INVX1_8/gnd DFFSR_144/D DFFSR_7/S
+ OAI21X1
XFILL_6_NAND2X1_222 INVX1_23/gnd DFFSR_186/S FILL
XFILL_16_CLKBUF1_3 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_3_INVX1_359 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_13_DFFSR_30 INVX1_89/gnd DFFSR_36/S FILL
XFILL_5_NAND3X1_120 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_46_DFFSR_126 BUFX2_17/gnd DFFSR_57/S FILL
XNAND2X1_258 DFFSR_9/S din[3] DFFSR_9/gnd OAI21X1_247/C DFFSR_9/S NAND2X1
XFILL_36_DFFSR_129 INVX1_2/gnd DFFSR_1/S FILL
XFILL_4_OAI21X1_204 BUFX2_36/A DFFSR_6/S FILL
XFILL_26_DFFSR_132 INVX1_2/gnd DFFSR_51/S FILL
XFILL_16_DFFSR_135 BUFX2_43/A DFFSR_97/S FILL
XFILL_2_INVX1_179 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_48_DFFSR_47 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_37_DFFSR_87 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_19_DFFPOSX1_13 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_4_DFFSR_44 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_21_DFFSR_37 INVX1_89/gnd DFFSR_2/S FILL
XFILL_10_DFFSR_77 INVX1_89/gnd DFFSR_2/S FILL
XFILL_1_NOR2X1_14 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_5_OAI21X1_138 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_0_INVX1_396 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_27_DFFPOSX1_1 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_2_DFFSR_132 INVX1_2/gnd DFFSR_51/S FILL
XFILL_14_XOR2X1_7 INVX1_23/gnd DFFSR_91/S FILL
XFILL_5_NAND2X1_252 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_43_DFFSR_163 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_45_DFFSR_94 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_27_0_0 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_13_XOR2X1_14 INVX1_89/gnd DFFSR_2/S FILL
XFILL_26_DFFPOSX1_4 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_33_DFFSR_166 INVX1_4/gnd DFFSR_51/S FILL
XFILL_1_DFFSR_91 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_23_DFFSR_169 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_1_INVX1_38 INVX1_94/gnd DFFSR_52/S FILL
XFILL_25_DFFPOSX1_7 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_6_AND2X2_3 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_18_DFFSR_84 BUFX2_43/A DFFSR_23/S FILL
XFILL_13_DFFSR_172 BUFX2_37/A DFFSR_8/S FILL
XFILL_5_AOI22X1_4 INVX1_94/gnd DFFSR_25/S FILL
XOAI21X1_108 BUFX2_19/Y INVX1_122/Y NAND2X1_108/Y BUFX2_8/gnd DFFSR_108/D DFFSR_25/S
+ OAI21X1
XFILL_29_DFFSR_44 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_25_2_1 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_3_OAI21X1_234 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_9_DFFPOSX1_24 BUFX2_43/A DFFSR_23/S FILL
XFILL_6_NAND2X1_186 BUFX2_37/A DFFSR_81/S FILL
XFILL_3_INVX1_323 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_7_1_0 BUFX2_35/A DFFSR_97/S FILL
XFILL_0_BUFX2_29 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_23_4_2 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_9_DFFSR_166 INVX1_4/gnd DFFSR_51/S FILL
XNAND2X1_222 AND2X2_11/A DFFSR_175/Q INVX1_23/gnd XOR2X1_5/A DFFSR_186/S NAND2X1
XFILL_5_3_1 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_4_OAI21X1_168 BUFX2_36/A DFFSR_6/S FILL
XFILL_2_INVX1_143 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_3_5_2 INVX1_23/gnd DFFSR_91/S FILL
XFILL_26_DFFSR_91 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_5_AND2X2_10 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_9_DFFSR_98 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_37_DFFSR_51 INVX1_2/gnd DFFSR_51/S FILL
XFILL_48_DFFSR_11 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_4_NAND2X1_282 INVX1_89/gnd DFFSR_2/S FILL
XFILL_10_DFFSR_41 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_5_OAI21X1_102 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_0_INVX1_360 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_13_CLKBUF1_4 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_43_DFFSR_127 BUFX2_43/A DFFSR_97/S FILL
XFILL_2_OAI21X1_264 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_5_NAND2X1_216 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_34_DFFSR_98 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_33_DFFSR_130 INVX1_4/gnd DFFSR_51/S FILL
XFILL_45_DFFSR_58 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_23_DFFSR_133 BUFX2_37/A DFFSR_81/S FILL
XFILL_4_NAND3X1_114 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_1_DFFSR_55 INVX1_89/gnd DFFSR_36/S FILL
XFILL_13_DFFSR_136 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_18_DFFSR_48 INVX1_4/gnd DFFSR_4/S FILL
XFILL_8_XNOR2X1_3 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_6_NAND2X1_150 BUFX2_37/A DFFSR_81/S FILL
XFILL_3_OAI21X1_198 INVX1_8/gnd DFFSR_7/S FILL
XFILL_3_INVX1_287 INVX1_4/gnd DFFSR_51/S FILL
XNAND2X1_186 AND2X2_4/Y AND2X2_5/Y BUFX2_37/A NAND3X1_7/C DFFSR_81/S NAND2X1
XFILL_9_DFFSR_130 INVX1_4/gnd DFFSR_51/S FILL
XFILL_26_DFFSR_4 INVX1_4/gnd DFFSR_4/S FILL
XFILL_50_DFFSR_161 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_4_OAI21X1_132 INVX1_4/gnd DFFSR_4/S FILL
XFILL_9_DFFSR_62 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_15_DFFSR_95 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_26_DFFSR_55 INVX1_89/gnd DFFSR_36/S FILL
XFILL_2_INVX1_107 INVX1_89/gnd DFFSR_36/S FILL
XFILL_40_DFFSR_164 INVX1_89/gnd DFFSR_2/S FILL
XFILL_37_DFFSR_15 INVX1_8/gnd DFFSR_7/S FILL
XFILL_30_DFFSR_167 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_10_XOR2X1_15 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_20_DFFSR_170 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_4_NAND2X1_246 INVX1_94/gnd DFFSR_25/S FILL
XFILL_10_DFFSR_173 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_15_DFFPOSX1_1 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_2_AOI22X1_5 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_5_NOR2X1_49 INVX1_89/gnd DFFSR_36/S FILL
XINVX1_434 XOR2X1_16/Y INVX1_8/gnd INVX1_434/Y DFFSR_5/S INVX1
XFILL_0_INVX1_324 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_14_DFFPOSX1_4 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_8_DFFPOSX1_18 BUFX2_37/A DFFSR_8/S FILL
XFILL_34_DFFSR_62 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_5_NAND2X1_180 INVX1_94/gnd DFFSR_52/S FILL
XFILL_45_DFFSR_22 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_2_OAI21X1_228 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_13_DFFPOSX1_7 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_6_DFFSR_167 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_1_DFFSR_19 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_13_DFFSR_100 INVX1_23/gnd DFFSR_186/S FILL
XFILL_18_DFFSR_12 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_2_AND2X2_11 BUFX2_35/A DFFSR_14/S FILL
XFILL_3_OAI21X1_162 INVX1_23/gnd DFFSR_91/S FILL
XFILL_3_INVX1_251 BUFX2_36/A DFFSR_8/S FILL
XFILL_6_NAND2X1_114 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_2_INVX1_2 INVX1_2/gnd DFFSR_51/S FILL
XFILL_42_DFFSR_69 BUFX2_43/A DFFSR_23/S FILL
XFILL_9_AOI21X1_39 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_20_CLKBUF1_2 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_50_DFFSR_125 BUFX2_6/gnd DFFSR_91/S FILL
XNAND2X1_150 DFFPOSX1_1/Q DFFSR_8/S BUFX2_37/A NAND2X1_150/Y DFFSR_81/S NAND2X1
XFILL_3_NAND2X1_276 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_10_CLKBUF1_5 INVX1_89/gnd DFFSR_2/S FILL
XFILL_8_AOI21X1_42 INVX1_23/gnd DFFSR_91/S FILL
XFILL_27_DFFPOSX1_26 BUFX2_37/A DFFSR_81/S FILL
XFILL_40_DFFSR_128 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_24_5_0 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_7_AOI21X1_45 INVX1_89/gnd DFFSR_36/S FILL
XFILL_30_DFFSR_131 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_26_DFFSR_19 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_9_DFFSR_26 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_15_DFFSR_59 INVX1_4/gnd DFFSR_51/S FILL
XFILL_6_AOI21X1_48 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_20_DFFSR_134 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_1_OAI21X1_258 INVX1_2/gnd DFFSR_51/S FILL
XFILL_4_NAND2X1_210 BUFX2_35/A DFFSR_97/S FILL
XAOI21X1_48 AOI21X1_48/A AOI21X1_48/B BUFX2_10/Y DFFSR_71/gnd AOI21X1_48/Y DFFSR_45/S
+ AOI21X1
XFILL_10_DFFSR_137 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_50_DFFSR_76 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_5_XNOR2X1_4 INVX1_8/gnd DFFSR_7/S FILL
XFILL_3_NAND3X1_108 BUFX2_37/A DFFSR_81/S FILL
XINVX1_398 INVX1_331/A DFFSR_5/gnd INVX1_398/Y DFFSR_2/S INVX1
XFILL_5_NOR2X1_13 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_0_INVX1_288 INVX1_4/gnd DFFSR_4/S FILL
XFILL_2_OAI21X1_192 BUFX2_37/A DFFSR_81/S FILL
XFILL_5_NAND2X1_144 INVX1_8/gnd DFFSR_7/S FILL
XFILL_6_DFFSR_131 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_34_DFFSR_26 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_23_DFFSR_66 INVX1_2/gnd DFFSR_51/S FILL
XFILL_6_DFFSR_73 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_47_DFFSR_162 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_37_DFFSR_165 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_27_DFFSR_168 BUFX2_36/A DFFSR_8/S FILL
XFILL_5_BUFX2_11 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_3_OAI21X1_126 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_9_OAI21X1_87 INVX1_4/gnd DFFSR_4/S FILL
XFILL_3_INVX1_215 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_9_AOI22X1_3 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_17_DFFSR_171 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_8_OAI21X1_90 DFFSR_1/gnd DFFSR_1/S FILL
XOAI21X1_1 DFFSR_51/S INVX1_2/Y OAI21X1_1/C INVX1_2/gnd DFFSR_1/D DFFSR_51/S OAI21X1
XFILL_7_OAI21X1_93 INVX1_4/gnd DFFSR_51/S FILL
XFILL_42_DFFSR_33 INVX1_94/gnd DFFSR_52/S FILL
XFILL_2_NOR2X1_50 INVX1_89/gnd DFFSR_36/S FILL
XNAND2X1_114 BUFX2_17/Y INVX1_342/A DFFSR_5/gnd OAI21X1_114/C DFFSR_5/S NAND2X1
XFILL_6_OAI21X1_96 INVX1_4/gnd DFFSR_51/S FILL
XFILL_3_INVX1_67 INVX1_4/gnd DFFSR_51/S FILL
XFILL_3_XOR2X1_10 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_31_DFFSR_73 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_3_NAND2X1_240 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_34_0_0 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_5_OAI21X1_99 BUFX2_43/A DFFSR_97/S FILL
XFILL_15_DFFSR_23 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_1_INVX1_432 DFFSR_71/gnd DFFSR_45/S FILL
XOAI21X1_96 BUFX2_15/Y INVX1_108/Y OAI21X1_96/C INVX1_4/gnd DFFSR_96/D DFFSR_51/S
+ OAI21X1
XFILL_3_DFFSR_168 BUFX2_36/A DFFSR_8/S FILL
XFILL_6_AOI21X1_12 INVX1_8/gnd DFFSR_7/S FILL
XFILL_1_OAI21X1_222 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_4_NAND2X1_174 BUFX2_43/A DFFSR_97/S FILL
XFILL_5_AOI21X1_15 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_32_2_1 INVX1_8/gnd DFFSR_5/S FILL
XFILL_7_DFFPOSX1_12 INVX1_8/gnd DFFSR_5/S FILL
XFILL_3_DFFPOSX1_1 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_4_AOI21X1_18 BUFX2_8/gnd DFFSR_10/S FILL
XAOI21X1_12 AOI21X1_12/A XOR2X1_3/B INVX1_236/Y INVX1_8/gnd AOI21X1_12/Y DFFSR_7/S
+ AOI21X1
XFILL_38_DFFSR_7 INVX1_8/gnd DFFSR_7/S FILL
XFILL_10_DFFSR_101 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_3_AOI21X1_21 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_0_INVX1_252 BUFX2_36/A DFFSR_6/S FILL
XINVX1_362 INVX1_362/A DFFSR_71/gnd INVX1_362/Y DFFSR_10/S INVX1
XFILL_30_4_2 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_50_DFFSR_40 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_2_DFFPOSX1_4 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_39_DFFSR_80 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_2_AOI21X1_24 BUFX2_43/A DFFSR_97/S FILL
XFILL_1_DFFPOSX1_7 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_16_DFFPOSX1_31 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_2_OAI21X1_156 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_5_NAND2X1_108 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_17_CLKBUF1_3 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_23_DFFSR_30 INVX1_89/gnd DFFSR_36/S FILL
XFILL_6_DFFSR_37 INVX1_89/gnd DFFSR_2/S FILL
XFILL_12_DFFSR_70 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_1_AOI21X1_27 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_47_DFFSR_126 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_0_AOI21X1_30 INVX1_23/gnd DFFSR_91/S FILL
XFILL_37_DFFSR_129 INVX1_2/gnd DFFSR_1/S FILL
XFILL_2_NAND2X1_270 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_27_DFFSR_132 INVX1_2/gnd DFFSR_51/S FILL
XBUFX2_15 INVX1_1/Y BUFX2_16/gnd BUFX2_15/Y DFFSR_65/S BUFX2
XFILL_17_DFFSR_135 BUFX2_43/A DFFSR_97/S FILL
XFILL_3_INVX1_179 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_26_DFFPOSX1_20 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_47_DFFSR_87 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_8_OAI21X1_54 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_3_DFFSR_84 BUFX2_43/A DFFSR_23/S FILL
XFILL_31_DFFSR_37 INVX1_89/gnd DFFSR_2/S FILL
XFILL_3_INVX1_31 INVX1_2/gnd DFFSR_1/S FILL
XFILL_6_NAND2X1_75 INVX1_4/gnd DFFSR_4/S FILL
XFILL_7_OAI21X1_57 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_3_NAND2X1_204 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_6_OAI21X1_60 BUFX2_37/A DFFSR_81/S FILL
XFILL_20_DFFSR_77 INVX1_89/gnd DFFSR_2/S FILL
XFILL_0_OAI21X1_252 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_2_NOR2X1_14 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_5_NAND2X1_78 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_5_OAI21X1_63 INVX1_94/gnd DFFSR_25/S FILL
XFILL_4_NAND2X1_81 INVX1_94/gnd DFFSR_25/S FILL
XFILL_1_INVX1_396 DFFSR_5/gnd DFFSR_5/S FILL
XNAND2X1_75 BUFX2_24/Y DFFSR_67/Q INVX1_4/gnd OAI21X1_75/C DFFSR_4/S NAND2X1
XFILL_2_NAND3X1_102 INVX1_23/gnd DFFSR_186/S FILL
XFILL_3_NAND2X1_84 BUFX2_36/A DFFSR_6/S FILL
XOAI21X1_60 DFFSR_8/S INVX1_68/Y OAI21X1_60/C BUFX2_37/A DFFSR_60/D DFFSR_81/S OAI21X1
XFILL_2_BUFX2_22 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_3_DFFSR_132 INVX1_2/gnd DFFSR_51/S FILL
XFILL_4_OAI21X1_66 INVX1_4/gnd DFFSR_51/S FILL
XFILL_1_OAI21X1_186 BUFX2_36/A DFFSR_8/S FILL
XFILL_3_OAI21X1_69 BUFX2_37/A DFFSR_8/S FILL
XFILL_2_NAND2X1_87 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_44_DFFSR_163 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_12_NOR3X1_1 INVX1_94/gnd DFFSR_52/S FILL
XFILL_14_XOR2X1_14 INVX1_89/gnd DFFSR_2/S FILL
XFILL_2_OAI21X1_72 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_1_NAND2X1_90 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_34_DFFSR_166 INVX1_4/gnd DFFSR_51/S FILL
XFILL_4_NAND2X1_138 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_24_DFFSR_169 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_1_OAI21X1_75 INVX1_4/gnd DFFSR_4/S FILL
XFILL_0_NAND2X1_93 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_28_DFFSR_84 BUFX2_43/A DFFSR_23/S FILL
XFILL_0_INVX1_216 BUFX2_36/A DFFSR_6/S FILL
XFILL_0_INVX1_78 BUFX2_36/A DFFSR_8/S FILL
XFILL_14_DFFSR_172 BUFX2_37/A DFFSR_8/S FILL
XFILL_39_DFFSR_44 BUFX2_8/gnd DFFSR_10/S FILL
XINVX1_326 INVX1_36/A BUFX2_17/gnd INVX1_326/Y DFFSR_7/S INVX1
XFILL_0_OAI21X1_78 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_6_AOI22X1_4 INVX1_94/gnd DFFSR_25/S FILL
XFILL_2_OAI21X1_120 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_4_INVX1_323 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_12_DFFSR_34 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_0_XOR2X1_11 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_3_INVX1_143 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_0_DFFSR_169 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_9_OAI21X1_15 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_25_DFFSR_1 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_2_NAND2X1_234 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_36_DFFSR_91 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_6_AND2X2_10 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_8_OAI21X1_18 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_47_DFFSR_51 INVX1_2/gnd DFFSR_51/S FILL
XFILL_6_NAND2X1_39 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_1_NAND3X1_132 INVX1_8/gnd DFFSR_7/S FILL
XFILL_7_OAI21X1_21 INVX1_2/gnd DFFSR_51/S FILL
XFILL_0_OAI21X1_216 BUFX2_35/A DFFSR_14/S FILL
XFILL_20_DFFSR_41 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_3_DFFSR_48 INVX1_4/gnd DFFSR_4/S FILL
XFILL_5_NAND2X1_42 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_6_OAI21X1_24 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_3_NAND2X1_168 BUFX2_36/A DFFSR_6/S FILL
XNAND2X1_39 DFFSR_10/S INVX1_35/A DFFSR_71/gnd NAND2X1_39/Y DFFSR_10/S NAND2X1
XFILL_4_NAND2X1_45 INVX1_89/gnd DFFSR_36/S FILL
XFILL_1_INVX1_360 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_14_CLKBUF1_4 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_5_OAI21X1_27 DFFSR_1/gnd DFFSR_1/S FILL
XOAI21X1_24 DFFSR_11/S INVX1_27/Y NAND2X1_24/Y DFFSR_73/gnd DFFSR_24/D DFFSR_11/S
+ OAI21X1
XFILL_44_DFFSR_127 BUFX2_43/A DFFSR_97/S FILL
XFILL_4_OAI21X1_30 INVX1_89/gnd DFFSR_36/S FILL
XFILL_3_NAND2X1_48 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_15_DFFPOSX1_25 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_3_OAI21X1_33 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_1_OAI21X1_150 INVX1_94/gnd DFFSR_52/S FILL
XFILL_4_NAND2X1_102 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_44_DFFSR_98 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_2_NAND2X1_51 INVX1_2/gnd DFFSR_51/S FILL
XFILL_34_DFFSR_130 INVX1_4/gnd DFFSR_51/S FILL
XFILL_24_DFFSR_133 BUFX2_37/A DFFSR_81/S FILL
XFILL_1_NAND2X1_54 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_2_OAI21X1_36 DFFSR_79/gnd DFFSR_45/S FILL
XINVX1_290 DFFSR_12/Q BUFX2_36/A INVX1_290/Y DFFSR_8/S INVX1
XFILL_0_INVX1_180 BUFX2_37/A DFFSR_8/S FILL
XFILL_5_AND2X2_7 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_1_OAI21X1_39 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_0_DFFSR_95 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_0_INVX1_42 INVX1_89/gnd DFFSR_36/S FILL
XFILL_0_NAND2X1_57 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_28_DFFSR_48 INVX1_4/gnd DFFSR_4/S FILL
XFILL_17_DFFSR_88 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_1_NAND2X1_264 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_9_XNOR2X1_3 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_19_2 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_0_CLKBUF1_1 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_14_DFFSR_136 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_0_OAI21X1_42 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_25_DFFPOSX1_14 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_8_AOI22X1_11 INVX1_23/gnd DFFSR_91/S FILL
XFILL_7_AOI22X1_14 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_31_5_0 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_51_DFFSR_161 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_0_DFFSR_133 BUFX2_37/A DFFSR_81/S FILL
XFILL_2_NAND2X1_198 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_25_DFFSR_95 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_36_DFFSR_55 INVX1_89/gnd DFFSR_36/S FILL
XFILL_3_INVX1_107 INVX1_89/gnd DFFSR_36/S FILL
XFILL_41_DFFSR_164 INVX1_89/gnd DFFSR_2/S FILL
XFILL_47_DFFSR_15 INVX1_8/gnd DFFSR_7/S FILL
XFILL_31_DFFSR_167 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_11_XOR2X1_15 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_3_DFFSR_12 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_21_DFFSR_170 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_11_DFFSR_173 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_0_OAI21X1_180 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_3_NAND2X1_132 INVX1_8/gnd DFFSR_5/S FILL
XFILL_3_AOI22X1_5 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_6_NOR2X1_49 INVX1_89/gnd DFFSR_36/S FILL
XFILL_1_INVX1_324 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_3_NAND2X1_12 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_11_OAI22X1_50 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_44_DFFSR_62 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_10_OAI22X1_53 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_1_OAI21X1_114 INVX1_89/gnd DFFSR_36/S FILL
XFILL_2_NAND2X1_15 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_7_DFFSR_167 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_1_NAND2X1_18 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_8_NAND3X1_74 BUFX2_35/A DFFSR_14/S FILL
XFILL_9_OAI22X1_56 BUFX2_37/A DFFSR_8/S FILL
XFILL_0_NAND2X1_21 INVX1_4/gnd DFFSR_4/S FILL
XFILL_14_DFFSR_100 INVX1_23/gnd DFFSR_186/S FILL
XINVX1_254 XOR2X1_6/Y BUFX2_6/gnd INVX1_254/Y DFFSR_14/S INVX1
XFILL_28_DFFSR_12 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_3_AND2X2_11 BUFX2_35/A DFFSR_14/S FILL
XFILL_7_NAND3X1_77 BUFX2_37/A DFFSR_81/S FILL
XFILL_17_DFFSR_52 INVX1_94/gnd DFFSR_52/S FILL
XFILL_0_INVX1_144 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_8_OAI22X1_59 INVX1_8/gnd DFFSR_7/S FILL
XFILL_0_DFFSR_59 INVX1_4/gnd DFFSR_51/S FILL
XFILL_1_NAND2X1_228 INVX1_23/gnd DFFSR_91/S FILL
XFILL_4_INVX1_251 BUFX2_36/A DFFSR_8/S FILL
XFILL_6_NAND3X1_80 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_7_OAI22X1_62 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_5_NAND3X1_83 BUFX2_37/A DFFSR_81/S FILL
XFILL_41_0_0 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_6_OAI22X1_65 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_16_DFFSR_8 BUFX2_36/A DFFSR_8/S FILL
XNAND3X1_80 NAND3X1_51/Y NAND3X1_83/B NAND3X1_79/Y BUFX2_7/gnd NAND3X1_80/Y DFFSR_54/S
+ NAND3X1
XFILL_4_NAND3X1_86 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_0_NAND3X1_126 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_5_OAI22X1_68 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_51_DFFSR_125 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_3_NAND3X1_89 BUFX2_43/A DFFSR_23/S FILL
XFILL_11_CLKBUF1_5 INVX1_89/gnd DFFSR_2/S FILL
XFILL_39_2_1 BUFX2_16/gnd DFFSR_65/S FILL
XOAI22X1_65 INVX1_388/Y OAI22X1_38/D INVX1_389/Y OAI22X1_49/D DFFSR_73/gnd NOR2X1_42/B
+ DFFSR_57/S OAI22X1
XFILL_8_OAI21X1_265 BUFX2_43/A DFFSR_97/S FILL
XFILL_2_NAND3X1_92 BUFX2_43/A DFFSR_23/S FILL
XFILL_41_DFFSR_128 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_2_NAND2X1_162 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_14_DFFSR_99 BUFX2_35/A DFFSR_97/S FILL
XFILL_31_DFFSR_131 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_36_DFFSR_19 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_8_DFFSR_66 INVX1_2/gnd DFFSR_51/S FILL
XFILL_25_DFFSR_59 INVX1_4/gnd DFFSR_51/S FILL
XFILL_37_4_2 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_1_NAND3X1_95 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_0_BUFX2_9 BUFX2_37/A DFFSR_8/S FILL
XFILL_21_DFFSR_134 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_0_NAND3X1_98 BUFX2_35/A DFFSR_14/S FILL
XFILL_0_OAI21X1_144 INVX1_8/gnd DFFSR_7/S FILL
XFILL_14_DFFPOSX1_19 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_11_DFFSR_137 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_6_XNOR2X1_4 INVX1_8/gnd DFFSR_7/S FILL
XFILL_9_OAI21X1_199 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_6_NOR2X1_13 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_1_INVX1_288 INVX1_4/gnd DFFSR_4/S FILL
XFILL_37_DFFSR_4 INVX1_4/gnd DFFSR_4/S FILL
XFILL_11_OAI22X1_14 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_10_OAI22X1_17 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_41_2 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_7_DFFSR_131 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_0_NAND2X1_258 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_44_DFFSR_26 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_33_DFFSR_66 INVX1_2/gnd DFFSR_51/S FILL
XFILL_48_DFFSR_162 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_38_DFFSR_165 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_0_DFFSR_23 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_8_NAND3X1_38 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_9_OAI22X1_20 BUFX2_8/gnd DFFSR_25/S FILL
XINVX1_218 INVX1_218/A DFFSR_71/gnd XOR2X1_2/B DFFSR_10/S INVX1
XFILL_17_DFFSR_16 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_0_INVX1_108 INVX1_2/gnd DFFSR_51/S FILL
XFILL_4_DFFPOSX1_30 BUFX2_43/A DFFSR_97/S FILL
XFILL_7_NAND3X1_41 BUFX2_43/A DFFSR_23/S FILL
XFILL_1_NAND2X1_192 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_28_DFFSR_168 BUFX2_36/A DFFSR_8/S FILL
XFILL_8_OAI22X1_23 INVX1_89/gnd DFFSR_2/S FILL
XFILL_4_INVX1_215 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_6_NAND3X1_44 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_18_DFFSR_171 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_7_OAI22X1_26 INVX1_94/gnd DFFSR_52/S FILL
XFILL_5_NAND3X1_47 BUFX2_43/A DFFSR_97/S FILL
XNAND3X1_44 OAI22X1_2/Y NAND3X1_48/B NAND3X1_42/Y BUFX2_5/gnd AOI22X1_7/D DFFSR_23/S
+ NAND3X1
XFILL_6_OAI22X1_29 INVX1_8/gnd DFFSR_5/S FILL
XXOR2X1_13 XOR2X1_13/A DFFSR_140/Q INVX1_8/gnd XOR2X1_13/Y DFFSR_7/S XOR2X1
XFILL_4_NAND3X1_50 BUFX2_37/A DFFSR_81/S FILL
XFILL_0_AOI22X1_6 BUFX2_37/A DFFSR_81/S FILL
XFILL_5_OAI22X1_32 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_3_NOR2X1_50 INVX1_89/gnd DFFSR_36/S FILL
XOAI22X1_29 INVX1_314/Y OAI22X1_9/B INVX1_313/Y OAI22X1_9/D INVX1_8/gnd NOR2X1_24/B
+ DFFSR_5/S OAI22X1
XFILL_4_XOR2X1_10 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_41_DFFSR_73 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_3_NAND3X1_53 BUFX2_37/A DFFSR_81/S FILL
XDFFSR_171 AND2X2_9/B CLKBUF1_15/Y DFFSR_175/R DFFSR_52/S DFFSR_171/D BUFX2_19/gnd
+ DFFSR_52/S DFFSR
XFILL_8_OAI21X1_229 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_4_OAI22X1_35 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_2_NAND2X1_126 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_25_DFFSR_23 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_2_NAND3X1_56 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_3_OAI22X1_38 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_14_DFFSR_63 INVX1_94/gnd DFFSR_52/S FILL
XFILL_2_INVX1_432 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_8_DFFSR_30 INVX1_89/gnd DFFSR_36/S FILL
XFILL_4_DFFSR_168 BUFX2_36/A DFFSR_8/S FILL
XFILL_1_NAND3X1_59 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_2_OAI22X1_41 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_0_NAND3X1_62 BUFX2_43/A DFFSR_23/S FILL
XFILL_1_OAI22X1_44 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_0_AND2X2_12 BUFX2_43/A DFFSR_97/S FILL
XFILL_0_OAI22X1_47 BUFX2_37/A DFFSR_8/S FILL
XFILL_0_OAI21X1_108 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_11_DFFSR_101 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_1_INVX1_252 BUFX2_36/A DFFSR_6/S FILL
XFILL_49_DFFSR_80 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_0_NAND2X1_222 INVX1_23/gnd DFFSR_186/S FILL
XINVX1_64 BUFX2_7/Y BUFX2_7/gnd DFFSR_54/R DFFSR_81/S INVX1
XFILL_18_CLKBUF1_3 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_33_DFFSR_30 INVX1_89/gnd DFFSR_36/S FILL
XFILL_5_DFFSR_77 INVX1_89/gnd DFFSR_2/S FILL
XFILL_22_DFFSR_70 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_48_DFFSR_126 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_13_0_1 BUFX2_36/A DFFSR_8/S FILL
XFILL_38_DFFSR_129 INVX1_2/gnd DFFSR_1/S FILL
XINVX1_182 DFFSR_154/Q BUFX2_37/A INVX1_182/Y DFFSR_8/S INVX1
XCLKBUF1_3 DFFSR_149/Q DFFSR_79/gnd CLKBUF1_3/Y DFFSR_36/S CLKBUF1
XFILL_28_DFFSR_132 INVX1_2/gnd DFFSR_51/S FILL
XFILL_4_BUFX2_15 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_7_OAI21X1_259 INVX1_23/gnd DFFSR_186/S FILL
XFILL_9_XOR2X1_7 INVX1_23/gnd DFFSR_91/S FILL
XFILL_4_INVX1_179 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_11_2_2 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_1_NAND2X1_156 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_4_DFFSR_7 INVX1_8/gnd DFFSR_7/S FILL
XFILL_18_DFFSR_135 BUFX2_43/A DFFSR_97/S FILL
XFILL_5_NAND3X1_11 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_4_NAND3X1_14 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_2_INVX1_71 INVX1_94/gnd DFFSR_25/S FILL
XFILL_41_DFFSR_37 INVX1_89/gnd DFFSR_2/S FILL
XFILL_13_DFFPOSX1_13 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_3_NAND3X1_17 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_30_DFFSR_77 INVX1_89/gnd DFFSR_2/S FILL
XFILL_3_NOR2X1_14 DFFSR_3/gnd DFFSR_4/S FILL
XDFFSR_135 DFFSR_135/Q CLKBUF1_11/Y DFFSR_135/R DFFSR_97/S DFFSR_135/D BUFX2_43/A
+ DFFSR_97/S DFFSR
XFILL_2_NAND3X1_20 BUFX2_37/A DFFSR_8/S FILL
XFILL_8_OAI21X1_193 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_2_INVX1_396 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_1_NAND3X1_23 BUFX2_37/A DFFSR_81/S FILL
XFILL_14_DFFSR_27 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_4_DFFSR_132 INVX1_2/gnd DFFSR_51/S FILL
XFILL_45_DFFSR_163 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_0_NAND3X1_26 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_15_XOR2X1_14 INVX1_89/gnd DFFSR_2/S FILL
XFILL_35_DFFSR_166 INVX1_4/gnd DFFSR_51/S FILL
XFILL_25_DFFSR_169 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_0_OAI22X1_11 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_38_DFFSR_84 BUFX2_43/A DFFSR_23/S FILL
XFILL_1_INVX1_216 BUFX2_36/A DFFSR_6/S FILL
XFILL_15_DFFSR_172 BUFX2_37/A DFFSR_8/S FILL
XFILL_49_DFFSR_44 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_38_5_0 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_3_DFFPOSX1_24 BUFX2_43/A DFFSR_23/S FILL
XFILL_7_AOI22X1_4 INVX1_94/gnd DFFSR_25/S FILL
XFILL_0_NAND2X1_186 BUFX2_37/A DFFSR_81/S FILL
XDFFSR_81 DFFSR_81/Q CLKBUF1_6/Y DFFSR_84/R DFFSR_81/S DFFSR_81/D BUFX2_7/gnd DFFSR_81/S
+ DFFSR
XINVX1_28 BUFX2_10/Y BUFX2_19/gnd DFFSR_20/R DFFSR_54/S INVX1
XFILL_0_NOR2X1_51 INVX1_89/gnd DFFSR_36/S FILL
XFILL_5_DFFSR_41 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_22_DFFSR_34 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_11_DFFSR_74 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_1_XOR2X1_11 DFFSR_73/gnd DFFSR_57/S FILL
XINVX1_146 XOR2X1_17/A INVX1_4/gnd INVX1_146/Y DFFSR_4/S INVX1
XFILL_15_XOR2X1_4 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_1_DFFSR_169 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_49_DFFSR_7 INVX1_8/gnd DFFSR_7/S FILL
XFILL_1_NAND2X1_120 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_7_OAI21X1_223 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_46_DFFSR_91 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_7_AND2X2_10 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_4_INVX1_143 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_2_INVX1_35 BUFX2_35/A DFFSR_97/S FILL
XFILL_19_DFFSR_81 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_30_DFFSR_41 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_2_DFFSR_88 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_8_OAI21X1_157 BUFX2_35/A DFFSR_97/S FILL
XFILL_2_INVX1_360 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_15_CLKBUF1_4 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_45_DFFSR_127 BUFX2_43/A DFFSR_97/S FILL
XFILL_1_BUFX2_26 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_35_DFFSR_130 INVX1_4/gnd DFFSR_51/S FILL
XFILL_25_DFFSR_133 BUFX2_37/A DFFSR_81/S FILL
XFILL_48_0_0 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_1_INVX1_180 BUFX2_37/A DFFSR_8/S FILL
XFILL_38_DFFSR_48 INVX1_4/gnd DFFSR_4/S FILL
XFILL_27_DFFSR_88 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_1_CLKBUF1_1 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_15_DFFSR_136 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_46_2_1 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_6_OAI21X1_253 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_0_NAND2X1_150 BUFX2_37/A DFFSR_81/S FILL
XDFFSR_45 DFFSR_45/Q DFFSR_52/CLK DFFSR_46/R DFFSR_45/S DFFSR_45/D DFFSR_79/gnd DFFSR_45/S
+ DFFSR
XFILL_11_DFFSR_38 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_44_4_2 INVX1_2/gnd DFFSR_51/S FILL
XFILL_0_NOR2X1_15 INVX1_4/gnd DFFSR_51/S FILL
XFILL_8_NAND3X1_103 INVX1_23/gnd DFFSR_186/S FILL
XINVX1_110 DFFSR_97/Q BUFX2_5/gnd INVX1_110/Y DFFSR_23/S INVX1
XFILL_1_DFFSR_133 BUFX2_37/A DFFSR_81/S FILL
XFILL_7_OAI21X1_187 BUFX2_37/A DFFSR_8/S FILL
XFILL_35_DFFSR_95 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_46_DFFSR_55 INVX1_89/gnd DFFSR_36/S FILL
XFILL_4_INVX1_107 INVX1_89/gnd DFFSR_36/S FILL
XFILL_42_DFFSR_164 INVX1_89/gnd DFFSR_2/S FILL
XFILL_15_DFFSR_5 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_32_DFFSR_167 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_12_XOR2X1_15 DFFSR_79/gnd DFFSR_36/S FILL
XAOI22X1_8 AOI22X1_8/A AOI22X1_8/B AOI22X1_8/C AOI22X1_8/D BUFX2_43/A AOI22X1_8/Y
+ DFFSR_97/S AOI22X1
XFILL_22_DFFSR_170 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_2_DFFSR_52 INVX1_94/gnd DFFSR_52/S FILL
XFILL_12_DFFSR_173 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_19_DFFSR_45 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_4_AOI22X1_5 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_12_3_0 BUFX2_36/A DFFSR_6/S FILL
XFILL_8_OAI21X1_121 BUFX2_36/A DFFSR_8/S FILL
XFILL_2_INVX1_324 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_10_5_1 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_2_DFFPOSX1_18 BUFX2_37/A DFFSR_8/S FILL
XFILL_36_DFFSR_1 DFFSR_1/gnd DFFSR_1/S FILL
XAND2X2_14 NOR2X1_44/A AND2X2_14/B BUFX2_35/A NOR2X1_45/A DFFSR_97/S AND2X2
XFILL_8_DFFSR_167 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_16_DFFSR_92 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_15_DFFSR_100 INVX1_23/gnd DFFSR_186/S FILL
XFILL_38_DFFSR_12 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_4_AND2X2_11 BUFX2_35/A DFFSR_14/S FILL
XFILL_27_DFFSR_52 INVX1_94/gnd DFFSR_52/S FILL
XFILL_1_INVX1_144 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_7_NAND3X1_133 INVX1_8/gnd DFFSR_5/S FILL
XFILL_6_OAI21X1_217 INVX1_23/gnd DFFSR_91/S FILL
XFILL_0_NAND2X1_114 DFFSR_5/gnd DFFSR_5/S FILL
XOAI21X1_253 DFFSR_92/S INVX1_416/Y OAI21X1_253/C DFFSR_89/gnd DFFSR_185/D DFFSR_92/S
+ OAI21X1
XFILL_12_CLKBUF1_5 INVX1_89/gnd DFFSR_2/S FILL
XFILL_21_DFFPOSX1_26 BUFX2_37/A DFFSR_81/S FILL
XFILL_7_OAI21X1_151 BUFX2_37/A DFFSR_81/S FILL
XFILL_42_DFFSR_128 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_24_DFFSR_99 BUFX2_35/A DFFSR_97/S FILL
XFILL_32_DFFSR_131 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_46_DFFSR_19 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_35_DFFSR_59 INVX1_4/gnd DFFSR_51/S FILL
XFILL_2_DFFSR_16 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_22_DFFSR_134 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_12_DFFSR_137 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_7_XNOR2X1_4 INVX1_8/gnd DFFSR_7/S FILL
XFILL_20_0_1 INVX1_94/gnd DFFSR_52/S FILL
XFILL_2_INVX1_288 INVX1_4/gnd DFFSR_4/S FILL
XFILL_18_2_2 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_5_OAI21X1_247 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_8_DFFSR_131 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_43_DFFSR_66 INVX1_2/gnd DFFSR_51/S FILL
XFILL_49_DFFSR_162 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_0_1_1 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_39_DFFSR_165 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_27_DFFSR_16 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_1_INVX1_108 INVX1_2/gnd DFFSR_51/S FILL
XFILL_16_DFFSR_56 INVX1_2/gnd DFFSR_51/S FILL
XFILL_29_DFFSR_168 BUFX2_36/A DFFSR_8/S FILL
XFILL_16_CLKBUF1_11 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_15_CLKBUF1_14 BUFX2_43/A DFFSR_23/S FILL
XFILL_19_DFFSR_171 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_6_OAI21X1_181 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_14_CLKBUF1_17 INVX1_94/gnd DFFSR_25/S FILL
XNOR2X1_53 INVX1_432/Y NOR2X1_53/B DFFSR_79/gnd NOR2X1_53/Y DFFSR_45/S NOR2X1
XFILL_3_DFFSR_4 INVX1_4/gnd DFFSR_4/S FILL
XFILL_1_AOI22X1_6 BUFX2_37/A DFFSR_81/S FILL
XFILL_4_NOR2X1_50 INVX1_89/gnd DFFSR_36/S FILL
XFILL_13_CLKBUF1_20 INVX1_4/gnd DFFSR_51/S FILL
XFILL_5_XOR2X1_10 BUFX2_16/gnd DFFSR_11/S FILL
XOAI21X1_217 XNOR2X1_3/A INVX1_247/Y OAI21X1_217/C INVX1_23/gnd OAI21X1_218/C DFFSR_91/S
+ OAI21X1
XFILL_12_CLKBUF1_23 INVX1_89/gnd DFFSR_2/S FILL
XFILL_35_DFFSR_23 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_7_OAI21X1_115 BUFX2_36/A DFFSR_6/S FILL
XFILL_24_DFFSR_63 INVX1_94/gnd DFFSR_52/S FILL
XFILL_3_INVX1_432 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_7_DFFSR_70 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_5_DFFSR_168 BUFX2_36/A DFFSR_8/S FILL
XFILL_45_5_0 INVX1_2/gnd DFFSR_1/S FILL
XFILL_1_AND2X2_12 BUFX2_43/A DFFSR_97/S FILL
XFILL_1_DFFPOSX1_12 INVX1_8/gnd DFFSR_5/S FILL
XFILL_12_DFFSR_101 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_2_INVX1_252 BUFX2_36/A DFFSR_6/S FILL
XFILL_27_DFFSR_8 BUFX2_36/A DFFSR_8/S FILL
XFILL_6_NAND3X1_127 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_4_INVX1_64 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_19_CLKBUF1_3 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_43_DFFSR_30 INVX1_89/gnd DFFSR_36/S FILL
XFILL_10_DFFPOSX1_31 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_32_DFFSR_70 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_5_OAI21X1_211 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_49_DFFSR_126 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_39_DFFSR_129 INVX1_2/gnd DFFSR_1/S FILL
XFILL_16_DFFSR_20 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_20_DFFPOSX1_20 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_29_DFFSR_132 INVX1_2/gnd DFFSR_51/S FILL
XFILL_6_OAI21X1_145 INVX1_23/gnd DFFSR_91/S FILL
XFILL_19_DFFSR_135 BUFX2_43/A DFFSR_97/S FILL
XFILL_7_NOR3X1_1 INVX1_94/gnd DFFSR_52/S FILL
XNOR2X1_17 NOR2X1_17/A NOR2X1_17/B INVX1_4/gnd NOR2X1_17/Y DFFSR_4/S NOR2X1
XFILL_48_DFFSR_4 INVX1_4/gnd DFFSR_4/S FILL
XFILL_40_DFFSR_77 INVX1_89/gnd DFFSR_2/S FILL
XOAI21X1_181 NOR2X1_6/Y AND2X2_3/Y NAND3X1_2/A BUFX2_17/gnd OAI21X1_182/C DFFSR_57/S
+ OAI21X1
XFILL_4_NOR2X1_14 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_3_INVX1_396 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_6_NAND2X1_259 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_24_DFFSR_27 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_7_DFFSR_34 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_13_DFFSR_67 INVX1_2/gnd DFFSR_51/S FILL
XFILL_5_DFFSR_132 INVX1_2/gnd DFFSR_51/S FILL
XFILL_46_DFFSR_163 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_16_XOR2X1_14 INVX1_89/gnd DFFSR_2/S FILL
XFILL_3_INVX1_6 INVX1_8/gnd DFFSR_5/S FILL
XFILL_36_DFFSR_166 INVX1_4/gnd DFFSR_51/S FILL
XFILL_0_XOR2X1_4 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_4_OAI21X1_241 BUFX2_35/A DFFSR_97/S FILL
XFILL_26_DFFSR_169 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_48_DFFSR_84 BUFX2_43/A DFFSR_23/S FILL
XFILL_2_INVX1_216 BUFX2_36/A DFFSR_6/S FILL
XFILL_16_DFFSR_172 BUFX2_37/A DFFSR_8/S FILL
XFILL_8_AOI22X1_4 INVX1_94/gnd DFFSR_25/S FILL
XFILL_5_OAI21X1_175 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_4_DFFSR_81 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_4_INVX1_28 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_1_NOR2X1_51 INVX1_89/gnd DFFSR_36/S FILL
XFILL_32_DFFSR_34 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_21_DFFSR_74 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_2_XOR2X1_11 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_4_CLKBUF1_11 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_0_INVX1_433 DFFSR_79/gnd DFFSR_45/S FILL
XNAND3X1_127 INVX1_397/Y INVX1_398/Y INVX1_399/Y DFFSR_5/gnd NAND3X1_127/Y DFFSR_2/S
+ NAND3X1
XFILL_2_DFFSR_169 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_3_BUFX2_19 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_3_CLKBUF1_14 BUFX2_43/A DFFSR_23/S FILL
XFILL_8_AND2X2_10 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_6_OAI21X1_109 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_19_3_0 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_2_CLKBUF1_17 INVX1_94/gnd DFFSR_25/S FILL
XFILL_14_DFFSR_2 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_29_DFFSR_81 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_17_5_1 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_40_DFFSR_41 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_1_INVX1_75 INVX1_4/gnd DFFSR_51/S FILL
XFILL_1_CLKBUF1_20 INVX1_4/gnd DFFSR_51/S FILL
XOAI21X1_145 OAI21X1_145/A INVX1_164/Y OAI21X1_145/C INVX1_23/gnd DFFSR_145/D DFFSR_91/S
+ OAI21X1
XFILL_0_CLKBUF1_23 INVX1_89/gnd DFFSR_2/S FILL
XFILL_6_NAND2X1_223 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_13_DFFSR_31 BUFX2_35/A DFFSR_97/S FILL
XFILL_3_INVX1_360 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_16_CLKBUF1_4 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_46_DFFSR_127 BUFX2_43/A DFFSR_97/S FILL
XFILL_5_NAND3X1_121 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_36_DFFSR_130 INVX1_4/gnd DFFSR_51/S FILL
XNAND2X1_259 DFFSR_11/S din[4] DFFSR_73/gnd OAI21X1_248/C DFFSR_11/S NAND2X1
XFILL_4_OAI21X1_205 BUFX2_36/A DFFSR_8/S FILL
XFILL_10_1 BUFX2_43/A DFFSR_23/S FILL
XFILL_2_INVX1_180 BUFX2_37/A DFFSR_8/S FILL
XFILL_26_DFFSR_133 BUFX2_37/A DFFSR_81/S FILL
XFILL_48_DFFSR_48 INVX1_4/gnd DFFSR_4/S FILL
XFILL_37_DFFSR_88 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_2_CLKBUF1_1 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_16_DFFSR_136 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_4_DFFSR_45 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_19_DFFPOSX1_14 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_21_DFFSR_38 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_10_DFFSR_78 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_1_NOR2X1_15 INVX1_4/gnd DFFSR_51/S FILL
XFILL_5_OAI21X1_139 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_0_INVX1_397 INVX1_89/gnd DFFSR_36/S FILL
XFILL_2_DFFSR_133 BUFX2_37/A DFFSR_81/S FILL
XFILL_14_XOR2X1_8 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_5_NAND2X1_253 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_45_DFFSR_95 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_27_DFFPOSX1_2 INVX1_89/gnd DFFSR_36/S FILL
XFILL_43_DFFSR_164 INVX1_89/gnd DFFSR_2/S FILL
XFILL_33_DFFSR_167 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_13_XOR2X1_15 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_27_0_1 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_26_DFFPOSX1_5 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_23_DFFSR_170 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_6_AND2X2_4 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_25_DFFPOSX1_8 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_1_DFFSR_92 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_13_DFFSR_173 BUFX2_6/gnd DFFSR_91/S FILL
XOAI21X1_109 BUFX2_20/Y INVX1_123/Y OAI21X1_109/C BUFX2_5/gnd DFFSR_109/D DFFSR_6/S
+ OAI21X1
XFILL_18_DFFSR_85 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_29_DFFSR_45 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_1_INVX1_39 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_3_OAI21X1_235 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_5_AOI22X1_5 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_6_NAND2X1_187 BUFX2_37/A DFFSR_8/S FILL
XFILL_9_DFFPOSX1_25 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_25_2_2 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_3_INVX1_324 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_7_1_1 BUFX2_35/A DFFSR_97/S FILL
XFILL_0_BUFX2_30 INVX1_4/gnd DFFSR_51/S FILL
XNAND2X1_223 AND2X2_8/A AND2X2_11/B BUFX2_6/gnd XOR2X1_5/B DFFSR_14/S NAND2X1
XFILL_5_3_2 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_9_DFFSR_167 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_4_OAI21X1_169 BUFX2_36/A DFFSR_8/S FILL
XFILL_26_DFFSR_92 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_16_DFFSR_100 INVX1_23/gnd DFFSR_186/S FILL
XFILL_48_DFFSR_12 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_5_AND2X2_11 BUFX2_35/A DFFSR_14/S FILL
XFILL_9_DFFSR_99 BUFX2_35/A DFFSR_97/S FILL
XFILL_37_DFFSR_52 INVX1_94/gnd DFFSR_52/S FILL
XFILL_2_INVX1_144 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_4_NAND2X1_283 INVX1_89/gnd DFFSR_36/S FILL
XFILL_5_OAI21X1_103 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_10_DFFSR_42 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_0_INVX1_361 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_13_CLKBUF1_5 INVX1_89/gnd DFFSR_2/S FILL
XFILL_2_OAI21X1_265 BUFX2_43/A DFFSR_97/S FILL
XFILL_43_DFFSR_128 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_2_DFFSR_1 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_34_DFFSR_99 BUFX2_35/A DFFSR_97/S FILL
XFILL_5_NAND2X1_217 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_45_DFFSR_59 INVX1_4/gnd DFFSR_51/S FILL
XFILL_33_DFFSR_131 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_4_NAND3X1_115 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_23_DFFSR_134 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_1_DFFSR_56 INVX1_2/gnd DFFSR_51/S FILL
XFILL_18_DFFSR_49 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_13_DFFSR_137 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_3_OAI21X1_199 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_6_NAND2X1_151 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_0_OR2X2_1 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_32_1 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_8_XNOR2X1_4 INVX1_8/gnd DFFSR_7/S FILL
XFILL_3_INVX1_288 INVX1_4/gnd DFFSR_4/S FILL
XNAND2X1_187 BUFX2_11/Y AND2X2_5/B BUFX2_37/A OAI22X1_2/A DFFSR_8/S NAND2X1
XFILL_26_DFFSR_5 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_9_DFFSR_131 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_50_DFFSR_162 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_4_OAI21X1_133 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_40_DFFSR_165 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_9_DFFSR_63 INVX1_94/gnd DFFSR_52/S FILL
XFILL_37_DFFSR_16 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_15_DFFSR_96 INVX1_2/gnd DFFSR_1/S FILL
XFILL_2_INVX1_108 INVX1_2/gnd DFFSR_51/S FILL
XFILL_26_DFFSR_56 INVX1_2/gnd DFFSR_51/S FILL
XFILL_30_DFFSR_168 BUFX2_36/A DFFSR_8/S FILL
XFILL_10_XOR2X1_16 INVX1_8/gnd DFFSR_5/S FILL
XFILL_20_DFFSR_171 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_10_DFFSR_174 BUFX2_43/A DFFSR_97/S FILL
XFILL_4_NAND2X1_247 INVX1_8/gnd DFFSR_5/S FILL
XFILL_2_AOI22X1_6 BUFX2_37/A DFFSR_81/S FILL
XFILL_15_DFFPOSX1_2 INVX1_89/gnd DFFSR_36/S FILL
XFILL_5_NOR2X1_50 INVX1_89/gnd DFFSR_36/S FILL
XINVX1_435 NOR2X1_53/Y INVX1_8/gnd INVX1_435/Y DFFSR_5/S INVX1
XFILL_0_INVX1_325 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_6_XOR2X1_10 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_47_DFFSR_1 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_14_DFFPOSX1_5 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_45_DFFSR_23 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_5_NAND2X1_181 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_34_DFFSR_63 INVX1_94/gnd DFFSR_52/S FILL
XFILL_2_OAI21X1_229 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_13_DFFPOSX1_8 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_8_DFFPOSX1_19 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_6_DFFSR_168 BUFX2_36/A DFFSR_8/S FILL
XFILL_1_DFFSR_20 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_2_AND2X2_12 BUFX2_43/A DFFSR_97/S FILL
XFILL_18_DFFSR_13 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_13_DFFSR_101 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_3_INVX1_252 BUFX2_36/A DFFSR_6/S FILL
XFILL_6_NAND2X1_115 BUFX2_36/A DFFSR_6/S FILL
XFILL_2_INVX1_3 INVX1_8/gnd DFFSR_5/S FILL
XFILL_3_OAI21X1_163 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_0_NOR2X1_1 BUFX2_36/A DFFSR_6/S FILL
XFILL_20_CLKBUF1_3 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_10_CLKBUF1_6 BUFX2_5/gnd DFFSR_23/S FILL
XNAND2X1_151 INVX1_174/A DFFSR_52/S BUFX2_19/gnd OAI21X1_151/C DFFSR_52/S NAND2X1
XFILL_3_NAND2X1_277 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_26_3_0 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_42_DFFSR_70 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_50_DFFSR_126 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_27_DFFPOSX1_27 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_8_AOI21X1_43 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_40_DFFSR_129 INVX1_2/gnd DFFSR_1/S FILL
XFILL_26_DFFSR_20 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_15_DFFSR_60 BUFX2_37/A DFFSR_8/S FILL
XFILL_7_AOI21X1_46 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_9_DFFSR_27 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_24_5_1 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_30_DFFSR_132 INVX1_2/gnd DFFSR_51/S FILL
XFILL_1_OAI21X1_259 INVX1_23/gnd DFFSR_186/S FILL
XFILL_4_NAND2X1_211 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_6_4_0 BUFX2_35/A DFFSR_14/S FILL
XFILL_20_DFFSR_135 BUFX2_43/A DFFSR_97/S FILL
XFILL_10_DFFSR_138 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_3_NAND3X1_109 BUFX2_36/A DFFSR_8/S FILL
XFILL_0_INVX1_289 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_50_DFFSR_77 INVX1_89/gnd DFFSR_2/S FILL
XINVX1_399 INVX1_332/A DFFSR_5/gnd INVX1_399/Y DFFSR_2/S INVX1
XFILL_5_NOR2X1_14 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_2_OAI21X1_193 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_4_INVX1_396 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_5_NAND2X1_145 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_34_DFFSR_27 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_6_DFFSR_74 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_23_DFFSR_67 INVX1_2/gnd DFFSR_51/S FILL
XFILL_6_DFFSR_132 INVX1_2/gnd DFFSR_51/S FILL
XFILL_47_DFFSR_163 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_37_DFFSR_166 INVX1_4/gnd DFFSR_51/S FILL
XFILL_3_OAI21X1_127 BUFX2_43/A DFFSR_23/S FILL
XFILL_27_DFFSR_169 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_5_BUFX2_12 BUFX2_37/A DFFSR_81/S FILL
XFILL_9_OAI21X1_88 INVX1_4/gnd DFFSR_4/S FILL
XFILL_3_INVX1_216 BUFX2_36/A DFFSR_6/S FILL
XFILL_17_DFFSR_172 BUFX2_37/A DFFSR_8/S FILL
XFILL_8_OAI21X1_91 BUFX2_43/A DFFSR_97/S FILL
XFILL_9_AOI22X1_4 INVX1_94/gnd DFFSR_25/S FILL
XOAI21X1_2 DFFSR_5/S INVX1_3/Y OAI21X1_2/C INVX1_8/gnd DFFSR_2/D DFFSR_5/S OAI21X1
XNAND2X1_115 BUFX2_25/Y INVX1_121/A BUFX2_36/A NAND2X1_115/Y DFFSR_6/S NAND2X1
XFILL_3_INVX1_68 BUFX2_37/A DFFSR_81/S FILL
XFILL_2_NOR2X1_51 INVX1_89/gnd DFFSR_36/S FILL
XFILL_42_DFFSR_34 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_31_DFFSR_74 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_7_OAI21X1_94 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_3_XOR2X1_11 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_6_OAI21X1_97 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_3_NAND2X1_241 BUFX2_17/gnd DFFSR_57/S FILL
XOAI21X1_97 BUFX2_20/Y INVX1_110/Y OAI21X1_97/C BUFX2_5/gnd DFFSR_97/D DFFSR_23/S
+ OAI21X1
XFILL_1_INVX1_433 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_34_0_1 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_7_AOI21X1_10 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_15_DFFSR_24 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_3_DFFSR_169 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_6_AOI21X1_13 INVX1_8/gnd DFFSR_7/S FILL
XFILL_1_OAI21X1_223 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_7_DFFPOSX1_13 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_4_NAND2X1_175 BUFX2_35/A DFFSR_14/S FILL
XFILL_5_AOI21X1_16 BUFX2_43/A DFFSR_23/S FILL
XFILL_9_AND2X2_10 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_32_2_2 INVX1_8/gnd DFFSR_5/S FILL
XFILL_38_DFFSR_8 BUFX2_36/A DFFSR_8/S FILL
XFILL_4_AOI21X1_19 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_3_DFFPOSX1_2 INVX1_89/gnd DFFSR_36/S FILL
XAOI21X1_13 NAND3X1_58/A AOI21X1_13/B INVX1_235/A INVX1_8/gnd AOI21X1_13/Y DFFSR_7/S
+ AOI21X1
XFILL_10_DFFSR_102 INVX1_8/gnd DFFSR_7/S FILL
XFILL_0_INVX1_253 BUFX2_35/A DFFSR_97/S FILL
XFILL_39_DFFSR_81 BUFX2_7/gnd DFFSR_81/S FILL
XINVX1_363 DFFSR_68/Q INVX1_94/gnd INVX1_363/Y DFFSR_25/S INVX1
XFILL_50_DFFSR_41 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_2_DFFPOSX1_5 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_3_AOI21X1_22 BUFX2_43/A DFFSR_97/S FILL
XFILL_23_DFFSR_31 BUFX2_35/A DFFSR_97/S FILL
XFILL_2_OAI21X1_157 BUFX2_35/A DFFSR_97/S FILL
XFILL_2_AOI21X1_25 BUFX2_43/A DFFSR_97/S FILL
XFILL_4_INVX1_360 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_5_NAND2X1_109 INVX1_94/gnd DFFSR_25/S FILL
XFILL_17_CLKBUF1_4 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_1_DFFPOSX1_8 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_6_DFFSR_38 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_47_DFFSR_127 BUFX2_43/A DFFSR_97/S FILL
XFILL_1_AOI21X1_28 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_12_DFFSR_71 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_0_AOI21X1_31 INVX1_23/gnd DFFSR_186/S FILL
XFILL_2_NAND2X1_271 INVX1_89/gnd DFFSR_2/S FILL
XFILL_37_DFFSR_130 INVX1_4/gnd DFFSR_51/S FILL
XBUFX2_16 INVX1_1/Y BUFX2_16/gnd BUFX2_16/Y DFFSR_65/S BUFX2
XFILL_26_DFFPOSX1_21 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_3_INVX1_180 BUFX2_37/A DFFSR_8/S FILL
XFILL_27_DFFSR_133 BUFX2_37/A DFFSR_81/S FILL
XFILL_47_DFFSR_88 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_3_CLKBUF1_1 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_8_OAI21X1_55 INVX1_89/gnd DFFSR_2/S FILL
XFILL_17_DFFSR_136 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_3_INVX1_32 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_6_NAND2X1_76 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_7_OAI21X1_58 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_0_OAI21X1_253 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_3_NAND2X1_205 BUFX2_36/A DFFSR_6/S FILL
XFILL_6_OAI21X1_61 BUFX2_36/A DFFSR_8/S FILL
XFILL_3_DFFSR_85 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_5_NAND2X1_79 INVX1_89/gnd DFFSR_36/S FILL
XFILL_31_DFFSR_38 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_20_DFFSR_78 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_2_NOR2X1_15 INVX1_4/gnd DFFSR_51/S FILL
XNAND2X1_76 BUFX2_19/Y DFFSR_68/Q BUFX2_19/gnd OAI21X1_76/C DFFSR_52/S NAND2X1
XFILL_1_INVX1_397 INVX1_89/gnd DFFSR_36/S FILL
XFILL_4_NAND2X1_82 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_5_OAI21X1_64 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_2_NAND3X1_103 INVX1_23/gnd DFFSR_186/S FILL
XOAI21X1_61 DFFSR_158/S INVX1_69/Y OAI21X1_61/C BUFX2_36/A DFFSR_61/D DFFSR_8/S OAI21X1
XFILL_3_DFFSR_133 BUFX2_37/A DFFSR_81/S FILL
XFILL_2_BUFX2_23 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_3_NAND2X1_85 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_4_OAI21X1_67 INVX1_2/gnd DFFSR_1/S FILL
XFILL_44_DFFSR_164 INVX1_89/gnd DFFSR_2/S FILL
XFILL_2_NAND2X1_88 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_3_OAI21X1_70 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_1_NAND2X1_91 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_1_OAI21X1_187 BUFX2_37/A DFFSR_8/S FILL
XFILL_34_DFFSR_167 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_14_XOR2X1_15 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_12_NOR3X1_2 INVX1_89/gnd DFFSR_2/S FILL
XFILL_4_NAND2X1_139 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_2_OAI21X1_73 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_24_DFFSR_170 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_1_OAI21X1_76 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_0_NAND2X1_94 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_14_DFFSR_173 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_0_INVX1_217 INVX1_94/gnd DFFSR_25/S FILL
XFILL_28_DFFSR_85 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_39_DFFSR_45 DFFSR_79/gnd DFFSR_45/S FILL
XINVX1_327 DFFSR_64/Q BUFX2_16/gnd INVX1_327/Y DFFSR_11/S INVX1
XFILL_0_INVX1_79 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_6_AOI22X1_5 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_2_OAI21X1_121 BUFX2_36/A DFFSR_8/S FILL
XFILL_0_OAI21X1_79 INVX1_89/gnd DFFSR_36/S FILL
XFILL_4_INVX1_324 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_12_DFFSR_35 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_0_XOR2X1_12 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_0_DFFSR_170 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_9_OAI21X1_16 INVX1_89/gnd DFFSR_36/S FILL
XFILL_25_DFFSR_2 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_2_NAND2X1_235 INVX1_4/gnd DFFSR_51/S FILL
XFILL_36_DFFSR_92 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_17_DFFSR_100 INVX1_23/gnd DFFSR_186/S FILL
XFILL_6_AND2X2_11 BUFX2_35/A DFFSR_14/S FILL
XFILL_47_DFFSR_52 INVX1_94/gnd DFFSR_52/S FILL
XFILL_3_INVX1_144 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_8_OAI21X1_19 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_1_NAND3X1_133 INVX1_8/gnd DFFSR_5/S FILL
XFILL_0_OAI21X1_217 INVX1_23/gnd DFFSR_91/S FILL
XFILL_7_OAI21X1_22 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_20_DFFSR_42 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_6_NAND2X1_40 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_3_DFFSR_49 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_3_NAND2X1_169 BUFX2_36/A DFFSR_8/S FILL
XFILL_6_OAI21X1_25 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_5_NAND2X1_43 INVX1_89/gnd DFFSR_2/S FILL
XNAND2X1_40 DFFSR_11/S INVX1_36/A DFFSR_73/gnd OAI21X1_40/C DFFSR_11/S NAND2X1
XFILL_5_OAI21X1_28 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_1_INVX1_361 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_4_NAND2X1_46 BUFX2_8/gnd DFFSR_25/S FILL
XOAI21X1_25 DFFSR_10/S INVX1_29/Y OAI21X1_25/C BUFX2_8/gnd DFFSR_25/D DFFSR_10/S OAI21X1
XFILL_14_CLKBUF1_5 INVX1_89/gnd DFFSR_2/S FILL
XFILL_4_OAI21X1_31 BUFX2_35/A DFFSR_97/S FILL
XFILL_44_DFFSR_128 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_3_NAND2X1_49 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_44_DFFSR_99 BUFX2_35/A DFFSR_97/S FILL
XFILL_15_DFFPOSX1_26 BUFX2_37/A DFFSR_81/S FILL
XFILL_1_OAI21X1_151 BUFX2_37/A DFFSR_81/S FILL
XFILL_2_NAND2X1_52 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_4_NAND2X1_103 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_3_OAI21X1_34 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_2_OAI21X1_37 INVX1_89/gnd DFFSR_2/S FILL
XFILL_1_NAND2X1_55 INVX1_89/gnd DFFSR_2/S FILL
XFILL_34_DFFSR_131 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_17_DFFSR_89 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_5_AND2X2_8 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_0_INVX1_181 BUFX2_37/A DFFSR_8/S FILL
XINVX1_291 DFFSR_52/Q BUFX2_8/gnd INVX1_291/Y DFFSR_25/S INVX1
XFILL_24_DFFSR_134 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_0_INVX1_43 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_1_OAI21X1_40 INVX1_8/gnd DFFSR_7/S FILL
XFILL_0_DFFSR_96 INVX1_2/gnd DFFSR_1/S FILL
XFILL_0_NAND2X1_58 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_28_DFFSR_49 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_14_DFFSR_137 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_19_3 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_0_OAI21X1_43 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_0_CLKBUF1_2 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_1_NAND2X1_265 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_25_DFFPOSX1_15 BUFX2_35/A DFFSR_14/S FILL
XFILL_33_3_0 INVX1_8/gnd DFFSR_7/S FILL
XFILL_9_XNOR2X1_4 INVX1_8/gnd DFFSR_7/S FILL
XFILL_4_INVX1_288 INVX1_4/gnd DFFSR_4/S FILL
XFILL_8_AOI22X1_12 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_31_5_1 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_2_NAND2X1_199 BUFX2_36/A DFFSR_8/S FILL
XFILL_0_DFFSR_134 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_41_DFFSR_165 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_47_DFFSR_16 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_25_DFFSR_96 INVX1_2/gnd DFFSR_1/S FILL
XFILL_3_INVX1_108 INVX1_2/gnd DFFSR_51/S FILL
XFILL_36_DFFSR_56 INVX1_2/gnd DFFSR_51/S FILL
XFILL_31_DFFSR_168 BUFX2_36/A DFFSR_8/S FILL
XFILL_11_XOR2X1_16 INVX1_8/gnd DFFSR_5/S FILL
XFILL_21_DFFSR_171 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_11_DFFSR_174 BUFX2_43/A DFFSR_97/S FILL
XFILL_3_NAND2X1_133 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_0_OAI21X1_181 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_3_DFFSR_13 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_3_AOI22X1_6 BUFX2_37/A DFFSR_81/S FILL
XFILL_6_NOR2X1_50 INVX1_89/gnd DFFSR_36/S FILL
XFILL_4_NAND2X1_10 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_1_INVX1_325 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_7_XOR2X1_10 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_11_OAI22X1_51 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_3_NAND2X1_13 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_44_DFFSR_63 INVX1_94/gnd DFFSR_52/S FILL
XFILL_10_OAI22X1_54 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_2_NAND2X1_16 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_1_OAI21X1_115 BUFX2_36/A DFFSR_6/S FILL
XFILL_7_DFFSR_168 BUFX2_36/A DFFSR_8/S FILL
XFILL_1_NAND2X1_19 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_8_NAND3X1_75 BUFX2_35/A DFFSR_97/S FILL
XFILL_0_NAND2X1_22 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_9_OAI22X1_57 BUFX2_17/gnd DFFSR_57/S FILL
XINVX1_255 INVX1_255/A BUFX2_6/gnd OR2X2_2/B DFFSR_91/S INVX1
XFILL_3_AND2X2_12 BUFX2_43/A DFFSR_97/S FILL
XFILL_0_INVX1_145 BUFX2_43/A DFFSR_97/S FILL
XFILL_0_DFFSR_60 BUFX2_37/A DFFSR_8/S FILL
XFILL_7_NAND3X1_78 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_17_DFFSR_53 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_8_OAI22X1_60 INVX1_8/gnd DFFSR_5/S FILL
XFILL_28_DFFSR_13 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_14_DFFSR_101 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_1_NAND2X1_229 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_4_INVX1_252 BUFX2_36/A DFFSR_6/S FILL
XFILL_6_NAND3X1_81 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_7_OAI22X1_63 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_5_NAND3X1_84 INVX1_94/gnd DFFSR_25/S FILL
XFILL_6_OAI22X1_66 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_41_0_1 DFFSR_3/gnd DFFSR_4/S FILL
XNAND3X1_81 AOI21X1_19/Y NAND3X1_77/Y NAND3X1_80/Y BUFX2_19/gnd NAND3X1_81/Y DFFSR_52/S
+ NAND3X1
XFILL_4_NAND3X1_87 INVX1_94/gnd DFFSR_52/S FILL
XFILL_21_CLKBUF1_3 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_0_NAND3X1_127 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_11_CLKBUF1_6 BUFX2_5/gnd DFFSR_23/S FILL
XOAI22X1_66 INVX1_390/Y OAI22X1_38/B INVX1_391/Y OAI22X1_40/D BUFX2_17/gnd NOR2X1_42/A
+ DFFSR_7/S OAI22X1
XFILL_16_DFFSR_9 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_39_2_2 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_3_NAND3X1_90 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_2_NAND2X1_163 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_36_DFFSR_20 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_2_NAND3X1_93 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_25_DFFSR_60 BUFX2_37/A DFFSR_8/S FILL
XFILL_41_DFFSR_129 INVX1_2/gnd DFFSR_1/S FILL
XFILL_8_DFFSR_67 INVX1_2/gnd DFFSR_51/S FILL
XFILL_1_NAND3X1_96 BUFX2_43/A DFFSR_97/S FILL
XFILL_31_DFFSR_132 INVX1_2/gnd DFFSR_51/S FILL
XFILL_0_OAI21X1_145 INVX1_23/gnd DFFSR_91/S FILL
XFILL_0_NAND3X1_99 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_21_DFFSR_135 BUFX2_43/A DFFSR_97/S FILL
XFILL_14_DFFPOSX1_20 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_9_OAI21X1_200 BUFX2_37/A DFFSR_8/S FILL
XFILL_11_DFFSR_138 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_1_INVX1_289 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_37_DFFSR_5 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_11_OAI22X1_15 INVX1_4/gnd DFFSR_4/S FILL
XFILL_6_NOR2X1_14 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_10_OAI22X1_18 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_41_3 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_44_DFFSR_27 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_33_DFFSR_67 INVX1_2/gnd DFFSR_51/S FILL
XFILL_7_DFFSR_132 INVX1_2/gnd DFFSR_51/S FILL
XFILL_0_NAND2X1_259 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_48_DFFSR_163 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_0_INVX1_109 BUFX2_35/A DFFSR_97/S FILL
XFILL_8_NAND3X1_39 BUFX2_5/gnd DFFSR_23/S FILL
XINVX1_219 INVX1_219/A INVX1_94/gnd NAND3X1_4/B DFFSR_52/S INVX1
XFILL_17_DFFSR_17 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_38_DFFSR_166 INVX1_4/gnd DFFSR_51/S FILL
XFILL_0_DFFSR_24 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_9_OAI22X1_21 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_7_NAND3X1_42 BUFX2_43/A DFFSR_23/S FILL
XFILL_28_DFFSR_169 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_8_OAI22X1_24 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_4_DFFPOSX1_31 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_6_NAND3X1_45 BUFX2_35/A DFFSR_97/S FILL
XFILL_4_INVX1_216 BUFX2_36/A DFFSR_6/S FILL
XFILL_18_DFFSR_172 BUFX2_37/A DFFSR_8/S FILL
XFILL_1_NAND2X1_193 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_7_OAI22X1_27 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_5_NAND3X1_48 BUFX2_43/A DFFSR_23/S FILL
XFILL_6_OAI22X1_30 INVX1_94/gnd DFFSR_25/S FILL
XXOR2X1_14 XOR2X1_14/A AND2X2_16/Y INVX1_89/gnd XOR2X1_14/Y DFFSR_2/S XOR2X1
XNAND3X1_45 INVX1_239/A NAND3X1_35/A NAND3X1_35/C BUFX2_35/A AOI22X1_8/A DFFSR_97/S
+ NAND3X1
XFILL_0_AOI22X1_7 BUFX2_43/A DFFSR_23/S FILL
XFILL_4_NAND3X1_51 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_3_NOR2X1_51 INVX1_89/gnd DFFSR_36/S FILL
XFILL_5_OAI22X1_33 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_41_DFFSR_74 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_4_XOR2X1_11 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_2_NAND2X1_127 BUFX2_5/gnd DFFSR_6/S FILL
XDFFSR_172 AND2X2_8/B CLKBUF1_15/Y DFFSR_175/R DFFSR_8/S DFFSR_172/D BUFX2_37/A DFFSR_8/S
+ DFFSR
XFILL_3_NAND3X1_54 BUFX2_7/gnd DFFSR_54/S FILL
XOAI22X1_30 INVX1_315/Y OAI22X1_6/B INVX1_316/Y OAI22X1_6/D INVX1_94/gnd NOR2X1_24/A
+ DFFSR_25/S OAI22X1
XFILL_4_OAI22X1_36 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_8_OAI21X1_230 INVX1_23/gnd DFFSR_186/S FILL
XFILL_8_DFFSR_31 BUFX2_35/A DFFSR_97/S FILL
XFILL_3_OAI22X1_39 BUFX2_37/A DFFSR_8/S FILL
XFILL_2_NAND3X1_57 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_2_INVX1_433 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_25_DFFSR_24 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_4_DFFSR_169 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_1_NAND3X1_60 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_2_OAI22X1_42 INVX1_8/gnd DFFSR_7/S FILL
XFILL_14_DFFSR_64 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_0_NAND3X1_63 BUFX2_43/A DFFSR_23/S FILL
XFILL_1_OAI22X1_45 INVX1_89/gnd DFFSR_2/S FILL
XFILL_0_OAI21X1_109 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_0_OAI22X1_48 BUFX2_37/A DFFSR_81/S FILL
XFILL_0_AND2X2_13 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_11_DFFSR_102 INVX1_8/gnd DFFSR_7/S FILL
XFILL_1_INVX1_253 BUFX2_35/A DFFSR_97/S FILL
XFILL_49_DFFSR_81 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_1_XOR2X1_1 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_0_NAND2X1_223 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_18_CLKBUF1_4 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_5_DFFSR_78 DFFSR_1/gnd DFFSR_1/S FILL
XINVX1_65 DFFSR_57/Q DFFSR_73/gnd INVX1_65/Y DFFSR_11/S INVX1
XFILL_33_DFFSR_31 BUFX2_35/A DFFSR_97/S FILL
XFILL_48_DFFSR_127 BUFX2_43/A DFFSR_97/S FILL
XFILL_22_DFFSR_71 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_13_0_2 BUFX2_36/A DFFSR_8/S FILL
XINVX1_183 BUFX2_9/Y BUFX2_37/A DFFSR_154/R DFFSR_8/S INVX1
XCLKBUF1_4 DFFSR_149/Q BUFX2_8/gnd CLKBUF1_4/Y DFFSR_10/S CLKBUF1
XFILL_38_DFFSR_130 INVX1_4/gnd DFFSR_51/S FILL
XFILL_4_BUFX2_16 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_1_NAND2X1_157 BUFX2_35/A DFFSR_97/S FILL
XFILL_9_XOR2X1_8 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_4_DFFSR_8 BUFX2_36/A DFFSR_8/S FILL
XFILL_4_INVX1_180 BUFX2_37/A DFFSR_8/S FILL
XFILL_28_DFFSR_133 BUFX2_37/A DFFSR_81/S FILL
XFILL_7_OAI21X1_260 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_5_NAND3X1_12 INVX1_94/gnd DFFSR_52/S FILL
XFILL_4_CLKBUF1_1 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_18_DFFSR_136 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_4_NAND3X1_15 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_13_DFFPOSX1_14 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_41_DFFSR_38 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_30_DFFSR_78 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_3_NOR2X1_15 INVX1_4/gnd DFFSR_51/S FILL
XFILL_2_INVX1_72 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_8_OAI21X1_194 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_2_INVX1_397 INVX1_89/gnd DFFSR_36/S FILL
XFILL_3_NAND3X1_18 DFFSR_5/gnd DFFSR_5/S FILL
XDFFSR_136 INVX1_153/A CLKBUF1_9/Y DFFSR_135/R DFFSR_5/S DFFSR_136/D DFFSR_5/gnd DFFSR_5/S
+ DFFSR
XFILL_4_DFFSR_133 BUFX2_37/A DFFSR_81/S FILL
XFILL_2_NAND3X1_21 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_14_DFFSR_28 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_1_NAND3X1_24 BUFX2_37/A DFFSR_8/S FILL
XFILL_45_DFFSR_164 INVX1_89/gnd DFFSR_2/S FILL
XFILL_0_NAND3X1_27 BUFX2_37/A DFFSR_81/S FILL
XFILL_35_DFFSR_167 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_15_XOR2X1_15 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_40_3_0 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_25_DFFSR_170 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_0_OAI22X1_12 INVX1_4/gnd DFFSR_51/S FILL
XFILL_15_DFFSR_173 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_1_INVX1_217 INVX1_94/gnd DFFSR_25/S FILL
XFILL_38_DFFSR_85 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_49_DFFSR_45 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_38_5_1 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_7_AOI22X1_5 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_3_DFFPOSX1_25 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_0_NAND2X1_187 BUFX2_37/A DFFSR_8/S FILL
XINVX1_29 DFFSR_25/Q BUFX2_8/gnd INVX1_29/Y DFFSR_10/S INVX1
XFILL_0_NOR2X1_52 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_22_DFFSR_35 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_1_XOR2X1_12 BUFX2_17/gnd DFFSR_7/S FILL
XDFFSR_82 DFFSR_82/Q CLKBUF1_2/Y DFFSR_84/R DFFSR_9/S DFFSR_82/D DFFSR_1/gnd DFFSR_9/S
+ DFFSR
XFILL_11_DFFSR_75 INVX1_4/gnd DFFSR_51/S FILL
XFILL_5_DFFSR_42 DFFSR_3/gnd DFFSR_65/S FILL
XINVX1_147 NOR2X1_46/A INVX1_4/gnd INVX1_147/Y DFFSR_4/S INVX1
XFILL_15_XOR2X1_5 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_1_DFFSR_170 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_46_DFFSR_92 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_18_DFFSR_100 INVX1_23/gnd DFFSR_186/S FILL
XFILL_7_OAI21X1_224 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_7_AND2X2_11 BUFX2_35/A DFFSR_14/S FILL
XFILL_49_DFFSR_8 BUFX2_36/A DFFSR_8/S FILL
XFILL_1_NAND2X1_121 BUFX2_36/A DFFSR_8/S FILL
XFILL_4_INVX1_144 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_2_DFFSR_89 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_7_AND2X2_1 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_19_DFFSR_82 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_2_INVX1_36 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_30_DFFSR_42 DFFSR_3/gnd DFFSR_65/S FILL
XDFFSR_100 DFFSR_100/Q INVX1_172/A DFFSR_97/R DFFSR_186/S DFFSR_100/D INVX1_23/gnd
+ DFFSR_186/S DFFSR
XFILL_8_OAI21X1_158 BUFX2_43/A DFFSR_97/S FILL
XFILL_2_INVX1_361 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_15_CLKBUF1_5 INVX1_89/gnd DFFSR_2/S FILL
XFILL_1_BUFX2_27 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_45_DFFSR_128 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_35_DFFSR_131 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_48_0_1 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_27_DFFSR_89 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_1_INVX1_181 BUFX2_37/A DFFSR_8/S FILL
XFILL_25_DFFSR_134 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_38_DFFSR_49 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_15_DFFSR_137 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_1_CLKBUF1_2 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_46_2_2 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_6_OAI21X1_254 INVX1_23/gnd DFFSR_91/S FILL
XDFFSR_46 DFFSR_46/Q INVX1_1/A DFFSR_46/R DFFSR_6/S DFFSR_46/D BUFX2_36/A DFFSR_6/S
+ DFFSR
XFILL_0_NAND2X1_151 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_11_DFFSR_39 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_0_NOR2X1_16 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_8_NAND3X1_104 INVX1_23/gnd DFFSR_186/S FILL
XFILL_1_DFFSR_134 DFFSR_79/gnd DFFSR_45/S FILL
XINVX1_111 DFFSR_98/Q DFFSR_1/gnd INVX1_111/Y DFFSR_9/S INVX1
XFILL_42_DFFSR_165 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_15_DFFSR_6 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_7_OAI21X1_188 INVX1_89/gnd DFFSR_2/S FILL
XFILL_35_DFFSR_96 INVX1_2/gnd DFFSR_1/S FILL
XFILL_4_INVX1_108 INVX1_2/gnd DFFSR_51/S FILL
XFILL_46_DFFSR_56 INVX1_2/gnd DFFSR_51/S FILL
XFILL_32_DFFSR_168 BUFX2_36/A DFFSR_8/S FILL
XFILL_12_XOR2X1_16 INVX1_8/gnd DFFSR_5/S FILL
XAOI22X1_9 BUFX2_11/Y AOI22X1_9/B AND2X2_6/A AND2X2_10/B BUFX2_5/gnd INVX1_249/A DFFSR_23/S
+ AOI22X1
XFILL_14_1_0 BUFX2_37/A DFFSR_8/S FILL
XFILL_22_DFFSR_171 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_12_DFFSR_174 BUFX2_43/A DFFSR_97/S FILL
XFILL_19_DFFSR_46 BUFX2_36/A DFFSR_6/S FILL
XFILL_2_DFFSR_53 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_12_3_1 BUFX2_36/A DFFSR_6/S FILL
XFILL_4_AOI22X1_6 BUFX2_37/A DFFSR_81/S FILL
XFILL_8_OAI21X1_122 INVX1_94/gnd DFFSR_25/S FILL
XFILL_2_INVX1_325 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_8_XOR2X1_10 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_10_5_2 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_8_DFFSR_168 BUFX2_36/A DFFSR_8/S FILL
XFILL_36_DFFSR_2 DFFSR_5/gnd DFFSR_2/S FILL
XAND2X2_15 XOR2X1_11/A XOR2X1_11/B DFFSR_3/gnd AND2X2_15/Y DFFSR_65/S AND2X2
XFILL_2_DFFPOSX1_19 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_4_AND2X2_12 BUFX2_43/A DFFSR_97/S FILL
XFILL_1_INVX1_145 BUFX2_43/A DFFSR_97/S FILL
XFILL_27_DFFSR_53 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_7_NAND3X1_134 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_16_DFFSR_93 INVX1_2/gnd DFFSR_51/S FILL
XFILL_38_DFFSR_13 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_15_DFFSR_101 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_6_OAI21X1_218 INVX1_23/gnd DFFSR_186/S FILL
XFILL_0_NAND2X1_115 BUFX2_36/A DFFSR_6/S FILL
XDFFSR_10 DFFSR_10/Q DFFSR_52/CLK DFFSR_9/R DFFSR_10/S DFFSR_10/D DFFSR_71/gnd DFFSR_10/S
+ DFFSR
XFILL_12_CLKBUF1_6 BUFX2_5/gnd DFFSR_23/S FILL
XOAI21X1_254 DFFSR_186/S INVX1_417/Y NAND2X1_265/Y INVX1_23/gnd DFFSR_186/D DFFSR_91/S
+ OAI21X1
XFILL_21_DFFPOSX1_27 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_46_DFFSR_20 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_7_OAI21X1_152 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_35_DFFSR_60 BUFX2_37/A DFFSR_8/S FILL
XFILL_42_DFFSR_129 INVX1_2/gnd DFFSR_1/S FILL
XFILL_32_DFFSR_132 INVX1_2/gnd DFFSR_51/S FILL
XFILL_22_DFFSR_135 BUFX2_43/A DFFSR_97/S FILL
XFILL_19_DFFSR_10 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_2_DFFSR_17 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_12_DFFSR_138 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_2_INVX1_289 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_20_0_2 INVX1_94/gnd DFFSR_52/S FILL
XFILL_43_DFFSR_67 INVX1_2/gnd DFFSR_51/S FILL
XFILL_8_DFFSR_132 INVX1_2/gnd DFFSR_51/S FILL
XFILL_5_OAI21X1_248 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_49_DFFSR_163 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_0_1_2 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_1_INVX1_109 BUFX2_35/A DFFSR_97/S FILL
XFILL_27_DFFSR_17 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_16_DFFSR_57 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_39_DFFSR_166 INVX1_4/gnd DFFSR_51/S FILL
XFILL_16_CLKBUF1_12 BUFX2_43/A DFFSR_23/S FILL
XFILL_29_DFFSR_169 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_19_DFFSR_172 BUFX2_37/A DFFSR_8/S FILL
XFILL_6_OAI21X1_182 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_15_CLKBUF1_15 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_14_CLKBUF1_18 BUFX2_8/gnd DFFSR_25/S FILL
XNOR2X1_54 NOR2X1_1/B BUFX2_8/Y DFFSR_1/gnd NOR2X1_54/Y DFFSR_9/S NOR2X1
XFILL_1_AOI22X1_7 BUFX2_43/A DFFSR_23/S FILL
XFILL_4_NOR2X1_51 INVX1_89/gnd DFFSR_36/S FILL
XFILL_3_DFFSR_5 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_13_CLKBUF1_21 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_51_DFFSR_74 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_5_XOR2X1_11 DFFSR_73/gnd DFFSR_57/S FILL
XOAI21X1_218 NOR2X1_7/A NOR2X1_7/B OAI21X1_218/C INVX1_23/gnd AOI22X1_13/B DFFSR_186/S
+ OAI21X1
XFILL_12_CLKBUF1_24 INVX1_23/gnd DFFSR_186/S FILL
XFILL_47_3_0 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_7_DFFSR_71 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_3_INVX1_433 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_7_OAI21X1_116 INVX1_89/gnd DFFSR_2/S FILL
XFILL_35_DFFSR_24 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_5_DFFSR_169 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_45_5_1 INVX1_2/gnd DFFSR_1/S FILL
XFILL_24_DFFSR_64 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_1_DFFPOSX1_13 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_1_AND2X2_13 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_12_DFFSR_102 INVX1_8/gnd DFFSR_7/S FILL
XFILL_2_INVX1_253 BUFX2_35/A DFFSR_97/S FILL
XFILL_6_NAND3X1_128 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_27_DFFSR_9 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_19_CLKBUF1_4 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_43_DFFSR_31 BUFX2_35/A DFFSR_97/S FILL
XFILL_5_OAI21X1_212 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_32_DFFSR_71 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_49_DFFSR_127 BUFX2_43/A DFFSR_97/S FILL
XFILL_16_DFFSR_21 INVX1_2/gnd DFFSR_1/S FILL
XFILL_39_DFFSR_130 INVX1_4/gnd DFFSR_51/S FILL
XFILL_29_DFFSR_133 BUFX2_37/A DFFSR_81/S FILL
XFILL_6_OAI21X1_146 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_20_DFFPOSX1_21 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_5_CLKBUF1_1 BUFX2_8/gnd DFFSR_25/S FILL
XNOR2X1_18 NOR2X1_18/A NOR2X1_18/B BUFX2_8/gnd NOR2X1_18/Y DFFSR_10/S NOR2X1
XFILL_7_NOR3X1_2 INVX1_89/gnd DFFSR_2/S FILL
XFILL_19_DFFSR_136 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_48_DFFSR_5 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_40_DFFSR_78 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_4_NOR2X1_15 INVX1_4/gnd DFFSR_51/S FILL
XFILL_6_NAND2X1_260 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_3_INVX1_397 INVX1_89/gnd DFFSR_36/S FILL
XOAI21X1_182 NAND3X1_2/A NAND2X1_183/Y OAI21X1_182/C BUFX2_17/gnd DFFPOSX1_4/D DFFSR_7/S
+ OAI21X1
XFILL_13_DFFSR_68 BUFX2_35/A DFFSR_14/S FILL
XFILL_5_DFFSR_133 BUFX2_37/A DFFSR_81/S FILL
XFILL_24_DFFSR_28 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_7_DFFSR_35 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_46_DFFSR_164 INVX1_89/gnd DFFSR_2/S FILL
XFILL_3_INVX1_7 BUFX2_36/A DFFSR_8/S FILL
XFILL_36_DFFSR_167 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_0_XOR2X1_5 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_4_OAI21X1_242 BUFX2_35/A DFFSR_97/S FILL
XFILL_26_DFFSR_170 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_16_DFFSR_173 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_2_INVX1_217 INVX1_94/gnd DFFSR_25/S FILL
XFILL_48_DFFSR_85 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_8_AOI22X1_5 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_4_INVX1_29 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_1_NOR2X1_52 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_32_DFFSR_35 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_2_XOR2X1_12 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_4_DFFSR_82 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_21_DFFSR_75 INVX1_4/gnd DFFSR_51/S FILL
XFILL_5_OAI21X1_176 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_21_1_0 INVX1_94/gnd DFFSR_25/S FILL
XNAND3X1_128 INVX1_396/Y NAND3X1_128/B NAND3X1_127/Y DFFSR_5/gnd NAND3X1_128/Y DFFSR_5/S
+ NAND3X1
XFILL_0_INVX1_434 INVX1_8/gnd DFFSR_5/S FILL
XFILL_4_CLKBUF1_12 BUFX2_43/A DFFSR_23/S FILL
XFILL_3_BUFX2_20 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_2_DFFSR_170 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_19_DFFSR_100 INVX1_23/gnd DFFSR_186/S FILL
XFILL_8_AND2X2_11 BUFX2_35/A DFFSR_14/S FILL
XFILL_19_3_1 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_3_CLKBUF1_15 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_6_OAI21X1_110 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_2_CLKBUF1_18 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_14_DFFSR_3 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_1_2_0 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_17_5_2 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_1_CLKBUF1_21 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_29_DFFSR_82 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_1_INVX1_76 INVX1_2/gnd DFFSR_1/S FILL
XFILL_40_DFFSR_42 DFFSR_3/gnd DFFSR_65/S FILL
XOAI21X1_146 DFFSR_186/S INVX1_166/Y OAI21X1_146/C DFFSR_89/gnd DFFSR_146/D DFFSR_186/S
+ OAI21X1
XFILL_0_CLKBUF1_24 INVX1_23/gnd DFFSR_186/S FILL
XFILL_3_INVX1_361 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_6_NAND2X1_224 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_16_CLKBUF1_5 INVX1_89/gnd DFFSR_2/S FILL
XFILL_13_DFFSR_32 INVX1_2/gnd DFFSR_1/S FILL
XFILL_46_DFFSR_128 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_5_NAND3X1_122 DFFSR_5/gnd DFFSR_5/S FILL
XNAND2X1_260 DFFSR_186/S din[5] DFFSR_89/gnd OAI21X1_249/C DFFSR_186/S NAND2X1
XFILL_4_OAI21X1_206 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_36_DFFSR_131 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_37_DFFSR_89 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_10_2 BUFX2_43/A DFFSR_23/S FILL
XFILL_2_INVX1_181 BUFX2_37/A DFFSR_8/S FILL
XFILL_26_DFFSR_134 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_48_DFFSR_49 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_16_DFFSR_137 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_2_CLKBUF1_2 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_19_DFFPOSX1_15 BUFX2_35/A DFFSR_14/S FILL
XFILL_4_DFFSR_46 BUFX2_36/A DFFSR_6/S FILL
XFILL_5_OAI21X1_140 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_21_DFFSR_39 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_10_DFFSR_79 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_1_NOR2X1_16 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_0_INVX1_398 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_2_DFFSR_134 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_43_DFFSR_165 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_5_NAND2X1_254 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_14_XOR2X1_9 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_27_DFFPOSX1_3 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_33_DFFSR_168 BUFX2_36/A DFFSR_8/S FILL
XFILL_27_0_2 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_13_XOR2X1_16 INVX1_8/gnd DFFSR_5/S FILL
XFILL_45_DFFSR_96 INVX1_2/gnd DFFSR_1/S FILL
XFILL_26_DFFPOSX1_6 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_25_DFFPOSX1_9 BUFX2_37/A DFFSR_8/S FILL
XFILL_6_AND2X2_5 BUFX2_37/A DFFSR_81/S FILL
XFILL_23_DFFSR_171 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_13_DFFSR_174 BUFX2_43/A DFFSR_97/S FILL
XFILL_29_DFFSR_46 BUFX2_36/A DFFSR_6/S FILL
XFILL_1_INVX1_40 INVX1_8/gnd DFFSR_5/S FILL
XFILL_18_DFFSR_86 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_1_DFFSR_93 INVX1_2/gnd DFFSR_51/S FILL
XFILL_3_OAI21X1_236 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_5_AOI22X1_6 BUFX2_37/A DFFSR_81/S FILL
XFILL_9_DFFPOSX1_26 BUFX2_37/A DFFSR_81/S FILL
XFILL_6_NAND2X1_188 INVX1_8/gnd DFFSR_7/S FILL
XFILL_3_INVX1_325 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_9_XOR2X1_10 BUFX2_16/gnd DFFSR_11/S FILL
XOAI21X1_110 BUFX2_24/Y INVX1_124/Y NAND2X1_110/Y DFFSR_73/gnd DFFSR_110/D DFFSR_11/S
+ OAI21X1
XFILL_7_1_2 BUFX2_35/A DFFSR_97/S FILL
XFILL_0_BUFX2_31 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_0_OAI21X1_1 INVX1_2/gnd DFFSR_51/S FILL
XFILL_9_DFFSR_168 BUFX2_36/A DFFSR_8/S FILL
XNAND2X1_224 BUFX2_12/Y NAND2X1_224/B BUFX2_19/gnd XNOR2X1_2/B DFFSR_52/S NAND2X1
XFILL_4_OAI21X1_170 INVX1_94/gnd DFFSR_25/S FILL
XFILL_5_AND2X2_12 BUFX2_43/A DFFSR_97/S FILL
XFILL_2_INVX1_145 BUFX2_43/A DFFSR_97/S FILL
XFILL_37_DFFSR_53 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_26_DFFSR_93 INVX1_2/gnd DFFSR_51/S FILL
XFILL_48_DFFSR_13 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_16_DFFSR_101 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_10_DFFSR_43 INVX1_94/gnd DFFSR_25/S FILL
XFILL_4_DFFSR_10 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_4_NAND2X1_284 INVX1_8/gnd DFFSR_5/S FILL
XFILL_5_OAI21X1_104 INVX1_4/gnd DFFSR_51/S FILL
XFILL_13_CLKBUF1_6 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_0_INVX1_362 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_2_DFFSR_2 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_45_DFFSR_60 BUFX2_37/A DFFSR_8/S FILL
XFILL_5_NAND2X1_218 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_43_DFFSR_129 INVX1_2/gnd DFFSR_1/S FILL
XFILL_33_DFFSR_132 INVX1_2/gnd DFFSR_51/S FILL
XFILL_23_DFFSR_135 BUFX2_43/A DFFSR_97/S FILL
XFILL_29_DFFSR_10 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_4_NAND3X1_116 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_1_DFFSR_57 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_18_DFFSR_50 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_3_OAI21X1_200 BUFX2_37/A DFFSR_8/S FILL
XFILL_13_DFFSR_138 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_0_OR2X2_2 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_6_NAND2X1_152 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_3_INVX1_289 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_32_2 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_26_DFFSR_6 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_9_DFFSR_132 INVX1_2/gnd DFFSR_51/S FILL
XFILL_4_OAI21X1_134 DFFSR_79/gnd DFFSR_36/S FILL
XNAND2X1_188 INVX1_236/A AOI21X1_12/A INVX1_8/gnd XOR2X1_3/A DFFSR_7/S NAND2X1
XFILL_50_DFFSR_163 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_2_INVX1_109 BUFX2_35/A DFFSR_97/S FILL
XFILL_37_DFFSR_17 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_26_DFFSR_57 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_40_DFFSR_166 INVX1_4/gnd DFFSR_51/S FILL
XFILL_9_DFFSR_64 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_15_DFFSR_97 BUFX2_35/A DFFSR_97/S FILL
XFILL_30_DFFSR_169 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_10_XOR2X1_17 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_20_DFFSR_172 BUFX2_37/A DFFSR_8/S FILL
XFILL_10_DFFSR_175 INVX1_23/gnd DFFSR_91/S FILL
XFILL_4_NAND2X1_248 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_2_AOI22X1_7 BUFX2_43/A DFFSR_23/S FILL
XFILL_15_DFFPOSX1_3 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_5_NOR2X1_51 INVX1_89/gnd DFFSR_36/S FILL
XINVX1_436 INVX1_436/A INVX1_89/gnd INVX1_436/Y DFFSR_36/S INVX1
XFILL_0_INVX1_326 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_6_XOR2X1_11 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_47_DFFSR_2 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_14_DFFPOSX1_6 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_2_OAI21X1_230 INVX1_23/gnd DFFSR_186/S FILL
XFILL_13_DFFPOSX1_9 BUFX2_37/A DFFSR_8/S FILL
XFILL_8_DFFPOSX1_20 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_5_NAND2X1_182 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_4_INVX1_433 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_6_DFFSR_169 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_45_DFFSR_24 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_34_DFFSR_64 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_18_DFFSR_14 BUFX2_35/A DFFSR_14/S FILL
XFILL_2_AND2X2_13 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_13_DFFSR_102 INVX1_8/gnd DFFSR_7/S FILL
XFILL_1_DFFSR_21 INVX1_2/gnd DFFSR_1/S FILL
XFILL_3_INVX1_253 BUFX2_35/A DFFSR_97/S FILL
XFILL_6_NAND2X1_116 INVX1_89/gnd DFFSR_36/S FILL
XFILL_3_OAI21X1_164 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_0_NOR2X1_2 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_28_1_0 INVX1_89/gnd DFFSR_36/S FILL
XFILL_2_INVX1_4 INVX1_4/gnd DFFSR_4/S FILL
XFILL_10_CLKBUF1_7 BUFX2_43/A DFFSR_97/S FILL
XNAND2X1_152 INVX1_176/A DFFSR_23/S BUFX2_5/gnd OAI21X1_152/C DFFSR_6/S NAND2X1
XFILL_42_DFFSR_71 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_26_3_1 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_3_NAND2X1_278 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_50_DFFSR_127 BUFX2_43/A DFFSR_97/S FILL
XFILL_8_AOI21X1_44 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_27_DFFPOSX1_28 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_8_2_0 BUFX2_43/A DFFSR_97/S FILL
XFILL_7_AOI21X1_47 BUFX2_43/A DFFSR_23/S FILL
XFILL_15_DFFSR_61 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_9_DFFSR_28 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_26_DFFSR_21 INVX1_2/gnd DFFSR_1/S FILL
XFILL_40_DFFSR_130 INVX1_4/gnd DFFSR_51/S FILL
XFILL_30_DFFSR_133 BUFX2_37/A DFFSR_81/S FILL
XFILL_24_5_2 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_4_NAND2X1_212 INVX1_23/gnd DFFSR_186/S FILL
XFILL_6_4_1 BUFX2_35/A DFFSR_14/S FILL
XFILL_6_CLKBUF1_1 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_20_DFFSR_136 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_1_OAI21X1_260 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_10_DFFSR_139 DFFSR_3/gnd DFFSR_4/S FILL
XINVX1_400 BUFX2_6/Y BUFX2_35/A INVX1_400/Y DFFSR_97/S INVX1
XFILL_0_INVX1_290 BUFX2_36/A DFFSR_8/S FILL
XFILL_3_NAND3X1_110 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_50_DFFSR_78 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_5_NOR2X1_15 INVX1_4/gnd DFFSR_51/S FILL
XFILL_5_NAND2X1_146 INVX1_23/gnd DFFSR_91/S FILL
XFILL_23_DFFSR_68 BUFX2_35/A DFFSR_14/S FILL
XFILL_6_DFFSR_133 BUFX2_37/A DFFSR_81/S FILL
XFILL_2_OAI21X1_194 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_34_DFFSR_28 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_6_DFFSR_75 INVX1_4/gnd DFFSR_51/S FILL
XFILL_47_DFFSR_164 INVX1_89/gnd DFFSR_2/S FILL
XFILL_37_DFFSR_167 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_27_DFFSR_170 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_5_BUFX2_13 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_3_OAI21X1_128 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_17_DFFSR_173 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_3_INVX1_217 INVX1_94/gnd DFFSR_25/S FILL
XFILL_8_OAI21X1_92 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_9_AOI22X1_5 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_3_INVX1_69 BUFX2_36/A DFFSR_8/S FILL
XFILL_7_OAI21X1_95 INVX1_89/gnd DFFSR_36/S FILL
XFILL_42_DFFSR_35 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_3_XOR2X1_12 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_31_DFFSR_75 INVX1_4/gnd DFFSR_51/S FILL
XOAI21X1_3 DFFSR_51/S INVX1_4/Y NAND2X1_3/Y INVX1_4/gnd DFFSR_3/D DFFSR_51/S OAI21X1
XFILL_3_NAND2X1_242 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_2_NOR2X1_52 DFFSR_79/gnd DFFSR_36/S FILL
XNAND2X1_116 BUFX2_17/Y INVX1_122/A INVX1_89/gnd NAND2X1_116/Y DFFSR_36/S NAND2X1
XFILL_6_OAI21X1_98 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_7_AOI21X1_11 INVX1_8/gnd DFFSR_5/S FILL
XFILL_1_INVX1_434 INVX1_8/gnd DFFSR_5/S FILL
XFILL_34_0_2 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_6_AOI21X1_14 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_3_DFFSR_170 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_15_DFFSR_25 BUFX2_8/gnd DFFSR_25/S FILL
XOAI21X1_98 BUFX2_24/Y INVX1_111/Y NAND2X1_98/Y DFFSR_1/gnd DFFSR_98/D DFFSR_9/S OAI21X1
XFILL_20_DFFSR_100 INVX1_23/gnd DFFSR_186/S FILL
XFILL_1_OAI21X1_224 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_7_DFFPOSX1_14 BUFX2_6/gnd DFFSR_14/S FILL
XAOI21X1_14 INVX1_233/Y NAND3X1_27/C AOI21X1_4/Y BUFX2_7/gnd AOI21X1_26/C DFFSR_81/S
+ AOI21X1
XFILL_4_NAND2X1_176 INVX1_94/gnd DFFSR_25/S FILL
XFILL_5_AOI21X1_17 INVX1_8/gnd DFFSR_5/S FILL
XFILL_10_DFFSR_103 INVX1_8/gnd DFFSR_7/S FILL
XFILL_38_DFFSR_9 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_0_INVX1_254 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_4_AOI21X1_20 BUFX2_7/gnd DFFSR_81/S FILL
XINVX1_364 DFFSR_69/Q DFFSR_71/gnd INVX1_364/Y DFFSR_10/S INVX1
XFILL_3_DFFPOSX1_3 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_39_DFFSR_82 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_50_DFFSR_42 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_3_AOI21X1_23 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_2_DFFPOSX1_6 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_2_OAI21X1_158 BUFX2_43/A DFFSR_97/S FILL
XFILL_2_AOI21X1_26 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_1_DFFPOSX1_9 BUFX2_37/A DFFSR_8/S FILL
XFILL_6_DFFSR_39 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_17_CLKBUF1_5 INVX1_89/gnd DFFSR_2/S FILL
XFILL_5_NAND2X1_110 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_1_AOI21X1_29 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_12_DFFSR_72 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_23_DFFSR_32 INVX1_2/gnd DFFSR_1/S FILL
XFILL_0_AOI21X1_32 BUFX2_43/A DFFSR_23/S FILL
XFILL_47_DFFSR_128 BUFX2_19/gnd DFFSR_52/S FILL
XBUFX2_17 INVX1_1/Y BUFX2_17/gnd BUFX2_17/Y DFFSR_57/S BUFX2
XFILL_37_DFFSR_131 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_47_DFFSR_89 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_3_INVX1_181 BUFX2_37/A DFFSR_8/S FILL
XFILL_16_XOR2X1_2 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_27_DFFSR_134 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_2_NAND2X1_272 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_26_DFFPOSX1_22 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_17_DFFSR_137 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_3_CLKBUF1_2 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_8_OAI21X1_56 INVX1_2/gnd DFFSR_51/S FILL
XFILL_6_NAND2X1_77 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_7_OAI21X1_59 INVX1_4/gnd DFFSR_51/S FILL
XFILL_0_OAI21X1_254 INVX1_23/gnd DFFSR_91/S FILL
XFILL_3_NAND2X1_206 BUFX2_43/A DFFSR_97/S FILL
XFILL_6_OAI21X1_62 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_31_DFFSR_39 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_20_DFFSR_79 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_5_NAND2X1_80 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_3_DFFSR_86 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_2_NOR2X1_16 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_3_INVX1_33 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_4_NAND2X1_83 BUFX2_8/gnd DFFSR_25/S FILL
XNAND2X1_77 BUFX2_23/Y DFFSR_69/Q DFFSR_79/gnd NAND2X1_77/Y DFFSR_36/S NAND2X1
XFILL_1_INVX1_398 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_5_OAI21X1_65 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_2_NAND3X1_104 INVX1_23/gnd DFFSR_186/S FILL
XFILL_4_OAI21X1_68 BUFX2_37/A DFFSR_81/S FILL
XOAI21X1_62 DFFSR_25/S INVX1_70/Y NAND2X1_62/Y BUFX2_19/gnd DFFSR_62/D DFFSR_54/S
+ OAI21X1
XFILL_3_DFFSR_134 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_3_NAND2X1_86 INVX1_4/gnd DFFSR_51/S FILL
XFILL_44_DFFSR_165 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_2_NAND2X1_89 BUFX2_37/A DFFSR_8/S FILL
XFILL_3_OAI21X1_71 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_2_BUFX2_24 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_34_DFFSR_168 BUFX2_36/A DFFSR_8/S FILL
XFILL_4_NAND2X1_140 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_1_OAI21X1_188 INVX1_89/gnd DFFSR_2/S FILL
XFILL_14_XOR2X1_16 INVX1_8/gnd DFFSR_5/S FILL
XFILL_1_NAND2X1_92 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_24_DFFSR_171 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_2_OAI21X1_74 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_14_DFFSR_174 BUFX2_43/A DFFSR_97/S FILL
XFILL_39_DFFSR_46 BUFX2_36/A DFFSR_6/S FILL
XFILL_0_INVX1_80 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_0_INVX1_218 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_1_OAI21X1_77 INVX1_89/gnd DFFSR_36/S FILL
XFILL_0_NAND2X1_95 INVX1_89/gnd DFFSR_36/S FILL
XINVX1_328 INVX1_9/A INVX1_8/gnd INVX1_328/Y DFFSR_7/S INVX1
XFILL_28_DFFSR_86 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_6_AOI22X1_6 BUFX2_37/A DFFSR_81/S FILL
XFILL_4_INVX1_325 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_0_OAI21X1_80 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_2_OAI21X1_122 INVX1_94/gnd DFFSR_25/S FILL
XFILL_12_DFFSR_36 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_0_XOR2X1_13 INVX1_8/gnd DFFSR_7/S FILL
XFILL_1_OAI21X1_1 INVX1_2/gnd DFFSR_51/S FILL
XFILL_0_DFFSR_171 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_2_NAND2X1_236 INVX1_2/gnd DFFSR_1/S FILL
XFILL_25_DFFSR_3 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_6_AND2X2_12 BUFX2_43/A DFFSR_97/S FILL
XFILL_3_INVX1_145 BUFX2_43/A DFFSR_97/S FILL
XFILL_47_DFFSR_53 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_36_DFFSR_93 INVX1_2/gnd DFFSR_51/S FILL
XFILL_17_DFFSR_101 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_8_OAI21X1_20 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_1_NAND3X1_134 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_0_OAI21X1_218 INVX1_23/gnd DFFSR_186/S FILL
XFILL_7_OAI21X1_23 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_20_DFFSR_43 INVX1_94/gnd DFFSR_25/S FILL
XFILL_6_NAND2X1_41 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_3_DFFSR_50 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_5_NAND2X1_44 DFFSR_71/gnd DFFSR_45/S FILL
XNAND2X1_41 DFFSR_33/Q DFFSR_2/S DFFSR_5/gnd NAND2X1_41/Y DFFSR_5/S NAND2X1
XFILL_6_OAI21X1_26 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_3_NAND2X1_170 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_14_CLKBUF1_6 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_1_INVX1_362 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_4_NAND2X1_47 DFFSR_79/gnd DFFSR_45/S FILL
XOAI21X1_26 DFFSR_51/S INVX1_30/Y OAI21X1_26/C DFFSR_1/gnd DFFSR_26/D DFFSR_9/S OAI21X1
XFILL_5_OAI21X1_29 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_3_NAND2X1_50 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_4_OAI21X1_32 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_1_OAI21X1_152 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_15_DFFPOSX1_27 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_2_NAND2X1_53 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_3_OAI21X1_35 INVX1_8/gnd DFFSR_5/S FILL
XFILL_44_DFFSR_129 INVX1_2/gnd DFFSR_1/S FILL
XFILL_2_OAI21X1_38 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_35_1_0 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_34_DFFSR_132 INVX1_2/gnd DFFSR_51/S FILL
XFILL_4_NAND2X1_104 INVX1_4/gnd DFFSR_51/S FILL
XFILL_1_NAND2X1_56 INVX1_4/gnd DFFSR_51/S FILL
XFILL_5_AND2X2_9 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_0_DFFSR_97 BUFX2_35/A DFFSR_97/S FILL
XFILL_24_DFFSR_135 BUFX2_43/A DFFSR_97/S FILL
XFILL_0_INVX1_182 BUFX2_37/A DFFSR_8/S FILL
XINVX1_292 INVX1_50/A BUFX2_8/gnd INVX1_292/Y DFFSR_10/S INVX1
XFILL_39_DFFSR_10 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_0_INVX1_44 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_1_OAI21X1_41 INVX1_8/gnd DFFSR_7/S FILL
XFILL_0_NAND2X1_59 INVX1_2/gnd DFFSR_1/S FILL
XFILL_28_DFFSR_50 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_19_4 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_0_OAI21X1_44 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_0_CLKBUF1_3 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_17_DFFSR_90 INVX1_2/gnd DFFSR_1/S FILL
XFILL_14_DFFSR_138 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_25_DFFPOSX1_16 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_4_INVX1_289 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_33_3_1 INVX1_8/gnd DFFSR_7/S FILL
XFILL_1_NAND2X1_266 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_9_AOI22X1_10 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_8_AOI22X1_13 INVX1_23/gnd DFFSR_186/S FILL
XFILL_1_INVX1_1 BUFX2_37/A DFFSR_81/S FILL
XFILL_31_5_2 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_0_DFFSR_135 BUFX2_43/A DFFSR_97/S FILL
XFILL_2_NAND2X1_200 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_3_INVX1_109 BUFX2_35/A DFFSR_97/S FILL
XFILL_47_DFFSR_17 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_41_DFFSR_166 INVX1_4/gnd DFFSR_51/S FILL
XFILL_25_DFFSR_97 BUFX2_35/A DFFSR_97/S FILL
XFILL_31_DFFSR_169 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_11_XOR2X1_17 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_36_DFFSR_57 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_21_DFFSR_172 BUFX2_37/A DFFSR_8/S FILL
XFILL_11_DFFSR_175 INVX1_23/gnd DFFSR_91/S FILL
XFILL_3_DFFSR_14 BUFX2_35/A DFFSR_14/S FILL
XFILL_3_NAND2X1_134 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_0_OAI21X1_182 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_3_AOI22X1_7 BUFX2_43/A DFFSR_23/S FILL
XFILL_1_INVX1_326 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_4_NAND2X1_11 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_7_XOR2X1_11 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_3_NAND2X1_14 BUFX2_43/A DFFSR_23/S FILL
XFILL_11_OAI22X1_52 INVX1_94/gnd DFFSR_25/S FILL
XFILL_6_NOR2X1_51 INVX1_89/gnd DFFSR_36/S FILL
XFILL_10_OAI22X1_55 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_2_NAND2X1_17 INVX1_8/gnd DFFSR_7/S FILL
XFILL_1_NAND2X1_20 INVX1_23/gnd DFFSR_186/S FILL
XFILL_9_NAND3X1_73 BUFX2_43/A DFFSR_23/S FILL
XFILL_7_DFFSR_169 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_1_OAI21X1_116 INVX1_89/gnd DFFSR_2/S FILL
XFILL_44_DFFSR_64 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_8_NAND3X1_76 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_9_OAI22X1_58 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_28_DFFSR_14 BUFX2_35/A DFFSR_14/S FILL
XFILL_0_NAND2X1_23 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_0_DFFSR_61 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_7_NAND3X1_79 BUFX2_36/A DFFSR_6/S FILL
XINVX1_256 INVX1_256/A BUFX2_36/A NOR2X1_10/A DFFSR_8/S INVX1
XFILL_17_DFFSR_54 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_3_AND2X2_13 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_8_OAI22X1_61 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_14_DFFSR_102 INVX1_8/gnd DFFSR_7/S FILL
XFILL_0_INVX1_146 INVX1_4/gnd DFFSR_4/S FILL
XFILL_1_NAND2X1_230 BUFX2_36/A DFFSR_6/S FILL
XFILL_6_NAND3X1_82 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_7_OAI22X1_64 INVX1_94/gnd DFFSR_25/S FILL
XFILL_41_0_2 DFFSR_3/gnd DFFSR_4/S FILL
XNAND3X1_82 NAND3X1_51/Y NAND3X1_76/Y XOR2X1_8/A BUFX2_7/gnd NAND3X1_82/Y DFFSR_81/S
+ NAND3X1
XFILL_5_NAND3X1_85 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_0_NAND3X1_128 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_6_OAI22X1_67 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_11_CLKBUF1_7 BUFX2_43/A DFFSR_97/S FILL
XFILL_4_NAND3X1_88 INVX1_94/gnd DFFSR_52/S FILL
XOAI22X1_67 INVX1_393/Y OAI22X1_39/B INVX1_392/Y OAI22X1_39/D DFFSR_3/gnd NOR2X1_43/A
+ DFFSR_65/S OAI22X1
XFILL_3_NAND3X1_91 BUFX2_43/A DFFSR_97/S FILL
XFILL_2_NAND2X1_164 INVX1_8/gnd DFFSR_5/S FILL
XFILL_8_DFFSR_68 BUFX2_35/A DFFSR_14/S FILL
XFILL_2_NAND3X1_94 BUFX2_35/A DFFSR_97/S FILL
XFILL_25_DFFSR_61 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_36_DFFSR_21 INVX1_2/gnd DFFSR_1/S FILL
XFILL_41_DFFSR_130 INVX1_4/gnd DFFSR_51/S FILL
XFILL_1_NAND3X1_97 BUFX2_35/A DFFSR_97/S FILL
XFILL_31_DFFSR_133 BUFX2_37/A DFFSR_81/S FILL
XFILL_0_OAI21X1_146 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_14_DFFPOSX1_21 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_7_CLKBUF1_1 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_21_DFFSR_136 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_9_OAI21X1_201 BUFX2_35/A DFFSR_97/S FILL
XFILL_11_DFFSR_139 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_1_INVX1_290 BUFX2_36/A DFFSR_8/S FILL
XFILL_6_NOR2X1_15 INVX1_4/gnd DFFSR_51/S FILL
XFILL_37_DFFSR_6 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_11_OAI22X1_16 INVX1_4/gnd DFFSR_4/S FILL
XFILL_41_4 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_0_NAND2X1_260 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_33_DFFSR_68 BUFX2_35/A DFFSR_14/S FILL
XFILL_7_DFFSR_133 BUFX2_37/A DFFSR_81/S FILL
XFILL_44_DFFSR_28 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_10_OAI22X1_19 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_48_DFFSR_164 INVX1_89/gnd DFFSR_2/S FILL
XFILL_24_DFFPOSX1_10 INVX1_8/gnd DFFSR_5/S FILL
XFILL_8_NAND3X1_40 BUFX2_43/A DFFSR_23/S FILL
XFILL_0_INVX1_110 BUFX2_5/gnd DFFSR_23/S FILL
XINVX1_220 AOI22X1_1/Y INVX1_94/gnd NAND3X1_4/A DFFSR_52/S INVX1
XFILL_0_DFFSR_25 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_38_DFFSR_167 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_17_DFFSR_18 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_9_OAI22X1_22 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_7_NAND3X1_43 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_28_DFFSR_170 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_8_OAI22X1_25 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_18_DFFSR_173 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_6_NAND3X1_46 BUFX2_35/A DFFSR_97/S FILL
XFILL_1_NAND2X1_194 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_4_INVX1_217 INVX1_94/gnd DFFSR_25/S FILL
XFILL_7_OAI22X1_28 INVX1_94/gnd DFFSR_25/S FILL
XFILL_5_NAND3X1_49 BUFX2_37/A DFFSR_8/S FILL
XFILL_6_OAI22X1_31 DFFSR_71/gnd DFFSR_45/S FILL
XXOR2X1_15 XOR2X1_15/A XOR2X1_15/B DFFSR_79/gnd XOR2X1_15/Y DFFSR_36/S XOR2X1
XNAND3X1_46 INVX1_239/Y NAND3X1_36/B NAND3X1_36/C BUFX2_35/A AOI22X1_8/B DFFSR_97/S
+ NAND3X1
XFILL_0_AOI22X1_8 BUFX2_43/A DFFSR_97/S FILL
XFILL_4_NAND3X1_52 BUFX2_36/A DFFSR_8/S FILL
XFILL_4_XOR2X1_12 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_41_DFFSR_75 INVX1_4/gnd DFFSR_51/S FILL
XFILL_5_OAI22X1_34 BUFX2_16/gnd DFFSR_11/S FILL
XDFFSR_173 INVX1_246/A CLKBUF1_14/Y DFFSR_175/R DFFSR_91/S DFFSR_173/D BUFX2_6/gnd
+ DFFSR_91/S DFFSR
XFILL_3_NAND3X1_55 BUFX2_7/gnd DFFSR_54/S FILL
XOAI22X1_31 INVX1_318/Y OAI22X1_7/B INVX1_317/Y OAI22X1_7/D DFFSR_71/gnd NOR2X1_25/B
+ DFFSR_45/S OAI22X1
XFILL_4_OAI22X1_37 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_3_NOR2X1_52 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_2_NAND2X1_128 INVX1_89/gnd DFFSR_2/S FILL
XFILL_8_OAI21X1_231 BUFX2_36/A DFFSR_6/S FILL
XFILL_3_OAI22X1_40 BUFX2_37/A DFFSR_8/S FILL
XFILL_2_NAND3X1_58 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_2_INVX1_434 INVX1_8/gnd DFFSR_5/S FILL
XFILL_8_DFFSR_32 INVX1_2/gnd DFFSR_1/S FILL
XFILL_4_DFFSR_170 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_25_DFFSR_25 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_2_OAI22X1_43 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_1_NAND3X1_61 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_14_DFFSR_65 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_21_DFFSR_100 INVX1_23/gnd DFFSR_186/S FILL
XFILL_0_NAND3X1_64 BUFX2_35/A DFFSR_14/S FILL
XFILL_1_OAI22X1_46 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_0_AND2X2_14 BUFX2_35/A DFFSR_97/S FILL
XFILL_0_OAI22X1_49 INVX1_94/gnd DFFSR_25/S FILL
XFILL_11_DFFSR_103 INVX1_8/gnd DFFSR_7/S FILL
XFILL_0_OAI21X1_110 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_1_INVX1_254 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_1_XOR2X1_2 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_49_DFFSR_82 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_0_NAND2X1_224 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_18_CLKBUF1_5 INVX1_89/gnd DFFSR_2/S FILL
XINVX1_66 INVX1_66/A DFFSR_3/gnd INVX1_66/Y DFFSR_65/S INVX1
XFILL_5_DFFSR_79 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_22_DFFSR_72 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_33_DFFSR_32 INVX1_2/gnd DFFSR_1/S FILL
XFILL_48_DFFSR_128 BUFX2_19/gnd DFFSR_52/S FILL
XINVX1_184 INVX1_184/A BUFX2_7/gnd INVX1_184/Y DFFSR_81/S INVX1
XCLKBUF1_5 DFFSR_149/Q INVX1_89/gnd CLKBUF1_5/Y DFFSR_2/S CLKBUF1
XFILL_38_DFFSR_131 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_1_NAND2X1_158 BUFX2_35/A DFFSR_97/S FILL
XFILL_4_INVX1_181 BUFX2_37/A DFFSR_8/S FILL
XFILL_6_NAND3X1_10 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_9_XOR2X1_9 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_28_DFFSR_134 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_7_OAI21X1_261 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_4_BUFX2_17 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_18_DFFSR_137 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_4_CLKBUF1_2 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_4_DFFSR_9 DFFSR_9/gnd DFFSR_9/S FILL
XNAND3X1_10 NAND3X1_8/A AOI22X1_3/C NAND3X1_7/C BUFX2_7/gnd AOI21X1_8/A DFFSR_54/S
+ NAND3X1
XFILL_5_NAND3X1_13 INVX1_94/gnd DFFSR_25/S FILL
XFILL_13_DFFPOSX1_15 BUFX2_35/A DFFSR_14/S FILL
XFILL_2_INVX1_73 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_4_NAND3X1_16 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_41_DFFSR_39 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_30_DFFSR_79 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_3_NOR2X1_16 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_8_OAI21X1_195 BUFX2_7/gnd DFFSR_81/S FILL
XDFFSR_137 DFFSR_137/Q CLKBUF1_11/Y DFFSR_137/R DFFSR_54/S DFFSR_137/D BUFX2_7/gnd
+ DFFSR_54/S DFFSR
XFILL_3_NAND3X1_19 INVX1_8/gnd DFFSR_5/S FILL
XFILL_2_NAND3X1_22 BUFX2_37/A DFFSR_81/S FILL
XFILL_4_DFFSR_134 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_2_INVX1_398 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_42_1_0 INVX1_4/gnd DFFSR_4/S FILL
XFILL_14_DFFSR_29 INVX1_4/gnd DFFSR_4/S FILL
XFILL_45_DFFSR_165 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_1_NAND3X1_25 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_35_DFFSR_168 BUFX2_36/A DFFSR_8/S FILL
XFILL_0_NAND3X1_28 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_15_XOR2X1_16 INVX1_8/gnd DFFSR_5/S FILL
XFILL_1_OAI22X1_10 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_40_3_1 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_25_DFFSR_171 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_9_OAI21X1_129 INVX1_4/gnd DFFSR_4/S FILL
XFILL_0_OAI22X1_13 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_15_DFFSR_174 BUFX2_43/A DFFSR_97/S FILL
XFILL_49_DFFSR_46 BUFX2_36/A DFFSR_6/S FILL
XFILL_1_INVX1_218 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_38_DFFSR_86 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_38_5_2 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_7_AOI22X1_6 BUFX2_37/A DFFSR_81/S FILL
XFILL_3_DFFPOSX1_26 BUFX2_37/A DFFSR_81/S FILL
XFILL_11_DFFSR_76 BUFX2_7/gnd DFFSR_54/S FILL
XDFFSR_83 DFFSR_83/Q CLKBUF1_6/Y DFFSR_84/R DFFSR_52/S DFFSR_83/D BUFX2_19/gnd DFFSR_54/S
+ DFFSR
XFILL_5_DFFSR_43 INVX1_94/gnd DFFSR_25/S FILL
XFILL_22_DFFSR_36 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_0_NAND2X1_188 INVX1_8/gnd DFFSR_7/S FILL
XINVX1_30 INVX1_30/A DFFSR_1/gnd INVX1_30/Y DFFSR_9/S INVX1
XFILL_0_NOR2X1_53 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_1_XOR2X1_13 INVX1_8/gnd DFFSR_7/S FILL
XFILL_2_OAI21X1_1 INVX1_2/gnd DFFSR_51/S FILL
XINVX1_148 XOR2X1_11/A DFFSR_1/gnd INVX1_148/Y DFFSR_9/S INVX1
XFILL_1_DFFSR_171 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_15_XOR2X1_6 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_7_OAI21X1_225 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_7_AND2X2_12 BUFX2_43/A DFFSR_97/S FILL
XFILL_4_INVX1_145 BUFX2_43/A DFFSR_97/S FILL
XFILL_1_NAND2X1_122 INVX1_94/gnd DFFSR_25/S FILL
XFILL_49_DFFSR_9 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_46_DFFSR_93 INVX1_2/gnd DFFSR_51/S FILL
XFILL_18_DFFSR_101 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_7_AND2X2_2 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_19_DFFSR_83 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_2_INVX1_37 INVX1_94/gnd DFFSR_52/S FILL
XFILL_30_DFFSR_43 INVX1_94/gnd DFFSR_25/S FILL
XFILL_2_DFFSR_90 INVX1_2/gnd DFFSR_1/S FILL
XDFFSR_101 INVX1_368/A CLKBUF1_4/Y DFFSR_97/R DFFSR_57/S DFFSR_101/D DFFSR_73/gnd
+ DFFSR_57/S DFFSR
XFILL_8_OAI21X1_159 BUFX2_43/A DFFSR_97/S FILL
XFILL_15_CLKBUF1_6 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_2_INVX1_362 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_1_BUFX2_28 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_45_DFFSR_129 INVX1_2/gnd DFFSR_1/S FILL
XFILL_48_0_2 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_35_DFFSR_132 INVX1_2/gnd DFFSR_51/S FILL
XFILL_25_DFFSR_135 BUFX2_43/A DFFSR_97/S FILL
XFILL_1_INVX1_182 BUFX2_37/A DFFSR_8/S FILL
XFILL_49_DFFSR_10 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_38_DFFSR_50 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_23_1 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_1_CLKBUF1_3 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_27_DFFSR_90 INVX1_2/gnd DFFSR_1/S FILL
XFILL_15_DFFSR_138 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_0_NAND2X1_152 BUFX2_5/gnd DFFSR_6/S FILL
XDFFSR_47 INVX1_53/A DFFSR_28/CLK DFFSR_46/R DFFSR_2/S DFFSR_47/D DFFSR_5/gnd DFFSR_2/S
+ DFFSR
XFILL_11_DFFSR_40 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_0_NOR2X1_17 INVX1_4/gnd DFFSR_4/S FILL
XFILL_6_OAI21X1_255 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_8_NAND3X1_105 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_1_DFFSR_135 BUFX2_43/A DFFSR_97/S FILL
XINVX1_112 DFFSR_99/Q BUFX2_43/A INVX1_112/Y DFFSR_97/S INVX1
XFILL_4_INVX1_109 BUFX2_35/A DFFSR_97/S FILL
XFILL_15_DFFSR_7 INVX1_8/gnd DFFSR_7/S FILL
XFILL_7_OAI21X1_189 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_42_DFFSR_166 INVX1_4/gnd DFFSR_51/S FILL
XFILL_35_DFFSR_97 BUFX2_35/A DFFSR_97/S FILL
XFILL_32_DFFSR_169 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_12_XOR2X1_17 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_46_DFFSR_57 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_22_DFFSR_172 BUFX2_37/A DFFSR_8/S FILL
XFILL_14_1_1 BUFX2_37/A DFFSR_8/S FILL
XFILL_12_DFFSR_175 INVX1_23/gnd DFFSR_91/S FILL
XFILL_2_DFFSR_54 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_19_DFFSR_47 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_8_OAI21X1_123 INVX1_23/gnd DFFSR_91/S FILL
XFILL_4_AOI22X1_7 BUFX2_43/A DFFSR_23/S FILL
XFILL_12_3_2 BUFX2_36/A DFFSR_6/S FILL
XFILL_2_INVX1_326 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_8_XOR2X1_11 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_8_DFFSR_169 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_2_DFFPOSX1_20 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_36_DFFSR_3 DFFSR_3/gnd DFFSR_4/S FILL
XAND2X2_16 AND2X2_16/A AND2X2_16/B DFFSR_79/gnd AND2X2_16/Y DFFSR_45/S AND2X2
XFILL_38_DFFSR_14 BUFX2_35/A DFFSR_14/S FILL
XFILL_27_DFFSR_54 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_4_AND2X2_13 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_15_DFFSR_102 INVX1_8/gnd DFFSR_7/S FILL
XFILL_1_INVX1_146 INVX1_4/gnd DFFSR_4/S FILL
XFILL_16_DFFSR_94 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_6_OAI21X1_219 BUFX2_35/A DFFSR_97/S FILL
XFILL_0_NAND2X1_116 INVX1_89/gnd DFFSR_36/S FILL
XDFFSR_11 DFFSR_11/Q DFFSR_3/CLK DFFSR_9/R DFFSR_11/S DFFSR_11/D BUFX2_16/gnd DFFSR_11/S
+ DFFSR
XFILL_12_CLKBUF1_7 BUFX2_43/A DFFSR_97/S FILL
XOAI21X1_255 DFFSR_4/S INVX1_418/Y NAND2X1_266/Y DFFSR_3/gnd DFFSR_187/D DFFSR_4/S
+ OAI21X1
XFILL_35_DFFSR_61 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_7_OAI21X1_153 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_46_DFFSR_21 INVX1_2/gnd DFFSR_1/S FILL
XFILL_42_DFFSR_130 INVX1_4/gnd DFFSR_51/S FILL
XFILL_21_DFFPOSX1_28 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_32_DFFSR_133 BUFX2_37/A DFFSR_81/S FILL
XFILL_8_CLKBUF1_1 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_22_DFFSR_136 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_2_DFFSR_18 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_19_DFFSR_11 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_12_DFFSR_139 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_2_INVX1_290 BUFX2_36/A DFFSR_8/S FILL
XFILL_45_1 INVX1_2/gnd DFFSR_51/S FILL
XFILL_43_DFFSR_68 BUFX2_35/A DFFSR_14/S FILL
XFILL_8_DFFSR_133 BUFX2_37/A DFFSR_81/S FILL
XFILL_5_OAI21X1_249 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_49_DFFSR_164 INVX1_89/gnd DFFSR_2/S FILL
XFILL_1_INVX1_110 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_39_DFFSR_167 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_17_CLKBUF1_10 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_29_DFFSR_170 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_27_DFFSR_18 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_16_CLKBUF1_13 INVX1_4/gnd DFFSR_51/S FILL
XFILL_16_DFFSR_58 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_19_DFFSR_173 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_15_CLKBUF1_16 BUFX2_36/A DFFSR_6/S FILL
XFILL_6_OAI21X1_183 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_14_CLKBUF1_19 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_1_AOI22X1_8 BUFX2_43/A DFFSR_97/S FILL
XFILL_3_DFFSR_6 BUFX2_5/gnd DFFSR_6/S FILL
XOAI21X1_219 INVX1_249/A NOR2X1_9/Y INVX1_248/A BUFX2_35/A NAND3X1_68/B DFFSR_97/S
+ OAI21X1
XFILL_13_CLKBUF1_22 INVX1_94/gnd DFFSR_25/S FILL
XFILL_4_NOR2X1_52 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_5_XOR2X1_12 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_47_3_1 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_12_CLKBUF1_25 INVX1_23/gnd DFFSR_186/S FILL
XFILL_7_OAI21X1_117 BUFX2_35/A DFFSR_97/S FILL
XFILL_3_INVX1_434 INVX1_8/gnd DFFSR_5/S FILL
XFILL_5_DFFSR_170 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_35_DFFSR_25 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_7_DFFSR_72 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_24_DFFSR_65 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_22_DFFSR_100 INVX1_23/gnd DFFSR_186/S FILL
XFILL_45_5_2 INVX1_2/gnd DFFSR_1/S FILL
XFILL_1_DFFPOSX1_14 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_1_AND2X2_14 BUFX2_35/A DFFSR_97/S FILL
XFILL_6_BUFX2_10 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_12_DFFSR_103 INVX1_8/gnd DFFSR_7/S FILL
XFILL_2_INVX1_254 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_6_NAND3X1_129 BUFX2_35/A DFFSR_14/S FILL
XFILL_19_CLKBUF1_5 INVX1_89/gnd DFFSR_2/S FILL
XFILL_5_OAI21X1_213 BUFX2_36/A DFFSR_6/S FILL
XFILL_32_DFFSR_72 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_43_DFFSR_32 INVX1_2/gnd DFFSR_1/S FILL
XFILL_13_4_0 BUFX2_36/A DFFSR_8/S FILL
XFILL_49_DFFSR_128 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_16_DFFSR_22 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_39_DFFSR_131 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_29_DFFSR_134 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_6_OAI21X1_147 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_19_DFFSR_137 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_5_CLKBUF1_2 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_20_DFFPOSX1_22 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_48_DFFSR_6 BUFX2_5/gnd DFFSR_6/S FILL
XNOR2X1_19 NOR2X1_19/A NOR2X1_19/B BUFX2_8/gnd NOR2X1_19/Y DFFSR_10/S NOR2X1
XFILL_51_DFFSR_39 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_40_DFFSR_79 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_4_NOR2X1_16 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_6_NAND2X1_261 BUFX2_8/gnd DFFSR_10/S FILL
XOAI21X1_183 NOR2X1_5/A AND2X2_3/B NAND3X1_6/Y BUFX2_17/gnd XOR2X1_3/B DFFSR_7/S OAI21X1
XFILL_13_DFFSR_69 BUFX2_43/A DFFSR_23/S FILL
XFILL_5_DFFSR_134 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_7_DFFSR_36 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_3_INVX1_398 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_24_DFFSR_29 INVX1_4/gnd DFFSR_4/S FILL
XFILL_46_DFFSR_165 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_36_DFFSR_168 BUFX2_36/A DFFSR_8/S FILL
XFILL_0_XOR2X1_6 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_4_OAI21X1_243 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_26_DFFSR_171 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_3_INVX1_8 INVX1_8/gnd DFFSR_5/S FILL
XFILL_16_DFFSR_174 BUFX2_43/A DFFSR_97/S FILL
XFILL_2_INVX1_218 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_48_DFFSR_86 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_8_AOI22X1_6 BUFX2_37/A DFFSR_81/S FILL
XFILL_21_DFFSR_76 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_4_DFFSR_83 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_32_DFFSR_36 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_4_INVX1_30 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_5_OAI21X1_177 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_1_NOR2X1_53 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_2_XOR2X1_13 INVX1_8/gnd DFFSR_7/S FILL
XFILL_3_OAI21X1_1 INVX1_2/gnd DFFSR_51/S FILL
XNAND3X1_129 INVX1_1/A INVX1_401/A NOR2X1_45/A BUFX2_35/A AOI21X1_42/A DFFSR_14/S
+ NAND3X1
XFILL_21_1_1 INVX1_94/gnd DFFSR_25/S FILL
XFILL_0_INVX1_435 INVX1_8/gnd DFFSR_5/S FILL
XFILL_5_CLKBUF1_10 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_3_0_0 INVX1_23/gnd DFFSR_91/S FILL
XFILL_3_BUFX2_21 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_2_DFFSR_171 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_4_CLKBUF1_13 INVX1_4/gnd DFFSR_51/S FILL
XFILL_8_AND2X2_12 BUFX2_43/A DFFSR_97/S FILL
XFILL_3_CLKBUF1_16 BUFX2_36/A DFFSR_6/S FILL
XFILL_19_3_2 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_6_OAI21X1_111 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_19_DFFSR_101 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_2_CLKBUF1_19 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_14_DFFSR_4 INVX1_4/gnd DFFSR_4/S FILL
XFILL_1_2_1 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_1_INVX1_77 BUFX2_37/A DFFSR_81/S FILL
XFILL_29_DFFSR_83 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_40_DFFSR_43 INVX1_94/gnd DFFSR_25/S FILL
XFILL_1_CLKBUF1_22 INVX1_94/gnd DFFSR_25/S FILL
XOAI21X1_147 DFFSR_186/S INVX1_168/Y NAND2X1_147/Y DFFSR_89/gnd DFFSR_147/D DFFSR_186/S
+ OAI21X1
XFILL_0_CLKBUF1_25 INVX1_23/gnd DFFSR_186/S FILL
XFILL_16_CLKBUF1_6 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_6_NAND2X1_225 BUFX2_36/A DFFSR_8/S FILL
XFILL_3_INVX1_362 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_13_DFFSR_33 INVX1_94/gnd DFFSR_52/S FILL
XFILL_5_NAND3X1_123 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_46_DFFSR_129 INVX1_2/gnd DFFSR_1/S FILL
XFILL_4_OAI21X1_207 BUFX2_37/A DFFSR_8/S FILL
XNAND2X1_261 DFFSR_10/S din[6] BUFX2_8/gnd NAND2X1_261/Y DFFSR_10/S NAND2X1
XFILL_36_DFFSR_132 INVX1_2/gnd DFFSR_51/S FILL
XFILL_26_DFFSR_135 BUFX2_43/A DFFSR_97/S FILL
XFILL_10_3 BUFX2_43/A DFFSR_23/S FILL
XFILL_2_INVX1_182 BUFX2_37/A DFFSR_8/S FILL
XFILL_48_DFFSR_50 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_2_CLKBUF1_3 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_37_DFFSR_90 INVX1_2/gnd DFFSR_1/S FILL
XFILL_16_DFFSR_138 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_19_DFFPOSX1_16 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_5_OAI21X1_141 INVX1_94/gnd DFFSR_52/S FILL
XFILL_4_DFFSR_47 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_21_DFFSR_40 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_1_NOR2X1_17 INVX1_4/gnd DFFSR_4/S FILL
XFILL_10_DFFSR_80 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_2_DFFSR_135 BUFX2_43/A DFFSR_97/S FILL
XFILL_0_INVX1_399 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_27_DFFPOSX1_4 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_43_DFFSR_166 INVX1_4/gnd DFFSR_51/S FILL
XFILL_45_DFFSR_97 BUFX2_35/A DFFSR_97/S FILL
XFILL_33_DFFSR_169 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_13_XOR2X1_17 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_26_DFFPOSX1_7 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_5_NAND2X1_255 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_6_AND2X2_6 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_23_DFFSR_172 BUFX2_37/A DFFSR_8/S FILL
XFILL_13_DFFSR_175 INVX1_23/gnd DFFSR_91/S FILL
XFILL_1_INVX1_41 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_29_DFFSR_47 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_18_DFFSR_87 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_1_DFFSR_94 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_5_AOI22X1_7 BUFX2_43/A DFFSR_23/S FILL
XFILL_6_NAND2X1_189 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_3_OAI21X1_237 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_9_DFFPOSX1_27 DFFSR_71/gnd DFFSR_45/S FILL
XOAI21X1_111 BUFX2_22/Y INVX1_125/Y NAND2X1_111/Y DFFSR_5/gnd DFFSR_111/D DFFSR_5/S
+ OAI21X1
XFILL_3_INVX1_326 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_9_XOR2X1_11 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_0_OAI21X1_2 INVX1_8/gnd DFFSR_5/S FILL
XFILL_0_BUFX2_32 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_9_DFFSR_169 BUFX2_5/gnd DFFSR_6/S FILL
XNAND2X1_225 NOR2X1_10/Y INVX1_257/Y BUFX2_36/A NAND3X1_92/C DFFSR_8/S NAND2X1
XFILL_4_OAI21X1_171 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_48_DFFSR_14 BUFX2_35/A DFFSR_14/S FILL
XFILL_37_DFFSR_54 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_5_AND2X2_13 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_16_DFFSR_102 INVX1_8/gnd DFFSR_7/S FILL
XFILL_2_INVX1_146 INVX1_4/gnd DFFSR_4/S FILL
XFILL_26_DFFSR_94 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_10_DFFSR_44 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_4_NAND2X1_285 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_4_DFFSR_11 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_5_OAI21X1_105 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_13_CLKBUF1_7 BUFX2_43/A DFFSR_97/S FILL
XFILL_0_INVX1_363 INVX1_94/gnd DFFSR_25/S FILL
XFILL_2_DFFSR_3 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_45_DFFSR_61 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_5_NAND2X1_219 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_43_DFFSR_130 INVX1_4/gnd DFFSR_51/S FILL
XFILL_33_DFFSR_133 BUFX2_37/A DFFSR_81/S FILL
XFILL_4_NAND3X1_117 INVX1_94/gnd DFFSR_25/S FILL
XFILL_9_CLKBUF1_1 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_23_DFFSR_136 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_1_DFFSR_58 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_29_DFFSR_11 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_18_DFFSR_51 INVX1_2/gnd DFFSR_51/S FILL
XFILL_13_DFFSR_139 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_3_OAI21X1_201 BUFX2_35/A DFFSR_97/S FILL
XFILL_0_OR2X2_3 BUFX2_43/A DFFSR_23/S FILL
XFILL_6_NAND2X1_153 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_3_INVX1_290 BUFX2_36/A DFFSR_8/S FILL
XFILL_20_4_0 INVX1_94/gnd DFFSR_52/S FILL
XFILL_9_DFFSR_133 BUFX2_37/A DFFSR_81/S FILL
XFILL_26_DFFSR_7 INVX1_8/gnd DFFSR_7/S FILL
XFILL_4_OAI21X1_135 BUFX2_5/gnd DFFSR_23/S FILL
XNAND2X1_189 AND2X2_8/A AND2X2_8/B BUFX2_5/gnd OAI21X1_201/C DFFSR_6/S NAND2X1
XFILL_50_DFFSR_164 INVX1_89/gnd DFFSR_2/S FILL
XFILL_18_DFFPOSX1_10 INVX1_8/gnd DFFSR_5/S FILL
XFILL_0_5_0 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_2_INVX1_110 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_40_DFFSR_167 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_9_DFFSR_65 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_30_DFFSR_170 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_15_DFFSR_98 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_37_DFFSR_18 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_26_DFFSR_58 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_20_DFFSR_173 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_16_DFFPOSX1_1 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_4_NAND2X1_249 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_10_DFFSR_176 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_2_AOI22X1_8 BUFX2_43/A DFFSR_97/S FILL
XFILL_15_DFFPOSX1_4 BUFX2_17/gnd DFFSR_7/S FILL
XINVX1_437 BUFX2_6/Y BUFX2_35/A INVX1_437/Y DFFSR_97/S INVX1
XFILL_14_DFFPOSX1_7 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_5_NOR2X1_52 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_6_XOR2X1_12 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_47_DFFSR_3 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_0_INVX1_327 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_8_DFFPOSX1_21 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_2_OAI21X1_231 BUFX2_36/A DFFSR_6/S FILL
XFILL_4_INVX1_434 INVX1_8/gnd DFFSR_5/S FILL
XFILL_6_DFFSR_170 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_45_DFFSR_25 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_5_NAND2X1_183 INVX1_8/gnd DFFSR_7/S FILL
XFILL_34_DFFSR_65 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_23_DFFSR_100 INVX1_23/gnd DFFSR_186/S FILL
XFILL_2_AND2X2_14 BUFX2_35/A DFFSR_97/S FILL
XFILL_1_DFFSR_22 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_18_DFFSR_15 INVX1_8/gnd DFFSR_7/S FILL
XFILL_13_DFFSR_103 INVX1_8/gnd DFFSR_7/S FILL
XFILL_3_INVX1_254 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_6_NAND2X1_117 BUFX2_35/A DFFSR_14/S FILL
XFILL_3_OAI21X1_165 BUFX2_35/A DFFSR_97/S FILL
XFILL_28_1_1 INVX1_89/gnd DFFSR_36/S FILL
XFILL_2_INVX1_5 INVX1_4/gnd DFFSR_51/S FILL
XFILL_0_NOR2X1_3 INVX1_94/gnd DFFSR_25/S FILL
XFILL_20_CLKBUF1_5 INVX1_89/gnd DFFSR_2/S FILL
XFILL_9_AOI21X1_42 INVX1_23/gnd DFFSR_91/S FILL
XNAND2X1_153 DFFSR_152/Q DFFSR_8/S BUFX2_5/gnd NAND2X1_153/Y DFFSR_6/S NAND2X1
XFILL_10_CLKBUF1_8 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_42_DFFSR_72 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_50_DFFSR_128 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_26_3_2 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_8_AOI21X1_45 INVX1_89/gnd DFFSR_36/S FILL
XFILL_3_NAND2X1_279 INVX1_89/gnd DFFSR_2/S FILL
XFILL_27_DFFPOSX1_29 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_8_2_1 BUFX2_43/A DFFSR_97/S FILL
XFILL_15_DFFSR_62 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_26_DFFSR_22 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_7_AOI21X1_48 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_40_DFFSR_131 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_9_DFFSR_29 INVX1_4/gnd DFFSR_4/S FILL
XFILL_30_DFFSR_134 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_6_4_2 BUFX2_35/A DFFSR_14/S FILL
XFILL_4_NAND2X1_213 BUFX2_35/A DFFSR_97/S FILL
XFILL_20_DFFSR_137 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_6_CLKBUF1_2 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_1_OAI21X1_261 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_10_DFFSR_140 DFFSR_71/gnd DFFSR_10/S FILL
XINVX1_401 INVX1_401/A BUFX2_35/A INVX1_401/Y DFFSR_14/S INVX1
XFILL_0_INVX1_291 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_3_NAND3X1_111 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_50_DFFSR_79 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_13_DFFSR_1 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_5_NOR2X1_16 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_5_NAND2X1_147 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_23_DFFSR_69 BUFX2_43/A DFFSR_23/S FILL
XFILL_2_OAI21X1_195 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_6_DFFSR_76 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_6_DFFSR_134 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_4_INVX1_398 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_34_DFFSR_29 INVX1_4/gnd DFFSR_4/S FILL
XFILL_47_DFFSR_165 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_37_DFFSR_168 BUFX2_36/A DFFSR_8/S FILL
XFILL_5_BUFX2_14 BUFX2_37/A DFFSR_81/S FILL
XFILL_27_DFFSR_171 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_17_DFFSR_174 BUFX2_43/A DFFSR_97/S FILL
XFILL_3_INVX1_218 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_3_OAI21X1_129 INVX1_4/gnd DFFSR_4/S FILL
XFILL_9_AOI22X1_6 BUFX2_37/A DFFSR_81/S FILL
XFILL_8_OAI21X1_93 INVX1_4/gnd DFFSR_51/S FILL
XFILL_31_DFFSR_76 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_3_INVX1_70 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_42_DFFSR_36 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_7_OAI21X1_96 INVX1_4/gnd DFFSR_51/S FILL
XOAI21X1_4 DFFSR_3/S INVX1_5/Y OAI21X1_4/C INVX1_4/gnd DFFSR_4/D DFFSR_51/S OAI21X1
XNAND2X1_117 BUFX2_21/Y DFFSR_109/Q BUFX2_35/A NAND2X1_117/Y DFFSR_14/S NAND2X1
XFILL_6_OAI21X1_99 BUFX2_43/A DFFSR_97/S FILL
XFILL_2_NOR2X1_53 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_3_XOR2X1_13 INVX1_8/gnd DFFSR_7/S FILL
XFILL_4_OAI21X1_1 INVX1_2/gnd DFFSR_51/S FILL
XFILL_3_NAND2X1_243 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_1_INVX1_435 INVX1_8/gnd DFFSR_5/S FILL
XOAI21X1_99 BUFX2_25/Y INVX1_112/Y NAND2X1_99/Y BUFX2_43/A DFFSR_99/D DFFSR_97/S OAI21X1
XFILL_3_DFFSR_171 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_7_AOI21X1_12 INVX1_8/gnd DFFSR_7/S FILL
XFILL_15_DFFSR_26 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_1_OAI21X1_225 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_7_DFFPOSX1_15 BUFX2_35/A DFFSR_14/S FILL
XFILL_9_AND2X2_12 BUFX2_43/A DFFSR_97/S FILL
XFILL_6_AOI21X1_15 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_20_DFFSR_101 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_4_DFFPOSX1_1 BUFX2_6/gnd DFFSR_14/S FILL
XAOI21X1_15 AOI22X1_7/C AOI22X1_7/D NAND3X1_73/B BUFX2_5/gnd AOI21X1_15/Y DFFSR_23/S
+ AOI21X1
XFILL_5_AOI21X1_18 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_4_NAND2X1_177 INVX1_89/gnd DFFSR_36/S FILL
XFILL_10_DFFSR_104 INVX1_4/gnd DFFSR_4/S FILL
XFILL_4_AOI21X1_21 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_50_DFFSR_43 INVX1_94/gnd DFFSR_25/S FILL
XFILL_3_DFFPOSX1_4 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_0_INVX1_255 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_3_AOI21X1_24 BUFX2_43/A DFFSR_97/S FILL
XFILL_39_DFFSR_83 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_2_DFFPOSX1_7 DFFSR_71/gnd DFFSR_45/S FILL
XINVX1_365 INVX1_87/A DFFSR_79/gnd INVX1_365/Y DFFSR_45/S INVX1
XFILL_2_OAI21X1_159 BUFX2_43/A DFFSR_97/S FILL
XFILL_17_CLKBUF1_6 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_2_AOI21X1_27 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_4_INVX1_362 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_1_AOI21X1_30 INVX1_23/gnd DFFSR_91/S FILL
XFILL_23_DFFSR_33 INVX1_94/gnd DFFSR_52/S FILL
XFILL_6_DFFSR_40 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_5_NAND2X1_111 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_12_DFFSR_73 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_0_AOI21X1_33 BUFX2_35/A DFFSR_14/S FILL
XFILL_47_DFFSR_129 INVX1_2/gnd DFFSR_1/S FILL
XFILL_37_DFFSR_132 INVX1_2/gnd DFFSR_51/S FILL
XBUFX2_18 INVX1_1/Y DFFSR_3/gnd BUFX2_18/Y DFFSR_65/S BUFX2
XFILL_26_DFFPOSX1_23 INVX1_23/gnd DFFSR_91/S FILL
XFILL_27_DFFSR_135 BUFX2_43/A DFFSR_97/S FILL
XFILL_3_INVX1_182 BUFX2_37/A DFFSR_8/S FILL
XFILL_2_NAND2X1_273 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_3_CLKBUF1_3 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_47_DFFSR_90 INVX1_2/gnd DFFSR_1/S FILL
XFILL_17_DFFSR_138 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_8_OAI21X1_57 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_7_OAI21X1_60 BUFX2_37/A DFFSR_81/S FILL
XFILL_6_NAND2X1_78 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_3_NAND2X1_207 BUFX2_43/A DFFSR_97/S FILL
XFILL_6_OAI21X1_63 INVX1_94/gnd DFFSR_25/S FILL
XFILL_5_NAND2X1_81 INVX1_94/gnd DFFSR_25/S FILL
XFILL_3_INVX1_34 INVX1_89/gnd DFFSR_36/S FILL
XFILL_31_DFFSR_40 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_2_NOR2X1_17 INVX1_4/gnd DFFSR_4/S FILL
XFILL_3_DFFSR_87 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_0_OAI21X1_255 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_20_DFFSR_80 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_4_NAND2X1_84 BUFX2_36/A DFFSR_6/S FILL
XFILL_5_OAI21X1_66 INVX1_4/gnd DFFSR_51/S FILL
XNAND2X1_78 BUFX2_16/Y DFFSR_70/Q DFFSR_73/gnd NAND2X1_78/Y DFFSR_11/S NAND2X1
XFILL_2_NAND3X1_105 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_3_DFFSR_135 BUFX2_43/A DFFSR_97/S FILL
XOAI21X1_63 DFFSR_25/S INVX1_71/Y OAI21X1_63/C INVX1_94/gnd DFFSR_63/D DFFSR_25/S
+ OAI21X1
XFILL_1_INVX1_399 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_2_BUFX2_25 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_4_OAI21X1_69 BUFX2_37/A DFFSR_8/S FILL
XFILL_3_NAND2X1_87 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_44_DFFSR_166 INVX1_4/gnd DFFSR_51/S FILL
XFILL_34_DFFSR_169 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_14_XOR2X1_17 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_4_NAND2X1_141 INVX1_94/gnd DFFSR_25/S FILL
XFILL_27_4_0 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_3_OAI21X1_72 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_1_OAI21X1_189 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_2_NAND2X1_90 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_24_DFFSR_172 BUFX2_37/A DFFSR_8/S FILL
XFILL_2_OAI21X1_75 INVX1_4/gnd DFFSR_4/S FILL
XFILL_1_NAND2X1_93 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_0_INVX1_219 INVX1_94/gnd DFFSR_52/S FILL
XINVX1_329 DFFSR_65/Q DFFSR_79/gnd INVX1_329/Y DFFSR_45/S INVX1
XFILL_39_DFFSR_47 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_0_INVX1_81 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_1_OAI21X1_78 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_0_NAND2X1_96 INVX1_4/gnd DFFSR_51/S FILL
XFILL_28_DFFSR_87 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_14_DFFSR_175 INVX1_23/gnd DFFSR_91/S FILL
XFILL_6_AOI22X1_7 BUFX2_43/A DFFSR_23/S FILL
XFILL_0_OAI21X1_81 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_2_OAI21X1_123 INVX1_23/gnd DFFSR_91/S FILL
XFILL_7_5_0 BUFX2_35/A DFFSR_97/S FILL
XFILL_12_DFFSR_37 INVX1_89/gnd DFFSR_2/S FILL
XFILL_4_INVX1_326 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_0_XOR2X1_14 INVX1_89/gnd DFFSR_2/S FILL
XFILL_1_OAI21X1_2 INVX1_8/gnd DFFSR_5/S FILL
XFILL_0_DFFSR_172 BUFX2_37/A DFFSR_8/S FILL
XFILL_2_NAND2X1_237 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_25_DFFSR_4 INVX1_4/gnd DFFSR_4/S FILL
XFILL_47_DFFSR_54 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_6_AND2X2_13 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_17_DFFSR_102 INVX1_8/gnd DFFSR_7/S FILL
XFILL_3_INVX1_146 INVX1_4/gnd DFFSR_4/S FILL
XFILL_36_DFFSR_94 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_8_OAI21X1_21 INVX1_2/gnd DFFSR_51/S FILL
XFILL_20_DFFSR_44 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_3_DFFSR_51 INVX1_2/gnd DFFSR_51/S FILL
XFILL_6_NAND2X1_42 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_7_OAI21X1_24 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_0_OAI21X1_219 BUFX2_35/A DFFSR_97/S FILL
XFILL_3_NAND2X1_171 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_5_NAND2X1_45 INVX1_89/gnd DFFSR_36/S FILL
XFILL_6_OAI21X1_27 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_14_CLKBUF1_7 BUFX2_43/A DFFSR_97/S FILL
XFILL_1_INVX1_363 INVX1_94/gnd DFFSR_25/S FILL
XFILL_5_OAI21X1_30 INVX1_89/gnd DFFSR_36/S FILL
XNAND2X1_42 DFFSR_51/S INVX1_39/A DFFSR_3/gnd OAI21X1_42/C DFFSR_4/S NAND2X1
XFILL_4_NAND2X1_48 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_4_OAI21X1_33 BUFX2_19/gnd DFFSR_52/S FILL
XOAI21X1_27 DFFSR_1/S INVX1_31/Y OAI21X1_27/C DFFSR_1/gnd DFFSR_27/D DFFSR_1/S OAI21X1
XFILL_3_NAND2X1_51 INVX1_2/gnd DFFSR_51/S FILL
XFILL_1_OAI21X1_153 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_2_NAND2X1_54 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_3_OAI21X1_36 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_44_DFFSR_130 INVX1_4/gnd DFFSR_51/S FILL
XFILL_15_DFFPOSX1_28 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_4_NAND2X1_105 BUFX2_35/A DFFSR_14/S FILL
XFILL_34_DFFSR_133 BUFX2_37/A DFFSR_81/S FILL
XFILL_2_OAI21X1_39 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_1_NAND2X1_57 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_0_INVX1_183 BUFX2_37/A DFFSR_8/S FILL
XFILL_0_NAND2X1_60 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_24_DFFSR_136 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_0_INVX1_45 INVX1_8/gnd DFFSR_5/S FILL
XFILL_35_1_1 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_1_OAI21X1_42 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_39_DFFSR_11 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_17_DFFSR_91 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_19_5 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_0_CLKBUF1_4 BUFX2_8/gnd DFFSR_10/S FILL
XINVX1_293 INVX1_41/A DFFSR_71/gnd INVX1_293/Y DFFSR_45/S INVX1
XFILL_0_OAI21X1_45 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_0_DFFSR_98 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_28_DFFSR_51 INVX1_2/gnd DFFSR_51/S FILL
XFILL_14_DFFSR_139 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_4_INVX1_290 BUFX2_36/A DFFSR_8/S FILL
XFILL_33_3_2 INVX1_8/gnd DFFSR_7/S FILL
XFILL_1_NAND2X1_267 INVX1_4/gnd DFFSR_4/S FILL
XFILL_9_AOI22X1_11 INVX1_23/gnd DFFSR_91/S FILL
XFILL_25_DFFPOSX1_17 BUFX2_37/A DFFSR_8/S FILL
XFILL_8_AOI22X1_14 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_1_INVX1_2 INVX1_2/gnd DFFSR_51/S FILL
XFILL_51_DFFSR_164 INVX1_89/gnd DFFSR_2/S FILL
XFILL_0_DFFSR_136 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_2_NAND2X1_201 BUFX2_35/A DFFSR_14/S FILL
XFILL_3_INVX1_110 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_41_DFFSR_167 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_31_DFFSR_170 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_25_DFFSR_98 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_47_DFFSR_18 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_36_DFFSR_58 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_21_DFFSR_173 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_3_NAND2X1_135 BUFX2_36/A DFFSR_6/S FILL
XFILL_3_DFFSR_15 INVX1_8/gnd DFFSR_7/S FILL
XFILL_0_OAI21X1_183 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_3_AOI22X1_8 BUFX2_43/A DFFSR_97/S FILL
XFILL_4_NAND2X1_12 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_11_DFFSR_176 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_11_OAI22X1_53 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_6_NOR2X1_52 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_7_XOR2X1_12 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_1_INVX1_327 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_10_OAI22X1_56 BUFX2_37/A DFFSR_8/S FILL
XFILL_3_NAND2X1_15 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_1_OAI21X1_117 BUFX2_35/A DFFSR_97/S FILL
XFILL_7_DFFSR_170 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_2_NAND2X1_18 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_44_DFFSR_65 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_24_DFFSR_100 INVX1_23/gnd DFFSR_186/S FILL
XFILL_8_NAND3X1_77 BUFX2_37/A DFFSR_81/S FILL
XFILL_1_NAND2X1_21 INVX1_4/gnd DFFSR_4/S FILL
XFILL_3_AND2X2_14 BUFX2_35/A DFFSR_97/S FILL
XINVX1_257 XNOR2X1_2/Y BUFX2_36/A INVX1_257/Y DFFSR_8/S INVX1
XFILL_0_DFFSR_62 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_17_DFFSR_55 INVX1_89/gnd DFFSR_36/S FILL
XFILL_28_DFFSR_15 INVX1_8/gnd DFFSR_7/S FILL
XFILL_9_OAI22X1_59 INVX1_8/gnd DFFSR_7/S FILL
XFILL_14_DFFSR_103 INVX1_8/gnd DFFSR_7/S FILL
XFILL_0_NAND2X1_24 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_0_INVX1_147 INVX1_4/gnd DFFSR_4/S FILL
XFILL_1_NAND2X1_231 BUFX2_37/A DFFSR_81/S FILL
XFILL_7_NAND3X1_80 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_8_OAI22X1_62 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_4_INVX1_254 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_6_NAND3X1_83 BUFX2_37/A DFFSR_81/S FILL
XFILL_7_OAI22X1_65 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_0_NAND3X1_129 BUFX2_35/A DFFSR_14/S FILL
XNAND3X1_83 NAND3X1_83/A NAND3X1_83/B NAND3X1_79/Y BUFX2_37/A NAND3X1_83/Y DFFSR_81/S
+ NAND3X1
XFILL_5_NAND3X1_86 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_6_OAI22X1_68 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_4_NAND3X1_89 BUFX2_43/A DFFSR_23/S FILL
XFILL_11_CLKBUF1_8 BUFX2_5/gnd DFFSR_6/S FILL
XOAI22X1_68 INVX1_394/Y OAI22X1_40/B INVX1_395/Y OAI22X1_52/D DFFSR_5/gnd NOR2X1_43/B
+ DFFSR_5/S OAI22X1
XFILL_0_DFFSR_100 INVX1_23/gnd DFFSR_186/S FILL
XFILL_3_NAND3X1_92 BUFX2_43/A DFFSR_23/S FILL
XFILL_51_DFFSR_128 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_2_NAND2X1_165 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_2_NAND3X1_95 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_8_DFFSR_69 BUFX2_43/A DFFSR_23/S FILL
XFILL_25_DFFSR_62 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_36_DFFSR_22 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_41_DFFSR_131 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_1_NAND3X1_98 BUFX2_35/A DFFSR_14/S FILL
XFILL_31_DFFSR_134 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_21_DFFSR_137 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_7_CLKBUF1_2 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_14_DFFPOSX1_22 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_0_OAI21X1_147 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_11_DFFSR_140 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_1_INVX1_291 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_6_NOR2X1_16 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_37_DFFSR_7 INVX1_8/gnd DFFSR_7/S FILL
XFILL_41_5 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_33_DFFSR_69 BUFX2_43/A DFFSR_23/S FILL
XFILL_10_OAI22X1_20 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_0_NAND2X1_261 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_7_DFFSR_134 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_44_DFFSR_29 INVX1_4/gnd DFFSR_4/S FILL
XFILL_48_DFFSR_165 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_24_DFFPOSX1_11 INVX1_4/gnd DFFSR_4/S FILL
XFILL_8_NAND3X1_41 BUFX2_43/A DFFSR_23/S FILL
XFILL_38_DFFSR_168 BUFX2_36/A DFFSR_8/S FILL
XFILL_9_OAI22X1_23 INVX1_89/gnd DFFSR_2/S FILL
XFILL_0_INVX1_111 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_0_DFFSR_26 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_7_NAND3X1_44 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_28_DFFSR_171 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_8_OAI22X1_26 INVX1_94/gnd DFFSR_52/S FILL
XINVX1_221 INVX1_221/A BUFX2_17/gnd AND2X2_3/B DFFSR_7/S INVX1
XFILL_17_DFFSR_19 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_6_NAND3X1_47 BUFX2_43/A DFFSR_97/S FILL
XFILL_1_NAND2X1_195 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_7_OAI22X1_29 INVX1_8/gnd DFFSR_5/S FILL
XFILL_18_DFFSR_174 BUFX2_43/A DFFSR_97/S FILL
XFILL_5_NAND3X1_50 BUFX2_37/A DFFSR_81/S FILL
XFILL_6_OAI22X1_32 DFFSR_71/gnd DFFSR_10/S FILL
XXOR2X1_16 INVX1_153/A DFFSR_144/Q INVX1_8/gnd XOR2X1_16/Y DFFSR_5/S XOR2X1
XNAND3X1_47 OAI22X1_2/Y NAND3X1_47/B NAND3X1_37/Y BUFX2_43/A AOI22X1_8/C DFFSR_97/S
+ NAND3X1
XFILL_0_AOI22X1_9 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_4_NAND3X1_53 BUFX2_37/A DFFSR_81/S FILL
XFILL_41_DFFSR_76 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_5_OAI22X1_35 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_3_NAND3X1_56 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_4_OAI22X1_38 BUFX2_19/gnd DFFSR_52/S FILL
XOAI22X1_32 INVX1_319/Y OAI22X1_8/B INVX1_320/Y OAI22X1_8/D DFFSR_71/gnd NOR2X1_25/A
+ DFFSR_10/S OAI22X1
XFILL_3_NOR2X1_53 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_4_XOR2X1_13 INVX1_8/gnd DFFSR_7/S FILL
XFILL_5_OAI21X1_1 INVX1_2/gnd DFFSR_51/S FILL
XFILL_8_OAI21X1_232 BUFX2_35/A DFFSR_97/S FILL
XDFFSR_174 AND2X2_11/B CLKBUF1_14/Y DFFSR_175/R DFFSR_97/S DFFSR_174/D BUFX2_43/A
+ DFFSR_97/S DFFSR
XFILL_2_NAND3X1_59 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_2_INVX1_435 INVX1_8/gnd DFFSR_5/S FILL
XFILL_34_4_0 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_2_NAND2X1_129 INVX1_4/gnd DFFSR_4/S FILL
XFILL_3_OAI22X1_41 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_1_NAND3X1_62 BUFX2_43/A DFFSR_23/S FILL
XFILL_4_DFFSR_171 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_8_DFFSR_33 INVX1_94/gnd DFFSR_52/S FILL
XFILL_25_DFFSR_26 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_14_DFFSR_66 INVX1_2/gnd DFFSR_51/S FILL
XFILL_2_OAI22X1_44 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_21_DFFSR_101 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_0_NAND3X1_65 BUFX2_35/A DFFSR_14/S FILL
XFILL_1_OAI22X1_47 BUFX2_37/A DFFSR_8/S FILL
XFILL_0_OAI21X1_111 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_0_AND2X2_15 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_0_OAI22X1_50 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_1_XOR2X1_3 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_11_DFFSR_104 INVX1_4/gnd DFFSR_4/S FILL
XFILL_1_INVX1_255 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_49_DFFSR_83 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_18_CLKBUF1_6 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_0_NAND2X1_225 BUFX2_36/A DFFSR_8/S FILL
XFILL_33_DFFSR_33 INVX1_94/gnd DFFSR_52/S FILL
XINVX1_67 INVX1_67/A INVX1_4/gnd INVX1_67/Y DFFSR_51/S INVX1
XFILL_5_DFFSR_80 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_22_DFFSR_73 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_48_DFFSR_129 INVX1_2/gnd DFFSR_1/S FILL
XCLKBUF1_6 DFFSR_149/Q BUFX2_5/gnd CLKBUF1_6/Y DFFSR_23/S CLKBUF1
XINVX1_185 BUFX2_9/Y BUFX2_19/gnd DFFSR_155/R DFFSR_52/S INVX1
XFILL_38_DFFSR_132 INVX1_2/gnd DFFSR_51/S FILL
XFILL_1_NAND2X1_159 BUFX2_43/A DFFSR_97/S FILL
XFILL_28_DFFSR_135 BUFX2_43/A DFFSR_97/S FILL
XFILL_4_INVX1_182 BUFX2_37/A DFFSR_8/S FILL
XFILL_7_OAI21X1_262 INVX1_89/gnd DFFSR_36/S FILL
XFILL_4_BUFX2_18 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_6_NAND3X1_11 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_4_CLKBUF1_3 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_18_DFFSR_138 DFFSR_73/gnd DFFSR_11/S FILL
XNAND3X1_11 AOI22X1_3/D NAND3X1_8/B NAND3X1_8/C BUFX2_19/gnd AOI21X1_8/B DFFSR_54/S
+ NAND3X1
XFILL_5_NAND3X1_14 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_24_DFFSR_1 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_13_DFFPOSX1_16 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_4_NAND3X1_17 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_41_DFFSR_40 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_3_NOR2X1_17 INVX1_4/gnd DFFSR_4/S FILL
XFILL_2_INVX1_74 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_30_DFFSR_80 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_3_NAND3X1_20 BUFX2_37/A DFFSR_8/S FILL
XFILL_8_OAI21X1_196 INVX1_94/gnd DFFSR_25/S FILL
XDFFSR_138 INVX1_156/A CLKBUF1_13/Y DFFSR_137/R DFFSR_11/S DFFSR_138/D DFFSR_73/gnd
+ DFFSR_11/S DFFSR
XFILL_4_DFFSR_135 BUFX2_43/A DFFSR_97/S FILL
XFILL_2_NAND3X1_23 BUFX2_37/A DFFSR_81/S FILL
XFILL_14_DFFSR_30 INVX1_89/gnd DFFSR_36/S FILL
XFILL_2_INVX1_399 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_42_1_1 INVX1_4/gnd DFFSR_4/S FILL
XFILL_1_NAND3X1_26 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_45_DFFSR_166 INVX1_4/gnd DFFSR_51/S FILL
XFILL_35_DFFSR_169 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_0_NAND3X1_29 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_15_XOR2X1_17 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_1_OAI22X1_11 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_40_3_2 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_25_DFFSR_172 BUFX2_37/A DFFSR_8/S FILL
XFILL_9_OAI21X1_130 INVX1_4/gnd DFFSR_4/S FILL
XFILL_0_OAI22X1_14 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_1_INVX1_219 INVX1_94/gnd DFFSR_52/S FILL
XFILL_49_DFFSR_47 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_38_DFFSR_87 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_15_DFFSR_175 INVX1_23/gnd DFFSR_91/S FILL
XFILL_7_AOI22X1_7 BUFX2_43/A DFFSR_23/S FILL
XDFFSR_84 DFFSR_84/Q CLKBUF1_6/Y DFFSR_84/R DFFSR_97/S DFFSR_84/D BUFX2_43/A DFFSR_23/S
+ DFFSR
XFILL_0_NAND2X1_189 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_5_DFFSR_44 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_3_DFFPOSX1_27 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_22_DFFSR_37 INVX1_89/gnd DFFSR_2/S FILL
XFILL_11_DFFSR_77 INVX1_89/gnd DFFSR_2/S FILL
XINVX1_31 INVX1_31/A INVX1_2/gnd INVX1_31/Y DFFSR_1/S INVX1
XFILL_1_XOR2X1_14 INVX1_89/gnd DFFSR_2/S FILL
XFILL_2_OAI21X1_2 INVX1_8/gnd DFFSR_5/S FILL
XFILL_0_NOR2X1_54 DFFSR_1/gnd DFFSR_9/S FILL
XINVX1_149 XOR2X1_13/A INVX1_4/gnd INVX1_149/Y DFFSR_51/S INVX1
XFILL_1_1 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_1_DFFSR_172 BUFX2_37/A DFFSR_8/S FILL
XFILL_15_XOR2X1_7 INVX1_23/gnd DFFSR_91/S FILL
XFILL_7_OAI21X1_226 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_1_NAND2X1_123 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_7_AND2X2_13 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_18_DFFSR_102 INVX1_8/gnd DFFSR_7/S FILL
XFILL_46_DFFSR_94 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_2_DFFSR_91 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_2_INVX1_38 INVX1_94/gnd DFFSR_52/S FILL
XFILL_7_AND2X2_3 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_19_DFFSR_84 BUFX2_43/A DFFSR_23/S FILL
XFILL_30_DFFSR_44 BUFX2_8/gnd DFFSR_10/S FILL
XDFFSR_102 INVX1_376/A CLKBUF1_3/Y DFFSR_97/R DFFSR_7/S DFFSR_102/D INVX1_8/gnd DFFSR_7/S
+ DFFSR
XFILL_2_INVX1_363 INVX1_94/gnd DFFSR_25/S FILL
XFILL_8_OAI21X1_160 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_15_CLKBUF1_7 BUFX2_43/A DFFSR_97/S FILL
XFILL_1_BUFX2_29 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_45_DFFSR_130 INVX1_4/gnd DFFSR_51/S FILL
XFILL_35_DFFSR_133 BUFX2_37/A DFFSR_81/S FILL
XFILL_25_DFFSR_136 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_27_DFFSR_91 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_1_INVX1_183 BUFX2_37/A DFFSR_8/S FILL
XFILL_23_2 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_1_CLKBUF1_4 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_38_DFFSR_51 INVX1_2/gnd DFFSR_51/S FILL
XFILL_15_DFFSR_139 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_49_DFFSR_11 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_0_NAND2X1_153 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_0_NOR2X1_18 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_11_DFFSR_41 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_6_OAI21X1_256 INVX1_2/gnd DFFSR_51/S FILL
XDFFSR_48 INVX1_54/A DFFSR_24/CLK DFFSR_46/R DFFSR_4/S DFFSR_48/D INVX1_4/gnd DFFSR_4/S
+ DFFSR
XINVX1_113 DFFSR_100/Q INVX1_23/gnd INVX1_113/Y DFFSR_91/S INVX1
XFILL_8_NAND3X1_106 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_7_OAI21X1_190 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_15_DFFSR_8 BUFX2_36/A DFFSR_8/S FILL
XFILL_42_DFFSR_167 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_1_DFFSR_136 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_12_DFFPOSX1_10 INVX1_8/gnd DFFSR_5/S FILL
XFILL_32_DFFSR_170 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_35_DFFSR_98 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_46_DFFSR_58 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_14_1_2 BUFX2_37/A DFFSR_8/S FILL
XFILL_22_DFFSR_173 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_2_DFFSR_55 INVX1_89/gnd DFFSR_36/S FILL
XFILL_19_DFFSR_48 INVX1_4/gnd DFFSR_4/S FILL
XFILL_4_AOI22X1_8 BUFX2_43/A DFFSR_97/S FILL
XFILL_8_OAI21X1_124 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_12_DFFSR_176 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_8_XOR2X1_12 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_2_INVX1_327 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_2_DFFPOSX1_21 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_8_DFFSR_170 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_36_DFFSR_4 INVX1_4/gnd DFFSR_4/S FILL
XFILL_25_DFFSR_100 INVX1_23/gnd DFFSR_186/S FILL
XAND2X2_17 AND2X2_17/A AND2X2_17/B DFFSR_5/gnd AND2X2_17/Y DFFSR_5/S AND2X2
XFILL_4_AND2X2_14 BUFX2_35/A DFFSR_97/S FILL
XFILL_16_DFFSR_95 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_27_DFFSR_55 INVX1_89/gnd DFFSR_36/S FILL
XFILL_38_DFFSR_15 INVX1_8/gnd DFFSR_7/S FILL
XFILL_1_INVX1_147 INVX1_4/gnd DFFSR_4/S FILL
XFILL_15_DFFSR_103 INVX1_8/gnd DFFSR_7/S FILL
XDFFSR_12 DFFSR_12/Q DFFSR_20/CLK DFFSR_9/R DFFSR_12/S DFFSR_12/D BUFX2_6/gnd DFFSR_14/S
+ DFFSR
XFILL_0_NAND2X1_117 BUFX2_35/A DFFSR_14/S FILL
XFILL_6_OAI21X1_220 BUFX2_43/A DFFSR_97/S FILL
XFILL_41_4_0 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_1_DFFSR_100 INVX1_23/gnd DFFSR_186/S FILL
XFILL_12_CLKBUF1_8 BUFX2_5/gnd DFFSR_6/S FILL
XOAI21X1_256 DFFSR_1/S INVX1_419/Y NAND2X1_267/Y INVX1_2/gnd DFFSR_188/D DFFSR_51/S
+ OAI21X1
XFILL_7_OAI21X1_154 BUFX2_37/A DFFSR_8/S FILL
XFILL_35_DFFSR_62 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_46_DFFSR_22 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_42_DFFSR_131 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_21_DFFPOSX1_29 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_32_DFFSR_134 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_22_DFFSR_137 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_8_CLKBUF1_2 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_2_DFFSR_19 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_19_DFFSR_12 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_12_DFFSR_140 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_2_INVX1_291 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_45_2 INVX1_2/gnd DFFSR_51/S FILL
XFILL_43_DFFSR_69 BUFX2_43/A DFFSR_23/S FILL
XFILL_49_DFFSR_165 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_8_DFFSR_134 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_5_OAI21X1_250 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_39_DFFSR_168 BUFX2_36/A DFFSR_8/S FILL
XFILL_17_CLKBUF1_11 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_7_NAND3X1_100 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_16_CLKBUF1_14 BUFX2_43/A DFFSR_23/S FILL
XFILL_29_DFFSR_171 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_27_DFFSR_19 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_1_INVX1_111 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_16_DFFSR_59 INVX1_4/gnd DFFSR_51/S FILL
XFILL_19_DFFSR_174 BUFX2_43/A DFFSR_97/S FILL
XFILL_6_OAI21X1_184 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_15_CLKBUF1_17 INVX1_94/gnd DFFSR_25/S FILL
XFILL_1_AOI22X1_9 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_3_DFFSR_7 INVX1_8/gnd DFFSR_7/S FILL
XFILL_14_CLKBUF1_20 INVX1_4/gnd DFFSR_51/S FILL
XOAI21X1_220 INVX1_241/A AND2X2_12/Y NAND3X1_37/C BUFX2_43/A NAND3X1_67/C DFFSR_97/S
+ OAI21X1
XFILL_4_NOR2X1_53 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_13_CLKBUF1_23 INVX1_89/gnd DFFSR_2/S FILL
XFILL_5_XOR2X1_13 INVX1_8/gnd DFFSR_7/S FILL
XFILL_47_3_2 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_6_OAI21X1_1 INVX1_2/gnd DFFSR_51/S FILL
XFILL_3_INVX1_435 INVX1_8/gnd DFFSR_5/S FILL
XFILL_7_OAI21X1_118 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_5_DFFSR_171 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_35_DFFSR_26 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_24_DFFSR_66 INVX1_2/gnd DFFSR_51/S FILL
XFILL_7_DFFSR_73 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_22_DFFSR_101 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_1_DFFPOSX1_15 BUFX2_35/A DFFSR_14/S FILL
XFILL_1_AND2X2_15 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_6_BUFX2_11 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_12_DFFSR_104 INVX1_4/gnd DFFSR_4/S FILL
XFILL_2_INVX1_255 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_15_2_0 BUFX2_37/A DFFSR_81/S FILL
XFILL_6_NAND3X1_130 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_5_OAI21X1_214 BUFX2_35/A DFFSR_97/S FILL
XFILL_19_CLKBUF1_6 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_43_DFFSR_33 INVX1_94/gnd DFFSR_52/S FILL
XFILL_32_DFFSR_73 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_13_4_1 BUFX2_36/A DFFSR_8/S FILL
XFILL_49_DFFSR_129 INVX1_2/gnd DFFSR_1/S FILL
XFILL_16_DFFSR_23 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_39_DFFSR_132 INVX1_2/gnd DFFSR_51/S FILL
XFILL_29_DFFSR_135 BUFX2_43/A DFFSR_97/S FILL
XFILL_6_OAI21X1_148 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_20_DFFPOSX1_23 INVX1_23/gnd DFFSR_91/S FILL
XFILL_5_CLKBUF1_3 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_19_DFFSR_138 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_48_DFFSR_7 INVX1_8/gnd DFFSR_7/S FILL
XNOR2X1_20 NOR2X1_20/A NOR2X1_20/B BUFX2_16/gnd NOR2X1_20/Y DFFSR_11/S NOR2X1
XFILL_4_NOR2X1_17 INVX1_4/gnd DFFSR_4/S FILL
XFILL_40_DFFSR_80 BUFX2_16/gnd DFFSR_65/S FILL
XOAI21X1_184 INVX1_219/A AOI22X1_1/Y NAND3X1_3/Y BUFX2_19/gnd AOI21X1_6/C DFFSR_52/S
+ OAI21X1
XFILL_6_NAND2X1_262 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_24_DFFSR_30 INVX1_89/gnd DFFSR_36/S FILL
XFILL_7_DFFSR_37 INVX1_89/gnd DFFSR_2/S FILL
XFILL_3_INVX1_399 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_13_DFFSR_70 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_5_DFFSR_135 BUFX2_43/A DFFSR_97/S FILL
XFILL_46_DFFSR_166 INVX1_4/gnd DFFSR_51/S FILL
XFILL_36_DFFSR_169 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_3_INVX1_9 BUFX2_36/A DFFSR_6/S FILL
XFILL_4_OAI21X1_244 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_0_XOR2X1_7 INVX1_23/gnd DFFSR_91/S FILL
XFILL_26_DFFSR_172 BUFX2_37/A DFFSR_8/S FILL
XFILL_2_INVX1_219 INVX1_94/gnd DFFSR_52/S FILL
XFILL_48_DFFSR_87 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_16_DFFSR_175 INVX1_23/gnd DFFSR_91/S FILL
XFILL_8_AOI22X1_7 BUFX2_43/A DFFSR_23/S FILL
XFILL_4_DFFSR_84 BUFX2_43/A DFFSR_23/S FILL
XFILL_32_DFFSR_37 INVX1_89/gnd DFFSR_2/S FILL
XFILL_4_INVX1_31 INVX1_2/gnd DFFSR_1/S FILL
XFILL_5_OAI21X1_178 INVX1_94/gnd DFFSR_25/S FILL
XFILL_2_XOR2X1_14 INVX1_89/gnd DFFSR_2/S FILL
XFILL_21_DFFSR_77 INVX1_89/gnd DFFSR_2/S FILL
XFILL_3_OAI21X1_2 INVX1_8/gnd DFFSR_5/S FILL
XFILL_1_NOR2X1_54 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_5_CLKBUF1_11 BUFX2_7/gnd DFFSR_54/S FILL
XNAND3X1_130 NOR2X1_1/B NOR2X1_1/A INVX1_404/Y BUFX2_19/gnd NAND3X1_130/Y DFFSR_52/S
+ NAND3X1
XFILL_21_1_2 INVX1_94/gnd DFFSR_25/S FILL
XFILL_0_INVX1_436 INVX1_89/gnd DFFSR_36/S FILL
XFILL_4_CLKBUF1_14 BUFX2_43/A DFFSR_23/S FILL
XFILL_2_DFFSR_172 BUFX2_37/A DFFSR_8/S FILL
XFILL_3_BUFX2_22 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_3_0_1 INVX1_23/gnd DFFSR_91/S FILL
XFILL_8_AND2X2_13 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_3_CLKBUF1_17 INVX1_94/gnd DFFSR_25/S FILL
XFILL_13_NOR3X1_1 INVX1_94/gnd DFFSR_52/S FILL
XFILL_14_DFFSR_5 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_19_DFFSR_102 INVX1_8/gnd DFFSR_7/S FILL
XFILL_2_CLKBUF1_20 INVX1_4/gnd DFFSR_51/S FILL
XFILL_6_OAI21X1_112 INVX1_4/gnd DFFSR_4/S FILL
XFILL_1_2_2 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_1_CLKBUF1_23 INVX1_89/gnd DFFSR_2/S FILL
XOAI21X1_148 OAI21X1_148/A INVX1_170/Y NAND2X1_148/Y DFFSR_89/gnd DFFSR_148/D DFFSR_186/S
+ OAI21X1
XFILL_29_DFFSR_84 BUFX2_43/A DFFSR_23/S FILL
XFILL_1_INVX1_78 BUFX2_36/A DFFSR_8/S FILL
XFILL_40_DFFSR_44 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_6_NAND2X1_226 BUFX2_36/A DFFSR_6/S FILL
XFILL_3_INVX1_363 INVX1_94/gnd DFFSR_25/S FILL
XFILL_16_CLKBUF1_7 BUFX2_43/A DFFSR_97/S FILL
XFILL_13_DFFSR_34 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_5_NAND3X1_124 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_46_DFFSR_130 INVX1_4/gnd DFFSR_51/S FILL
XNAND2X1_262 DFFSR_186/S din[7] DFFSR_89/gnd NAND2X1_262/Y DFFSR_92/S NAND2X1
XFILL_36_DFFSR_133 BUFX2_37/A DFFSR_81/S FILL
XFILL_48_4_0 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_10_4 BUFX2_43/A DFFSR_23/S FILL
XFILL_4_OAI21X1_208 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_26_DFFSR_136 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_35_DFFSR_1 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_37_DFFSR_91 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_2_INVX1_183 BUFX2_37/A DFFSR_8/S FILL
XFILL_2_CLKBUF1_4 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_48_DFFSR_51 INVX1_2/gnd DFFSR_51/S FILL
XFILL_16_DFFSR_139 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_19_DFFPOSX1_17 BUFX2_37/A DFFSR_8/S FILL
XFILL_10_DFFSR_81 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_5_OAI21X1_142 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_1_NOR2X1_18 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_21_DFFSR_41 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_4_DFFSR_48 INVX1_4/gnd DFFSR_4/S FILL
XFILL_0_INVX1_400 BUFX2_35/A DFFSR_97/S FILL
XFILL_43_DFFSR_167 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_2_DFFSR_136 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_27_DFFPOSX1_5 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_33_DFFSR_170 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_26_DFFPOSX1_8 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_5_NAND2X1_256 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_45_DFFSR_98 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_23_DFFSR_173 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_6_AND2X2_7 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_1_DFFSR_95 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_1_INVX1_42 INVX1_89/gnd DFFSR_36/S FILL
XFILL_29_DFFSR_48 INVX1_4/gnd DFFSR_4/S FILL
XFILL_18_DFFSR_88 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_5_AOI22X1_8 BUFX2_43/A DFFSR_97/S FILL
XFILL_3_OAI21X1_238 BUFX2_19/gnd DFFSR_52/S FILL
XOAI21X1_112 BUFX2_15/Y INVX1_126/Y OAI21X1_112/C INVX1_4/gnd DFFSR_112/D DFFSR_4/S
+ OAI21X1
XFILL_9_DFFPOSX1_28 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_13_DFFSR_176 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_6_NAND2X1_190 BUFX2_35/A DFFSR_97/S FILL
XFILL_9_XOR2X1_12 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_3_INVX1_327 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_0_BUFX2_33 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_0_OAI21X1_3 INVX1_4/gnd DFFSR_51/S FILL
XNAND2X1_226 NOR2X1_10/Y XNOR2X1_2/Y BUFX2_36/A NAND3X1_90/B DFFSR_6/S NAND2X1
XFILL_9_DFFSR_170 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_26_DFFSR_100 INVX1_23/gnd DFFSR_186/S FILL
XFILL_4_OAI21X1_172 BUFX2_36/A DFFSR_6/S FILL
XFILL_5_AND2X2_14 BUFX2_35/A DFFSR_97/S FILL
XFILL_26_DFFSR_95 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_37_DFFSR_55 INVX1_89/gnd DFFSR_36/S FILL
XFILL_48_DFFSR_15 INVX1_8/gnd DFFSR_7/S FILL
XFILL_2_INVX1_147 INVX1_4/gnd DFFSR_4/S FILL
XFILL_16_DFFSR_103 INVX1_8/gnd DFFSR_7/S FILL
XFILL_4_DFFSR_12 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_4_NAND2X1_286 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_10_DFFSR_45 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_5_OAI21X1_106 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_0_INVX1_364 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_2_DFFSR_100 INVX1_23/gnd DFFSR_186/S FILL
XFILL_13_CLKBUF1_8 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_2_DFFSR_4 INVX1_4/gnd DFFSR_4/S FILL
XFILL_5_NAND2X1_220 BUFX2_35/A DFFSR_14/S FILL
XFILL_45_DFFSR_62 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_43_DFFSR_131 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_33_DFFSR_134 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_23_DFFSR_137 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_22_2_0 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_4_NAND3X1_118 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_9_CLKBUF1_2 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_29_DFFSR_12 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_18_DFFSR_52 INVX1_94/gnd DFFSR_52/S FILL
XFILL_13_DFFSR_140 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_1_DFFSR_59 INVX1_4/gnd DFFSR_51/S FILL
XFILL_3_OAI21X1_202 BUFX2_35/A DFFSR_14/S FILL
XFILL_6_NAND2X1_154 BUFX2_37/A DFFSR_8/S FILL
XFILL_20_4_1 INVX1_94/gnd DFFSR_52/S FILL
XFILL_3_INVX1_291 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_2_3_0 INVX1_23/gnd DFFSR_186/S FILL
XFILL_26_DFFSR_8 BUFX2_36/A DFFSR_8/S FILL
XFILL_50_DFFSR_165 BUFX2_6/gnd DFFSR_14/S FILL
XNAND2X1_190 AND2X2_8/A AND2X2_9/B BUFX2_35/A NAND2X1_190/Y DFFSR_97/S NAND2X1
XFILL_9_DFFSR_134 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_4_OAI21X1_136 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_18_DFFPOSX1_11 INVX1_4/gnd DFFSR_4/S FILL
XFILL_0_5_1 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_40_DFFSR_168 BUFX2_36/A DFFSR_8/S FILL
XFILL_15_DFFSR_99 BUFX2_35/A DFFSR_97/S FILL
XFILL_37_DFFSR_19 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_2_INVX1_111 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_9_DFFSR_66 INVX1_2/gnd DFFSR_51/S FILL
XFILL_26_DFFSR_59 INVX1_4/gnd DFFSR_51/S FILL
XFILL_30_DFFSR_171 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_20_DFFSR_174 BUFX2_43/A DFFSR_97/S FILL
XFILL_16_DFFPOSX1_2 INVX1_89/gnd DFFSR_36/S FILL
XFILL_4_NAND2X1_250 INVX1_8/gnd DFFSR_5/S FILL
XFILL_2_AOI22X1_9 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_10_DFFSR_177 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_15_DFFPOSX1_5 DFFSR_73/gnd DFFSR_11/S FILL
XINVX1_438 NOR2X1_2/A DFFSR_71/gnd INVX1_438/Y DFFSR_10/S INVX1
XFILL_5_NOR2X1_53 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_14_DFFPOSX1_8 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_0_INVX1_328 INVX1_8/gnd DFFSR_7/S FILL
XFILL_6_XOR2X1_13 INVX1_8/gnd DFFSR_7/S FILL
XFILL_7_OAI21X1_1 INVX1_2/gnd DFFSR_51/S FILL
XFILL_47_DFFSR_4 INVX1_4/gnd DFFSR_4/S FILL
XFILL_2_OAI21X1_232 BUFX2_35/A DFFSR_97/S FILL
XFILL_4_INVX1_435 INVX1_8/gnd DFFSR_5/S FILL
XFILL_8_DFFPOSX1_22 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_5_NAND2X1_184 BUFX2_37/A DFFSR_8/S FILL
XFILL_6_DFFSR_171 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_45_DFFSR_26 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_34_DFFSR_66 INVX1_2/gnd DFFSR_51/S FILL
XFILL_1_DFFSR_23 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_18_DFFSR_16 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_2_AND2X2_15 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_23_DFFSR_101 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_13_DFFSR_104 INVX1_4/gnd DFFSR_4/S FILL
XFILL_3_OAI21X1_166 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_3_INVX1_255 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_28_1_2 INVX1_89/gnd DFFSR_36/S FILL
XFILL_2_INVX1_6 INVX1_8/gnd DFFSR_5/S FILL
XFILL_6_NAND2X1_118 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_0_NOR2X1_4 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_20_CLKBUF1_6 BUFX2_5/gnd DFFSR_23/S FILL
XNAND2X1_154 DFFSR_153/Q DFFSR_8/S BUFX2_37/A OAI21X1_154/C DFFSR_8/S NAND2X1
XFILL_42_DFFSR_73 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_4_OAI21X1_100 INVX1_23/gnd DFFSR_91/S FILL
XFILL_27_DFFPOSX1_30 BUFX2_43/A DFFSR_97/S FILL
XFILL_3_NAND2X1_280 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_8_AOI21X1_46 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_10_CLKBUF1_9 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_50_DFFSR_129 INVX1_2/gnd DFFSR_1/S FILL
XFILL_8_2_2 BUFX2_43/A DFFSR_97/S FILL
XFILL_26_DFFSR_23 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_15_DFFSR_63 INVX1_94/gnd DFFSR_52/S FILL
XFILL_9_DFFSR_30 INVX1_89/gnd DFFSR_36/S FILL
XFILL_40_DFFSR_132 INVX1_2/gnd DFFSR_51/S FILL
XFILL_30_DFFSR_135 BUFX2_43/A DFFSR_97/S FILL
XFILL_4_NAND2X1_214 BUFX2_35/A DFFSR_97/S FILL
XFILL_6_CLKBUF1_3 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_1_OAI21X1_262 INVX1_89/gnd DFFSR_36/S FILL
XFILL_20_DFFSR_138 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_10_DFFSR_141 INVX1_94/gnd DFFSR_25/S FILL
XINVX1_402 INVX1_402/A BUFX2_6/gnd INVX1_402/Y DFFSR_14/S INVX1
XFILL_0_INVX1_292 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_3_NAND3X1_112 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_13_DFFSR_2 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_5_NOR2X1_17 INVX1_4/gnd DFFSR_4/S FILL
XFILL_50_DFFSR_80 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_5_NAND2X1_148 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_2_OAI21X1_196 INVX1_94/gnd DFFSR_25/S FILL
XFILL_34_DFFSR_30 INVX1_89/gnd DFFSR_36/S FILL
XFILL_6_DFFSR_77 INVX1_89/gnd DFFSR_2/S FILL
XFILL_4_INVX1_399 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_23_DFFSR_70 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_6_DFFSR_135 BUFX2_43/A DFFSR_97/S FILL
XFILL_47_DFFSR_166 INVX1_4/gnd DFFSR_51/S FILL
XFILL_37_DFFSR_169 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_5_BUFX2_15 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_27_DFFSR_172 BUFX2_37/A DFFSR_8/S FILL
XFILL_3_INVX1_219 INVX1_94/gnd DFFSR_52/S FILL
XFILL_3_OAI21X1_130 INVX1_4/gnd DFFSR_4/S FILL
XFILL_17_DFFSR_175 INVX1_23/gnd DFFSR_91/S FILL
XFILL_9_AOI22X1_7 BUFX2_43/A DFFSR_23/S FILL
XFILL_8_OAI21X1_94 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_7_OAI21X1_97 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_3_INVX1_71 INVX1_94/gnd DFFSR_25/S FILL
XFILL_42_DFFSR_37 INVX1_89/gnd DFFSR_2/S FILL
XOAI21X1_5 DFFSR_5/S INVX1_6/Y OAI21X1_5/C INVX1_8/gnd DFFSR_5/D DFFSR_5/S OAI21X1
XFILL_3_NAND2X1_244 INVX1_94/gnd DFFSR_52/S FILL
XFILL_3_XOR2X1_14 INVX1_89/gnd DFFSR_2/S FILL
XFILL_31_DFFSR_77 INVX1_89/gnd DFFSR_2/S FILL
XFILL_4_OAI21X1_2 INVX1_8/gnd DFFSR_5/S FILL
XFILL_2_NOR2X1_54 DFFSR_1/gnd DFFSR_9/S FILL
XNAND2X1_118 BUFX2_24/Y DFFSR_110/Q DFFSR_73/gnd OAI21X1_118/C DFFSR_11/S NAND2X1
XFILL_1_INVX1_436 INVX1_89/gnd DFFSR_36/S FILL
XFILL_8_AOI21X1_10 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_3_DFFSR_172 BUFX2_37/A DFFSR_8/S FILL
XFILL_7_AOI21X1_13 INVX1_8/gnd DFFSR_7/S FILL
XFILL_15_DFFSR_27 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_6_AOI21X1_16 BUFX2_43/A DFFSR_23/S FILL
XFILL_1_OAI21X1_226 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_7_DFFPOSX1_16 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_5_AOI21X1_19 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_4_NAND2X1_178 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_4_DFFPOSX1_2 INVX1_89/gnd DFFSR_36/S FILL
XFILL_20_DFFSR_102 INVX1_8/gnd DFFSR_7/S FILL
XFILL_10_DFFSR_105 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_4_AOI21X1_22 BUFX2_43/A DFFSR_97/S FILL
XAOI21X1_16 AOI22X1_8/C AOI22X1_8/D AOI21X1_25/A BUFX2_43/A AOI21X1_16/Y DFFSR_23/S
+ AOI21X1
XFILL_3_DFFPOSX1_5 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_3_AOI21X1_25 BUFX2_43/A DFFSR_97/S FILL
XFILL_39_DFFSR_84 BUFX2_43/A DFFSR_23/S FILL
XFILL_0_INVX1_256 BUFX2_36/A DFFSR_8/S FILL
XINVX1_366 DFFSR_117/Q BUFX2_37/A INVX1_366/Y DFFSR_81/S INVX1
XFILL_50_DFFSR_44 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_2_DFFPOSX1_8 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_2_AOI21X1_28 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_2_OAI21X1_160 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_1_AOI21X1_31 INVX1_23/gnd DFFSR_186/S FILL
XFILL_17_CLKBUF1_7 BUFX2_43/A DFFSR_97/S FILL
XFILL_6_DFFSR_41 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_23_DFFSR_34 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_12_DFFSR_74 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_5_NAND2X1_112 INVX1_4/gnd DFFSR_4/S FILL
XFILL_0_AOI21X1_34 INVX1_94/gnd DFFSR_25/S FILL
XFILL_47_DFFSR_130 INVX1_4/gnd DFFSR_51/S FILL
XFILL_37_DFFSR_133 BUFX2_37/A DFFSR_81/S FILL
XFILL_26_DFFPOSX1_24 BUFX2_43/A DFFSR_23/S FILL
XFILL_14_1 BUFX2_36/A DFFSR_8/S FILL
XBUFX2_19 INVX1_1/Y BUFX2_19/gnd BUFX2_19/Y DFFSR_54/S BUFX2
XFILL_27_DFFSR_136 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_2_NAND2X1_274 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_47_DFFSR_91 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_3_INVX1_183 BUFX2_37/A DFFSR_8/S FILL
XFILL_3_CLKBUF1_4 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_17_DFFSR_139 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_8_OAI21X1_58 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_6_NAND2X1_79 INVX1_89/gnd DFFSR_36/S FILL
XFILL_3_INVX1_35 BUFX2_35/A DFFSR_97/S FILL
XFILL_7_OAI21X1_61 BUFX2_36/A DFFSR_8/S FILL
XFILL_20_DFFSR_81 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_2_NOR2X1_18 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_31_DFFSR_41 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_0_OAI21X1_256 INVX1_2/gnd DFFSR_51/S FILL
XFILL_3_DFFSR_88 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_3_NAND2X1_208 BUFX2_8/gnd DFFSR_10/S FILL
XNAND2X1_79 BUFX2_22/Y INVX1_80/A INVX1_89/gnd NAND2X1_79/Y DFFSR_36/S NAND2X1
XFILL_5_NAND2X1_82 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_6_OAI21X1_64 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_1_INVX1_400 BUFX2_35/A DFFSR_97/S FILL
XFILL_2_NAND3X1_106 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_4_NAND2X1_85 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_29_2_0 INVX1_89/gnd DFFSR_2/S FILL
XFILL_5_OAI21X1_67 INVX1_2/gnd DFFSR_1/S FILL
XOAI21X1_64 DFFSR_65/S INVX1_72/Y NAND2X1_64/Y BUFX2_16/gnd DFFSR_64/D DFFSR_65/S
+ OAI21X1
XFILL_44_DFFSR_167 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_3_DFFSR_136 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_2_BUFX2_26 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_3_NAND2X1_88 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_4_OAI21X1_70 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_2_NAND2X1_91 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_1_OAI21X1_190 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_4_NAND2X1_142 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_1_DFFSR_1 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_3_OAI21X1_73 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_34_DFFSR_170 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_2_OAI21X1_76 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_27_4_1 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_1_NAND2X1_94 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_24_DFFSR_173 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_0_INVX1_82 BUFX2_35/A DFFSR_97/S FILL
XFILL_9_3_0 BUFX2_43/A DFFSR_23/S FILL
XFILL_0_NAND2X1_97 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_0_INVX1_220 INVX1_94/gnd DFFSR_52/S FILL
XINVX1_330 DFFSR_73/Q DFFSR_71/gnd INVX1_330/Y DFFSR_45/S INVX1
XFILL_1_OAI21X1_79 INVX1_89/gnd DFFSR_36/S FILL
XFILL_39_DFFSR_48 INVX1_4/gnd DFFSR_4/S FILL
XFILL_28_DFFSR_88 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_6_AOI22X1_8 BUFX2_43/A DFFSR_97/S FILL
XFILL_0_OAI21X1_82 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_14_DFFSR_176 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_7_5_1 BUFX2_35/A DFFSR_97/S FILL
XFILL_2_OAI21X1_124 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_4_INVX1_327 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_0_XOR2X1_15 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_12_DFFSR_38 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_1_OAI21X1_3 INVX1_4/gnd DFFSR_51/S FILL
XFILL_0_DFFSR_173 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_2_NAND2X1_238 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_27_DFFSR_100 INVX1_23/gnd DFFSR_186/S FILL
XFILL_6_AND2X2_14 BUFX2_35/A DFFSR_97/S FILL
XFILL_36_DFFSR_95 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_47_DFFSR_55 INVX1_89/gnd DFFSR_36/S FILL
XFILL_25_DFFSR_5 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_3_INVX1_147 INVX1_4/gnd DFFSR_4/S FILL
XFILL_8_OAI21X1_22 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_17_DFFSR_103 INVX1_8/gnd DFFSR_7/S FILL
XFILL_3_DFFSR_52 INVX1_94/gnd DFFSR_52/S FILL
XFILL_7_OAI21X1_25 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_6_NAND2X1_43 INVX1_89/gnd DFFSR_2/S FILL
XFILL_0_OAI21X1_220 BUFX2_43/A DFFSR_97/S FILL
XFILL_3_NAND2X1_172 BUFX2_36/A DFFSR_6/S FILL
XFILL_6_OAI21X1_28 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_5_NAND2X1_46 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_20_DFFSR_45 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_6_DFFPOSX1_10 INVX1_8/gnd DFFSR_5/S FILL
XFILL_5_OAI21X1_31 BUFX2_35/A DFFSR_97/S FILL
XFILL_1_INVX1_364 DFFSR_71/gnd DFFSR_10/S FILL
XNAND2X1_43 DFFSR_2/S DFFSR_35/Q INVX1_89/gnd OAI21X1_43/C DFFSR_2/S NAND2X1
XFILL_4_NAND2X1_49 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_3_DFFSR_100 INVX1_23/gnd DFFSR_186/S FILL
XFILL_14_CLKBUF1_8 BUFX2_5/gnd DFFSR_6/S FILL
XOAI21X1_28 DFFSR_54/S INVX1_32/Y OAI21X1_28/C BUFX2_7/gnd DFFSR_28/D DFFSR_81/S OAI21X1
XFILL_3_NAND2X1_52 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_4_OAI21X1_34 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_3_OAI21X1_37 INVX1_89/gnd DFFSR_2/S FILL
XFILL_2_NAND2X1_55 INVX1_89/gnd DFFSR_2/S FILL
XFILL_46_DFFSR_1 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_44_DFFSR_131 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_15_DFFPOSX1_29 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_1_OAI21X1_154 BUFX2_37/A DFFSR_8/S FILL
XFILL_34_DFFSR_134 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_2_OAI21X1_40 INVX1_8/gnd DFFSR_7/S FILL
XFILL_4_NAND2X1_106 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_1_NAND2X1_58 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_0_NAND2X1_61 BUFX2_37/A DFFSR_81/S FILL
XFILL_24_DFFSR_137 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_1_OAI21X1_43 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_35_1_2 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_17_DFFSR_92 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_39_DFFSR_12 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_0_DFFSR_99 BUFX2_35/A DFFSR_97/S FILL
XFILL_0_OAI21X1_46 BUFX2_37/A DFFSR_81/S FILL
XFILL_0_INVX1_184 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_19_6 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_28_DFFSR_52 INVX1_94/gnd DFFSR_52/S FILL
XINVX1_294 INVX1_32/A DFFSR_71/gnd INVX1_294/Y DFFSR_10/S INVX1
XFILL_14_DFFSR_140 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_0_INVX1_46 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_0_CLKBUF1_5 INVX1_89/gnd DFFSR_2/S FILL
XFILL_1_NAND2X1_268 BUFX2_37/A DFFSR_8/S FILL
XFILL_4_INVX1_291 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_36_1 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_9_AOI22X1_12 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_25_DFFPOSX1_18 BUFX2_37/A DFFSR_8/S FILL
XFILL_1_INVX1_3 INVX1_8/gnd DFFSR_5/S FILL
XFILL_2_NAND2X1_202 BUFX2_35/A DFFSR_97/S FILL
XFILL_41_DFFSR_168 BUFX2_36/A DFFSR_8/S FILL
XFILL_0_DFFSR_137 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_25_DFFSR_99 BUFX2_35/A DFFSR_97/S FILL
XFILL_47_DFFSR_19 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_3_INVX1_111 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_36_DFFSR_59 INVX1_4/gnd DFFSR_51/S FILL
XFILL_1_NAND3X1_100 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_31_DFFSR_171 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_21_DFFSR_174 BUFX2_43/A DFFSR_97/S FILL
XFILL_0_OAI21X1_184 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_3_DFFSR_16 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_3_AOI22X1_9 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_3_NAND2X1_136 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_11_DFFSR_177 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_5_NAND2X1_10 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_11_OAI22X1_54 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_6_NOR2X1_53 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_1_INVX1_328 INVX1_8/gnd DFFSR_7/S FILL
XFILL_7_XOR2X1_13 INVX1_8/gnd DFFSR_7/S FILL
XFILL_8_OAI21X1_1 INVX1_2/gnd DFFSR_51/S FILL
XFILL_4_NAND2X1_13 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_3_NAND2X1_16 DFFSR_79/gnd DFFSR_36/S FILL
XDFFPOSX1_10 INVX1_397/A CLKBUF1_9/Y NAND2X1_250/Y INVX1_8/gnd DFFSR_5/S DFFPOSX1
XFILL_10_OAI22X1_57 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_7_DFFSR_171 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_2_NAND2X1_19 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_44_DFFSR_66 INVX1_2/gnd DFFSR_51/S FILL
XFILL_1_OAI21X1_118 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_1_NAND2X1_22 BUFX2_19/gnd DFFSR_52/S FILL
XINVX1_258 INVX1_258/A BUFX2_43/A INVX1_258/Y DFFSR_23/S INVX1
XFILL_0_INVX1_10 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_8_NAND3X1_78 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_0_DFFSR_63 INVX1_94/gnd DFFSR_52/S FILL
XFILL_28_DFFSR_16 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_0_NAND2X1_25 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_9_OAI22X1_60 INVX1_8/gnd DFFSR_5/S FILL
XFILL_0_INVX1_148 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_17_DFFSR_56 INVX1_2/gnd DFFSR_51/S FILL
XFILL_3_AND2X2_15 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_24_DFFSR_101 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_7_NAND3X1_81 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_8_OAI22X1_63 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_0_OAI21X1_10 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_14_DFFSR_104 INVX1_4/gnd DFFSR_4/S FILL
XFILL_4_INVX1_255 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_1_NAND2X1_232 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_6_NAND3X1_84 INVX1_94/gnd DFFSR_25/S FILL
XFILL_7_OAI22X1_66 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_0_NAND3X1_130 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_5_NAND3X1_87 INVX1_94/gnd DFFSR_52/S FILL
XFILL_4_NAND3X1_90 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_21_CLKBUF1_6 BUFX2_5/gnd DFFSR_23/S FILL
XNAND3X1_84 NAND3X1_55/Y NAND3X1_82/Y NAND3X1_83/Y INVX1_94/gnd NAND3X1_84/Y DFFSR_25/S
+ NAND3X1
XFILL_3_NAND3X1_93 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_11_CLKBUF1_9 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_51_DFFSR_129 INVX1_2/gnd DFFSR_1/S FILL
XFILL_2_NAND2X1_166 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_0_DFFSR_101 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_2_NAND3X1_96 BUFX2_43/A DFFSR_97/S FILL
XFILL_36_DFFSR_23 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_25_DFFSR_63 INVX1_94/gnd DFFSR_52/S FILL
XFILL_8_DFFSR_70 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_41_DFFSR_132 INVX1_2/gnd DFFSR_51/S FILL
XFILL_1_NAND3X1_99 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_31_DFFSR_135 BUFX2_43/A DFFSR_97/S FILL
XFILL_14_DFFPOSX1_23 INVX1_23/gnd DFFSR_91/S FILL
XFILL_7_CLKBUF1_3 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_21_DFFSR_138 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_0_OAI21X1_148 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_3_NAND2X1_100 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_9_OAI21X1_203 BUFX2_35/A DFFSR_14/S FILL
XFILL_11_DFFSR_141 INVX1_94/gnd DFFSR_25/S FILL
XFILL_1_INVX1_292 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_6_NOR2X1_17 INVX1_4/gnd DFFSR_4/S FILL
XFILL_37_DFFSR_8 BUFX2_36/A DFFSR_8/S FILL
XFILL_41_6 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_0_NAND2X1_262 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_44_DFFSR_30 INVX1_89/gnd DFFSR_36/S FILL
XFILL_10_OAI22X1_21 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_7_DFFSR_135 BUFX2_43/A DFFSR_97/S FILL
XFILL_9_NAND3X1_39 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_24_DFFPOSX1_12 INVX1_8/gnd DFFSR_5/S FILL
XFILL_33_DFFSR_70 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_48_DFFSR_166 INVX1_4/gnd DFFSR_51/S FILL
XFILL_8_NAND3X1_42 BUFX2_43/A DFFSR_23/S FILL
XFILL_9_OAI22X1_24 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_17_DFFSR_20 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_7_NAND3X1_45 BUFX2_35/A DFFSR_97/S FILL
XFILL_0_INVX1_112 BUFX2_43/A DFFSR_97/S FILL
XFILL_38_DFFSR_169 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_8_OAI22X1_27 DFFSR_79/gnd DFFSR_36/S FILL
XINVX1_222 NAND3X1_6/Y BUFX2_17/gnd NOR2X1_5/B DFFSR_7/S INVX1
XFILL_0_DFFSR_27 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_6_NAND3X1_48 BUFX2_43/A DFFSR_23/S FILL
XFILL_28_DFFSR_172 BUFX2_37/A DFFSR_8/S FILL
XFILL_1_NAND2X1_196 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_7_OAI22X1_30 INVX1_94/gnd DFFSR_25/S FILL
XFILL_18_DFFSR_175 INVX1_23/gnd DFFSR_91/S FILL
XFILL_5_NAND3X1_51 BUFX2_7/gnd DFFSR_81/S FILL
XXOR2X1_17 XOR2X1_17/A DFFSR_137/Q BUFX2_19/gnd XOR2X1_17/Y DFFSR_52/S XOR2X1
XFILL_8_NOR3X1_1 INVX1_94/gnd DFFSR_52/S FILL
XFILL_6_OAI22X1_33 DFFSR_73/gnd DFFSR_57/S FILL
XNAND3X1_48 AOI22X1_5/Y NAND3X1_48/B NAND3X1_42/Y BUFX2_43/A AOI22X1_8/D DFFSR_23/S
+ NAND3X1
XFILL_4_NAND3X1_54 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_5_OAI22X1_36 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_36_2_0 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_3_NAND3X1_57 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_4_XOR2X1_14 INVX1_89/gnd DFFSR_2/S FILL
XFILL_41_DFFSR_77 INVX1_89/gnd DFFSR_2/S FILL
XFILL_5_OAI21X1_2 INVX1_8/gnd DFFSR_5/S FILL
XOAI22X1_33 INVX1_321/Y OAI22X1_6/D INVX1_322/Y OAI22X1_9/B DFFSR_73/gnd NOR2X1_26/B
+ DFFSR_57/S OAI22X1
XFILL_3_NOR2X1_54 DFFSR_1/gnd DFFSR_9/S FILL
XDFFSR_175 DFFSR_175/Q CLKBUF1_14/Y DFFSR_175/R DFFSR_91/S DFFSR_175/D INVX1_23/gnd
+ DFFSR_91/S DFFSR
XFILL_8_OAI21X1_233 BUFX2_36/A DFFSR_8/S FILL
XFILL_4_OAI22X1_39 BUFX2_37/A DFFSR_8/S FILL
XFILL_2_INVX1_436 INVX1_89/gnd DFFSR_36/S FILL
XFILL_34_4_1 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_2_NAND2X1_130 INVX1_4/gnd DFFSR_4/S FILL
XFILL_4_DFFSR_172 BUFX2_37/A DFFSR_8/S FILL
XFILL_2_NAND3X1_60 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_3_OAI22X1_42 INVX1_8/gnd DFFSR_7/S FILL
XFILL_25_DFFSR_27 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_8_DFFSR_34 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_14_DFFSR_67 INVX1_2/gnd DFFSR_51/S FILL
XFILL_1_NAND3X1_63 BUFX2_43/A DFFSR_23/S FILL
XFILL_2_OAI22X1_45 INVX1_89/gnd DFFSR_2/S FILL
XFILL_0_NAND3X1_66 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_1_OAI22X1_48 BUFX2_37/A DFFSR_81/S FILL
XFILL_0_AND2X2_16 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_21_DFFSR_102 INVX1_8/gnd DFFSR_7/S FILL
XFILL_0_OAI21X1_112 INVX1_4/gnd DFFSR_4/S FILL
XFILL_1_XOR2X1_4 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_11_DFFSR_105 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_0_OAI22X1_51 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_49_DFFSR_84 BUFX2_43/A DFFSR_23/S FILL
XFILL_1_INVX1_256 BUFX2_36/A DFFSR_8/S FILL
XFILL_18_CLKBUF1_7 BUFX2_43/A DFFSR_97/S FILL
XFILL_0_NAND2X1_226 BUFX2_36/A DFFSR_6/S FILL
XINVX1_68 DFFSR_60/Q BUFX2_37/A INVX1_68/Y DFFSR_81/S INVX1
XFILL_5_DFFSR_81 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_33_DFFSR_34 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_22_DFFSR_74 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_48_DFFSR_130 INVX1_4/gnd DFFSR_51/S FILL
XINVX1_186 DFFSR_156/Q BUFX2_6/gnd INVX1_186/Y DFFSR_14/S INVX1
XFILL_38_DFFSR_133 BUFX2_37/A DFFSR_81/S FILL
XCLKBUF1_7 DFFSR_149/Q BUFX2_43/A CLKBUF1_7/Y DFFSR_97/S CLKBUF1
XFILL_4_BUFX2_19 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_28_DFFSR_136 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_1_NAND2X1_160 INVX1_8/gnd DFFSR_5/S FILL
XFILL_4_INVX1_183 BUFX2_37/A DFFSR_8/S FILL
XFILL_6_NAND3X1_12 INVX1_94/gnd DFFSR_52/S FILL
XFILL_4_CLKBUF1_4 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_7_OAI21X1_263 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_18_DFFSR_139 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_5_NAND3X1_15 BUFX2_19/gnd DFFSR_52/S FILL
XNAND3X1_12 AOI21X1_8/A AOI21X1_8/B AOI21X1_2/Y INVX1_94/gnd AOI21X1_9/B DFFSR_52/S
+ NAND3X1
XFILL_24_DFFSR_2 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_30_DFFSR_81 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_3_NOR2X1_18 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_4_NAND3X1_18 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_41_DFFSR_41 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_2_INVX1_75 INVX1_4/gnd DFFSR_51/S FILL
XFILL_13_DFFPOSX1_17 BUFX2_37/A DFFSR_8/S FILL
XFILL_3_NAND3X1_21 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_8_OAI21X1_197 INVX1_8/gnd DFFSR_7/S FILL
XDFFSR_139 XOR2X1_11/B CLKBUF1_13/Y DFFSR_137/R DFFSR_4/S DFFSR_139/D DFFSR_3/gnd
+ DFFSR_4/S DFFSR
XFILL_14_DFFSR_31 BUFX2_35/A DFFSR_97/S FILL
XFILL_2_INVX1_400 BUFX2_35/A DFFSR_97/S FILL
XFILL_2_NAND3X1_24 BUFX2_37/A DFFSR_8/S FILL
XFILL_42_1_2 INVX1_4/gnd DFFSR_4/S FILL
XFILL_1_NAND3X1_27 BUFX2_37/A DFFSR_81/S FILL
XFILL_45_DFFSR_167 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_4_DFFSR_136 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_0_NAND3X1_30 INVX1_94/gnd DFFSR_52/S FILL
XFILL_1_OAI22X1_12 INVX1_4/gnd DFFSR_51/S FILL
XFILL_35_DFFSR_170 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_9_OAI21X1_131 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_0_OAI22X1_15 INVX1_4/gnd DFFSR_4/S FILL
XFILL_25_DFFSR_173 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_1_INVX1_220 INVX1_94/gnd DFFSR_52/S FILL
XFILL_49_DFFSR_48 INVX1_4/gnd DFFSR_4/S FILL
XFILL_38_DFFSR_88 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_7_AOI22X1_8 BUFX2_43/A DFFSR_97/S FILL
XFILL_15_DFFSR_176 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_0_NAND2X1_190 BUFX2_35/A DFFSR_97/S FILL
XFILL_10_0_0 BUFX2_5/gnd DFFSR_23/S FILL
XINVX1_32 INVX1_32/A BUFX2_7/gnd INVX1_32/Y DFFSR_54/S INVX1
XDFFSR_85 DFFSR_85/Q CLKBUF1_2/Y DFFSR_84/R DFFSR_45/S DFFSR_85/D DFFSR_71/gnd DFFSR_45/S
+ DFFSR
XFILL_5_DFFSR_45 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_3_DFFPOSX1_28 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_1_XOR2X1_15 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_22_DFFSR_38 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_11_DFFSR_78 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_2_OAI21X1_3 INVX1_4/gnd DFFSR_51/S FILL
XFILL_1_2 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_1_DFFSR_173 BUFX2_6/gnd DFFSR_91/S FILL
XINVX1_150 DFFSR_133/Q BUFX2_7/gnd INVX1_150/Y DFFSR_54/S INVX1
XFILL_28_DFFSR_100 INVX1_23/gnd DFFSR_186/S FILL
XFILL_7_AND2X2_14 BUFX2_35/A DFFSR_97/S FILL
XFILL_7_OAI21X1_227 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_15_XOR2X1_8 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_46_DFFSR_95 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_1_NAND2X1_124 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_18_DFFSR_103 INVX1_8/gnd DFFSR_7/S FILL
XFILL_7_AND2X2_4 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_2_DFFSR_92 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_19_DFFSR_85 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_30_DFFSR_45 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_2_INVX1_39 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_8_OAI21X1_161 INVX1_23/gnd DFFSR_186/S FILL
XFILL_2_INVX1_364 DFFSR_71/gnd DFFSR_10/S FILL
XDFFSR_103 INVX1_116/A CLKBUF1_4/Y DFFSR_97/R DFFSR_7/S DFFSR_103/D INVX1_8/gnd DFFSR_7/S
+ DFFSR
XFILL_4_DFFSR_100 INVX1_23/gnd DFFSR_186/S FILL
XFILL_15_CLKBUF1_8 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_1_BUFX2_30 INVX1_4/gnd DFFSR_51/S FILL
XFILL_45_DFFSR_131 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_35_DFFSR_134 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_25_DFFSR_137 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_27_DFFSR_92 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_49_DFFSR_12 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_1_INVX1_184 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_38_DFFSR_52 INVX1_94/gnd DFFSR_52/S FILL
XFILL_23_3 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_15_DFFSR_140 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_1_CLKBUF1_5 INVX1_89/gnd DFFSR_2/S FILL
XFILL_0_NAND2X1_154 BUFX2_37/A DFFSR_8/S FILL
XFILL_0_NOR2X1_19 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_6_OAI21X1_257 INVX1_2/gnd DFFSR_51/S FILL
XFILL_11_DFFSR_42 DFFSR_3/gnd DFFSR_65/S FILL
XDFFSR_49 DFFSR_49/Q DFFSR_2/CLK DFFSR_54/R DFFSR_49/S DFFSR_49/D DFFSR_73/gnd DFFSR_11/S
+ DFFSR
XFILL_8_NAND3X1_107 BUFX2_43/A DFFSR_97/S FILL
XINVX1_114 INVX1_368/A BUFX2_17/gnd INVX1_114/Y DFFSR_7/S INVX1
XFILL_1_DFFSR_137 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_15_DFFSR_9 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_12_DFFPOSX1_11 INVX1_4/gnd DFFSR_4/S FILL
XFILL_35_DFFSR_99 BUFX2_35/A DFFSR_97/S FILL
XFILL_42_DFFSR_168 BUFX2_36/A DFFSR_8/S FILL
XFILL_7_OAI21X1_191 BUFX2_37/A DFFSR_8/S FILL
XFILL_46_DFFSR_59 INVX1_4/gnd DFFSR_51/S FILL
XFILL_32_DFFSR_171 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_22_DFFSR_174 BUFX2_43/A DFFSR_97/S FILL
XFILL_2_DFFSR_56 INVX1_2/gnd DFFSR_51/S FILL
XFILL_19_DFFSR_49 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_8_OAI21X1_125 BUFX2_35/A DFFSR_14/S FILL
XFILL_4_AOI22X1_9 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_12_DFFSR_177 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_2_INVX1_328 INVX1_8/gnd DFFSR_7/S FILL
XFILL_8_XOR2X1_13 INVX1_8/gnd DFFSR_7/S FILL
XFILL_8_DFFSR_171 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_36_DFFSR_5 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_2_DFFPOSX1_22 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_38_DFFSR_16 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_16_DFFSR_96 INVX1_2/gnd DFFSR_1/S FILL
XFILL_1_INVX1_148 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_27_DFFSR_56 INVX1_2/gnd DFFSR_51/S FILL
XFILL_43_2_0 INVX1_4/gnd DFFSR_51/S FILL
XFILL_4_AND2X2_15 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_25_DFFSR_101 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_15_DFFSR_104 INVX1_4/gnd DFFSR_4/S FILL
XFILL_6_OAI21X1_221 BUFX2_35/A DFFSR_14/S FILL
XFILL_41_4_1 DFFSR_3/gnd DFFSR_4/S FILL
XDFFSR_13 DFFSR_13/Q DFFSR_3/CLK DFFSR_9/R DFFSR_13/S DFFSR_13/D BUFX2_16/gnd DFFSR_65/S
+ DFFSR
XFILL_0_NAND2X1_118 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_12_CLKBUF1_9 BUFX2_17/gnd DFFSR_7/S FILL
XOAI21X1_257 DFFSR_166/S INVX1_420/Y NAND2X1_268/Y INVX1_2/gnd DFFSR_189/D DFFSR_51/S
+ OAI21X1
XFILL_1_DFFSR_101 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_21_DFFPOSX1_30 BUFX2_43/A DFFSR_97/S FILL
XFILL_46_DFFSR_23 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_7_OAI21X1_155 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_35_DFFSR_63 INVX1_94/gnd DFFSR_52/S FILL
XFILL_42_DFFSR_132 INVX1_2/gnd DFFSR_51/S FILL
XFILL_32_DFFSR_135 BUFX2_43/A DFFSR_97/S FILL
XFILL_8_CLKBUF1_3 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_22_DFFSR_138 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_2_DFFSR_20 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_12_DFFSR_141 INVX1_94/gnd DFFSR_25/S FILL
XFILL_19_DFFSR_13 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_2_INVX1_292 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_1_NOR2X1_1 BUFX2_36/A DFFSR_6/S FILL
XFILL_45_3 INVX1_2/gnd DFFSR_51/S FILL
XFILL_5_OAI21X1_251 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_8_DFFSR_135 BUFX2_43/A DFFSR_97/S FILL
XFILL_43_DFFSR_70 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_49_DFFSR_166 INVX1_4/gnd DFFSR_51/S FILL
XFILL_27_DFFSR_20 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_7_NAND3X1_101 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_1_INVX1_112 BUFX2_43/A DFFSR_97/S FILL
XFILL_17_CLKBUF1_12 BUFX2_43/A DFFSR_23/S FILL
XFILL_39_DFFSR_169 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_16_DFFSR_60 BUFX2_37/A DFFSR_8/S FILL
XFILL_29_DFFSR_172 BUFX2_37/A DFFSR_8/S FILL
XFILL_16_CLKBUF1_15 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_19_DFFSR_175 INVX1_23/gnd DFFSR_91/S FILL
XFILL_6_OAI21X1_185 BUFX2_36/A DFFSR_8/S FILL
XFILL_15_CLKBUF1_18 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_3_DFFSR_8 BUFX2_36/A DFFSR_8/S FILL
XFILL_14_CLKBUF1_21 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_13_CLKBUF1_24 INVX1_23/gnd DFFSR_186/S FILL
XFILL_5_XOR2X1_14 INVX1_89/gnd DFFSR_2/S FILL
XFILL_51_DFFSR_77 INVX1_89/gnd DFFSR_2/S FILL
XFILL_4_NOR2X1_54 DFFSR_1/gnd DFFSR_9/S FILL
XOAI21X1_221 INVX1_249/A NOR2X1_9/Y INVX1_248/Y BUFX2_35/A NAND3X1_67/B DFFSR_14/S
+ OAI21X1
XFILL_3_INVX1_436 INVX1_89/gnd DFFSR_36/S FILL
XFILL_6_OAI21X1_2 INVX1_8/gnd DFFSR_5/S FILL
XFILL_5_DFFSR_172 BUFX2_37/A DFFSR_8/S FILL
XFILL_7_OAI21X1_119 BUFX2_37/A DFFSR_8/S FILL
XFILL_35_DFFSR_27 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_7_DFFSR_74 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_24_DFFSR_67 INVX1_2/gnd DFFSR_51/S FILL
XFILL_1_DFFPOSX1_16 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_1_AND2X2_16 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_22_DFFSR_102 INVX1_8/gnd DFFSR_7/S FILL
XFILL_12_DFFSR_105 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_6_BUFX2_12 BUFX2_37/A DFFSR_81/S FILL
XFILL_17_0_0 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_2_INVX1_256 BUFX2_36/A DFFSR_8/S FILL
XFILL_15_2_1 BUFX2_37/A DFFSR_81/S FILL
XFILL_6_NAND3X1_131 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_5_OAI21X1_215 BUFX2_43/A DFFSR_97/S FILL
XFILL_19_CLKBUF1_7 BUFX2_43/A DFFSR_97/S FILL
XFILL_43_DFFSR_34 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_32_DFFSR_74 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_13_4_2 BUFX2_36/A DFFSR_8/S FILL
XFILL_49_DFFSR_130 INVX1_4/gnd DFFSR_51/S FILL
XFILL_39_DFFSR_133 BUFX2_37/A DFFSR_81/S FILL
XFILL_16_DFFSR_24 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_29_DFFSR_136 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_6_OAI21X1_149 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_20_DFFPOSX1_24 BUFX2_43/A DFFSR_23/S FILL
XFILL_5_CLKBUF1_4 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_19_DFFSR_139 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_48_DFFSR_8 BUFX2_36/A DFFSR_8/S FILL
XNOR2X1_21 NOR2X1_21/A NOR2X1_21/B DFFSR_79/gnd NOR2X1_21/Y DFFSR_36/S NOR2X1
XFILL_40_DFFSR_81 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_4_NOR2X1_18 BUFX2_8/gnd DFFSR_10/S FILL
XOAI21X1_185 INVX1_216/Y INVX1_226/Y OAI22X1_2/A BUFX2_36/A AOI22X1_3/C DFFSR_8/S
+ OAI21X1
XFILL_24_DFFSR_31 BUFX2_35/A DFFSR_97/S FILL
XFILL_3_INVX1_400 BUFX2_35/A DFFSR_97/S FILL
XFILL_7_DFFSR_38 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_6_NAND2X1_263 INVX1_2/gnd DFFSR_51/S FILL
XFILL_13_DFFSR_71 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_5_DFFSR_136 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_46_DFFSR_167 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_36_DFFSR_170 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_4_OAI21X1_245 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_26_DFFSR_173 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_0_XOR2X1_8 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_2_INVX1_220 INVX1_94/gnd DFFSR_52/S FILL
XFILL_48_DFFSR_88 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_8_AOI22X1_8 BUFX2_43/A DFFSR_97/S FILL
XFILL_16_DFFSR_176 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_4_INVX1_32 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_5_OAI21X1_179 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_4_DFFSR_85 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_2_XOR2X1_15 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_32_DFFSR_38 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_21_DFFSR_78 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_0_INVX1_437 BUFX2_35/A DFFSR_97/S FILL
XFILL_5_CLKBUF1_12 BUFX2_43/A DFFSR_23/S FILL
XNAND3X1_131 NOR2X1_1/B NOR2X1_1/A NOR2X1_2/A BUFX2_7/gnd INVX1_405/A DFFSR_54/S NAND3X1
XFILL_3_OAI21X1_3 INVX1_4/gnd DFFSR_51/S FILL
XFILL_2_DFFSR_173 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_3_BUFX2_23 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_4_CLKBUF1_15 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_29_DFFSR_100 INVX1_23/gnd DFFSR_186/S FILL
XFILL_3_0_2 INVX1_23/gnd DFFSR_91/S FILL
XFILL_8_AND2X2_14 BUFX2_35/A DFFSR_97/S FILL
XFILL_3_CLKBUF1_18 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_6_OAI21X1_113 INVX1_23/gnd DFFSR_91/S FILL
XFILL_14_DFFSR_6 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_13_NOR3X1_2 INVX1_89/gnd DFFSR_2/S FILL
XFILL_19_DFFSR_103 INVX1_8/gnd DFFSR_7/S FILL
XFILL_2_CLKBUF1_21 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_1_CLKBUF1_24 INVX1_23/gnd DFFSR_186/S FILL
XFILL_29_DFFSR_85 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_40_DFFSR_45 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_0_DFFPOSX1_10 INVX1_8/gnd DFFSR_5/S FILL
XFILL_1_INVX1_79 DFFSR_73/gnd DFFSR_57/S FILL
XOAI21X1_149 DFFSR_91/S INVX1_172/Y OAI21X1_149/C DFFSR_89/gnd DFFSR_149/D DFFSR_186/S
+ OAI21X1
XFILL_6_NAND2X1_227 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_3_INVX1_364 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_5_DFFSR_100 INVX1_23/gnd DFFSR_186/S FILL
XFILL_16_CLKBUF1_8 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_13_DFFSR_35 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_5_NAND3X1_125 INVX1_8/gnd DFFSR_5/S FILL
XFILL_46_DFFSR_131 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_36_DFFSR_134 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_48_4_1 DFFSR_9/gnd DFFSR_9/S FILL
XNAND2X1_263 DFFSR_160/Q DFFSR_1/S INVX1_2/gnd NAND2X1_263/Y DFFSR_51/S NAND2X1
XFILL_10_5 BUFX2_43/A DFFSR_23/S FILL
XFILL_26_DFFSR_137 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_35_DFFSR_2 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_4_OAI21X1_209 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_37_DFFSR_92 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_2_INVX1_184 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_48_DFFSR_52 INVX1_94/gnd DFFSR_52/S FILL
XFILL_16_DFFSR_140 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_2_CLKBUF1_5 INVX1_89/gnd DFFSR_2/S FILL
XFILL_19_DFFPOSX1_18 BUFX2_37/A DFFSR_8/S FILL
XFILL_1_NOR2X1_19 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_5_OAI21X1_143 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_10_DFFSR_82 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_21_DFFSR_42 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_4_DFFSR_49 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_0_INVX1_401 BUFX2_35/A DFFSR_14/S FILL
XFILL_2_DFFSR_137 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_27_DFFPOSX1_6 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_45_DFFSR_99 BUFX2_35/A DFFSR_97/S FILL
XFILL_43_DFFSR_168 BUFX2_36/A DFFSR_8/S FILL
XFILL_26_DFFPOSX1_9 BUFX2_37/A DFFSR_8/S FILL
XFILL_5_NAND2X1_257 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_14_5_0 BUFX2_37/A DFFSR_8/S FILL
XFILL_33_DFFSR_171 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_18_DFFSR_89 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_23_DFFSR_174 BUFX2_43/A DFFSR_97/S FILL
XFILL_6_AND2X2_8 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_1_INVX1_43 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_1_DFFSR_96 INVX1_2/gnd DFFSR_1/S FILL
XFILL_29_DFFSR_49 DFFSR_73/gnd DFFSR_11/S FILL
XOAI21X1_113 BUFX2_21/Y INVX1_128/Y NAND2X1_113/Y INVX1_23/gnd DFFSR_113/D DFFSR_91/S
+ OAI21X1
XFILL_5_AOI22X1_9 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_13_DFFSR_177 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_9_DFFPOSX1_29 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_3_OAI21X1_239 INVX1_4/gnd DFFSR_4/S FILL
XFILL_6_NAND2X1_191 BUFX2_37/A DFFSR_8/S FILL
XFILL_3_INVX1_328 INVX1_8/gnd DFFSR_7/S FILL
XFILL_9_XOR2X1_13 INVX1_8/gnd DFFSR_7/S FILL
XFILL_0_BUFX2_34 BUFX2_37/A DFFSR_81/S FILL
XFILL_9_DFFSR_171 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_0_OAI21X1_4 INVX1_4/gnd DFFSR_51/S FILL
XNAND2X1_227 AND2X2_9/B AND2X2_6/B BUFX2_6/gnd XNOR2X1_3/B DFFSR_91/S NAND2X1
XFILL_4_OAI21X1_173 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_48_DFFSR_16 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_26_DFFSR_96 INVX1_2/gnd DFFSR_1/S FILL
XFILL_2_INVX1_148 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_37_DFFSR_56 INVX1_2/gnd DFFSR_51/S FILL
XFILL_5_AND2X2_15 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_26_DFFSR_101 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_16_DFFSR_104 INVX1_4/gnd DFFSR_4/S FILL
XFILL_10_DFFSR_46 BUFX2_36/A DFFSR_6/S FILL
XFILL_5_OAI21X1_107 BUFX2_36/A DFFSR_6/S FILL
XFILL_4_DFFSR_13 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_0_INVX1_365 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_2_DFFSR_5 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_13_CLKBUF1_9 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_2_DFFSR_101 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_5_NAND2X1_221 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_45_DFFSR_63 INVX1_94/gnd DFFSR_52/S FILL
XFILL_24_0_0 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_43_DFFSR_132 INVX1_2/gnd DFFSR_51/S FILL
XFILL_33_DFFSR_135 BUFX2_43/A DFFSR_97/S FILL
XFILL_22_2_1 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_9_CLKBUF1_3 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_4_NAND3X1_119 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_23_DFFSR_138 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_4_1_0 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_1_DFFSR_60 BUFX2_37/A DFFSR_8/S FILL
XFILL_13_DFFSR_141 INVX1_94/gnd DFFSR_25/S FILL
XFILL_18_DFFSR_53 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_29_DFFSR_13 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_3_OAI21X1_203 BUFX2_35/A DFFSR_14/S FILL
XFILL_6_NAND2X1_155 BUFX2_37/A DFFSR_81/S FILL
XFILL_20_4_2 INVX1_94/gnd DFFSR_52/S FILL
XFILL_3_INVX1_292 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_2_3_1 INVX1_23/gnd DFFSR_186/S FILL
XFILL_9_DFFSR_135 BUFX2_43/A DFFSR_97/S FILL
XNAND2X1_191 AND2X2_9/A INVX1_256/A BUFX2_37/A OAI22X1_2/C DFFSR_8/S NAND2X1
XFILL_18_DFFPOSX1_12 INVX1_8/gnd DFFSR_5/S FILL
XFILL_26_DFFSR_9 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_0_5_2 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_4_OAI21X1_137 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_50_DFFSR_166 INVX1_4/gnd DFFSR_51/S FILL
XFILL_37_DFFSR_20 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_2_INVX1_112 BUFX2_43/A DFFSR_97/S FILL
XFILL_40_DFFSR_169 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_26_DFFSR_60 BUFX2_37/A DFFSR_8/S FILL
XFILL_9_DFFSR_67 INVX1_2/gnd DFFSR_51/S FILL
XFILL_30_DFFSR_172 BUFX2_37/A DFFSR_8/S FILL
XFILL_20_DFFSR_175 INVX1_23/gnd DFFSR_91/S FILL
XFILL_4_NAND2X1_251 BUFX2_35/A DFFSR_97/S FILL
XFILL_10_DFFSR_10 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_16_DFFPOSX1_3 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_10_DFFSR_178 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_0_INVX1_329 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_6_XOR2X1_14 INVX1_89/gnd DFFSR_2/S FILL
XFILL_47_DFFSR_5 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_5_NOR2X1_54 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_15_DFFPOSX1_6 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_14_DFFPOSX1_9 BUFX2_37/A DFFSR_8/S FILL
XFILL_4_INVX1_436 INVX1_89/gnd DFFSR_36/S FILL
XFILL_7_OAI21X1_2 INVX1_8/gnd DFFSR_5/S FILL
XFILL_8_DFFPOSX1_23 INVX1_23/gnd DFFSR_91/S FILL
XFILL_2_OAI21X1_233 BUFX2_36/A DFFSR_8/S FILL
XFILL_6_DFFSR_172 BUFX2_37/A DFFSR_8/S FILL
XFILL_5_NAND2X1_185 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_45_DFFSR_27 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_34_DFFSR_67 INVX1_2/gnd DFFSR_51/S FILL
XFILL_2_AND2X2_16 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_18_DFFSR_17 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_23_DFFSR_102 INVX1_8/gnd DFFSR_7/S FILL
XFILL_1_DFFSR_24 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_13_DFFSR_105 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_3_OAI21X1_167 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_3_INVX1_256 BUFX2_36/A DFFSR_8/S FILL
XFILL_2_INVX1_7 BUFX2_36/A DFFSR_8/S FILL
XFILL_6_NAND2X1_119 BUFX2_37/A DFFSR_8/S FILL
XFILL_0_NOR2X1_5 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_9_AOI21X1_44 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_42_DFFSR_74 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_8_AOI21X1_47 BUFX2_43/A DFFSR_23/S FILL
XNAND2X1_155 DFFSR_154/Q DFFSR_81/S BUFX2_37/A NAND2X1_155/Y DFFSR_81/S NAND2X1
XFILL_3_NAND2X1_281 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_4_OAI21X1_101 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_27_DFFPOSX1_31 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_50_DFFSR_130 INVX1_4/gnd DFFSR_51/S FILL
XFILL_9_DFFSR_31 BUFX2_35/A DFFSR_97/S FILL
XFILL_40_DFFSR_133 BUFX2_37/A DFFSR_81/S FILL
XFILL_26_DFFSR_24 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_30_DFFSR_136 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_15_DFFSR_64 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_6_CLKBUF1_4 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_1_OAI21X1_263 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_20_DFFSR_139 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_4_NAND2X1_215 BUFX2_43/A DFFSR_23/S FILL
XFILL_10_DFFSR_142 BUFX2_19/gnd DFFSR_54/S FILL
XINVX1_403 NOR2X1_1/B BUFX2_37/A INVX1_403/Y DFFSR_8/S INVX1
XFILL_50_DFFSR_81 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_5_NOR2X1_18 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_3_NAND3X1_113 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_0_INVX1_293 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_2_XOR2X1_1 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_13_DFFSR_3 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_5_NAND2X1_149 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_2_OAI21X1_197 INVX1_8/gnd DFFSR_7/S FILL
XFILL_6_DFFSR_78 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_34_DFFSR_31 BUFX2_35/A DFFSR_97/S FILL
XFILL_23_DFFSR_71 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_6_DFFSR_136 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_47_DFFSR_167 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_37_DFFSR_170 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_5_BUFX2_16 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_27_DFFSR_173 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_3_INVX1_220 INVX1_94/gnd DFFSR_52/S FILL
XFILL_3_OAI21X1_131 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_9_AOI22X1_8 BUFX2_43/A DFFSR_97/S FILL
XFILL_8_OAI21X1_95 INVX1_89/gnd DFFSR_36/S FILL
XFILL_17_DFFSR_176 BUFX2_16/gnd DFFSR_65/S FILL
XOAI21X1_6 DFFSR_8/S INVX1_7/Y NAND2X1_6/Y BUFX2_36/A DFFSR_6/D DFFSR_6/S OAI21X1
XFILL_7_OAI21X1_98 DFFSR_1/gnd DFFSR_9/S FILL
XNAND2X1_119 BUFX2_20/Y INVX1_387/A BUFX2_37/A OAI21X1_119/C DFFSR_8/S NAND2X1
XFILL_3_NAND2X1_245 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_3_XOR2X1_15 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_42_DFFSR_38 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_31_DFFSR_78 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_3_INVX1_72 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_1_INVX1_437 BUFX2_35/A DFFSR_97/S FILL
XFILL_21_5_0 INVX1_94/gnd DFFSR_25/S FILL
XFILL_8_AOI21X1_11 INVX1_8/gnd DFFSR_5/S FILL
XFILL_4_OAI21X1_3 INVX1_4/gnd DFFSR_51/S FILL
XFILL_3_DFFSR_173 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_7_AOI21X1_14 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_15_DFFSR_28 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_30_DFFSR_100 INVX1_23/gnd DFFSR_186/S FILL
XFILL_9_AND2X2_14 BUFX2_35/A DFFSR_97/S FILL
XFILL_6_AOI21X1_17 INVX1_8/gnd DFFSR_5/S FILL
XFILL_1_OAI21X1_227 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_7_DFFPOSX1_17 BUFX2_37/A DFFSR_8/S FILL
XFILL_5_AOI21X1_20 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_4_NAND2X1_179 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_4_DFFPOSX1_3 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_20_DFFSR_103 INVX1_8/gnd DFFSR_7/S FILL
XFILL_4_AOI21X1_23 BUFX2_5/gnd DFFSR_6/S FILL
XAOI21X1_17 AOI21X1_17/A AOI21X1_17/B INVX1_237/Y INVX1_8/gnd AOI21X1_17/Y DFFSR_5/S
+ AOI21X1
XFILL_10_DFFSR_106 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_3_DFFPOSX1_6 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_3_AOI21X1_26 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_0_INVX1_257 BUFX2_36/A DFFSR_8/S FILL
XFILL_2_DFFPOSX1_9 BUFX2_37/A DFFSR_8/S FILL
XINVX1_367 DFFSR_85/Q DFFSR_71/gnd INVX1_367/Y DFFSR_10/S INVX1
XFILL_39_DFFSR_85 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_50_DFFSR_45 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_2_OAI21X1_161 INVX1_23/gnd DFFSR_186/S FILL
XFILL_4_INVX1_364 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_2_AOI21X1_29 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_6_DFFSR_100 INVX1_23/gnd DFFSR_186/S FILL
XFILL_5_NAND2X1_113 INVX1_23/gnd DFFSR_91/S FILL
XFILL_1_AOI21X1_32 BUFX2_43/A DFFSR_23/S FILL
XFILL_17_CLKBUF1_8 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_23_DFFSR_35 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_12_DFFSR_75 INVX1_4/gnd DFFSR_51/S FILL
XFILL_6_DFFSR_42 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_0_AOI21X1_35 INVX1_94/gnd DFFSR_25/S FILL
XFILL_47_DFFSR_131 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_37_DFFSR_134 DFFSR_79/gnd DFFSR_45/S FILL
XBUFX2_20 INVX1_1/Y BUFX2_5/gnd BUFX2_20/Y DFFSR_6/S BUFX2
XFILL_14_2 BUFX2_36/A DFFSR_8/S FILL
XFILL_27_DFFSR_137 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_2_NAND2X1_275 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_47_DFFSR_92 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_3_INVX1_184 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_26_DFFPOSX1_25 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_17_DFFSR_140 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_3_CLKBUF1_5 INVX1_89/gnd DFFSR_2/S FILL
XFILL_8_OAI21X1_59 INVX1_4/gnd DFFSR_51/S FILL
XFILL_3_DFFSR_89 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_8_AND2X2_1 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_7_OAI21X1_62 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_2_NOR2X1_19 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_31_0_0 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_6_NAND2X1_80 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_20_DFFSR_82 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_0_OAI21X1_257 INVX1_2/gnd DFFSR_51/S FILL
XFILL_3_INVX1_36 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_31_DFFSR_42 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_5_NAND2X1_83 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_3_NAND2X1_209 DFFSR_71/gnd DFFSR_10/S FILL
XNAND2X1_80 BUFX2_16/Y INVX1_81/A BUFX2_17/gnd NAND2X1_80/Y DFFSR_57/S NAND2X1
XFILL_6_OAI21X1_65 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_1_INVX1_401 BUFX2_35/A DFFSR_14/S FILL
XFILL_5_OAI21X1_68 BUFX2_37/A DFFSR_81/S FILL
XFILL_29_2_1 INVX1_89/gnd DFFSR_2/S FILL
XFILL_4_NAND2X1_86 INVX1_4/gnd DFFSR_51/S FILL
XOAI21X1_65 BUFX2_24/Y INVX1_74/Y OAI21X1_65/C DFFSR_3/gnd DFFSR_65/D DFFSR_4/S OAI21X1
XFILL_2_BUFX2_27 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_2_NAND3X1_107 BUFX2_43/A DFFSR_97/S FILL
XFILL_3_NAND2X1_89 BUFX2_37/A DFFSR_8/S FILL
XFILL_3_DFFSR_137 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_4_OAI21X1_71 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_2_NAND2X1_92 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_44_DFFSR_168 BUFX2_36/A DFFSR_8/S FILL
XFILL_1_OAI21X1_191 BUFX2_37/A DFFSR_8/S FILL
XFILL_1_DFFSR_2 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_3_OAI21X1_74 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_34_DFFSR_171 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_4_NAND2X1_143 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_27_4_2 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_2_OAI21X1_77 INVX1_89/gnd DFFSR_36/S FILL
XFILL_1_NAND2X1_95 INVX1_89/gnd DFFSR_36/S FILL
XFILL_28_DFFSR_89 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_24_DFFSR_174 BUFX2_43/A DFFSR_97/S FILL
XFILL_9_3_1 BUFX2_43/A DFFSR_23/S FILL
XINVX1_331 INVX1_331/A DFFSR_5/gnd INVX1_331/Y DFFSR_2/S INVX1
XFILL_0_INVX1_221 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_0_NAND2X1_98 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_0_INVX1_83 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_1_OAI21X1_80 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_39_DFFSR_49 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_6_AOI22X1_9 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_0_OAI21X1_83 INVX1_94/gnd DFFSR_52/S FILL
XFILL_14_DFFSR_177 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_2_OAI21X1_125 BUFX2_35/A DFFSR_14/S FILL
XFILL_7_5_2 BUFX2_35/A DFFSR_97/S FILL
XFILL_4_INVX1_328 INVX1_8/gnd DFFSR_7/S FILL
XFILL_12_DFFSR_39 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_0_XOR2X1_16 INVX1_8/gnd DFFSR_5/S FILL
XFILL_1_OAI21X1_4 INVX1_4/gnd DFFSR_51/S FILL
XFILL_0_DFFSR_174 BUFX2_43/A DFFSR_97/S FILL
XFILL_2_NAND2X1_239 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_25_DFFSR_6 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_36_DFFSR_96 INVX1_2/gnd DFFSR_1/S FILL
XFILL_3_INVX1_148 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_47_DFFSR_56 INVX1_2/gnd DFFSR_51/S FILL
XFILL_6_AND2X2_15 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_27_DFFSR_101 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_8_OAI21X1_23 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_17_DFFSR_104 INVX1_4/gnd DFFSR_4/S FILL
XFILL_6_NAND2X1_44 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_7_OAI21X1_26 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_0_OAI21X1_221 BUFX2_35/A DFFSR_14/S FILL
XFILL_3_NAND2X1_173 BUFX2_35/A DFFSR_14/S FILL
XFILL_20_DFFSR_46 BUFX2_36/A DFFSR_6/S FILL
XFILL_3_DFFSR_53 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_5_NAND2X1_47 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_6_DFFPOSX1_11 INVX1_4/gnd DFFSR_4/S FILL
XFILL_6_OAI21X1_29 DFFSR_3/gnd DFFSR_65/S FILL
XNAND2X1_44 DFFSR_44/S INVX1_41/A DFFSR_71/gnd OAI21X1_44/C DFFSR_45/S NAND2X1
XFILL_1_INVX1_365 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_4_NAND2X1_50 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_5_OAI21X1_32 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_3_NAND2X1_53 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_4_OAI21X1_35 INVX1_8/gnd DFFSR_5/S FILL
XFILL_14_CLKBUF1_9 BUFX2_17/gnd DFFSR_7/S FILL
XOAI21X1_29 DFFSR_65/S INVX1_33/Y OAI21X1_29/C DFFSR_3/gnd DFFSR_29/D DFFSR_65/S OAI21X1
XFILL_3_DFFSR_101 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_15_DFFPOSX1_30 BUFX2_43/A DFFSR_97/S FILL
XFILL_3_OAI21X1_38 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_44_DFFSR_132 INVX1_2/gnd DFFSR_51/S FILL
XFILL_2_NAND2X1_56 INVX1_4/gnd DFFSR_51/S FILL
XFILL_34_DFFSR_135 BUFX2_43/A DFFSR_97/S FILL
XFILL_4_NAND2X1_107 BUFX2_36/A DFFSR_6/S FILL
XFILL_1_OAI21X1_155 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_46_DFFSR_2 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_2_OAI21X1_41 INVX1_8/gnd DFFSR_7/S FILL
XFILL_1_NAND2X1_59 INVX1_2/gnd DFFSR_1/S FILL
XFILL_24_DFFSR_138 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_10_AOI22X1_10 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_0_CLKBUF1_6 BUFX2_5/gnd DFFSR_23/S FILL
XINVX1_295 DFFSR_60/Q BUFX2_7/gnd INVX1_295/Y DFFSR_54/S INVX1
XFILL_19_7 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_0_NAND2X1_62 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_0_INVX1_185 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_14_DFFSR_141 INVX1_94/gnd DFFSR_25/S FILL
XFILL_28_DFFSR_53 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_1_OAI21X1_44 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_0_INVX1_47 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_17_DFFSR_93 INVX1_2/gnd DFFSR_51/S FILL
XFILL_39_DFFSR_13 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_4_INVX1_292 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_0_OAI21X1_47 INVX1_89/gnd DFFSR_2/S FILL
XFILL_36_2 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_1_NAND2X1_269 INVX1_4/gnd DFFSR_4/S FILL
XFILL_9_AOI22X1_13 INVX1_23/gnd DFFSR_186/S FILL
XFILL_25_DFFPOSX1_19 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_1_INVX1_4 INVX1_4/gnd DFFSR_4/S FILL
XFILL_2_NAND2X1_203 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_0_DFFSR_138 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_47_DFFSR_20 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_3_INVX1_112 BUFX2_43/A DFFSR_97/S FILL
XFILL_41_DFFSR_169 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_36_DFFSR_60 BUFX2_37/A DFFSR_8/S FILL
XFILL_1_NAND3X1_101 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_31_DFFSR_172 BUFX2_37/A DFFSR_8/S FILL
XFILL_21_DFFSR_175 INVX1_23/gnd DFFSR_91/S FILL
XFILL_0_OAI21X1_185 BUFX2_36/A DFFSR_8/S FILL
XFILL_20_DFFSR_10 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_3_DFFSR_17 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_3_NAND2X1_137 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_9_OAI21X1_240 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_11_DFFSR_178 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_5_NAND2X1_11 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_4_NAND2X1_14 BUFX2_43/A DFFSR_23/S FILL
XFILL_1_INVX1_329 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_7_XOR2X1_14 INVX1_89/gnd DFFSR_2/S FILL
XFILL_6_NOR2X1_54 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_11_OAI22X1_55 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_8_OAI21X1_2 INVX1_8/gnd DFFSR_5/S FILL
XFILL_3_NAND2X1_17 INVX1_8/gnd DFFSR_7/S FILL
XDFFPOSX1_11 INVX1_331/A CLKBUF1_13/Y DFFPOSX1_11/D INVX1_4/gnd DFFSR_4/S DFFPOSX1
XFILL_2_NAND2X1_20 INVX1_23/gnd DFFSR_186/S FILL
XFILL_7_DFFSR_172 BUFX2_37/A DFFSR_8/S FILL
XFILL_1_OAI21X1_119 BUFX2_37/A DFFSR_8/S FILL
XFILL_10_OAI22X1_58 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_44_DFFSR_67 INVX1_2/gnd DFFSR_51/S FILL
XFILL_9_NAND3X1_76 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_1_NAND2X1_23 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_8_NAND3X1_79 BUFX2_36/A DFFSR_6/S FILL
XINVX1_259 XOR2X1_7/Y BUFX2_37/A INVX1_259/Y DFFSR_81/S INVX1
XFILL_9_OAI22X1_61 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_28_DFFSR_17 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_24_DFFSR_102 INVX1_8/gnd DFFSR_7/S FILL
XFILL_17_DFFSR_57 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_0_INVX1_11 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_0_NAND2X1_26 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_0_INVX1_149 INVX1_4/gnd DFFSR_51/S FILL
XFILL_0_DFFSR_64 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_14_DFFSR_105 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_7_NAND3X1_82 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_8_OAI22X1_64 INVX1_94/gnd DFFSR_25/S FILL
XFILL_3_AND2X2_16 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_0_OAI21X1_11 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_4_INVX1_256 BUFX2_36/A DFFSR_8/S FILL
XFILL_1_NAND2X1_233 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_6_NAND3X1_85 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_28_5_0 INVX1_89/gnd DFFSR_36/S FILL
XFILL_7_OAI22X1_67 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_0_NAND3X1_131 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_5_NAND3X1_88 INVX1_94/gnd DFFSR_52/S FILL
XFILL_4_NAND3X1_91 BUFX2_43/A DFFSR_97/S FILL
XNAND3X1_85 INVX1_250/A NAND3X1_81/Y NAND3X1_84/Y BUFX2_8/gnd NAND3X1_85/Y DFFSR_10/S
+ NAND3X1
XFILL_3_NAND3X1_94 BUFX2_35/A DFFSR_97/S FILL
XFILL_0_DFFSR_102 INVX1_8/gnd DFFSR_7/S FILL
XFILL_2_NAND2X1_167 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_2_NAND3X1_97 BUFX2_35/A DFFSR_97/S FILL
XFILL_41_DFFSR_133 BUFX2_37/A DFFSR_81/S FILL
XFILL_8_DFFSR_71 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_36_DFFSR_24 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_31_DFFSR_136 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_25_DFFSR_64 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_7_CLKBUF1_4 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_21_DFFSR_139 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_0_OAI21X1_149 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_14_DFFPOSX1_24 BUFX2_43/A DFFSR_23/S FILL
XFILL_9_OAI21X1_204 BUFX2_36/A DFFSR_6/S FILL
XFILL_11_DFFSR_142 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_3_NAND2X1_101 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_6_NOR2X1_18 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_1_INVX1_293 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_37_DFFSR_9 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_0_NAND2X1_263 INVX1_2/gnd DFFSR_51/S FILL
XFILL_10_OAI22X1_22 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_24_DFFPOSX1_13 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_44_DFFSR_31 BUFX2_35/A DFFSR_97/S FILL
XFILL_33_DFFSR_71 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_7_DFFSR_136 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_8_NAND3X1_43 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_9_OAI22X1_25 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_48_DFFSR_167 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_0_INVX1_113 INVX1_23/gnd DFFSR_91/S FILL
XINVX1_223 INVX1_223/A BUFX2_35/A INVX1_223/Y DFFSR_97/S INVX1
XFILL_7_NAND3X1_46 BUFX2_35/A DFFSR_97/S FILL
XFILL_38_DFFSR_170 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_0_DFFSR_28 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_8_OAI22X1_28 INVX1_94/gnd DFFSR_25/S FILL
XFILL_17_DFFSR_21 INVX1_2/gnd DFFSR_1/S FILL
XFILL_38_0_0 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_28_DFFSR_173 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_6_NAND3X1_49 BUFX2_37/A DFFSR_8/S FILL
XFILL_7_OAI22X1_31 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_1_NAND2X1_197 INVX1_8/gnd DFFSR_5/S FILL
XFILL_5_NAND3X1_52 BUFX2_36/A DFFSR_8/S FILL
XFILL_8_NOR3X1_2 INVX1_89/gnd DFFSR_2/S FILL
XFILL_18_DFFSR_176 BUFX2_16/gnd DFFSR_65/S FILL
XNAND3X1_49 INVX1_238/Y NAND3X1_52/B AOI21X1_27/B BUFX2_37/A NAND3X1_49/Y DFFSR_8/S
+ NAND3X1
XFILL_6_OAI22X1_34 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_36_2_1 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_4_NAND3X1_55 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_5_OAI22X1_37 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_4_XOR2X1_15 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_41_DFFSR_78 DFFSR_1/gnd DFFSR_1/S FILL
XOAI22X1_34 INVX1_323/Y OAI22X1_6/B INVX1_324/Y OAI22X1_8/D BUFX2_16/gnd NOR2X1_26/A
+ DFFSR_11/S OAI22X1
XFILL_8_OAI21X1_234 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_2_INVX1_437 BUFX2_35/A DFFSR_97/S FILL
XFILL_4_OAI22X1_40 BUFX2_37/A DFFSR_8/S FILL
XFILL_3_NAND3X1_58 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_34_4_2 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_2_NAND2X1_131 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_5_OAI21X1_3 INVX1_4/gnd DFFSR_51/S FILL
XDFFSR_176 DFFSR_176/Q DFFSR_3/CLK DFFSR_183/R DFFSR_65/S DFFSR_176/D BUFX2_16/gnd
+ DFFSR_65/S DFFSR
XFILL_4_DFFSR_173 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_14_DFFSR_68 BUFX2_35/A DFFSR_14/S FILL
XFILL_25_DFFSR_28 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_3_OAI22X1_43 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_2_NAND3X1_61 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_8_DFFSR_35 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_31_DFFSR_100 INVX1_23/gnd DFFSR_186/S FILL
XFILL_1_NAND3X1_64 BUFX2_35/A DFFSR_14/S FILL
XFILL_2_OAI22X1_46 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_0_OAI21X1_113 INVX1_23/gnd DFFSR_91/S FILL
XFILL_0_NAND3X1_67 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_1_OAI22X1_49 INVX1_94/gnd DFFSR_25/S FILL
XFILL_21_DFFSR_103 INVX1_8/gnd DFFSR_7/S FILL
XFILL_1_XOR2X1_5 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_9_OAI21X1_168 BUFX2_36/A DFFSR_6/S FILL
XFILL_0_OAI22X1_52 INVX1_94/gnd DFFSR_25/S FILL
XFILL_0_AND2X2_17 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_11_DFFSR_106 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_1_INVX1_257 BUFX2_36/A DFFSR_8/S FILL
XFILL_49_DFFSR_85 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_7_DFFSR_100 INVX1_23/gnd DFFSR_186/S FILL
XFILL_0_NAND2X1_227 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_18_CLKBUF1_8 BUFX2_5/gnd DFFSR_6/S FILL
XINVX1_69 DFFSR_61/Q BUFX2_36/A INVX1_69/Y DFFSR_8/S INVX1
XFILL_33_DFFSR_35 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_5_DFFSR_82 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_22_DFFSR_75 INVX1_4/gnd DFFSR_51/S FILL
XFILL_48_DFFSR_131 DFFSR_1/gnd DFFSR_1/S FILL
XINVX1_187 BUFX2_6/Y INVX1_23/gnd INVX1_187/Y DFFSR_186/S INVX1
XFILL_38_DFFSR_134 DFFSR_79/gnd DFFSR_45/S FILL
XCLKBUF1_8 DFFSR_149/Q BUFX2_5/gnd INVX1_172/A DFFSR_6/S CLKBUF1
XFILL_4_BUFX2_20 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_7_NAND3X1_10 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_28_DFFSR_137 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_1_NAND2X1_161 INVX1_23/gnd DFFSR_186/S FILL
XFILL_4_INVX1_184 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_6_NAND3X1_13 INVX1_94/gnd DFFSR_25/S FILL
XFILL_18_DFFSR_140 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_4_CLKBUF1_5 INVX1_89/gnd DFFSR_2/S FILL
XFILL_7_OAI21X1_264 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_5_NAND3X1_16 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_24_DFFSR_3 DFFSR_3/gnd DFFSR_4/S FILL
XNAND3X1_13 INVX1_224/Y NAND3X1_9/Y AOI21X1_9/B INVX1_94/gnd AOI22X1_4/B DFFSR_25/S
+ NAND3X1
XFILL_9_NAND3X1_114 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_4_NAND3X1_19 INVX1_8/gnd DFFSR_5/S FILL
XFILL_30_DFFSR_82 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_2_INVX1_76 INVX1_2/gnd DFFSR_1/S FILL
XFILL_41_DFFSR_42 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_13_DFFPOSX1_18 BUFX2_37/A DFFSR_8/S FILL
XFILL_3_NAND3X1_22 BUFX2_37/A DFFSR_81/S FILL
XFILL_3_NOR2X1_19 BUFX2_8/gnd DFFSR_10/S FILL
XDFFSR_140 DFFSR_140/Q CLKBUF1_9/Y DFFSR_137/R DFFSR_10/S DFFSR_140/D DFFSR_71/gnd
+ DFFSR_10/S DFFSR
XFILL_2_INVX1_401 BUFX2_35/A DFFSR_14/S FILL
XFILL_2_NAND3X1_25 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_8_OAI21X1_198 INVX1_8/gnd DFFSR_7/S FILL
XFILL_1_NAND3X1_28 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_4_DFFSR_137 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_14_DFFSR_32 INVX1_2/gnd DFFSR_1/S FILL
XFILL_2_OAI22X1_10 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_45_DFFSR_168 BUFX2_36/A DFFSR_8/S FILL
XFILL_0_NAND3X1_31 INVX1_94/gnd DFFSR_52/S FILL
XFILL_1_OAI22X1_13 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_35_DFFSR_171 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_9_OAI21X1_132 INVX1_4/gnd DFFSR_4/S FILL
XFILL_0_OAI22X1_16 INVX1_4/gnd DFFSR_4/S FILL
XFILL_38_DFFSR_89 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_25_DFFSR_174 BUFX2_43/A DFFSR_97/S FILL
XFILL_1_INVX1_221 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_49_DFFSR_49 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_7_AOI22X1_9 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_15_DFFSR_177 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_10_0_1 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_0_NAND2X1_191 BUFX2_37/A DFFSR_8/S FILL
XFILL_3_DFFPOSX1_29 DFFSR_1/gnd DFFSR_9/S FILL
XDFFSR_86 INVX1_97/A CLKBUF1_5/Y DFFSR_84/R DFFSR_9/S DFFSR_86/D DFFSR_1/gnd DFFSR_9/S
+ DFFSR
XINVX1_33 INVX1_33/A DFFSR_3/gnd INVX1_33/Y DFFSR_65/S INVX1
XFILL_5_DFFSR_46 BUFX2_36/A DFFSR_6/S FILL
XFILL_22_DFFSR_39 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_11_DFFSR_79 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_1_XOR2X1_16 INVX1_8/gnd DFFSR_5/S FILL
XFILL_2_OAI21X1_4 INVX1_4/gnd DFFSR_51/S FILL
XFILL_1_3 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_1_DFFSR_174 BUFX2_43/A DFFSR_97/S FILL
XFILL_0_INVX1_1 BUFX2_37/A DFFSR_81/S FILL
XINVX1_151 DFFSR_134/Q DFFSR_79/gnd INVX1_151/Y DFFSR_36/S INVX1
XFILL_1_NAND2X1_125 BUFX2_35/A DFFSR_14/S FILL
XFILL_15_XOR2X1_9 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_7_OAI21X1_228 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_28_DFFSR_101 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_46_DFFSR_96 INVX1_2/gnd DFFSR_1/S FILL
XFILL_18_DFFSR_104 INVX1_4/gnd DFFSR_4/S FILL
XFILL_7_AND2X2_15 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_7_AND2X2_5 BUFX2_37/A DFFSR_81/S FILL
XFILL_30_DFFSR_46 BUFX2_36/A DFFSR_6/S FILL
XFILL_2_INVX1_40 INVX1_8/gnd DFFSR_5/S FILL
XFILL_19_DFFSR_86 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_2_DFFSR_93 INVX1_2/gnd DFFSR_51/S FILL
XFILL_8_OAI21X1_162 INVX1_23/gnd DFFSR_91/S FILL
XFILL_2_INVX1_365 DFFSR_79/gnd DFFSR_45/S FILL
XDFFSR_104 INVX1_392/A CLKBUF1_5/Y DFFSR_97/R DFFSR_4/S DFFSR_104/D INVX1_4/gnd DFFSR_4/S
+ DFFSR
XFILL_15_CLKBUF1_9 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_4_DFFSR_101 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_1_BUFX2_31 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_45_DFFSR_132 INVX1_2/gnd DFFSR_51/S FILL
XFILL_35_DFFSR_135 BUFX2_43/A DFFSR_97/S FILL
XFILL_35_5_0 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_25_DFFSR_138 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_1_CLKBUF1_6 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_1_INVX1_185 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_15_DFFSR_141 INVX1_94/gnd DFFSR_25/S FILL
XFILL_23_4 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_38_DFFSR_53 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_27_DFFSR_93 INVX1_2/gnd DFFSR_51/S FILL
XFILL_49_DFFSR_13 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_0_NAND2X1_155 BUFX2_37/A DFFSR_81/S FILL
XFILL_11_DFFSR_43 INVX1_94/gnd DFFSR_25/S FILL
XFILL_5_DFFSR_10 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_6_OAI21X1_258 INVX1_2/gnd DFFSR_51/S FILL
XDFFSR_50 INVX1_57/A DFFSR_15/CLK DFFSR_54/R DFFSR_11/S DFFSR_50/D DFFSR_73/gnd DFFSR_11/S
+ DFFSR
XFILL_0_NOR2X1_20 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_8_NAND3X1_108 BUFX2_37/A DFFSR_81/S FILL
XINVX1_115 INVX1_376/A BUFX2_17/gnd INVX1_115/Y DFFSR_57/S INVX1
XFILL_12_DFFPOSX1_12 INVX1_8/gnd DFFSR_5/S FILL
XFILL_1_DFFSR_138 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_42_DFFSR_169 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_46_DFFSR_60 BUFX2_37/A DFFSR_8/S FILL
XFILL_7_OAI21X1_192 BUFX2_37/A DFFSR_81/S FILL
XFILL_32_DFFSR_172 BUFX2_37/A DFFSR_8/S FILL
XFILL_22_DFFSR_175 INVX1_23/gnd DFFSR_91/S FILL
XFILL_30_DFFSR_10 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_2_DFFSR_57 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_19_DFFSR_50 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_12_DFFSR_178 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_2_INVX1_329 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_8_XOR2X1_14 INVX1_89/gnd DFFSR_2/S FILL
XFILL_8_OAI21X1_126 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_2_DFFPOSX1_23 INVX1_23/gnd DFFSR_91/S FILL
XFILL_36_DFFSR_6 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_8_DFFSR_172 BUFX2_37/A DFFSR_8/S FILL
XFILL_45_0_0 INVX1_2/gnd DFFSR_1/S FILL
XFILL_38_DFFSR_17 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_25_DFFSR_102 INVX1_8/gnd DFFSR_7/S FILL
XFILL_27_DFFSR_57 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_43_2_1 INVX1_4/gnd DFFSR_51/S FILL
XFILL_1_INVX1_149 INVX1_4/gnd DFFSR_51/S FILL
XFILL_15_DFFSR_105 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_16_DFFSR_97 BUFX2_35/A DFFSR_97/S FILL
XFILL_4_AND2X2_16 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_6_OAI21X1_222 DFFSR_89/gnd DFFSR_92/S FILL
XDFFSR_14 DFFSR_14/Q INVX1_1/A DFFSR_9/R DFFSR_14/S DFFSR_14/D BUFX2_35/A DFFSR_14/S
+ DFFSR
XFILL_0_NAND2X1_119 BUFX2_37/A DFFSR_8/S FILL
XFILL_41_4_2 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_1_DFFSR_102 INVX1_8/gnd DFFSR_7/S FILL
XOAI21X1_258 DFFSR_166/S INVX1_421/Y NAND2X1_269/Y INVX1_2/gnd DFFSR_190/D DFFSR_51/S
+ OAI21X1
XFILL_7_OAI21X1_156 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_42_DFFSR_133 BUFX2_37/A DFFSR_81/S FILL
XFILL_21_DFFPOSX1_31 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_32_DFFSR_136 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_46_DFFSR_24 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_35_DFFSR_64 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_8_CLKBUF1_4 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_22_DFFSR_139 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_19_DFFSR_14 BUFX2_35/A DFFSR_14/S FILL
XFILL_12_DFFSR_142 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_2_DFFSR_21 INVX1_2/gnd DFFSR_1/S FILL
XFILL_2_INVX1_293 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_1_NOR2X1_2 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_45_4 INVX1_2/gnd DFFSR_51/S FILL
XFILL_43_DFFSR_71 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_8_DFFSR_136 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_5_OAI21X1_252 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_49_DFFSR_167 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_18_CLKBUF1_10 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_7_NAND3X1_102 INVX1_23/gnd DFFSR_186/S FILL
XFILL_1_INVX1_113 INVX1_23/gnd DFFSR_91/S FILL
XFILL_16_DFFSR_61 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_39_DFFSR_170 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_27_DFFSR_21 INVX1_2/gnd DFFSR_1/S FILL
XFILL_17_CLKBUF1_13 INVX1_4/gnd DFFSR_51/S FILL
XFILL_29_DFFSR_173 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_16_CLKBUF1_16 BUFX2_36/A DFFSR_6/S FILL
XFILL_6_OAI21X1_186 BUFX2_36/A DFFSR_8/S FILL
XFILL_15_CLKBUF1_19 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_19_DFFSR_176 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_14_CLKBUF1_22 INVX1_94/gnd DFFSR_25/S FILL
XFILL_3_DFFSR_9 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_13_CLKBUF1_25 INVX1_23/gnd DFFSR_186/S FILL
XFILL_5_XOR2X1_15 DFFSR_79/gnd DFFSR_36/S FILL
XOAI21X1_222 NOR2X1_7/A NOR2X1_7/B XOR2X1_4/Y DFFSR_89/gnd AOI22X1_11/A DFFSR_92/S
+ OAI21X1
XFILL_6_OAI21X1_3 INVX1_4/gnd DFFSR_51/S FILL
XFILL_5_DFFSR_173 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_24_DFFSR_68 BUFX2_35/A DFFSR_14/S FILL
XFILL_3_INVX1_437 BUFX2_35/A DFFSR_97/S FILL
XFILL_35_DFFSR_28 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_7_DFFSR_75 INVX1_4/gnd DFFSR_51/S FILL
XFILL_7_OAI21X1_120 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_32_DFFSR_100 INVX1_23/gnd DFFSR_186/S FILL
XFILL_1_DFFPOSX1_17 BUFX2_37/A DFFSR_8/S FILL
XFILL_22_DFFSR_103 INVX1_8/gnd DFFSR_7/S FILL
XFILL_6_BUFX2_13 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_17_0_1 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_1_AND2X2_17 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_12_DFFSR_106 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_2_INVX1_257 BUFX2_36/A DFFSR_8/S FILL
XFILL_15_2_2 BUFX2_37/A DFFSR_81/S FILL
XFILL_6_NAND3X1_132 INVX1_8/gnd DFFSR_7/S FILL
XFILL_8_DFFSR_100 INVX1_23/gnd DFFSR_186/S FILL
XFILL_19_CLKBUF1_8 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_43_DFFSR_35 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_32_DFFSR_75 INVX1_4/gnd DFFSR_51/S FILL
XFILL_5_OAI21X1_216 BUFX2_35/A DFFSR_14/S FILL
XFILL_49_DFFSR_131 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_39_DFFSR_134 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_29_DFFSR_137 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_16_DFFSR_25 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_20_DFFPOSX1_25 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_6_OAI21X1_150 INVX1_94/gnd DFFSR_52/S FILL
XFILL_19_DFFSR_140 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_5_CLKBUF1_5 INVX1_89/gnd DFFSR_2/S FILL
XNOR2X1_22 NOR2X1_22/A NOR2X1_22/B BUFX2_8/gnd NOR2X1_22/Y DFFSR_25/S NOR2X1
XFILL_48_DFFSR_9 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_40_DFFSR_82 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_51_DFFSR_42 DFFSR_3/gnd DFFSR_65/S FILL
XOAI21X1_186 INVX1_216/Y INVX1_226/Y AND2X2_5/Y BUFX2_36/A NAND3X1_8/B DFFSR_8/S OAI21X1
XFILL_4_NOR2X1_19 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_6_NAND2X1_264 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_3_INVX1_401 BUFX2_35/A DFFSR_14/S FILL
XFILL_42_5_0 INVX1_4/gnd DFFSR_4/S FILL
XFILL_5_DFFSR_137 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_7_DFFSR_39 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_13_DFFSR_72 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_24_DFFSR_32 INVX1_2/gnd DFFSR_1/S FILL
XFILL_46_DFFSR_168 BUFX2_36/A DFFSR_8/S FILL
XFILL_36_DFFSR_171 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_4_OAI21X1_246 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_48_DFFSR_89 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_26_DFFSR_174 BUFX2_43/A DFFSR_97/S FILL
XFILL_0_XOR2X1_9 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_2_INVX1_221 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_8_AOI22X1_9 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_16_DFFSR_177 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_5_OAI21X1_180 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_32_DFFSR_39 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_21_DFFSR_79 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_2_XOR2X1_16 INVX1_8/gnd DFFSR_5/S FILL
XFILL_6_CLKBUF1_10 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_4_DFFSR_86 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_4_INVX1_33 DFFSR_3/gnd DFFSR_65/S FILL
XNAND3X1_132 XOR2X1_12/B XOR2X1_13/Y XOR2X1_12/A INVX1_8/gnd AND2X2_17/A DFFSR_7/S
+ NAND3X1
XFILL_5_CLKBUF1_13 INVX1_4/gnd DFFSR_51/S FILL
XFILL_3_OAI21X1_4 INVX1_4/gnd DFFSR_51/S FILL
XFILL_2_DFFSR_174 BUFX2_43/A DFFSR_97/S FILL
XFILL_4_CLKBUF1_16 BUFX2_36/A DFFSR_6/S FILL
XFILL_0_INVX1_438 DFFSR_71/gnd DFFSR_10/S FILL
XCLKBUF1_10 clk DFFSR_73/gnd CLKBUF1_10/Y DFFSR_57/S CLKBUF1
XFILL_3_CLKBUF1_19 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_3_BUFX2_24 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_29_DFFSR_101 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_2_CLKBUF1_22 INVX1_94/gnd DFFSR_25/S FILL
XFILL_6_OAI21X1_114 INVX1_89/gnd DFFSR_36/S FILL
XFILL_14_DFFSR_7 INVX1_8/gnd DFFSR_7/S FILL
XFILL_19_DFFSR_104 INVX1_4/gnd DFFSR_4/S FILL
XFILL_8_AND2X2_15 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_1_CLKBUF1_25 INVX1_23/gnd DFFSR_186/S FILL
XFILL_40_DFFSR_46 BUFX2_36/A DFFSR_6/S FILL
XFILL_1_INVX1_80 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_29_DFFSR_86 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_0_DFFPOSX1_11 INVX1_4/gnd DFFSR_4/S FILL
XFILL_6_NAND2X1_228 INVX1_23/gnd DFFSR_91/S FILL
XOAI21X1_150 DFFSR_52/S INVX1_174/Y NAND2X1_150/Y INVX1_94/gnd DFFSR_150/D DFFSR_52/S
+ OAI21X1
XFILL_3_INVX1_365 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_13_DFFSR_36 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_16_CLKBUF1_9 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_5_DFFSR_101 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_5_NAND3X1_126 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_46_DFFSR_132 INVX1_2/gnd DFFSR_51/S FILL
XNAND2X1_264 DFFSR_186/S DFFSR_161/Q DFFSR_89/gnd OAI21X1_253/C DFFSR_186/S NAND2X1
XFILL_36_DFFSR_135 BUFX2_43/A DFFSR_97/S FILL
XFILL_10_6 BUFX2_43/A DFFSR_23/S FILL
XFILL_4_OAI21X1_210 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_48_4_2 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_35_DFFSR_3 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_26_DFFSR_138 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_2_CLKBUF1_6 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_2_INVX1_185 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_16_DFFSR_141 INVX1_94/gnd DFFSR_25/S FILL
XFILL_48_DFFSR_53 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_27_1 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_37_DFFSR_93 INVX1_2/gnd DFFSR_51/S FILL
XFILL_10_DFFSR_83 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_21_DFFSR_43 INVX1_94/gnd DFFSR_25/S FILL
XFILL_19_DFFPOSX1_19 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_4_DFFSR_50 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_5_OAI21X1_144 INVX1_8/gnd DFFSR_7/S FILL
XFILL_1_NOR2X1_20 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_0_INVX1_402 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_16_3_0 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_27_DFFPOSX1_7 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_2_DFFSR_138 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_43_DFFSR_169 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_5_NAND2X1_258 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_14_5_1 BUFX2_37/A DFFSR_8/S FILL
XFILL_33_DFFSR_172 BUFX2_37/A DFFSR_8/S FILL
XFILL_23_DFFSR_175 INVX1_23/gnd DFFSR_91/S FILL
XFILL_6_AND2X2_9 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_1_DFFSR_97 BUFX2_35/A DFFSR_97/S FILL
XFILL_40_DFFSR_10 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_1_INVX1_44 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_29_DFFSR_50 DFFSR_73/gnd DFFSR_11/S FILL
XOAI21X1_114 BUFX2_22/Y INVX1_129/Y OAI21X1_114/C INVX1_89/gnd DFFSR_114/D DFFSR_36/S
+ OAI21X1
XFILL_13_DFFSR_178 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_18_DFFSR_90 INVX1_2/gnd DFFSR_1/S FILL
XFILL_9_DFFPOSX1_30 BUFX2_43/A DFFSR_97/S FILL
XFILL_6_NAND2X1_192 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_3_INVX1_329 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_9_XOR2X1_14 INVX1_89/gnd DFFSR_2/S FILL
XFILL_3_OAI21X1_240 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_0_BUFX2_35 BUFX2_35/A DFFSR_14/S FILL
XFILL_9_DFFSR_172 BUFX2_37/A DFFSR_8/S FILL
XFILL_0_OAI21X1_5 INVX1_8/gnd DFFSR_5/S FILL
XNAND2X1_228 AND2X2_9/A INVX1_246/A INVX1_23/gnd XOR2X1_7/B DFFSR_91/S NAND2X1
XFILL_4_OAI21X1_174 BUFX2_43/A DFFSR_23/S FILL
XFILL_48_DFFSR_17 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_26_DFFSR_102 INVX1_8/gnd DFFSR_7/S FILL
XFILL_2_INVX1_149 INVX1_4/gnd DFFSR_51/S FILL
XFILL_16_DFFSR_105 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_26_DFFSR_97 BUFX2_35/A DFFSR_97/S FILL
XFILL_5_AND2X2_16 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_37_DFFSR_57 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_4_DFFSR_14 BUFX2_35/A DFFSR_14/S FILL
XFILL_5_OAI21X1_108 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_10_DFFSR_47 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_2_DFFSR_6 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_0_INVX1_366 BUFX2_37/A DFFSR_81/S FILL
XFILL_2_DFFSR_102 INVX1_8/gnd DFFSR_7/S FILL
XFILL_43_DFFSR_133 BUFX2_37/A DFFSR_81/S FILL
XFILL_24_0_1 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_5_NAND2X1_222 INVX1_23/gnd DFFSR_186/S FILL
XFILL_33_DFFSR_136 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_45_DFFSR_64 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_22_2_2 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_9_CLKBUF1_4 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_4_NAND3X1_120 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_23_DFFSR_139 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_29_DFFSR_14 BUFX2_35/A DFFSR_14/S FILL
XFILL_1_DFFSR_61 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_18_DFFSR_54 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_13_DFFSR_142 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_4_1_1 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_6_NAND2X1_156 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_3_OAI21X1_204 BUFX2_36/A DFFSR_6/S FILL
XFILL_3_INVX1_293 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_2_3_2 INVX1_23/gnd DFFSR_186/S FILL
XNAND2X1_192 AND2X2_5/Y AND2X2_6/Y BUFX2_5/gnd NAND3X1_24/C DFFSR_6/S NAND2X1
XFILL_9_DFFSR_136 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_18_DFFPOSX1_13 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_50_DFFSR_167 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_4_OAI21X1_138 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_2_INVX1_113 INVX1_23/gnd DFFSR_91/S FILL
XFILL_9_DFFSR_68 BUFX2_35/A DFFSR_14/S FILL
XFILL_26_DFFSR_61 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_40_DFFSR_170 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_37_DFFSR_21 INVX1_2/gnd DFFSR_1/S FILL
XFILL_30_DFFSR_173 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_17_DFFPOSX1_1 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_4_NAND2X1_252 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_20_DFFSR_176 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_10_DFFSR_11 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_16_DFFPOSX1_4 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_10_DFFSR_179 INVX1_2/gnd DFFSR_1/S FILL
XFILL_15_DFFPOSX1_7 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_0_INVX1_330 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_6_XOR2X1_15 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_47_DFFSR_6 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_7_OAI21X1_3 INVX1_4/gnd DFFSR_51/S FILL
XFILL_2_OAI21X1_234 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_6_DFFSR_173 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_34_DFFSR_68 BUFX2_35/A DFFSR_14/S FILL
XFILL_4_INVX1_437 BUFX2_35/A DFFSR_97/S FILL
XFILL_8_DFFPOSX1_24 BUFX2_43/A DFFSR_23/S FILL
XFILL_5_NAND2X1_186 BUFX2_37/A DFFSR_81/S FILL
XFILL_45_DFFSR_28 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_33_DFFSR_100 INVX1_23/gnd DFFSR_186/S FILL
XFILL_1_DFFSR_25 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_23_DFFSR_103 INVX1_8/gnd DFFSR_7/S FILL
XFILL_18_DFFSR_18 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_3_OAI21X1_168 BUFX2_36/A DFFSR_6/S FILL
XFILL_2_AND2X2_17 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_13_DFFSR_106 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_3_INVX1_257 BUFX2_36/A DFFSR_8/S FILL
XFILL_2_INVX1_8 INVX1_8/gnd DFFSR_5/S FILL
XFILL_6_NAND2X1_120 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_0_NOR2X1_6 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_9_DFFSR_100 INVX1_23/gnd DFFSR_186/S FILL
XFILL_20_CLKBUF1_8 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_9_AOI21X1_45 INVX1_89/gnd DFFSR_36/S FILL
XFILL_42_DFFSR_75 INVX1_4/gnd DFFSR_51/S FILL
XNAND2X1_156 INVX1_184/A DFFSR_6/S BUFX2_5/gnd OAI21X1_156/C DFFSR_6/S NAND2X1
XFILL_8_AOI21X1_48 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_3_NAND2X1_282 INVX1_89/gnd DFFSR_2/S FILL
XFILL_4_OAI21X1_102 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_50_DFFSR_131 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_40_DFFSR_134 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_9_DFFSR_32 INVX1_2/gnd DFFSR_1/S FILL
XFILL_30_DFFSR_137 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_26_DFFSR_25 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_15_DFFSR_65 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_20_DFFSR_140 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_6_CLKBUF1_5 INVX1_89/gnd DFFSR_2/S FILL
XFILL_1_OAI21X1_264 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_4_NAND2X1_216 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_10_DFFSR_143 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_2_XOR2X1_2 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_0_INVX1_294 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_50_DFFSR_82 DFFSR_1/gnd DFFSR_9/S FILL
XINVX1_404 NOR2X1_2/A BUFX2_19/gnd INVX1_404/Y DFFSR_52/S INVX1
XFILL_5_NOR2X1_19 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_3_NAND3X1_114 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_13_DFFSR_4 INVX1_4/gnd DFFSR_4/S FILL
XFILL_2_OAI21X1_198 INVX1_8/gnd DFFSR_7/S FILL
XFILL_5_NAND2X1_150 BUFX2_37/A DFFSR_81/S FILL
XFILL_6_DFFSR_137 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_6_DFFSR_79 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_23_DFFSR_72 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_34_DFFSR_32 INVX1_2/gnd DFFSR_1/S FILL
XFILL_47_DFFSR_168 BUFX2_36/A DFFSR_8/S FILL
XFILL_37_DFFSR_171 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_27_DFFSR_174 BUFX2_43/A DFFSR_97/S FILL
XFILL_3_INVX1_221 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_5_BUFX2_17 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_3_OAI21X1_132 INVX1_4/gnd DFFSR_4/S FILL
XFILL_9_AOI22X1_9 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_17_DFFSR_177 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_8_OAI21X1_96 INVX1_4/gnd DFFSR_51/S FILL
XFILL_7_OAI21X1_99 BUFX2_43/A DFFSR_97/S FILL
XFILL_23_3_0 BUFX2_8/gnd DFFSR_10/S FILL
XOAI21X1_7 DFFSR_37/S INVX1_8/Y NAND2X1_7/Y INVX1_8/gnd DFFSR_7/D DFFSR_5/S OAI21X1
XFILL_3_INVX1_73 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_3_NAND2X1_246 INVX1_94/gnd DFFSR_25/S FILL
XFILL_42_DFFSR_39 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_31_DFFSR_79 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_3_XOR2X1_16 INVX1_8/gnd DFFSR_5/S FILL
XNAND2X1_120 BUFX2_15/Y INVX1_391/A BUFX2_16/gnd OAI21X1_120/C DFFSR_65/S NAND2X1
XFILL_21_5_1 INVX1_94/gnd DFFSR_25/S FILL
XFILL_8_AOI21X1_12 INVX1_8/gnd DFFSR_7/S FILL
XFILL_4_OAI21X1_4 INVX1_4/gnd DFFSR_51/S FILL
XFILL_3_DFFSR_174 BUFX2_43/A DFFSR_97/S FILL
XFILL_7_AOI21X1_15 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_1_INVX1_438 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_15_DFFSR_29 INVX1_4/gnd DFFSR_4/S FILL
XFILL_3_4_0 INVX1_23/gnd DFFSR_91/S FILL
XFILL_5_DFFPOSX1_1 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_6_AOI21X1_18 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_30_DFFSR_101 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_5_AOI21X1_21 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_7_DFFPOSX1_18 BUFX2_37/A DFFSR_8/S FILL
XFILL_4_NAND2X1_180 INVX1_94/gnd DFFSR_52/S FILL
XFILL_1_OAI21X1_228 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_4_DFFPOSX1_4 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_20_DFFSR_104 INVX1_4/gnd DFFSR_4/S FILL
XFILL_9_AND2X2_15 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_4_AOI21X1_24 BUFX2_43/A DFFSR_97/S FILL
XFILL_10_DFFSR_107 BUFX2_36/A DFFSR_8/S FILL
XAOI21X1_18 NAND3X1_55/Y NAND3X1_58/Y INVX1_243/A BUFX2_8/gnd AOI21X1_18/Y DFFSR_10/S
+ AOI21X1
XFILL_3_DFFPOSX1_7 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_0_INVX1_258 BUFX2_43/A DFFSR_23/S FILL
XFILL_3_AOI21X1_27 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_50_DFFSR_46 BUFX2_36/A DFFSR_6/S FILL
XINVX1_368 INVX1_368/A DFFSR_79/gnd INVX1_368/Y DFFSR_36/S INVX1
XFILL_39_DFFSR_86 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_2_AOI21X1_30 INVX1_23/gnd DFFSR_91/S FILL
XFILL_2_OAI21X1_162 INVX1_23/gnd DFFSR_91/S FILL
XFILL_1_AOI21X1_33 BUFX2_35/A DFFSR_14/S FILL
XFILL_12_DFFSR_76 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_6_DFFSR_43 INVX1_94/gnd DFFSR_25/S FILL
XFILL_23_DFFSR_36 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_5_NAND2X1_114 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_17_CLKBUF1_9 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_6_DFFSR_101 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_47_DFFSR_132 INVX1_2/gnd DFFSR_51/S FILL
XFILL_37_DFFSR_135 BUFX2_43/A DFFSR_97/S FILL
XFILL_0_AOI21X1_36 BUFX2_8/gnd DFFSR_25/S FILL
XBUFX2_21 INVX1_1/Y BUFX2_5/gnd BUFX2_21/Y DFFSR_6/S BUFX2
XFILL_14_3 BUFX2_36/A DFFSR_8/S FILL
XFILL_2_NAND2X1_276 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_27_DFFSR_138 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_3_CLKBUF1_6 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_26_DFFPOSX1_26 BUFX2_37/A DFFSR_81/S FILL
XFILL_3_INVX1_185 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_17_DFFSR_141 INVX1_94/gnd DFFSR_25/S FILL
XFILL_47_DFFSR_93 INVX1_2/gnd DFFSR_51/S FILL
XFILL_9_OAI21X1_57 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_8_OAI21X1_60 BUFX2_37/A DFFSR_81/S FILL
XFILL_8_AND2X2_2 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_20_DFFSR_83 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_3_INVX1_37 INVX1_94/gnd DFFSR_52/S FILL
XFILL_31_DFFSR_43 INVX1_94/gnd DFFSR_25/S FILL
XFILL_7_OAI21X1_63 INVX1_94/gnd DFFSR_25/S FILL
XFILL_6_NAND2X1_81 INVX1_94/gnd DFFSR_25/S FILL
XFILL_31_0_1 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_3_DFFSR_90 INVX1_2/gnd DFFSR_1/S FILL
XFILL_3_NAND2X1_210 BUFX2_35/A DFFSR_97/S FILL
XFILL_5_NAND2X1_84 BUFX2_36/A DFFSR_6/S FILL
XFILL_0_OAI21X1_258 INVX1_2/gnd DFFSR_51/S FILL
XFILL_6_OAI21X1_66 INVX1_4/gnd DFFSR_51/S FILL
XFILL_2_NOR2X1_20 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_1_INVX1_402 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_5_OAI21X1_69 BUFX2_37/A DFFSR_8/S FILL
XNAND2X1_81 DFFSR_73/Q BUFX2_19/Y INVX1_94/gnd OAI21X1_81/C DFFSR_25/S NAND2X1
XFILL_4_NAND2X1_87 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_2_BUFX2_28 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_2_NAND3X1_108 BUFX2_37/A DFFSR_81/S FILL
XFILL_29_2_2 INVX1_89/gnd DFFSR_2/S FILL
XFILL_4_OAI21X1_72 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_3_NAND2X1_90 DFFSR_1/gnd DFFSR_1/S FILL
XOAI21X1_66 BUFX2_15/Y INVX1_75/Y OAI21X1_66/C INVX1_4/gnd DFFSR_66/D DFFSR_51/S OAI21X1
XFILL_3_DFFSR_138 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_44_DFFSR_169 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_1_OAI21X1_192 BUFX2_37/A DFFSR_81/S FILL
XFILL_3_OAI21X1_75 INVX1_4/gnd DFFSR_4/S FILL
XFILL_1_DFFSR_3 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_2_NAND2X1_93 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_34_DFFSR_172 BUFX2_37/A DFFSR_8/S FILL
XFILL_4_NAND2X1_144 INVX1_8/gnd DFFSR_7/S FILL
XFILL_2_OAI21X1_78 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_1_NAND2X1_96 INVX1_4/gnd DFFSR_51/S FILL
XFILL_24_DFFSR_175 INVX1_23/gnd DFFSR_91/S FILL
XFILL_0_NAND2X1_99 BUFX2_43/A DFFSR_97/S FILL
XFILL_9_3_2 BUFX2_43/A DFFSR_23/S FILL
XFILL_1_OAI21X1_81 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_50_DFFSR_10 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_0_INVX1_222 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_0_INVX1_84 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_39_DFFSR_50 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_0_OAI21X1_84 BUFX2_5/gnd DFFSR_6/S FILL
XINVX1_332 INVX1_332/A DFFSR_5/gnd INVX1_332/Y DFFSR_2/S INVX1
XFILL_14_DFFSR_178 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_28_DFFSR_90 INVX1_2/gnd DFFSR_1/S FILL
XFILL_4_INVX1_329 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_2_OAI21X1_126 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_0_XOR2X1_17 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_12_DFFSR_40 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_1_OAI21X1_5 INVX1_8/gnd DFFSR_5/S FILL
XFILL_0_DFFSR_175 INVX1_23/gnd DFFSR_91/S FILL
XFILL_2_NAND2X1_240 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_25_DFFSR_7 INVX1_8/gnd DFFSR_7/S FILL
XFILL_27_DFFSR_102 INVX1_8/gnd DFFSR_7/S FILL
XFILL_3_INVX1_149 INVX1_4/gnd DFFSR_51/S FILL
XFILL_17_DFFSR_105 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_36_DFFSR_97 BUFX2_35/A DFFSR_97/S FILL
XFILL_6_AND2X2_16 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_47_DFFSR_57 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_8_OAI21X1_24 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_6_NAND2X1_45 INVX1_89/gnd DFFSR_36/S FILL
XFILL_7_OAI21X1_27 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_0_OAI21X1_222 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_3_NAND2X1_174 BUFX2_43/A DFFSR_97/S FILL
XFILL_3_DFFSR_54 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_6_OAI21X1_30 INVX1_89/gnd DFFSR_36/S FILL
XFILL_20_DFFSR_47 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_6_DFFPOSX1_12 INVX1_8/gnd DFFSR_5/S FILL
XFILL_5_NAND2X1_48 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_5_OAI21X1_33 BUFX2_19/gnd DFFSR_52/S FILL
XNAND2X1_45 DFFSR_36/S INVX1_42/A INVX1_89/gnd OAI21X1_45/C DFFSR_36/S NAND2X1
XFILL_4_NAND2X1_51 INVX1_2/gnd DFFSR_51/S FILL
XFILL_1_INVX1_366 BUFX2_37/A DFFSR_81/S FILL
XFILL_3_NAND2X1_54 BUFX2_7/gnd DFFSR_54/S FILL
XOAI21X1_30 DFFSR_2/S INVX1_34/Y NAND2X1_30/Y INVX1_89/gnd DFFSR_30/D DFFSR_36/S OAI21X1
XFILL_3_DFFSR_102 INVX1_8/gnd DFFSR_7/S FILL
XFILL_44_DFFSR_133 BUFX2_37/A DFFSR_81/S FILL
XFILL_4_OAI21X1_36 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_1_OAI21X1_156 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_4_NAND2X1_108 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_3_OAI21X1_39 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_34_DFFSR_136 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_2_NAND2X1_57 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_15_DFFPOSX1_31 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_46_DFFSR_3 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_1_NAND2X1_60 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_24_DFFSR_139 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_2_OAI21X1_42 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_10_AOI22X1_11 INVX1_23/gnd DFFSR_91/S FILL
XFILL_0_INVX1_186 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_39_DFFSR_14 BUFX2_35/A DFFSR_14/S FILL
XFILL_0_CLKBUF1_7 BUFX2_43/A DFFSR_97/S FILL
XFILL_28_DFFSR_54 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_19_8 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_14_DFFSR_142 BUFX2_19/gnd DFFSR_54/S FILL
XINVX1_296 DFFSR_4/Q BUFX2_8/gnd INVX1_296/Y DFFSR_25/S INVX1
XFILL_0_NAND2X1_63 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_1_OAI21X1_45 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_17_DFFSR_94 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_0_INVX1_48 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_1_NAND2X1_270 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_4_INVX1_293 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_36_3 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_0_OAI21X1_48 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_25_DFFPOSX1_20 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_9_AOI22X1_14 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_1_INVX1_5 INVX1_4/gnd DFFSR_51/S FILL
XFILL_2_NAND2X1_204 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_51_DFFSR_167 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_0_DFFSR_139 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_3_INVX1_113 INVX1_23/gnd DFFSR_91/S FILL
XFILL_36_DFFSR_61 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_41_DFFSR_170 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_47_DFFSR_21 INVX1_2/gnd DFFSR_1/S FILL
XFILL_1_NAND3X1_102 INVX1_23/gnd DFFSR_186/S FILL
XFILL_31_DFFSR_173 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_3_DFFSR_18 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_21_DFFSR_176 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_20_DFFSR_11 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_9_OAI21X1_241 BUFX2_35/A DFFSR_97/S FILL
XFILL_0_OAI21X1_186 BUFX2_36/A DFFSR_8/S FILL
XFILL_5_NAND2X1_12 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_11_DFFSR_179 INVX1_2/gnd DFFSR_1/S FILL
XFILL_3_NAND2X1_138 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_1_INVX1_330 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_7_XOR2X1_15 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_4_NAND2X1_15 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_11_OAI22X1_56 BUFX2_37/A DFFSR_8/S FILL
XDFFPOSX1_12 INVX1_332/A CLKBUF1_9/Y NAND3X1_128/Y INVX1_8/gnd DFFSR_5/S DFFPOSX1
XFILL_3_NAND2X1_18 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_8_OAI21X1_3 INVX1_4/gnd DFFSR_51/S FILL
XFILL_7_DFFSR_173 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_44_DFFSR_68 BUFX2_35/A DFFSR_14/S FILL
XFILL_10_OAI22X1_59 INVX1_8/gnd DFFSR_7/S FILL
XFILL_12_DFFSR_1 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_2_NAND2X1_21 INVX1_4/gnd DFFSR_4/S FILL
XFILL_1_OAI21X1_120 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_34_DFFSR_100 INVX1_23/gnd DFFSR_186/S FILL
XFILL_1_NAND2X1_24 DFFSR_73/gnd DFFSR_57/S FILL
XINVX1_260 INVX1_260/A DFFSR_89/gnd INVX1_260/Y DFFSR_186/S INVX1
XFILL_8_NAND3X1_80 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_0_INVX1_150 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_9_OAI22X1_62 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_0_INVX1_12 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_30_3_0 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_24_DFFSR_103 INVX1_8/gnd DFFSR_7/S FILL
XFILL_0_NAND2X1_27 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_0_DFFSR_65 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_0_OAI21X1_12 BUFX2_35/A DFFSR_14/S FILL
XFILL_7_NAND3X1_83 BUFX2_37/A DFFSR_81/S FILL
XFILL_3_AND2X2_17 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_14_DFFSR_106 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_28_DFFSR_18 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_17_DFFSR_58 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_8_OAI22X1_65 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_4_INVX1_257 BUFX2_36/A DFFSR_8/S FILL
XFILL_6_NAND3X1_86 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_7_OAI22X1_68 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_1_NAND2X1_234 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_5_NAND3X1_89 BUFX2_43/A DFFSR_23/S FILL
XFILL_28_5_1 INVX1_89/gnd DFFSR_36/S FILL
XFILL_4_NAND3X1_92 BUFX2_43/A DFFSR_23/S FILL
XNAND3X1_86 NAND3X1_55/Y NAND3X1_77/Y NAND3X1_80/Y BUFX2_19/gnd NAND3X1_86/Y DFFSR_52/S
+ NAND3X1
XFILL_0_NAND3X1_132 INVX1_8/gnd DFFSR_7/S FILL
XFILL_3_NAND3X1_95 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_0_DFFSR_103 INVX1_8/gnd DFFSR_7/S FILL
XFILL_2_NAND3X1_98 BUFX2_35/A DFFSR_14/S FILL
XFILL_2_NAND2X1_168 BUFX2_36/A DFFSR_6/S FILL
XFILL_41_DFFSR_134 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_31_DFFSR_137 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_36_DFFSR_25 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_8_DFFSR_72 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_25_DFFSR_65 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_21_DFFSR_140 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_7_CLKBUF1_5 INVX1_89/gnd DFFSR_2/S FILL
XFILL_14_DFFPOSX1_25 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_0_OAI21X1_150 INVX1_94/gnd DFFSR_52/S FILL
XFILL_11_DFFSR_143 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_3_NAND2X1_102 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_9_OAI21X1_205 BUFX2_36/A DFFSR_8/S FILL
XFILL_6_NOR2X1_19 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_1_INVX1_294 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_0_NAND2X1_264 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_10_OAI22X1_23 INVX1_89/gnd DFFSR_2/S FILL
XFILL_24_DFFPOSX1_14 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_7_DFFSR_137 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_33_DFFSR_72 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_44_DFFSR_32 INVX1_2/gnd DFFSR_1/S FILL
XFILL_8_NAND3X1_44 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_48_DFFSR_168 BUFX2_36/A DFFSR_8/S FILL
XFILL_9_OAI22X1_26 INVX1_94/gnd DFFSR_52/S FILL
XINVX1_224 INVX1_224/A BUFX2_7/gnd INVX1_224/Y DFFSR_54/S INVX1
XFILL_38_DFFSR_171 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_17_DFFSR_22 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_0_INVX1_114 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_0_DFFSR_29 INVX1_4/gnd DFFSR_4/S FILL
XFILL_7_NAND3X1_47 BUFX2_43/A DFFSR_97/S FILL
XFILL_28_DFFSR_174 BUFX2_43/A DFFSR_97/S FILL
XFILL_8_OAI22X1_29 INVX1_8/gnd DFFSR_5/S FILL
XFILL_4_INVX1_221 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_1_NAND2X1_198 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_38_0_1 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_6_NAND3X1_50 BUFX2_37/A DFFSR_81/S FILL
XFILL_7_OAI22X1_32 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_18_DFFSR_177 DFFSR_5/gnd DFFSR_5/S FILL
XNAND3X1_50 INVX1_238/A NAND3X1_53/B NAND3X1_53/C BUFX2_37/A NAND3X1_50/Y DFFSR_81/S
+ NAND3X1
XFILL_5_NAND3X1_53 BUFX2_37/A DFFSR_81/S FILL
XFILL_6_OAI22X1_35 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_36_2_2 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_4_NAND3X1_56 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_5_OAI22X1_38 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_41_DFFSR_79 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_4_XOR2X1_16 INVX1_8/gnd DFFSR_5/S FILL
XOAI22X1_35 INVX1_326/Y OAI22X1_7/B INVX1_325/Y OAI22X1_7/D BUFX2_17/gnd NOR2X1_27/A
+ DFFSR_7/S OAI22X1
XFILL_8_OAI21X1_235 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_3_NAND3X1_59 BUFX2_8/gnd DFFSR_25/S FILL
XDFFSR_177 INVX1_407/A DFFSR_3/CLK DFFSR_183/R DFFSR_5/S DFFSR_177/D DFFSR_5/gnd DFFSR_5/S
+ DFFSR
XFILL_2_NAND2X1_132 INVX1_8/gnd DFFSR_5/S FILL
XFILL_5_OAI21X1_4 INVX1_4/gnd DFFSR_51/S FILL
XFILL_4_OAI22X1_41 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_4_DFFSR_174 BUFX2_43/A DFFSR_97/S FILL
XFILL_2_NAND3X1_62 BUFX2_43/A DFFSR_23/S FILL
XFILL_14_DFFSR_69 BUFX2_43/A DFFSR_23/S FILL
XFILL_2_INVX1_438 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_8_DFFSR_36 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_25_DFFSR_29 INVX1_4/gnd DFFSR_4/S FILL
XFILL_3_OAI22X1_44 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_1_NAND3X1_65 BUFX2_35/A DFFSR_14/S FILL
XFILL_2_OAI22X1_47 BUFX2_37/A DFFSR_8/S FILL
XFILL_31_DFFSR_101 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_0_NAND3X1_68 BUFX2_35/A DFFSR_14/S FILL
XFILL_1_OAI22X1_50 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_0_OAI21X1_114 INVX1_89/gnd DFFSR_36/S FILL
XFILL_21_DFFSR_104 INVX1_4/gnd DFFSR_4/S FILL
XFILL_1_XOR2X1_6 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_9_OAI21X1_169 BUFX2_36/A DFFSR_8/S FILL
XFILL_11_DFFSR_107 BUFX2_36/A DFFSR_8/S FILL
XFILL_0_OAI22X1_53 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_1_INVX1_258 BUFX2_43/A DFFSR_23/S FILL
XFILL_49_DFFSR_86 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_0_NAND2X1_228 INVX1_23/gnd DFFSR_91/S FILL
XFILL_22_DFFSR_76 BUFX2_7/gnd DFFSR_54/S FILL
XINVX1_70 INVX1_70/A BUFX2_19/gnd INVX1_70/Y DFFSR_54/S INVX1
XFILL_5_DFFSR_83 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_33_DFFSR_36 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_18_CLKBUF1_9 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_7_DFFSR_101 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_48_DFFSR_132 INVX1_2/gnd DFFSR_51/S FILL
XINVX1_188 DFFSR_157/Q BUFX2_35/A INVX1_188/Y DFFSR_97/S INVX1
XFILL_38_DFFSR_135 BUFX2_43/A DFFSR_97/S FILL
XFILL_4_BUFX2_21 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_7_NAND3X1_11 BUFX2_19/gnd DFFSR_54/S FILL
XCLKBUF1_9 clk BUFX2_17/gnd CLKBUF1_9/Y DFFSR_7/S CLKBUF1
XFILL_28_DFFSR_138 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_7_OAI21X1_265 BUFX2_43/A DFFSR_97/S FILL
XFILL_4_CLKBUF1_6 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_6_NAND3X1_14 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_4_INVX1_185 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_18_DFFSR_141 INVX1_94/gnd DFFSR_25/S FILL
XFILL_1_NAND2X1_162 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_5_NAND3X1_17 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_24_DFFSR_4 INVX1_4/gnd DFFSR_4/S FILL
XFILL_4_NAND3X1_20 BUFX2_37/A DFFSR_8/S FILL
XFILL_2_INVX1_77 BUFX2_37/A DFFSR_81/S FILL
XFILL_30_DFFSR_83 BUFX2_19/gnd DFFSR_54/S FILL
XNAND3X1_14 NAND3X1_7/Y NAND3X1_8/Y AOI21X1_2/Y BUFX2_19/gnd NAND3X1_14/Y DFFSR_52/S
+ NAND3X1
XFILL_41_DFFSR_43 INVX1_94/gnd DFFSR_25/S FILL
XFILL_3_NAND3X1_23 BUFX2_37/A DFFSR_81/S FILL
XDFFSR_141 INVX1_159/A CLKBUF1_9/Y DFFSR_137/R DFFSR_25/S DFFSR_141/D INVX1_94/gnd
+ DFFSR_25/S DFFSR
XFILL_13_DFFPOSX1_19 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_3_NOR2X1_20 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_2_INVX1_402 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_2_NAND3X1_26 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_8_OAI21X1_199 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_1_NAND3X1_29 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_14_DFFSR_33 INVX1_94/gnd DFFSR_52/S FILL
XFILL_2_OAI22X1_11 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_4_DFFSR_138 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_45_DFFSR_169 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_0_NAND3X1_32 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_35_DFFSR_172 BUFX2_37/A DFFSR_8/S FILL
XFILL_1_OAI22X1_14 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_25_DFFSR_175 INVX1_23/gnd DFFSR_91/S FILL
XFILL_9_OAI21X1_133 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_0_OAI22X1_17 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_49_DFFSR_50 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_1_INVX1_222 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_15_DFFSR_178 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_38_DFFSR_90 INVX1_2/gnd DFFSR_1/S FILL
XFILL_3_DFFPOSX1_30 BUFX2_43/A DFFSR_97/S FILL
XFILL_0_NAND2X1_192 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_10_0_2 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_1_XOR2X1_17 BUFX2_19/gnd DFFSR_52/S FILL
XINVX1_34 DFFSR_30/Q INVX1_89/gnd INVX1_34/Y DFFSR_36/S INVX1
XFILL_5_DFFSR_47 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_22_DFFSR_40 DFFSR_5/gnd DFFSR_2/S FILL
XDFFSR_87 DFFSR_87/Q CLKBUF1_4/Y DFFSR_84/R DFFSR_4/S DFFSR_87/D DFFSR_3/gnd DFFSR_4/S
+ DFFSR
XFILL_11_DFFSR_80 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_2_OAI21X1_5 INVX1_8/gnd DFFSR_5/S FILL
XINVX1_152 DFFSR_135/Q BUFX2_5/gnd INVX1_152/Y DFFSR_23/S INVX1
XFILL_0_INVX1_2 INVX1_2/gnd DFFSR_51/S FILL
XFILL_1_DFFSR_175 INVX1_23/gnd DFFSR_91/S FILL
XFILL_7_OAI21X1_229 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_28_DFFSR_102 INVX1_8/gnd DFFSR_7/S FILL
XFILL_1_NAND2X1_126 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_18_DFFSR_105 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_46_DFFSR_97 BUFX2_35/A DFFSR_97/S FILL
XFILL_7_AND2X2_16 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_7_AND2X2_6 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_2_INVX1_41 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_30_DFFSR_47 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_19_DFFSR_87 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_2_DFFSR_94 BUFX2_16/gnd DFFSR_65/S FILL
XDFFSR_105 DFFSR_105/Q CLKBUF1_7/Y DFFSR_105/R DFFSR_186/S DFFSR_105/D DFFSR_89/gnd
+ DFFSR_186/S DFFSR
XFILL_8_OAI21X1_163 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_2_INVX1_366 BUFX2_37/A DFFSR_81/S FILL
XFILL_4_DFFSR_102 INVX1_8/gnd DFFSR_7/S FILL
XFILL_45_DFFSR_133 BUFX2_37/A DFFSR_81/S FILL
XFILL_1_BUFX2_32 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_37_3_0 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_35_DFFSR_136 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_35_5_1 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_25_DFFSR_139 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_1_INVX1_186 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_49_DFFSR_14 BUFX2_35/A DFFSR_14/S FILL
XFILL_1_CLKBUF1_7 BUFX2_43/A DFFSR_97/S FILL
XFILL_38_DFFSR_54 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_15_DFFSR_142 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_23_5 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_27_DFFSR_94 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_6_OAI21X1_259 INVX1_23/gnd DFFSR_186/S FILL
XFILL_0_NAND2X1_156 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_11_DFFSR_44 BUFX2_8/gnd DFFSR_10/S FILL
XDFFSR_51 INVX1_58/A DFFSR_15/CLK DFFSR_54/R DFFSR_51/S DFFSR_51/D INVX1_2/gnd DFFSR_51/S
+ DFFSR
XFILL_5_DFFSR_11 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_0_NOR2X1_21 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_8_NAND3X1_109 BUFX2_36/A DFFSR_8/S FILL
XINVX1_116 INVX1_116/A DFFSR_5/gnd INVX1_116/Y DFFSR_5/S INVX1
XFILL_12_DFFPOSX1_13 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_1_DFFSR_139 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_46_DFFSR_61 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_42_DFFSR_170 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_7_OAI21X1_193 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_32_DFFSR_173 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_2_DFFSR_58 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_22_DFFSR_176 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_30_DFFSR_11 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_12_DFFSR_179 INVX1_2/gnd DFFSR_1/S FILL
XFILL_19_DFFSR_51 INVX1_2/gnd DFFSR_51/S FILL
XFILL_8_OAI21X1_127 BUFX2_43/A DFFSR_23/S FILL
XFILL_2_INVX1_330 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_8_XOR2X1_15 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_8_DFFSR_173 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_2_DFFPOSX1_24 BUFX2_43/A DFFSR_23/S FILL
XFILL_36_DFFSR_7 INVX1_8/gnd DFFSR_7/S FILL
XFILL_45_0_1 INVX1_2/gnd DFFSR_1/S FILL
XFILL_35_DFFSR_100 INVX1_23/gnd DFFSR_186/S FILL
XFILL_1_INVX1_150 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_25_DFFSR_103 INVX1_8/gnd DFFSR_7/S FILL
XFILL_43_2_2 INVX1_4/gnd DFFSR_51/S FILL
XFILL_4_AND2X2_17 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_15_DFFSR_106 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_16_DFFSR_98 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_38_DFFSR_18 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_27_DFFSR_58 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_0_NAND2X1_120 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_6_OAI21X1_223 BUFX2_6/gnd DFFSR_91/S FILL
XDFFSR_15 DFFSR_15/Q DFFSR_15/CLK DFFSR_9/R DFFSR_15/S DFFSR_15/D INVX1_8/gnd DFFSR_7/S
+ DFFSR
XOAI21X1_259 DFFSR_91/S INVX1_422/Y OAI21X1_259/C INVX1_23/gnd DFFSR_191/D DFFSR_186/S
+ OAI21X1
XFILL_1_DFFSR_103 INVX1_8/gnd DFFSR_7/S FILL
XFILL_7_OAI21X1_157 BUFX2_35/A DFFSR_97/S FILL
XFILL_11_1_0 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_42_DFFSR_134 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_32_DFFSR_137 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_46_DFFSR_25 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_35_DFFSR_65 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_22_DFFSR_140 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_8_CLKBUF1_5 INVX1_89/gnd DFFSR_2/S FILL
XFILL_2_DFFSR_22 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_19_DFFSR_15 INVX1_8/gnd DFFSR_7/S FILL
XFILL_12_DFFSR_143 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_2_INVX1_294 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_45_5 INVX1_2/gnd DFFSR_51/S FILL
XFILL_1_NOR2X1_3 INVX1_94/gnd DFFSR_25/S FILL
XFILL_5_OAI21X1_253 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_8_DFFSR_137 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_43_DFFSR_72 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_49_DFFSR_168 BUFX2_36/A DFFSR_8/S FILL
XFILL_18_CLKBUF1_11 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_17_CLKBUF1_14 BUFX2_43/A DFFSR_23/S FILL
XFILL_39_DFFSR_171 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_16_DFFSR_62 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_27_DFFSR_22 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_1_INVX1_114 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_7_NAND3X1_103 INVX1_23/gnd DFFSR_186/S FILL
XFILL_29_DFFSR_174 BUFX2_43/A DFFSR_97/S FILL
XFILL_16_CLKBUF1_17 INVX1_94/gnd DFFSR_25/S FILL
XFILL_6_OAI21X1_187 BUFX2_37/A DFFSR_8/S FILL
XFILL_19_DFFSR_177 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_15_CLKBUF1_20 INVX1_4/gnd DFFSR_51/S FILL
XFILL_14_CLKBUF1_23 INVX1_89/gnd DFFSR_2/S FILL
XFILL_5_XOR2X1_16 INVX1_8/gnd DFFSR_5/S FILL
XFILL_23_DFFSR_1 DFFSR_1/gnd DFFSR_1/S FILL
XOAI21X1_223 AOI22X1_10/Y AOI22X1_11/Y OAI21X1_223/C BUFX2_6/gnd NAND3X1_70/A DFFSR_91/S
+ OAI21X1
XFILL_6_OAI21X1_4 INVX1_4/gnd DFFSR_51/S FILL
XFILL_24_DFFSR_69 BUFX2_43/A DFFSR_23/S FILL
XFILL_7_OAI21X1_121 BUFX2_36/A DFFSR_8/S FILL
XFILL_7_DFFSR_76 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_3_INVX1_438 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_35_DFFSR_29 INVX1_4/gnd DFFSR_4/S FILL
XFILL_5_DFFSR_174 BUFX2_43/A DFFSR_97/S FILL
XFILL_32_DFFSR_101 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_1_DFFPOSX1_18 BUFX2_37/A DFFSR_8/S FILL
XFILL_22_DFFSR_104 INVX1_4/gnd DFFSR_4/S FILL
XFILL_12_DFFSR_107 BUFX2_36/A DFFSR_8/S FILL
XFILL_6_BUFX2_14 BUFX2_37/A DFFSR_81/S FILL
XFILL_17_0_2 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_2_INVX1_258 BUFX2_43/A DFFSR_23/S FILL
XFILL_6_NAND3X1_133 INVX1_8/gnd DFFSR_5/S FILL
XFILL_32_DFFSR_76 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_43_DFFSR_36 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_19_CLKBUF1_9 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_8_DFFSR_101 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_5_OAI21X1_217 INVX1_23/gnd DFFSR_91/S FILL
XFILL_49_DFFSR_132 INVX1_2/gnd DFFSR_51/S FILL
XFILL_39_DFFSR_135 BUFX2_43/A DFFSR_97/S FILL
XFILL_16_DFFSR_26 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_29_DFFSR_138 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_5_CLKBUF1_6 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_20_DFFPOSX1_26 BUFX2_37/A DFFSR_81/S FILL
XFILL_19_DFFSR_141 INVX1_94/gnd DFFSR_25/S FILL
XFILL_6_OAI21X1_151 BUFX2_37/A DFFSR_81/S FILL
XNOR2X1_23 NOR2X1_23/A NOR2X1_23/B DFFSR_79/gnd NOR2X1_23/Y DFFSR_45/S NOR2X1
XFILL_44_3_0 INVX1_2/gnd DFFSR_51/S FILL
XOAI21X1_187 INVX1_213/Y INVX1_227/Y AND2X2_4/Y BUFX2_37/A NAND3X1_8/C DFFSR_8/S OAI21X1
XFILL_40_DFFSR_83 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_4_NOR2X1_20 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_6_NAND2X1_265 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_3_INVX1_402 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_42_5_1 INVX1_4/gnd DFFSR_4/S FILL
XFILL_24_DFFSR_33 INVX1_94/gnd DFFSR_52/S FILL
XFILL_7_DFFSR_40 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_13_DFFSR_73 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_5_DFFSR_138 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_46_DFFSR_169 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_36_DFFSR_172 BUFX2_37/A DFFSR_8/S FILL
XFILL_4_OAI21X1_247 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_26_DFFSR_175 INVX1_23/gnd DFFSR_91/S FILL
XFILL_2_INVX1_222 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_16_DFFSR_178 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_48_DFFSR_90 INVX1_2/gnd DFFSR_1/S FILL
XFILL_6_CLKBUF1_11 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_2_XOR2X1_17 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_4_INVX1_34 INVX1_89/gnd DFFSR_36/S FILL
XFILL_32_DFFSR_40 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_5_OAI21X1_181 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_4_DFFSR_87 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_21_DFFSR_80 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_5_CLKBUF1_14 BUFX2_43/A DFFSR_23/S FILL
XFILL_3_OAI21X1_5 INVX1_8/gnd DFFSR_5/S FILL
XNAND3X1_133 INVX1_435/Y XOR2X1_16/Y OAI21X1_264/Y INVX1_8/gnd NAND3X1_133/Y DFFSR_5/S
+ NAND3X1
XFILL_5_1 BUFX2_6/gnd DFFSR_91/S FILL
XCLKBUF1_11 clk BUFX2_7/gnd CLKBUF1_11/Y DFFSR_54/S CLKBUF1
XFILL_4_CLKBUF1_17 INVX1_94/gnd DFFSR_25/S FILL
XFILL_2_DFFSR_175 INVX1_23/gnd DFFSR_91/S FILL
XFILL_3_BUFX2_25 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_29_DFFSR_102 INVX1_8/gnd DFFSR_7/S FILL
XFILL_3_CLKBUF1_20 INVX1_4/gnd DFFSR_51/S FILL
XFILL_19_DFFSR_105 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_6_OAI21X1_115 BUFX2_36/A DFFSR_6/S FILL
XFILL_8_AND2X2_16 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_14_DFFSR_8 BUFX2_36/A DFFSR_8/S FILL
XFILL_2_CLKBUF1_23 INVX1_89/gnd DFFSR_2/S FILL
XFILL_40_DFFSR_47 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_1_INVX1_81 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_29_DFFSR_87 DFFSR_3/gnd DFFSR_4/S FILL
XOAI21X1_151 DFFSR_8/S INVX1_176/Y OAI21X1_151/C BUFX2_37/A DFFSR_151/D DFFSR_81/S
+ OAI21X1
XFILL_0_DFFPOSX1_12 INVX1_8/gnd DFFSR_5/S FILL
XFILL_6_NAND2X1_229 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_3_INVX1_366 BUFX2_37/A DFFSR_81/S FILL
XFILL_13_DFFSR_37 INVX1_89/gnd DFFSR_2/S FILL
XFILL_5_DFFSR_102 INVX1_8/gnd DFFSR_7/S FILL
XFILL_46_DFFSR_133 BUFX2_37/A DFFSR_81/S FILL
XFILL_5_NAND3X1_127 DFFSR_5/gnd DFFSR_2/S FILL
XNAND2X1_265 DFFSR_186/S DFFSR_162/Q DFFSR_89/gnd NAND2X1_265/Y DFFSR_186/S NAND2X1
XFILL_36_DFFSR_136 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_10_7 BUFX2_43/A DFFSR_23/S FILL
XFILL_4_OAI21X1_211 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_35_DFFSR_4 INVX1_4/gnd DFFSR_4/S FILL
XFILL_26_DFFSR_139 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_2_INVX1_186 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_48_DFFSR_54 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_37_DFFSR_94 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_2_CLKBUF1_7 BUFX2_43/A DFFSR_97/S FILL
XFILL_16_DFFSR_142 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_21_DFFSR_44 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_4_DFFSR_51 INVX1_2/gnd DFFSR_51/S FILL
XFILL_5_OAI21X1_145 INVX1_23/gnd DFFSR_91/S FILL
XFILL_10_DFFSR_84 BUFX2_43/A DFFSR_23/S FILL
XFILL_19_DFFPOSX1_20 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_18_1_0 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_1_NOR2X1_21 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_0_INVX1_403 BUFX2_37/A DFFSR_8/S FILL
XFILL_16_3_1 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_2_DFFSR_139 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_43_DFFSR_170 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_27_DFFPOSX1_8 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_5_NAND2X1_259 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_33_DFFSR_173 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_14_5_2 BUFX2_37/A DFFSR_8/S FILL
XFILL_1_INVX1_45 INVX1_8/gnd DFFSR_5/S FILL
XFILL_23_DFFSR_176 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_40_DFFSR_11 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_18_DFFSR_91 BUFX2_6/gnd DFFSR_91/S FILL
XOAI21X1_115 BUFX2_25/Y INVX1_130/Y NAND2X1_115/Y BUFX2_36/A DFFSR_115/D DFFSR_6/S
+ OAI21X1
XFILL_1_DFFSR_98 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_13_DFFSR_179 INVX1_2/gnd DFFSR_1/S FILL
XFILL_29_DFFSR_51 INVX1_2/gnd DFFSR_51/S FILL
XFILL_3_OAI21X1_241 BUFX2_35/A DFFSR_97/S FILL
XFILL_6_NAND2X1_193 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_3_INVX1_330 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_9_XOR2X1_15 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_9_DFFPOSX1_31 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_0_BUFX2_36 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_0_OAI21X1_6 BUFX2_36/A DFFSR_6/S FILL
XFILL_36_DFFSR_100 INVX1_23/gnd DFFSR_186/S FILL
XFILL_9_DFFSR_173 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_4_OAI21X1_175 BUFX2_6/gnd DFFSR_91/S FILL
XNAND2X1_229 AOI21X1_32/B AOI21X1_32/A BUFX2_5/gnd OR2X2_3/A DFFSR_23/S NAND2X1
XFILL_26_DFFSR_103 INVX1_8/gnd DFFSR_7/S FILL
XFILL_2_INVX1_150 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_5_AND2X2_17 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_16_DFFSR_106 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_26_DFFSR_98 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_48_DFFSR_18 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_37_DFFSR_58 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_5_OAI21X1_109 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_4_DFFSR_15 INVX1_8/gnd DFFSR_7/S FILL
XFILL_10_DFFSR_48 INVX1_4/gnd DFFSR_4/S FILL
XFILL_0_INVX1_367 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_2_DFFSR_7 INVX1_8/gnd DFFSR_7/S FILL
XFILL_24_0_2 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_43_DFFSR_134 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_2_DFFSR_103 INVX1_8/gnd DFFSR_7/S FILL
XFILL_5_NAND2X1_223 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_33_DFFSR_137 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_45_DFFSR_65 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_23_DFFSR_140 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_9_CLKBUF1_5 INVX1_89/gnd DFFSR_2/S FILL
XFILL_1_DFFSR_62 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_18_DFFSR_55 INVX1_89/gnd DFFSR_36/S FILL
XFILL_4_NAND3X1_121 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_29_DFFSR_15 INVX1_8/gnd DFFSR_7/S FILL
XFILL_4_1_2 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_3_OAI21X1_205 BUFX2_36/A DFFSR_8/S FILL
XFILL_13_DFFSR_143 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_6_NAND2X1_157 BUFX2_35/A DFFSR_97/S FILL
XFILL_3_INVX1_294 DFFSR_71/gnd DFFSR_10/S FILL
XNAND2X1_193 AND2X2_6/A AND2X2_5/B BUFX2_7/gnd NAND3X1_21/C DFFSR_81/S NAND2X1
XFILL_9_DFFSR_137 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_18_DFFPOSX1_14 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_50_DFFSR_168 BUFX2_36/A DFFSR_8/S FILL
XFILL_4_OAI21X1_139 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_9_DFFSR_69 BUFX2_43/A DFFSR_23/S FILL
XFILL_40_DFFSR_171 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_26_DFFSR_62 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_37_DFFSR_22 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_2_INVX1_114 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_30_DFFSR_174 BUFX2_43/A DFFSR_97/S FILL
XFILL_4_NAND2X1_253 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_17_DFFPOSX1_2 INVX1_89/gnd DFFSR_36/S FILL
XFILL_20_DFFSR_177 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_10_DFFSR_12 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_10_DFFSR_180 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_16_DFFPOSX1_5 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_15_DFFPOSX1_8 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_0_INVX1_331 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_6_XOR2X1_16 INVX1_8/gnd DFFSR_5/S FILL
XFILL_47_DFFSR_7 INVX1_8/gnd DFFSR_7/S FILL
XFILL_7_OAI21X1_4 INVX1_4/gnd DFFSR_51/S FILL
XFILL_2_OAI21X1_235 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_34_DFFSR_69 BUFX2_43/A DFFSR_23/S FILL
XFILL_5_NAND2X1_187 BUFX2_37/A DFFSR_8/S FILL
XFILL_8_DFFPOSX1_25 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_4_INVX1_438 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_45_DFFSR_29 INVX1_4/gnd DFFSR_4/S FILL
XFILL_6_DFFSR_174 BUFX2_43/A DFFSR_97/S FILL
XFILL_33_DFFSR_101 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_1_DFFSR_26 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_23_DFFSR_104 INVX1_4/gnd DFFSR_4/S FILL
XFILL_13_DFFSR_107 BUFX2_36/A DFFSR_8/S FILL
XFILL_18_DFFSR_19 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_3_INVX1_258 BUFX2_43/A DFFSR_23/S FILL
XFILL_2_INVX1_9 BUFX2_36/A DFFSR_6/S FILL
XFILL_3_OAI21X1_169 BUFX2_36/A DFFSR_8/S FILL
XFILL_6_NAND2X1_121 BUFX2_36/A DFFSR_8/S FILL
XFILL_0_NOR2X1_7 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_42_DFFSR_76 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_20_CLKBUF1_9 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_9_DFFSR_101 DFFSR_73/gnd DFFSR_57/S FILL
XNAND2X1_157 DFFSR_156/Q DFFSR_97/S BUFX2_35/A OAI21X1_157/C DFFSR_97/S NAND2X1
XFILL_3_NAND2X1_283 INVX1_89/gnd DFFSR_36/S FILL
XFILL_4_OAI21X1_103 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_50_DFFSR_132 INVX1_2/gnd DFFSR_51/S FILL
XFILL_40_DFFSR_135 BUFX2_43/A DFFSR_97/S FILL
XFILL_9_DFFSR_33 INVX1_94/gnd DFFSR_52/S FILL
XFILL_26_DFFSR_26 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_15_DFFSR_66 INVX1_2/gnd DFFSR_51/S FILL
XFILL_30_DFFSR_138 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_1_OAI21X1_265 BUFX2_43/A DFFSR_97/S FILL
XFILL_6_CLKBUF1_6 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_20_DFFSR_141 INVX1_94/gnd DFFSR_25/S FILL
XFILL_4_NAND2X1_217 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_10_DFFSR_144 INVX1_8/gnd DFFSR_5/S FILL
XFILL_2_XOR2X1_3 BUFX2_17/gnd DFFSR_7/S FILL
XINVX1_405 INVX1_405/A BUFX2_7/gnd INVX1_405/Y DFFSR_54/S INVX1
XFILL_0_INVX1_295 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_50_DFFSR_83 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_3_NAND3X1_115 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_13_DFFSR_5 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_5_NOR2X1_20 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_4_INVX1_402 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_2_OAI21X1_199 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_5_NAND2X1_151 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_34_DFFSR_33 INVX1_94/gnd DFFSR_52/S FILL
XFILL_6_DFFSR_80 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_23_DFFSR_73 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_6_DFFSR_138 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_47_DFFSR_169 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_37_DFFSR_172 BUFX2_37/A DFFSR_8/S FILL
XFILL_27_DFFSR_175 INVX1_23/gnd DFFSR_91/S FILL
XFILL_3_OAI21X1_133 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_25_1_0 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_5_BUFX2_18 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_8_OAI21X1_97 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_3_INVX1_222 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_17_DFFSR_178 DFFSR_1/gnd DFFSR_9/S FILL
XOAI21X1_8 DFFSR_6/S INVX1_9/Y NAND2X1_8/Y BUFX2_36/A DFFSR_8/D DFFSR_6/S OAI21X1
XFILL_23_3_1 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_34_DFFSR_1 DFFSR_1/gnd DFFSR_1/S FILL
XNAND2X1_121 DFFSR_113/Q BUFX2_20/Y BUFX2_36/A NAND2X1_121/Y DFFSR_8/S NAND2X1
XFILL_3_XOR2X1_17 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_42_DFFSR_40 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_9_AOI21X1_10 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_3_INVX1_74 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_31_DFFSR_80 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_5_2_0 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_21_5_2 INVX1_94/gnd DFFSR_25/S FILL
XFILL_4_OAI21X1_5 INVX1_8/gnd DFFSR_5/S FILL
XFILL_3_NAND2X1_247 INVX1_8/gnd DFFSR_5/S FILL
XFILL_8_AOI21X1_13 INVX1_8/gnd DFFSR_7/S FILL
XFILL_7_AOI21X1_16 BUFX2_43/A DFFSR_23/S FILL
XFILL_15_DFFSR_30 INVX1_89/gnd DFFSR_36/S FILL
XFILL_3_4_1 INVX1_23/gnd DFFSR_91/S FILL
XFILL_3_DFFSR_175 INVX1_23/gnd DFFSR_91/S FILL
XFILL_6_AOI21X1_19 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_5_DFFPOSX1_2 INVX1_89/gnd DFFSR_36/S FILL
XFILL_30_DFFSR_102 INVX1_8/gnd DFFSR_7/S FILL
XFILL_20_DFFSR_105 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_5_AOI21X1_22 BUFX2_43/A DFFSR_97/S FILL
XFILL_4_NAND2X1_181 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_1_OAI21X1_229 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_7_DFFPOSX1_19 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_4_DFFPOSX1_5 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_4_AOI21X1_25 BUFX2_43/A DFFSR_97/S FILL
XAOI21X1_19 NAND3X1_56/Y NAND3X1_57/Y NAND3X1_58/A BUFX2_19/gnd AOI21X1_19/Y DFFSR_54/S
+ AOI21X1
XFILL_3_DFFPOSX1_8 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_10_DFFSR_108 INVX1_89/gnd DFFSR_2/S FILL
XFILL_0_INVX1_259 BUFX2_37/A DFFSR_81/S FILL
XFILL_3_AOI21X1_28 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_50_DFFSR_47 DFFSR_5/gnd DFFSR_2/S FILL
XINVX1_369 DFFSR_93/Q DFFSR_5/gnd INVX1_369/Y DFFSR_2/S INVX1
XFILL_39_DFFSR_87 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_2_AOI21X1_31 INVX1_23/gnd DFFSR_186/S FILL
XFILL_5_NAND2X1_115 BUFX2_36/A DFFSR_6/S FILL
XFILL_4_INVX1_366 BUFX2_37/A DFFSR_81/S FILL
XFILL_6_DFFSR_44 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_23_DFFSR_37 INVX1_89/gnd DFFSR_2/S FILL
XFILL_12_DFFSR_77 INVX1_89/gnd DFFSR_2/S FILL
XFILL_2_OAI21X1_163 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_47_DFFSR_133 BUFX2_37/A DFFSR_81/S FILL
XFILL_1_AOI21X1_34 INVX1_94/gnd DFFSR_25/S FILL
XFILL_6_DFFSR_102 INVX1_8/gnd DFFSR_7/S FILL
XFILL_0_AOI21X1_37 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_37_DFFSR_136 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_14_4 BUFX2_36/A DFFSR_8/S FILL
XFILL_2_NAND2X1_277 DFFSR_71/gnd DFFSR_10/S FILL
XBUFX2_22 INVX1_1/Y DFFSR_5/gnd BUFX2_22/Y DFFSR_2/S BUFX2
XFILL_27_DFFSR_139 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_16_XOR2X1_7 INVX1_23/gnd DFFSR_91/S FILL
XFILL_3_INVX1_186 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_26_DFFPOSX1_27 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_9_OAI21X1_58 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_47_DFFSR_94 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_3_CLKBUF1_7 BUFX2_43/A DFFSR_97/S FILL
XFILL_8_OAI21X1_61 BUFX2_36/A DFFSR_8/S FILL
XFILL_17_DFFSR_142 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_3_DFFSR_91 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_3_INVX1_38 INVX1_94/gnd DFFSR_52/S FILL
XFILL_31_0_2 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_8_AND2X2_3 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_6_NAND2X1_82 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_7_OAI21X1_64 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_0_OAI21X1_259 INVX1_23/gnd DFFSR_186/S FILL
XFILL_3_NAND2X1_211 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_20_DFFSR_84 BUFX2_43/A DFFSR_23/S FILL
XFILL_31_DFFSR_44 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_5_NAND2X1_85 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_2_NOR2X1_21 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_6_OAI21X1_67 INVX1_2/gnd DFFSR_1/S FILL
XFILL_1_INVX1_403 BUFX2_37/A DFFSR_8/S FILL
XNAND2X1_82 BUFX2_18/Y DFFSR_74/Q DFFSR_9/gnd NAND2X1_82/Y DFFSR_9/S NAND2X1
XFILL_4_NAND2X1_88 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_5_OAI21X1_70 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_3_NAND2X1_91 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_2_NAND3X1_109 BUFX2_36/A DFFSR_8/S FILL
XOAI21X1_67 BUFX2_24/Y INVX1_76/Y NAND2X1_67/Y INVX1_2/gnd DFFSR_67/D DFFSR_1/S OAI21X1
XFILL_3_DFFSR_139 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_2_BUFX2_29 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_4_OAI21X1_73 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_44_DFFSR_170 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_1_OAI21X1_193 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_3_OAI21X1_76 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_2_NAND2X1_94 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_34_DFFSR_173 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_4_NAND2X1_145 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_1_NAND2X1_97 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_2_OAI21X1_79 INVX1_89/gnd DFFSR_36/S FILL
XFILL_1_DFFSR_4 INVX1_4/gnd DFFSR_4/S FILL
XFILL_1_OAI21X1_82 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_24_DFFSR_176 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_28_DFFSR_91 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_0_INVX1_223 BUFX2_35/A DFFSR_97/S FILL
XFILL_0_OAI21X1_85 DFFSR_79/gnd DFFSR_45/S FILL
XINVX1_333 INVX1_397/A DFFSR_5/gnd INVX1_333/Y DFFSR_2/S INVX1
XFILL_14_DFFSR_179 INVX1_2/gnd DFFSR_1/S FILL
XFILL_39_DFFSR_51 INVX1_2/gnd DFFSR_51/S FILL
XFILL_0_INVX1_85 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_50_DFFSR_11 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_2_OAI21X1_127 BUFX2_43/A DFFSR_23/S FILL
XFILL_4_INVX1_330 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_12_DFFSR_41 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_1_OAI21X1_6 BUFX2_36/A DFFSR_6/S FILL
XFILL_37_DFFSR_100 INVX1_23/gnd DFFSR_186/S FILL
XFILL_25_DFFSR_8 BUFX2_36/A DFFSR_8/S FILL
XFILL_27_DFFSR_103 INVX1_8/gnd DFFSR_7/S FILL
XFILL_2_NAND2X1_241 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_0_DFFSR_176 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_3_INVX1_150 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_8_OAI21X1_25 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_6_AND2X2_17 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_17_DFFSR_106 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_36_DFFSR_98 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_47_DFFSR_58 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_7_OAI21X1_28 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_6_NAND2X1_46 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_0_OAI21X1_223 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_6_DFFPOSX1_13 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_3_DFFSR_55 INVX1_89/gnd DFFSR_36/S FILL
XFILL_20_DFFSR_48 INVX1_4/gnd DFFSR_4/S FILL
XFILL_5_NAND2X1_49 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_3_NAND2X1_175 BUFX2_35/A DFFSR_14/S FILL
XFILL_6_OAI21X1_31 BUFX2_35/A DFFSR_97/S FILL
XNAND2X1_46 DFFSR_10/S INVX1_43/A BUFX2_8/gnd OAI21X1_46/C DFFSR_25/S NAND2X1
XOAI21X1_31 DFFSR_97/S INVX1_35/Y OAI21X1_31/C BUFX2_35/A DFFSR_31/D DFFSR_97/S OAI21X1
XFILL_4_NAND2X1_52 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_1_INVX1_367 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_5_OAI21X1_34 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_44_DFFSR_134 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_4_OAI21X1_37 INVX1_89/gnd DFFSR_2/S FILL
XFILL_3_NAND2X1_55 INVX1_89/gnd DFFSR_2/S FILL
XFILL_3_DFFSR_103 INVX1_8/gnd DFFSR_7/S FILL
XFILL_1_OAI21X1_157 BUFX2_35/A DFFSR_97/S FILL
XFILL_34_DFFSR_137 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_4_NAND2X1_109 INVX1_94/gnd DFFSR_25/S FILL
XFILL_3_OAI21X1_40 INVX1_8/gnd DFFSR_7/S FILL
XFILL_46_DFFSR_4 INVX1_4/gnd DFFSR_4/S FILL
XFILL_2_NAND2X1_58 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_1_NAND2X1_61 BUFX2_37/A DFFSR_81/S FILL
XFILL_2_OAI21X1_43 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_0_INVX1_187 INVX1_23/gnd DFFSR_186/S FILL
XFILL_10_AOI22X1_12 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_1_OAI21X1_46 BUFX2_37/A DFFSR_81/S FILL
XFILL_0_INVX1_49 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_24_DFFSR_140 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_17_DFFSR_95 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_28_DFFSR_55 INVX1_89/gnd DFFSR_36/S FILL
XFILL_39_DFFSR_15 INVX1_8/gnd DFFSR_7/S FILL
XFILL_0_NAND2X1_64 BUFX2_16/gnd DFFSR_65/S FILL
XINVX1_297 DFFSR_5/Q DFFSR_73/gnd INVX1_297/Y DFFSR_11/S INVX1
XFILL_0_CLKBUF1_8 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_14_DFFSR_143 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_1_NAND2X1_271 INVX1_89/gnd DFFSR_2/S FILL
XFILL_0_OAI21X1_49 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_25_DFFPOSX1_21 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_4_INVX1_294 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_1_INVX1_6 INVX1_8/gnd DFFSR_5/S FILL
XFILL_2_NAND2X1_205 BUFX2_36/A DFFSR_6/S FILL
XFILL_51_DFFSR_168 BUFX2_36/A DFFSR_8/S FILL
XFILL_0_DFFSR_140 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_41_DFFSR_171 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_36_DFFSR_62 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_47_DFFSR_22 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_3_INVX1_114 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_1_NAND3X1_103 INVX1_23/gnd DFFSR_186/S FILL
XFILL_31_DFFSR_174 BUFX2_43/A DFFSR_97/S FILL
XFILL_21_DFFSR_177 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_6_NAND2X1_10 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_3_DFFSR_19 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_20_DFFSR_12 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_9_OAI21X1_242 BUFX2_35/A DFFSR_97/S FILL
XFILL_0_OAI21X1_187 BUFX2_37/A DFFSR_8/S FILL
XFILL_11_DFFSR_180 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_3_NAND2X1_139 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_5_NAND2X1_13 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_4_NAND2X1_16 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_1_INVX1_331 DFFSR_5/gnd DFFSR_2/S FILL
XNAND2X1_10 DFFSR_37/S DFFSR_2/Q DFFSR_5/gnd OAI21X1_10/C DFFSR_5/S NAND2X1
XFILL_7_XOR2X1_16 INVX1_8/gnd DFFSR_5/S FILL
XDFFPOSX1_13 NOR2X1_44/A CLKBUF1_12/Y NOR2X1_44/Y BUFX2_6/gnd DFFSR_91/S DFFPOSX1
XFILL_11_OAI22X1_57 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_3_NAND2X1_19 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_8_OAI21X1_4 INVX1_4/gnd DFFSR_51/S FILL
XFILL_44_DFFSR_69 BUFX2_43/A DFFSR_23/S FILL
XFILL_1_OAI21X1_121 BUFX2_36/A DFFSR_8/S FILL
XFILL_2_NAND2X1_22 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_12_DFFSR_2 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_32_1_0 INVX1_8/gnd DFFSR_5/S FILL
XFILL_10_OAI22X1_60 INVX1_8/gnd DFFSR_5/S FILL
XFILL_7_DFFSR_174 BUFX2_43/A DFFSR_97/S FILL
XFILL_1_NAND2X1_25 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_34_DFFSR_101 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_0_NAND2X1_28 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_8_NAND3X1_81 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_9_OAI22X1_63 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_1_OAI21X1_10 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_30_3_1 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_24_DFFSR_104 INVX1_4/gnd DFFSR_4/S FILL
XFILL_14_DFFSR_107 BUFX2_36/A DFFSR_8/S FILL
XINVX1_261 INVX1_261/A BUFX2_19/gnd AND2X2_13/B DFFSR_52/S INVX1
XFILL_7_NAND3X1_84 INVX1_94/gnd DFFSR_25/S FILL
XFILL_0_INVX1_151 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_8_OAI22X1_66 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_28_DFFSR_19 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_0_DFFSR_66 INVX1_2/gnd DFFSR_51/S FILL
XFILL_17_DFFSR_59 INVX1_4/gnd DFFSR_51/S FILL
XFILL_0_OAI21X1_13 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_0_INVX1_13 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_4_INVX1_258 BUFX2_43/A DFFSR_23/S FILL
XFILL_6_NAND3X1_87 INVX1_94/gnd DFFSR_52/S FILL
XFILL_1_NAND2X1_235 INVX1_4/gnd DFFSR_51/S FILL
XFILL_5_NAND3X1_90 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_28_5_2 INVX1_89/gnd DFFSR_36/S FILL
XFILL_4_NAND3X1_93 BUFX2_5/gnd DFFSR_23/S FILL
XNAND3X1_87 AOI21X1_19/Y NAND3X1_82/Y NAND3X1_83/Y INVX1_94/gnd NAND3X1_87/Y DFFSR_52/S
+ NAND3X1
XFILL_0_NAND3X1_133 INVX1_8/gnd DFFSR_5/S FILL
XFILL_3_NAND3X1_96 BUFX2_43/A DFFSR_97/S FILL
XFILL_51_DFFSR_132 INVX1_2/gnd DFFSR_51/S FILL
XFILL_41_DFFSR_135 BUFX2_43/A DFFSR_97/S FILL
XFILL_2_NAND2X1_169 BUFX2_36/A DFFSR_8/S FILL
XFILL_0_DFFSR_104 INVX1_4/gnd DFFSR_4/S FILL
XFILL_2_NAND3X1_99 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_36_DFFSR_26 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_25_DFFSR_66 INVX1_2/gnd DFFSR_51/S FILL
XFILL_8_DFFSR_73 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_31_DFFSR_138 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_7_CLKBUF1_6 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_14_DFFPOSX1_26 BUFX2_37/A DFFSR_81/S FILL
XFILL_0_OAI21X1_151 BUFX2_37/A DFFSR_81/S FILL
XFILL_21_DFFSR_141 INVX1_94/gnd DFFSR_25/S FILL
XFILL_3_NAND2X1_103 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_11_DFFSR_144 INVX1_8/gnd DFFSR_5/S FILL
XFILL_1_INVX1_295 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_6_NOR2X1_20 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_10_OAI22X1_24 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_0_NAND2X1_265 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_24_DFFPOSX1_15 BUFX2_35/A DFFSR_14/S FILL
XFILL_44_DFFSR_33 INVX1_94/gnd DFFSR_52/S FILL
XFILL_33_DFFSR_73 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_7_DFFSR_138 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_48_DFFSR_169 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_8_NAND3X1_45 BUFX2_35/A DFFSR_97/S FILL
XFILL_17_DFFSR_23 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_38_DFFSR_172 BUFX2_37/A DFFSR_8/S FILL
XINVX1_225 NAND3X1_8/A BUFX2_19/gnd AOI22X1_3/D DFFSR_54/S INVX1
XFILL_9_OAI22X1_27 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_0_DFFSR_30 INVX1_89/gnd DFFSR_36/S FILL
XFILL_0_INVX1_115 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_28_DFFSR_175 INVX1_23/gnd DFFSR_91/S FILL
XFILL_7_NAND3X1_48 BUFX2_43/A DFFSR_23/S FILL
XFILL_1_NAND2X1_199 BUFX2_36/A DFFSR_8/S FILL
XFILL_8_OAI22X1_30 INVX1_94/gnd DFFSR_25/S FILL
XFILL_38_0_2 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_6_NAND3X1_51 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_4_INVX1_222 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_7_OAI22X1_33 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_18_DFFSR_178 DFFSR_1/gnd DFFSR_9/S FILL
XNAND3X1_51 NOR3X1_1/B NAND3X1_49/Y NAND3X1_50/Y BUFX2_7/gnd NAND3X1_51/Y DFFSR_81/S
+ NAND3X1
XFILL_5_NAND3X1_54 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_6_OAI22X1_36 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_5_OAI22X1_39 BUFX2_37/A DFFSR_8/S FILL
XFILL_4_NAND3X1_57 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_4_XOR2X1_17 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_41_DFFSR_80 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_8_OAI21X1_236 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_2_NAND2X1_133 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_3_NAND3X1_60 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_5_OAI21X1_5 INVX1_8/gnd DFFSR_5/S FILL
XFILL_4_OAI22X1_42 INVX1_8/gnd DFFSR_7/S FILL
XOAI22X1_36 INVX1_327/Y OAI22X1_8/B INVX1_328/Y OAI22X1_9/D BUFX2_17/gnd NOR2X1_27/B
+ DFFSR_57/S OAI22X1
XDFFSR_178 NAND2X1_3/B DFFSR_1/CLK DFFSR_183/R DFFSR_9/S DFFSR_178/D DFFSR_1/gnd DFFSR_9/S
+ DFFSR
XFILL_2_NAND3X1_63 BUFX2_43/A DFFSR_23/S FILL
XFILL_25_DFFSR_30 INVX1_89/gnd DFFSR_36/S FILL
XFILL_8_DFFSR_37 INVX1_89/gnd DFFSR_2/S FILL
XFILL_3_OAI22X1_45 INVX1_89/gnd DFFSR_2/S FILL
XFILL_14_DFFSR_70 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_4_DFFSR_175 INVX1_23/gnd DFFSR_91/S FILL
XFILL_1_NAND3X1_66 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_2_OAI22X1_48 BUFX2_37/A DFFSR_81/S FILL
XFILL_31_DFFSR_102 INVX1_8/gnd DFFSR_7/S FILL
XFILL_21_DFFSR_105 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_0_NAND3X1_69 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_1_OAI22X1_51 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_0_OAI21X1_115 BUFX2_36/A DFFSR_6/S FILL
XFILL_9_OAI21X1_170 INVX1_94/gnd DFFSR_25/S FILL
XFILL_0_OAI22X1_54 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_11_DFFSR_108 INVX1_89/gnd DFFSR_2/S FILL
XFILL_1_XOR2X1_7 INVX1_23/gnd DFFSR_91/S FILL
XFILL_1_INVX1_259 BUFX2_37/A DFFSR_81/S FILL
XFILL_0_DFFSR_1 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_49_DFFSR_87 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_5_DFFSR_84 BUFX2_43/A DFFSR_23/S FILL
XFILL_0_NAND2X1_229 BUFX2_5/gnd DFFSR_23/S FILL
XINVX1_71 DFFSR_63/Q INVX1_94/gnd INVX1_71/Y DFFSR_25/S INVX1
XFILL_33_DFFSR_37 INVX1_89/gnd DFFSR_2/S FILL
XFILL_48_DFFSR_133 BUFX2_37/A DFFSR_81/S FILL
XFILL_22_DFFSR_77 INVX1_89/gnd DFFSR_2/S FILL
XFILL_7_DFFSR_102 INVX1_8/gnd DFFSR_7/S FILL
XFILL_38_DFFSR_136 DFFSR_5/gnd DFFSR_5/S FILL
XINVX1_189 BUFX2_5/Y BUFX2_35/A DFFSR_157/R DFFSR_14/S INVX1
XFILL_7_NAND3X1_12 INVX1_94/gnd DFFSR_52/S FILL
XFILL_4_BUFX2_22 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_4_INVX1_186 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_6_NAND3X1_15 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_1_NAND2X1_163 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_28_DFFSR_139 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_4_CLKBUF1_7 BUFX2_43/A DFFSR_97/S FILL
XFILL_18_DFFSR_142 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_14_NOR3X1_1 INVX1_94/gnd DFFSR_52/S FILL
XFILL_5_NAND3X1_18 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_24_DFFSR_5 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_4_NAND3X1_21 BUFX2_7/gnd DFFSR_81/S FILL
XNAND3X1_15 AOI21X1_8/A AOI21X1_6/C AOI21X1_8/B BUFX2_19/gnd NAND3X1_15/Y DFFSR_52/S
+ NAND3X1
XFILL_30_DFFSR_84 BUFX2_43/A DFFSR_23/S FILL
XFILL_2_INVX1_78 BUFX2_36/A DFFSR_8/S FILL
XFILL_3_NAND3X1_24 BUFX2_37/A DFFSR_8/S FILL
XFILL_13_DFFPOSX1_20 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_41_DFFSR_44 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_3_NOR2X1_21 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_8_OAI21X1_200 BUFX2_37/A DFFSR_8/S FILL
XFILL_2_INVX1_403 BUFX2_37/A DFFSR_8/S FILL
XFILL_2_NAND3X1_27 BUFX2_37/A DFFSR_81/S FILL
XDFFSR_142 DFFSR_142/Q CLKBUF1_9/Y DFFSR_137/R DFFSR_54/S DFFSR_142/D BUFX2_19/gnd
+ DFFSR_54/S DFFSR
XFILL_14_DFFSR_34 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_4_DFFSR_139 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_45_DFFSR_170 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_1_NAND3X1_30 INVX1_94/gnd DFFSR_52/S FILL
XFILL_2_OAI22X1_12 INVX1_4/gnd DFFSR_51/S FILL
XFILL_35_DFFSR_173 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_0_NAND3X1_33 INVX1_8/gnd DFFSR_7/S FILL
XFILL_1_OAI22X1_15 INVX1_4/gnd DFFSR_4/S FILL
XFILL_0_OAI22X1_18 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_9_OAI21X1_134 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_45_DFFSR_1 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_25_DFFSR_176 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_38_DFFSR_91 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_1_INVX1_223 BUFX2_35/A DFFSR_97/S FILL
XFILL_15_DFFSR_179 INVX1_2/gnd DFFSR_1/S FILL
XFILL_49_DFFSR_51 INVX1_2/gnd DFFSR_51/S FILL
XFILL_3_DFFPOSX1_31 BUFX2_17/gnd DFFSR_57/S FILL
XINVX1_35 INVX1_35/A BUFX2_35/A INVX1_35/Y DFFSR_97/S INVX1
XFILL_0_NAND2X1_193 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_11_DFFSR_81 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_22_DFFSR_41 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_5_DFFSR_48 INVX1_4/gnd DFFSR_4/S FILL
XDFFSR_88 DFFSR_88/Q CLKBUF1_2/Y DFFSR_84/R DFFSR_4/S DFFSR_88/D DFFSR_3/gnd DFFSR_4/S
+ DFFSR
XFILL_2_OAI21X1_6 BUFX2_36/A DFFSR_6/S FILL
XFILL_38_DFFSR_100 INVX1_23/gnd DFFSR_186/S FILL
XINVX1_153 INVX1_153/A DFFSR_5/gnd INVX1_153/Y DFFSR_2/S INVX1
XFILL_1_NAND2X1_127 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_0_INVX1_3 INVX1_8/gnd DFFSR_5/S FILL
XFILL_28_DFFSR_103 INVX1_8/gnd DFFSR_7/S FILL
XFILL_1_DFFSR_176 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_7_OAI21X1_230 INVX1_23/gnd DFFSR_186/S FILL
XFILL_7_AND2X2_17 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_18_DFFSR_106 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_46_DFFSR_98 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_7_AND2X2_7 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_2_DFFSR_95 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_2_INVX1_42 INVX1_89/gnd DFFSR_36/S FILL
XFILL_30_DFFSR_48 INVX1_4/gnd DFFSR_4/S FILL
XFILL_19_DFFSR_88 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_39_1_0 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_8_OAI21X1_164 DFFSR_5/gnd DFFSR_2/S FILL
XDFFSR_106 INVX1_342/A CLKBUF1_2/Y DFFSR_105/R DFFSR_1/S DFFSR_106/D DFFSR_1/gnd DFFSR_1/S
+ DFFSR
XFILL_2_INVX1_367 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_1_BUFX2_33 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_45_DFFSR_134 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_4_DFFSR_103 INVX1_8/gnd DFFSR_7/S FILL
XFILL_37_3_1 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_35_DFFSR_137 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_35_5_2 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_1_INVX1_187 INVX1_23/gnd DFFSR_186/S FILL
XFILL_25_DFFSR_140 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_27_DFFSR_95 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_38_DFFSR_55 INVX1_89/gnd DFFSR_36/S FILL
XFILL_49_DFFSR_15 INVX1_8/gnd DFFSR_7/S FILL
XFILL_1_CLKBUF1_8 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_15_DFFSR_143 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_40_1 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_5_DFFSR_12 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_0_NAND2X1_157 BUFX2_35/A DFFSR_97/S FILL
XDFFSR_52 DFFSR_52/Q DFFSR_52/CLK DFFSR_54/R DFFSR_52/S DFFSR_52/D INVX1_94/gnd DFFSR_52/S
+ DFFSR
XFILL_6_OAI21X1_260 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_0_NOR2X1_22 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_11_DFFSR_45 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_12_DFFPOSX1_14 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_8_NAND3X1_110 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_1_DFFSR_140 DFFSR_71/gnd DFFSR_10/S FILL
XINVX1_117 INVX1_392/A INVX1_4/gnd INVX1_117/Y DFFSR_51/S INVX1
XFILL_7_OAI21X1_194 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_42_DFFSR_171 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_46_DFFSR_62 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_32_DFFSR_174 BUFX2_43/A DFFSR_97/S FILL
XFILL_22_DFFSR_177 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_30_DFFSR_12 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_19_DFFSR_52 INVX1_94/gnd DFFSR_52/S FILL
XFILL_12_DFFSR_180 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_2_DFFSR_59 INVX1_4/gnd DFFSR_51/S FILL
XFILL_8_OAI21X1_128 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_2_INVX1_331 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_8_XOR2X1_16 INVX1_8/gnd DFFSR_5/S FILL
XFILL_36_DFFSR_8 BUFX2_36/A DFFSR_8/S FILL
XFILL_2_DFFPOSX1_25 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_45_0_2 INVX1_2/gnd DFFSR_1/S FILL
XFILL_8_DFFSR_174 BUFX2_43/A DFFSR_97/S FILL
XFILL_35_DFFSR_101 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_25_DFFSR_104 INVX1_4/gnd DFFSR_4/S FILL
XFILL_16_DFFSR_99 BUFX2_35/A DFFSR_97/S FILL
XFILL_15_DFFSR_107 BUFX2_36/A DFFSR_8/S FILL
XFILL_1_INVX1_151 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_38_DFFSR_19 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_27_DFFSR_59 INVX1_4/gnd DFFSR_51/S FILL
XFILL_6_OAI21X1_224 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_0_NAND2X1_121 BUFX2_36/A DFFSR_8/S FILL
XDFFSR_16 DFFSR_16/Q DFFSR_28/CLK DFFSR_9/R DFFSR_45/S DFFSR_16/D DFFSR_71/gnd DFFSR_45/S
+ DFFSR
XFILL_42_DFFSR_135 BUFX2_43/A DFFSR_97/S FILL
XFILL_1_DFFSR_104 INVX1_4/gnd DFFSR_4/S FILL
XOAI21X1_260 XOR2X1_10/B INVX1_424/A NAND2X1_272/Y BUFX2_16/gnd XOR2X1_12/A DFFSR_11/S
+ OAI21X1
XFILL_7_OAI21X1_158 BUFX2_43/A DFFSR_97/S FILL
XFILL_11_1_1 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_46_DFFSR_26 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_35_DFFSR_66 INVX1_2/gnd DFFSR_51/S FILL
XFILL_32_DFFSR_138 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_2_DFFSR_23 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_8_CLKBUF1_6 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_22_DFFSR_141 INVX1_94/gnd DFFSR_25/S FILL
XFILL_19_DFFSR_16 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_12_DFFSR_144 INVX1_8/gnd DFFSR_5/S FILL
XFILL_2_INVX1_295 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_45_6 INVX1_2/gnd DFFSR_51/S FILL
XFILL_1_NOR2X1_4 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_5_OAI21X1_254 INVX1_23/gnd DFFSR_91/S FILL
XFILL_43_DFFSR_73 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_8_DFFSR_138 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_18_CLKBUF1_12 BUFX2_43/A DFFSR_23/S FILL
XFILL_49_DFFSR_169 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_27_DFFSR_23 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_39_DFFSR_172 BUFX2_37/A DFFSR_8/S FILL
XFILL_16_DFFSR_63 INVX1_94/gnd DFFSR_52/S FILL
XFILL_17_CLKBUF1_15 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_1_INVX1_115 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_7_NAND3X1_104 INVX1_23/gnd DFFSR_186/S FILL
XFILL_29_DFFSR_175 INVX1_23/gnd DFFSR_91/S FILL
XFILL_16_CLKBUF1_18 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_6_OAI21X1_188 INVX1_89/gnd DFFSR_2/S FILL
XFILL_15_CLKBUF1_21 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_19_DFFSR_178 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_14_CLKBUF1_24 INVX1_23/gnd DFFSR_186/S FILL
XFILL_5_XOR2X1_17 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_23_DFFSR_2 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_51_DFFSR_80 BUFX2_16/gnd DFFSR_65/S FILL
XOAI21X1_224 OR2X2_2/A AOI22X1_13/Y AOI21X1_25/Y BUFX2_6/gnd NAND3X1_70/C DFFSR_91/S
+ OAI21X1
XFILL_6_OAI21X1_5 INVX1_8/gnd DFFSR_5/S FILL
XFILL_7_OAI21X1_122 INVX1_94/gnd DFFSR_25/S FILL
XFILL_35_DFFSR_30 INVX1_89/gnd DFFSR_36/S FILL
XFILL_7_DFFSR_77 INVX1_89/gnd DFFSR_2/S FILL
XFILL_24_DFFSR_70 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_5_DFFSR_175 INVX1_23/gnd DFFSR_91/S FILL
XFILL_32_DFFSR_102 INVX1_8/gnd DFFSR_7/S FILL
XFILL_22_DFFSR_105 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_12_DFFSR_108 INVX1_89/gnd DFFSR_2/S FILL
XFILL_6_BUFX2_15 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_1_DFFPOSX1_19 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_2_INVX1_259 BUFX2_37/A DFFSR_81/S FILL
XFILL_6_NAND3X1_134 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_43_DFFSR_37 INVX1_89/gnd DFFSR_2/S FILL
XFILL_5_OAI21X1_218 INVX1_23/gnd DFFSR_186/S FILL
XFILL_49_DFFSR_133 BUFX2_37/A DFFSR_81/S FILL
XFILL_32_DFFSR_77 INVX1_89/gnd DFFSR_2/S FILL
XFILL_8_DFFSR_102 INVX1_8/gnd DFFSR_7/S FILL
XFILL_39_DFFSR_136 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_16_DFFSR_27 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_46_1_0 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_29_DFFSR_139 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_5_CLKBUF1_7 BUFX2_43/A DFFSR_97/S FILL
XFILL_6_OAI21X1_152 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_19_DFFSR_142 BUFX2_19/gnd DFFSR_54/S FILL
XNOR2X1_24 NOR2X1_24/A NOR2X1_24/B BUFX2_8/gnd NOR2X1_24/Y DFFSR_10/S NOR2X1
XFILL_20_DFFPOSX1_27 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_44_3_1 INVX1_2/gnd DFFSR_51/S FILL
XFILL_40_DFFSR_84 BUFX2_43/A DFFSR_23/S FILL
XFILL_4_NOR2X1_21 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_3_INVX1_403 BUFX2_37/A DFFSR_8/S FILL
XOAI21X1_188 AOI21X1_3/Y INVX1_230/Y INVX1_229/Y INVX1_89/gnd AOI21X1_12/A DFFSR_2/S
+ OAI21X1
XFILL_42_5_2 INVX1_4/gnd DFFSR_4/S FILL
XFILL_6_NAND2X1_266 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_7_DFFSR_41 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_24_DFFSR_34 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_13_DFFSR_74 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_5_DFFSR_139 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_46_DFFSR_170 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_36_DFFSR_173 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_4_OAI21X1_248 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_26_DFFSR_176 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_48_DFFSR_91 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_2_INVX1_223 BUFX2_35/A DFFSR_97/S FILL
XFILL_16_DFFSR_179 INVX1_2/gnd DFFSR_1/S FILL
XFILL_4_INVX1_35 BUFX2_35/A DFFSR_97/S FILL
XFILL_6_CLKBUF1_12 BUFX2_43/A DFFSR_23/S FILL
XFILL_10_4_0 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_21_DFFSR_81 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_5_OAI21X1_182 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_32_DFFSR_41 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_4_DFFSR_88 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_3_OAI21X1_6 BUFX2_36/A DFFSR_6/S FILL
XFILL_39_DFFSR_100 INVX1_23/gnd DFFSR_186/S FILL
XCLKBUF1_12 clk BUFX2_43/A CLKBUF1_12/Y DFFSR_23/S CLKBUF1
XNAND3X1_134 NOR2X1_1/B NOR2X1_1/A INVX1_438/Y DFFSR_71/gnd AOI21X1_48/A DFFSR_10/S
+ NAND3X1
XFILL_5_CLKBUF1_15 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_5_2 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_4_CLKBUF1_18 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_29_DFFSR_103 INVX1_8/gnd DFFSR_7/S FILL
XFILL_3_BUFX2_26 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_2_DFFSR_176 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_6_OAI21X1_116 INVX1_89/gnd DFFSR_2/S FILL
XFILL_8_AND2X2_17 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_3_CLKBUF1_21 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_19_DFFSR_106 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_2_CLKBUF1_24 INVX1_23/gnd DFFSR_186/S FILL
XFILL_14_DFFSR_9 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_1_INVX1_82 BUFX2_35/A DFFSR_97/S FILL
XFILL_40_DFFSR_48 INVX1_4/gnd DFFSR_4/S FILL
XFILL_29_DFFSR_88 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_0_DFFPOSX1_13 BUFX2_6/gnd DFFSR_91/S FILL
XOAI21X1_152 DFFSR_23/S INVX1_178/Y OAI21X1_152/C BUFX2_5/gnd DFFSR_152/D DFFSR_6/S
+ OAI21X1
XFILL_6_NAND2X1_230 BUFX2_36/A DFFSR_6/S FILL
XFILL_3_INVX1_367 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_46_DFFSR_134 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_5_DFFSR_103 INVX1_8/gnd DFFSR_7/S FILL
XFILL_13_DFFSR_38 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_5_NAND3X1_128 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_4_OAI21X1_212 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_36_DFFSR_137 BUFX2_7/gnd DFFSR_54/S FILL
XNAND2X1_266 DFFSR_4/S DFFSR_163/Q DFFSR_3/gnd NAND2X1_266/Y DFFSR_4/S NAND2X1
XFILL_2_INVX1_187 INVX1_23/gnd DFFSR_186/S FILL
XFILL_26_DFFSR_140 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_37_DFFSR_95 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_48_DFFSR_55 INVX1_89/gnd DFFSR_36/S FILL
XFILL_35_DFFSR_5 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_2_CLKBUF1_8 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_16_DFFSR_143 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_4_DFFSR_52 INVX1_94/gnd DFFSR_52/S FILL
XFILL_5_OAI21X1_146 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_19_DFFPOSX1_21 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_18_1_1 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_1_NOR2X1_22 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_10_DFFSR_85 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_21_DFFSR_45 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_0_0_0 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_0_INVX1_404 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_16_3_2 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_2_DFFSR_140 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_5_NAND2X1_260 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_27_DFFPOSX1_9 BUFX2_37/A DFFSR_8/S FILL
XFILL_43_DFFSR_171 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_33_DFFSR_174 BUFX2_43/A DFFSR_97/S FILL
XFILL_23_DFFSR_177 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_18_DFFSR_92 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_40_DFFSR_12 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_1_DFFSR_99 BUFX2_35/A DFFSR_97/S FILL
XFILL_29_DFFSR_52 INVX1_94/gnd DFFSR_52/S FILL
XFILL_1_INVX1_46 DFFSR_71/gnd DFFSR_45/S FILL
XOAI21X1_116 BUFX2_17/Y INVX1_131/Y NAND2X1_116/Y INVX1_89/gnd DFFSR_116/D DFFSR_2/S
+ OAI21X1
XFILL_13_DFFSR_180 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_3_OAI21X1_242 BUFX2_35/A DFFSR_97/S FILL
XFILL_6_NAND2X1_194 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_3_INVX1_331 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_9_XOR2X1_16 INVX1_8/gnd DFFSR_5/S FILL
XFILL_0_BUFX2_37 BUFX2_37/A DFFSR_81/S FILL
XFILL_0_OAI21X1_7 INVX1_8/gnd DFFSR_5/S FILL
XFILL_9_DFFSR_174 BUFX2_43/A DFFSR_97/S FILL
XNAND2X1_230 OR2X2_3/B OR2X2_3/A BUFX2_36/A AOI21X1_38/B DFFSR_6/S NAND2X1
XFILL_36_DFFSR_101 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_4_OAI21X1_176 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_26_DFFSR_104 INVX1_4/gnd DFFSR_4/S FILL
XFILL_26_DFFSR_99 BUFX2_35/A DFFSR_97/S FILL
XFILL_16_DFFSR_107 BUFX2_36/A DFFSR_8/S FILL
XFILL_2_INVX1_151 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_48_DFFSR_19 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_37_DFFSR_59 INVX1_4/gnd DFFSR_51/S FILL
XFILL_4_DFFSR_16 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_5_OAI21X1_110 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_10_DFFSR_49 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_0_INVX1_368 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_2_DFFSR_8 BUFX2_36/A DFFSR_8/S FILL
XFILL_2_DFFSR_104 INVX1_4/gnd DFFSR_4/S FILL
XFILL_43_DFFSR_135 BUFX2_43/A DFFSR_97/S FILL
XFILL_5_NAND2X1_224 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_45_DFFSR_66 INVX1_2/gnd DFFSR_51/S FILL
XFILL_33_DFFSR_138 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_9_CLKBUF1_6 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_1_INVX1_10 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_1_DFFSR_63 INVX1_94/gnd DFFSR_52/S FILL
XFILL_23_DFFSR_141 INVX1_94/gnd DFFSR_25/S FILL
XFILL_29_DFFSR_16 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_4_NAND3X1_122 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_18_DFFSR_56 INVX1_2/gnd DFFSR_51/S FILL
XFILL_3_OAI21X1_206 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_13_DFFSR_144 INVX1_8/gnd DFFSR_5/S FILL
XFILL_6_NAND2X1_158 BUFX2_35/A DFFSR_97/S FILL
XFILL_3_INVX1_295 BUFX2_7/gnd DFFSR_54/S FILL
XNAND2X1_194 BUFX2_13/Y AND2X2_6/B BUFX2_7/gnd NAND2X1_195/B DFFSR_54/S NAND2X1
XFILL_9_DFFSR_138 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_18_DFFPOSX1_15 BUFX2_35/A DFFSR_14/S FILL
XFILL_50_DFFSR_169 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_4_OAI21X1_140 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_37_DFFSR_23 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_40_DFFSR_172 BUFX2_37/A DFFSR_8/S FILL
XFILL_26_DFFSR_63 INVX1_94/gnd DFFSR_52/S FILL
XFILL_9_DFFSR_70 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_2_INVX1_115 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_30_DFFSR_175 INVX1_23/gnd DFFSR_91/S FILL
XFILL_17_DFFPOSX1_3 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_20_DFFSR_178 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_10_DFFSR_181 INVX1_23/gnd DFFSR_186/S FILL
XFILL_4_NAND2X1_254 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_16_DFFPOSX1_6 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_10_DFFSR_13 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_15_DFFPOSX1_9 BUFX2_37/A DFFSR_8/S FILL
XFILL_6_XOR2X1_17 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_0_INVX1_332 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_47_DFFSR_8 BUFX2_36/A DFFSR_8/S FILL
XFILL_7_OAI21X1_5 INVX1_8/gnd DFFSR_5/S FILL
XFILL_2_OAI21X1_236 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_8_DFFPOSX1_26 BUFX2_37/A DFFSR_81/S FILL
XFILL_45_DFFSR_30 INVX1_89/gnd DFFSR_36/S FILL
XFILL_5_NAND2X1_188 INVX1_8/gnd DFFSR_7/S FILL
XFILL_6_DFFSR_175 INVX1_23/gnd DFFSR_91/S FILL
XFILL_33_DFFSR_102 INVX1_8/gnd DFFSR_7/S FILL
XFILL_34_DFFSR_70 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_23_DFFSR_105 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_18_DFFSR_20 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_17_4_0 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_13_DFFSR_108 INVX1_89/gnd DFFSR_2/S FILL
XFILL_1_DFFSR_27 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_10_OAI22X1_1 BUFX2_36/A DFFSR_8/S FILL
XFILL_3_INVX1_259 BUFX2_37/A DFFSR_81/S FILL
XFILL_3_OAI21X1_170 INVX1_94/gnd DFFSR_25/S FILL
XFILL_6_NAND2X1_122 INVX1_94/gnd DFFSR_25/S FILL
XFILL_0_NOR2X1_8 BUFX2_43/A DFFSR_23/S FILL
XFILL_9_NOR3X1_1 INVX1_94/gnd DFFSR_52/S FILL
XNAND2X1_158 DFFSR_157/Q DFFSR_97/S BUFX2_35/A NAND2X1_158/Y DFFSR_97/S NAND2X1
XFILL_50_DFFSR_133 BUFX2_37/A DFFSR_81/S FILL
XFILL_42_DFFSR_77 INVX1_89/gnd DFFSR_2/S FILL
XFILL_3_NAND2X1_284 INVX1_8/gnd DFFSR_5/S FILL
XFILL_9_DFFSR_102 INVX1_8/gnd DFFSR_7/S FILL
XFILL_4_OAI21X1_104 INVX1_4/gnd DFFSR_51/S FILL
XFILL_40_DFFSR_136 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_26_DFFSR_27 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_9_DFFSR_34 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_15_DFFSR_67 INVX1_2/gnd DFFSR_51/S FILL
XFILL_30_DFFSR_139 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_6_CLKBUF1_7 BUFX2_43/A DFFSR_97/S FILL
XFILL_20_DFFSR_142 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_4_NAND2X1_218 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_2_XOR2X1_4 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_10_DFFSR_145 INVX1_23/gnd DFFSR_186/S FILL
XFILL_50_DFFSR_84 BUFX2_43/A DFFSR_23/S FILL
XFILL_13_DFFSR_6 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_0_INVX1_296 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_3_NAND3X1_116 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_5_NOR2X1_21 DFFSR_79/gnd DFFSR_36/S FILL
XINVX1_406 DFFSR_176/Q DFFSR_3/gnd INVX1_406/Y DFFSR_65/S INVX1
XFILL_2_OAI21X1_200 BUFX2_37/A DFFSR_8/S FILL
XFILL_5_NAND2X1_152 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_6_DFFSR_81 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_34_DFFSR_34 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_23_DFFSR_74 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_6_DFFSR_139 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_47_DFFSR_170 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_37_DFFSR_173 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_5_BUFX2_19 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_25_1_1 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_3_OAI21X1_134 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_27_DFFSR_176 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_3_INVX1_223 BUFX2_35/A DFFSR_97/S FILL
XFILL_7_0_0 BUFX2_35/A DFFSR_97/S FILL
XFILL_17_DFFSR_179 INVX1_2/gnd DFFSR_1/S FILL
XFILL_23_3_2 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_34_DFFSR_2 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_8_OAI21X1_98 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_31_DFFSR_81 BUFX2_7/gnd DFFSR_81/S FILL
XNAND2X1_122 BUFX2_19/Y INVX1_344/A INVX1_94/gnd NAND2X1_122/Y DFFSR_25/S NAND2X1
XFILL_42_DFFSR_41 BUFX2_17/gnd DFFSR_57/S FILL
XOAI21X1_9 DFFSR_9/S INVX1_11/Y NAND2X1_9/Y DFFSR_1/gnd DFFSR_9/D DFFSR_9/S OAI21X1
XFILL_3_INVX1_75 INVX1_4/gnd DFFSR_51/S FILL
XFILL_5_2_1 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_4_OAI21X1_6 BUFX2_36/A DFFSR_6/S FILL
XFILL_8_AOI21X1_14 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_3_NAND2X1_248 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_40_DFFSR_100 INVX1_23/gnd DFFSR_186/S FILL
XFILL_15_DFFSR_31 BUFX2_35/A DFFSR_97/S FILL
XFILL_7_AOI21X1_17 INVX1_8/gnd DFFSR_5/S FILL
XFILL_3_4_2 INVX1_23/gnd DFFSR_91/S FILL
XFILL_6_AOI21X1_20 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_5_DFFPOSX1_3 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_30_DFFSR_103 INVX1_8/gnd DFFSR_7/S FILL
XFILL_3_DFFSR_176 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_1_OAI21X1_230 INVX1_23/gnd DFFSR_186/S FILL
XFILL_5_AOI21X1_23 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_7_DFFPOSX1_20 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_20_DFFSR_106 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_4_DFFPOSX1_6 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_10_DFFSR_109 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_3_DFFPOSX1_9 BUFX2_37/A DFFSR_8/S FILL
XAOI21X1_20 NAND3X1_53/Y NAND3X1_52/Y NAND3X1_56/A BUFX2_7/gnd NAND3X1_83/A DFFSR_81/S
+ AOI21X1
XFILL_4_NAND2X1_182 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_0_INVX1_260 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_4_AOI21X1_26 BUFX2_5/gnd DFFSR_23/S FILL
XINVX1_370 DFFSR_125/Q BUFX2_36/A INVX1_370/Y DFFSR_8/S INVX1
XFILL_50_DFFSR_48 INVX1_4/gnd DFFSR_4/S FILL
XFILL_39_DFFSR_88 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_3_AOI21X1_29 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_2_AOI21X1_32 BUFX2_43/A DFFSR_23/S FILL
XFILL_6_DFFSR_45 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_5_NAND2X1_116 INVX1_89/gnd DFFSR_36/S FILL
XFILL_2_OAI21X1_164 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_1_AOI21X1_35 INVX1_94/gnd DFFSR_25/S FILL
XFILL_6_DFFSR_103 INVX1_8/gnd DFFSR_7/S FILL
XFILL_23_DFFSR_38 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_12_DFFSR_78 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_0_AOI21X1_38 BUFX2_36/A DFFSR_8/S FILL
XFILL_47_DFFSR_134 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_14_5 BUFX2_36/A DFFSR_8/S FILL
XFILL_37_DFFSR_137 BUFX2_7/gnd DFFSR_54/S FILL
XBUFX2_23 INVX1_1/Y BUFX2_19/gnd BUFX2_23/Y DFFSR_54/S BUFX2
XFILL_2_NAND2X1_278 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_3_INVX1_187 INVX1_23/gnd DFFSR_186/S FILL
XFILL_16_XOR2X1_8 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_27_DFFSR_140 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_47_DFFSR_95 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_9_OAI21X1_59 INVX1_4/gnd DFFSR_51/S FILL
XFILL_26_DFFPOSX1_28 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_3_CLKBUF1_8 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_8_OAI21X1_62 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_17_DFFSR_143 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_8_AND2X2_4 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_6_NAND2X1_83 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_7_OAI21X1_65 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_3_DFFSR_92 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_3_NAND2X1_212 INVX1_23/gnd DFFSR_186/S FILL
XFILL_6_OAI21X1_68 BUFX2_37/A DFFSR_81/S FILL
XFILL_2_NOR2X1_22 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_20_DFFSR_85 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_31_DFFSR_45 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_3_INVX1_39 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_5_NAND2X1_86 INVX1_4/gnd DFFSR_51/S FILL
XFILL_0_OAI21X1_260 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_4_NAND2X1_89 BUFX2_37/A DFFSR_8/S FILL
XFILL_1_INVX1_404 BUFX2_19/gnd DFFSR_52/S FILL
XNAND2X1_83 BUFX2_19/Y INVX1_85/A BUFX2_8/gnd OAI21X1_83/C DFFSR_25/S NAND2X1
XFILL_5_OAI21X1_71 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_3_NAND2X1_92 BUFX2_5/gnd DFFSR_23/S FILL
XOAI21X1_68 BUFX2_23/Y INVX1_77/Y OAI21X1_68/C BUFX2_37/A DFFSR_68/D DFFSR_81/S OAI21X1
XFILL_2_NAND3X1_110 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_3_DFFSR_140 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_4_OAI21X1_74 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_2_BUFX2_30 INVX1_4/gnd DFFSR_51/S FILL
XFILL_44_DFFSR_171 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_3_OAI21X1_77 INVX1_89/gnd DFFSR_36/S FILL
XFILL_2_NAND2X1_95 INVX1_89/gnd DFFSR_36/S FILL
XFILL_4_NAND2X1_146 INVX1_23/gnd DFFSR_91/S FILL
XFILL_34_DFFSR_174 BUFX2_43/A DFFSR_97/S FILL
XFILL_1_OAI21X1_194 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_1_DFFSR_5 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_1_NAND2X1_98 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_2_OAI21X1_80 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_24_DFFSR_177 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_28_DFFSR_92 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_50_DFFSR_12 BUFX2_6/gnd DFFSR_14/S FILL
XINVX1_334 DFFSR_113/Q BUFX2_7/gnd INVX1_334/Y DFFSR_81/S INVX1
XFILL_0_INVX1_224 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_0_INVX1_86 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_39_DFFSR_52 INVX1_94/gnd DFFSR_52/S FILL
XFILL_1_OAI21X1_83 INVX1_94/gnd DFFSR_52/S FILL
XFILL_14_DFFSR_180 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_2_OAI21X1_128 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_0_OAI21X1_86 INVX1_4/gnd DFFSR_51/S FILL
XBUFX2_1 BUFX2_2/A DFFSR_5/gnd BUFX2_1/Y DFFSR_2/S BUFX2
XFILL_12_DFFSR_42 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_1_OAI21X1_7 INVX1_8/gnd DFFSR_5/S FILL
XFILL_37_DFFSR_101 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_2_NAND2X1_242 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_0_DFFSR_177 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_25_DFFSR_9 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_27_DFFSR_104 INVX1_4/gnd DFFSR_4/S FILL
XFILL_36_DFFSR_99 BUFX2_35/A DFFSR_97/S FILL
XFILL_17_DFFSR_107 BUFX2_36/A DFFSR_8/S FILL
XFILL_3_INVX1_151 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_47_DFFSR_59 INVX1_4/gnd DFFSR_51/S FILL
XFILL_8_OAI21X1_26 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_0_OAI21X1_224 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_6_DFFPOSX1_14 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_6_NAND2X1_47 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_3_DFFSR_56 INVX1_2/gnd DFFSR_51/S FILL
XFILL_7_OAI21X1_29 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_20_DFFSR_49 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_3_NAND2X1_176 INVX1_94/gnd DFFSR_25/S FILL
XNAND2X1_47 DFFSR_36/S DFFSR_39/Q DFFSR_79/gnd NAND2X1_47/Y DFFSR_45/S NAND2X1
XFILL_5_NAND2X1_50 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_6_OAI21X1_32 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_4_NAND2X1_53 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_1_INVX1_368 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_5_OAI21X1_35 INVX1_8/gnd DFFSR_5/S FILL
XOAI21X1_32 DFFSR_51/S INVX1_36/Y NAND2X1_32/Y DFFSR_3/gnd DFFSR_32/D DFFSR_4/S OAI21X1
XFILL_24_4_0 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_4_OAI21X1_38 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_3_NAND2X1_56 INVX1_4/gnd DFFSR_51/S FILL
XFILL_3_DFFSR_104 INVX1_4/gnd DFFSR_4/S FILL
XFILL_1_OAI21X1_158 BUFX2_43/A DFFSR_97/S FILL
XFILL_44_DFFSR_135 BUFX2_43/A DFFSR_97/S FILL
XFILL_46_DFFSR_5 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_3_OAI21X1_41 INVX1_8/gnd DFFSR_7/S FILL
XFILL_2_NAND2X1_59 INVX1_2/gnd DFFSR_1/S FILL
XFILL_11_AOI22X1_10 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_1_NAND2X1_62 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_2_OAI21X1_44 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_4_NAND2X1_110 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_34_DFFSR_138 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_10_AOI22X1_13 INVX1_23/gnd DFFSR_186/S FILL
XFILL_0_INVX1_188 BUFX2_35/A DFFSR_97/S FILL
XFILL_24_DFFSR_141 INVX1_94/gnd DFFSR_25/S FILL
XFILL_0_INVX1_50 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_39_DFFSR_16 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_1_OAI21X1_47 INVX1_89/gnd DFFSR_2/S FILL
XFILL_17_DFFSR_96 INVX1_2/gnd DFFSR_1/S FILL
XFILL_28_DFFSR_56 INVX1_2/gnd DFFSR_51/S FILL
XFILL_0_NAND2X1_65 DFFSR_3/gnd DFFSR_4/S FILL
XINVX1_298 DFFSR_13/Q DFFSR_3/gnd INVX1_298/Y DFFSR_65/S INVX1
XFILL_4_5_0 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_14_DFFSR_144 INVX1_8/gnd DFFSR_5/S FILL
XFILL_0_OAI21X1_50 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_0_CLKBUF1_9 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_4_INVX1_295 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_1_NAND2X1_272 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_25_DFFPOSX1_22 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_1_INVX1_7 BUFX2_36/A DFFSR_8/S FILL
XFILL_2_NAND2X1_206 BUFX2_43/A DFFSR_97/S FILL
XFILL_0_DFFSR_141 INVX1_94/gnd DFFSR_25/S FILL
XFILL_47_DFFSR_23 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_41_DFFSR_172 BUFX2_37/A DFFSR_8/S FILL
XFILL_36_DFFSR_63 INVX1_94/gnd DFFSR_52/S FILL
XFILL_3_INVX1_115 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_1_NAND3X1_104 INVX1_23/gnd DFFSR_186/S FILL
XFILL_31_DFFSR_175 INVX1_23/gnd DFFSR_91/S FILL
XFILL_21_DFFSR_178 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_6_NAND2X1_11 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_3_DFFSR_20 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_11_DFFSR_181 INVX1_23/gnd DFFSR_186/S FILL
XFILL_5_NAND2X1_14 BUFX2_43/A DFFSR_23/S FILL
XFILL_3_NAND2X1_140 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_0_OAI21X1_188 INVX1_89/gnd DFFSR_2/S FILL
XFILL_20_DFFSR_13 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_7_XOR2X1_17 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_1_INVX1_332 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_4_NAND2X1_17 INVX1_8/gnd DFFSR_7/S FILL
XNAND2X1_11 DFFSR_11/S DFFSR_3/Q BUFX2_16/gnd OAI21X1_11/C DFFSR_65/S NAND2X1
XFILL_3_NAND2X1_20 INVX1_23/gnd DFFSR_186/S FILL
XFILL_2_NOR2X1_1 BUFX2_36/A DFFSR_6/S FILL
XFILL_8_OAI21X1_5 INVX1_8/gnd DFFSR_5/S FILL
XFILL_11_OAI22X1_58 BUFX2_17/gnd DFFSR_7/S FILL
XDFFPOSX1_14 AND2X2_14/B CLKBUF1_12/Y NOR2X1_45/Y BUFX2_6/gnd DFFSR_14/S DFFPOSX1
XFILL_2_NAND2X1_23 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_10_OAI22X1_61 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_32_1_1 INVX1_8/gnd DFFSR_5/S FILL
XFILL_12_DFFSR_3 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_7_DFFSR_175 INVX1_23/gnd DFFSR_91/S FILL
XFILL_9_NAND3X1_79 BUFX2_36/A DFFSR_6/S FILL
XFILL_1_OAI21X1_122 INVX1_94/gnd DFFSR_25/S FILL
XFILL_34_DFFSR_102 INVX1_8/gnd DFFSR_7/S FILL
XFILL_44_DFFSR_70 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_1_NAND2X1_26 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_24_DFFSR_105 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_8_NAND3X1_82 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_9_OAI22X1_64 INVX1_94/gnd DFFSR_25/S FILL
XFILL_0_NAND2X1_29 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_28_DFFSR_20 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_0_INVX1_14 BUFX2_35/A DFFSR_14/S FILL
XFILL_0_INVX1_152 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_17_DFFSR_60 BUFX2_37/A DFFSR_8/S FILL
XFILL_7_NAND3X1_85 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_14_DFFSR_108 INVX1_89/gnd DFFSR_2/S FILL
XFILL_30_3_2 DFFSR_5/gnd DFFSR_2/S FILL
XINVX1_262 INVX1_2/A INVX1_2/gnd OAI22X1_5/C DFFSR_1/S INVX1
XFILL_0_DFFSR_67 INVX1_2/gnd DFFSR_51/S FILL
XFILL_8_OAI22X1_67 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_1_OAI21X1_11 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_0_OAI21X1_14 BUFX2_43/A DFFSR_23/S FILL
XFILL_6_NAND3X1_88 INVX1_94/gnd DFFSR_52/S FILL
XFILL_1_NAND2X1_236 INVX1_2/gnd DFFSR_1/S FILL
XFILL_5_NAND3X1_91 BUFX2_43/A DFFSR_97/S FILL
XNAND3X1_88 INVX1_250/Y NAND3X1_86/Y NAND3X1_87/Y INVX1_94/gnd NAND3X1_88/Y DFFSR_52/S
+ NAND3X1
XFILL_0_NAND3X1_134 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_4_NAND3X1_94 BUFX2_35/A DFFSR_97/S FILL
XFILL_0_DFFSR_105 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_3_NAND3X1_97 BUFX2_35/A DFFSR_97/S FILL
XFILL_2_NAND2X1_170 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_41_DFFSR_136 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_36_DFFSR_27 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_8_DFFSR_74 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_25_DFFSR_67 INVX1_2/gnd DFFSR_51/S FILL
XFILL_31_DFFSR_139 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_7_CLKBUF1_7 BUFX2_43/A DFFSR_97/S FILL
XFILL_0_OAI21X1_152 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_21_DFFSR_142 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_14_DFFPOSX1_27 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_11_DFFSR_145 INVX1_23/gnd DFFSR_186/S FILL
XFILL_9_OAI21X1_207 BUFX2_37/A DFFSR_8/S FILL
XFILL_3_NAND2X1_104 INVX1_4/gnd DFFSR_51/S FILL
XFILL_1_INVX1_296 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_6_NOR2X1_21 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_24_DFFPOSX1_16 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_10_OAI22X1_25 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_44_DFFSR_34 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_33_DFFSR_74 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_7_DFFSR_139 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_0_NAND2X1_266 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_48_DFFSR_170 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_38_DFFSR_173 BUFX2_6/gnd DFFSR_91/S FILL
XINVX1_226 AND2X2_9/A BUFX2_35/A INVX1_226/Y DFFSR_14/S INVX1
XFILL_8_NAND3X1_46 BUFX2_35/A DFFSR_97/S FILL
XFILL_0_DFFSR_31 BUFX2_35/A DFFSR_97/S FILL
XFILL_9_OAI22X1_28 INVX1_94/gnd DFFSR_25/S FILL
XFILL_0_INVX1_116 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_17_DFFSR_24 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_7_NAND3X1_49 BUFX2_37/A DFFSR_8/S FILL
XFILL_8_OAI22X1_31 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_28_DFFSR_176 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_1_NAND2X1_200 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_4_INVX1_223 BUFX2_35/A DFFSR_97/S FILL
XFILL_6_NAND3X1_52 BUFX2_36/A DFFSR_8/S FILL
XFILL_18_DFFSR_179 INVX1_2/gnd DFFSR_1/S FILL
XFILL_7_OAI22X1_34 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_5_NAND3X1_55 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_6_OAI22X1_37 DFFSR_71/gnd DFFSR_45/S FILL
XNAND3X1_52 INVX1_238/A NAND3X1_52/B AOI21X1_27/B BUFX2_36/A NAND3X1_52/Y DFFSR_8/S
+ NAND3X1
XFILL_5_OAI22X1_40 BUFX2_37/A DFFSR_8/S FILL
XFILL_41_DFFSR_81 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_4_NAND3X1_58 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_5_OAI21X1_6 BUFX2_36/A DFFSR_6/S FILL
XFILL_4_OAI22X1_43 BUFX2_8/gnd DFFSR_25/S FILL
XOAI22X1_37 INVX1_330/Y OAI22X1_49/D INVX1_329/Y OAI22X1_52/D DFFSR_71/gnd NOR2X1_28/B
+ DFFSR_45/S OAI22X1
XFILL_3_NAND3X1_61 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_2_NAND2X1_134 DFFSR_79/gnd DFFSR_36/S FILL
XDFFSR_179 NAND2X1_4/B DFFSR_1/CLK DFFSR_183/R DFFSR_1/S DFFSR_179/D INVX1_2/gnd DFFSR_1/S
+ DFFSR
XFILL_41_DFFSR_100 INVX1_23/gnd DFFSR_186/S FILL
XFILL_2_NAND3X1_64 BUFX2_35/A DFFSR_14/S FILL
XFILL_25_DFFSR_31 BUFX2_35/A DFFSR_97/S FILL
XFILL_3_OAI22X1_46 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_8_OAI21X1_237 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_8_DFFSR_38 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_1_NAND3X1_67 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_2_OAI22X1_49 INVX1_94/gnd DFFSR_25/S FILL
XFILL_14_DFFSR_71 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_31_DFFSR_103 INVX1_8/gnd DFFSR_7/S FILL
XFILL_4_DFFSR_176 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_0_NAND3X1_70 BUFX2_35/A DFFSR_14/S FILL
XFILL_1_OAI22X1_52 INVX1_94/gnd DFFSR_25/S FILL
XFILL_21_DFFSR_106 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_11_DFFSR_109 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_9_OAI21X1_171 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_0_OAI22X1_55 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_0_OAI21X1_116 INVX1_89/gnd DFFSR_2/S FILL
XFILL_1_INVX1_260 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_1_XOR2X1_8 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_0_DFFSR_2 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_49_DFFSR_88 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_0_NAND2X1_230 BUFX2_36/A DFFSR_6/S FILL
XINVX1_72 DFFSR_64/Q BUFX2_16/gnd INVX1_72/Y DFFSR_11/S INVX1
XFILL_5_DFFSR_85 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_7_DFFSR_103 INVX1_8/gnd DFFSR_7/S FILL
XFILL_33_DFFSR_38 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_22_DFFSR_78 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_8_NAND3X1_10 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_48_DFFSR_134 DFFSR_79/gnd DFFSR_45/S FILL
XINVX1_190 INVX1_190/A BUFX2_43/A INVX1_190/Y DFFSR_97/S INVX1
XFILL_38_DFFSR_137 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_4_BUFX2_23 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_7_NAND3X1_13 INVX1_94/gnd DFFSR_25/S FILL
XFILL_4_INVX1_187 INVX1_23/gnd DFFSR_186/S FILL
XFILL_6_NAND3X1_16 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_28_DFFSR_140 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_1_NAND2X1_164 INVX1_8/gnd DFFSR_5/S FILL
XFILL_24_DFFSR_6 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_4_CLKBUF1_8 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_18_DFFSR_143 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_14_NOR3X1_2 INVX1_89/gnd DFFSR_2/S FILL
XFILL_5_NAND3X1_19 INVX1_8/gnd DFFSR_5/S FILL
XNAND3X1_16 INVX1_224/A NAND3X1_15/Y NAND3X1_14/Y BUFX2_19/gnd AOI21X1_3/B DFFSR_52/S
+ NAND3X1
XFILL_9_NAND3X1_117 INVX1_94/gnd DFFSR_25/S FILL
XFILL_31_4_0 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_13_DFFPOSX1_21 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_4_NAND3X1_22 BUFX2_37/A DFFSR_81/S FILL
XFILL_3_NOR2X1_22 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_30_DFFSR_85 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_41_DFFSR_45 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_2_INVX1_79 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_8_OAI21X1_201 BUFX2_35/A DFFSR_97/S FILL
XFILL_3_NAND3X1_25 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_2_INVX1_404 BUFX2_19/gnd DFFSR_52/S FILL
XDFFSR_143 DFFSR_143/Q CLKBUF1_9/Y DFFSR_137/R DFFSR_10/S DFFSR_143/D BUFX2_8/gnd
+ DFFSR_25/S DFFSR
XFILL_2_NAND3X1_28 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_4_DFFSR_140 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_14_DFFSR_35 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_3_OAI22X1_10 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_45_DFFSR_171 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_1_NAND3X1_31 INVX1_94/gnd DFFSR_52/S FILL
XFILL_2_OAI22X1_13 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_35_DFFSR_174 BUFX2_43/A DFFSR_97/S FILL
XFILL_0_NAND3X1_34 INVX1_2/gnd DFFSR_1/S FILL
XFILL_1_OAI22X1_16 INVX1_4/gnd DFFSR_4/S FILL
XFILL_9_OAI21X1_135 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_0_OAI22X1_19 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_45_DFFSR_2 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_25_DFFSR_177 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_23_DFFPOSX1_10 INVX1_8/gnd DFFSR_5/S FILL
XFILL_38_DFFSR_92 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_1_INVX1_224 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_49_DFFSR_52 INVX1_94/gnd DFFSR_52/S FILL
XFILL_15_DFFSR_180 BUFX2_17/gnd DFFSR_7/S FILL
XDFFSR_89 DFFSR_89/Q CLKBUF1_7/Y DFFSR_89/R DFFSR_92/S DFFSR_89/D DFFSR_89/gnd DFFSR_92/S
+ DFFSR
XFILL_0_NAND2X1_194 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_11_DFFSR_82 DFFSR_1/gnd DFFSR_9/S FILL
XINVX1_36 INVX1_36/A DFFSR_3/gnd INVX1_36/Y DFFSR_65/S INVX1
XFILL_22_DFFSR_42 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_5_DFFSR_49 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_2_OAI21X1_7 INVX1_8/gnd DFFSR_5/S FILL
XINVX1_154 BUFX2_8/Y INVX1_8/gnd DFFSR_135/R DFFSR_7/S INVX1
XFILL_38_DFFSR_101 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_1_DFFSR_177 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_28_DFFSR_104 INVX1_4/gnd DFFSR_4/S FILL
XFILL_0_INVX1_4 INVX1_4/gnd DFFSR_4/S FILL
XFILL_46_DFFSR_99 BUFX2_35/A DFFSR_97/S FILL
XFILL_7_OAI21X1_231 BUFX2_36/A DFFSR_6/S FILL
XFILL_18_DFFSR_107 BUFX2_36/A DFFSR_8/S FILL
XFILL_1_NAND2X1_128 INVX1_89/gnd DFFSR_2/S FILL
XFILL_19_DFFSR_89 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_7_AND2X2_8 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_2_INVX1_43 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_2_DFFSR_96 INVX1_2/gnd DFFSR_1/S FILL
XFILL_30_DFFSR_49 DFFSR_73/gnd DFFSR_11/S FILL
XDFFSR_107 INVX1_121/A CLKBUF1_6/Y DFFSR_105/R DFFSR_8/S DFFSR_107/D BUFX2_36/A DFFSR_8/S
+ DFFSR
XFILL_39_1_1 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_8_OAI21X1_165 BUFX2_35/A DFFSR_97/S FILL
XFILL_2_INVX1_368 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_1_BUFX2_34 BUFX2_37/A DFFSR_81/S FILL
XFILL_4_DFFSR_104 INVX1_4/gnd DFFSR_4/S FILL
XFILL_37_3_2 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_45_DFFSR_135 BUFX2_43/A DFFSR_97/S FILL
XFILL_35_DFFSR_138 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_1_INVX1_188 BUFX2_35/A DFFSR_97/S FILL
XFILL_25_DFFSR_141 INVX1_94/gnd DFFSR_25/S FILL
XFILL_49_DFFSR_16 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_27_DFFSR_96 INVX1_2/gnd DFFSR_1/S FILL
XFILL_38_DFFSR_56 INVX1_2/gnd DFFSR_51/S FILL
XFILL_15_DFFSR_144 INVX1_8/gnd DFFSR_5/S FILL
XFILL_1_CLKBUF1_9 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_40_2 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_0_NAND2X1_158 BUFX2_35/A DFFSR_97/S FILL
XDFFSR_53 DFFSR_53/Q DFFSR_52/CLK DFFSR_54/R DFFSR_10/S DFFSR_53/D DFFSR_71/gnd DFFSR_10/S
+ DFFSR
XFILL_6_OAI21X1_261 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_11_DFFSR_46 BUFX2_36/A DFFSR_6/S FILL
XFILL_0_NOR2X1_23 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_5_DFFSR_13 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_12_DFFPOSX1_15 BUFX2_35/A DFFSR_14/S FILL
XINVX1_118 BUFX2_9/Y BUFX2_37/A DFFSR_97/R DFFSR_8/S INVX1
XFILL_1_DFFSR_141 INVX1_94/gnd DFFSR_25/S FILL
XFILL_8_NAND3X1_111 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_42_DFFSR_172 BUFX2_37/A DFFSR_8/S FILL
XFILL_7_OAI21X1_195 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_46_DFFSR_63 INVX1_94/gnd DFFSR_52/S FILL
XFILL_32_DFFSR_175 INVX1_23/gnd DFFSR_91/S FILL
XFILL_22_DFFSR_178 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_12_DFFSR_181 INVX1_23/gnd DFFSR_186/S FILL
XFILL_2_DFFSR_60 BUFX2_37/A DFFSR_8/S FILL
XFILL_19_DFFSR_53 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_30_DFFSR_13 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_8_XOR2X1_17 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_2_INVX1_332 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_8_OAI21X1_129 INVX1_4/gnd DFFSR_4/S FILL
XFILL_8_DFFSR_175 INVX1_23/gnd DFFSR_91/S FILL
XFILL_2_DFFPOSX1_26 BUFX2_37/A DFFSR_81/S FILL
XFILL_35_DFFSR_102 INVX1_8/gnd DFFSR_7/S FILL
XFILL_36_DFFSR_9 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_25_DFFSR_105 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_38_DFFSR_20 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_1_INVX1_152 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_27_DFFSR_60 BUFX2_37/A DFFSR_8/S FILL
XFILL_15_DFFSR_108 INVX1_89/gnd DFFSR_2/S FILL
XFILL_6_OAI21X1_225 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_0_NAND2X1_122 INVX1_94/gnd DFFSR_25/S FILL
XFILL_11_DFFSR_10 DFFSR_71/gnd DFFSR_10/S FILL
XDFFSR_17 DFFSR_17/Q DFFSR_2/CLK DFFSR_20/R DFFSR_17/S DFFSR_17/D DFFSR_5/gnd DFFSR_5/S
+ DFFSR
XFILL_1_DFFSR_105 DFFSR_89/gnd DFFSR_186/S FILL
XOAI21X1_261 NOR3X1_2/C AND2X2_17/Y AND2X2_16/B DFFSR_79/gnd XOR2X1_15/A DFFSR_36/S
+ OAI21X1
XFILL_7_OAI21X1_159 BUFX2_43/A DFFSR_97/S FILL
XFILL_11_1_2 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_42_DFFSR_136 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_46_DFFSR_27 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_35_DFFSR_67 INVX1_2/gnd DFFSR_51/S FILL
XFILL_32_DFFSR_139 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_8_CLKBUF1_7 BUFX2_43/A DFFSR_97/S FILL
XFILL_22_DFFSR_142 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_19_DFFSR_17 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_2_DFFSR_24 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_12_DFFSR_145 INVX1_23/gnd DFFSR_186/S FILL
XFILL_2_INVX1_296 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_1_NOR2X1_5 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_45_7 INVX1_2/gnd DFFSR_51/S FILL
XFILL_19_CLKBUF1_10 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_43_DFFSR_74 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_8_DFFSR_139 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_49_DFFSR_170 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_18_CLKBUF1_13 INVX1_4/gnd DFFSR_51/S FILL
XFILL_5_OAI21X1_255 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_39_DFFSR_173 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_17_CLKBUF1_16 BUFX2_36/A DFFSR_6/S FILL
XFILL_1_INVX1_116 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_27_DFFSR_24 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_7_NAND3X1_105 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_16_CLKBUF1_19 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_29_DFFSR_176 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_16_DFFSR_64 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_38_4_0 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_15_CLKBUF1_22 INVX1_94/gnd DFFSR_25/S FILL
XFILL_6_OAI21X1_189 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_19_DFFSR_179 INVX1_2/gnd DFFSR_1/S FILL
XFILL_14_CLKBUF1_25 INVX1_23/gnd DFFSR_186/S FILL
XFILL_51_DFFSR_81 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_3_XOR2X1_1 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_23_DFFSR_3 DFFSR_3/gnd DFFSR_4/S FILL
XOAI21X1_225 AOI22X1_10/Y AOI22X1_11/Y AOI21X1_25/Y BUFX2_6/gnd NAND3X1_71/B DFFSR_91/S
+ OAI21X1
XFILL_6_OAI21X1_6 BUFX2_36/A DFFSR_6/S FILL
XFILL_42_DFFSR_100 INVX1_23/gnd DFFSR_186/S FILL
XFILL_7_OAI21X1_123 INVX1_23/gnd DFFSR_91/S FILL
XFILL_7_DFFSR_78 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_35_DFFSR_31 BUFX2_35/A DFFSR_97/S FILL
XFILL_24_DFFSR_71 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_32_DFFSR_103 INVX1_8/gnd DFFSR_7/S FILL
XFILL_5_DFFSR_176 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_22_DFFSR_106 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_12_DFFSR_109 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_1_DFFPOSX1_20 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_6_BUFX2_16 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_2_INVX1_260 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_5_OAI21X1_219 BUFX2_35/A DFFSR_97/S FILL
XFILL_8_DFFSR_103 INVX1_8/gnd DFFSR_7/S FILL
XFILL_43_DFFSR_38 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_32_DFFSR_78 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_49_DFFSR_134 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_39_DFFSR_137 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_16_DFFSR_28 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_29_DFFSR_140 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_46_1_1 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_6_OAI21X1_153 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_5_CLKBUF1_8 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_19_DFFSR_143 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_20_DFFPOSX1_28 DFFSR_3/gnd DFFSR_65/S FILL
XNOR2X1_25 NOR2X1_25/A NOR2X1_25/B DFFSR_71/gnd NOR2X1_25/Y DFFSR_45/S NOR2X1
XFILL_44_3_2 INVX1_2/gnd DFFSR_51/S FILL
XFILL_4_NOR2X1_22 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_40_DFFSR_85 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_51_DFFSR_45 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_3_INVX1_404 BUFX2_19/gnd DFFSR_52/S FILL
XOAI21X1_189 BUFX2_1/Y XOR2X1_3/Y NAND3X1_19/Y DFFSR_73/gnd DFFPOSX1_5/D DFFSR_57/S
+ OAI21X1
XFILL_6_NAND2X1_267 INVX1_4/gnd DFFSR_4/S FILL
XFILL_5_DFFSR_140 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_24_DFFSR_35 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_13_DFFSR_75 INVX1_4/gnd DFFSR_51/S FILL
XFILL_7_DFFSR_42 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_46_DFFSR_171 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_36_DFFSR_174 BUFX2_43/A DFFSR_97/S FILL
XFILL_4_OAI21X1_249 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_12_2_0 BUFX2_36/A DFFSR_6/S FILL
XFILL_26_DFFSR_177 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_48_DFFSR_92 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_2_INVX1_224 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_16_DFFSR_180 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_4_DFFSR_89 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_10_4_1 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_9_AND2X2_1 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_7_CLKBUF1_10 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_21_DFFSR_82 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_4_INVX1_36 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_32_DFFSR_42 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_3_OAI21X1_7 INVX1_8/gnd DFFSR_5/S FILL
XFILL_5_OAI21X1_183 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_6_CLKBUF1_13 INVX1_4/gnd DFFSR_51/S FILL
XFILL_5_CLKBUF1_16 BUFX2_36/A DFFSR_6/S FILL
XCLKBUF1_13 clk INVX1_4/gnd CLKBUF1_13/Y DFFSR_51/S CLKBUF1
XFILL_39_DFFSR_101 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_3_BUFX2_27 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_5_3 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_2_DFFSR_177 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_4_CLKBUF1_19 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_29_DFFSR_104 INVX1_4/gnd DFFSR_4/S FILL
XFILL_6_OAI21X1_117 BUFX2_35/A DFFSR_97/S FILL
XFILL_19_DFFSR_107 BUFX2_36/A DFFSR_8/S FILL
XFILL_3_CLKBUF1_22 INVX1_94/gnd DFFSR_25/S FILL
XFILL_2_CLKBUF1_25 INVX1_23/gnd DFFSR_186/S FILL
XFILL_29_DFFSR_89 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_1_INVX1_83 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_40_DFFSR_49 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_0_DFFPOSX1_14 BUFX2_6/gnd DFFSR_14/S FILL
XOAI21X1_153 DFFSR_23/S INVX1_180/Y NAND2X1_153/Y BUFX2_5/gnd DFFSR_153/D DFFSR_6/S
+ OAI21X1
XFILL_6_NAND2X1_231 BUFX2_37/A DFFSR_81/S FILL
XFILL_3_INVX1_368 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_13_DFFSR_39 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_5_DFFSR_104 INVX1_4/gnd DFFSR_4/S FILL
XFILL_5_NAND3X1_129 BUFX2_35/A DFFSR_14/S FILL
XFILL_46_DFFSR_135 BUFX2_43/A DFFSR_97/S FILL
XFILL_4_OAI21X1_213 BUFX2_36/A DFFSR_6/S FILL
XNAND2X1_267 DFFSR_51/S DFFSR_164/Q INVX1_4/gnd NAND2X1_267/Y DFFSR_4/S NAND2X1
XFILL_36_DFFSR_138 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_2_INVX1_188 BUFX2_35/A DFFSR_97/S FILL
XFILL_35_DFFSR_6 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_26_DFFSR_141 INVX1_94/gnd DFFSR_25/S FILL
XFILL_37_DFFSR_96 INVX1_2/gnd DFFSR_1/S FILL
XFILL_48_DFFSR_56 INVX1_2/gnd DFFSR_51/S FILL
XFILL_16_DFFSR_144 INVX1_8/gnd DFFSR_5/S FILL
XFILL_2_CLKBUF1_9 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_5_OAI21X1_147 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_21_DFFSR_46 BUFX2_36/A DFFSR_6/S FILL
XFILL_18_1_2 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_4_DFFSR_53 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_1_NOR2X1_23 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_10_DFFSR_86 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_19_DFFPOSX1_22 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_0_0_1 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_0_INVX1_405 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_2_DFFSR_141 INVX1_94/gnd DFFSR_25/S FILL
XFILL_43_DFFSR_172 BUFX2_37/A DFFSR_8/S FILL
XFILL_33_DFFSR_175 INVX1_23/gnd DFFSR_91/S FILL
XFILL_5_NAND2X1_261 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_23_DFFSR_178 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_13_DFFSR_181 INVX1_23/gnd DFFSR_186/S FILL
XFILL_29_DFFSR_53 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_1_INVX1_47 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_18_DFFSR_93 INVX1_2/gnd DFFSR_51/S FILL
XFILL_40_DFFSR_13 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_3_OAI21X1_243 BUFX2_6/gnd DFFSR_14/S FILL
XOAI21X1_117 BUFX2_21/Y INVX1_132/Y NAND2X1_117/Y BUFX2_35/A DFFSR_117/D DFFSR_97/S
+ OAI21X1
XFILL_6_NAND2X1_195 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_9_XOR2X1_17 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_3_INVX1_332 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_0_OAI21X1_8 BUFX2_36/A DFFSR_6/S FILL
XFILL_0_BUFX2_38 BUFX2_37/A DFFSR_81/S FILL
XFILL_45_4_0 INVX1_2/gnd DFFSR_1/S FILL
XFILL_9_DFFSR_175 INVX1_23/gnd DFFSR_91/S FILL
XNAND2X1_231 NAND3X1_109/Y NAND2X1_231/B BUFX2_37/A NAND2X1_231/Y DFFSR_81/S NAND2X1
XFILL_36_DFFSR_102 INVX1_8/gnd DFFSR_7/S FILL
XFILL_26_DFFSR_105 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_4_OAI21X1_177 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_48_DFFSR_20 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_2_INVX1_152 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_37_DFFSR_60 BUFX2_37/A DFFSR_8/S FILL
XFILL_16_DFFSR_108 INVX1_89/gnd DFFSR_2/S FILL
XFILL_21_DFFSR_10 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_4_DFFSR_17 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_10_DFFSR_50 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_5_OAI21X1_111 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_0_INVX1_369 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_2_DFFSR_105 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_2_DFFSR_9 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_5_NAND2X1_225 BUFX2_36/A DFFSR_8/S FILL
XFILL_43_DFFSR_136 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_45_DFFSR_67 INVX1_2/gnd DFFSR_51/S FILL
XFILL_33_DFFSR_139 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_9_CLKBUF1_7 BUFX2_43/A DFFSR_97/S FILL
XFILL_23_DFFSR_142 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_4_NAND3X1_123 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_29_DFFSR_17 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_18_DFFSR_57 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_1_INVX1_11 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_1_DFFSR_64 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_13_DFFSR_145 INVX1_23/gnd DFFSR_186/S FILL
XFILL_3_OAI21X1_207 BUFX2_37/A DFFSR_8/S FILL
XFILL_6_BUFX2_1 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_6_NAND2X1_159 BUFX2_43/A DFFSR_97/S FILL
XFILL_3_INVX1_296 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_9_DFFSR_139 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_18_DFFPOSX1_16 BUFX2_6/gnd DFFSR_91/S FILL
XNAND2X1_195 NAND3X1_21/C NAND2X1_195/B BUFX2_7/gnd AOI22X1_5/C DFFSR_81/S NAND2X1
XFILL_50_DFFSR_170 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_4_OAI21X1_141 INVX1_94/gnd DFFSR_52/S FILL
XFILL_40_DFFSR_173 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_9_DFFSR_71 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_2_INVX1_116 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_37_DFFSR_24 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_18_DFFPOSX1_1 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_30_DFFSR_176 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_26_DFFSR_64 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_17_DFFPOSX1_4 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_20_DFFSR_179 INVX1_2/gnd DFFSR_1/S FILL
XFILL_10_DFFSR_14 BUFX2_35/A DFFSR_14/S FILL
XFILL_16_DFFPOSX1_7 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_10_DFFSR_182 INVX1_89/gnd DFFSR_36/S FILL
XFILL_4_NAND2X1_255 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_0_INVX1_333 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_7_OAI21X1_6 BUFX2_36/A DFFSR_6/S FILL
XFILL_47_DFFSR_9 DFFSR_9/gnd DFFSR_9/S FILL
XFILL_43_DFFSR_100 INVX1_23/gnd DFFSR_186/S FILL
XFILL_2_OAI21X1_237 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_8_DFFPOSX1_27 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_45_DFFSR_31 BUFX2_35/A DFFSR_97/S FILL
XFILL_5_NAND2X1_189 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_19_2_0 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_34_DFFSR_71 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_33_DFFSR_103 INVX1_8/gnd DFFSR_7/S FILL
XFILL_6_DFFSR_176 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_23_DFFSR_106 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_13_DFFSR_109 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_17_4_1 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_1_DFFSR_28 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_18_DFFSR_21 INVX1_2/gnd DFFSR_1/S FILL
XFILL_3_INVX1_260 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_6_NAND2X1_123 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_10_OAI22X1_2 BUFX2_36/A DFFSR_8/S FILL
XFILL_3_OAI21X1_171 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_0_NOR2X1_9 BUFX2_43/A DFFSR_97/S FILL
XFILL_9_NOR3X1_2 INVX1_89/gnd DFFSR_2/S FILL
XNAND2X1_159 INVX1_190/A DFFSR_23/S BUFX2_43/A NAND2X1_159/Y DFFSR_97/S NAND2X1
XFILL_3_NAND2X1_285 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_9_AOI21X1_48 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_9_DFFSR_103 INVX1_8/gnd DFFSR_7/S FILL
XFILL_42_DFFSR_78 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_4_OAI21X1_105 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_50_DFFSR_134 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_15_DFFSR_68 BUFX2_35/A DFFSR_14/S FILL
XFILL_40_DFFSR_137 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_26_DFFSR_28 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_9_DFFSR_35 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_30_DFFSR_140 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_6_CLKBUF1_8 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_4_NAND2X1_219 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_20_DFFSR_143 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_10_DFFSR_146 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_2_XOR2X1_5 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_3_NAND3X1_117 INVX1_94/gnd DFFSR_25/S FILL
XFILL_5_NOR2X1_22 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_50_DFFSR_85 DFFSR_71/gnd DFFSR_45/S FILL
XINVX1_407 INVX1_407/A DFFSR_5/gnd INVX1_407/Y DFFSR_2/S INVX1
XFILL_13_DFFSR_7 INVX1_8/gnd DFFSR_7/S FILL
XFILL_0_INVX1_297 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_2_OAI21X1_201 BUFX2_35/A DFFSR_97/S FILL
XFILL_5_NAND2X1_153 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_4_INVX1_404 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_6_DFFSR_140 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_34_DFFSR_35 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_6_DFFSR_82 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_23_DFFSR_75 INVX1_4/gnd DFFSR_51/S FILL
XFILL_47_DFFSR_171 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_37_DFFSR_174 BUFX2_43/A DFFSR_97/S FILL
XFILL_3_OAI21X1_135 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_5_BUFX2_20 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_25_1_2 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_27_DFFSR_177 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_17_DFFPOSX1_10 INVX1_8/gnd DFFSR_5/S FILL
XFILL_3_INVX1_224 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_17_DFFSR_180 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_7_0_1 BUFX2_35/A DFFSR_97/S FILL
XFILL_8_OAI21X1_99 BUFX2_43/A DFFSR_97/S FILL
XFILL_34_DFFSR_3 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_9_AOI21X1_12 INVX1_8/gnd DFFSR_7/S FILL
XFILL_31_DFFSR_82 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_3_INVX1_76 INVX1_2/gnd DFFSR_1/S FILL
XFILL_42_DFFSR_42 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_5_2_2 BUFX2_6/gnd DFFSR_14/S FILL
XNAND2X1_123 BUFX2_25/Y DFFSR_115/Q BUFX2_6/gnd OAI21X1_123/C DFFSR_14/S NAND2X1
XFILL_8_AOI21X1_15 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_4_OAI21X1_7 INVX1_8/gnd DFFSR_5/S FILL
XFILL_3_NAND2X1_249 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_6_DFFPOSX1_1 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_7_AOI21X1_18 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_40_DFFSR_101 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_3_DFFSR_177 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_5_DFFPOSX1_4 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_15_DFFSR_32 INVX1_2/gnd DFFSR_1/S FILL
XFILL_30_DFFSR_104 INVX1_4/gnd DFFSR_4/S FILL
XDFFPOSX1_1 DFFPOSX1_1/Q CLKBUF1_12/Y AND2X2_1/Y BUFX2_6/gnd DFFSR_14/S DFFPOSX1
XFILL_6_AOI21X1_21 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_7_DFFPOSX1_21 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_1_OAI21X1_231 BUFX2_36/A DFFSR_6/S FILL
XFILL_20_DFFSR_107 BUFX2_36/A DFFSR_8/S FILL
XFILL_5_AOI21X1_24 BUFX2_43/A DFFSR_97/S FILL
XAOI21X1_21 NAND3X1_42/Y NAND3X1_48/B AOI22X1_5/Y BUFX2_5/gnd AOI21X1_25/C DFFSR_23/S
+ AOI21X1
XFILL_4_DFFPOSX1_7 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_4_NAND2X1_183 INVX1_8/gnd DFFSR_7/S FILL
XFILL_10_DFFSR_110 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_39_DFFSR_89 DFFSR_89/gnd DFFSR_92/S FILL
XINVX1_371 DFFSR_109/Q BUFX2_5/gnd INVX1_371/Y DFFSR_23/S INVX1
XFILL_4_AOI21X1_27 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_0_INVX1_261 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_50_DFFSR_49 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_3_AOI21X1_30 INVX1_23/gnd DFFSR_91/S FILL
XFILL_2_AOI21X1_33 BUFX2_35/A DFFSR_14/S FILL
XFILL_2_OAI21X1_165 BUFX2_35/A DFFSR_97/S FILL
XFILL_4_INVX1_368 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_5_NAND2X1_117 BUFX2_35/A DFFSR_14/S FILL
XFILL_6_DFFSR_46 BUFX2_36/A DFFSR_6/S FILL
XFILL_1_AOI21X1_36 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_23_DFFSR_39 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_12_DFFSR_79 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_6_DFFSR_104 INVX1_4/gnd DFFSR_4/S FILL
XFILL_47_DFFSR_135 BUFX2_43/A DFFSR_97/S FILL
XFILL_0_AOI21X1_39 BUFX2_7/gnd DFFSR_81/S FILL
XBUFX2_24 INVX1_1/Y DFFSR_73/gnd BUFX2_24/Y DFFSR_11/S BUFX2
XFILL_37_DFFSR_138 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_3_INVX1_188 BUFX2_35/A DFFSR_97/S FILL
XFILL_14_6 BUFX2_36/A DFFSR_8/S FILL
XFILL_9_OAI21X1_60 BUFX2_37/A DFFSR_81/S FILL
XFILL_16_XOR2X1_9 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_27_DFFSR_141 INVX1_94/gnd DFFSR_25/S FILL
XFILL_2_NAND2X1_279 INVX1_89/gnd DFFSR_2/S FILL
XFILL_31_1 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_26_DFFPOSX1_29 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_8_OAI21X1_63 INVX1_94/gnd DFFSR_25/S FILL
XFILL_17_DFFSR_144 INVX1_8/gnd DFFSR_5/S FILL
XFILL_3_CLKBUF1_9 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_47_DFFSR_96 INVX1_2/gnd DFFSR_1/S FILL
XFILL_6_NAND2X1_84 BUFX2_36/A DFFSR_6/S FILL
XFILL_8_AND2X2_5 BUFX2_37/A DFFSR_81/S FILL
XFILL_7_OAI21X1_66 INVX1_4/gnd DFFSR_51/S FILL
XFILL_3_NAND2X1_213 BUFX2_35/A DFFSR_97/S FILL
XFILL_31_DFFSR_46 BUFX2_36/A DFFSR_6/S FILL
XFILL_6_OAI21X1_69 BUFX2_37/A DFFSR_8/S FILL
XFILL_2_NOR2X1_23 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_0_OAI21X1_261 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_5_NAND2X1_87 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_3_INVX1_40 INVX1_8/gnd DFFSR_5/S FILL
XFILL_20_DFFSR_86 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_3_DFFSR_93 INVX1_2/gnd DFFSR_51/S FILL
XNAND2X1_84 BUFX2_20/Y DFFSR_76/Q BUFX2_36/A OAI21X1_84/C DFFSR_6/S NAND2X1
XFILL_5_OAI21X1_72 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_4_NAND2X1_90 DFFSR_1/gnd DFFSR_1/S FILL
XOAI21X1_69 BUFX2_23/Y INVX1_78/Y OAI21X1_69/C BUFX2_37/A DFFSR_69/D DFFSR_8/S OAI21X1
XFILL_1_INVX1_405 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_3_DFFSR_141 INVX1_94/gnd DFFSR_25/S FILL
XFILL_2_NAND3X1_111 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_4_OAI21X1_75 INVX1_4/gnd DFFSR_4/S FILL
XFILL_3_NAND2X1_93 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_44_DFFSR_172 BUFX2_37/A DFFSR_8/S FILL
XFILL_2_BUFX2_31 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_4_NAND2X1_147 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_34_DFFSR_175 INVX1_23/gnd DFFSR_91/S FILL
XFILL_1_DFFSR_6 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_1_OAI21X1_195 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_3_OAI21X1_78 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_2_NAND2X1_96 INVX1_4/gnd DFFSR_51/S FILL
XFILL_1_NAND2X1_99 BUFX2_43/A DFFSR_97/S FILL
XFILL_2_OAI21X1_81 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_24_DFFSR_178 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_14_DFFSR_181 INVX1_23/gnd DFFSR_186/S FILL
XFILL_1_OAI21X1_84 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_0_INVX1_225 BUFX2_19/gnd DFFSR_54/S FILL
XINVX1_335 DFFSR_81/Q BUFX2_19/gnd INVX1_335/Y DFFSR_54/S INVX1
XFILL_39_DFFSR_53 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_0_INVX1_87 INVX1_89/gnd DFFSR_36/S FILL
XFILL_28_DFFSR_93 INVX1_2/gnd DFFSR_51/S FILL
XFILL_50_DFFSR_13 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_4_INVX1_332 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_0_OAI21X1_87 INVX1_4/gnd DFFSR_4/S FILL
XBUFX2_2 BUFX2_2/A BUFX2_43/A BUFX2_2/Y DFFSR_23/S BUFX2
XFILL_12_DFFSR_43 INVX1_94/gnd DFFSR_25/S FILL
XFILL_6_DFFSR_10 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_2_OAI21X1_129 INVX1_4/gnd DFFSR_4/S FILL
XFILL_1_OAI21X1_8 BUFX2_36/A DFFSR_6/S FILL
XFILL_37_DFFSR_102 INVX1_8/gnd DFFSR_7/S FILL
XFILL_27_DFFSR_105 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_0_DFFSR_178 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_2_NAND2X1_243 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_3_INVX1_152 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_47_DFFSR_60 BUFX2_37/A DFFSR_8/S FILL
XFILL_17_DFFSR_108 INVX1_89/gnd DFFSR_2/S FILL
XFILL_8_OAI21X1_27 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_0_OAI21X1_225 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_31_DFFSR_10 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_7_OAI21X1_30 INVX1_89/gnd DFFSR_36/S FILL
XFILL_3_DFFSR_57 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_6_NAND2X1_48 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_20_DFFSR_50 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_6_DFFPOSX1_15 BUFX2_35/A DFFSR_14/S FILL
XFILL_6_OAI21X1_33 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_26_2_0 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_3_NAND2X1_177 INVX1_89/gnd DFFSR_36/S FILL
XFILL_5_NAND2X1_51 INVX1_2/gnd DFFSR_51/S FILL
XNAND2X1_48 DFFSR_11/S DFFSR_40/Q BUFX2_16/gnd NAND2X1_48/Y DFFSR_11/S NAND2X1
XFILL_4_NAND2X1_54 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_5_OAI21X1_36 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_1_INVX1_369 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_3_DFFSR_105 DFFSR_89/gnd DFFSR_186/S FILL
XOAI21X1_33 DFFSR_52/S INVX1_38/Y OAI21X1_33/C BUFX2_19/gnd DFFSR_33/D DFFSR_52/S
+ OAI21X1
XFILL_24_4_1 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_4_OAI21X1_39 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_3_NAND2X1_57 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_1_OAI21X1_159 BUFX2_43/A DFFSR_97/S FILL
XFILL_46_DFFSR_6 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_2_NAND2X1_60 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_44_DFFSR_136 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_3_OAI21X1_42 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_6_3_0 BUFX2_35/A DFFSR_14/S FILL
XFILL_1_NAND2X1_63 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_2_OAI21X1_45 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_4_NAND2X1_111 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_34_DFFSR_139 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_0_INVX1_189 BUFX2_35/A DFFSR_14/S FILL
XFILL_24_DFFSR_142 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_0_INVX1_51 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_10_AOI22X1_14 DFFSR_79/gnd DFFSR_36/S FILL
XINVX1_299 DFFSR_53/Q INVX1_89/gnd INVX1_299/Y DFFSR_36/S INVX1
XFILL_39_DFFSR_17 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_28_DFFSR_57 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_0_NAND2X1_66 INVX1_4/gnd DFFSR_51/S FILL
XFILL_1_OAI21X1_48 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_14_DFFSR_145 INVX1_23/gnd DFFSR_186/S FILL
XFILL_4_5_1 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_17_DFFSR_97 BUFX2_35/A DFFSR_97/S FILL
XFILL_0_OAI21X1_51 INVX1_2/gnd DFFSR_51/S FILL
XFILL_25_DFFPOSX1_23 INVX1_23/gnd DFFSR_91/S FILL
XFILL_4_INVX1_296 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_1_NAND2X1_273 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_1_INVX1_8 INVX1_8/gnd DFFSR_5/S FILL
XFILL_0_DFFSR_142 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_41_DFFSR_173 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_2_NAND2X1_207 BUFX2_43/A DFFSR_97/S FILL
XFILL_3_INVX1_116 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_1_NAND3X1_105 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_47_DFFSR_24 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_31_DFFSR_176 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_36_DFFSR_64 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_6_NAND2X1_12 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_21_DFFSR_179 INVX1_2/gnd DFFSR_1/S FILL
XFILL_20_DFFSR_14 BUFX2_35/A DFFSR_14/S FILL
XFILL_3_NAND2X1_141 INVX1_94/gnd DFFSR_25/S FILL
XFILL_11_DFFSR_182 INVX1_89/gnd DFFSR_36/S FILL
XFILL_5_NAND2X1_15 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_0_OAI21X1_189 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_3_DFFSR_21 INVX1_2/gnd DFFSR_1/S FILL
XNAND2X1_12 DFFSR_10/S DFFSR_4/Q BUFX2_8/gnd OAI21X1_12/C DFFSR_10/S NAND2X1
XFILL_4_NAND2X1_18 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_9_OAI21X1_244 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_8_OAI21X1_6 BUFX2_36/A DFFSR_6/S FILL
XFILL_2_NOR2X1_2 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_1_INVX1_333 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_11_OAI22X1_59 INVX1_8/gnd DFFSR_7/S FILL
XFILL_3_NAND2X1_21 INVX1_4/gnd DFFSR_4/S FILL
XFILL_44_DFFSR_100 INVX1_23/gnd DFFSR_186/S FILL
XDFFPOSX1_15 INVX1_401/A CLKBUF1_14/Y AOI21X1_41/Y BUFX2_35/A DFFSR_14/S DFFPOSX1
XFILL_10_OAI22X1_62 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_32_1_2 INVX1_8/gnd DFFSR_5/S FILL
XFILL_2_NAND2X1_24 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_12_DFFSR_4 INVX1_4/gnd DFFSR_4/S FILL
XFILL_1_OAI21X1_123 INVX1_23/gnd DFFSR_91/S FILL
XFILL_44_DFFSR_71 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_34_DFFSR_103 INVX1_8/gnd DFFSR_7/S FILL
XFILL_7_DFFSR_176 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_8_NAND3X1_83 BUFX2_37/A DFFSR_81/S FILL
XFILL_1_NAND2X1_27 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_24_DFFSR_106 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_9_OAI22X1_65 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_14_DFFSR_109 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_1_OAI21X1_12 BUFX2_35/A DFFSR_14/S FILL
XFILL_0_DFFSR_68 BUFX2_35/A DFFSR_14/S FILL
XFILL_17_DFFSR_61 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_7_NAND3X1_86 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_0_NAND2X1_30 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_0_INVX1_153 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_28_DFFSR_21 INVX1_2/gnd DFFSR_1/S FILL
XFILL_0_INVX1_15 DFFSR_3/gnd DFFSR_65/S FILL
XINVX1_263 DFFSR_9/Q BUFX2_16/gnd OAI22X1_5/A DFFSR_65/S INVX1
XFILL_11_OAI22X1_2 BUFX2_36/A DFFSR_8/S FILL
XFILL_1_NAND2X1_237 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_8_OAI22X1_68 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_0_OAI21X1_15 BUFX2_17/gnd DFFSR_57/S FILL
XFILL_6_NAND3X1_89 BUFX2_43/A DFFSR_23/S FILL
XNAND3X1_89 NAND3X1_92/A INVX1_258/Y NAND3X1_92/C BUFX2_43/A NAND3X1_97/B DFFSR_23/S
+ NAND3X1
XFILL_5_NAND3X1_92 BUFX2_43/A DFFSR_23/S FILL
XFILL_4_NAND3X1_95 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_3_NAND3X1_98 BUFX2_35/A DFFSR_14/S FILL
XFILL_2_NAND2X1_171 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_0_DFFSR_106 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_25_DFFSR_68 BUFX2_35/A DFFSR_14/S FILL
XFILL_41_DFFSR_137 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_36_DFFSR_28 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_8_DFFSR_75 INVX1_4/gnd DFFSR_51/S FILL
XFILL_31_DFFSR_140 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_0_OAI21X1_153 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_7_CLKBUF1_8 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_21_DFFSR_143 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_14_DFFPOSX1_28 DFFSR_3/gnd DFFSR_65/S FILL
XFILL_11_DFFSR_146 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_3_NAND2X1_105 BUFX2_35/A DFFSR_14/S FILL
XFILL_6_NOR2X1_22 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_1_INVX1_297 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_10_OAI22X1_26 INVX1_94/gnd DFFSR_52/S FILL
XFILL_7_DFFSR_140 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_44_DFFSR_35 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_33_DFFSR_75 INVX1_4/gnd DFFSR_51/S FILL
XFILL_0_NAND2X1_267 INVX1_4/gnd DFFSR_4/S FILL
XFILL_9_NAND3X1_44 BUFX2_5/gnd DFFSR_23/S FILL
XFILL_24_DFFPOSX1_17 BUFX2_37/A DFFSR_8/S FILL
XFILL_48_DFFSR_171 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_8_NAND3X1_47 BUFX2_43/A DFFSR_97/S FILL
XFILL_38_DFFSR_174 BUFX2_43/A DFFSR_97/S FILL
XINVX1_227 AND2X2_5/B BUFX2_5/gnd INVX1_227/Y DFFSR_6/S INVX1
XFILL_9_OAI22X1_29 INVX1_8/gnd DFFSR_5/S FILL
XFILL_0_DFFSR_32 INVX1_2/gnd DFFSR_1/S FILL
XFILL_0_INVX1_117 INVX1_4/gnd DFFSR_51/S FILL
XFILL_7_NAND3X1_50 BUFX2_37/A DFFSR_81/S FILL
XFILL_17_DFFSR_25 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_8_OAI22X1_32 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_28_DFFSR_177 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_1_NAND2X1_201 BUFX2_35/A DFFSR_14/S FILL
XFILL_6_NAND3X1_53 BUFX2_37/A DFFSR_81/S FILL
XFILL_4_INVX1_224 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_18_DFFSR_180 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_7_OAI22X1_35 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_5_NAND3X1_56 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_6_OAI22X1_38 BUFX2_19/gnd DFFSR_52/S FILL
XNAND3X1_53 INVX1_238/Y NAND3X1_53/B NAND3X1_53/C BUFX2_37/A NAND3X1_53/Y DFFSR_81/S
+ NAND3X1
XFILL_4_NAND3X1_59 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_41_DFFSR_82 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_5_OAI22X1_41 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_3_NAND3X1_62 BUFX2_43/A DFFSR_23/S FILL
XOAI22X1_38 INVX1_334/Y OAI22X1_38/B INVX1_335/Y OAI22X1_38/D BUFX2_19/gnd NOR2X1_28/A
+ DFFSR_52/S OAI22X1
XFILL_5_OAI21X1_7 INVX1_8/gnd DFFSR_5/S FILL
XDFFSR_180 NAND2X1_5/B DFFSR_3/CLK DFFSR_183/R DFFSR_7/S DFFSR_180/D BUFX2_17/gnd
+ DFFSR_7/S DFFSR
XFILL_4_OAI22X1_44 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_2_NAND3X1_65 BUFX2_35/A DFFSR_14/S FILL
XFILL_2_NAND2X1_135 BUFX2_36/A DFFSR_6/S FILL
XFILL_3_OAI22X1_47 BUFX2_37/A DFFSR_8/S FILL
XFILL_8_OAI21X1_238 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_41_DFFSR_101 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_1_NAND3X1_68 BUFX2_35/A DFFSR_14/S FILL
XFILL_8_DFFSR_39 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_2_OAI22X1_50 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_4_DFFSR_177 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_14_DFFSR_72 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_25_DFFSR_32 INVX1_2/gnd DFFSR_1/S FILL
XFILL_31_DFFSR_104 INVX1_4/gnd DFFSR_4/S FILL
XFILL_0_NAND3X1_71 BUFX2_35/A DFFSR_14/S FILL
XFILL_21_DFFSR_107 BUFX2_36/A DFFSR_8/S FILL
XFILL_1_OAI22X1_53 DFFSR_71/gnd DFFSR_10/S FILL
XNAND2X1_1 DFFSR_176/Q DFFSR_166/S INVX1_2/gnd OAI21X1_1/C DFFSR_51/S NAND2X1
XFILL_0_OAI21X1_117 BUFX2_35/A DFFSR_97/S FILL
XFILL_11_DFFSR_110 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_49_DFFSR_89 DFFSR_89/gnd DFFSR_92/S FILL
XFILL_9_OAI21X1_172 BUFX2_36/A DFFSR_6/S FILL
XFILL_0_OAI22X1_56 BUFX2_37/A DFFSR_8/S FILL
XFILL_1_INVX1_261 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_1_XOR2X1_9 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_0_DFFSR_3 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_0_NAND2X1_231 BUFX2_37/A DFFSR_81/S FILL
XINVX1_73 BUFX2_10/Y BUFX2_19/gnd DFFSR_61/R DFFSR_54/S INVX1
XFILL_33_DFFSR_39 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_22_DFFSR_79 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_5_DFFSR_86 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_7_DFFSR_104 INVX1_4/gnd DFFSR_4/S FILL
XFILL_48_DFFSR_135 BUFX2_43/A DFFSR_97/S FILL
XFILL_8_NAND3X1_11 BUFX2_19/gnd DFFSR_54/S FILL
XINVX1_191 BUFX2_7/Y BUFX2_5/gnd DFFSR_158/R DFFSR_23/S INVX1
XFILL_7_NAND3X1_14 BUFX2_19/gnd DFFSR_52/S FILL
XFILL_38_DFFSR_138 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_4_INVX1_188 BUFX2_35/A DFFSR_97/S FILL
XFILL_28_DFFSR_141 INVX1_94/gnd DFFSR_25/S FILL
XFILL_1_NAND2X1_165 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_33_2_0 INVX1_8/gnd DFFSR_7/S FILL
XFILL_4_BUFX2_24 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_6_NAND3X1_17 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_18_DFFSR_144 INVX1_8/gnd DFFSR_5/S FILL
XFILL_24_DFFSR_7 INVX1_8/gnd DFFSR_7/S FILL
XFILL_4_CLKBUF1_9 BUFX2_17/gnd DFFSR_7/S FILL
XFILL_5_NAND3X1_20 BUFX2_37/A DFFSR_8/S FILL
XNAND3X1_17 INVX1_223/Y AOI22X1_4/B AOI21X1_3/B DFFSR_79/gnd NOR3X1_1/A DFFSR_45/S
+ NAND3X1
XFILL_41_DFFSR_46 BUFX2_36/A DFFSR_6/S FILL
XFILL_4_NAND3X1_23 BUFX2_37/A DFFSR_81/S FILL
XFILL_2_INVX1_80 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_3_NOR2X1_23 DFFSR_79/gnd DFFSR_45/S FILL
XFILL_31_4_1 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_30_DFFSR_86 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_13_DFFPOSX1_22 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_8_OAI21X1_202 BUFX2_35/A DFFSR_14/S FILL
XFILL_3_NAND3X1_26 BUFX2_7/gnd DFFSR_81/S FILL
XDFFSR_144 DFFSR_144/Q CLKBUF1_9/Y DFFSR_137/R DFFSR_5/S DFFSR_144/D INVX1_8/gnd DFFSR_5/S
+ DFFSR
XFILL_2_NAND3X1_29 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_2_INVX1_405 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_4_DFFSR_141 INVX1_94/gnd DFFSR_25/S FILL
XFILL_14_DFFSR_36 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_3_OAI22X1_11 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_45_DFFSR_172 BUFX2_37/A DFFSR_8/S FILL
XFILL_1_NAND3X1_32 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_2_OAI22X1_14 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_35_DFFSR_175 INVX1_23/gnd DFFSR_91/S FILL
XFILL_0_NAND3X1_35 BUFX2_35/A DFFSR_97/S FILL
XFILL_1_OAI22X1_17 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_0_OAI22X1_20 BUFX2_8/gnd DFFSR_25/S FILL
XFILL_9_OAI21X1_136 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_25_DFFSR_178 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_23_DFFPOSX1_11 INVX1_4/gnd DFFSR_4/S FILL
XFILL_45_DFFSR_3 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_15_DFFSR_181 INVX1_23/gnd DFFSR_186/S FILL
XFILL_1_INVX1_225 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_49_DFFSR_53 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_38_DFFSR_93 INVX1_2/gnd DFFSR_51/S FILL
XFILL_0_NAND2X1_195 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_11_DFFSR_83 BUFX2_19/gnd DFFSR_54/S FILL
XINVX1_37 BUFX2_10/Y INVX1_94/gnd DFFSR_31/R DFFSR_52/S INVX1
XFILL_22_DFFSR_43 INVX1_94/gnd DFFSR_25/S FILL
XDFFSR_90 DFFSR_90/Q CLKBUF1_2/Y DFFSR_89/R DFFSR_1/S DFFSR_90/D INVX1_2/gnd DFFSR_1/S
+ DFFSR
XFILL_5_DFFSR_50 DFFSR_73/gnd DFFSR_11/S FILL
XFILL_2_OAI21X1_8 BUFX2_36/A DFFSR_6/S FILL
XINVX1_155 DFFSR_137/Q INVX1_94/gnd INVX1_155/Y DFFSR_52/S INVX1
XFILL_38_DFFSR_102 INVX1_8/gnd DFFSR_7/S FILL
XFILL_28_DFFSR_105 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_1_DFFSR_178 DFFSR_1/gnd DFFSR_9/S FILL
XFILL_0_INVX1_5 INVX1_4/gnd DFFSR_51/S FILL
XFILL_7_OAI21X1_232 BUFX2_35/A DFFSR_97/S FILL
XFILL_18_DFFSR_108 INVX1_89/gnd DFFSR_2/S FILL
XFILL_1_NAND2X1_129 INVX1_4/gnd DFFSR_4/S FILL
XFILL_7_AND2X2_9 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_2_DFFSR_97 BUFX2_35/A DFFSR_97/S FILL
XFILL_41_DFFSR_10 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_2_INVX1_44 DFFSR_79/gnd DFFSR_36/S FILL
XFILL_30_DFFSR_50 DFFSR_73/gnd DFFSR_11/S FILL
XDFFSR_108 INVX1_122/A CLKBUF1_1/Y DFFSR_105/R DFFSR_2/S DFFSR_108/D INVX1_89/gnd
+ DFFSR_2/S DFFSR
XFILL_19_DFFSR_90 INVX1_2/gnd DFFSR_1/S FILL
XFILL_39_1_2 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_2_INVX1_369 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_8_OAI21X1_166 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_4_DFFSR_105 DFFSR_89/gnd DFFSR_186/S FILL
XFILL_1_BUFX2_35 BUFX2_35/A DFFSR_14/S FILL
XFILL_45_DFFSR_136 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_9_OAI21X1_100 INVX1_23/gnd DFFSR_91/S FILL
XFILL_11_DFFSR_1 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_35_DFFSR_139 DFFSR_3/gnd DFFSR_4/S FILL
XFILL_1_INVX1_189 BUFX2_35/A DFFSR_14/S FILL
XFILL_25_DFFSR_142 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_49_DFFSR_17 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_15_DFFSR_145 INVX1_23/gnd DFFSR_186/S FILL
XFILL_27_DFFSR_97 BUFX2_35/A DFFSR_97/S FILL
XFILL_38_DFFSR_57 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_40_3 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_0_NAND2X1_159 BUFX2_43/A DFFSR_97/S FILL
XDFFSR_54 DFFSR_54/Q INVX1_1/A DFFSR_54/R DFFSR_54/S DFFSR_54/D BUFX2_7/gnd DFFSR_81/S
+ DFFSR
XFILL_5_DFFSR_14 BUFX2_35/A DFFSR_14/S FILL
XFILL_0_NOR2X1_24 BUFX2_8/gnd DFFSR_10/S FILL
XFILL_6_OAI21X1_262 INVX1_89/gnd DFFSR_36/S FILL
XFILL_11_DFFSR_47 DFFSR_5/gnd DFFSR_2/S FILL
XINVX1_119 DFFSR_105/Q BUFX2_6/gnd INVX1_119/Y DFFSR_14/S INVX1
XFILL_1_DFFSR_142 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_8_NAND3X1_112 DFFSR_71/gnd DFFSR_10/S FILL
XFILL_42_DFFSR_173 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_12_DFFPOSX1_16 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_7_OAI21X1_196 INVX1_94/gnd DFFSR_25/S FILL
XFILL_32_DFFSR_176 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_46_DFFSR_64 BUFX2_16/gnd DFFSR_11/S FILL
XFILL_22_DFFSR_179 INVX1_2/gnd DFFSR_1/S FILL
XFILL_30_DFFSR_14 BUFX2_35/A DFFSR_14/S FILL
XFILL_2_DFFSR_61 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_19_DFFSR_54 BUFX2_7/gnd DFFSR_81/S FILL
XFILL_12_DFFSR_182 INVX1_89/gnd DFFSR_36/S FILL
XFILL_8_OAI21X1_130 INVX1_4/gnd DFFSR_4/S FILL
XFILL_2_INVX1_333 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_45_DFFSR_100 INVX1_23/gnd DFFSR_186/S FILL
XFILL_2_DFFPOSX1_27 DFFSR_71/gnd DFFSR_45/S FILL
XFILL_35_DFFSR_103 INVX1_8/gnd DFFSR_7/S FILL
XFILL_8_DFFSR_176 BUFX2_16/gnd DFFSR_65/S FILL
XFILL_25_DFFSR_106 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_15_DFFSR_109 BUFX2_6/gnd DFFSR_14/S FILL
XFILL_27_DFFSR_61 BUFX2_5/gnd DFFSR_6/S FILL
XFILL_1_INVX1_153 DFFSR_5/gnd DFFSR_2/S FILL
XFILL_38_DFFSR_21 INVX1_2/gnd DFFSR_1/S FILL
XFILL_6_OAI21X1_226 BUFX2_6/gnd DFFSR_91/S FILL
XFILL_0_NAND2X1_123 BUFX2_6/gnd DFFSR_14/S FILL
XDFFSR_18 INVX1_21/A DFFSR_24/CLK DFFSR_20/R DFFSR_9/S DFFSR_18/D DFFSR_9/gnd DFFSR_9/S
+ DFFSR
XFILL_11_DFFSR_11 BUFX2_16/gnd DFFSR_11/S FILL
XOAI21X1_262 AOI21X1_46/C AND2X2_17/Y INVX1_436/A INVX1_89/gnd NOR2X1_51/B DFFSR_36/S
+ OAI21X1
XFILL_1_DFFSR_106 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_35_DFFSR_68 BUFX2_35/A DFFSR_14/S FILL
XFILL_42_DFFSR_137 BUFX2_7/gnd DFFSR_54/S FILL
XFILL_46_DFFSR_28 BUFX2_19/gnd DFFSR_54/S FILL
XFILL_7_OAI21X1_160 DFFSR_73/gnd DFFSR_57/S FILL
XFILL_32_DFFSR_140 DFFSR_71/gnd DFFSR_10/S FILL
.ends

