module mips (clk, rst, MemData, MemWrite, MemRead, MemWriteData, MemAddr);

input clk;
input rst;
output MemWrite;
output MemRead;
input [31:0] MemData;
output [31:0] MemWriteData;
output [31:0] MemAddr;

wire vdd = 1'b1;
wire gnd = 1'b0;

BUFX2 BUFX2_1 ( .A(datapath_1_Instr_23_bF_buf10_), .Y(datapath_1_Instr_23_bF_buf10_bF_buf3_) );
BUFX2 BUFX2_2 ( .A(datapath_1_Instr_23_bF_buf10_), .Y(datapath_1_Instr_23_bF_buf10_bF_buf2_) );
BUFX2 BUFX2_3 ( .A(datapath_1_Instr_23_bF_buf10_), .Y(datapath_1_Instr_23_bF_buf10_bF_buf1_) );
BUFX2 BUFX2_4 ( .A(datapath_1_Instr_23_bF_buf10_), .Y(datapath_1_Instr_23_bF_buf10_bF_buf0_) );
BUFX2 BUFX2_5 ( .A(datapath_1_Instr_17_), .Y(datapath_1_Instr_17__hier0_bF_buf6) );
BUFX2 BUFX2_6 ( .A(datapath_1_Instr_17_), .Y(datapath_1_Instr_17__hier0_bF_buf5) );
BUFX2 BUFX2_7 ( .A(datapath_1_Instr_17_), .Y(datapath_1_Instr_17__hier0_bF_buf4) );
BUFX2 BUFX2_8 ( .A(datapath_1_Instr_17_), .Y(datapath_1_Instr_17__hier0_bF_buf3) );
BUFX2 BUFX2_9 ( .A(datapath_1_Instr_17_), .Y(datapath_1_Instr_17__hier0_bF_buf2) );
BUFX2 BUFX2_10 ( .A(datapath_1_Instr_17_), .Y(datapath_1_Instr_17__hier0_bF_buf1) );
BUFX2 BUFX2_11 ( .A(datapath_1_Instr_17_), .Y(datapath_1_Instr_17__hier0_bF_buf0) );
BUFX2 BUFX2_12 ( .A(clk), .Y(clk_hier0_bF_buf9) );
BUFX2 BUFX2_13 ( .A(clk), .Y(clk_hier0_bF_buf8) );
BUFX2 BUFX2_14 ( .A(clk), .Y(clk_hier0_bF_buf7) );
BUFX2 BUFX2_15 ( .A(clk), .Y(clk_hier0_bF_buf6) );
BUFX2 BUFX2_16 ( .A(clk), .Y(clk_hier0_bF_buf5) );
BUFX2 BUFX2_17 ( .A(clk), .Y(clk_hier0_bF_buf4) );
BUFX2 BUFX2_18 ( .A(clk), .Y(clk_hier0_bF_buf3) );
BUFX2 BUFX2_19 ( .A(clk), .Y(clk_hier0_bF_buf2) );
BUFX2 BUFX2_20 ( .A(clk), .Y(clk_hier0_bF_buf1) );
BUFX2 BUFX2_21 ( .A(clk), .Y(clk_hier0_bF_buf0) );
BUFX2 BUFX2_22 ( .A(datapath_1_Instr_23_bF_buf9_), .Y(datapath_1_Instr_23_bF_buf9_bF_buf3_) );
BUFX2 BUFX2_23 ( .A(datapath_1_Instr_23_bF_buf9_), .Y(datapath_1_Instr_23_bF_buf9_bF_buf2_) );
BUFX2 BUFX2_24 ( .A(datapath_1_Instr_23_bF_buf9_), .Y(datapath_1_Instr_23_bF_buf9_bF_buf1_) );
BUFX2 BUFX2_25 ( .A(datapath_1_Instr_23_bF_buf9_), .Y(datapath_1_Instr_23_bF_buf9_bF_buf0_) );
BUFX2 BUFX2_26 ( .A(datapath_1_Instr_23_bF_buf6_), .Y(datapath_1_Instr_23_bF_buf6_bF_buf3_) );
BUFX2 BUFX2_27 ( .A(datapath_1_Instr_23_bF_buf6_), .Y(datapath_1_Instr_23_bF_buf6_bF_buf2_) );
BUFX2 BUFX2_28 ( .A(datapath_1_Instr_23_bF_buf6_), .Y(datapath_1_Instr_23_bF_buf6_bF_buf1_) );
BUFX2 BUFX2_29 ( .A(datapath_1_Instr_23_bF_buf6_), .Y(datapath_1_Instr_23_bF_buf6_bF_buf0_) );
BUFX2 BUFX2_30 ( .A(datapath_1_Instr_23_bF_buf3_), .Y(datapath_1_Instr_23_bF_buf3_bF_buf3_) );
BUFX2 BUFX2_31 ( .A(datapath_1_Instr_23_bF_buf3_), .Y(datapath_1_Instr_23_bF_buf3_bF_buf2_) );
BUFX2 BUFX2_32 ( .A(datapath_1_Instr_23_bF_buf3_), .Y(datapath_1_Instr_23_bF_buf3_bF_buf1_) );
BUFX2 BUFX2_33 ( .A(datapath_1_Instr_23_bF_buf3_), .Y(datapath_1_Instr_23_bF_buf3_bF_buf0_) );
BUFX2 BUFX2_34 ( .A(datapath_1_Instr_23_bF_buf15_), .Y(datapath_1_Instr_23_bF_buf15_bF_buf3_) );
BUFX2 BUFX2_35 ( .A(datapath_1_Instr_23_bF_buf15_), .Y(datapath_1_Instr_23_bF_buf15_bF_buf2_) );
BUFX2 BUFX2_36 ( .A(datapath_1_Instr_23_bF_buf15_), .Y(datapath_1_Instr_23_bF_buf15_bF_buf1_) );
BUFX2 BUFX2_37 ( .A(datapath_1_Instr_23_bF_buf15_), .Y(datapath_1_Instr_23_bF_buf15_bF_buf0_) );
BUFX2 BUFX2_38 ( .A(datapath_1_Instr_23_bF_buf12_), .Y(datapath_1_Instr_23_bF_buf12_bF_buf3_) );
BUFX2 BUFX2_39 ( .A(datapath_1_Instr_23_bF_buf12_), .Y(datapath_1_Instr_23_bF_buf12_bF_buf2_) );
BUFX2 BUFX2_40 ( .A(datapath_1_Instr_23_bF_buf12_), .Y(datapath_1_Instr_23_bF_buf12_bF_buf1_) );
BUFX2 BUFX2_41 ( .A(datapath_1_Instr_23_bF_buf12_), .Y(datapath_1_Instr_23_bF_buf12_bF_buf0_) );
BUFX2 BUFX2_42 ( .A(datapath_1_Instr_22_), .Y(datapath_1_Instr_22__hier0_bF_buf6) );
BUFX2 BUFX2_43 ( .A(datapath_1_Instr_22_), .Y(datapath_1_Instr_22__hier0_bF_buf5) );
BUFX2 BUFX2_44 ( .A(datapath_1_Instr_22_), .Y(datapath_1_Instr_22__hier0_bF_buf4) );
BUFX2 BUFX2_45 ( .A(datapath_1_Instr_22_), .Y(datapath_1_Instr_22__hier0_bF_buf3) );
BUFX2 BUFX2_46 ( .A(datapath_1_Instr_22_), .Y(datapath_1_Instr_22__hier0_bF_buf2) );
BUFX2 BUFX2_47 ( .A(datapath_1_Instr_22_), .Y(datapath_1_Instr_22__hier0_bF_buf1) );
BUFX2 BUFX2_48 ( .A(datapath_1_Instr_22_), .Y(datapath_1_Instr_22__hier0_bF_buf0) );
BUFX2 BUFX2_49 ( .A(datapath_1_Instr_16_), .Y(datapath_1_Instr_16__hier0_bF_buf6) );
BUFX2 BUFX2_50 ( .A(datapath_1_Instr_16_), .Y(datapath_1_Instr_16__hier0_bF_buf5) );
BUFX2 BUFX2_51 ( .A(datapath_1_Instr_16_), .Y(datapath_1_Instr_16__hier0_bF_buf4) );
BUFX2 BUFX2_52 ( .A(datapath_1_Instr_16_), .Y(datapath_1_Instr_16__hier0_bF_buf3) );
BUFX2 BUFX2_53 ( .A(datapath_1_Instr_16_), .Y(datapath_1_Instr_16__hier0_bF_buf2) );
BUFX2 BUFX2_54 ( .A(datapath_1_Instr_16_), .Y(datapath_1_Instr_16__hier0_bF_buf1) );
BUFX2 BUFX2_55 ( .A(datapath_1_Instr_16_), .Y(datapath_1_Instr_16__hier0_bF_buf0) );
BUFX2 BUFX2_56 ( .A(_5265_), .Y(_5265__hier0_bF_buf8) );
BUFX2 BUFX2_57 ( .A(_5265_), .Y(_5265__hier0_bF_buf7) );
BUFX2 BUFX2_58 ( .A(_5265_), .Y(_5265__hier0_bF_buf6) );
BUFX2 BUFX2_59 ( .A(_5265_), .Y(_5265__hier0_bF_buf5) );
BUFX2 BUFX2_60 ( .A(_5265_), .Y(_5265__hier0_bF_buf4) );
BUFX2 BUFX2_61 ( .A(_5265_), .Y(_5265__hier0_bF_buf3) );
BUFX2 BUFX2_62 ( .A(_5265_), .Y(_5265__hier0_bF_buf2) );
BUFX2 BUFX2_63 ( .A(_5265_), .Y(_5265__hier0_bF_buf1) );
BUFX2 BUFX2_64 ( .A(_5265_), .Y(_5265__hier0_bF_buf0) );
BUFX2 BUFX2_65 ( .A(_1890_), .Y(_1890__hier0_bF_buf5) );
BUFX2 BUFX2_66 ( .A(_1890_), .Y(_1890__hier0_bF_buf4) );
BUFX2 BUFX2_67 ( .A(_1890_), .Y(_1890__hier0_bF_buf3) );
BUFX2 BUFX2_68 ( .A(_1890_), .Y(_1890__hier0_bF_buf2) );
BUFX2 BUFX2_69 ( .A(_1890_), .Y(_1890__hier0_bF_buf1) );
BUFX2 BUFX2_70 ( .A(_1890_), .Y(_1890__hier0_bF_buf0) );
BUFX2 BUFX2_71 ( .A(datapath_1_Instr_23_bF_buf8_), .Y(datapath_1_Instr_23_bF_buf8_bF_buf3_) );
BUFX2 BUFX2_72 ( .A(datapath_1_Instr_23_bF_buf8_), .Y(datapath_1_Instr_23_bF_buf8_bF_buf2_) );
BUFX2 BUFX2_73 ( .A(datapath_1_Instr_23_bF_buf8_), .Y(datapath_1_Instr_23_bF_buf8_bF_buf1_) );
BUFX2 BUFX2_74 ( .A(datapath_1_Instr_23_bF_buf8_), .Y(datapath_1_Instr_23_bF_buf8_bF_buf0_) );
BUFX2 BUFX2_75 ( .A(datapath_1_Instr_23_bF_buf5_), .Y(datapath_1_Instr_23_bF_buf5_bF_buf3_) );
BUFX2 BUFX2_76 ( .A(datapath_1_Instr_23_bF_buf5_), .Y(datapath_1_Instr_23_bF_buf5_bF_buf2_) );
BUFX2 BUFX2_77 ( .A(datapath_1_Instr_23_bF_buf5_), .Y(datapath_1_Instr_23_bF_buf5_bF_buf1_) );
BUFX2 BUFX2_78 ( .A(datapath_1_Instr_23_bF_buf5_), .Y(datapath_1_Instr_23_bF_buf5_bF_buf0_) );
BUFX2 BUFX2_79 ( .A(datapath_1_Instr_23_bF_buf2_), .Y(datapath_1_Instr_23_bF_buf2_bF_buf3_) );
BUFX2 BUFX2_80 ( .A(datapath_1_Instr_23_bF_buf2_), .Y(datapath_1_Instr_23_bF_buf2_bF_buf2_) );
BUFX2 BUFX2_81 ( .A(datapath_1_Instr_23_bF_buf2_), .Y(datapath_1_Instr_23_bF_buf2_bF_buf1_) );
BUFX2 BUFX2_82 ( .A(datapath_1_Instr_23_bF_buf2_), .Y(datapath_1_Instr_23_bF_buf2_bF_buf0_) );
BUFX2 BUFX2_83 ( .A(datapath_1_Instr_23_bF_buf14_), .Y(datapath_1_Instr_23_bF_buf14_bF_buf3_) );
BUFX2 BUFX2_84 ( .A(datapath_1_Instr_23_bF_buf14_), .Y(datapath_1_Instr_23_bF_buf14_bF_buf2_) );
BUFX2 BUFX2_85 ( .A(datapath_1_Instr_23_bF_buf14_), .Y(datapath_1_Instr_23_bF_buf14_bF_buf1_) );
BUFX2 BUFX2_86 ( .A(datapath_1_Instr_23_bF_buf14_), .Y(datapath_1_Instr_23_bF_buf14_bF_buf0_) );
BUFX2 BUFX2_87 ( .A(datapath_1_Instr_23_bF_buf11_), .Y(datapath_1_Instr_23_bF_buf11_bF_buf3_) );
BUFX2 BUFX2_88 ( .A(datapath_1_Instr_23_bF_buf11_), .Y(datapath_1_Instr_23_bF_buf11_bF_buf2_) );
BUFX2 BUFX2_89 ( .A(datapath_1_Instr_23_bF_buf11_), .Y(datapath_1_Instr_23_bF_buf11_bF_buf1_) );
BUFX2 BUFX2_90 ( .A(datapath_1_Instr_23_bF_buf11_), .Y(datapath_1_Instr_23_bF_buf11_bF_buf0_) );
BUFX2 BUFX2_91 ( .A(datapath_1_Instr_21_), .Y(datapath_1_Instr_21__hier0_bF_buf6) );
BUFX2 BUFX2_92 ( .A(datapath_1_Instr_21_), .Y(datapath_1_Instr_21__hier0_bF_buf5) );
BUFX2 BUFX2_93 ( .A(datapath_1_Instr_21_), .Y(datapath_1_Instr_21__hier0_bF_buf4) );
BUFX2 BUFX2_94 ( .A(datapath_1_Instr_21_), .Y(datapath_1_Instr_21__hier0_bF_buf3) );
BUFX2 BUFX2_95 ( .A(datapath_1_Instr_21_), .Y(datapath_1_Instr_21__hier0_bF_buf2) );
BUFX2 BUFX2_96 ( .A(datapath_1_Instr_21_), .Y(datapath_1_Instr_21__hier0_bF_buf1) );
BUFX2 BUFX2_97 ( .A(datapath_1_Instr_21_), .Y(datapath_1_Instr_21__hier0_bF_buf0) );
BUFX2 BUFX2_98 ( .A(datapath_1_Instr_18_), .Y(datapath_1_Instr_18__hier0_bF_buf5) );
BUFX2 BUFX2_99 ( .A(datapath_1_Instr_18_), .Y(datapath_1_Instr_18__hier0_bF_buf4) );
BUFX2 BUFX2_100 ( .A(datapath_1_Instr_18_), .Y(datapath_1_Instr_18__hier0_bF_buf3) );
BUFX2 BUFX2_101 ( .A(datapath_1_Instr_18_), .Y(datapath_1_Instr_18__hier0_bF_buf2) );
BUFX2 BUFX2_102 ( .A(datapath_1_Instr_18_), .Y(datapath_1_Instr_18__hier0_bF_buf1) );
BUFX2 BUFX2_103 ( .A(datapath_1_Instr_18_), .Y(datapath_1_Instr_18__hier0_bF_buf0) );
BUFX2 BUFX2_104 ( .A(_3588_), .Y(_3588__hier0_bF_buf5) );
BUFX2 BUFX2_105 ( .A(_3588_), .Y(_3588__hier0_bF_buf4) );
BUFX2 BUFX2_106 ( .A(_3588_), .Y(_3588__hier0_bF_buf3) );
BUFX2 BUFX2_107 ( .A(_3588_), .Y(_3588__hier0_bF_buf2) );
BUFX2 BUFX2_108 ( .A(_3588_), .Y(_3588__hier0_bF_buf1) );
BUFX2 BUFX2_109 ( .A(_3588_), .Y(_3588__hier0_bF_buf0) );
BUFX2 BUFX2_110 ( .A(datapath_1_Instr_23_bF_buf7_), .Y(datapath_1_Instr_23_bF_buf7_bF_buf3_) );
BUFX2 BUFX2_111 ( .A(datapath_1_Instr_23_bF_buf7_), .Y(datapath_1_Instr_23_bF_buf7_bF_buf2_) );
BUFX2 BUFX2_112 ( .A(datapath_1_Instr_23_bF_buf7_), .Y(datapath_1_Instr_23_bF_buf7_bF_buf1_) );
BUFX2 BUFX2_113 ( .A(datapath_1_Instr_23_bF_buf7_), .Y(datapath_1_Instr_23_bF_buf7_bF_buf0_) );
BUFX2 BUFX2_114 ( .A(datapath_1_Instr_23_bF_buf4_), .Y(datapath_1_Instr_23_bF_buf4_bF_buf3_) );
BUFX2 BUFX2_115 ( .A(datapath_1_Instr_23_bF_buf4_), .Y(datapath_1_Instr_23_bF_buf4_bF_buf2_) );
BUFX2 BUFX2_116 ( .A(datapath_1_Instr_23_bF_buf4_), .Y(datapath_1_Instr_23_bF_buf4_bF_buf1_) );
BUFX2 BUFX2_117 ( .A(datapath_1_Instr_23_bF_buf4_), .Y(datapath_1_Instr_23_bF_buf4_bF_buf0_) );
BUFX2 BUFX2_118 ( .A(datapath_1_Instr_23_bF_buf13_), .Y(datapath_1_Instr_23_bF_buf13_bF_buf3_) );
BUFX2 BUFX2_119 ( .A(datapath_1_Instr_23_bF_buf13_), .Y(datapath_1_Instr_23_bF_buf13_bF_buf2_) );
BUFX2 BUFX2_120 ( .A(datapath_1_Instr_23_bF_buf13_), .Y(datapath_1_Instr_23_bF_buf13_bF_buf1_) );
BUFX2 BUFX2_121 ( .A(datapath_1_Instr_23_bF_buf13_), .Y(datapath_1_Instr_23_bF_buf13_bF_buf0_) );
BUFX2 BUFX2_122 ( .A(_5278_), .Y(_5278__bF_buf4) );
BUFX2 BUFX2_123 ( .A(_5278_), .Y(_5278__bF_buf3) );
BUFX2 BUFX2_124 ( .A(_5278_), .Y(_5278__bF_buf2) );
BUFX2 BUFX2_125 ( .A(_5278_), .Y(_5278__bF_buf1) );
BUFX2 BUFX2_126 ( .A(_5278_), .Y(_5278__bF_buf0) );
BUFX2 BUFX2_127 ( .A(_5334_), .Y(_5334__bF_buf4) );
BUFX2 BUFX2_128 ( .A(_5334_), .Y(_5334__bF_buf3) );
BUFX2 BUFX2_129 ( .A(_5334_), .Y(_5334__bF_buf2) );
BUFX2 BUFX2_130 ( .A(_5334_), .Y(_5334__bF_buf1) );
BUFX2 BUFX2_131 ( .A(_5334_), .Y(_5334__bF_buf0) );
BUFX2 BUFX2_132 ( .A(_5275_), .Y(_5275__bF_buf7) );
BUFX2 BUFX2_133 ( .A(_5275_), .Y(_5275__bF_buf6) );
BUFX2 BUFX2_134 ( .A(_5275_), .Y(_5275__bF_buf5) );
BUFX2 BUFX2_135 ( .A(_5275_), .Y(_5275__bF_buf4) );
BUFX2 BUFX2_136 ( .A(_5275_), .Y(_5275__bF_buf3) );
BUFX2 BUFX2_137 ( .A(_5275_), .Y(_5275__bF_buf2) );
BUFX2 BUFX2_138 ( .A(_5275_), .Y(_5275__bF_buf1) );
BUFX2 BUFX2_139 ( .A(_5275_), .Y(_5275__bF_buf0) );
BUFX2 BUFX2_140 ( .A(_3570_), .Y(_3570__bF_buf4) );
BUFX2 BUFX2_141 ( .A(_3570_), .Y(_3570__bF_buf3) );
BUFX2 BUFX2_142 ( .A(_3570_), .Y(_3570__bF_buf2) );
BUFX2 BUFX2_143 ( .A(_3570_), .Y(_3570__bF_buf1) );
BUFX2 BUFX2_144 ( .A(_3570_), .Y(_3570__bF_buf0) );
BUFX2 BUFX2_145 ( .A(datapath_1_Instr_23_), .Y(datapath_1_Instr_23_bF_buf15_) );
BUFX2 BUFX2_146 ( .A(datapath_1_Instr_23_), .Y(datapath_1_Instr_23_bF_buf14_) );
BUFX2 BUFX2_147 ( .A(datapath_1_Instr_23_), .Y(datapath_1_Instr_23_bF_buf13_) );
BUFX2 BUFX2_148 ( .A(datapath_1_Instr_23_), .Y(datapath_1_Instr_23_bF_buf12_) );
BUFX2 BUFX2_149 ( .A(datapath_1_Instr_23_), .Y(datapath_1_Instr_23_bF_buf11_) );
BUFX2 BUFX2_150 ( .A(datapath_1_Instr_23_), .Y(datapath_1_Instr_23_bF_buf10_) );
BUFX2 BUFX2_151 ( .A(datapath_1_Instr_23_), .Y(datapath_1_Instr_23_bF_buf9_) );
BUFX2 BUFX2_152 ( .A(datapath_1_Instr_23_), .Y(datapath_1_Instr_23_bF_buf8_) );
BUFX2 BUFX2_153 ( .A(datapath_1_Instr_23_), .Y(datapath_1_Instr_23_bF_buf7_) );
BUFX2 BUFX2_154 ( .A(datapath_1_Instr_23_), .Y(datapath_1_Instr_23_bF_buf6_) );
BUFX2 BUFX2_155 ( .A(datapath_1_Instr_23_), .Y(datapath_1_Instr_23_bF_buf5_) );
BUFX2 BUFX2_156 ( .A(datapath_1_Instr_23_), .Y(datapath_1_Instr_23_bF_buf4_) );
BUFX2 BUFX2_157 ( .A(datapath_1_Instr_23_), .Y(datapath_1_Instr_23_bF_buf3_) );
BUFX2 BUFX2_158 ( .A(datapath_1_Instr_23_), .Y(datapath_1_Instr_23_bF_buf2_) );
BUFX2 BUFX2_159 ( .A(datapath_1_Instr_23_), .Y(datapath_1_Instr_23_bF_buf1_) );
BUFX2 BUFX2_160 ( .A(datapath_1_Instr_23_), .Y(datapath_1_Instr_23_bF_buf0_) );
BUFX2 BUFX2_161 ( .A(_3567_), .Y(_3567__bF_buf10) );
BUFX2 BUFX2_162 ( .A(_3567_), .Y(_3567__bF_buf9) );
BUFX2 BUFX2_163 ( .A(_3567_), .Y(_3567__bF_buf8) );
BUFX2 BUFX2_164 ( .A(_3567_), .Y(_3567__bF_buf7) );
BUFX2 BUFX2_165 ( .A(_3567_), .Y(_3567__bF_buf6) );
BUFX2 BUFX2_166 ( .A(_3567_), .Y(_3567__bF_buf5) );
BUFX2 BUFX2_167 ( .A(_3567_), .Y(_3567__bF_buf4) );
BUFX2 BUFX2_168 ( .A(_3567_), .Y(_3567__bF_buf3) );
BUFX2 BUFX2_169 ( .A(_3567_), .Y(_3567__bF_buf2) );
BUFX2 BUFX2_170 ( .A(_3567_), .Y(_3567__bF_buf1) );
BUFX2 BUFX2_171 ( .A(_3567_), .Y(_3567__bF_buf0) );
BUFX2 BUFX2_172 ( .A(_5713_), .Y(_5713__bF_buf7) );
BUFX2 BUFX2_173 ( .A(_5713_), .Y(_5713__bF_buf6) );
BUFX2 BUFX2_174 ( .A(_5713_), .Y(_5713__bF_buf5) );
BUFX2 BUFX2_175 ( .A(_5713_), .Y(_5713__bF_buf4) );
BUFX2 BUFX2_176 ( .A(_5713_), .Y(_5713__bF_buf3) );
BUFX2 BUFX2_177 ( .A(_5713_), .Y(_5713__bF_buf2) );
BUFX2 BUFX2_178 ( .A(_5713_), .Y(_5713__bF_buf1) );
BUFX2 BUFX2_179 ( .A(_5713_), .Y(_5713__bF_buf0) );
BUFX2 BUFX2_180 ( .A(_6918_), .Y(_6918__bF_buf4) );
BUFX2 BUFX2_181 ( .A(_6918_), .Y(_6918__bF_buf3) );
BUFX2 BUFX2_182 ( .A(_6918_), .Y(_6918__bF_buf2) );
BUFX2 BUFX2_183 ( .A(_6918_), .Y(_6918__bF_buf1) );
BUFX2 BUFX2_184 ( .A(_6918_), .Y(_6918__bF_buf0) );
BUFX2 BUFX2_185 ( .A(_6116_), .Y(_6116__bF_buf7) );
BUFX2 BUFX2_186 ( .A(_6116_), .Y(_6116__bF_buf6) );
BUFX2 BUFX2_187 ( .A(_6116_), .Y(_6116__bF_buf5) );
BUFX2 BUFX2_188 ( .A(_6116_), .Y(_6116__bF_buf4) );
BUFX2 BUFX2_189 ( .A(_6116_), .Y(_6116__bF_buf3) );
BUFX2 BUFX2_190 ( .A(_6116_), .Y(_6116__bF_buf2) );
BUFX2 BUFX2_191 ( .A(_6116_), .Y(_6116__bF_buf1) );
BUFX2 BUFX2_192 ( .A(_6116_), .Y(_6116__bF_buf0) );
BUFX2 BUFX2_193 ( .A(_5980_), .Y(_5980__bF_buf7) );
BUFX2 BUFX2_194 ( .A(_5980_), .Y(_5980__bF_buf6) );
BUFX2 BUFX2_195 ( .A(_5980_), .Y(_5980__bF_buf5) );
BUFX2 BUFX2_196 ( .A(_5980_), .Y(_5980__bF_buf4) );
BUFX2 BUFX2_197 ( .A(_5980_), .Y(_5980__bF_buf3) );
BUFX2 BUFX2_198 ( .A(_5980_), .Y(_5980__bF_buf2) );
BUFX2 BUFX2_199 ( .A(_5980_), .Y(_5980__bF_buf1) );
BUFX2 BUFX2_200 ( .A(_5980_), .Y(_5980__bF_buf0) );
BUFX2 BUFX2_201 ( .A(_256_), .Y(_256__bF_buf3) );
BUFX2 BUFX2_202 ( .A(_256_), .Y(_256__bF_buf2) );
BUFX2 BUFX2_203 ( .A(_256_), .Y(_256__bF_buf1) );
BUFX2 BUFX2_204 ( .A(_256_), .Y(_256__bF_buf0) );
BUFX2 BUFX2_205 ( .A(_6383_), .Y(_6383__bF_buf4) );
BUFX2 BUFX2_206 ( .A(_6383_), .Y(_6383__bF_buf3) );
BUFX2 BUFX2_207 ( .A(_6383_), .Y(_6383__bF_buf2) );
BUFX2 BUFX2_208 ( .A(_6383_), .Y(_6383__bF_buf1) );
BUFX2 BUFX2_209 ( .A(_6383_), .Y(_6383__bF_buf0) );
BUFX2 BUFX2_210 ( .A(_5272_), .Y(_5272__bF_buf5) );
BUFX2 BUFX2_211 ( .A(_5272_), .Y(_5272__bF_buf4) );
BUFX2 BUFX2_212 ( .A(_5272_), .Y(_5272__bF_buf3) );
BUFX2 BUFX2_213 ( .A(_5272_), .Y(_5272__bF_buf2) );
BUFX2 BUFX2_214 ( .A(_5272_), .Y(_5272__bF_buf1) );
BUFX2 BUFX2_215 ( .A(_5272_), .Y(_5272__bF_buf0) );
BUFX2 BUFX2_216 ( .A(_5328_), .Y(_5328__bF_buf4) );
BUFX2 BUFX2_217 ( .A(_5328_), .Y(_5328__bF_buf3) );
BUFX2 BUFX2_218 ( .A(_5328_), .Y(_5328__bF_buf2) );
BUFX2 BUFX2_219 ( .A(_5328_), .Y(_5328__bF_buf1) );
BUFX2 BUFX2_220 ( .A(_5328_), .Y(_5328__bF_buf0) );
BUFX2 BUFX2_221 ( .A(datapath_1_Instr_20_), .Y(datapath_1_Instr_20_bF_buf5_) );
BUFX2 BUFX2_222 ( .A(datapath_1_Instr_20_), .Y(datapath_1_Instr_20_bF_buf4_) );
BUFX2 BUFX2_223 ( .A(datapath_1_Instr_20_), .Y(datapath_1_Instr_20_bF_buf3_) );
BUFX2 BUFX2_224 ( .A(datapath_1_Instr_20_), .Y(datapath_1_Instr_20_bF_buf2_) );
BUFX2 BUFX2_225 ( .A(datapath_1_Instr_20_), .Y(datapath_1_Instr_20_bF_buf1_) );
BUFX2 BUFX2_226 ( .A(datapath_1_Instr_20_), .Y(datapath_1_Instr_20_bF_buf0_) );
BUFX2 BUFX2_227 ( .A(datapath_1_Instr_17__hier0_bF_buf3), .Y(datapath_1_Instr_17_bF_buf50_) );
BUFX2 BUFX2_228 ( .A(datapath_1_Instr_17__hier0_bF_buf1), .Y(datapath_1_Instr_17_bF_buf49_) );
BUFX2 BUFX2_229 ( .A(datapath_1_Instr_17__hier0_bF_buf1), .Y(datapath_1_Instr_17_bF_buf48_) );
BUFX2 BUFX2_230 ( .A(datapath_1_Instr_17__hier0_bF_buf1), .Y(datapath_1_Instr_17_bF_buf47_) );
BUFX2 BUFX2_231 ( .A(datapath_1_Instr_17__hier0_bF_buf4), .Y(datapath_1_Instr_17_bF_buf46_) );
BUFX2 BUFX2_232 ( .A(datapath_1_Instr_17__hier0_bF_buf5), .Y(datapath_1_Instr_17_bF_buf45_) );
BUFX2 BUFX2_233 ( .A(datapath_1_Instr_17__hier0_bF_buf5), .Y(datapath_1_Instr_17_bF_buf44_) );
BUFX2 BUFX2_234 ( .A(datapath_1_Instr_17__hier0_bF_buf1), .Y(datapath_1_Instr_17_bF_buf43_) );
BUFX2 BUFX2_235 ( .A(datapath_1_Instr_17__hier0_bF_buf5), .Y(datapath_1_Instr_17_bF_buf42_) );
BUFX2 BUFX2_236 ( .A(datapath_1_Instr_17__hier0_bF_buf4), .Y(datapath_1_Instr_17_bF_buf41_) );
BUFX2 BUFX2_237 ( .A(datapath_1_Instr_17__hier0_bF_buf5), .Y(datapath_1_Instr_17_bF_buf40_) );
BUFX2 BUFX2_238 ( .A(datapath_1_Instr_17__hier0_bF_buf5), .Y(datapath_1_Instr_17_bF_buf39_) );
BUFX2 BUFX2_239 ( .A(datapath_1_Instr_17__hier0_bF_buf1), .Y(datapath_1_Instr_17_bF_buf38_) );
BUFX2 BUFX2_240 ( .A(datapath_1_Instr_17__hier0_bF_buf4), .Y(datapath_1_Instr_17_bF_buf37_) );
BUFX2 BUFX2_241 ( .A(datapath_1_Instr_17__hier0_bF_buf4), .Y(datapath_1_Instr_17_bF_buf36_) );
BUFX2 BUFX2_242 ( .A(datapath_1_Instr_17__hier0_bF_buf4), .Y(datapath_1_Instr_17_bF_buf35_) );
BUFX2 BUFX2_243 ( .A(datapath_1_Instr_17__hier0_bF_buf1), .Y(datapath_1_Instr_17_bF_buf34_) );
BUFX2 BUFX2_244 ( .A(datapath_1_Instr_17__hier0_bF_buf5), .Y(datapath_1_Instr_17_bF_buf33_) );
BUFX2 BUFX2_245 ( .A(datapath_1_Instr_17__hier0_bF_buf3), .Y(datapath_1_Instr_17_bF_buf32_) );
BUFX2 BUFX2_246 ( .A(datapath_1_Instr_17__hier0_bF_buf4), .Y(datapath_1_Instr_17_bF_buf31_) );
BUFX2 BUFX2_247 ( .A(datapath_1_Instr_17__hier0_bF_buf6), .Y(datapath_1_Instr_17_bF_buf30_) );
BUFX2 BUFX2_248 ( .A(datapath_1_Instr_17__hier0_bF_buf5), .Y(datapath_1_Instr_17_bF_buf29_) );
BUFX2 BUFX2_249 ( .A(datapath_1_Instr_17__hier0_bF_buf3), .Y(datapath_1_Instr_17_bF_buf28_) );
BUFX2 BUFX2_250 ( .A(datapath_1_Instr_17__hier0_bF_buf6), .Y(datapath_1_Instr_17_bF_buf27_) );
BUFX2 BUFX2_251 ( .A(datapath_1_Instr_17__hier0_bF_buf5), .Y(datapath_1_Instr_17_bF_buf26_) );
BUFX2 BUFX2_252 ( .A(datapath_1_Instr_17__hier0_bF_buf3), .Y(datapath_1_Instr_17_bF_buf25_) );
BUFX2 BUFX2_253 ( .A(datapath_1_Instr_17__hier0_bF_buf3), .Y(datapath_1_Instr_17_bF_buf24_) );
BUFX2 BUFX2_254 ( .A(datapath_1_Instr_17__hier0_bF_buf3), .Y(datapath_1_Instr_17_bF_buf23_) );
BUFX2 BUFX2_255 ( .A(datapath_1_Instr_17__hier0_bF_buf6), .Y(datapath_1_Instr_17_bF_buf22_) );
BUFX2 BUFX2_256 ( .A(datapath_1_Instr_17__hier0_bF_buf2), .Y(datapath_1_Instr_17_bF_buf21_) );
BUFX2 BUFX2_257 ( .A(datapath_1_Instr_17__hier0_bF_buf2), .Y(datapath_1_Instr_17_bF_buf20_) );
BUFX2 BUFX2_258 ( .A(datapath_1_Instr_17__hier0_bF_buf0), .Y(datapath_1_Instr_17_bF_buf19_) );
BUFX2 BUFX2_259 ( .A(datapath_1_Instr_17__hier0_bF_buf6), .Y(datapath_1_Instr_17_bF_buf18_) );
BUFX2 BUFX2_260 ( .A(datapath_1_Instr_17__hier0_bF_buf0), .Y(datapath_1_Instr_17_bF_buf17_) );
BUFX2 BUFX2_261 ( .A(datapath_1_Instr_17__hier0_bF_buf2), .Y(datapath_1_Instr_17_bF_buf16_) );
BUFX2 BUFX2_262 ( .A(datapath_1_Instr_17__hier0_bF_buf0), .Y(datapath_1_Instr_17_bF_buf15_) );
BUFX2 BUFX2_263 ( .A(datapath_1_Instr_17__hier0_bF_buf0), .Y(datapath_1_Instr_17_bF_buf14_) );
BUFX2 BUFX2_264 ( .A(datapath_1_Instr_17__hier0_bF_buf2), .Y(datapath_1_Instr_17_bF_buf13_) );
BUFX2 BUFX2_265 ( .A(datapath_1_Instr_17__hier0_bF_buf0), .Y(datapath_1_Instr_17_bF_buf12_) );
BUFX2 BUFX2_266 ( .A(datapath_1_Instr_17__hier0_bF_buf2), .Y(datapath_1_Instr_17_bF_buf11_) );
BUFX2 BUFX2_267 ( .A(datapath_1_Instr_17__hier0_bF_buf2), .Y(datapath_1_Instr_17_bF_buf10_) );
BUFX2 BUFX2_268 ( .A(datapath_1_Instr_17__hier0_bF_buf0), .Y(datapath_1_Instr_17_bF_buf9_) );
BUFX2 BUFX2_269 ( .A(datapath_1_Instr_17__hier0_bF_buf0), .Y(datapath_1_Instr_17_bF_buf8_) );
BUFX2 BUFX2_270 ( .A(datapath_1_Instr_17__hier0_bF_buf4), .Y(datapath_1_Instr_17_bF_buf7_) );
BUFX2 BUFX2_271 ( .A(datapath_1_Instr_17__hier0_bF_buf6), .Y(datapath_1_Instr_17_bF_buf6_) );
BUFX2 BUFX2_272 ( .A(datapath_1_Instr_17__hier0_bF_buf2), .Y(datapath_1_Instr_17_bF_buf5_) );
BUFX2 BUFX2_273 ( .A(datapath_1_Instr_17__hier0_bF_buf3), .Y(datapath_1_Instr_17_bF_buf4_) );
BUFX2 BUFX2_274 ( .A(datapath_1_Instr_17__hier0_bF_buf6), .Y(datapath_1_Instr_17_bF_buf3_) );
BUFX2 BUFX2_275 ( .A(datapath_1_Instr_17__hier0_bF_buf6), .Y(datapath_1_Instr_17_bF_buf2_) );
BUFX2 BUFX2_276 ( .A(datapath_1_Instr_17__hier0_bF_buf1), .Y(datapath_1_Instr_17_bF_buf1_) );
BUFX2 BUFX2_277 ( .A(datapath_1_Instr_17__hier0_bF_buf6), .Y(datapath_1_Instr_17_bF_buf0_) );
BUFX2 BUFX2_278 ( .A(_5613_), .Y(_5613__bF_buf7) );
BUFX2 BUFX2_279 ( .A(_5613_), .Y(_5613__bF_buf6) );
BUFX2 BUFX2_280 ( .A(_5613_), .Y(_5613__bF_buf5) );
BUFX2 BUFX2_281 ( .A(_5613_), .Y(_5613__bF_buf4) );
BUFX2 BUFX2_282 ( .A(_5613_), .Y(_5613__bF_buf3) );
BUFX2 BUFX2_283 ( .A(_5613_), .Y(_5613__bF_buf2) );
BUFX2 BUFX2_284 ( .A(_5613_), .Y(_5613__bF_buf1) );
BUFX2 BUFX2_285 ( .A(_5613_), .Y(_5613__bF_buf0) );
BUFX2 BUFX2_286 ( .A(_5880_), .Y(_5880__bF_buf7) );
BUFX2 BUFX2_287 ( .A(_5880_), .Y(_5880__bF_buf6) );
BUFX2 BUFX2_288 ( .A(_5880_), .Y(_5880__bF_buf5) );
BUFX2 BUFX2_289 ( .A(_5880_), .Y(_5880__bF_buf4) );
BUFX2 BUFX2_290 ( .A(_5880_), .Y(_5880__bF_buf3) );
BUFX2 BUFX2_291 ( .A(_5880_), .Y(_5880__bF_buf2) );
BUFX2 BUFX2_292 ( .A(_5880_), .Y(_5880__bF_buf1) );
BUFX2 BUFX2_293 ( .A(_5880_), .Y(_5880__bF_buf0) );
BUFX2 BUFX2_294 ( .A(_6283_), .Y(_6283__bF_buf7) );
BUFX2 BUFX2_295 ( .A(_6283_), .Y(_6283__bF_buf6) );
BUFX2 BUFX2_296 ( .A(_6283_), .Y(_6283__bF_buf5) );
BUFX2 BUFX2_297 ( .A(_6283_), .Y(_6283__bF_buf4) );
BUFX2 BUFX2_298 ( .A(_6283_), .Y(_6283__bF_buf3) );
BUFX2 BUFX2_299 ( .A(_6283_), .Y(_6283__bF_buf2) );
BUFX2 BUFX2_300 ( .A(_6283_), .Y(_6283__bF_buf1) );
BUFX2 BUFX2_301 ( .A(_6283_), .Y(_6283__bF_buf0) );
BUFX2 BUFX2_302 ( .A(_6013_), .Y(_6013__bF_buf7) );
BUFX2 BUFX2_303 ( .A(_6013_), .Y(_6013__bF_buf6) );
BUFX2 BUFX2_304 ( .A(_6013_), .Y(_6013__bF_buf5) );
BUFX2 BUFX2_305 ( .A(_6013_), .Y(_6013__bF_buf4) );
BUFX2 BUFX2_306 ( .A(_6013_), .Y(_6013__bF_buf3) );
BUFX2 BUFX2_307 ( .A(_6013_), .Y(_6013__bF_buf2) );
BUFX2 BUFX2_308 ( .A(_6013_), .Y(_6013__bF_buf1) );
BUFX2 BUFX2_309 ( .A(_6013_), .Y(_6013__bF_buf0) );
BUFX2 BUFX2_310 ( .A(_5322_), .Y(_5322__bF_buf4) );
BUFX2 BUFX2_311 ( .A(_5322_), .Y(_5322__bF_buf3) );
BUFX2 BUFX2_312 ( .A(_5322_), .Y(_5322__bF_buf2) );
BUFX2 BUFX2_313 ( .A(_5322_), .Y(_5322__bF_buf1) );
BUFX2 BUFX2_314 ( .A(_5322_), .Y(_5322__bF_buf0) );
BUFX2 BUFX2_315 ( .A(_1888_), .Y(_1888__bF_buf7) );
BUFX2 BUFX2_316 ( .A(_1888_), .Y(_1888__bF_buf6) );
BUFX2 BUFX2_317 ( .A(_1888_), .Y(_1888__bF_buf5) );
BUFX2 BUFX2_318 ( .A(_1888_), .Y(_1888__bF_buf4) );
BUFX2 BUFX2_319 ( .A(_1888_), .Y(_1888__bF_buf3) );
BUFX2 BUFX2_320 ( .A(_1888_), .Y(_1888__bF_buf2) );
BUFX2 BUFX2_321 ( .A(_1888_), .Y(_1888__bF_buf1) );
BUFX2 BUFX2_322 ( .A(_1888_), .Y(_1888__bF_buf0) );
BUFX2 BUFX2_323 ( .A(_5298_), .Y(_5298__bF_buf4) );
BUFX2 BUFX2_324 ( .A(_5298_), .Y(_5298__bF_buf3) );
BUFX2 BUFX2_325 ( .A(_5298_), .Y(_5298__bF_buf2) );
BUFX2 BUFX2_326 ( .A(_5298_), .Y(_5298__bF_buf1) );
BUFX2 BUFX2_327 ( .A(_5298_), .Y(_5298__bF_buf0) );
BUFX2 BUFX2_328 ( .A(IorD), .Y(IorD_bF_buf7) );
BUFX2 BUFX2_329 ( .A(IorD), .Y(IorD_bF_buf6) );
BUFX2 BUFX2_330 ( .A(IorD), .Y(IorD_bF_buf5) );
BUFX2 BUFX2_331 ( .A(IorD), .Y(IorD_bF_buf4) );
BUFX2 BUFX2_332 ( .A(IorD), .Y(IorD_bF_buf3) );
BUFX2 BUFX2_333 ( .A(IorD), .Y(IorD_bF_buf2) );
BUFX2 BUFX2_334 ( .A(IorD), .Y(IorD_bF_buf1) );
BUFX2 BUFX2_335 ( .A(IorD), .Y(IorD_bF_buf0) );
CLKBUF1 CLKBUF1_1 ( .A(clk_hier0_bF_buf7), .Y(clk_bF_buf113) );
CLKBUF1 CLKBUF1_2 ( .A(clk_hier0_bF_buf2), .Y(clk_bF_buf112) );
CLKBUF1 CLKBUF1_3 ( .A(clk_hier0_bF_buf1), .Y(clk_bF_buf111) );
CLKBUF1 CLKBUF1_4 ( .A(clk_hier0_bF_buf5), .Y(clk_bF_buf110) );
CLKBUF1 CLKBUF1_5 ( .A(clk_hier0_bF_buf2), .Y(clk_bF_buf109) );
CLKBUF1 CLKBUF1_6 ( .A(clk_hier0_bF_buf4), .Y(clk_bF_buf108) );
CLKBUF1 CLKBUF1_7 ( .A(clk_hier0_bF_buf1), .Y(clk_bF_buf107) );
CLKBUF1 CLKBUF1_8 ( .A(clk_hier0_bF_buf7), .Y(clk_bF_buf106) );
CLKBUF1 CLKBUF1_9 ( .A(clk_hier0_bF_buf6), .Y(clk_bF_buf105) );
CLKBUF1 CLKBUF1_10 ( .A(clk_hier0_bF_buf3), .Y(clk_bF_buf104) );
CLKBUF1 CLKBUF1_11 ( .A(clk_hier0_bF_buf7), .Y(clk_bF_buf103) );
CLKBUF1 CLKBUF1_12 ( .A(clk_hier0_bF_buf2), .Y(clk_bF_buf102) );
CLKBUF1 CLKBUF1_13 ( .A(clk_hier0_bF_buf8), .Y(clk_bF_buf101) );
CLKBUF1 CLKBUF1_14 ( .A(clk_hier0_bF_buf9), .Y(clk_bF_buf100) );
CLKBUF1 CLKBUF1_15 ( .A(clk_hier0_bF_buf5), .Y(clk_bF_buf99) );
CLKBUF1 CLKBUF1_16 ( .A(clk_hier0_bF_buf8), .Y(clk_bF_buf98) );
CLKBUF1 CLKBUF1_17 ( .A(clk_hier0_bF_buf3), .Y(clk_bF_buf97) );
CLKBUF1 CLKBUF1_18 ( .A(clk_hier0_bF_buf7), .Y(clk_bF_buf96) );
CLKBUF1 CLKBUF1_19 ( .A(clk_hier0_bF_buf3), .Y(clk_bF_buf95) );
CLKBUF1 CLKBUF1_20 ( .A(clk_hier0_bF_buf1), .Y(clk_bF_buf94) );
CLKBUF1 CLKBUF1_21 ( .A(clk_hier0_bF_buf5), .Y(clk_bF_buf93) );
CLKBUF1 CLKBUF1_22 ( .A(clk_hier0_bF_buf1), .Y(clk_bF_buf92) );
CLKBUF1 CLKBUF1_23 ( .A(clk_hier0_bF_buf4), .Y(clk_bF_buf91) );
CLKBUF1 CLKBUF1_24 ( .A(clk_hier0_bF_buf9), .Y(clk_bF_buf90) );
CLKBUF1 CLKBUF1_25 ( .A(clk_hier0_bF_buf8), .Y(clk_bF_buf89) );
CLKBUF1 CLKBUF1_26 ( .A(clk_hier0_bF_buf4), .Y(clk_bF_buf88) );
CLKBUF1 CLKBUF1_27 ( .A(clk_hier0_bF_buf9), .Y(clk_bF_buf87) );
CLKBUF1 CLKBUF1_28 ( .A(clk_hier0_bF_buf9), .Y(clk_bF_buf86) );
CLKBUF1 CLKBUF1_29 ( .A(clk_hier0_bF_buf0), .Y(clk_bF_buf85) );
CLKBUF1 CLKBUF1_30 ( .A(clk_hier0_bF_buf5), .Y(clk_bF_buf84) );
CLKBUF1 CLKBUF1_31 ( .A(clk_hier0_bF_buf3), .Y(clk_bF_buf83) );
CLKBUF1 CLKBUF1_32 ( .A(clk_hier0_bF_buf7), .Y(clk_bF_buf82) );
CLKBUF1 CLKBUF1_33 ( .A(clk_hier0_bF_buf5), .Y(clk_bF_buf81) );
CLKBUF1 CLKBUF1_34 ( .A(clk_hier0_bF_buf6), .Y(clk_bF_buf80) );
CLKBUF1 CLKBUF1_35 ( .A(clk_hier0_bF_buf9), .Y(clk_bF_buf79) );
CLKBUF1 CLKBUF1_36 ( .A(clk_hier0_bF_buf3), .Y(clk_bF_buf78) );
CLKBUF1 CLKBUF1_37 ( .A(clk_hier0_bF_buf7), .Y(clk_bF_buf77) );
CLKBUF1 CLKBUF1_38 ( .A(clk_hier0_bF_buf4), .Y(clk_bF_buf76) );
CLKBUF1 CLKBUF1_39 ( .A(clk_hier0_bF_buf0), .Y(clk_bF_buf75) );
CLKBUF1 CLKBUF1_40 ( .A(clk_hier0_bF_buf1), .Y(clk_bF_buf74) );
CLKBUF1 CLKBUF1_41 ( .A(clk_hier0_bF_buf8), .Y(clk_bF_buf73) );
CLKBUF1 CLKBUF1_42 ( .A(clk_hier0_bF_buf2), .Y(clk_bF_buf72) );
CLKBUF1 CLKBUF1_43 ( .A(clk_hier0_bF_buf4), .Y(clk_bF_buf71) );
CLKBUF1 CLKBUF1_44 ( .A(clk_hier0_bF_buf8), .Y(clk_bF_buf70) );
CLKBUF1 CLKBUF1_45 ( .A(clk_hier0_bF_buf6), .Y(clk_bF_buf69) );
CLKBUF1 CLKBUF1_46 ( .A(clk_hier0_bF_buf6), .Y(clk_bF_buf68) );
CLKBUF1 CLKBUF1_47 ( .A(clk_hier0_bF_buf7), .Y(clk_bF_buf67) );
CLKBUF1 CLKBUF1_48 ( .A(clk_hier0_bF_buf4), .Y(clk_bF_buf66) );
CLKBUF1 CLKBUF1_49 ( .A(clk_hier0_bF_buf7), .Y(clk_bF_buf65) );
CLKBUF1 CLKBUF1_50 ( .A(clk_hier0_bF_buf8), .Y(clk_bF_buf64) );
CLKBUF1 CLKBUF1_51 ( .A(clk_hier0_bF_buf0), .Y(clk_bF_buf63) );
CLKBUF1 CLKBUF1_52 ( .A(clk_hier0_bF_buf5), .Y(clk_bF_buf62) );
CLKBUF1 CLKBUF1_53 ( .A(clk_hier0_bF_buf8), .Y(clk_bF_buf61) );
CLKBUF1 CLKBUF1_54 ( .A(clk_hier0_bF_buf4), .Y(clk_bF_buf60) );
CLKBUF1 CLKBUF1_55 ( .A(clk_hier0_bF_buf3), .Y(clk_bF_buf59) );
CLKBUF1 CLKBUF1_56 ( .A(clk_hier0_bF_buf3), .Y(clk_bF_buf58) );
CLKBUF1 CLKBUF1_57 ( .A(clk_hier0_bF_buf3), .Y(clk_bF_buf57) );
CLKBUF1 CLKBUF1_58 ( .A(clk_hier0_bF_buf9), .Y(clk_bF_buf56) );
CLKBUF1 CLKBUF1_59 ( .A(clk_hier0_bF_buf8), .Y(clk_bF_buf55) );
CLKBUF1 CLKBUF1_60 ( .A(clk_hier0_bF_buf8), .Y(clk_bF_buf54) );
CLKBUF1 CLKBUF1_61 ( .A(clk_hier0_bF_buf1), .Y(clk_bF_buf53) );
CLKBUF1 CLKBUF1_62 ( .A(clk_hier0_bF_buf3), .Y(clk_bF_buf52) );
CLKBUF1 CLKBUF1_63 ( .A(clk_hier0_bF_buf7), .Y(clk_bF_buf51) );
CLKBUF1 CLKBUF1_64 ( .A(clk_hier0_bF_buf4), .Y(clk_bF_buf50) );
CLKBUF1 CLKBUF1_65 ( .A(clk_hier0_bF_buf8), .Y(clk_bF_buf49) );
CLKBUF1 CLKBUF1_66 ( .A(clk_hier0_bF_buf9), .Y(clk_bF_buf48) );
CLKBUF1 CLKBUF1_67 ( .A(clk_hier0_bF_buf4), .Y(clk_bF_buf47) );
CLKBUF1 CLKBUF1_68 ( .A(clk_hier0_bF_buf2), .Y(clk_bF_buf46) );
CLKBUF1 CLKBUF1_69 ( .A(clk_hier0_bF_buf2), .Y(clk_bF_buf45) );
CLKBUF1 CLKBUF1_70 ( .A(clk_hier0_bF_buf6), .Y(clk_bF_buf44) );
CLKBUF1 CLKBUF1_71 ( .A(clk_hier0_bF_buf4), .Y(clk_bF_buf43) );
CLKBUF1 CLKBUF1_72 ( .A(clk_hier0_bF_buf0), .Y(clk_bF_buf42) );
CLKBUF1 CLKBUF1_73 ( .A(clk_hier0_bF_buf0), .Y(clk_bF_buf41) );
CLKBUF1 CLKBUF1_74 ( .A(clk_hier0_bF_buf0), .Y(clk_bF_buf40) );
CLKBUF1 CLKBUF1_75 ( .A(clk_hier0_bF_buf5), .Y(clk_bF_buf39) );
CLKBUF1 CLKBUF1_76 ( .A(clk_hier0_bF_buf0), .Y(clk_bF_buf38) );
CLKBUF1 CLKBUF1_77 ( .A(clk_hier0_bF_buf1), .Y(clk_bF_buf37) );
CLKBUF1 CLKBUF1_78 ( .A(clk_hier0_bF_buf2), .Y(clk_bF_buf36) );
CLKBUF1 CLKBUF1_79 ( .A(clk_hier0_bF_buf8), .Y(clk_bF_buf35) );
CLKBUF1 CLKBUF1_80 ( .A(clk_hier0_bF_buf9), .Y(clk_bF_buf34) );
CLKBUF1 CLKBUF1_81 ( .A(clk_hier0_bF_buf5), .Y(clk_bF_buf33) );
CLKBUF1 CLKBUF1_82 ( .A(clk_hier0_bF_buf8), .Y(clk_bF_buf32) );
CLKBUF1 CLKBUF1_83 ( .A(clk_hier0_bF_buf3), .Y(clk_bF_buf31) );
CLKBUF1 CLKBUF1_84 ( .A(clk_hier0_bF_buf1), .Y(clk_bF_buf30) );
CLKBUF1 CLKBUF1_85 ( .A(clk_hier0_bF_buf9), .Y(clk_bF_buf29) );
CLKBUF1 CLKBUF1_86 ( .A(clk_hier0_bF_buf5), .Y(clk_bF_buf28) );
CLKBUF1 CLKBUF1_87 ( .A(clk_hier0_bF_buf6), .Y(clk_bF_buf27) );
CLKBUF1 CLKBUF1_88 ( .A(clk_hier0_bF_buf4), .Y(clk_bF_buf26) );
CLKBUF1 CLKBUF1_89 ( .A(clk_hier0_bF_buf0), .Y(clk_bF_buf25) );
CLKBUF1 CLKBUF1_90 ( .A(clk_hier0_bF_buf6), .Y(clk_bF_buf24) );
CLKBUF1 CLKBUF1_91 ( .A(clk_hier0_bF_buf9), .Y(clk_bF_buf23) );
CLKBUF1 CLKBUF1_92 ( .A(clk_hier0_bF_buf9), .Y(clk_bF_buf22) );
CLKBUF1 CLKBUF1_93 ( .A(clk_hier0_bF_buf7), .Y(clk_bF_buf21) );
CLKBUF1 CLKBUF1_94 ( .A(clk_hier0_bF_buf2), .Y(clk_bF_buf20) );
CLKBUF1 CLKBUF1_95 ( .A(clk_hier0_bF_buf1), .Y(clk_bF_buf19) );
CLKBUF1 CLKBUF1_96 ( .A(clk_hier0_bF_buf6), .Y(clk_bF_buf18) );
CLKBUF1 CLKBUF1_97 ( .A(clk_hier0_bF_buf5), .Y(clk_bF_buf17) );
CLKBUF1 CLKBUF1_98 ( .A(clk_hier0_bF_buf2), .Y(clk_bF_buf16) );
CLKBUF1 CLKBUF1_99 ( .A(clk_hier0_bF_buf1), .Y(clk_bF_buf15) );
CLKBUF1 CLKBUF1_100 ( .A(clk_hier0_bF_buf0), .Y(clk_bF_buf14) );
CLKBUF1 CLKBUF1_101 ( .A(clk_hier0_bF_buf9), .Y(clk_bF_buf13) );
CLKBUF1 CLKBUF1_102 ( .A(clk_hier0_bF_buf5), .Y(clk_bF_buf12) );
CLKBUF1 CLKBUF1_103 ( .A(clk_hier0_bF_buf2), .Y(clk_bF_buf11) );
CLKBUF1 CLKBUF1_104 ( .A(clk_hier0_bF_buf3), .Y(clk_bF_buf10) );
CLKBUF1 CLKBUF1_105 ( .A(clk_hier0_bF_buf6), .Y(clk_bF_buf9) );
CLKBUF1 CLKBUF1_106 ( .A(clk_hier0_bF_buf6), .Y(clk_bF_buf8) );
CLKBUF1 CLKBUF1_107 ( .A(clk_hier0_bF_buf2), .Y(clk_bF_buf7) );
CLKBUF1 CLKBUF1_108 ( .A(clk_hier0_bF_buf0), .Y(clk_bF_buf6) );
CLKBUF1 CLKBUF1_109 ( .A(clk_hier0_bF_buf1), .Y(clk_bF_buf5) );
CLKBUF1 CLKBUF1_110 ( .A(clk_hier0_bF_buf6), .Y(clk_bF_buf4) );
CLKBUF1 CLKBUF1_111 ( .A(clk_hier0_bF_buf0), .Y(clk_bF_buf3) );
CLKBUF1 CLKBUF1_112 ( .A(clk_hier0_bF_buf7), .Y(clk_bF_buf2) );
CLKBUF1 CLKBUF1_113 ( .A(clk_hier0_bF_buf7), .Y(clk_bF_buf1) );
CLKBUF1 CLKBUF1_114 ( .A(clk_hier0_bF_buf6), .Y(clk_bF_buf0) );
BUFX2 BUFX2_336 ( .A(_5316_), .Y(_5316__bF_buf4) );
BUFX2 BUFX2_337 ( .A(_5316_), .Y(_5316__bF_buf3) );
BUFX2 BUFX2_338 ( .A(_5316_), .Y(_5316__bF_buf2) );
BUFX2 BUFX2_339 ( .A(_5316_), .Y(_5316__bF_buf1) );
BUFX2 BUFX2_340 ( .A(_5316_), .Y(_5316__bF_buf0) );
BUFX2 BUFX2_341 ( .A(_5545_), .Y(_5545__bF_buf7) );
BUFX2 BUFX2_342 ( .A(_5545_), .Y(_5545__bF_buf6) );
BUFX2 BUFX2_343 ( .A(_5545_), .Y(_5545__bF_buf5) );
BUFX2 BUFX2_344 ( .A(_5545_), .Y(_5545__bF_buf4) );
BUFX2 BUFX2_345 ( .A(_5545_), .Y(_5545__bF_buf3) );
BUFX2 BUFX2_346 ( .A(_5545_), .Y(_5545__bF_buf2) );
BUFX2 BUFX2_347 ( .A(_5545_), .Y(_5545__bF_buf1) );
BUFX2 BUFX2_348 ( .A(_5545_), .Y(_5545__bF_buf0) );
BUFX2 BUFX2_349 ( .A(_1885_), .Y(_1885__bF_buf11) );
BUFX2 BUFX2_350 ( .A(_1885_), .Y(_1885__bF_buf10) );
BUFX2 BUFX2_351 ( .A(_1885_), .Y(_1885__bF_buf9) );
BUFX2 BUFX2_352 ( .A(_1885_), .Y(_1885__bF_buf8) );
BUFX2 BUFX2_353 ( .A(_1885_), .Y(_1885__bF_buf7) );
BUFX2 BUFX2_354 ( .A(_1885_), .Y(_1885__bF_buf6) );
BUFX2 BUFX2_355 ( .A(_1885_), .Y(_1885__bF_buf5) );
BUFX2 BUFX2_356 ( .A(_1885_), .Y(_1885__bF_buf4) );
BUFX2 BUFX2_357 ( .A(_1885_), .Y(_1885__bF_buf3) );
BUFX2 BUFX2_358 ( .A(_1885_), .Y(_1885__bF_buf2) );
BUFX2 BUFX2_359 ( .A(_1885_), .Y(_1885__bF_buf1) );
BUFX2 BUFX2_360 ( .A(_1885_), .Y(_1885__bF_buf0) );
BUFX2 BUFX2_361 ( .A(datapath_1_PCEn), .Y(datapath_1_PCEn_bF_buf4) );
BUFX2 BUFX2_362 ( .A(datapath_1_PCEn), .Y(datapath_1_PCEn_bF_buf3) );
BUFX2 BUFX2_363 ( .A(datapath_1_PCEn), .Y(datapath_1_PCEn_bF_buf2) );
BUFX2 BUFX2_364 ( .A(datapath_1_PCEn), .Y(datapath_1_PCEn_bF_buf1) );
BUFX2 BUFX2_365 ( .A(datapath_1_PCEn), .Y(datapath_1_PCEn_bF_buf0) );
BUFX2 BUFX2_366 ( .A(_5580_), .Y(_5580__bF_buf7) );
BUFX2 BUFX2_367 ( .A(_5580_), .Y(_5580__bF_buf6) );
BUFX2 BUFX2_368 ( .A(_5580_), .Y(_5580__bF_buf5) );
BUFX2 BUFX2_369 ( .A(_5580_), .Y(_5580__bF_buf4) );
BUFX2 BUFX2_370 ( .A(_5580_), .Y(_5580__bF_buf3) );
BUFX2 BUFX2_371 ( .A(_5580_), .Y(_5580__bF_buf2) );
BUFX2 BUFX2_372 ( .A(_5580_), .Y(_5580__bF_buf1) );
BUFX2 BUFX2_373 ( .A(_5580_), .Y(_5580__bF_buf0) );
BUFX2 BUFX2_374 ( .A(_5292_), .Y(_5292__bF_buf4) );
BUFX2 BUFX2_375 ( .A(_5292_), .Y(_5292__bF_buf3) );
BUFX2 BUFX2_376 ( .A(_5292_), .Y(_5292__bF_buf2) );
BUFX2 BUFX2_377 ( .A(_5292_), .Y(_5292__bF_buf1) );
BUFX2 BUFX2_378 ( .A(_5292_), .Y(_5292__bF_buf0) );
BUFX2 BUFX2_379 ( .A(_5310_), .Y(_5310__bF_buf4) );
BUFX2 BUFX2_380 ( .A(_5310_), .Y(_5310__bF_buf3) );
BUFX2 BUFX2_381 ( .A(_5310_), .Y(_5310__bF_buf2) );
BUFX2 BUFX2_382 ( .A(_5310_), .Y(_5310__bF_buf1) );
BUFX2 BUFX2_383 ( .A(_5310_), .Y(_5310__bF_buf0) );
BUFX2 BUFX2_384 ( .A(_5286_), .Y(_5286__bF_buf4) );
BUFX2 BUFX2_385 ( .A(_5286_), .Y(_5286__bF_buf3) );
BUFX2 BUFX2_386 ( .A(_5286_), .Y(_5286__bF_buf2) );
BUFX2 BUFX2_387 ( .A(_5286_), .Y(_5286__bF_buf1) );
BUFX2 BUFX2_388 ( .A(_5286_), .Y(_5286__bF_buf0) );
BUFX2 BUFX2_389 ( .A(_7050_), .Y(_7050__bF_buf4) );
BUFX2 BUFX2_390 ( .A(_7050_), .Y(_7050__bF_buf3) );
BUFX2 BUFX2_391 ( .A(_7050_), .Y(_7050__bF_buf2) );
BUFX2 BUFX2_392 ( .A(_7050_), .Y(_7050__bF_buf1) );
BUFX2 BUFX2_393 ( .A(_7050_), .Y(_7050__bF_buf0) );
BUFX2 BUFX2_394 ( .A(ALUSrcB_0_), .Y(ALUSrcB_0_bF_buf4_) );
BUFX2 BUFX2_395 ( .A(ALUSrcB_0_), .Y(ALUSrcB_0_bF_buf3_) );
BUFX2 BUFX2_396 ( .A(ALUSrcB_0_), .Y(ALUSrcB_0_bF_buf2_) );
BUFX2 BUFX2_397 ( .A(ALUSrcB_0_), .Y(ALUSrcB_0_bF_buf1_) );
BUFX2 BUFX2_398 ( .A(ALUSrcB_0_), .Y(ALUSrcB_0_bF_buf0_) );
BUFX2 BUFX2_399 ( .A(_5304_), .Y(_5304__bF_buf4) );
BUFX2 BUFX2_400 ( .A(_5304_), .Y(_5304__bF_buf3) );
BUFX2 BUFX2_401 ( .A(_5304_), .Y(_5304__bF_buf2) );
BUFX2 BUFX2_402 ( .A(_5304_), .Y(_5304__bF_buf1) );
BUFX2 BUFX2_403 ( .A(_5304_), .Y(_5304__bF_buf0) );
BUFX2 BUFX2_404 ( .A(_5342_), .Y(_5342__bF_buf7) );
BUFX2 BUFX2_405 ( .A(_5342_), .Y(_5342__bF_buf6) );
BUFX2 BUFX2_406 ( .A(_5342_), .Y(_5342__bF_buf5) );
BUFX2 BUFX2_407 ( .A(_5342_), .Y(_5342__bF_buf4) );
BUFX2 BUFX2_408 ( .A(_5342_), .Y(_5342__bF_buf3) );
BUFX2 BUFX2_409 ( .A(_5342_), .Y(_5342__bF_buf2) );
BUFX2 BUFX2_410 ( .A(_5342_), .Y(_5342__bF_buf1) );
BUFX2 BUFX2_411 ( .A(_5342_), .Y(_5342__bF_buf0) );
BUFX2 BUFX2_412 ( .A(_6547_), .Y(_6547__bF_buf4) );
BUFX2 BUFX2_413 ( .A(_6547_), .Y(_6547__bF_buf3) );
BUFX2 BUFX2_414 ( .A(_6547_), .Y(_6547__bF_buf2) );
BUFX2 BUFX2_415 ( .A(_6547_), .Y(_6547__bF_buf1) );
BUFX2 BUFX2_416 ( .A(_6547_), .Y(_6547__bF_buf0) );
BUFX2 BUFX2_417 ( .A(_5377_), .Y(_5377__bF_buf7) );
BUFX2 BUFX2_418 ( .A(_5377_), .Y(_5377__bF_buf6) );
BUFX2 BUFX2_419 ( .A(_5377_), .Y(_5377__bF_buf5) );
BUFX2 BUFX2_420 ( .A(_5377_), .Y(_5377__bF_buf4) );
BUFX2 BUFX2_421 ( .A(_5377_), .Y(_5377__bF_buf3) );
BUFX2 BUFX2_422 ( .A(_5377_), .Y(_5377__bF_buf2) );
BUFX2 BUFX2_423 ( .A(_5377_), .Y(_5377__bF_buf1) );
BUFX2 BUFX2_424 ( .A(_5377_), .Y(_5377__bF_buf0) );
BUFX2 BUFX2_425 ( .A(_5280_), .Y(_5280__bF_buf4) );
BUFX2 BUFX2_426 ( .A(_5280_), .Y(_5280__bF_buf3) );
BUFX2 BUFX2_427 ( .A(_5280_), .Y(_5280__bF_buf2) );
BUFX2 BUFX2_428 ( .A(_5280_), .Y(_5280__bF_buf1) );
BUFX2 BUFX2_429 ( .A(_5280_), .Y(_5280__bF_buf0) );
BUFX2 BUFX2_430 ( .A(_5336_), .Y(_5336__bF_buf4) );
BUFX2 BUFX2_431 ( .A(_5336_), .Y(_5336__bF_buf3) );
BUFX2 BUFX2_432 ( .A(_5336_), .Y(_5336__bF_buf2) );
BUFX2 BUFX2_433 ( .A(_5336_), .Y(_5336__bF_buf1) );
BUFX2 BUFX2_434 ( .A(_5336_), .Y(_5336__bF_buf0) );
BUFX2 BUFX2_435 ( .A(_6388_), .Y(_6388__bF_buf4) );
BUFX2 BUFX2_436 ( .A(_6388_), .Y(_6388__bF_buf3) );
BUFX2 BUFX2_437 ( .A(_6388_), .Y(_6388__bF_buf2) );
BUFX2 BUFX2_438 ( .A(_6388_), .Y(_6388__bF_buf1) );
BUFX2 BUFX2_439 ( .A(_6388_), .Y(_6388__bF_buf0) );
BUFX2 BUFX2_440 ( .A(datapath_1_Instr_25_), .Y(datapath_1_Instr_25_bF_buf5_) );
BUFX2 BUFX2_441 ( .A(datapath_1_Instr_25_), .Y(datapath_1_Instr_25_bF_buf4_) );
BUFX2 BUFX2_442 ( .A(datapath_1_Instr_25_), .Y(datapath_1_Instr_25_bF_buf3_) );
BUFX2 BUFX2_443 ( .A(datapath_1_Instr_25_), .Y(datapath_1_Instr_25_bF_buf2_) );
BUFX2 BUFX2_444 ( .A(datapath_1_Instr_25_), .Y(datapath_1_Instr_25_bF_buf1_) );
BUFX2 BUFX2_445 ( .A(datapath_1_Instr_25_), .Y(datapath_1_Instr_25_bF_buf0_) );
BUFX2 BUFX2_446 ( .A(_5812_), .Y(_5812__bF_buf7) );
BUFX2 BUFX2_447 ( .A(_5812_), .Y(_5812__bF_buf6) );
BUFX2 BUFX2_448 ( .A(_5812_), .Y(_5812__bF_buf5) );
BUFX2 BUFX2_449 ( .A(_5812_), .Y(_5812__bF_buf4) );
BUFX2 BUFX2_450 ( .A(_5812_), .Y(_5812__bF_buf3) );
BUFX2 BUFX2_451 ( .A(_5812_), .Y(_5812__bF_buf2) );
BUFX2 BUFX2_452 ( .A(_5812_), .Y(_5812__bF_buf1) );
BUFX2 BUFX2_453 ( .A(_5812_), .Y(_5812__bF_buf0) );
BUFX2 BUFX2_454 ( .A(_6350_), .Y(_6350__bF_buf7) );
BUFX2 BUFX2_455 ( .A(_6350_), .Y(_6350__bF_buf6) );
BUFX2 BUFX2_456 ( .A(_6350_), .Y(_6350__bF_buf5) );
BUFX2 BUFX2_457 ( .A(_6350_), .Y(_6350__bF_buf4) );
BUFX2 BUFX2_458 ( .A(_6350_), .Y(_6350__bF_buf3) );
BUFX2 BUFX2_459 ( .A(_6350_), .Y(_6350__bF_buf2) );
BUFX2 BUFX2_460 ( .A(_6350_), .Y(_6350__bF_buf1) );
BUFX2 BUFX2_461 ( .A(_6350_), .Y(_6350__bF_buf0) );
BUFX2 BUFX2_462 ( .A(_6215_), .Y(_6215__bF_buf7) );
BUFX2 BUFX2_463 ( .A(_6215_), .Y(_6215__bF_buf6) );
BUFX2 BUFX2_464 ( .A(_6215_), .Y(_6215__bF_buf5) );
BUFX2 BUFX2_465 ( .A(_6215_), .Y(_6215__bF_buf4) );
BUFX2 BUFX2_466 ( .A(_6215_), .Y(_6215__bF_buf3) );
BUFX2 BUFX2_467 ( .A(_6215_), .Y(_6215__bF_buf2) );
BUFX2 BUFX2_468 ( .A(_6215_), .Y(_6215__bF_buf1) );
BUFX2 BUFX2_469 ( .A(_6215_), .Y(_6215__bF_buf0) );
BUFX2 BUFX2_470 ( .A(_3569_), .Y(_3569__bF_buf4) );
BUFX2 BUFX2_471 ( .A(_3569_), .Y(_3569__bF_buf3) );
BUFX2 BUFX2_472 ( .A(_3569_), .Y(_3569__bF_buf2) );
BUFX2 BUFX2_473 ( .A(_3569_), .Y(_3569__bF_buf1) );
BUFX2 BUFX2_474 ( .A(_3569_), .Y(_3569__bF_buf0) );
BUFX2 BUFX2_475 ( .A(_5847_), .Y(_5847__bF_buf7) );
BUFX2 BUFX2_476 ( .A(_5847_), .Y(_5847__bF_buf6) );
BUFX2 BUFX2_477 ( .A(_5847_), .Y(_5847__bF_buf5) );
BUFX2 BUFX2_478 ( .A(_5847_), .Y(_5847__bF_buf4) );
BUFX2 BUFX2_479 ( .A(_5847_), .Y(_5847__bF_buf3) );
BUFX2 BUFX2_480 ( .A(_5847_), .Y(_5847__bF_buf2) );
BUFX2 BUFX2_481 ( .A(_5847_), .Y(_5847__bF_buf1) );
BUFX2 BUFX2_482 ( .A(_5847_), .Y(_5847__bF_buf0) );
BUFX2 BUFX2_483 ( .A(_6385_), .Y(_6385__bF_buf4) );
BUFX2 BUFX2_484 ( .A(_6385_), .Y(_6385__bF_buf3) );
BUFX2 BUFX2_485 ( .A(_6385_), .Y(_6385__bF_buf2) );
BUFX2 BUFX2_486 ( .A(_6385_), .Y(_6385__bF_buf1) );
BUFX2 BUFX2_487 ( .A(_6385_), .Y(_6385__bF_buf0) );
BUFX2 BUFX2_488 ( .A(datapath_1_Instr_22__hier0_bF_buf3), .Y(datapath_1_Instr_22_bF_buf50_) );
BUFX2 BUFX2_489 ( .A(datapath_1_Instr_22__hier0_bF_buf3), .Y(datapath_1_Instr_22_bF_buf49_) );
BUFX2 BUFX2_490 ( .A(datapath_1_Instr_22__hier0_bF_buf2), .Y(datapath_1_Instr_22_bF_buf48_) );
BUFX2 BUFX2_491 ( .A(datapath_1_Instr_22__hier0_bF_buf0), .Y(datapath_1_Instr_22_bF_buf47_) );
BUFX2 BUFX2_492 ( .A(datapath_1_Instr_22__hier0_bF_buf2), .Y(datapath_1_Instr_22_bF_buf46_) );
BUFX2 BUFX2_493 ( .A(datapath_1_Instr_22__hier0_bF_buf0), .Y(datapath_1_Instr_22_bF_buf45_) );
BUFX2 BUFX2_494 ( .A(datapath_1_Instr_22__hier0_bF_buf2), .Y(datapath_1_Instr_22_bF_buf44_) );
BUFX2 BUFX2_495 ( .A(datapath_1_Instr_22__hier0_bF_buf2), .Y(datapath_1_Instr_22_bF_buf43_) );
BUFX2 BUFX2_496 ( .A(datapath_1_Instr_22__hier0_bF_buf2), .Y(datapath_1_Instr_22_bF_buf42_) );
BUFX2 BUFX2_497 ( .A(datapath_1_Instr_22__hier0_bF_buf0), .Y(datapath_1_Instr_22_bF_buf41_) );
BUFX2 BUFX2_498 ( .A(datapath_1_Instr_22__hier0_bF_buf0), .Y(datapath_1_Instr_22_bF_buf40_) );
BUFX2 BUFX2_499 ( .A(datapath_1_Instr_22__hier0_bF_buf2), .Y(datapath_1_Instr_22_bF_buf39_) );
BUFX2 BUFX2_500 ( .A(datapath_1_Instr_22__hier0_bF_buf2), .Y(datapath_1_Instr_22_bF_buf38_) );
BUFX2 BUFX2_501 ( .A(datapath_1_Instr_22__hier0_bF_buf0), .Y(datapath_1_Instr_22_bF_buf37_) );
BUFX2 BUFX2_502 ( .A(datapath_1_Instr_22__hier0_bF_buf0), .Y(datapath_1_Instr_22_bF_buf36_) );
BUFX2 BUFX2_503 ( .A(datapath_1_Instr_22__hier0_bF_buf3), .Y(datapath_1_Instr_22_bF_buf35_) );
BUFX2 BUFX2_504 ( .A(datapath_1_Instr_22__hier0_bF_buf0), .Y(datapath_1_Instr_22_bF_buf34_) );
BUFX2 BUFX2_505 ( .A(datapath_1_Instr_22__hier0_bF_buf5), .Y(datapath_1_Instr_22_bF_buf33_) );
BUFX2 BUFX2_506 ( .A(datapath_1_Instr_22__hier0_bF_buf5), .Y(datapath_1_Instr_22_bF_buf32_) );
BUFX2 BUFX2_507 ( .A(datapath_1_Instr_22__hier0_bF_buf1), .Y(datapath_1_Instr_22_bF_buf31_) );
BUFX2 BUFX2_508 ( .A(datapath_1_Instr_22__hier0_bF_buf4), .Y(datapath_1_Instr_22_bF_buf30_) );
BUFX2 BUFX2_509 ( .A(datapath_1_Instr_22__hier0_bF_buf6), .Y(datapath_1_Instr_22_bF_buf29_) );
BUFX2 BUFX2_510 ( .A(datapath_1_Instr_22__hier0_bF_buf6), .Y(datapath_1_Instr_22_bF_buf28_) );
BUFX2 BUFX2_511 ( .A(datapath_1_Instr_22__hier0_bF_buf6), .Y(datapath_1_Instr_22_bF_buf27_) );
BUFX2 BUFX2_512 ( .A(datapath_1_Instr_22__hier0_bF_buf1), .Y(datapath_1_Instr_22_bF_buf26_) );
BUFX2 BUFX2_513 ( .A(datapath_1_Instr_22__hier0_bF_buf1), .Y(datapath_1_Instr_22_bF_buf25_) );
BUFX2 BUFX2_514 ( .A(datapath_1_Instr_22__hier0_bF_buf6), .Y(datapath_1_Instr_22_bF_buf24_) );
BUFX2 BUFX2_515 ( .A(datapath_1_Instr_22__hier0_bF_buf4), .Y(datapath_1_Instr_22_bF_buf23_) );
BUFX2 BUFX2_516 ( .A(datapath_1_Instr_22__hier0_bF_buf1), .Y(datapath_1_Instr_22_bF_buf22_) );
BUFX2 BUFX2_517 ( .A(datapath_1_Instr_22__hier0_bF_buf1), .Y(datapath_1_Instr_22_bF_buf21_) );
BUFX2 BUFX2_518 ( .A(datapath_1_Instr_22__hier0_bF_buf4), .Y(datapath_1_Instr_22_bF_buf20_) );
BUFX2 BUFX2_519 ( .A(datapath_1_Instr_22__hier0_bF_buf4), .Y(datapath_1_Instr_22_bF_buf19_) );
BUFX2 BUFX2_520 ( .A(datapath_1_Instr_22__hier0_bF_buf4), .Y(datapath_1_Instr_22_bF_buf18_) );
BUFX2 BUFX2_521 ( .A(datapath_1_Instr_22__hier0_bF_buf6), .Y(datapath_1_Instr_22_bF_buf17_) );
BUFX2 BUFX2_522 ( .A(datapath_1_Instr_22__hier0_bF_buf1), .Y(datapath_1_Instr_22_bF_buf16_) );
BUFX2 BUFX2_523 ( .A(datapath_1_Instr_22__hier0_bF_buf4), .Y(datapath_1_Instr_22_bF_buf15_) );
BUFX2 BUFX2_524 ( .A(datapath_1_Instr_22__hier0_bF_buf6), .Y(datapath_1_Instr_22_bF_buf14_) );
BUFX2 BUFX2_525 ( .A(datapath_1_Instr_22__hier0_bF_buf4), .Y(datapath_1_Instr_22_bF_buf13_) );
BUFX2 BUFX2_526 ( .A(datapath_1_Instr_22__hier0_bF_buf1), .Y(datapath_1_Instr_22_bF_buf12_) );
BUFX2 BUFX2_527 ( .A(datapath_1_Instr_22__hier0_bF_buf3), .Y(datapath_1_Instr_22_bF_buf11_) );
BUFX2 BUFX2_528 ( .A(datapath_1_Instr_22__hier0_bF_buf5), .Y(datapath_1_Instr_22_bF_buf10_) );
BUFX2 BUFX2_529 ( .A(datapath_1_Instr_22__hier0_bF_buf6), .Y(datapath_1_Instr_22_bF_buf9_) );
BUFX2 BUFX2_530 ( .A(datapath_1_Instr_22__hier0_bF_buf5), .Y(datapath_1_Instr_22_bF_buf8_) );
BUFX2 BUFX2_531 ( .A(datapath_1_Instr_22__hier0_bF_buf6), .Y(datapath_1_Instr_22_bF_buf7_) );
BUFX2 BUFX2_532 ( .A(datapath_1_Instr_22__hier0_bF_buf5), .Y(datapath_1_Instr_22_bF_buf6_) );
BUFX2 BUFX2_533 ( .A(datapath_1_Instr_22__hier0_bF_buf5), .Y(datapath_1_Instr_22_bF_buf5_) );
BUFX2 BUFX2_534 ( .A(datapath_1_Instr_22__hier0_bF_buf3), .Y(datapath_1_Instr_22_bF_buf4_) );
BUFX2 BUFX2_535 ( .A(datapath_1_Instr_22__hier0_bF_buf5), .Y(datapath_1_Instr_22_bF_buf3_) );
BUFX2 BUFX2_536 ( .A(datapath_1_Instr_22__hier0_bF_buf3), .Y(datapath_1_Instr_22_bF_buf2_) );
BUFX2 BUFX2_537 ( .A(datapath_1_Instr_22__hier0_bF_buf5), .Y(datapath_1_Instr_22_bF_buf1_) );
BUFX2 BUFX2_538 ( .A(datapath_1_Instr_22__hier0_bF_buf3), .Y(datapath_1_Instr_22_bF_buf0_) );
BUFX2 BUFX2_539 ( .A(_3566_), .Y(_3566__bF_buf10) );
BUFX2 BUFX2_540 ( .A(_3566_), .Y(_3566__bF_buf9) );
BUFX2 BUFX2_541 ( .A(_3566_), .Y(_3566__bF_buf8) );
BUFX2 BUFX2_542 ( .A(_3566_), .Y(_3566__bF_buf7) );
BUFX2 BUFX2_543 ( .A(_3566_), .Y(_3566__bF_buf6) );
BUFX2 BUFX2_544 ( .A(_3566_), .Y(_3566__bF_buf5) );
BUFX2 BUFX2_545 ( .A(_3566_), .Y(_3566__bF_buf4) );
BUFX2 BUFX2_546 ( .A(_3566_), .Y(_3566__bF_buf3) );
BUFX2 BUFX2_547 ( .A(_3566_), .Y(_3566__bF_buf2) );
BUFX2 BUFX2_548 ( .A(_3566_), .Y(_3566__bF_buf1) );
BUFX2 BUFX2_549 ( .A(_3566_), .Y(_3566__bF_buf0) );
BUFX2 BUFX2_550 ( .A(datapath_1_Instr_19_), .Y(datapath_1_Instr_19_bF_buf6_) );
BUFX2 BUFX2_551 ( .A(datapath_1_Instr_19_), .Y(datapath_1_Instr_19_bF_buf5_) );
BUFX2 BUFX2_552 ( .A(datapath_1_Instr_19_), .Y(datapath_1_Instr_19_bF_buf4_) );
BUFX2 BUFX2_553 ( .A(datapath_1_Instr_19_), .Y(datapath_1_Instr_19_bF_buf3_) );
BUFX2 BUFX2_554 ( .A(datapath_1_Instr_19_), .Y(datapath_1_Instr_19_bF_buf2_) );
BUFX2 BUFX2_555 ( .A(datapath_1_Instr_19_), .Y(datapath_1_Instr_19_bF_buf1_) );
BUFX2 BUFX2_556 ( .A(datapath_1_Instr_19_), .Y(datapath_1_Instr_19_bF_buf0_) );
BUFX2 BUFX2_557 ( .A(_6250_), .Y(_6250__bF_buf7) );
BUFX2 BUFX2_558 ( .A(_6250_), .Y(_6250__bF_buf6) );
BUFX2 BUFX2_559 ( .A(_6250_), .Y(_6250__bF_buf5) );
BUFX2 BUFX2_560 ( .A(_6250_), .Y(_6250__bF_buf4) );
BUFX2 BUFX2_561 ( .A(_6250_), .Y(_6250__bF_buf3) );
BUFX2 BUFX2_562 ( .A(_6250_), .Y(_6250__bF_buf2) );
BUFX2 BUFX2_563 ( .A(_6250_), .Y(_6250__bF_buf1) );
BUFX2 BUFX2_564 ( .A(_6250_), .Y(_6250__bF_buf0) );
BUFX2 BUFX2_565 ( .A(_1917_), .Y(_1917__bF_buf4) );
BUFX2 BUFX2_566 ( .A(_1917_), .Y(_1917__bF_buf3) );
BUFX2 BUFX2_567 ( .A(_1917_), .Y(_1917__bF_buf2) );
BUFX2 BUFX2_568 ( .A(_1917_), .Y(_1917__bF_buf1) );
BUFX2 BUFX2_569 ( .A(_1917_), .Y(_1917__bF_buf0) );
BUFX2 BUFX2_570 ( .A(_5330_), .Y(_5330__bF_buf4) );
BUFX2 BUFX2_571 ( .A(_5330_), .Y(_5330__bF_buf3) );
BUFX2 BUFX2_572 ( .A(_5330_), .Y(_5330__bF_buf2) );
BUFX2 BUFX2_573 ( .A(_5330_), .Y(_5330__bF_buf1) );
BUFX2 BUFX2_574 ( .A(_5330_), .Y(_5330__bF_buf0) );
BUFX2 BUFX2_575 ( .A(datapath_1_Instr_16__hier0_bF_buf5), .Y(datapath_1_Instr_16_bF_buf55_) );
BUFX2 BUFX2_576 ( .A(datapath_1_Instr_16__hier0_bF_buf6), .Y(datapath_1_Instr_16_bF_buf54_) );
BUFX2 BUFX2_577 ( .A(datapath_1_Instr_16__hier0_bF_buf2), .Y(datapath_1_Instr_16_bF_buf53_) );
BUFX2 BUFX2_578 ( .A(datapath_1_Instr_16__hier0_bF_buf5), .Y(datapath_1_Instr_16_bF_buf52_) );
BUFX2 BUFX2_579 ( .A(datapath_1_Instr_16__hier0_bF_buf0), .Y(datapath_1_Instr_16_bF_buf51_) );
BUFX2 BUFX2_580 ( .A(datapath_1_Instr_16__hier0_bF_buf1), .Y(datapath_1_Instr_16_bF_buf50_) );
BUFX2 BUFX2_581 ( .A(datapath_1_Instr_16__hier0_bF_buf4), .Y(datapath_1_Instr_16_bF_buf49_) );
BUFX2 BUFX2_582 ( .A(datapath_1_Instr_16__hier0_bF_buf3), .Y(datapath_1_Instr_16_bF_buf48_) );
BUFX2 BUFX2_583 ( .A(datapath_1_Instr_16__hier0_bF_buf4), .Y(datapath_1_Instr_16_bF_buf47_) );
BUFX2 BUFX2_584 ( .A(datapath_1_Instr_16__hier0_bF_buf3), .Y(datapath_1_Instr_16_bF_buf46_) );
BUFX2 BUFX2_585 ( .A(datapath_1_Instr_16__hier0_bF_buf3), .Y(datapath_1_Instr_16_bF_buf45_) );
BUFX2 BUFX2_586 ( .A(datapath_1_Instr_16__hier0_bF_buf1), .Y(datapath_1_Instr_16_bF_buf44_) );
BUFX2 BUFX2_587 ( .A(datapath_1_Instr_16__hier0_bF_buf4), .Y(datapath_1_Instr_16_bF_buf43_) );
BUFX2 BUFX2_588 ( .A(datapath_1_Instr_16__hier0_bF_buf3), .Y(datapath_1_Instr_16_bF_buf42_) );
BUFX2 BUFX2_589 ( .A(datapath_1_Instr_16__hier0_bF_buf5), .Y(datapath_1_Instr_16_bF_buf41_) );
BUFX2 BUFX2_590 ( .A(datapath_1_Instr_16__hier0_bF_buf4), .Y(datapath_1_Instr_16_bF_buf40_) );
BUFX2 BUFX2_591 ( .A(datapath_1_Instr_16__hier0_bF_buf3), .Y(datapath_1_Instr_16_bF_buf39_) );
BUFX2 BUFX2_592 ( .A(datapath_1_Instr_16__hier0_bF_buf3), .Y(datapath_1_Instr_16_bF_buf38_) );
BUFX2 BUFX2_593 ( .A(datapath_1_Instr_16__hier0_bF_buf1), .Y(datapath_1_Instr_16_bF_buf37_) );
BUFX2 BUFX2_594 ( .A(datapath_1_Instr_16__hier0_bF_buf1), .Y(datapath_1_Instr_16_bF_buf36_) );
BUFX2 BUFX2_595 ( .A(datapath_1_Instr_16__hier0_bF_buf1), .Y(datapath_1_Instr_16_bF_buf35_) );
BUFX2 BUFX2_596 ( .A(datapath_1_Instr_16__hier0_bF_buf1), .Y(datapath_1_Instr_16_bF_buf34_) );
BUFX2 BUFX2_597 ( .A(datapath_1_Instr_16__hier0_bF_buf4), .Y(datapath_1_Instr_16_bF_buf33_) );
BUFX2 BUFX2_598 ( .A(datapath_1_Instr_16__hier0_bF_buf0), .Y(datapath_1_Instr_16_bF_buf32_) );
BUFX2 BUFX2_599 ( .A(datapath_1_Instr_16__hier0_bF_buf0), .Y(datapath_1_Instr_16_bF_buf31_) );
BUFX2 BUFX2_600 ( .A(datapath_1_Instr_16__hier0_bF_buf3), .Y(datapath_1_Instr_16_bF_buf30_) );
BUFX2 BUFX2_601 ( .A(datapath_1_Instr_16__hier0_bF_buf3), .Y(datapath_1_Instr_16_bF_buf29_) );
BUFX2 BUFX2_602 ( .A(datapath_1_Instr_16__hier0_bF_buf4), .Y(datapath_1_Instr_16_bF_buf28_) );
BUFX2 BUFX2_603 ( .A(datapath_1_Instr_16__hier0_bF_buf0), .Y(datapath_1_Instr_16_bF_buf27_) );
BUFX2 BUFX2_604 ( .A(datapath_1_Instr_16__hier0_bF_buf0), .Y(datapath_1_Instr_16_bF_buf26_) );
BUFX2 BUFX2_605 ( .A(datapath_1_Instr_16__hier0_bF_buf0), .Y(datapath_1_Instr_16_bF_buf25_) );
BUFX2 BUFX2_606 ( .A(datapath_1_Instr_16__hier0_bF_buf4), .Y(datapath_1_Instr_16_bF_buf24_) );
BUFX2 BUFX2_607 ( .A(datapath_1_Instr_16__hier0_bF_buf0), .Y(datapath_1_Instr_16_bF_buf23_) );
BUFX2 BUFX2_608 ( .A(datapath_1_Instr_16__hier0_bF_buf1), .Y(datapath_1_Instr_16_bF_buf22_) );
BUFX2 BUFX2_609 ( .A(datapath_1_Instr_16__hier0_bF_buf4), .Y(datapath_1_Instr_16_bF_buf21_) );
BUFX2 BUFX2_610 ( .A(datapath_1_Instr_16__hier0_bF_buf2), .Y(datapath_1_Instr_16_bF_buf20_) );
BUFX2 BUFX2_611 ( .A(datapath_1_Instr_16__hier0_bF_buf0), .Y(datapath_1_Instr_16_bF_buf19_) );
BUFX2 BUFX2_612 ( .A(datapath_1_Instr_16__hier0_bF_buf6), .Y(datapath_1_Instr_16_bF_buf18_) );
BUFX2 BUFX2_613 ( .A(datapath_1_Instr_16__hier0_bF_buf2), .Y(datapath_1_Instr_16_bF_buf17_) );
BUFX2 BUFX2_614 ( .A(datapath_1_Instr_16__hier0_bF_buf6), .Y(datapath_1_Instr_16_bF_buf16_) );
BUFX2 BUFX2_615 ( .A(datapath_1_Instr_16__hier0_bF_buf2), .Y(datapath_1_Instr_16_bF_buf15_) );
BUFX2 BUFX2_616 ( .A(datapath_1_Instr_16__hier0_bF_buf5), .Y(datapath_1_Instr_16_bF_buf14_) );
BUFX2 BUFX2_617 ( .A(datapath_1_Instr_16__hier0_bF_buf5), .Y(datapath_1_Instr_16_bF_buf13_) );
BUFX2 BUFX2_618 ( .A(datapath_1_Instr_16__hier0_bF_buf6), .Y(datapath_1_Instr_16_bF_buf12_) );
BUFX2 BUFX2_619 ( .A(datapath_1_Instr_16__hier0_bF_buf5), .Y(datapath_1_Instr_16_bF_buf11_) );
BUFX2 BUFX2_620 ( .A(datapath_1_Instr_16__hier0_bF_buf6), .Y(datapath_1_Instr_16_bF_buf10_) );
BUFX2 BUFX2_621 ( .A(datapath_1_Instr_16__hier0_bF_buf6), .Y(datapath_1_Instr_16_bF_buf9_) );
BUFX2 BUFX2_622 ( .A(datapath_1_Instr_16__hier0_bF_buf2), .Y(datapath_1_Instr_16_bF_buf8_) );
BUFX2 BUFX2_623 ( .A(datapath_1_Instr_16__hier0_bF_buf6), .Y(datapath_1_Instr_16_bF_buf7_) );
BUFX2 BUFX2_624 ( .A(datapath_1_Instr_16__hier0_bF_buf6), .Y(datapath_1_Instr_16_bF_buf6_) );
BUFX2 BUFX2_625 ( .A(datapath_1_Instr_16__hier0_bF_buf2), .Y(datapath_1_Instr_16_bF_buf5_) );
BUFX2 BUFX2_626 ( .A(datapath_1_Instr_16__hier0_bF_buf2), .Y(datapath_1_Instr_16_bF_buf4_) );
BUFX2 BUFX2_627 ( .A(datapath_1_Instr_16__hier0_bF_buf5), .Y(datapath_1_Instr_16_bF_buf3_) );
BUFX2 BUFX2_628 ( .A(datapath_1_Instr_16__hier0_bF_buf2), .Y(datapath_1_Instr_16_bF_buf2_) );
BUFX2 BUFX2_629 ( .A(datapath_1_Instr_16__hier0_bF_buf1), .Y(datapath_1_Instr_16_bF_buf1_) );
BUFX2 BUFX2_630 ( .A(datapath_1_Instr_16__hier0_bF_buf5), .Y(datapath_1_Instr_16_bF_buf0_) );
BUFX2 BUFX2_631 ( .A(rst), .Y(rst_bF_buf13) );
BUFX2 BUFX2_632 ( .A(rst), .Y(rst_bF_buf12) );
BUFX2 BUFX2_633 ( .A(rst), .Y(rst_bF_buf11) );
BUFX2 BUFX2_634 ( .A(rst), .Y(rst_bF_buf10) );
BUFX2 BUFX2_635 ( .A(rst), .Y(rst_bF_buf9) );
BUFX2 BUFX2_636 ( .A(rst), .Y(rst_bF_buf8) );
BUFX2 BUFX2_637 ( .A(rst), .Y(rst_bF_buf7) );
BUFX2 BUFX2_638 ( .A(rst), .Y(rst_bF_buf6) );
BUFX2 BUFX2_639 ( .A(rst), .Y(rst_bF_buf5) );
BUFX2 BUFX2_640 ( .A(rst), .Y(rst_bF_buf4) );
BUFX2 BUFX2_641 ( .A(rst), .Y(rst_bF_buf3) );
BUFX2 BUFX2_642 ( .A(rst), .Y(rst_bF_buf2) );
BUFX2 BUFX2_643 ( .A(rst), .Y(rst_bF_buf1) );
BUFX2 BUFX2_644 ( .A(rst), .Y(rst_bF_buf0) );
BUFX2 BUFX2_645 ( .A(_5324_), .Y(_5324__bF_buf4) );
BUFX2 BUFX2_646 ( .A(_5324_), .Y(_5324__bF_buf3) );
BUFX2 BUFX2_647 ( .A(_5324_), .Y(_5324__bF_buf2) );
BUFX2 BUFX2_648 ( .A(_5324_), .Y(_5324__bF_buf1) );
BUFX2 BUFX2_649 ( .A(_5324_), .Y(_5324__bF_buf0) );
BUFX2 BUFX2_650 ( .A(ALUOp_0_), .Y(ALUOp_0_bF_buf5_) );
BUFX2 BUFX2_651 ( .A(ALUOp_0_), .Y(ALUOp_0_bF_buf4_) );
BUFX2 BUFX2_652 ( .A(ALUOp_0_), .Y(ALUOp_0_bF_buf3_) );
BUFX2 BUFX2_653 ( .A(ALUOp_0_), .Y(ALUOp_0_bF_buf2_) );
BUFX2 BUFX2_654 ( .A(ALUOp_0_), .Y(ALUOp_0_bF_buf1_) );
BUFX2 BUFX2_655 ( .A(ALUOp_0_), .Y(ALUOp_0_bF_buf0_) );
BUFX2 BUFX2_656 ( .A(_5265__hier0_bF_buf3), .Y(_5265__bF_buf98) );
BUFX2 BUFX2_657 ( .A(_5265__hier0_bF_buf8), .Y(_5265__bF_buf97) );
BUFX2 BUFX2_658 ( .A(_5265__hier0_bF_buf4), .Y(_5265__bF_buf96) );
BUFX2 BUFX2_659 ( .A(_5265__hier0_bF_buf7), .Y(_5265__bF_buf95) );
BUFX2 BUFX2_660 ( .A(_5265__hier0_bF_buf4), .Y(_5265__bF_buf94) );
BUFX2 BUFX2_661 ( .A(_5265__hier0_bF_buf8), .Y(_5265__bF_buf93) );
BUFX2 BUFX2_662 ( .A(_5265__hier0_bF_buf8), .Y(_5265__bF_buf92) );
BUFX2 BUFX2_663 ( .A(_5265__hier0_bF_buf6), .Y(_5265__bF_buf91) );
BUFX2 BUFX2_664 ( .A(_5265__hier0_bF_buf1), .Y(_5265__bF_buf90) );
BUFX2 BUFX2_665 ( .A(_5265__hier0_bF_buf0), .Y(_5265__bF_buf89) );
BUFX2 BUFX2_666 ( .A(_5265__hier0_bF_buf0), .Y(_5265__bF_buf88) );
BUFX2 BUFX2_667 ( .A(_5265__hier0_bF_buf3), .Y(_5265__bF_buf87) );
BUFX2 BUFX2_668 ( .A(_5265__hier0_bF_buf4), .Y(_5265__bF_buf86) );
BUFX2 BUFX2_669 ( .A(_5265__hier0_bF_buf4), .Y(_5265__bF_buf85) );
BUFX2 BUFX2_670 ( .A(_5265__hier0_bF_buf4), .Y(_5265__bF_buf84) );
BUFX2 BUFX2_671 ( .A(_5265__hier0_bF_buf6), .Y(_5265__bF_buf83) );
BUFX2 BUFX2_672 ( .A(_5265__hier0_bF_buf7), .Y(_5265__bF_buf82) );
BUFX2 BUFX2_673 ( .A(_5265__hier0_bF_buf5), .Y(_5265__bF_buf81) );
BUFX2 BUFX2_674 ( .A(_5265__hier0_bF_buf2), .Y(_5265__bF_buf80) );
BUFX2 BUFX2_675 ( .A(_5265__hier0_bF_buf5), .Y(_5265__bF_buf79) );
BUFX2 BUFX2_676 ( .A(_5265__hier0_bF_buf0), .Y(_5265__bF_buf78) );
BUFX2 BUFX2_677 ( .A(_5265__hier0_bF_buf3), .Y(_5265__bF_buf77) );
BUFX2 BUFX2_678 ( .A(_5265__hier0_bF_buf4), .Y(_5265__bF_buf76) );
BUFX2 BUFX2_679 ( .A(_5265__hier0_bF_buf7), .Y(_5265__bF_buf75) );
BUFX2 BUFX2_680 ( .A(_5265__hier0_bF_buf6), .Y(_5265__bF_buf74) );
BUFX2 BUFX2_681 ( .A(_5265__hier0_bF_buf1), .Y(_5265__bF_buf73) );
BUFX2 BUFX2_682 ( .A(_5265__hier0_bF_buf8), .Y(_5265__bF_buf72) );
BUFX2 BUFX2_683 ( .A(_5265__hier0_bF_buf2), .Y(_5265__bF_buf71) );
BUFX2 BUFX2_684 ( .A(_5265__hier0_bF_buf4), .Y(_5265__bF_buf70) );
BUFX2 BUFX2_685 ( .A(_5265__hier0_bF_buf0), .Y(_5265__bF_buf69) );
BUFX2 BUFX2_686 ( .A(_5265__hier0_bF_buf3), .Y(_5265__bF_buf68) );
BUFX2 BUFX2_687 ( .A(_5265__hier0_bF_buf2), .Y(_5265__bF_buf67) );
BUFX2 BUFX2_688 ( .A(_5265__hier0_bF_buf7), .Y(_5265__bF_buf66) );
BUFX2 BUFX2_689 ( .A(_5265__hier0_bF_buf8), .Y(_5265__bF_buf65) );
BUFX2 BUFX2_690 ( .A(_5265__hier0_bF_buf1), .Y(_5265__bF_buf64) );
BUFX2 BUFX2_691 ( .A(_5265__hier0_bF_buf8), .Y(_5265__bF_buf63) );
BUFX2 BUFX2_692 ( .A(_5265__hier0_bF_buf4), .Y(_5265__bF_buf62) );
BUFX2 BUFX2_693 ( .A(_5265__hier0_bF_buf7), .Y(_5265__bF_buf61) );
BUFX2 BUFX2_694 ( .A(_5265__hier0_bF_buf1), .Y(_5265__bF_buf60) );
BUFX2 BUFX2_695 ( .A(_5265__hier0_bF_buf1), .Y(_5265__bF_buf59) );
BUFX2 BUFX2_696 ( .A(_5265__hier0_bF_buf5), .Y(_5265__bF_buf58) );
BUFX2 BUFX2_697 ( .A(_5265__hier0_bF_buf4), .Y(_5265__bF_buf57) );
BUFX2 BUFX2_698 ( .A(_5265__hier0_bF_buf6), .Y(_5265__bF_buf56) );
BUFX2 BUFX2_699 ( .A(_5265__hier0_bF_buf8), .Y(_5265__bF_buf55) );
BUFX2 BUFX2_700 ( .A(_5265__hier0_bF_buf7), .Y(_5265__bF_buf54) );
BUFX2 BUFX2_701 ( .A(_5265__hier0_bF_buf2), .Y(_5265__bF_buf53) );
BUFX2 BUFX2_702 ( .A(_5265__hier0_bF_buf3), .Y(_5265__bF_buf52) );
BUFX2 BUFX2_703 ( .A(_5265__hier0_bF_buf3), .Y(_5265__bF_buf51) );
BUFX2 BUFX2_704 ( .A(_5265__hier0_bF_buf6), .Y(_5265__bF_buf50) );
BUFX2 BUFX2_705 ( .A(_5265__hier0_bF_buf7), .Y(_5265__bF_buf49) );
BUFX2 BUFX2_706 ( .A(_5265__hier0_bF_buf1), .Y(_5265__bF_buf48) );
BUFX2 BUFX2_707 ( .A(_5265__hier0_bF_buf5), .Y(_5265__bF_buf47) );
BUFX2 BUFX2_708 ( .A(_5265__hier0_bF_buf7), .Y(_5265__bF_buf46) );
BUFX2 BUFX2_709 ( .A(_5265__hier0_bF_buf8), .Y(_5265__bF_buf45) );
BUFX2 BUFX2_710 ( .A(_5265__hier0_bF_buf8), .Y(_5265__bF_buf44) );
BUFX2 BUFX2_711 ( .A(_5265__hier0_bF_buf6), .Y(_5265__bF_buf43) );
BUFX2 BUFX2_712 ( .A(_5265__hier0_bF_buf3), .Y(_5265__bF_buf42) );
BUFX2 BUFX2_713 ( .A(_5265__hier0_bF_buf2), .Y(_5265__bF_buf41) );
BUFX2 BUFX2_714 ( .A(_5265__hier0_bF_buf2), .Y(_5265__bF_buf40) );
BUFX2 BUFX2_715 ( .A(_5265__hier0_bF_buf4), .Y(_5265__bF_buf39) );
BUFX2 BUFX2_716 ( .A(_5265__hier0_bF_buf1), .Y(_5265__bF_buf38) );
BUFX2 BUFX2_717 ( .A(_5265__hier0_bF_buf5), .Y(_5265__bF_buf37) );
BUFX2 BUFX2_718 ( .A(_5265__hier0_bF_buf0), .Y(_5265__bF_buf36) );
BUFX2 BUFX2_719 ( .A(_5265__hier0_bF_buf6), .Y(_5265__bF_buf35) );
BUFX2 BUFX2_720 ( .A(_5265__hier0_bF_buf2), .Y(_5265__bF_buf34) );
BUFX2 BUFX2_721 ( .A(_5265__hier0_bF_buf5), .Y(_5265__bF_buf33) );
BUFX2 BUFX2_722 ( .A(_5265__hier0_bF_buf2), .Y(_5265__bF_buf32) );
BUFX2 BUFX2_723 ( .A(_5265__hier0_bF_buf1), .Y(_5265__bF_buf31) );
BUFX2 BUFX2_724 ( .A(_5265__hier0_bF_buf4), .Y(_5265__bF_buf30) );
BUFX2 BUFX2_725 ( .A(_5265__hier0_bF_buf5), .Y(_5265__bF_buf29) );
BUFX2 BUFX2_726 ( .A(_5265__hier0_bF_buf7), .Y(_5265__bF_buf28) );
BUFX2 BUFX2_727 ( .A(_5265__hier0_bF_buf3), .Y(_5265__bF_buf27) );
BUFX2 BUFX2_728 ( .A(_5265__hier0_bF_buf6), .Y(_5265__bF_buf26) );
BUFX2 BUFX2_729 ( .A(_5265__hier0_bF_buf8), .Y(_5265__bF_buf25) );
BUFX2 BUFX2_730 ( .A(_5265__hier0_bF_buf2), .Y(_5265__bF_buf24) );
BUFX2 BUFX2_731 ( .A(_5265__hier0_bF_buf6), .Y(_5265__bF_buf23) );
BUFX2 BUFX2_732 ( .A(_5265__hier0_bF_buf1), .Y(_5265__bF_buf22) );
BUFX2 BUFX2_733 ( .A(_5265__hier0_bF_buf3), .Y(_5265__bF_buf21) );
BUFX2 BUFX2_734 ( .A(_5265__hier0_bF_buf0), .Y(_5265__bF_buf20) );
BUFX2 BUFX2_735 ( .A(_5265__hier0_bF_buf0), .Y(_5265__bF_buf19) );
BUFX2 BUFX2_736 ( .A(_5265__hier0_bF_buf1), .Y(_5265__bF_buf18) );
BUFX2 BUFX2_737 ( .A(_5265__hier0_bF_buf5), .Y(_5265__bF_buf17) );
BUFX2 BUFX2_738 ( .A(_5265__hier0_bF_buf2), .Y(_5265__bF_buf16) );
BUFX2 BUFX2_739 ( .A(_5265__hier0_bF_buf5), .Y(_5265__bF_buf15) );
BUFX2 BUFX2_740 ( .A(_5265__hier0_bF_buf0), .Y(_5265__bF_buf14) );
BUFX2 BUFX2_741 ( .A(_5265__hier0_bF_buf6), .Y(_5265__bF_buf13) );
BUFX2 BUFX2_742 ( .A(_5265__hier0_bF_buf1), .Y(_5265__bF_buf12) );
BUFX2 BUFX2_743 ( .A(_5265__hier0_bF_buf2), .Y(_5265__bF_buf11) );
BUFX2 BUFX2_744 ( .A(_5265__hier0_bF_buf0), .Y(_5265__bF_buf10) );
BUFX2 BUFX2_745 ( .A(_5265__hier0_bF_buf0), .Y(_5265__bF_buf9) );
BUFX2 BUFX2_746 ( .A(_5265__hier0_bF_buf7), .Y(_5265__bF_buf8) );
BUFX2 BUFX2_747 ( .A(_5265__hier0_bF_buf3), .Y(_5265__bF_buf7) );
BUFX2 BUFX2_748 ( .A(_5265__hier0_bF_buf3), .Y(_5265__bF_buf6) );
BUFX2 BUFX2_749 ( .A(_5265__hier0_bF_buf8), .Y(_5265__bF_buf5) );
BUFX2 BUFX2_750 ( .A(_5265__hier0_bF_buf7), .Y(_5265__bF_buf4) );
BUFX2 BUFX2_751 ( .A(_5265__hier0_bF_buf0), .Y(_5265__bF_buf3) );
BUFX2 BUFX2_752 ( .A(_5265__hier0_bF_buf5), .Y(_5265__bF_buf2) );
BUFX2 BUFX2_753 ( .A(_5265__hier0_bF_buf5), .Y(_5265__bF_buf1) );
BUFX2 BUFX2_754 ( .A(_5265__hier0_bF_buf6), .Y(_5265__bF_buf0) );
BUFX2 BUFX2_755 ( .A(_5779_), .Y(_5779__bF_buf7) );
BUFX2 BUFX2_756 ( .A(_5779_), .Y(_5779__bF_buf6) );
BUFX2 BUFX2_757 ( .A(_5779_), .Y(_5779__bF_buf5) );
BUFX2 BUFX2_758 ( .A(_5779_), .Y(_5779__bF_buf4) );
BUFX2 BUFX2_759 ( .A(_5779_), .Y(_5779__bF_buf3) );
BUFX2 BUFX2_760 ( .A(_5779_), .Y(_5779__bF_buf2) );
BUFX2 BUFX2_761 ( .A(_5779_), .Y(_5779__bF_buf1) );
BUFX2 BUFX2_762 ( .A(_5779_), .Y(_5779__bF_buf0) );
BUFX2 BUFX2_763 ( .A(_6852_), .Y(_6852__bF_buf4) );
BUFX2 BUFX2_764 ( .A(_6852_), .Y(_6852__bF_buf3) );
BUFX2 BUFX2_765 ( .A(_6852_), .Y(_6852__bF_buf2) );
BUFX2 BUFX2_766 ( .A(_6852_), .Y(_6852__bF_buf1) );
BUFX2 BUFX2_767 ( .A(_6852_), .Y(_6852__bF_buf0) );
BUFX2 BUFX2_768 ( .A(_5512_), .Y(_5512__bF_buf7) );
BUFX2 BUFX2_769 ( .A(_5512_), .Y(_5512__bF_buf6) );
BUFX2 BUFX2_770 ( .A(_5512_), .Y(_5512__bF_buf5) );
BUFX2 BUFX2_771 ( .A(_5512_), .Y(_5512__bF_buf4) );
BUFX2 BUFX2_772 ( .A(_5512_), .Y(_5512__bF_buf3) );
BUFX2 BUFX2_773 ( .A(_5512_), .Y(_5512__bF_buf2) );
BUFX2 BUFX2_774 ( .A(_5512_), .Y(_5512__bF_buf1) );
BUFX2 BUFX2_775 ( .A(_5512_), .Y(_5512__bF_buf0) );
BUFX2 BUFX2_776 ( .A(_1890__hier0_bF_buf5), .Y(_1890__bF_buf47) );
BUFX2 BUFX2_777 ( .A(_1890__hier0_bF_buf3), .Y(_1890__bF_buf46) );
BUFX2 BUFX2_778 ( .A(_1890__hier0_bF_buf3), .Y(_1890__bF_buf45) );
BUFX2 BUFX2_779 ( .A(_1890__hier0_bF_buf2), .Y(_1890__bF_buf44) );
BUFX2 BUFX2_780 ( .A(_1890__hier0_bF_buf2), .Y(_1890__bF_buf43) );
BUFX2 BUFX2_781 ( .A(_1890__hier0_bF_buf5), .Y(_1890__bF_buf42) );
BUFX2 BUFX2_782 ( .A(_1890__hier0_bF_buf4), .Y(_1890__bF_buf41) );
BUFX2 BUFX2_783 ( .A(_1890__hier0_bF_buf1), .Y(_1890__bF_buf40) );
BUFX2 BUFX2_784 ( .A(_1890__hier0_bF_buf1), .Y(_1890__bF_buf39) );
BUFX2 BUFX2_785 ( .A(_1890__hier0_bF_buf0), .Y(_1890__bF_buf38) );
BUFX2 BUFX2_786 ( .A(_1890__hier0_bF_buf1), .Y(_1890__bF_buf37) );
BUFX2 BUFX2_787 ( .A(_1890__hier0_bF_buf0), .Y(_1890__bF_buf36) );
BUFX2 BUFX2_788 ( .A(_1890__hier0_bF_buf2), .Y(_1890__bF_buf35) );
BUFX2 BUFX2_789 ( .A(_1890__hier0_bF_buf1), .Y(_1890__bF_buf34) );
BUFX2 BUFX2_790 ( .A(_1890__hier0_bF_buf3), .Y(_1890__bF_buf33) );
BUFX2 BUFX2_791 ( .A(_1890__hier0_bF_buf2), .Y(_1890__bF_buf32) );
BUFX2 BUFX2_792 ( .A(_1890__hier0_bF_buf2), .Y(_1890__bF_buf31) );
BUFX2 BUFX2_793 ( .A(_1890__hier0_bF_buf3), .Y(_1890__bF_buf30) );
BUFX2 BUFX2_794 ( .A(_1890__hier0_bF_buf5), .Y(_1890__bF_buf29) );
BUFX2 BUFX2_795 ( .A(_1890__hier0_bF_buf0), .Y(_1890__bF_buf28) );
BUFX2 BUFX2_796 ( .A(_1890__hier0_bF_buf0), .Y(_1890__bF_buf27) );
BUFX2 BUFX2_797 ( .A(_1890__hier0_bF_buf4), .Y(_1890__bF_buf26) );
BUFX2 BUFX2_798 ( .A(_1890__hier0_bF_buf2), .Y(_1890__bF_buf25) );
BUFX2 BUFX2_799 ( .A(_1890__hier0_bF_buf1), .Y(_1890__bF_buf24) );
BUFX2 BUFX2_800 ( .A(_1890__hier0_bF_buf5), .Y(_1890__bF_buf23) );
BUFX2 BUFX2_801 ( .A(_1890__hier0_bF_buf1), .Y(_1890__bF_buf22) );
BUFX2 BUFX2_802 ( .A(_1890__hier0_bF_buf4), .Y(_1890__bF_buf21) );
BUFX2 BUFX2_803 ( .A(_1890__hier0_bF_buf0), .Y(_1890__bF_buf20) );
BUFX2 BUFX2_804 ( .A(_1890__hier0_bF_buf5), .Y(_1890__bF_buf19) );
BUFX2 BUFX2_805 ( .A(_1890__hier0_bF_buf4), .Y(_1890__bF_buf18) );
BUFX2 BUFX2_806 ( .A(_1890__hier0_bF_buf5), .Y(_1890__bF_buf17) );
BUFX2 BUFX2_807 ( .A(_1890__hier0_bF_buf4), .Y(_1890__bF_buf16) );
BUFX2 BUFX2_808 ( .A(_1890__hier0_bF_buf3), .Y(_1890__bF_buf15) );
BUFX2 BUFX2_809 ( .A(_1890__hier0_bF_buf3), .Y(_1890__bF_buf14) );
BUFX2 BUFX2_810 ( .A(_1890__hier0_bF_buf3), .Y(_1890__bF_buf13) );
BUFX2 BUFX2_811 ( .A(_1890__hier0_bF_buf4), .Y(_1890__bF_buf12) );
BUFX2 BUFX2_812 ( .A(_1890__hier0_bF_buf2), .Y(_1890__bF_buf11) );
BUFX2 BUFX2_813 ( .A(_1890__hier0_bF_buf0), .Y(_1890__bF_buf10) );
BUFX2 BUFX2_814 ( .A(_1890__hier0_bF_buf1), .Y(_1890__bF_buf9) );
BUFX2 BUFX2_815 ( .A(_1890__hier0_bF_buf4), .Y(_1890__bF_buf8) );
BUFX2 BUFX2_816 ( .A(_1890__hier0_bF_buf0), .Y(_1890__bF_buf7) );
BUFX2 BUFX2_817 ( .A(_1890__hier0_bF_buf5), .Y(_1890__bF_buf6) );
BUFX2 BUFX2_818 ( .A(_1890__hier0_bF_buf3), .Y(_1890__bF_buf5) );
BUFX2 BUFX2_819 ( .A(_1890__hier0_bF_buf1), .Y(_1890__bF_buf4) );
BUFX2 BUFX2_820 ( .A(_1890__hier0_bF_buf4), .Y(_1890__bF_buf3) );
BUFX2 BUFX2_821 ( .A(_1890__hier0_bF_buf2), .Y(_1890__bF_buf2) );
BUFX2 BUFX2_822 ( .A(_1890__hier0_bF_buf0), .Y(_1890__bF_buf1) );
BUFX2 BUFX2_823 ( .A(_1890__hier0_bF_buf5), .Y(_1890__bF_buf0) );
BUFX2 BUFX2_824 ( .A(_6984_), .Y(_6984__bF_buf4) );
BUFX2 BUFX2_825 ( .A(_6984_), .Y(_6984__bF_buf3) );
BUFX2 BUFX2_826 ( .A(_6984_), .Y(_6984__bF_buf2) );
BUFX2 BUFX2_827 ( .A(_6984_), .Y(_6984__bF_buf1) );
BUFX2 BUFX2_828 ( .A(_6984_), .Y(_6984__bF_buf0) );
BUFX2 BUFX2_829 ( .A(_6182_), .Y(_6182__bF_buf7) );
BUFX2 BUFX2_830 ( .A(_6182_), .Y(_6182__bF_buf6) );
BUFX2 BUFX2_831 ( .A(_6182_), .Y(_6182__bF_buf5) );
BUFX2 BUFX2_832 ( .A(_6182_), .Y(_6182__bF_buf4) );
BUFX2 BUFX2_833 ( .A(_6182_), .Y(_6182__bF_buf3) );
BUFX2 BUFX2_834 ( .A(_6182_), .Y(_6182__bF_buf2) );
BUFX2 BUFX2_835 ( .A(_6182_), .Y(_6182__bF_buf1) );
BUFX2 BUFX2_836 ( .A(_6182_), .Y(_6182__bF_buf0) );
BUFX2 BUFX2_837 ( .A(_5318_), .Y(_5318__bF_buf4) );
BUFX2 BUFX2_838 ( .A(_5318_), .Y(_5318__bF_buf3) );
BUFX2 BUFX2_839 ( .A(_5318_), .Y(_5318__bF_buf2) );
BUFX2 BUFX2_840 ( .A(_5318_), .Y(_5318__bF_buf1) );
BUFX2 BUFX2_841 ( .A(_5318_), .Y(_5318__bF_buf0) );
BUFX2 BUFX2_842 ( .A(_1887_), .Y(_1887__bF_buf4) );
BUFX2 BUFX2_843 ( .A(_1887_), .Y(_1887__bF_buf3) );
BUFX2 BUFX2_844 ( .A(_1887_), .Y(_1887__bF_buf2) );
BUFX2 BUFX2_845 ( .A(_1887_), .Y(_1887__bF_buf1) );
BUFX2 BUFX2_846 ( .A(_1887_), .Y(_1887__bF_buf0) );
BUFX2 BUFX2_847 ( .A(_5679_), .Y(_5679__bF_buf7) );
BUFX2 BUFX2_848 ( .A(_5679_), .Y(_5679__bF_buf6) );
BUFX2 BUFX2_849 ( .A(_5679_), .Y(_5679__bF_buf5) );
BUFX2 BUFX2_850 ( .A(_5679_), .Y(_5679__bF_buf4) );
BUFX2 BUFX2_851 ( .A(_5679_), .Y(_5679__bF_buf3) );
BUFX2 BUFX2_852 ( .A(_5679_), .Y(_5679__bF_buf2) );
BUFX2 BUFX2_853 ( .A(_5679_), .Y(_5679__bF_buf1) );
BUFX2 BUFX2_854 ( .A(_5679_), .Y(_5679__bF_buf0) );
BUFX2 BUFX2_855 ( .A(PCSource_1_), .Y(PCSource_1_bF_buf5_) );
BUFX2 BUFX2_856 ( .A(PCSource_1_), .Y(PCSource_1_bF_buf4_) );
BUFX2 BUFX2_857 ( .A(PCSource_1_), .Y(PCSource_1_bF_buf3_) );
BUFX2 BUFX2_858 ( .A(PCSource_1_), .Y(PCSource_1_bF_buf2_) );
BUFX2 BUFX2_859 ( .A(PCSource_1_), .Y(PCSource_1_bF_buf1_) );
BUFX2 BUFX2_860 ( .A(PCSource_1_), .Y(PCSource_1_bF_buf0_) );
BUFX2 BUFX2_861 ( .A(_1884_), .Y(_1884__bF_buf9) );
BUFX2 BUFX2_862 ( .A(_1884_), .Y(_1884__bF_buf8) );
BUFX2 BUFX2_863 ( .A(_1884_), .Y(_1884__bF_buf7) );
BUFX2 BUFX2_864 ( .A(_1884_), .Y(_1884__bF_buf6) );
BUFX2 BUFX2_865 ( .A(_1884_), .Y(_1884__bF_buf5) );
BUFX2 BUFX2_866 ( .A(_1884_), .Y(_1884__bF_buf4) );
BUFX2 BUFX2_867 ( .A(_1884_), .Y(_1884__bF_buf3) );
BUFX2 BUFX2_868 ( .A(_1884_), .Y(_1884__bF_buf2) );
BUFX2 BUFX2_869 ( .A(_1884_), .Y(_1884__bF_buf1) );
BUFX2 BUFX2_870 ( .A(_1884_), .Y(_1884__bF_buf0) );
BUFX2 BUFX2_871 ( .A(_5294_), .Y(_5294__bF_buf4) );
BUFX2 BUFX2_872 ( .A(_5294_), .Y(_5294__bF_buf3) );
BUFX2 BUFX2_873 ( .A(_5294_), .Y(_5294__bF_buf2) );
BUFX2 BUFX2_874 ( .A(_5294_), .Y(_5294__bF_buf1) );
BUFX2 BUFX2_875 ( .A(_5294_), .Y(_5294__bF_buf0) );
BUFX2 BUFX2_876 ( .A(_6079_), .Y(_6079__bF_buf7) );
BUFX2 BUFX2_877 ( .A(_6079_), .Y(_6079__bF_buf6) );
BUFX2 BUFX2_878 ( .A(_6079_), .Y(_6079__bF_buf5) );
BUFX2 BUFX2_879 ( .A(_6079_), .Y(_6079__bF_buf4) );
BUFX2 BUFX2_880 ( .A(_6079_), .Y(_6079__bF_buf3) );
BUFX2 BUFX2_881 ( .A(_6079_), .Y(_6079__bF_buf2) );
BUFX2 BUFX2_882 ( .A(_6079_), .Y(_6079__bF_buf1) );
BUFX2 BUFX2_883 ( .A(_6079_), .Y(_6079__bF_buf0) );
BUFX2 BUFX2_884 ( .A(_240_), .Y(_240__bF_buf4) );
BUFX2 BUFX2_885 ( .A(_240_), .Y(_240__bF_buf3) );
BUFX2 BUFX2_886 ( .A(_240_), .Y(_240__bF_buf2) );
BUFX2 BUFX2_887 ( .A(_240_), .Y(_240__bF_buf1) );
BUFX2 BUFX2_888 ( .A(_240_), .Y(_240__bF_buf0) );
BUFX2 BUFX2_889 ( .A(_5312_), .Y(_5312__bF_buf4) );
BUFX2 BUFX2_890 ( .A(_5312_), .Y(_5312__bF_buf3) );
BUFX2 BUFX2_891 ( .A(_5312_), .Y(_5312__bF_buf2) );
BUFX2 BUFX2_892 ( .A(_5312_), .Y(_5312__bF_buf1) );
BUFX2 BUFX2_893 ( .A(_5312_), .Y(_5312__bF_buf0) );
BUFX2 BUFX2_894 ( .A(_237_), .Y(_237__bF_buf3) );
BUFX2 BUFX2_895 ( .A(_237_), .Y(_237__bF_buf2) );
BUFX2 BUFX2_896 ( .A(_237_), .Y(_237__bF_buf1) );
BUFX2 BUFX2_897 ( .A(_237_), .Y(_237__bF_buf0) );
BUFX2 BUFX2_898 ( .A(_5479_), .Y(_5479__bF_buf7) );
BUFX2 BUFX2_899 ( .A(_5479_), .Y(_5479__bF_buf6) );
BUFX2 BUFX2_900 ( .A(_5479_), .Y(_5479__bF_buf5) );
BUFX2 BUFX2_901 ( .A(_5479_), .Y(_5479__bF_buf4) );
BUFX2 BUFX2_902 ( .A(_5479_), .Y(_5479__bF_buf3) );
BUFX2 BUFX2_903 ( .A(_5479_), .Y(_5479__bF_buf2) );
BUFX2 BUFX2_904 ( .A(_5479_), .Y(_5479__bF_buf1) );
BUFX2 BUFX2_905 ( .A(_5479_), .Y(_5479__bF_buf0) );
BUFX2 BUFX2_906 ( .A(_5288_), .Y(_5288__bF_buf4) );
BUFX2 BUFX2_907 ( .A(_5288_), .Y(_5288__bF_buf3) );
BUFX2 BUFX2_908 ( .A(_5288_), .Y(_5288__bF_buf2) );
BUFX2 BUFX2_909 ( .A(_5288_), .Y(_5288__bF_buf1) );
BUFX2 BUFX2_910 ( .A(_5288_), .Y(_5288__bF_buf0) );
BUFX2 BUFX2_911 ( .A(MemtoReg), .Y(MemtoReg_bF_buf7) );
BUFX2 BUFX2_912 ( .A(MemtoReg), .Y(MemtoReg_bF_buf6) );
BUFX2 BUFX2_913 ( .A(MemtoReg), .Y(MemtoReg_bF_buf5) );
BUFX2 BUFX2_914 ( .A(MemtoReg), .Y(MemtoReg_bF_buf4) );
BUFX2 BUFX2_915 ( .A(MemtoReg), .Y(MemtoReg_bF_buf3) );
BUFX2 BUFX2_916 ( .A(MemtoReg), .Y(MemtoReg_bF_buf2) );
BUFX2 BUFX2_917 ( .A(MemtoReg), .Y(MemtoReg_bF_buf1) );
BUFX2 BUFX2_918 ( .A(MemtoReg), .Y(MemtoReg_bF_buf0) );
BUFX2 BUFX2_919 ( .A(_6552_), .Y(_6552__bF_buf4) );
BUFX2 BUFX2_920 ( .A(_6552_), .Y(_6552__bF_buf3) );
BUFX2 BUFX2_921 ( .A(_6552_), .Y(_6552__bF_buf2) );
BUFX2 BUFX2_922 ( .A(_6552_), .Y(_6552__bF_buf1) );
BUFX2 BUFX2_923 ( .A(_6552_), .Y(_6552__bF_buf0) );
BUFX2 BUFX2_924 ( .A(_5306_), .Y(_5306__bF_buf4) );
BUFX2 BUFX2_925 ( .A(_5306_), .Y(_5306__bF_buf3) );
BUFX2 BUFX2_926 ( .A(_5306_), .Y(_5306__bF_buf2) );
BUFX2 BUFX2_927 ( .A(_5306_), .Y(_5306__bF_buf1) );
BUFX2 BUFX2_928 ( .A(_5306_), .Y(_5306__bF_buf0) );
BUFX2 BUFX2_929 ( .A(_6549_), .Y(_6549__bF_buf4) );
BUFX2 BUFX2_930 ( .A(_6549_), .Y(_6549__bF_buf3) );
BUFX2 BUFX2_931 ( .A(_6549_), .Y(_6549__bF_buf2) );
BUFX2 BUFX2_932 ( .A(_6549_), .Y(_6549__bF_buf1) );
BUFX2 BUFX2_933 ( .A(_6549_), .Y(_6549__bF_buf0) );
BUFX2 BUFX2_934 ( .A(ALUSrcA), .Y(ALUSrcA_bF_buf7) );
BUFX2 BUFX2_935 ( .A(ALUSrcA), .Y(ALUSrcA_bF_buf6) );
BUFX2 BUFX2_936 ( .A(ALUSrcA), .Y(ALUSrcA_bF_buf5) );
BUFX2 BUFX2_937 ( .A(ALUSrcA), .Y(ALUSrcA_bF_buf4) );
BUFX2 BUFX2_938 ( .A(ALUSrcA), .Y(ALUSrcA_bF_buf3) );
BUFX2 BUFX2_939 ( .A(ALUSrcA), .Y(ALUSrcA_bF_buf2) );
BUFX2 BUFX2_940 ( .A(ALUSrcA), .Y(ALUSrcA_bF_buf1) );
BUFX2 BUFX2_941 ( .A(ALUSrcA), .Y(ALUSrcA_bF_buf0) );
BUFX2 BUFX2_942 ( .A(_5282_), .Y(_5282__bF_buf4) );
BUFX2 BUFX2_943 ( .A(_5282_), .Y(_5282__bF_buf3) );
BUFX2 BUFX2_944 ( .A(_5282_), .Y(_5282__bF_buf2) );
BUFX2 BUFX2_945 ( .A(_5282_), .Y(_5282__bF_buf1) );
BUFX2 BUFX2_946 ( .A(_5282_), .Y(_5282__bF_buf0) );
BUFX2 BUFX2_947 ( .A(_5338_), .Y(_5338__bF_buf4) );
BUFX2 BUFX2_948 ( .A(_5338_), .Y(_5338__bF_buf3) );
BUFX2 BUFX2_949 ( .A(_5338_), .Y(_5338__bF_buf2) );
BUFX2 BUFX2_950 ( .A(_5338_), .Y(_5338__bF_buf1) );
BUFX2 BUFX2_951 ( .A(_5338_), .Y(_5338__bF_buf0) );
BUFX2 BUFX2_952 ( .A(_5300_), .Y(_5300__bF_buf4) );
BUFX2 BUFX2_953 ( .A(_5300_), .Y(_5300__bF_buf3) );
BUFX2 BUFX2_954 ( .A(_5300_), .Y(_5300__bF_buf2) );
BUFX2 BUFX2_955 ( .A(_5300_), .Y(_5300__bF_buf1) );
BUFX2 BUFX2_956 ( .A(_5300_), .Y(_5300__bF_buf0) );
BUFX2 BUFX2_957 ( .A(_5946_), .Y(_5946__bF_buf7) );
BUFX2 BUFX2_958 ( .A(_5946_), .Y(_5946__bF_buf6) );
BUFX2 BUFX2_959 ( .A(_5946_), .Y(_5946__bF_buf5) );
BUFX2 BUFX2_960 ( .A(_5946_), .Y(_5946__bF_buf4) );
BUFX2 BUFX2_961 ( .A(_5946_), .Y(_5946__bF_buf3) );
BUFX2 BUFX2_962 ( .A(_5946_), .Y(_5946__bF_buf2) );
BUFX2 BUFX2_963 ( .A(_5946_), .Y(_5946__bF_buf1) );
BUFX2 BUFX2_964 ( .A(_5946_), .Y(_5946__bF_buf0) );
BUFX2 BUFX2_965 ( .A(_6387_), .Y(_6387__bF_buf4) );
BUFX2 BUFX2_966 ( .A(_6387_), .Y(_6387__bF_buf3) );
BUFX2 BUFX2_967 ( .A(_6387_), .Y(_6387__bF_buf2) );
BUFX2 BUFX2_968 ( .A(_6387_), .Y(_6387__bF_buf1) );
BUFX2 BUFX2_969 ( .A(_6387_), .Y(_6387__bF_buf0) );
BUFX2 BUFX2_970 ( .A(_5276_), .Y(_5276__bF_buf4) );
BUFX2 BUFX2_971 ( .A(_5276_), .Y(_5276__bF_buf3) );
BUFX2 BUFX2_972 ( .A(_5276_), .Y(_5276__bF_buf2) );
BUFX2 BUFX2_973 ( .A(_5276_), .Y(_5276__bF_buf1) );
BUFX2 BUFX2_974 ( .A(_5276_), .Y(_5276__bF_buf0) );
BUFX2 BUFX2_975 ( .A(_3571_), .Y(_3571__bF_buf7) );
BUFX2 BUFX2_976 ( .A(_3571_), .Y(_3571__bF_buf6) );
BUFX2 BUFX2_977 ( .A(_3571_), .Y(_3571__bF_buf5) );
BUFX2 BUFX2_978 ( .A(_3571_), .Y(_3571__bF_buf4) );
BUFX2 BUFX2_979 ( .A(_3571_), .Y(_3571__bF_buf3) );
BUFX2 BUFX2_980 ( .A(_3571_), .Y(_3571__bF_buf2) );
BUFX2 BUFX2_981 ( .A(_3571_), .Y(_3571__bF_buf1) );
BUFX2 BUFX2_982 ( .A(_3571_), .Y(_3571__bF_buf0) );
BUFX2 BUFX2_983 ( .A(datapath_1_Instr_24_), .Y(datapath_1_Instr_24_bF_buf6_) );
BUFX2 BUFX2_984 ( .A(datapath_1_Instr_24_), .Y(datapath_1_Instr_24_bF_buf5_) );
BUFX2 BUFX2_985 ( .A(datapath_1_Instr_24_), .Y(datapath_1_Instr_24_bF_buf4_) );
BUFX2 BUFX2_986 ( .A(datapath_1_Instr_24_), .Y(datapath_1_Instr_24_bF_buf3_) );
BUFX2 BUFX2_987 ( .A(datapath_1_Instr_24_), .Y(datapath_1_Instr_24_bF_buf2_) );
BUFX2 BUFX2_988 ( .A(datapath_1_Instr_24_), .Y(datapath_1_Instr_24_bF_buf1_) );
BUFX2 BUFX2_989 ( .A(datapath_1_Instr_24_), .Y(datapath_1_Instr_24_bF_buf0_) );
BUFX2 BUFX2_990 ( .A(_5332_), .Y(_5332__bF_buf4) );
BUFX2 BUFX2_991 ( .A(_5332_), .Y(_5332__bF_buf3) );
BUFX2 BUFX2_992 ( .A(_5332_), .Y(_5332__bF_buf2) );
BUFX2 BUFX2_993 ( .A(_5332_), .Y(_5332__bF_buf1) );
BUFX2 BUFX2_994 ( .A(_5332_), .Y(_5332__bF_buf0) );
BUFX2 BUFX2_995 ( .A(datapath_1_Instr_21__hier0_bF_buf6), .Y(datapath_1_Instr_21_bF_buf55_) );
BUFX2 BUFX2_996 ( .A(datapath_1_Instr_21__hier0_bF_buf0), .Y(datapath_1_Instr_21_bF_buf54_) );
BUFX2 BUFX2_997 ( .A(datapath_1_Instr_21__hier0_bF_buf5), .Y(datapath_1_Instr_21_bF_buf53_) );
BUFX2 BUFX2_998 ( .A(datapath_1_Instr_21__hier0_bF_buf1), .Y(datapath_1_Instr_21_bF_buf52_) );
BUFX2 BUFX2_999 ( .A(datapath_1_Instr_21__hier0_bF_buf1), .Y(datapath_1_Instr_21_bF_buf51_) );
BUFX2 BUFX2_1000 ( .A(datapath_1_Instr_21__hier0_bF_buf0), .Y(datapath_1_Instr_21_bF_buf50_) );
BUFX2 BUFX2_1001 ( .A(datapath_1_Instr_21__hier0_bF_buf1), .Y(datapath_1_Instr_21_bF_buf49_) );
BUFX2 BUFX2_1002 ( .A(datapath_1_Instr_21__hier0_bF_buf5), .Y(datapath_1_Instr_21_bF_buf48_) );
BUFX2 BUFX2_1003 ( .A(datapath_1_Instr_21__hier0_bF_buf0), .Y(datapath_1_Instr_21_bF_buf47_) );
BUFX2 BUFX2_1004 ( .A(datapath_1_Instr_21__hier0_bF_buf3), .Y(datapath_1_Instr_21_bF_buf46_) );
BUFX2 BUFX2_1005 ( .A(datapath_1_Instr_21__hier0_bF_buf1), .Y(datapath_1_Instr_21_bF_buf45_) );
BUFX2 BUFX2_1006 ( .A(datapath_1_Instr_21__hier0_bF_buf1), .Y(datapath_1_Instr_21_bF_buf44_) );
BUFX2 BUFX2_1007 ( .A(datapath_1_Instr_21__hier0_bF_buf3), .Y(datapath_1_Instr_21_bF_buf43_) );
BUFX2 BUFX2_1008 ( .A(datapath_1_Instr_21__hier0_bF_buf3), .Y(datapath_1_Instr_21_bF_buf42_) );
BUFX2 BUFX2_1009 ( .A(datapath_1_Instr_21__hier0_bF_buf3), .Y(datapath_1_Instr_21_bF_buf41_) );
BUFX2 BUFX2_1010 ( .A(datapath_1_Instr_21__hier0_bF_buf3), .Y(datapath_1_Instr_21_bF_buf40_) );
BUFX2 BUFX2_1011 ( .A(datapath_1_Instr_21__hier0_bF_buf3), .Y(datapath_1_Instr_21_bF_buf39_) );
BUFX2 BUFX2_1012 ( .A(datapath_1_Instr_21__hier0_bF_buf3), .Y(datapath_1_Instr_21_bF_buf38_) );
BUFX2 BUFX2_1013 ( .A(datapath_1_Instr_21__hier0_bF_buf5), .Y(datapath_1_Instr_21_bF_buf37_) );
BUFX2 BUFX2_1014 ( .A(datapath_1_Instr_21__hier0_bF_buf5), .Y(datapath_1_Instr_21_bF_buf36_) );
BUFX2 BUFX2_1015 ( .A(datapath_1_Instr_21__hier0_bF_buf1), .Y(datapath_1_Instr_21_bF_buf35_) );
BUFX2 BUFX2_1016 ( .A(datapath_1_Instr_21__hier0_bF_buf5), .Y(datapath_1_Instr_21_bF_buf34_) );
BUFX2 BUFX2_1017 ( .A(datapath_1_Instr_21__hier0_bF_buf0), .Y(datapath_1_Instr_21_bF_buf33_) );
BUFX2 BUFX2_1018 ( .A(datapath_1_Instr_21__hier0_bF_buf1), .Y(datapath_1_Instr_21_bF_buf32_) );
BUFX2 BUFX2_1019 ( .A(datapath_1_Instr_21__hier0_bF_buf5), .Y(datapath_1_Instr_21_bF_buf31_) );
BUFX2 BUFX2_1020 ( .A(datapath_1_Instr_21__hier0_bF_buf0), .Y(datapath_1_Instr_21_bF_buf30_) );
BUFX2 BUFX2_1021 ( .A(datapath_1_Instr_21__hier0_bF_buf0), .Y(datapath_1_Instr_21_bF_buf29_) );
BUFX2 BUFX2_1022 ( .A(datapath_1_Instr_21__hier0_bF_buf3), .Y(datapath_1_Instr_21_bF_buf28_) );
BUFX2 BUFX2_1023 ( .A(datapath_1_Instr_21__hier0_bF_buf2), .Y(datapath_1_Instr_21_bF_buf27_) );
BUFX2 BUFX2_1024 ( .A(datapath_1_Instr_21__hier0_bF_buf0), .Y(datapath_1_Instr_21_bF_buf26_) );
BUFX2 BUFX2_1025 ( .A(datapath_1_Instr_21__hier0_bF_buf0), .Y(datapath_1_Instr_21_bF_buf25_) );
BUFX2 BUFX2_1026 ( .A(datapath_1_Instr_21__hier0_bF_buf5), .Y(datapath_1_Instr_21_bF_buf24_) );
BUFX2 BUFX2_1027 ( .A(datapath_1_Instr_21__hier0_bF_buf4), .Y(datapath_1_Instr_21_bF_buf23_) );
BUFX2 BUFX2_1028 ( .A(datapath_1_Instr_21__hier0_bF_buf6), .Y(datapath_1_Instr_21_bF_buf22_) );
BUFX2 BUFX2_1029 ( .A(datapath_1_Instr_21__hier0_bF_buf2), .Y(datapath_1_Instr_21_bF_buf21_) );
BUFX2 BUFX2_1030 ( .A(datapath_1_Instr_21__hier0_bF_buf2), .Y(datapath_1_Instr_21_bF_buf20_) );
BUFX2 BUFX2_1031 ( .A(datapath_1_Instr_21__hier0_bF_buf4), .Y(datapath_1_Instr_21_bF_buf19_) );
BUFX2 BUFX2_1032 ( .A(datapath_1_Instr_21__hier0_bF_buf4), .Y(datapath_1_Instr_21_bF_buf18_) );
BUFX2 BUFX2_1033 ( .A(datapath_1_Instr_21__hier0_bF_buf4), .Y(datapath_1_Instr_21_bF_buf17_) );
BUFX2 BUFX2_1034 ( .A(datapath_1_Instr_21__hier0_bF_buf4), .Y(datapath_1_Instr_21_bF_buf16_) );
BUFX2 BUFX2_1035 ( .A(datapath_1_Instr_21__hier0_bF_buf6), .Y(datapath_1_Instr_21_bF_buf15_) );
BUFX2 BUFX2_1036 ( .A(datapath_1_Instr_21__hier0_bF_buf4), .Y(datapath_1_Instr_21_bF_buf14_) );
BUFX2 BUFX2_1037 ( .A(datapath_1_Instr_21__hier0_bF_buf4), .Y(datapath_1_Instr_21_bF_buf13_) );
BUFX2 BUFX2_1038 ( .A(datapath_1_Instr_21__hier0_bF_buf4), .Y(datapath_1_Instr_21_bF_buf12_) );
BUFX2 BUFX2_1039 ( .A(datapath_1_Instr_21__hier0_bF_buf6), .Y(datapath_1_Instr_21_bF_buf11_) );
BUFX2 BUFX2_1040 ( .A(datapath_1_Instr_21__hier0_bF_buf6), .Y(datapath_1_Instr_21_bF_buf10_) );
BUFX2 BUFX2_1041 ( .A(datapath_1_Instr_21__hier0_bF_buf6), .Y(datapath_1_Instr_21_bF_buf9_) );
BUFX2 BUFX2_1042 ( .A(datapath_1_Instr_21__hier0_bF_buf6), .Y(datapath_1_Instr_21_bF_buf8_) );
BUFX2 BUFX2_1043 ( .A(datapath_1_Instr_21__hier0_bF_buf2), .Y(datapath_1_Instr_21_bF_buf7_) );
BUFX2 BUFX2_1044 ( .A(datapath_1_Instr_21__hier0_bF_buf6), .Y(datapath_1_Instr_21_bF_buf6_) );
BUFX2 BUFX2_1045 ( .A(datapath_1_Instr_21__hier0_bF_buf2), .Y(datapath_1_Instr_21_bF_buf5_) );
BUFX2 BUFX2_1046 ( .A(datapath_1_Instr_21__hier0_bF_buf2), .Y(datapath_1_Instr_21_bF_buf4_) );
BUFX2 BUFX2_1047 ( .A(datapath_1_Instr_21__hier0_bF_buf1), .Y(datapath_1_Instr_21_bF_buf3_) );
BUFX2 BUFX2_1048 ( .A(datapath_1_Instr_21__hier0_bF_buf2), .Y(datapath_1_Instr_21_bF_buf2_) );
BUFX2 BUFX2_1049 ( .A(datapath_1_Instr_21__hier0_bF_buf2), .Y(datapath_1_Instr_21_bF_buf1_) );
BUFX2 BUFX2_1050 ( .A(datapath_1_Instr_21__hier0_bF_buf5), .Y(datapath_1_Instr_21_bF_buf0_) );
BUFX2 BUFX2_1051 ( .A(_3565_), .Y(_3565__bF_buf4) );
BUFX2 BUFX2_1052 ( .A(_3565_), .Y(_3565__bF_buf3) );
BUFX2 BUFX2_1053 ( .A(_3565_), .Y(_3565__bF_buf2) );
BUFX2 BUFX2_1054 ( .A(_3565_), .Y(_3565__bF_buf1) );
BUFX2 BUFX2_1055 ( .A(_3565_), .Y(_3565__bF_buf0) );
BUFX2 BUFX2_1056 ( .A(datapath_1_Instr_18__hier0_bF_buf4), .Y(datapath_1_Instr_18_bF_buf44_) );
BUFX2 BUFX2_1057 ( .A(datapath_1_Instr_18__hier0_bF_buf3), .Y(datapath_1_Instr_18_bF_buf43_) );
BUFX2 BUFX2_1058 ( .A(datapath_1_Instr_18__hier0_bF_buf5), .Y(datapath_1_Instr_18_bF_buf42_) );
BUFX2 BUFX2_1059 ( .A(datapath_1_Instr_18__hier0_bF_buf3), .Y(datapath_1_Instr_18_bF_buf41_) );
BUFX2 BUFX2_1060 ( .A(datapath_1_Instr_18__hier0_bF_buf4), .Y(datapath_1_Instr_18_bF_buf40_) );
BUFX2 BUFX2_1061 ( .A(datapath_1_Instr_18__hier0_bF_buf4), .Y(datapath_1_Instr_18_bF_buf39_) );
BUFX2 BUFX2_1062 ( .A(datapath_1_Instr_18__hier0_bF_buf0), .Y(datapath_1_Instr_18_bF_buf38_) );
BUFX2 BUFX2_1063 ( .A(datapath_1_Instr_18__hier0_bF_buf4), .Y(datapath_1_Instr_18_bF_buf37_) );
BUFX2 BUFX2_1064 ( .A(datapath_1_Instr_18__hier0_bF_buf3), .Y(datapath_1_Instr_18_bF_buf36_) );
BUFX2 BUFX2_1065 ( .A(datapath_1_Instr_18__hier0_bF_buf1), .Y(datapath_1_Instr_18_bF_buf35_) );
BUFX2 BUFX2_1066 ( .A(datapath_1_Instr_18__hier0_bF_buf2), .Y(datapath_1_Instr_18_bF_buf34_) );
BUFX2 BUFX2_1067 ( .A(datapath_1_Instr_18__hier0_bF_buf1), .Y(datapath_1_Instr_18_bF_buf33_) );
BUFX2 BUFX2_1068 ( .A(datapath_1_Instr_18__hier0_bF_buf0), .Y(datapath_1_Instr_18_bF_buf32_) );
BUFX2 BUFX2_1069 ( .A(datapath_1_Instr_18__hier0_bF_buf5), .Y(datapath_1_Instr_18_bF_buf31_) );
BUFX2 BUFX2_1070 ( .A(datapath_1_Instr_18__hier0_bF_buf0), .Y(datapath_1_Instr_18_bF_buf30_) );
BUFX2 BUFX2_1071 ( .A(datapath_1_Instr_18__hier0_bF_buf4), .Y(datapath_1_Instr_18_bF_buf29_) );
BUFX2 BUFX2_1072 ( .A(datapath_1_Instr_18__hier0_bF_buf5), .Y(datapath_1_Instr_18_bF_buf28_) );
BUFX2 BUFX2_1073 ( .A(datapath_1_Instr_18__hier0_bF_buf2), .Y(datapath_1_Instr_18_bF_buf27_) );
BUFX2 BUFX2_1074 ( .A(datapath_1_Instr_18__hier0_bF_buf1), .Y(datapath_1_Instr_18_bF_buf26_) );
BUFX2 BUFX2_1075 ( .A(datapath_1_Instr_18__hier0_bF_buf0), .Y(datapath_1_Instr_18_bF_buf25_) );
BUFX2 BUFX2_1076 ( .A(datapath_1_Instr_18__hier0_bF_buf0), .Y(datapath_1_Instr_18_bF_buf24_) );
BUFX2 BUFX2_1077 ( .A(datapath_1_Instr_18__hier0_bF_buf3), .Y(datapath_1_Instr_18_bF_buf23_) );
BUFX2 BUFX2_1078 ( .A(datapath_1_Instr_18__hier0_bF_buf5), .Y(datapath_1_Instr_18_bF_buf22_) );
BUFX2 BUFX2_1079 ( .A(datapath_1_Instr_18__hier0_bF_buf1), .Y(datapath_1_Instr_18_bF_buf21_) );
BUFX2 BUFX2_1080 ( .A(datapath_1_Instr_18__hier0_bF_buf0), .Y(datapath_1_Instr_18_bF_buf20_) );
BUFX2 BUFX2_1081 ( .A(datapath_1_Instr_18__hier0_bF_buf5), .Y(datapath_1_Instr_18_bF_buf19_) );
BUFX2 BUFX2_1082 ( .A(datapath_1_Instr_18__hier0_bF_buf2), .Y(datapath_1_Instr_18_bF_buf18_) );
BUFX2 BUFX2_1083 ( .A(datapath_1_Instr_18__hier0_bF_buf0), .Y(datapath_1_Instr_18_bF_buf17_) );
BUFX2 BUFX2_1084 ( .A(datapath_1_Instr_18__hier0_bF_buf2), .Y(datapath_1_Instr_18_bF_buf16_) );
BUFX2 BUFX2_1085 ( .A(datapath_1_Instr_18__hier0_bF_buf2), .Y(datapath_1_Instr_18_bF_buf15_) );
BUFX2 BUFX2_1086 ( .A(datapath_1_Instr_18__hier0_bF_buf5), .Y(datapath_1_Instr_18_bF_buf14_) );
BUFX2 BUFX2_1087 ( .A(datapath_1_Instr_18__hier0_bF_buf5), .Y(datapath_1_Instr_18_bF_buf13_) );
BUFX2 BUFX2_1088 ( .A(datapath_1_Instr_18__hier0_bF_buf3), .Y(datapath_1_Instr_18_bF_buf12_) );
BUFX2 BUFX2_1089 ( .A(datapath_1_Instr_18__hier0_bF_buf5), .Y(datapath_1_Instr_18_bF_buf11_) );
BUFX2 BUFX2_1090 ( .A(datapath_1_Instr_18__hier0_bF_buf2), .Y(datapath_1_Instr_18_bF_buf10_) );
BUFX2 BUFX2_1091 ( .A(datapath_1_Instr_18__hier0_bF_buf1), .Y(datapath_1_Instr_18_bF_buf9_) );
BUFX2 BUFX2_1092 ( .A(datapath_1_Instr_18__hier0_bF_buf1), .Y(datapath_1_Instr_18_bF_buf8_) );
BUFX2 BUFX2_1093 ( .A(datapath_1_Instr_18__hier0_bF_buf2), .Y(datapath_1_Instr_18_bF_buf7_) );
BUFX2 BUFX2_1094 ( .A(datapath_1_Instr_18__hier0_bF_buf1), .Y(datapath_1_Instr_18_bF_buf6_) );
BUFX2 BUFX2_1095 ( .A(datapath_1_Instr_18__hier0_bF_buf4), .Y(datapath_1_Instr_18_bF_buf5_) );
BUFX2 BUFX2_1096 ( .A(datapath_1_Instr_18__hier0_bF_buf3), .Y(datapath_1_Instr_18_bF_buf4_) );
BUFX2 BUFX2_1097 ( .A(datapath_1_Instr_18__hier0_bF_buf4), .Y(datapath_1_Instr_18_bF_buf3_) );
BUFX2 BUFX2_1098 ( .A(datapath_1_Instr_18__hier0_bF_buf3), .Y(datapath_1_Instr_18_bF_buf2_) );
BUFX2 BUFX2_1099 ( .A(datapath_1_Instr_18__hier0_bF_buf3), .Y(datapath_1_Instr_18_bF_buf1_) );
BUFX2 BUFX2_1100 ( .A(datapath_1_Instr_18__hier0_bF_buf4), .Y(datapath_1_Instr_18_bF_buf0_) );
BUFX2 BUFX2_1101 ( .A(_5746_), .Y(_5746__bF_buf7) );
BUFX2 BUFX2_1102 ( .A(_5746_), .Y(_5746__bF_buf6) );
BUFX2 BUFX2_1103 ( .A(_5746_), .Y(_5746__bF_buf5) );
BUFX2 BUFX2_1104 ( .A(_5746_), .Y(_5746__bF_buf4) );
BUFX2 BUFX2_1105 ( .A(_5746_), .Y(_5746__bF_buf3) );
BUFX2 BUFX2_1106 ( .A(_5746_), .Y(_5746__bF_buf2) );
BUFX2 BUFX2_1107 ( .A(_5746_), .Y(_5746__bF_buf1) );
BUFX2 BUFX2_1108 ( .A(_5746_), .Y(_5746__bF_buf0) );
BUFX2 BUFX2_1109 ( .A(_5326_), .Y(_5326__bF_buf4) );
BUFX2 BUFX2_1110 ( .A(_5326_), .Y(_5326__bF_buf3) );
BUFX2 BUFX2_1111 ( .A(_5326_), .Y(_5326__bF_buf2) );
BUFX2 BUFX2_1112 ( .A(_5326_), .Y(_5326__bF_buf1) );
BUFX2 BUFX2_1113 ( .A(_5326_), .Y(_5326__bF_buf0) );
BUFX2 BUFX2_1114 ( .A(_6149_), .Y(_6149__bF_buf7) );
BUFX2 BUFX2_1115 ( .A(_6149_), .Y(_6149__bF_buf6) );
BUFX2 BUFX2_1116 ( .A(_6149_), .Y(_6149__bF_buf5) );
BUFX2 BUFX2_1117 ( .A(_6149_), .Y(_6149__bF_buf4) );
BUFX2 BUFX2_1118 ( .A(_6149_), .Y(_6149__bF_buf3) );
BUFX2 BUFX2_1119 ( .A(_6149_), .Y(_6149__bF_buf2) );
BUFX2 BUFX2_1120 ( .A(_6149_), .Y(_6149__bF_buf1) );
BUFX2 BUFX2_1121 ( .A(_6149_), .Y(_6149__bF_buf0) );
BUFX2 BUFX2_1122 ( .A(datapath_1_Instr_15_), .Y(datapath_1_Instr_15_bF_buf4_) );
BUFX2 BUFX2_1123 ( .A(datapath_1_Instr_15_), .Y(datapath_1_Instr_15_bF_buf3_) );
BUFX2 BUFX2_1124 ( .A(datapath_1_Instr_15_), .Y(datapath_1_Instr_15_bF_buf2_) );
BUFX2 BUFX2_1125 ( .A(datapath_1_Instr_15_), .Y(datapath_1_Instr_15_bF_buf1_) );
BUFX2 BUFX2_1126 ( .A(datapath_1_Instr_15_), .Y(datapath_1_Instr_15_bF_buf0_) );
BUFX2 BUFX2_1127 ( .A(_248_), .Y(_248__bF_buf3) );
BUFX2 BUFX2_1128 ( .A(_248_), .Y(_248__bF_buf2) );
BUFX2 BUFX2_1129 ( .A(_248_), .Y(_248__bF_buf1) );
BUFX2 BUFX2_1130 ( .A(_248_), .Y(_248__bF_buf0) );
BUFX2 BUFX2_1131 ( .A(_5646_), .Y(_5646__bF_buf7) );
BUFX2 BUFX2_1132 ( .A(_5646_), .Y(_5646__bF_buf6) );
BUFX2 BUFX2_1133 ( .A(_5646_), .Y(_5646__bF_buf5) );
BUFX2 BUFX2_1134 ( .A(_5646_), .Y(_5646__bF_buf4) );
BUFX2 BUFX2_1135 ( .A(_5646_), .Y(_5646__bF_buf3) );
BUFX2 BUFX2_1136 ( .A(_5646_), .Y(_5646__bF_buf2) );
BUFX2 BUFX2_1137 ( .A(_5646_), .Y(_5646__bF_buf1) );
BUFX2 BUFX2_1138 ( .A(_5646_), .Y(_5646__bF_buf0) );
BUFX2 BUFX2_1139 ( .A(IRWrite), .Y(IRWrite_bF_buf4) );
BUFX2 BUFX2_1140 ( .A(IRWrite), .Y(IRWrite_bF_buf3) );
BUFX2 BUFX2_1141 ( .A(IRWrite), .Y(IRWrite_bF_buf2) );
BUFX2 BUFX2_1142 ( .A(IRWrite), .Y(IRWrite_bF_buf1) );
BUFX2 BUFX2_1143 ( .A(IRWrite), .Y(IRWrite_bF_buf0) );
BUFX2 BUFX2_1144 ( .A(_5320_), .Y(_5320__bF_buf4) );
BUFX2 BUFX2_1145 ( .A(_5320_), .Y(_5320__bF_buf3) );
BUFX2 BUFX2_1146 ( .A(_5320_), .Y(_5320__bF_buf2) );
BUFX2 BUFX2_1147 ( .A(_5320_), .Y(_5320__bF_buf1) );
BUFX2 BUFX2_1148 ( .A(_5320_), .Y(_5320__bF_buf0) );
BUFX2 BUFX2_1149 ( .A(_245_), .Y(_245__bF_buf3) );
BUFX2 BUFX2_1150 ( .A(_245_), .Y(_245__bF_buf2) );
BUFX2 BUFX2_1151 ( .A(_245_), .Y(_245__bF_buf1) );
BUFX2 BUFX2_1152 ( .A(_245_), .Y(_245__bF_buf0) );
BUFX2 BUFX2_1153 ( .A(_6046_), .Y(_6046__bF_buf7) );
BUFX2 BUFX2_1154 ( .A(_6046_), .Y(_6046__bF_buf6) );
BUFX2 BUFX2_1155 ( .A(_6046_), .Y(_6046__bF_buf5) );
BUFX2 BUFX2_1156 ( .A(_6046_), .Y(_6046__bF_buf4) );
BUFX2 BUFX2_1157 ( .A(_6046_), .Y(_6046__bF_buf3) );
BUFX2 BUFX2_1158 ( .A(_6046_), .Y(_6046__bF_buf2) );
BUFX2 BUFX2_1159 ( .A(_6046_), .Y(_6046__bF_buf1) );
BUFX2 BUFX2_1160 ( .A(_6046_), .Y(_6046__bF_buf0) );
BUFX2 BUFX2_1161 ( .A(_5296_), .Y(_5296__bF_buf4) );
BUFX2 BUFX2_1162 ( .A(_5296_), .Y(_5296__bF_buf3) );
BUFX2 BUFX2_1163 ( .A(_5296_), .Y(_5296__bF_buf2) );
BUFX2 BUFX2_1164 ( .A(_5296_), .Y(_5296__bF_buf1) );
BUFX2 BUFX2_1165 ( .A(_5296_), .Y(_5296__bF_buf0) );
BUFX2 BUFX2_1166 ( .A(_7116_), .Y(_7116__bF_buf4) );
BUFX2 BUFX2_1167 ( .A(_7116_), .Y(_7116__bF_buf3) );
BUFX2 BUFX2_1168 ( .A(_7116_), .Y(_7116__bF_buf2) );
BUFX2 BUFX2_1169 ( .A(_7116_), .Y(_7116__bF_buf1) );
BUFX2 BUFX2_1170 ( .A(_7116_), .Y(_7116__bF_buf0) );
BUFX2 BUFX2_1171 ( .A(_5411_), .Y(_5411__bF_buf7) );
BUFX2 BUFX2_1172 ( .A(_5411_), .Y(_5411__bF_buf6) );
BUFX2 BUFX2_1173 ( .A(_5411_), .Y(_5411__bF_buf5) );
BUFX2 BUFX2_1174 ( .A(_5411_), .Y(_5411__bF_buf4) );
BUFX2 BUFX2_1175 ( .A(_5411_), .Y(_5411__bF_buf3) );
BUFX2 BUFX2_1176 ( .A(_5411_), .Y(_5411__bF_buf2) );
BUFX2 BUFX2_1177 ( .A(_5411_), .Y(_5411__bF_buf1) );
BUFX2 BUFX2_1178 ( .A(_5411_), .Y(_5411__bF_buf0) );
BUFX2 BUFX2_1179 ( .A(_3588__hier0_bF_buf5), .Y(_3588__bF_buf44) );
BUFX2 BUFX2_1180 ( .A(_3588__hier0_bF_buf4), .Y(_3588__bF_buf43) );
BUFX2 BUFX2_1181 ( .A(_3588__hier0_bF_buf4), .Y(_3588__bF_buf42) );
BUFX2 BUFX2_1182 ( .A(_3588__hier0_bF_buf3), .Y(_3588__bF_buf41) );
BUFX2 BUFX2_1183 ( .A(_3588__hier0_bF_buf4), .Y(_3588__bF_buf40) );
BUFX2 BUFX2_1184 ( .A(_3588__hier0_bF_buf1), .Y(_3588__bF_buf39) );
BUFX2 BUFX2_1185 ( .A(_3588__hier0_bF_buf0), .Y(_3588__bF_buf38) );
BUFX2 BUFX2_1186 ( .A(_3588__hier0_bF_buf3), .Y(_3588__bF_buf37) );
BUFX2 BUFX2_1187 ( .A(_3588__hier0_bF_buf4), .Y(_3588__bF_buf36) );
BUFX2 BUFX2_1188 ( .A(_3588__hier0_bF_buf5), .Y(_3588__bF_buf35) );
BUFX2 BUFX2_1189 ( .A(_3588__hier0_bF_buf2), .Y(_3588__bF_buf34) );
BUFX2 BUFX2_1190 ( .A(_3588__hier0_bF_buf3), .Y(_3588__bF_buf33) );
BUFX2 BUFX2_1191 ( .A(_3588__hier0_bF_buf0), .Y(_3588__bF_buf32) );
BUFX2 BUFX2_1192 ( .A(_3588__hier0_bF_buf1), .Y(_3588__bF_buf31) );
BUFX2 BUFX2_1193 ( .A(_3588__hier0_bF_buf5), .Y(_3588__bF_buf30) );
BUFX2 BUFX2_1194 ( .A(_3588__hier0_bF_buf0), .Y(_3588__bF_buf29) );
BUFX2 BUFX2_1195 ( .A(_3588__hier0_bF_buf2), .Y(_3588__bF_buf28) );
BUFX2 BUFX2_1196 ( .A(_3588__hier0_bF_buf0), .Y(_3588__bF_buf27) );
BUFX2 BUFX2_1197 ( .A(_3588__hier0_bF_buf1), .Y(_3588__bF_buf26) );
BUFX2 BUFX2_1198 ( .A(_3588__hier0_bF_buf4), .Y(_3588__bF_buf25) );
BUFX2 BUFX2_1199 ( .A(_3588__hier0_bF_buf3), .Y(_3588__bF_buf24) );
BUFX2 BUFX2_1200 ( .A(_3588__hier0_bF_buf0), .Y(_3588__bF_buf23) );
BUFX2 BUFX2_1201 ( .A(_3588__hier0_bF_buf2), .Y(_3588__bF_buf22) );
BUFX2 BUFX2_1202 ( .A(_3588__hier0_bF_buf0), .Y(_3588__bF_buf21) );
BUFX2 BUFX2_1203 ( .A(_3588__hier0_bF_buf0), .Y(_3588__bF_buf20) );
BUFX2 BUFX2_1204 ( .A(_3588__hier0_bF_buf1), .Y(_3588__bF_buf19) );
BUFX2 BUFX2_1205 ( .A(_3588__hier0_bF_buf5), .Y(_3588__bF_buf18) );
BUFX2 BUFX2_1206 ( .A(_3588__hier0_bF_buf2), .Y(_3588__bF_buf17) );
BUFX2 BUFX2_1207 ( .A(_3588__hier0_bF_buf3), .Y(_3588__bF_buf16) );
BUFX2 BUFX2_1208 ( .A(_3588__hier0_bF_buf1), .Y(_3588__bF_buf15) );
BUFX2 BUFX2_1209 ( .A(_3588__hier0_bF_buf1), .Y(_3588__bF_buf14) );
BUFX2 BUFX2_1210 ( .A(_3588__hier0_bF_buf1), .Y(_3588__bF_buf13) );
BUFX2 BUFX2_1211 ( .A(_3588__hier0_bF_buf2), .Y(_3588__bF_buf12) );
BUFX2 BUFX2_1212 ( .A(_3588__hier0_bF_buf2), .Y(_3588__bF_buf11) );
BUFX2 BUFX2_1213 ( .A(_3588__hier0_bF_buf5), .Y(_3588__bF_buf10) );
BUFX2 BUFX2_1214 ( .A(_3588__hier0_bF_buf4), .Y(_3588__bF_buf9) );
BUFX2 BUFX2_1215 ( .A(_3588__hier0_bF_buf4), .Y(_3588__bF_buf8) );
BUFX2 BUFX2_1216 ( .A(_3588__hier0_bF_buf5), .Y(_3588__bF_buf7) );
BUFX2 BUFX2_1217 ( .A(_3588__hier0_bF_buf3), .Y(_3588__bF_buf6) );
BUFX2 BUFX2_1218 ( .A(_3588__hier0_bF_buf3), .Y(_3588__bF_buf5) );
BUFX2 BUFX2_1219 ( .A(_3588__hier0_bF_buf5), .Y(_3588__bF_buf4) );
BUFX2 BUFX2_1220 ( .A(_3588__hier0_bF_buf5), .Y(_3588__bF_buf3) );
BUFX2 BUFX2_1221 ( .A(_3588__hier0_bF_buf3), .Y(_3588__bF_buf2) );
BUFX2 BUFX2_1222 ( .A(_3588__hier0_bF_buf4), .Y(_3588__bF_buf1) );
BUFX2 BUFX2_1223 ( .A(_3588__hier0_bF_buf2), .Y(_3588__bF_buf0) );
BUFX2 BUFX2_1224 ( .A(_5314_), .Y(_5314__bF_buf4) );
BUFX2 BUFX2_1225 ( .A(_5314_), .Y(_5314__bF_buf3) );
BUFX2 BUFX2_1226 ( .A(_5314_), .Y(_5314__bF_buf2) );
BUFX2 BUFX2_1227 ( .A(_5314_), .Y(_5314__bF_buf1) );
BUFX2 BUFX2_1228 ( .A(_5314_), .Y(_5314__bF_buf0) );
BUFX2 BUFX2_1229 ( .A(_1883_), .Y(_1883__bF_buf4) );
BUFX2 BUFX2_1230 ( .A(_1883_), .Y(_1883__bF_buf3) );
BUFX2 BUFX2_1231 ( .A(_1883_), .Y(_1883__bF_buf2) );
BUFX2 BUFX2_1232 ( .A(_1883_), .Y(_1883__bF_buf1) );
BUFX2 BUFX2_1233 ( .A(_1883_), .Y(_1883__bF_buf0) );
BUFX2 BUFX2_1234 ( .A(_6786_), .Y(_6786__bF_buf4) );
BUFX2 BUFX2_1235 ( .A(_6786_), .Y(_6786__bF_buf3) );
BUFX2 BUFX2_1236 ( .A(_6786_), .Y(_6786__bF_buf2) );
BUFX2 BUFX2_1237 ( .A(_6786_), .Y(_6786__bF_buf1) );
BUFX2 BUFX2_1238 ( .A(_6786_), .Y(_6786__bF_buf0) );
BUFX2 BUFX2_1239 ( .A(_5446_), .Y(_5446__bF_buf7) );
BUFX2 BUFX2_1240 ( .A(_5446_), .Y(_5446__bF_buf6) );
BUFX2 BUFX2_1241 ( .A(_5446_), .Y(_5446__bF_buf5) );
BUFX2 BUFX2_1242 ( .A(_5446_), .Y(_5446__bF_buf4) );
BUFX2 BUFX2_1243 ( .A(_5446_), .Y(_5446__bF_buf3) );
BUFX2 BUFX2_1244 ( .A(_5446_), .Y(_5446__bF_buf2) );
BUFX2 BUFX2_1245 ( .A(_5446_), .Y(_5446__bF_buf1) );
BUFX2 BUFX2_1246 ( .A(_5446_), .Y(_5446__bF_buf0) );
BUFX2 BUFX2_1247 ( .A(_277_), .Y(_277__bF_buf3) );
BUFX2 BUFX2_1248 ( .A(_277_), .Y(_277__bF_buf2) );
BUFX2 BUFX2_1249 ( .A(_277_), .Y(_277__bF_buf1) );
BUFX2 BUFX2_1250 ( .A(_277_), .Y(_277__bF_buf0) );
BUFX2 BUFX2_1251 ( .A(_5308_), .Y(_5308__bF_buf4) );
BUFX2 BUFX2_1252 ( .A(_5308_), .Y(_5308__bF_buf3) );
BUFX2 BUFX2_1253 ( .A(_5308_), .Y(_5308__bF_buf2) );
BUFX2 BUFX2_1254 ( .A(_5308_), .Y(_5308__bF_buf1) );
BUFX2 BUFX2_1255 ( .A(_5308_), .Y(_5308__bF_buf0) );
BUFX2 BUFX2_1256 ( .A(_5290_), .Y(_5290__bF_buf4) );
BUFX2 BUFX2_1257 ( .A(_5290_), .Y(_5290__bF_buf3) );
BUFX2 BUFX2_1258 ( .A(_5290_), .Y(_5290__bF_buf2) );
BUFX2 BUFX2_1259 ( .A(_5290_), .Y(_5290__bF_buf1) );
BUFX2 BUFX2_1260 ( .A(_5290_), .Y(_5290__bF_buf0) );
BUFX2 BUFX2_1261 ( .A(ALUSrcB_1_), .Y(ALUSrcB_1_bF_buf4_) );
BUFX2 BUFX2_1262 ( .A(ALUSrcB_1_), .Y(ALUSrcB_1_bF_buf3_) );
BUFX2 BUFX2_1263 ( .A(ALUSrcB_1_), .Y(ALUSrcB_1_bF_buf2_) );
BUFX2 BUFX2_1264 ( .A(ALUSrcB_1_), .Y(ALUSrcB_1_bF_buf1_) );
BUFX2 BUFX2_1265 ( .A(ALUSrcB_1_), .Y(ALUSrcB_1_bF_buf0_) );
BUFX2 BUFX2_1266 ( .A(_6551_), .Y(_6551__bF_buf4) );
BUFX2 BUFX2_1267 ( .A(_6551_), .Y(_6551__bF_buf3) );
BUFX2 BUFX2_1268 ( .A(_6551_), .Y(_6551__bF_buf2) );
BUFX2 BUFX2_1269 ( .A(_6551_), .Y(_6551__bF_buf1) );
BUFX2 BUFX2_1270 ( .A(_6551_), .Y(_6551__bF_buf0) );
BUFX2 BUFX2_1271 ( .A(_5284_), .Y(_5284__bF_buf4) );
BUFX2 BUFX2_1272 ( .A(_5284_), .Y(_5284__bF_buf3) );
BUFX2 BUFX2_1273 ( .A(_5284_), .Y(_5284__bF_buf2) );
BUFX2 BUFX2_1274 ( .A(_5284_), .Y(_5284__bF_buf1) );
BUFX2 BUFX2_1275 ( .A(_5284_), .Y(_5284__bF_buf0) );
BUFX2 BUFX2_1276 ( .A(_5913_), .Y(_5913__bF_buf7) );
BUFX2 BUFX2_1277 ( .A(_5913_), .Y(_5913__bF_buf6) );
BUFX2 BUFX2_1278 ( .A(_5913_), .Y(_5913__bF_buf5) );
BUFX2 BUFX2_1279 ( .A(_5913_), .Y(_5913__bF_buf4) );
BUFX2 BUFX2_1280 ( .A(_5913_), .Y(_5913__bF_buf3) );
BUFX2 BUFX2_1281 ( .A(_5913_), .Y(_5913__bF_buf2) );
BUFX2 BUFX2_1282 ( .A(_5913_), .Y(_5913__bF_buf1) );
BUFX2 BUFX2_1283 ( .A(_5913_), .Y(_5913__bF_buf0) );
BUFX2 BUFX2_1284 ( .A(_5302_), .Y(_5302__bF_buf4) );
BUFX2 BUFX2_1285 ( .A(_5302_), .Y(_5302__bF_buf3) );
BUFX2 BUFX2_1286 ( .A(_5302_), .Y(_5302__bF_buf2) );
BUFX2 BUFX2_1287 ( .A(_5302_), .Y(_5302__bF_buf1) );
BUFX2 BUFX2_1288 ( .A(_5302_), .Y(_5302__bF_buf0) );
BUFX2 BUFX2_1289 ( .A(_6316_), .Y(_6316__bF_buf7) );
BUFX2 BUFX2_1290 ( .A(_6316_), .Y(_6316__bF_buf6) );
BUFX2 BUFX2_1291 ( .A(_6316_), .Y(_6316__bF_buf5) );
BUFX2 BUFX2_1292 ( .A(_6316_), .Y(_6316__bF_buf4) );
BUFX2 BUFX2_1293 ( .A(_6316_), .Y(_6316__bF_buf3) );
BUFX2 BUFX2_1294 ( .A(_6316_), .Y(_6316__bF_buf2) );
BUFX2 BUFX2_1295 ( .A(_6316_), .Y(_6316__bF_buf1) );
BUFX2 BUFX2_1296 ( .A(_6316_), .Y(_6316__bF_buf0) );
OAI22X1 OAI22X1_1 ( .A(_3686_), .B(_3685_), .C(datapath_1_Instr_17_bF_buf50_), .D(_3684_), .Y(_3687_) );
INVX1 INVX1_1 ( .A(datapath_1_RegisterFile_regfile_mem_15__2_), .Y(_3688_) );
AOI21X1 AOI21X1_1 ( .A(_3588__bF_buf43), .B(datapath_1_RegisterFile_regfile_mem_14__2_), .C(_3566__bF_buf1), .Y(_3689_) );
OAI21X1 OAI21X1_1 ( .A(_3688_), .B(_3588__bF_buf43), .C(_3689_), .Y(_3690_) );
NAND2X1 NAND2X1_1 ( .A(datapath_1_RegisterFile_regfile_mem_12__2_), .B(_3588__bF_buf1), .Y(_3691_) );
AOI21X1 AOI21X1_2 ( .A(datapath_1_RegisterFile_regfile_mem_13__2_), .B(datapath_1_Instr_16_bF_buf55_), .C(datapath_1_Instr_17_bF_buf49_), .Y(_3692_) );
AOI21X1 AOI21X1_3 ( .A(_3691_), .B(_3692_), .C(_3567__bF_buf4), .Y(_3693_) );
AOI22X1 AOI22X1_1 ( .A(_3690_), .B(_3693_), .C(_3567__bF_buf4), .D(_3687_), .Y(_3694_) );
NOR2X1 NOR2X1_1 ( .A(datapath_1_RegisterFile_regfile_mem_0__2_), .B(datapath_1_Instr_16_bF_buf54_), .Y(_3695_) );
OAI21X1 OAI21X1_2 ( .A(datapath_1_RegisterFile_regfile_mem_1__2_), .B(_3588__bF_buf43), .C(_3566__bF_buf1), .Y(_3696_) );
NOR2X1 NOR2X1_2 ( .A(datapath_1_RegisterFile_regfile_mem_3__2_), .B(_3588__bF_buf43), .Y(_3697_) );
OAI21X1 OAI21X1_3 ( .A(datapath_1_RegisterFile_regfile_mem_2__2_), .B(datapath_1_Instr_16_bF_buf53_), .C(datapath_1_Instr_17_bF_buf48_), .Y(_3698_) );
OAI22X1 OAI22X1_2 ( .A(_3697_), .B(_3698_), .C(_3695_), .D(_3696_), .Y(_3699_) );
NOR2X1 NOR2X1_3 ( .A(datapath_1_Instr_18_bF_buf44_), .B(_3699_), .Y(_3700_) );
MUX2X1 MUX2X1_1 ( .A(datapath_1_RegisterFile_regfile_mem_5__2_), .B(datapath_1_RegisterFile_regfile_mem_4__2_), .S(datapath_1_Instr_16_bF_buf52_), .Y(_3701_) );
NOR2X1 NOR2X1_4 ( .A(datapath_1_RegisterFile_regfile_mem_7__2_), .B(_3588__bF_buf9), .Y(_3702_) );
OAI21X1 OAI21X1_4 ( .A(datapath_1_RegisterFile_regfile_mem_6__2_), .B(datapath_1_Instr_16_bF_buf51_), .C(datapath_1_Instr_17_bF_buf47_), .Y(_3703_) );
OAI22X1 OAI22X1_3 ( .A(_3703_), .B(_3702_), .C(datapath_1_Instr_17_bF_buf46_), .D(_3701_), .Y(_3704_) );
OAI21X1 OAI21X1_5 ( .A(_3567__bF_buf4), .B(_3704_), .C(_3571__bF_buf1), .Y(_3705_) );
OAI22X1 OAI22X1_4 ( .A(_3571__bF_buf1), .B(_3694_), .C(_3700_), .D(_3705_), .Y(_3706_) );
NAND2X1 NAND2X1_2 ( .A(_3570__bF_buf2), .B(_3706_), .Y(_3707_) );
INVX1 INVX1_2 ( .A(datapath_1_RegisterFile_regfile_mem_27__2_), .Y(_3708_) );
AOI21X1 AOI21X1_4 ( .A(datapath_1_RegisterFile_regfile_mem_31__2_), .B(datapath_1_Instr_18_bF_buf43_), .C(_3588__bF_buf31), .Y(_3709_) );
OAI21X1 OAI21X1_6 ( .A(_3708_), .B(datapath_1_Instr_18_bF_buf42_), .C(_3709_), .Y(_3710_) );
INVX1 INVX1_3 ( .A(datapath_1_RegisterFile_regfile_mem_26__2_), .Y(_3711_) );
AOI21X1 AOI21X1_5 ( .A(datapath_1_RegisterFile_regfile_mem_30__2_), .B(datapath_1_Instr_18_bF_buf41_), .C(datapath_1_Instr_16_bF_buf50_), .Y(_3712_) );
OAI21X1 OAI21X1_7 ( .A(_3711_), .B(datapath_1_Instr_18_bF_buf40_), .C(_3712_), .Y(_3713_) );
NAND3X1 NAND3X1_1 ( .A(datapath_1_Instr_17_bF_buf45_), .B(_3713_), .C(_3710_), .Y(_3714_) );
INVX1 INVX1_4 ( .A(datapath_1_RegisterFile_regfile_mem_25__2_), .Y(_3715_) );
AOI21X1 AOI21X1_6 ( .A(datapath_1_RegisterFile_regfile_mem_29__2_), .B(datapath_1_Instr_18_bF_buf39_), .C(_3588__bF_buf31), .Y(_3716_) );
OAI21X1 OAI21X1_8 ( .A(_3715_), .B(datapath_1_Instr_18_bF_buf38_), .C(_3716_), .Y(_3717_) );
INVX1 INVX1_5 ( .A(datapath_1_RegisterFile_regfile_mem_24__2_), .Y(_3718_) );
AOI21X1 AOI21X1_7 ( .A(datapath_1_RegisterFile_regfile_mem_28__2_), .B(datapath_1_Instr_18_bF_buf37_), .C(datapath_1_Instr_16_bF_buf49_), .Y(_3719_) );
OAI21X1 OAI21X1_9 ( .A(_3718_), .B(datapath_1_Instr_18_bF_buf36_), .C(_3719_), .Y(_3720_) );
NAND3X1 NAND3X1_2 ( .A(_3566__bF_buf10), .B(_3720_), .C(_3717_), .Y(_3721_) );
AOI21X1 AOI21X1_8 ( .A(_3714_), .B(_3721_), .C(_3571__bF_buf7), .Y(_3722_) );
MUX2X1 MUX2X1_2 ( .A(datapath_1_RegisterFile_regfile_mem_18__2_), .B(datapath_1_RegisterFile_regfile_mem_16__2_), .S(datapath_1_Instr_17_bF_buf44_), .Y(_3723_) );
NAND2X1 NAND2X1_3 ( .A(_3588__bF_buf15), .B(_3723_), .Y(_3724_) );
MUX2X1 MUX2X1_3 ( .A(datapath_1_RegisterFile_regfile_mem_19__2_), .B(datapath_1_RegisterFile_regfile_mem_17__2_), .S(datapath_1_Instr_17_bF_buf43_), .Y(_3725_) );
NAND2X1 NAND2X1_4 ( .A(datapath_1_Instr_16_bF_buf48_), .B(_3725_), .Y(_3726_) );
NAND3X1 NAND3X1_3 ( .A(_3567__bF_buf0), .B(_3724_), .C(_3726_), .Y(_3727_) );
MUX2X1 MUX2X1_4 ( .A(datapath_1_RegisterFile_regfile_mem_22__2_), .B(datapath_1_RegisterFile_regfile_mem_20__2_), .S(datapath_1_Instr_17_bF_buf42_), .Y(_3728_) );
NAND2X1 NAND2X1_5 ( .A(_3588__bF_buf31), .B(_3728_), .Y(_3729_) );
MUX2X1 MUX2X1_5 ( .A(datapath_1_RegisterFile_regfile_mem_23__2_), .B(datapath_1_RegisterFile_regfile_mem_21__2_), .S(datapath_1_Instr_17_bF_buf41_), .Y(_3730_) );
NAND2X1 NAND2X1_6 ( .A(datapath_1_Instr_16_bF_buf47_), .B(_3730_), .Y(_3731_) );
NAND3X1 NAND3X1_4 ( .A(datapath_1_Instr_18_bF_buf35_), .B(_3729_), .C(_3731_), .Y(_3732_) );
AOI21X1 AOI21X1_9 ( .A(_3727_), .B(_3732_), .C(datapath_1_Instr_19_bF_buf6_), .Y(_3733_) );
OAI21X1 OAI21X1_10 ( .A(_3722_), .B(_3733_), .C(datapath_1_Instr_20_bF_buf5_), .Y(_3734_) );
AOI22X1 AOI22X1_2 ( .A(_3565__bF_buf1), .B(_3569__bF_buf1), .C(_3734_), .D(_3707_), .Y(datapath_1_RD2_2_) );
NAND2X1 NAND2X1_7 ( .A(datapath_1_RegisterFile_regfile_mem_27__3_), .B(datapath_1_Instr_16_bF_buf46_), .Y(_3735_) );
NAND2X1 NAND2X1_8 ( .A(datapath_1_RegisterFile_regfile_mem_26__3_), .B(_3588__bF_buf11), .Y(_3736_) );
NAND3X1 NAND3X1_5 ( .A(datapath_1_Instr_17_bF_buf40_), .B(_3735_), .C(_3736_), .Y(_3737_) );
NAND2X1 NAND2X1_9 ( .A(datapath_1_RegisterFile_regfile_mem_25__3_), .B(datapath_1_Instr_16_bF_buf45_), .Y(_3738_) );
AOI21X1 AOI21X1_10 ( .A(_3588__bF_buf0), .B(datapath_1_RegisterFile_regfile_mem_24__3_), .C(datapath_1_Instr_17_bF_buf39_), .Y(_3739_) );
NAND2X1 NAND2X1_10 ( .A(_3738_), .B(_3739_), .Y(_3740_) );
NAND3X1 NAND3X1_6 ( .A(_3567__bF_buf10), .B(_3737_), .C(_3740_), .Y(_3741_) );
NAND2X1 NAND2X1_11 ( .A(datapath_1_RegisterFile_regfile_mem_31__3_), .B(datapath_1_Instr_16_bF_buf44_), .Y(_3742_) );
AOI21X1 AOI21X1_11 ( .A(_3588__bF_buf14), .B(datapath_1_RegisterFile_regfile_mem_30__3_), .C(_3566__bF_buf9), .Y(_3743_) );
NAND2X1 NAND2X1_12 ( .A(_3742_), .B(_3743_), .Y(_3744_) );
AOI21X1 AOI21X1_12 ( .A(datapath_1_RegisterFile_regfile_mem_29__3_), .B(datapath_1_Instr_16_bF_buf43_), .C(datapath_1_Instr_17_bF_buf38_), .Y(_3745_) );
OAI21X1 OAI21X1_11 ( .A(_2059_), .B(datapath_1_Instr_16_bF_buf42_), .C(_3745_), .Y(_3746_) );
NAND3X1 NAND3X1_7 ( .A(datapath_1_Instr_18_bF_buf34_), .B(_3746_), .C(_3744_), .Y(_3747_) );
AOI21X1 AOI21X1_13 ( .A(_3741_), .B(_3747_), .C(_3571__bF_buf4), .Y(_3748_) );
MUX2X1 MUX2X1_6 ( .A(datapath_1_RegisterFile_regfile_mem_18__3_), .B(datapath_1_RegisterFile_regfile_mem_16__3_), .S(datapath_1_Instr_17_bF_buf37_), .Y(_3749_) );
NAND2X1 NAND2X1_13 ( .A(_3588__bF_buf14), .B(_3749_), .Y(_3750_) );
MUX2X1 MUX2X1_7 ( .A(datapath_1_RegisterFile_regfile_mem_19__3_), .B(datapath_1_RegisterFile_regfile_mem_17__3_), .S(datapath_1_Instr_17_bF_buf36_), .Y(_3751_) );
NAND2X1 NAND2X1_14 ( .A(datapath_1_Instr_16_bF_buf41_), .B(_3751_), .Y(_3752_) );
NAND3X1 NAND3X1_8 ( .A(_3567__bF_buf5), .B(_3750_), .C(_3752_), .Y(_3753_) );
MUX2X1 MUX2X1_8 ( .A(datapath_1_RegisterFile_regfile_mem_22__3_), .B(datapath_1_RegisterFile_regfile_mem_20__3_), .S(datapath_1_Instr_17_bF_buf35_), .Y(_3754_) );
NAND2X1 NAND2X1_15 ( .A(_3588__bF_buf14), .B(_3754_), .Y(_3755_) );
MUX2X1 MUX2X1_9 ( .A(datapath_1_RegisterFile_regfile_mem_23__3_), .B(datapath_1_RegisterFile_regfile_mem_21__3_), .S(datapath_1_Instr_17_bF_buf34_), .Y(_3756_) );
NAND2X1 NAND2X1_16 ( .A(datapath_1_Instr_16_bF_buf40_), .B(_3756_), .Y(_3757_) );
NAND3X1 NAND3X1_9 ( .A(datapath_1_Instr_18_bF_buf33_), .B(_3755_), .C(_3757_), .Y(_3758_) );
AOI21X1 AOI21X1_14 ( .A(_3753_), .B(_3758_), .C(datapath_1_Instr_19_bF_buf5_), .Y(_3759_) );
OAI21X1 OAI21X1_12 ( .A(_3759_), .B(_3748_), .C(datapath_1_Instr_20_bF_buf4_), .Y(_3760_) );
INVX1 INVX1_6 ( .A(datapath_1_RegisterFile_regfile_mem_9__3_), .Y(_3761_) );
AOI21X1 AOI21X1_15 ( .A(datapath_1_RegisterFile_regfile_mem_13__3_), .B(datapath_1_Instr_18_bF_buf32_), .C(_3588__bF_buf36), .Y(_3762_) );
OAI21X1 OAI21X1_13 ( .A(_3761_), .B(datapath_1_Instr_18_bF_buf31_), .C(_3762_), .Y(_3763_) );
INVX1 INVX1_7 ( .A(datapath_1_RegisterFile_regfile_mem_8__3_), .Y(_3764_) );
AOI21X1 AOI21X1_16 ( .A(datapath_1_RegisterFile_regfile_mem_12__3_), .B(datapath_1_Instr_18_bF_buf30_), .C(datapath_1_Instr_16_bF_buf39_), .Y(_3765_) );
OAI21X1 OAI21X1_14 ( .A(_3764_), .B(datapath_1_Instr_18_bF_buf29_), .C(_3765_), .Y(_3766_) );
NAND3X1 NAND3X1_10 ( .A(_3566__bF_buf1), .B(_3766_), .C(_3763_), .Y(_3767_) );
INVX1 INVX1_8 ( .A(datapath_1_RegisterFile_regfile_mem_11__3_), .Y(_3768_) );
AOI21X1 AOI21X1_17 ( .A(datapath_1_RegisterFile_regfile_mem_15__3_), .B(datapath_1_Instr_18_bF_buf28_), .C(_3588__bF_buf43), .Y(_3769_) );
OAI21X1 OAI21X1_15 ( .A(_3768_), .B(datapath_1_Instr_18_bF_buf27_), .C(_3769_), .Y(_3770_) );
INVX1 INVX1_9 ( .A(datapath_1_RegisterFile_regfile_mem_10__3_), .Y(_3771_) );
AOI21X1 AOI21X1_18 ( .A(datapath_1_RegisterFile_regfile_mem_14__3_), .B(datapath_1_Instr_18_bF_buf26_), .C(datapath_1_Instr_16_bF_buf38_), .Y(_3772_) );
OAI21X1 OAI21X1_16 ( .A(_3771_), .B(datapath_1_Instr_18_bF_buf25_), .C(_3772_), .Y(_3773_) );
NAND3X1 NAND3X1_11 ( .A(datapath_1_Instr_17_bF_buf33_), .B(_3773_), .C(_3770_), .Y(_3774_) );
AOI21X1 AOI21X1_19 ( .A(_3767_), .B(_3774_), .C(_3571__bF_buf1), .Y(_3775_) );
MUX2X1 MUX2X1_10 ( .A(datapath_1_RegisterFile_regfile_mem_1__3_), .B(datapath_1_RegisterFile_regfile_mem_0__3_), .S(datapath_1_Instr_16_bF_buf37_), .Y(_3776_) );
NOR2X1 NOR2X1_5 ( .A(datapath_1_RegisterFile_regfile_mem_3__3_), .B(_3588__bF_buf9), .Y(_3777_) );
OAI21X1 OAI21X1_17 ( .A(datapath_1_RegisterFile_regfile_mem_2__3_), .B(datapath_1_Instr_16_bF_buf36_), .C(datapath_1_Instr_17_bF_buf32_), .Y(_3778_) );
OAI22X1 OAI22X1_5 ( .A(_3778_), .B(_3777_), .C(datapath_1_Instr_17_bF_buf31_), .D(_3776_), .Y(_3779_) );
NAND2X1 NAND2X1_17 ( .A(_3567__bF_buf4), .B(_3779_), .Y(_3780_) );
MUX2X1 MUX2X1_11 ( .A(datapath_1_RegisterFile_regfile_mem_5__3_), .B(datapath_1_RegisterFile_regfile_mem_4__3_), .S(datapath_1_Instr_16_bF_buf35_), .Y(_3781_) );
NOR2X1 NOR2X1_6 ( .A(datapath_1_RegisterFile_regfile_mem_7__3_), .B(_3588__bF_buf42), .Y(_3782_) );
OAI21X1 OAI21X1_18 ( .A(datapath_1_RegisterFile_regfile_mem_6__3_), .B(datapath_1_Instr_16_bF_buf34_), .C(datapath_1_Instr_17_bF_buf30_), .Y(_3783_) );
OAI22X1 OAI22X1_6 ( .A(_3783_), .B(_3782_), .C(datapath_1_Instr_17_bF_buf29_), .D(_3781_), .Y(_3784_) );
NAND2X1 NAND2X1_18 ( .A(datapath_1_Instr_18_bF_buf24_), .B(_3784_), .Y(_3785_) );
AOI21X1 AOI21X1_20 ( .A(_3780_), .B(_3785_), .C(datapath_1_Instr_19_bF_buf4_), .Y(_3786_) );
OAI21X1 OAI21X1_19 ( .A(_3775_), .B(_3786_), .C(_3570__bF_buf2), .Y(_3787_) );
AOI22X1 AOI22X1_3 ( .A(_3565__bF_buf1), .B(_3569__bF_buf1), .C(_3760_), .D(_3787_), .Y(datapath_1_RD2_3_) );
NAND2X1 NAND2X1_19 ( .A(datapath_1_RegisterFile_regfile_mem_27__4_), .B(datapath_1_Instr_16_bF_buf33_), .Y(_3788_) );
NAND2X1 NAND2X1_20 ( .A(datapath_1_RegisterFile_regfile_mem_26__4_), .B(_3588__bF_buf24), .Y(_3789_) );
NAND3X1 NAND3X1_12 ( .A(datapath_1_Instr_17_bF_buf28_), .B(_3788_), .C(_3789_), .Y(_3790_) );
NAND2X1 NAND2X1_21 ( .A(datapath_1_RegisterFile_regfile_mem_25__4_), .B(datapath_1_Instr_16_bF_buf32_), .Y(_3791_) );
AOI21X1 AOI21X1_21 ( .A(_3588__bF_buf2), .B(datapath_1_RegisterFile_regfile_mem_24__4_), .C(datapath_1_Instr_17_bF_buf27_), .Y(_3792_) );
NAND2X1 NAND2X1_22 ( .A(_3791_), .B(_3792_), .Y(_3793_) );
NAND3X1 NAND3X1_13 ( .A(_3567__bF_buf2), .B(_3790_), .C(_3793_), .Y(_3794_) );
NAND2X1 NAND2X1_23 ( .A(datapath_1_RegisterFile_regfile_mem_31__4_), .B(datapath_1_Instr_16_bF_buf31_), .Y(_3795_) );
AOI21X1 AOI21X1_22 ( .A(_3588__bF_buf24), .B(datapath_1_RegisterFile_regfile_mem_30__4_), .C(_3566__bF_buf10), .Y(_3796_) );
NAND2X1 NAND2X1_24 ( .A(_3795_), .B(_3796_), .Y(_3797_) );
INVX1 INVX1_10 ( .A(datapath_1_RegisterFile_regfile_mem_28__4_), .Y(_3798_) );
AOI21X1 AOI21X1_23 ( .A(datapath_1_RegisterFile_regfile_mem_29__4_), .B(datapath_1_Instr_16_bF_buf30_), .C(datapath_1_Instr_17_bF_buf26_), .Y(_3799_) );
OAI21X1 OAI21X1_20 ( .A(_3798_), .B(datapath_1_Instr_16_bF_buf29_), .C(_3799_), .Y(_3800_) );
NAND3X1 NAND3X1_14 ( .A(datapath_1_Instr_18_bF_buf23_), .B(_3800_), .C(_3797_), .Y(_3801_) );
AOI21X1 AOI21X1_24 ( .A(_3794_), .B(_3801_), .C(_3571__bF_buf7), .Y(_3802_) );
MUX2X1 MUX2X1_12 ( .A(datapath_1_RegisterFile_regfile_mem_17__4_), .B(datapath_1_RegisterFile_regfile_mem_16__4_), .S(datapath_1_Instr_16_bF_buf28_), .Y(_3803_) );
NOR2X1 NOR2X1_7 ( .A(datapath_1_RegisterFile_regfile_mem_19__4_), .B(_3588__bF_buf16), .Y(_3804_) );
OAI21X1 OAI21X1_21 ( .A(datapath_1_RegisterFile_regfile_mem_18__4_), .B(datapath_1_Instr_16_bF_buf27_), .C(datapath_1_Instr_17_bF_buf25_), .Y(_3805_) );
OAI22X1 OAI22X1_7 ( .A(_3805_), .B(_3804_), .C(datapath_1_Instr_17_bF_buf24_), .D(_3803_), .Y(_3806_) );
NAND2X1 NAND2X1_25 ( .A(_3567__bF_buf3), .B(_3806_), .Y(_3807_) );
MUX2X1 MUX2X1_13 ( .A(datapath_1_RegisterFile_regfile_mem_21__4_), .B(datapath_1_RegisterFile_regfile_mem_20__4_), .S(datapath_1_Instr_16_bF_buf26_), .Y(_3808_) );
NOR2X1 NOR2X1_8 ( .A(datapath_1_RegisterFile_regfile_mem_23__4_), .B(_3588__bF_buf16), .Y(_3809_) );
OAI21X1 OAI21X1_22 ( .A(datapath_1_RegisterFile_regfile_mem_22__4_), .B(datapath_1_Instr_16_bF_buf25_), .C(datapath_1_Instr_17_bF_buf23_), .Y(_3810_) );
OAI22X1 OAI22X1_8 ( .A(_3810_), .B(_3809_), .C(datapath_1_Instr_17_bF_buf22_), .D(_3808_), .Y(_3811_) );
NAND2X1 NAND2X1_26 ( .A(datapath_1_Instr_18_bF_buf22_), .B(_3811_), .Y(_3812_) );
AOI21X1 AOI21X1_25 ( .A(_3807_), .B(_3812_), .C(datapath_1_Instr_19_bF_buf3_), .Y(_3813_) );
OAI21X1 OAI21X1_23 ( .A(_3802_), .B(_3813_), .C(datapath_1_Instr_20_bF_buf3_), .Y(_3814_) );
NAND2X1 NAND2X1_27 ( .A(datapath_1_RegisterFile_regfile_mem_11__4_), .B(datapath_1_Instr_17_bF_buf21_), .Y(_3815_) );
NAND2X1 NAND2X1_28 ( .A(datapath_1_RegisterFile_regfile_mem_9__4_), .B(_3566__bF_buf8), .Y(_3816_) );
NAND3X1 NAND3X1_15 ( .A(datapath_1_Instr_16_bF_buf24_), .B(_3815_), .C(_3816_), .Y(_3817_) );
NAND2X1 NAND2X1_29 ( .A(datapath_1_RegisterFile_regfile_mem_10__4_), .B(datapath_1_Instr_17_bF_buf20_), .Y(_3818_) );
AOI21X1 AOI21X1_26 ( .A(_3566__bF_buf7), .B(datapath_1_RegisterFile_regfile_mem_8__4_), .C(datapath_1_Instr_16_bF_buf23_), .Y(_3819_) );
NAND2X1 NAND2X1_30 ( .A(_3818_), .B(_3819_), .Y(_3820_) );
NAND3X1 NAND3X1_16 ( .A(_3567__bF_buf8), .B(_3817_), .C(_3820_), .Y(_3821_) );
NAND2X1 NAND2X1_31 ( .A(datapath_1_RegisterFile_regfile_mem_15__4_), .B(datapath_1_Instr_17_bF_buf19_), .Y(_3822_) );
NAND2X1 NAND2X1_32 ( .A(datapath_1_RegisterFile_regfile_mem_13__4_), .B(_3566__bF_buf8), .Y(_3823_) );
NAND3X1 NAND3X1_17 ( .A(datapath_1_Instr_16_bF_buf22_), .B(_3822_), .C(_3823_), .Y(_3824_) );
NAND2X1 NAND2X1_33 ( .A(datapath_1_RegisterFile_regfile_mem_14__4_), .B(datapath_1_Instr_17_bF_buf18_), .Y(_3825_) );
AOI21X1 AOI21X1_27 ( .A(_3566__bF_buf8), .B(datapath_1_RegisterFile_regfile_mem_12__4_), .C(datapath_1_Instr_16_bF_buf21_), .Y(_3826_) );
NAND2X1 NAND2X1_34 ( .A(_3825_), .B(_3826_), .Y(_3827_) );
NAND3X1 NAND3X1_18 ( .A(datapath_1_Instr_18_bF_buf21_), .B(_3824_), .C(_3827_), .Y(_3828_) );
AOI21X1 AOI21X1_28 ( .A(_3821_), .B(_3828_), .C(_3571__bF_buf3), .Y(_3829_) );
INVX1 INVX1_11 ( .A(datapath_1_RegisterFile_regfile_mem_1__4_), .Y(_3830_) );
AOI21X1 AOI21X1_29 ( .A(datapath_1_RegisterFile_regfile_mem_5__4_), .B(datapath_1_Instr_18_bF_buf20_), .C(_3588__bF_buf25), .Y(_3831_) );
OAI21X1 OAI21X1_24 ( .A(_3830_), .B(datapath_1_Instr_18_bF_buf19_), .C(_3831_), .Y(_3832_) );
INVX1 INVX1_12 ( .A(datapath_1_RegisterFile_regfile_mem_0__4_), .Y(_3833_) );
AOI21X1 AOI21X1_30 ( .A(datapath_1_RegisterFile_regfile_mem_4__4_), .B(datapath_1_Instr_18_bF_buf18_), .C(datapath_1_Instr_16_bF_buf20_), .Y(_3834_) );
OAI21X1 OAI21X1_25 ( .A(_3833_), .B(datapath_1_Instr_18_bF_buf17_), .C(_3834_), .Y(_3835_) );
NAND3X1 NAND3X1_19 ( .A(_3566__bF_buf7), .B(_3835_), .C(_3832_), .Y(_3836_) );
INVX1 INVX1_13 ( .A(datapath_1_RegisterFile_regfile_mem_3__4_), .Y(_3837_) );
AOI21X1 AOI21X1_31 ( .A(datapath_1_RegisterFile_regfile_mem_7__4_), .B(datapath_1_Instr_18_bF_buf16_), .C(_3588__bF_buf18), .Y(_3838_) );
OAI21X1 OAI21X1_26 ( .A(_3837_), .B(datapath_1_Instr_18_bF_buf15_), .C(_3838_), .Y(_3839_) );
INVX1 INVX1_14 ( .A(datapath_1_RegisterFile_regfile_mem_2__4_), .Y(_3840_) );
AOI21X1 AOI21X1_32 ( .A(datapath_1_RegisterFile_regfile_mem_6__4_), .B(datapath_1_Instr_18_bF_buf14_), .C(datapath_1_Instr_16_bF_buf19_), .Y(_3841_) );
OAI21X1 OAI21X1_27 ( .A(_3840_), .B(datapath_1_Instr_18_bF_buf13_), .C(_3841_), .Y(_3842_) );
NAND3X1 NAND3X1_20 ( .A(datapath_1_Instr_17_bF_buf17_), .B(_3842_), .C(_3839_), .Y(_3843_) );
AOI21X1 AOI21X1_33 ( .A(_3836_), .B(_3843_), .C(datapath_1_Instr_19_bF_buf2_), .Y(_3844_) );
OAI21X1 OAI21X1_28 ( .A(_3844_), .B(_3829_), .C(_3570__bF_buf3), .Y(_3845_) );
AOI22X1 AOI22X1_4 ( .A(_3565__bF_buf4), .B(_3569__bF_buf4), .C(_3845_), .D(_3814_), .Y(datapath_1_RD2_4_) );
NAND2X1 NAND2X1_35 ( .A(datapath_1_RegisterFile_regfile_mem_27__5_), .B(datapath_1_Instr_16_bF_buf18_), .Y(_3846_) );
NAND2X1 NAND2X1_36 ( .A(datapath_1_RegisterFile_regfile_mem_26__5_), .B(_3588__bF_buf23), .Y(_3847_) );
NAND3X1 NAND3X1_21 ( .A(datapath_1_Instr_17_bF_buf16_), .B(_3846_), .C(_3847_), .Y(_3848_) );
NAND2X1 NAND2X1_37 ( .A(datapath_1_RegisterFile_regfile_mem_25__5_), .B(datapath_1_Instr_16_bF_buf17_), .Y(_3849_) );
AOI21X1 AOI21X1_34 ( .A(_3588__bF_buf23), .B(datapath_1_RegisterFile_regfile_mem_24__5_), .C(datapath_1_Instr_17_bF_buf15_), .Y(_3850_) );
NAND2X1 NAND2X1_38 ( .A(_3849_), .B(_3850_), .Y(_3851_) );
NAND3X1 NAND3X1_22 ( .A(_3567__bF_buf9), .B(_3848_), .C(_3851_), .Y(_3852_) );
NAND2X1 NAND2X1_39 ( .A(datapath_1_RegisterFile_regfile_mem_31__5_), .B(datapath_1_Instr_16_bF_buf16_), .Y(_3853_) );
AOI21X1 AOI21X1_35 ( .A(_3588__bF_buf38), .B(datapath_1_RegisterFile_regfile_mem_30__5_), .C(_3566__bF_buf6), .Y(_3854_) );
NAND2X1 NAND2X1_40 ( .A(_3853_), .B(_3854_), .Y(_3855_) );
INVX1 INVX1_15 ( .A(datapath_1_RegisterFile_regfile_mem_28__5_), .Y(_3856_) );
AOI21X1 AOI21X1_36 ( .A(datapath_1_RegisterFile_regfile_mem_29__5_), .B(datapath_1_Instr_16_bF_buf15_), .C(datapath_1_Instr_17_bF_buf14_), .Y(_3857_) );
OAI21X1 OAI21X1_29 ( .A(_3856_), .B(datapath_1_Instr_16_bF_buf14_), .C(_3857_), .Y(_3858_) );
NAND3X1 NAND3X1_23 ( .A(datapath_1_Instr_18_bF_buf12_), .B(_3858_), .C(_3855_), .Y(_3859_) );
AOI21X1 AOI21X1_37 ( .A(_3852_), .B(_3859_), .C(_3571__bF_buf5), .Y(_3860_) );
MUX2X1 MUX2X1_14 ( .A(datapath_1_RegisterFile_regfile_mem_18__5_), .B(datapath_1_RegisterFile_regfile_mem_16__5_), .S(datapath_1_Instr_17_bF_buf13_), .Y(_3861_) );
NAND2X1 NAND2X1_41 ( .A(_3588__bF_buf27), .B(_3861_), .Y(_3862_) );
MUX2X1 MUX2X1_15 ( .A(datapath_1_RegisterFile_regfile_mem_19__5_), .B(datapath_1_RegisterFile_regfile_mem_17__5_), .S(datapath_1_Instr_17_bF_buf12_), .Y(_3863_) );
NAND2X1 NAND2X1_42 ( .A(datapath_1_Instr_16_bF_buf13_), .B(_3863_), .Y(_3864_) );
NAND3X1 NAND3X1_24 ( .A(_3567__bF_buf9), .B(_3862_), .C(_3864_), .Y(_3865_) );
MUX2X1 MUX2X1_16 ( .A(datapath_1_RegisterFile_regfile_mem_22__5_), .B(datapath_1_RegisterFile_regfile_mem_20__5_), .S(datapath_1_Instr_17_bF_buf11_), .Y(_3866_) );
NAND2X1 NAND2X1_43 ( .A(_3588__bF_buf27), .B(_3866_), .Y(_3867_) );
MUX2X1 MUX2X1_17 ( .A(datapath_1_RegisterFile_regfile_mem_23__5_), .B(datapath_1_RegisterFile_regfile_mem_21__5_), .S(datapath_1_Instr_17_bF_buf10_), .Y(_3868_) );
NAND2X1 NAND2X1_44 ( .A(datapath_1_Instr_16_bF_buf12_), .B(_3868_), .Y(_3869_) );
NAND3X1 NAND3X1_25 ( .A(datapath_1_Instr_18_bF_buf11_), .B(_3867_), .C(_3869_), .Y(_3870_) );
AOI21X1 AOI21X1_38 ( .A(_3865_), .B(_3870_), .C(datapath_1_Instr_19_bF_buf1_), .Y(_3871_) );
OAI21X1 OAI21X1_30 ( .A(_3871_), .B(_3860_), .C(datapath_1_Instr_20_bF_buf2_), .Y(_3872_) );
MUX2X1 MUX2X1_18 ( .A(datapath_1_RegisterFile_regfile_mem_9__5_), .B(datapath_1_RegisterFile_regfile_mem_8__5_), .S(datapath_1_Instr_16_bF_buf11_), .Y(_3873_) );
NOR2X1 NOR2X1_9 ( .A(datapath_1_RegisterFile_regfile_mem_11__5_), .B(_3588__bF_buf10), .Y(_3874_) );
OAI21X1 OAI21X1_31 ( .A(datapath_1_RegisterFile_regfile_mem_10__5_), .B(datapath_1_Instr_16_bF_buf10_), .C(datapath_1_Instr_17_bF_buf9_), .Y(_3875_) );
OAI22X1 OAI22X1_9 ( .A(_3875_), .B(_3874_), .C(datapath_1_Instr_17_bF_buf8_), .D(_3873_), .Y(_3876_) );
AOI21X1 AOI21X1_39 ( .A(_3588__bF_buf10), .B(datapath_1_RegisterFile_regfile_mem_14__5_), .C(_3566__bF_buf3), .Y(_3877_) );
OAI21X1 OAI21X1_32 ( .A(_2162_), .B(_3588__bF_buf10), .C(_3877_), .Y(_3878_) );
NAND2X1 NAND2X1_45 ( .A(datapath_1_RegisterFile_regfile_mem_12__5_), .B(_3588__bF_buf10), .Y(_3879_) );
AOI21X1 AOI21X1_40 ( .A(datapath_1_RegisterFile_regfile_mem_13__5_), .B(datapath_1_Instr_16_bF_buf9_), .C(datapath_1_Instr_17_bF_buf7_), .Y(_3880_) );
AOI21X1 AOI21X1_41 ( .A(_3879_), .B(_3880_), .C(_3567__bF_buf6), .Y(_3881_) );
AOI22X1 AOI22X1_5 ( .A(_3878_), .B(_3881_), .C(_3567__bF_buf6), .D(_3876_), .Y(_3882_) );
NOR2X1 NOR2X1_10 ( .A(datapath_1_RegisterFile_regfile_mem_0__5_), .B(datapath_1_Instr_16_bF_buf8_), .Y(_3883_) );
OAI21X1 OAI21X1_33 ( .A(datapath_1_RegisterFile_regfile_mem_1__5_), .B(_3588__bF_buf44), .C(_3566__bF_buf6), .Y(_3884_) );
NOR2X1 NOR2X1_11 ( .A(datapath_1_RegisterFile_regfile_mem_3__5_), .B(_3588__bF_buf44), .Y(_3885_) );
OAI21X1 OAI21X1_34 ( .A(datapath_1_RegisterFile_regfile_mem_2__5_), .B(datapath_1_Instr_16_bF_buf7_), .C(datapath_1_Instr_17_bF_buf6_), .Y(_3886_) );
OAI22X1 OAI22X1_10 ( .A(_3885_), .B(_3886_), .C(_3883_), .D(_3884_), .Y(_3887_) );
NOR2X1 NOR2X1_12 ( .A(datapath_1_Instr_18_bF_buf10_), .B(_3887_), .Y(_3888_) );
MUX2X1 MUX2X1_19 ( .A(datapath_1_RegisterFile_regfile_mem_5__5_), .B(datapath_1_RegisterFile_regfile_mem_4__5_), .S(datapath_1_Instr_16_bF_buf6_), .Y(_3889_) );
NOR2X1 NOR2X1_13 ( .A(datapath_1_RegisterFile_regfile_mem_7__5_), .B(_3588__bF_buf4), .Y(_3890_) );
OAI21X1 OAI21X1_35 ( .A(datapath_1_RegisterFile_regfile_mem_6__5_), .B(datapath_1_Instr_16_bF_buf5_), .C(datapath_1_Instr_17_bF_buf5_), .Y(_3891_) );
OAI22X1 OAI22X1_11 ( .A(_3891_), .B(_3890_), .C(datapath_1_Instr_17_bF_buf4_), .D(_3889_), .Y(_3892_) );
OAI21X1 OAI21X1_36 ( .A(_3567__bF_buf1), .B(_3892_), .C(_3571__bF_buf6), .Y(_3893_) );
OAI22X1 OAI22X1_12 ( .A(_3571__bF_buf6), .B(_3882_), .C(_3888_), .D(_3893_), .Y(_3894_) );
NAND2X1 NAND2X1_46 ( .A(_3570__bF_buf4), .B(_3894_), .Y(_3895_) );
AOI22X1 AOI22X1_6 ( .A(_3565__bF_buf3), .B(_3569__bF_buf3), .C(_3872_), .D(_3895_), .Y(datapath_1_RD2_5_) );
MUX2X1 MUX2X1_20 ( .A(datapath_1_RegisterFile_regfile_mem_9__6_), .B(datapath_1_RegisterFile_regfile_mem_8__6_), .S(datapath_1_Instr_16_bF_buf4_), .Y(_3896_) );
NOR2X1 NOR2X1_14 ( .A(datapath_1_RegisterFile_regfile_mem_11__6_), .B(_3588__bF_buf25), .Y(_3897_) );
OAI21X1 OAI21X1_37 ( .A(datapath_1_RegisterFile_regfile_mem_10__6_), .B(datapath_1_Instr_16_bF_buf3_), .C(datapath_1_Instr_17_bF_buf3_), .Y(_3898_) );
OAI22X1 OAI22X1_13 ( .A(_3898_), .B(_3897_), .C(datapath_1_Instr_17_bF_buf2_), .D(_3896_), .Y(_3899_) );
INVX1 INVX1_16 ( .A(datapath_1_RegisterFile_regfile_mem_15__6_), .Y(_3900_) );
AOI21X1 AOI21X1_42 ( .A(_3588__bF_buf1), .B(datapath_1_RegisterFile_regfile_mem_14__6_), .C(_3566__bF_buf0), .Y(_3901_) );
OAI21X1 OAI21X1_38 ( .A(_3900_), .B(_3588__bF_buf1), .C(_3901_), .Y(_3902_) );
NAND2X1 NAND2X1_47 ( .A(datapath_1_RegisterFile_regfile_mem_12__6_), .B(_3588__bF_buf1), .Y(_3903_) );
AOI21X1 AOI21X1_43 ( .A(datapath_1_RegisterFile_regfile_mem_13__6_), .B(datapath_1_Instr_16_bF_buf2_), .C(datapath_1_Instr_17_bF_buf1_), .Y(_3904_) );
AOI21X1 AOI21X1_44 ( .A(_3903_), .B(_3904_), .C(_3567__bF_buf4), .Y(_3905_) );
AOI22X1 AOI22X1_7 ( .A(_3902_), .B(_3905_), .C(_3567__bF_buf8), .D(_3899_), .Y(_3906_) );
NOR2X1 NOR2X1_15 ( .A(datapath_1_RegisterFile_regfile_mem_0__6_), .B(datapath_1_Instr_16_bF_buf1_), .Y(_3907_) );
OAI21X1 OAI21X1_39 ( .A(datapath_1_RegisterFile_regfile_mem_1__6_), .B(_3588__bF_buf25), .C(_3566__bF_buf7), .Y(_3908_) );
NOR2X1 NOR2X1_16 ( .A(datapath_1_RegisterFile_regfile_mem_3__6_), .B(_3588__bF_buf25), .Y(_3909_) );
OAI21X1 OAI21X1_40 ( .A(datapath_1_RegisterFile_regfile_mem_2__6_), .B(datapath_1_Instr_16_bF_buf0_), .C(datapath_1_Instr_17_bF_buf0_), .Y(_3910_) );
OAI22X1 OAI22X1_14 ( .A(_3909_), .B(_3910_), .C(_3907_), .D(_3908_), .Y(_3911_) );
NOR2X1 NOR2X1_17 ( .A(datapath_1_Instr_18_bF_buf9_), .B(_3911_), .Y(_3912_) );
MUX2X1 MUX2X1_21 ( .A(datapath_1_RegisterFile_regfile_mem_5__6_), .B(datapath_1_RegisterFile_regfile_mem_4__6_), .S(datapath_1_Instr_16_bF_buf55_), .Y(_3913_) );
NOR2X1 NOR2X1_18 ( .A(datapath_1_RegisterFile_regfile_mem_7__6_), .B(_3588__bF_buf25), .Y(_3914_) );
OAI21X1 OAI21X1_41 ( .A(datapath_1_RegisterFile_regfile_mem_6__6_), .B(datapath_1_Instr_16_bF_buf54_), .C(datapath_1_Instr_17_bF_buf50_), .Y(_3915_) );
OAI22X1 OAI22X1_15 ( .A(_3915_), .B(_3914_), .C(datapath_1_Instr_17_bF_buf49_), .D(_3913_), .Y(_3916_) );
OAI21X1 OAI21X1_42 ( .A(_3567__bF_buf4), .B(_3916_), .C(_3571__bF_buf1), .Y(_3917_) );
OAI22X1 OAI22X1_16 ( .A(_3571__bF_buf3), .B(_3906_), .C(_3912_), .D(_3917_), .Y(_3918_) );
NAND2X1 NAND2X1_48 ( .A(_3570__bF_buf3), .B(_3918_), .Y(_3919_) );
INVX1 INVX1_17 ( .A(datapath_1_RegisterFile_regfile_mem_27__6_), .Y(_3920_) );
AOI21X1 AOI21X1_45 ( .A(datapath_1_RegisterFile_regfile_mem_31__6_), .B(datapath_1_Instr_18_bF_buf8_), .C(_3588__bF_buf5), .Y(_3921_) );
OAI21X1 OAI21X1_43 ( .A(_3920_), .B(datapath_1_Instr_18_bF_buf7_), .C(_3921_), .Y(_3922_) );
INVX1 INVX1_18 ( .A(datapath_1_RegisterFile_regfile_mem_26__6_), .Y(_3923_) );
AOI21X1 AOI21X1_46 ( .A(datapath_1_RegisterFile_regfile_mem_30__6_), .B(datapath_1_Instr_18_bF_buf6_), .C(datapath_1_Instr_16_bF_buf53_), .Y(_3924_) );
OAI21X1 OAI21X1_44 ( .A(_3923_), .B(datapath_1_Instr_18_bF_buf5_), .C(_3924_), .Y(_3925_) );
NAND3X1 NAND3X1_26 ( .A(datapath_1_Instr_17_bF_buf48_), .B(_3925_), .C(_3922_), .Y(_3926_) );
INVX1 INVX1_19 ( .A(datapath_1_RegisterFile_regfile_mem_25__6_), .Y(_3927_) );
AOI21X1 AOI21X1_47 ( .A(datapath_1_RegisterFile_regfile_mem_29__6_), .B(datapath_1_Instr_18_bF_buf4_), .C(_3588__bF_buf37), .Y(_3928_) );
OAI21X1 OAI21X1_45 ( .A(_3927_), .B(datapath_1_Instr_18_bF_buf3_), .C(_3928_), .Y(_3929_) );
INVX1 INVX1_20 ( .A(datapath_1_RegisterFile_regfile_mem_24__6_), .Y(_3930_) );
AOI21X1 AOI21X1_48 ( .A(datapath_1_RegisterFile_regfile_mem_28__6_), .B(datapath_1_Instr_18_bF_buf2_), .C(datapath_1_Instr_16_bF_buf52_), .Y(_3931_) );
OAI21X1 OAI21X1_46 ( .A(_3930_), .B(datapath_1_Instr_18_bF_buf1_), .C(_3931_), .Y(_3932_) );
NAND3X1 NAND3X1_27 ( .A(_3566__bF_buf4), .B(_3932_), .C(_3929_), .Y(_3933_) );
AOI21X1 AOI21X1_49 ( .A(_3926_), .B(_3933_), .C(_3571__bF_buf7), .Y(_3934_) );
MUX2X1 MUX2X1_22 ( .A(datapath_1_RegisterFile_regfile_mem_18__6_), .B(datapath_1_RegisterFile_regfile_mem_16__6_), .S(datapath_1_Instr_17_bF_buf47_), .Y(_3935_) );
NAND2X1 NAND2X1_49 ( .A(_3588__bF_buf2), .B(_3935_), .Y(_3936_) );
MUX2X1 MUX2X1_23 ( .A(datapath_1_RegisterFile_regfile_mem_19__6_), .B(datapath_1_RegisterFile_regfile_mem_17__6_), .S(datapath_1_Instr_17_bF_buf46_), .Y(_3937_) );
NAND2X1 NAND2X1_50 ( .A(datapath_1_Instr_16_bF_buf51_), .B(_3937_), .Y(_3938_) );
NAND3X1 NAND3X1_28 ( .A(_3567__bF_buf2), .B(_3936_), .C(_3938_), .Y(_3939_) );
MUX2X1 MUX2X1_24 ( .A(datapath_1_RegisterFile_regfile_mem_22__6_), .B(datapath_1_RegisterFile_regfile_mem_20__6_), .S(datapath_1_Instr_17_bF_buf45_), .Y(_3940_) );
NAND2X1 NAND2X1_51 ( .A(_3588__bF_buf33), .B(_3940_), .Y(_3941_) );
MUX2X1 MUX2X1_25 ( .A(datapath_1_RegisterFile_regfile_mem_23__6_), .B(datapath_1_RegisterFile_regfile_mem_21__6_), .S(datapath_1_Instr_17_bF_buf44_), .Y(_3942_) );
NAND2X1 NAND2X1_52 ( .A(datapath_1_Instr_16_bF_buf50_), .B(_3942_), .Y(_3943_) );
NAND3X1 NAND3X1_29 ( .A(datapath_1_Instr_18_bF_buf0_), .B(_3941_), .C(_3943_), .Y(_3944_) );
AOI21X1 AOI21X1_50 ( .A(_3939_), .B(_3944_), .C(datapath_1_Instr_19_bF_buf0_), .Y(_3945_) );
OAI21X1 OAI21X1_47 ( .A(_3934_), .B(_3945_), .C(datapath_1_Instr_20_bF_buf1_), .Y(_3946_) );
AOI22X1 AOI22X1_8 ( .A(_3565__bF_buf4), .B(_3569__bF_buf4), .C(_3946_), .D(_3919_), .Y(datapath_1_RD2_6_) );
MUX2X1 MUX2X1_26 ( .A(datapath_1_RegisterFile_regfile_mem_9__7_), .B(datapath_1_RegisterFile_regfile_mem_8__7_), .S(datapath_1_Instr_16_bF_buf49_), .Y(_3947_) );
NOR2X1 NOR2X1_19 ( .A(datapath_1_RegisterFile_regfile_mem_11__7_), .B(_3588__bF_buf22), .Y(_3948_) );
OAI21X1 OAI21X1_48 ( .A(datapath_1_RegisterFile_regfile_mem_10__7_), .B(datapath_1_Instr_16_bF_buf48_), .C(datapath_1_Instr_17_bF_buf43_), .Y(_3949_) );
OAI22X1 OAI22X1_17 ( .A(_3949_), .B(_3948_), .C(datapath_1_Instr_17_bF_buf42_), .D(_3947_), .Y(_3950_) );
AOI21X1 AOI21X1_51 ( .A(_3588__bF_buf22), .B(datapath_1_RegisterFile_regfile_mem_14__7_), .C(_3566__bF_buf2), .Y(_3951_) );
OAI21X1 OAI21X1_49 ( .A(_2297_), .B(_3588__bF_buf22), .C(_3951_), .Y(_3952_) );
NAND2X1 NAND2X1_53 ( .A(datapath_1_RegisterFile_regfile_mem_12__7_), .B(_3588__bF_buf17), .Y(_3953_) );
AOI21X1 AOI21X1_52 ( .A(datapath_1_RegisterFile_regfile_mem_13__7_), .B(datapath_1_Instr_16_bF_buf47_), .C(datapath_1_Instr_17_bF_buf41_), .Y(_3954_) );
AOI21X1 AOI21X1_53 ( .A(_3953_), .B(_3954_), .C(_3567__bF_buf7), .Y(_3955_) );
AOI22X1 AOI22X1_9 ( .A(_3952_), .B(_3955_), .C(_3567__bF_buf7), .D(_3950_), .Y(_3956_) );
NOR2X1 NOR2X1_20 ( .A(datapath_1_RegisterFile_regfile_mem_0__7_), .B(datapath_1_Instr_16_bF_buf46_), .Y(_3957_) );
OAI21X1 OAI21X1_50 ( .A(datapath_1_RegisterFile_regfile_mem_1__7_), .B(_3588__bF_buf34), .C(_3566__bF_buf2), .Y(_3958_) );
NOR2X1 NOR2X1_21 ( .A(datapath_1_RegisterFile_regfile_mem_3__7_), .B(_3588__bF_buf34), .Y(_3959_) );
OAI21X1 OAI21X1_51 ( .A(datapath_1_RegisterFile_regfile_mem_2__7_), .B(datapath_1_Instr_16_bF_buf45_), .C(datapath_1_Instr_17_bF_buf40_), .Y(_3960_) );
OAI22X1 OAI22X1_18 ( .A(_3959_), .B(_3960_), .C(_3957_), .D(_3958_), .Y(_3961_) );
NOR2X1 NOR2X1_22 ( .A(datapath_1_Instr_18_bF_buf44_), .B(_3961_), .Y(_3962_) );
MUX2X1 MUX2X1_27 ( .A(datapath_1_RegisterFile_regfile_mem_5__7_), .B(datapath_1_RegisterFile_regfile_mem_4__7_), .S(datapath_1_Instr_16_bF_buf44_), .Y(_3963_) );
NOR2X1 NOR2X1_23 ( .A(datapath_1_RegisterFile_regfile_mem_7__7_), .B(_3588__bF_buf17), .Y(_3964_) );
OAI21X1 OAI21X1_52 ( .A(datapath_1_RegisterFile_regfile_mem_6__7_), .B(datapath_1_Instr_16_bF_buf43_), .C(datapath_1_Instr_17_bF_buf39_), .Y(_3965_) );
OAI22X1 OAI22X1_19 ( .A(_3965_), .B(_3964_), .C(datapath_1_Instr_17_bF_buf38_), .D(_3963_), .Y(_3966_) );
OAI21X1 OAI21X1_53 ( .A(_3567__bF_buf10), .B(_3966_), .C(_3571__bF_buf0), .Y(_3967_) );
OAI22X1 OAI22X1_20 ( .A(_3571__bF_buf0), .B(_3956_), .C(_3962_), .D(_3967_), .Y(_3968_) );
NAND2X1 NAND2X1_54 ( .A(_3570__bF_buf1), .B(_3968_), .Y(_3969_) );
INVX1 INVX1_21 ( .A(datapath_1_RegisterFile_regfile_mem_19__7_), .Y(_3970_) );
AOI21X1 AOI21X1_54 ( .A(datapath_1_RegisterFile_regfile_mem_23__7_), .B(datapath_1_Instr_18_bF_buf43_), .C(_3588__bF_buf26), .Y(_3971_) );
OAI21X1 OAI21X1_54 ( .A(_3970_), .B(datapath_1_Instr_18_bF_buf42_), .C(_3971_), .Y(_3972_) );
NAND2X1 NAND2X1_55 ( .A(datapath_1_RegisterFile_regfile_mem_18__7_), .B(_3567__bF_buf5), .Y(_3973_) );
AOI21X1 AOI21X1_55 ( .A(datapath_1_RegisterFile_regfile_mem_22__7_), .B(datapath_1_Instr_18_bF_buf41_), .C(datapath_1_Instr_16_bF_buf42_), .Y(_3974_) );
AOI21X1 AOI21X1_56 ( .A(_3973_), .B(_3974_), .C(_3566__bF_buf9), .Y(_3975_) );
INVX1 INVX1_22 ( .A(datapath_1_RegisterFile_regfile_mem_17__7_), .Y(_3976_) );
AOI21X1 AOI21X1_57 ( .A(datapath_1_RegisterFile_regfile_mem_21__7_), .B(datapath_1_Instr_18_bF_buf40_), .C(_3588__bF_buf26), .Y(_3977_) );
OAI21X1 OAI21X1_55 ( .A(_3976_), .B(datapath_1_Instr_18_bF_buf39_), .C(_3977_), .Y(_3978_) );
NAND2X1 NAND2X1_56 ( .A(datapath_1_RegisterFile_regfile_mem_16__7_), .B(_3567__bF_buf5), .Y(_3979_) );
AOI21X1 AOI21X1_58 ( .A(datapath_1_RegisterFile_regfile_mem_20__7_), .B(datapath_1_Instr_18_bF_buf38_), .C(datapath_1_Instr_16_bF_buf41_), .Y(_3980_) );
AOI21X1 AOI21X1_59 ( .A(_3979_), .B(_3980_), .C(datapath_1_Instr_17_bF_buf37_), .Y(_3981_) );
AOI22X1 AOI22X1_10 ( .A(_3975_), .B(_3972_), .C(_3978_), .D(_3981_), .Y(_3982_) );
NOR2X1 NOR2X1_24 ( .A(datapath_1_RegisterFile_regfile_mem_24__7_), .B(datapath_1_Instr_16_bF_buf40_), .Y(_3983_) );
OAI21X1 OAI21X1_56 ( .A(datapath_1_RegisterFile_regfile_mem_25__7_), .B(_3588__bF_buf0), .C(_3566__bF_buf9), .Y(_3984_) );
NOR2X1 NOR2X1_25 ( .A(datapath_1_RegisterFile_regfile_mem_27__7_), .B(_3588__bF_buf0), .Y(_3985_) );
OAI21X1 OAI21X1_57 ( .A(datapath_1_RegisterFile_regfile_mem_26__7_), .B(datapath_1_Instr_16_bF_buf39_), .C(datapath_1_Instr_17_bF_buf36_), .Y(_3986_) );
OAI22X1 OAI22X1_21 ( .A(_3985_), .B(_3986_), .C(_3983_), .D(_3984_), .Y(_3987_) );
NOR2X1 NOR2X1_26 ( .A(datapath_1_Instr_18_bF_buf37_), .B(_3987_), .Y(_3988_) );
MUX2X1 MUX2X1_28 ( .A(datapath_1_RegisterFile_regfile_mem_29__7_), .B(datapath_1_RegisterFile_regfile_mem_28__7_), .S(datapath_1_Instr_16_bF_buf38_), .Y(_3989_) );
NOR2X1 NOR2X1_27 ( .A(datapath_1_RegisterFile_regfile_mem_31__7_), .B(_3588__bF_buf11), .Y(_3990_) );
OAI21X1 OAI21X1_58 ( .A(datapath_1_RegisterFile_regfile_mem_30__7_), .B(datapath_1_Instr_16_bF_buf37_), .C(datapath_1_Instr_17_bF_buf35_), .Y(_3991_) );
OAI22X1 OAI22X1_22 ( .A(_3991_), .B(_3990_), .C(datapath_1_Instr_17_bF_buf34_), .D(_3989_), .Y(_3992_) );
OAI21X1 OAI21X1_59 ( .A(_3567__bF_buf5), .B(_3992_), .C(datapath_1_Instr_19_bF_buf6_), .Y(_3993_) );
OAI22X1 OAI22X1_23 ( .A(datapath_1_Instr_19_bF_buf5_), .B(_3982_), .C(_3988_), .D(_3993_), .Y(_3994_) );
NAND2X1 NAND2X1_57 ( .A(datapath_1_Instr_20_bF_buf0_), .B(_3994_), .Y(_3995_) );
AOI22X1 AOI22X1_11 ( .A(_3565__bF_buf1), .B(_3569__bF_buf1), .C(_3995_), .D(_3969_), .Y(datapath_1_RD2_7_) );
NAND2X1 NAND2X1_58 ( .A(datapath_1_RegisterFile_regfile_mem_27__8_), .B(datapath_1_Instr_16_bF_buf36_), .Y(_3996_) );
NAND2X1 NAND2X1_59 ( .A(datapath_1_RegisterFile_regfile_mem_26__8_), .B(_3588__bF_buf2), .Y(_3997_) );
NAND3X1 NAND3X1_30 ( .A(datapath_1_Instr_17_bF_buf33_), .B(_3996_), .C(_3997_), .Y(_3998_) );
NAND2X1 NAND2X1_60 ( .A(datapath_1_RegisterFile_regfile_mem_25__8_), .B(datapath_1_Instr_16_bF_buf35_), .Y(_3999_) );
AOI21X1 AOI21X1_60 ( .A(_3588__bF_buf2), .B(datapath_1_RegisterFile_regfile_mem_24__8_), .C(datapath_1_Instr_17_bF_buf32_), .Y(_4000_) );
NAND2X1 NAND2X1_61 ( .A(_3999_), .B(_4000_), .Y(_4001_) );
NAND3X1 NAND3X1_31 ( .A(_3567__bF_buf2), .B(_3998_), .C(_4001_), .Y(_4002_) );
NAND2X1 NAND2X1_62 ( .A(datapath_1_RegisterFile_regfile_mem_31__8_), .B(datapath_1_Instr_16_bF_buf34_), .Y(_4003_) );
AOI21X1 AOI21X1_61 ( .A(_3588__bF_buf24), .B(datapath_1_RegisterFile_regfile_mem_30__8_), .C(_3566__bF_buf10), .Y(_4004_) );
NAND2X1 NAND2X1_63 ( .A(_4003_), .B(_4004_), .Y(_4005_) );
INVX1 INVX1_23 ( .A(datapath_1_RegisterFile_regfile_mem_28__8_), .Y(_4006_) );
AOI21X1 AOI21X1_62 ( .A(datapath_1_RegisterFile_regfile_mem_29__8_), .B(datapath_1_Instr_16_bF_buf33_), .C(datapath_1_Instr_17_bF_buf31_), .Y(_4007_) );
OAI21X1 OAI21X1_60 ( .A(_4006_), .B(datapath_1_Instr_16_bF_buf32_), .C(_4007_), .Y(_4008_) );
NAND3X1 NAND3X1_32 ( .A(datapath_1_Instr_18_bF_buf36_), .B(_4008_), .C(_4005_), .Y(_4009_) );
AOI21X1 AOI21X1_63 ( .A(_4002_), .B(_4009_), .C(_3571__bF_buf7), .Y(_4010_) );
MUX2X1 MUX2X1_29 ( .A(datapath_1_RegisterFile_regfile_mem_18__8_), .B(datapath_1_RegisterFile_regfile_mem_16__8_), .S(datapath_1_Instr_17_bF_buf30_), .Y(_4011_) );
NAND2X1 NAND2X1_64 ( .A(_3588__bF_buf2), .B(_4011_), .Y(_4012_) );
MUX2X1 MUX2X1_30 ( .A(datapath_1_RegisterFile_regfile_mem_19__8_), .B(datapath_1_RegisterFile_regfile_mem_17__8_), .S(datapath_1_Instr_17_bF_buf29_), .Y(_4013_) );
NAND2X1 NAND2X1_65 ( .A(datapath_1_Instr_16_bF_buf31_), .B(_4013_), .Y(_4014_) );
NAND3X1 NAND3X1_33 ( .A(_3567__bF_buf2), .B(_4012_), .C(_4014_), .Y(_4015_) );
MUX2X1 MUX2X1_31 ( .A(datapath_1_RegisterFile_regfile_mem_22__8_), .B(datapath_1_RegisterFile_regfile_mem_20__8_), .S(datapath_1_Instr_17_bF_buf28_), .Y(_4016_) );
NAND2X1 NAND2X1_66 ( .A(_3588__bF_buf24), .B(_4016_), .Y(_4017_) );
MUX2X1 MUX2X1_32 ( .A(datapath_1_RegisterFile_regfile_mem_23__8_), .B(datapath_1_RegisterFile_regfile_mem_21__8_), .S(datapath_1_Instr_17_bF_buf27_), .Y(_4018_) );
NAND2X1 NAND2X1_67 ( .A(datapath_1_Instr_16_bF_buf30_), .B(_4018_), .Y(_4019_) );
NAND3X1 NAND3X1_34 ( .A(datapath_1_Instr_18_bF_buf35_), .B(_4017_), .C(_4019_), .Y(_4020_) );
AOI21X1 AOI21X1_64 ( .A(_4015_), .B(_4020_), .C(datapath_1_Instr_19_bF_buf4_), .Y(_4021_) );
OAI21X1 OAI21X1_61 ( .A(_4021_), .B(_4010_), .C(datapath_1_Instr_20_bF_buf5_), .Y(_4022_) );
MUX2X1 MUX2X1_33 ( .A(datapath_1_RegisterFile_regfile_mem_9__8_), .B(datapath_1_RegisterFile_regfile_mem_8__8_), .S(datapath_1_Instr_16_bF_buf29_), .Y(_4023_) );
NOR2X1 NOR2X1_28 ( .A(datapath_1_RegisterFile_regfile_mem_11__8_), .B(_3588__bF_buf8), .Y(_4024_) );
OAI21X1 OAI21X1_62 ( .A(datapath_1_RegisterFile_regfile_mem_10__8_), .B(datapath_1_Instr_16_bF_buf28_), .C(datapath_1_Instr_17_bF_buf26_), .Y(_4025_) );
OAI22X1 OAI22X1_24 ( .A(_4025_), .B(_4024_), .C(datapath_1_Instr_17_bF_buf25_), .D(_4023_), .Y(_4026_) );
AOI21X1 AOI21X1_65 ( .A(_3588__bF_buf8), .B(datapath_1_RegisterFile_regfile_mem_14__8_), .C(_3566__bF_buf0), .Y(_4027_) );
OAI21X1 OAI21X1_63 ( .A(_2321_), .B(_3588__bF_buf8), .C(_4027_), .Y(_4028_) );
NAND2X1 NAND2X1_68 ( .A(datapath_1_RegisterFile_regfile_mem_12__8_), .B(_3588__bF_buf8), .Y(_4029_) );
AOI21X1 AOI21X1_66 ( .A(datapath_1_RegisterFile_regfile_mem_13__8_), .B(datapath_1_Instr_16_bF_buf27_), .C(datapath_1_Instr_17_bF_buf24_), .Y(_4030_) );
AOI21X1 AOI21X1_67 ( .A(_4029_), .B(_4030_), .C(_3567__bF_buf8), .Y(_4031_) );
AOI22X1 AOI22X1_12 ( .A(_4028_), .B(_4031_), .C(_3567__bF_buf8), .D(_4026_), .Y(_4032_) );
NOR2X1 NOR2X1_29 ( .A(datapath_1_RegisterFile_regfile_mem_0__8_), .B(datapath_1_Instr_16_bF_buf26_), .Y(_4033_) );
OAI21X1 OAI21X1_64 ( .A(datapath_1_RegisterFile_regfile_mem_1__8_), .B(_3588__bF_buf25), .C(_3566__bF_buf7), .Y(_4034_) );
NOR2X1 NOR2X1_30 ( .A(datapath_1_RegisterFile_regfile_mem_3__8_), .B(_3588__bF_buf9), .Y(_4035_) );
OAI21X1 OAI21X1_65 ( .A(datapath_1_RegisterFile_regfile_mem_2__8_), .B(datapath_1_Instr_16_bF_buf25_), .C(datapath_1_Instr_17_bF_buf23_), .Y(_4036_) );
OAI22X1 OAI22X1_25 ( .A(_4035_), .B(_4036_), .C(_4033_), .D(_4034_), .Y(_4037_) );
NOR2X1 NOR2X1_31 ( .A(datapath_1_Instr_18_bF_buf34_), .B(_4037_), .Y(_4038_) );
MUX2X1 MUX2X1_34 ( .A(datapath_1_RegisterFile_regfile_mem_5__8_), .B(datapath_1_RegisterFile_regfile_mem_4__8_), .S(datapath_1_Instr_16_bF_buf24_), .Y(_4039_) );
NOR2X1 NOR2X1_32 ( .A(datapath_1_RegisterFile_regfile_mem_7__8_), .B(_3588__bF_buf25), .Y(_4040_) );
OAI21X1 OAI21X1_66 ( .A(datapath_1_RegisterFile_regfile_mem_6__8_), .B(datapath_1_Instr_16_bF_buf23_), .C(datapath_1_Instr_17_bF_buf22_), .Y(_4041_) );
OAI22X1 OAI22X1_26 ( .A(_4041_), .B(_4040_), .C(datapath_1_Instr_17_bF_buf21_), .D(_4039_), .Y(_4042_) );
OAI21X1 OAI21X1_67 ( .A(_3567__bF_buf8), .B(_4042_), .C(_3571__bF_buf3), .Y(_4043_) );
OAI22X1 OAI22X1_27 ( .A(_3571__bF_buf3), .B(_4032_), .C(_4038_), .D(_4043_), .Y(_4044_) );
NAND2X1 NAND2X1_69 ( .A(_3570__bF_buf3), .B(_4044_), .Y(_4045_) );
AOI22X1 AOI22X1_13 ( .A(_3565__bF_buf4), .B(_3569__bF_buf4), .C(_4022_), .D(_4045_), .Y(datapath_1_RD2_8_) );
NAND2X1 NAND2X1_70 ( .A(datapath_1_RegisterFile_regfile_mem_27__9_), .B(datapath_1_Instr_16_bF_buf22_), .Y(_4046_) );
NAND2X1 NAND2X1_71 ( .A(datapath_1_RegisterFile_regfile_mem_26__9_), .B(_3588__bF_buf21), .Y(_4047_) );
NAND3X1 NAND3X1_35 ( .A(datapath_1_Instr_17_bF_buf20_), .B(_4046_), .C(_4047_), .Y(_4048_) );
NAND2X1 NAND2X1_72 ( .A(datapath_1_RegisterFile_regfile_mem_25__9_), .B(datapath_1_Instr_16_bF_buf21_), .Y(_4049_) );
AOI21X1 AOI21X1_68 ( .A(_3588__bF_buf21), .B(datapath_1_RegisterFile_regfile_mem_24__9_), .C(datapath_1_Instr_17_bF_buf19_), .Y(_4050_) );
NAND2X1 NAND2X1_73 ( .A(_4049_), .B(_4050_), .Y(_4051_) );
NAND3X1 NAND3X1_36 ( .A(_3567__bF_buf3), .B(_4048_), .C(_4051_), .Y(_4052_) );
NAND2X1 NAND2X1_74 ( .A(datapath_1_RegisterFile_regfile_mem_31__9_), .B(datapath_1_Instr_16_bF_buf20_), .Y(_4053_) );
AOI21X1 AOI21X1_69 ( .A(_3588__bF_buf21), .B(datapath_1_RegisterFile_regfile_mem_30__9_), .C(_3566__bF_buf4), .Y(_4054_) );
NAND2X1 NAND2X1_75 ( .A(_4053_), .B(_4054_), .Y(_4055_) );
INVX1 INVX1_24 ( .A(datapath_1_RegisterFile_regfile_mem_28__9_), .Y(_4056_) );
AOI21X1 AOI21X1_70 ( .A(datapath_1_RegisterFile_regfile_mem_29__9_), .B(datapath_1_Instr_16_bF_buf19_), .C(datapath_1_Instr_17_bF_buf18_), .Y(_4057_) );
OAI21X1 OAI21X1_68 ( .A(_4056_), .B(datapath_1_Instr_16_bF_buf18_), .C(_4057_), .Y(_4058_) );
NAND3X1 NAND3X1_37 ( .A(datapath_1_Instr_18_bF_buf33_), .B(_4058_), .C(_4055_), .Y(_4059_) );
AOI21X1 AOI21X1_71 ( .A(_4052_), .B(_4059_), .C(_3571__bF_buf5), .Y(_4060_) );
MUX2X1 MUX2X1_35 ( .A(datapath_1_RegisterFile_regfile_mem_17__9_), .B(datapath_1_RegisterFile_regfile_mem_16__9_), .S(datapath_1_Instr_16_bF_buf17_), .Y(_4061_) );
NOR2X1 NOR2X1_33 ( .A(datapath_1_RegisterFile_regfile_mem_19__9_), .B(_3588__bF_buf32), .Y(_4062_) );
OAI21X1 OAI21X1_69 ( .A(datapath_1_RegisterFile_regfile_mem_18__9_), .B(datapath_1_Instr_16_bF_buf16_), .C(datapath_1_Instr_17_bF_buf17_), .Y(_4063_) );
OAI22X1 OAI22X1_28 ( .A(_4063_), .B(_4062_), .C(datapath_1_Instr_17_bF_buf16_), .D(_4061_), .Y(_4064_) );
NAND2X1 NAND2X1_76 ( .A(_3567__bF_buf9), .B(_4064_), .Y(_4065_) );
MUX2X1 MUX2X1_36 ( .A(datapath_1_RegisterFile_regfile_mem_21__9_), .B(datapath_1_RegisterFile_regfile_mem_20__9_), .S(datapath_1_Instr_16_bF_buf15_), .Y(_4066_) );
NOR2X1 NOR2X1_34 ( .A(datapath_1_RegisterFile_regfile_mem_23__9_), .B(_3588__bF_buf23), .Y(_4067_) );
OAI21X1 OAI21X1_70 ( .A(datapath_1_RegisterFile_regfile_mem_22__9_), .B(datapath_1_Instr_16_bF_buf14_), .C(datapath_1_Instr_17_bF_buf15_), .Y(_4068_) );
OAI22X1 OAI22X1_29 ( .A(_4068_), .B(_4067_), .C(datapath_1_Instr_17_bF_buf14_), .D(_4066_), .Y(_4069_) );
NAND2X1 NAND2X1_77 ( .A(datapath_1_Instr_18_bF_buf32_), .B(_4069_), .Y(_4070_) );
AOI21X1 AOI21X1_72 ( .A(_4065_), .B(_4070_), .C(datapath_1_Instr_19_bF_buf3_), .Y(_4071_) );
OAI21X1 OAI21X1_71 ( .A(_4060_), .B(_4071_), .C(datapath_1_Instr_20_bF_buf4_), .Y(_4072_) );
NAND2X1 NAND2X1_78 ( .A(datapath_1_RegisterFile_regfile_mem_11__9_), .B(datapath_1_Instr_17_bF_buf13_), .Y(_4073_) );
NAND2X1 NAND2X1_79 ( .A(datapath_1_RegisterFile_regfile_mem_9__9_), .B(_3566__bF_buf3), .Y(_4074_) );
NAND3X1 NAND3X1_38 ( .A(datapath_1_Instr_16_bF_buf13_), .B(_4073_), .C(_4074_), .Y(_4075_) );
NAND2X1 NAND2X1_80 ( .A(datapath_1_RegisterFile_regfile_mem_10__9_), .B(datapath_1_Instr_17_bF_buf12_), .Y(_4076_) );
AOI21X1 AOI21X1_73 ( .A(_3566__bF_buf3), .B(datapath_1_RegisterFile_regfile_mem_8__9_), .C(datapath_1_Instr_16_bF_buf12_), .Y(_4077_) );
NAND2X1 NAND2X1_81 ( .A(_4076_), .B(_4077_), .Y(_4078_) );
NAND3X1 NAND3X1_39 ( .A(_3567__bF_buf6), .B(_4075_), .C(_4078_), .Y(_4079_) );
NAND2X1 NAND2X1_82 ( .A(datapath_1_RegisterFile_regfile_mem_15__9_), .B(datapath_1_Instr_17_bF_buf11_), .Y(_4080_) );
NAND2X1 NAND2X1_83 ( .A(datapath_1_RegisterFile_regfile_mem_13__9_), .B(_3566__bF_buf8), .Y(_4081_) );
NAND3X1 NAND3X1_40 ( .A(datapath_1_Instr_16_bF_buf11_), .B(_4080_), .C(_4081_), .Y(_4082_) );
NAND2X1 NAND2X1_84 ( .A(datapath_1_RegisterFile_regfile_mem_14__9_), .B(datapath_1_Instr_17_bF_buf10_), .Y(_4083_) );
AOI21X1 AOI21X1_74 ( .A(_3566__bF_buf3), .B(datapath_1_RegisterFile_regfile_mem_12__9_), .C(datapath_1_Instr_16_bF_buf10_), .Y(_4084_) );
NAND2X1 NAND2X1_85 ( .A(_4083_), .B(_4084_), .Y(_4085_) );
NAND3X1 NAND3X1_41 ( .A(datapath_1_Instr_18_bF_buf31_), .B(_4082_), .C(_4085_), .Y(_4086_) );
AOI21X1 AOI21X1_75 ( .A(_4079_), .B(_4086_), .C(_3571__bF_buf6), .Y(_4087_) );
AOI21X1 AOI21X1_76 ( .A(datapath_1_RegisterFile_regfile_mem_5__9_), .B(datapath_1_Instr_18_bF_buf30_), .C(_3588__bF_buf18), .Y(_4088_) );
OAI21X1 OAI21X1_72 ( .A(_2367_), .B(datapath_1_Instr_18_bF_buf29_), .C(_4088_), .Y(_4089_) );
AOI21X1 AOI21X1_77 ( .A(datapath_1_RegisterFile_regfile_mem_4__9_), .B(datapath_1_Instr_18_bF_buf28_), .C(datapath_1_Instr_16_bF_buf9_), .Y(_4090_) );
OAI21X1 OAI21X1_73 ( .A(_2370_), .B(datapath_1_Instr_18_bF_buf27_), .C(_4090_), .Y(_4091_) );
NAND3X1 NAND3X1_42 ( .A(_3566__bF_buf8), .B(_4091_), .C(_4089_), .Y(_4092_) );
AOI21X1 AOI21X1_78 ( .A(datapath_1_RegisterFile_regfile_mem_7__9_), .B(datapath_1_Instr_18_bF_buf26_), .C(_3588__bF_buf18), .Y(_4093_) );
OAI21X1 OAI21X1_74 ( .A(_2374_), .B(datapath_1_Instr_18_bF_buf25_), .C(_4093_), .Y(_4094_) );
AOI21X1 AOI21X1_79 ( .A(datapath_1_RegisterFile_regfile_mem_6__9_), .B(datapath_1_Instr_18_bF_buf24_), .C(datapath_1_Instr_16_bF_buf8_), .Y(_4095_) );
OAI21X1 OAI21X1_75 ( .A(_2377_), .B(datapath_1_Instr_18_bF_buf23_), .C(_4095_), .Y(_4096_) );
NAND3X1 NAND3X1_43 ( .A(datapath_1_Instr_17_bF_buf9_), .B(_4096_), .C(_4094_), .Y(_4097_) );
AOI21X1 AOI21X1_80 ( .A(_4092_), .B(_4097_), .C(datapath_1_Instr_19_bF_buf2_), .Y(_4098_) );
OAI21X1 OAI21X1_76 ( .A(_4098_), .B(_4087_), .C(_3570__bF_buf0), .Y(_4099_) );
AOI22X1 AOI22X1_14 ( .A(_3565__bF_buf3), .B(_3569__bF_buf3), .C(_4099_), .D(_4072_), .Y(datapath_1_RD2_9_) );
NAND2X1 NAND2X1_86 ( .A(datapath_1_RegisterFile_regfile_mem_27__10_), .B(datapath_1_Instr_16_bF_buf7_), .Y(_4100_) );
NAND2X1 NAND2X1_87 ( .A(datapath_1_RegisterFile_regfile_mem_26__10_), .B(_3588__bF_buf21), .Y(_4101_) );
NAND3X1 NAND3X1_44 ( .A(datapath_1_Instr_17_bF_buf8_), .B(_4100_), .C(_4101_), .Y(_4102_) );
NAND2X1 NAND2X1_88 ( .A(datapath_1_RegisterFile_regfile_mem_25__10_), .B(datapath_1_Instr_16_bF_buf6_), .Y(_4103_) );
AOI21X1 AOI21X1_81 ( .A(_3588__bF_buf21), .B(datapath_1_RegisterFile_regfile_mem_24__10_), .C(datapath_1_Instr_17_bF_buf7_), .Y(_4104_) );
NAND2X1 NAND2X1_89 ( .A(_4103_), .B(_4104_), .Y(_4105_) );
NAND3X1 NAND3X1_45 ( .A(_3567__bF_buf1), .B(_4102_), .C(_4105_), .Y(_4106_) );
NAND2X1 NAND2X1_90 ( .A(datapath_1_RegisterFile_regfile_mem_31__10_), .B(datapath_1_Instr_16_bF_buf5_), .Y(_4107_) );
AOI21X1 AOI21X1_82 ( .A(_3588__bF_buf20), .B(datapath_1_RegisterFile_regfile_mem_30__10_), .C(_3566__bF_buf6), .Y(_4108_) );
NAND2X1 NAND2X1_91 ( .A(_4107_), .B(_4108_), .Y(_4109_) );
AOI21X1 AOI21X1_83 ( .A(datapath_1_RegisterFile_regfile_mem_29__10_), .B(datapath_1_Instr_16_bF_buf4_), .C(datapath_1_Instr_17_bF_buf6_), .Y(_4110_) );
OAI21X1 OAI21X1_77 ( .A(_2435_), .B(datapath_1_Instr_16_bF_buf3_), .C(_4110_), .Y(_4111_) );
NAND3X1 NAND3X1_46 ( .A(datapath_1_Instr_18_bF_buf22_), .B(_4111_), .C(_4109_), .Y(_4112_) );
AOI21X1 AOI21X1_84 ( .A(_4106_), .B(_4112_), .C(_3571__bF_buf5), .Y(_4113_) );
MUX2X1 MUX2X1_37 ( .A(datapath_1_RegisterFile_regfile_mem_17__10_), .B(datapath_1_RegisterFile_regfile_mem_16__10_), .S(datapath_1_Instr_16_bF_buf2_), .Y(_4114_) );
NOR2X1 NOR2X1_35 ( .A(datapath_1_RegisterFile_regfile_mem_19__10_), .B(_3588__bF_buf27), .Y(_4115_) );
OAI21X1 OAI21X1_78 ( .A(datapath_1_RegisterFile_regfile_mem_18__10_), .B(datapath_1_Instr_16_bF_buf1_), .C(datapath_1_Instr_17_bF_buf5_), .Y(_4116_) );
OAI22X1 OAI22X1_30 ( .A(_4116_), .B(_4115_), .C(datapath_1_Instr_17_bF_buf4_), .D(_4114_), .Y(_4117_) );
NAND2X1 NAND2X1_92 ( .A(_3567__bF_buf3), .B(_4117_), .Y(_4118_) );
MUX2X1 MUX2X1_38 ( .A(datapath_1_RegisterFile_regfile_mem_21__10_), .B(datapath_1_RegisterFile_regfile_mem_20__10_), .S(datapath_1_Instr_16_bF_buf0_), .Y(_4119_) );
NOR2X1 NOR2X1_36 ( .A(datapath_1_RegisterFile_regfile_mem_23__10_), .B(_3588__bF_buf29), .Y(_4120_) );
OAI21X1 OAI21X1_79 ( .A(datapath_1_RegisterFile_regfile_mem_22__10_), .B(datapath_1_Instr_16_bF_buf55_), .C(datapath_1_Instr_17_bF_buf3_), .Y(_4121_) );
OAI22X1 OAI22X1_31 ( .A(_4121_), .B(_4120_), .C(datapath_1_Instr_17_bF_buf2_), .D(_4119_), .Y(_4122_) );
NAND2X1 NAND2X1_93 ( .A(datapath_1_Instr_18_bF_buf21_), .B(_4122_), .Y(_4123_) );
AOI21X1 AOI21X1_85 ( .A(_4118_), .B(_4123_), .C(datapath_1_Instr_19_bF_buf1_), .Y(_4124_) );
OAI21X1 OAI21X1_80 ( .A(_4113_), .B(_4124_), .C(datapath_1_Instr_20_bF_buf3_), .Y(_4125_) );
NAND2X1 NAND2X1_94 ( .A(datapath_1_RegisterFile_regfile_mem_11__10_), .B(datapath_1_Instr_17_bF_buf1_), .Y(_4126_) );
NAND2X1 NAND2X1_95 ( .A(datapath_1_RegisterFile_regfile_mem_9__10_), .B(_3566__bF_buf0), .Y(_4127_) );
NAND3X1 NAND3X1_47 ( .A(datapath_1_Instr_16_bF_buf54_), .B(_4126_), .C(_4127_), .Y(_4128_) );
NAND2X1 NAND2X1_96 ( .A(datapath_1_RegisterFile_regfile_mem_10__10_), .B(datapath_1_Instr_17_bF_buf0_), .Y(_4129_) );
AOI21X1 AOI21X1_86 ( .A(_3566__bF_buf0), .B(datapath_1_RegisterFile_regfile_mem_8__10_), .C(datapath_1_Instr_16_bF_buf53_), .Y(_4130_) );
NAND2X1 NAND2X1_97 ( .A(_4129_), .B(_4130_), .Y(_4131_) );
NAND3X1 NAND3X1_48 ( .A(_3567__bF_buf8), .B(_4128_), .C(_4131_), .Y(_4132_) );
NAND2X1 NAND2X1_98 ( .A(datapath_1_RegisterFile_regfile_mem_15__10_), .B(datapath_1_Instr_17_bF_buf50_), .Y(_4133_) );
NAND2X1 NAND2X1_99 ( .A(datapath_1_RegisterFile_regfile_mem_13__10_), .B(_3566__bF_buf0), .Y(_4134_) );
NAND3X1 NAND3X1_49 ( .A(datapath_1_Instr_16_bF_buf52_), .B(_4133_), .C(_4134_), .Y(_4135_) );
NAND2X1 NAND2X1_100 ( .A(datapath_1_RegisterFile_regfile_mem_14__10_), .B(datapath_1_Instr_17_bF_buf49_), .Y(_4136_) );
AOI21X1 AOI21X1_87 ( .A(_3566__bF_buf0), .B(datapath_1_RegisterFile_regfile_mem_12__10_), .C(datapath_1_Instr_16_bF_buf51_), .Y(_4137_) );
NAND2X1 NAND2X1_101 ( .A(_4136_), .B(_4137_), .Y(_4138_) );
NAND3X1 NAND3X1_50 ( .A(datapath_1_Instr_18_bF_buf20_), .B(_4135_), .C(_4138_), .Y(_4139_) );
AOI21X1 AOI21X1_88 ( .A(_4132_), .B(_4139_), .C(_3571__bF_buf3), .Y(_4140_) );
INVX1 INVX1_25 ( .A(datapath_1_RegisterFile_regfile_mem_1__10_), .Y(_4141_) );
AOI21X1 AOI21X1_89 ( .A(datapath_1_RegisterFile_regfile_mem_5__10_), .B(datapath_1_Instr_18_bF_buf19_), .C(_3588__bF_buf6), .Y(_4142_) );
OAI21X1 OAI21X1_81 ( .A(_4141_), .B(datapath_1_Instr_18_bF_buf18_), .C(_4142_), .Y(_4143_) );
INVX1 INVX1_26 ( .A(datapath_1_RegisterFile_regfile_mem_0__10_), .Y(_4144_) );
AOI21X1 AOI21X1_90 ( .A(datapath_1_RegisterFile_regfile_mem_4__10_), .B(datapath_1_Instr_18_bF_buf17_), .C(datapath_1_Instr_16_bF_buf50_), .Y(_4145_) );
OAI21X1 OAI21X1_82 ( .A(_4144_), .B(datapath_1_Instr_18_bF_buf16_), .C(_4145_), .Y(_4146_) );
NAND3X1 NAND3X1_51 ( .A(_3566__bF_buf7), .B(_4146_), .C(_4143_), .Y(_4147_) );
INVX1 INVX1_27 ( .A(datapath_1_RegisterFile_regfile_mem_3__10_), .Y(_4148_) );
AOI21X1 AOI21X1_91 ( .A(datapath_1_RegisterFile_regfile_mem_7__10_), .B(datapath_1_Instr_18_bF_buf15_), .C(_3588__bF_buf6), .Y(_4149_) );
OAI21X1 OAI21X1_83 ( .A(_4148_), .B(datapath_1_Instr_18_bF_buf14_), .C(_4149_), .Y(_4150_) );
INVX1 INVX1_28 ( .A(datapath_1_RegisterFile_regfile_mem_2__10_), .Y(_4151_) );
AOI21X1 AOI21X1_92 ( .A(datapath_1_RegisterFile_regfile_mem_6__10_), .B(datapath_1_Instr_18_bF_buf13_), .C(datapath_1_Instr_16_bF_buf49_), .Y(_4152_) );
OAI21X1 OAI21X1_84 ( .A(_4151_), .B(datapath_1_Instr_18_bF_buf12_), .C(_4152_), .Y(_4153_) );
NAND3X1 NAND3X1_52 ( .A(datapath_1_Instr_17_bF_buf48_), .B(_4153_), .C(_4150_), .Y(_4154_) );
AOI21X1 AOI21X1_93 ( .A(_4147_), .B(_4154_), .C(datapath_1_Instr_19_bF_buf0_), .Y(_4155_) );
OAI21X1 OAI21X1_85 ( .A(_4155_), .B(_4140_), .C(_3570__bF_buf4), .Y(_4156_) );
AOI22X1 AOI22X1_15 ( .A(_3565__bF_buf2), .B(_3569__bF_buf2), .C(_4156_), .D(_4125_), .Y(datapath_1_RD2_10_) );
NAND2X1 NAND2X1_102 ( .A(datapath_1_RegisterFile_regfile_mem_27__11_), .B(datapath_1_Instr_16_bF_buf48_), .Y(_4157_) );
NAND2X1 NAND2X1_103 ( .A(datapath_1_RegisterFile_regfile_mem_26__11_), .B(_3588__bF_buf11), .Y(_4158_) );
NAND3X1 NAND3X1_53 ( .A(datapath_1_Instr_17_bF_buf47_), .B(_4157_), .C(_4158_), .Y(_4159_) );
NAND2X1 NAND2X1_104 ( .A(datapath_1_RegisterFile_regfile_mem_25__11_), .B(datapath_1_Instr_16_bF_buf47_), .Y(_4160_) );
AOI21X1 AOI21X1_94 ( .A(_3588__bF_buf14), .B(datapath_1_RegisterFile_regfile_mem_24__11_), .C(datapath_1_Instr_17_bF_buf46_), .Y(_4161_) );
NAND2X1 NAND2X1_105 ( .A(_4160_), .B(_4161_), .Y(_4162_) );
NAND3X1 NAND3X1_54 ( .A(_3567__bF_buf10), .B(_4159_), .C(_4162_), .Y(_4163_) );
NAND2X1 NAND2X1_106 ( .A(datapath_1_RegisterFile_regfile_mem_31__11_), .B(datapath_1_Instr_16_bF_buf46_), .Y(_4164_) );
AOI21X1 AOI21X1_95 ( .A(_3588__bF_buf11), .B(datapath_1_RegisterFile_regfile_mem_30__11_), .C(_3566__bF_buf9), .Y(_4165_) );
NAND2X1 NAND2X1_107 ( .A(_4164_), .B(_4165_), .Y(_4166_) );
INVX1 INVX1_29 ( .A(datapath_1_RegisterFile_regfile_mem_28__11_), .Y(_4167_) );
AOI21X1 AOI21X1_96 ( .A(datapath_1_RegisterFile_regfile_mem_29__11_), .B(datapath_1_Instr_16_bF_buf45_), .C(datapath_1_Instr_17_bF_buf45_), .Y(_4168_) );
OAI21X1 OAI21X1_86 ( .A(_4167_), .B(datapath_1_Instr_16_bF_buf44_), .C(_4168_), .Y(_4169_) );
NAND3X1 NAND3X1_55 ( .A(datapath_1_Instr_18_bF_buf11_), .B(_4169_), .C(_4166_), .Y(_4170_) );
AOI21X1 AOI21X1_97 ( .A(_4163_), .B(_4170_), .C(_3571__bF_buf4), .Y(_4171_) );
MUX2X1 MUX2X1_39 ( .A(datapath_1_RegisterFile_regfile_mem_18__11_), .B(datapath_1_RegisterFile_regfile_mem_16__11_), .S(datapath_1_Instr_17_bF_buf44_), .Y(_4172_) );
NAND2X1 NAND2X1_108 ( .A(_3588__bF_buf19), .B(_4172_), .Y(_4173_) );
MUX2X1 MUX2X1_40 ( .A(datapath_1_RegisterFile_regfile_mem_19__11_), .B(datapath_1_RegisterFile_regfile_mem_17__11_), .S(datapath_1_Instr_17_bF_buf43_), .Y(_4174_) );
NAND2X1 NAND2X1_109 ( .A(datapath_1_Instr_16_bF_buf43_), .B(_4174_), .Y(_4175_) );
NAND3X1 NAND3X1_56 ( .A(_3567__bF_buf0), .B(_4173_), .C(_4175_), .Y(_4176_) );
MUX2X1 MUX2X1_41 ( .A(datapath_1_RegisterFile_regfile_mem_22__11_), .B(datapath_1_RegisterFile_regfile_mem_20__11_), .S(datapath_1_Instr_17_bF_buf42_), .Y(_4177_) );
NAND2X1 NAND2X1_110 ( .A(_3588__bF_buf19), .B(_4177_), .Y(_4178_) );
MUX2X1 MUX2X1_42 ( .A(datapath_1_RegisterFile_regfile_mem_23__11_), .B(datapath_1_RegisterFile_regfile_mem_21__11_), .S(datapath_1_Instr_17_bF_buf41_), .Y(_4179_) );
NAND2X1 NAND2X1_111 ( .A(datapath_1_Instr_16_bF_buf42_), .B(_4179_), .Y(_4180_) );
NAND3X1 NAND3X1_57 ( .A(datapath_1_Instr_18_bF_buf10_), .B(_4178_), .C(_4180_), .Y(_4181_) );
AOI21X1 AOI21X1_98 ( .A(_4176_), .B(_4181_), .C(datapath_1_Instr_19_bF_buf6_), .Y(_4182_) );
OAI21X1 OAI21X1_87 ( .A(_4182_), .B(_4171_), .C(datapath_1_Instr_20_bF_buf2_), .Y(_4183_) );
MUX2X1 MUX2X1_43 ( .A(datapath_1_RegisterFile_regfile_mem_9__11_), .B(datapath_1_RegisterFile_regfile_mem_8__11_), .S(datapath_1_Instr_16_bF_buf41_), .Y(_4184_) );
NOR2X1 NOR2X1_37 ( .A(datapath_1_RegisterFile_regfile_mem_11__11_), .B(_3588__bF_buf28), .Y(_4185_) );
OAI21X1 OAI21X1_88 ( .A(datapath_1_RegisterFile_regfile_mem_10__11_), .B(datapath_1_Instr_16_bF_buf40_), .C(datapath_1_Instr_17_bF_buf40_), .Y(_4186_) );
OAI22X1 OAI22X1_32 ( .A(_4186_), .B(_4185_), .C(datapath_1_Instr_17_bF_buf39_), .D(_4184_), .Y(_4187_) );
INVX1 INVX1_30 ( .A(datapath_1_RegisterFile_regfile_mem_15__11_), .Y(_4188_) );
AOI21X1 AOI21X1_99 ( .A(_3588__bF_buf17), .B(datapath_1_RegisterFile_regfile_mem_14__11_), .C(_3566__bF_buf2), .Y(_4189_) );
OAI21X1 OAI21X1_89 ( .A(_4188_), .B(_3588__bF_buf17), .C(_4189_), .Y(_4190_) );
NAND2X1 NAND2X1_112 ( .A(datapath_1_RegisterFile_regfile_mem_12__11_), .B(_3588__bF_buf28), .Y(_4191_) );
AOI21X1 AOI21X1_100 ( .A(datapath_1_RegisterFile_regfile_mem_13__11_), .B(datapath_1_Instr_16_bF_buf39_), .C(datapath_1_Instr_17_bF_buf38_), .Y(_4192_) );
AOI21X1 AOI21X1_101 ( .A(_4191_), .B(_4192_), .C(_3567__bF_buf10), .Y(_4193_) );
AOI22X1 AOI22X1_16 ( .A(_4190_), .B(_4193_), .C(_3567__bF_buf10), .D(_4187_), .Y(_4194_) );
NOR2X1 NOR2X1_38 ( .A(datapath_1_RegisterFile_regfile_mem_0__11_), .B(datapath_1_Instr_16_bF_buf38_), .Y(_4195_) );
OAI21X1 OAI21X1_90 ( .A(datapath_1_RegisterFile_regfile_mem_1__11_), .B(_3588__bF_buf42), .C(_3566__bF_buf7), .Y(_4196_) );
NOR2X1 NOR2X1_39 ( .A(datapath_1_RegisterFile_regfile_mem_3__11_), .B(_3588__bF_buf42), .Y(_4197_) );
OAI21X1 OAI21X1_91 ( .A(datapath_1_RegisterFile_regfile_mem_2__11_), .B(datapath_1_Instr_16_bF_buf37_), .C(datapath_1_Instr_17_bF_buf37_), .Y(_4198_) );
OAI22X1 OAI22X1_33 ( .A(_4197_), .B(_4198_), .C(_4195_), .D(_4196_), .Y(_4199_) );
NOR2X1 NOR2X1_40 ( .A(datapath_1_Instr_18_bF_buf9_), .B(_4199_), .Y(_4200_) );
MUX2X1 MUX2X1_44 ( .A(datapath_1_RegisterFile_regfile_mem_5__11_), .B(datapath_1_RegisterFile_regfile_mem_4__11_), .S(datapath_1_Instr_16_bF_buf36_), .Y(_4201_) );
NOR2X1 NOR2X1_41 ( .A(datapath_1_RegisterFile_regfile_mem_7__11_), .B(_3588__bF_buf13), .Y(_4202_) );
OAI21X1 OAI21X1_92 ( .A(datapath_1_RegisterFile_regfile_mem_6__11_), .B(datapath_1_Instr_16_bF_buf35_), .C(datapath_1_Instr_17_bF_buf36_), .Y(_4203_) );
OAI22X1 OAI22X1_34 ( .A(_4203_), .B(_4202_), .C(datapath_1_Instr_17_bF_buf35_), .D(_4201_), .Y(_4204_) );
OAI21X1 OAI21X1_93 ( .A(_3567__bF_buf10), .B(_4204_), .C(_3571__bF_buf4), .Y(_4205_) );
OAI22X1 OAI22X1_35 ( .A(_3571__bF_buf4), .B(_4194_), .C(_4200_), .D(_4205_), .Y(_4206_) );
NAND2X1 NAND2X1_113 ( .A(_3570__bF_buf1), .B(_4206_), .Y(_4207_) );
AOI22X1 AOI22X1_17 ( .A(_3565__bF_buf0), .B(_3569__bF_buf0), .C(_4183_), .D(_4207_), .Y(datapath_1_RD2_11_) );
NAND2X1 NAND2X1_114 ( .A(datapath_1_RegisterFile_regfile_mem_27__12_), .B(datapath_1_Instr_16_bF_buf34_), .Y(_4208_) );
NAND2X1 NAND2X1_115 ( .A(datapath_1_RegisterFile_regfile_mem_26__12_), .B(_3588__bF_buf13), .Y(_4209_) );
NAND3X1 NAND3X1_58 ( .A(datapath_1_Instr_17_bF_buf34_), .B(_4208_), .C(_4209_), .Y(_4210_) );
NAND2X1 NAND2X1_116 ( .A(datapath_1_RegisterFile_regfile_mem_25__12_), .B(datapath_1_Instr_16_bF_buf33_), .Y(_4211_) );
AOI21X1 AOI21X1_102 ( .A(_3588__bF_buf13), .B(datapath_1_RegisterFile_regfile_mem_24__12_), .C(datapath_1_Instr_17_bF_buf33_), .Y(_4212_) );
NAND2X1 NAND2X1_117 ( .A(_4211_), .B(_4212_), .Y(_4213_) );
NAND3X1 NAND3X1_59 ( .A(_3567__bF_buf5), .B(_4210_), .C(_4213_), .Y(_4214_) );
NAND2X1 NAND2X1_118 ( .A(datapath_1_RegisterFile_regfile_mem_31__12_), .B(datapath_1_Instr_16_bF_buf32_), .Y(_4215_) );
AOI21X1 AOI21X1_103 ( .A(_3588__bF_buf6), .B(datapath_1_RegisterFile_regfile_mem_30__12_), .C(_3566__bF_buf10), .Y(_4216_) );
NAND2X1 NAND2X1_119 ( .A(_4215_), .B(_4216_), .Y(_4217_) );
AOI21X1 AOI21X1_104 ( .A(datapath_1_RegisterFile_regfile_mem_29__12_), .B(datapath_1_Instr_16_bF_buf31_), .C(datapath_1_Instr_17_bF_buf32_), .Y(_4218_) );
OAI21X1 OAI21X1_94 ( .A(_2543_), .B(datapath_1_Instr_16_bF_buf30_), .C(_4218_), .Y(_4219_) );
NAND3X1 NAND3X1_60 ( .A(datapath_1_Instr_18_bF_buf8_), .B(_4219_), .C(_4217_), .Y(_4220_) );
AOI21X1 AOI21X1_105 ( .A(_4214_), .B(_4220_), .C(_3571__bF_buf7), .Y(_4221_) );
MUX2X1 MUX2X1_45 ( .A(datapath_1_RegisterFile_regfile_mem_18__12_), .B(datapath_1_RegisterFile_regfile_mem_16__12_), .S(datapath_1_Instr_17_bF_buf31_), .Y(_4222_) );
NAND2X1 NAND2X1_120 ( .A(_3588__bF_buf13), .B(_4222_), .Y(_4223_) );
MUX2X1 MUX2X1_46 ( .A(datapath_1_RegisterFile_regfile_mem_19__12_), .B(datapath_1_RegisterFile_regfile_mem_17__12_), .S(datapath_1_Instr_17_bF_buf30_), .Y(_4224_) );
NAND2X1 NAND2X1_121 ( .A(datapath_1_Instr_16_bF_buf29_), .B(_4224_), .Y(_4225_) );
NAND3X1 NAND3X1_61 ( .A(_3567__bF_buf5), .B(_4223_), .C(_4225_), .Y(_4226_) );
MUX2X1 MUX2X1_47 ( .A(datapath_1_RegisterFile_regfile_mem_22__12_), .B(datapath_1_RegisterFile_regfile_mem_20__12_), .S(datapath_1_Instr_17_bF_buf29_), .Y(_4227_) );
NAND2X1 NAND2X1_122 ( .A(_3588__bF_buf31), .B(_4227_), .Y(_4228_) );
MUX2X1 MUX2X1_48 ( .A(datapath_1_RegisterFile_regfile_mem_23__12_), .B(datapath_1_RegisterFile_regfile_mem_21__12_), .S(datapath_1_Instr_17_bF_buf28_), .Y(_4229_) );
NAND2X1 NAND2X1_123 ( .A(datapath_1_Instr_16_bF_buf28_), .B(_4229_), .Y(_4230_) );
NAND3X1 NAND3X1_62 ( .A(datapath_1_Instr_18_bF_buf7_), .B(_4228_), .C(_4230_), .Y(_4231_) );
AOI21X1 AOI21X1_106 ( .A(_4226_), .B(_4231_), .C(datapath_1_Instr_19_bF_buf5_), .Y(_4232_) );
OAI21X1 OAI21X1_95 ( .A(_4232_), .B(_4221_), .C(datapath_1_Instr_20_bF_buf1_), .Y(_4233_) );
MUX2X1 MUX2X1_49 ( .A(datapath_1_RegisterFile_regfile_mem_9__12_), .B(datapath_1_RegisterFile_regfile_mem_8__12_), .S(datapath_1_Instr_16_bF_buf27_), .Y(_4234_) );
NOR2X1 NOR2X1_42 ( .A(datapath_1_RegisterFile_regfile_mem_11__12_), .B(_3588__bF_buf1), .Y(_4235_) );
OAI21X1 OAI21X1_96 ( .A(datapath_1_RegisterFile_regfile_mem_10__12_), .B(datapath_1_Instr_16_bF_buf26_), .C(datapath_1_Instr_17_bF_buf27_), .Y(_4236_) );
OAI22X1 OAI22X1_36 ( .A(_4236_), .B(_4235_), .C(datapath_1_Instr_17_bF_buf26_), .D(_4234_), .Y(_4237_) );
AOI21X1 AOI21X1_107 ( .A(_3588__bF_buf8), .B(datapath_1_RegisterFile_regfile_mem_14__12_), .C(_3566__bF_buf0), .Y(_4238_) );
OAI21X1 OAI21X1_97 ( .A(_2564_), .B(_3588__bF_buf8), .C(_4238_), .Y(_4239_) );
NAND2X1 NAND2X1_124 ( .A(datapath_1_RegisterFile_regfile_mem_12__12_), .B(_3588__bF_buf8), .Y(_4240_) );
AOI21X1 AOI21X1_108 ( .A(datapath_1_RegisterFile_regfile_mem_13__12_), .B(datapath_1_Instr_16_bF_buf25_), .C(datapath_1_Instr_17_bF_buf25_), .Y(_4241_) );
AOI21X1 AOI21X1_109 ( .A(_4240_), .B(_4241_), .C(_3567__bF_buf8), .Y(_4242_) );
AOI22X1 AOI22X1_18 ( .A(_4239_), .B(_4242_), .C(_3567__bF_buf4), .D(_4237_), .Y(_4243_) );
NOR2X1 NOR2X1_43 ( .A(datapath_1_RegisterFile_regfile_mem_0__12_), .B(datapath_1_Instr_16_bF_buf24_), .Y(_4244_) );
OAI21X1 OAI21X1_98 ( .A(datapath_1_RegisterFile_regfile_mem_1__12_), .B(_3588__bF_buf43), .C(_3566__bF_buf7), .Y(_4245_) );
NOR2X1 NOR2X1_44 ( .A(datapath_1_RegisterFile_regfile_mem_3__12_), .B(_3588__bF_buf43), .Y(_4246_) );
OAI21X1 OAI21X1_99 ( .A(datapath_1_RegisterFile_regfile_mem_2__12_), .B(datapath_1_Instr_16_bF_buf23_), .C(datapath_1_Instr_17_bF_buf24_), .Y(_4247_) );
OAI22X1 OAI22X1_37 ( .A(_4246_), .B(_4247_), .C(_4244_), .D(_4245_), .Y(_4248_) );
NOR2X1 NOR2X1_45 ( .A(datapath_1_Instr_18_bF_buf6_), .B(_4248_), .Y(_4249_) );
MUX2X1 MUX2X1_50 ( .A(datapath_1_RegisterFile_regfile_mem_5__12_), .B(datapath_1_RegisterFile_regfile_mem_4__12_), .S(datapath_1_Instr_16_bF_buf22_), .Y(_4250_) );
NOR2X1 NOR2X1_46 ( .A(datapath_1_RegisterFile_regfile_mem_7__12_), .B(_3588__bF_buf9), .Y(_4251_) );
OAI21X1 OAI21X1_100 ( .A(datapath_1_RegisterFile_regfile_mem_6__12_), .B(datapath_1_Instr_16_bF_buf21_), .C(datapath_1_Instr_17_bF_buf23_), .Y(_4252_) );
OAI22X1 OAI22X1_38 ( .A(_4252_), .B(_4251_), .C(datapath_1_Instr_17_bF_buf22_), .D(_4250_), .Y(_4253_) );
OAI21X1 OAI21X1_101 ( .A(_3567__bF_buf4), .B(_4253_), .C(_3571__bF_buf1), .Y(_4254_) );
OAI22X1 OAI22X1_39 ( .A(_3571__bF_buf1), .B(_4243_), .C(_4249_), .D(_4254_), .Y(_4255_) );
NAND2X1 NAND2X1_125 ( .A(_3570__bF_buf3), .B(_4255_), .Y(_4256_) );
AOI22X1 AOI22X1_19 ( .A(_3565__bF_buf1), .B(_3569__bF_buf1), .C(_4233_), .D(_4256_), .Y(datapath_1_RD2_12_) );
MUX2X1 MUX2X1_51 ( .A(datapath_1_RegisterFile_regfile_mem_9__13_), .B(datapath_1_RegisterFile_regfile_mem_8__13_), .S(datapath_1_Instr_16_bF_buf20_), .Y(_4257_) );
NOR2X1 NOR2X1_47 ( .A(datapath_1_RegisterFile_regfile_mem_11__13_), .B(_3588__bF_buf10), .Y(_4258_) );
OAI21X1 OAI21X1_102 ( .A(datapath_1_RegisterFile_regfile_mem_10__13_), .B(datapath_1_Instr_16_bF_buf19_), .C(datapath_1_Instr_17_bF_buf21_), .Y(_4259_) );
OAI22X1 OAI22X1_40 ( .A(_4259_), .B(_4258_), .C(datapath_1_Instr_17_bF_buf20_), .D(_4257_), .Y(_4260_) );
AOI21X1 AOI21X1_110 ( .A(_3588__bF_buf10), .B(datapath_1_RegisterFile_regfile_mem_14__13_), .C(_3566__bF_buf3), .Y(_4261_) );
OAI21X1 OAI21X1_103 ( .A(_2615_), .B(_3588__bF_buf10), .C(_4261_), .Y(_4262_) );
NAND2X1 NAND2X1_126 ( .A(datapath_1_RegisterFile_regfile_mem_12__13_), .B(_3588__bF_buf4), .Y(_4263_) );
AOI21X1 AOI21X1_111 ( .A(datapath_1_RegisterFile_regfile_mem_13__13_), .B(datapath_1_Instr_16_bF_buf18_), .C(datapath_1_Instr_17_bF_buf19_), .Y(_4264_) );
AOI21X1 AOI21X1_112 ( .A(_4263_), .B(_4264_), .C(_3567__bF_buf1), .Y(_4265_) );
AOI22X1 AOI22X1_20 ( .A(_4262_), .B(_4265_), .C(_3567__bF_buf1), .D(_4260_), .Y(_4266_) );
NOR2X1 NOR2X1_48 ( .A(datapath_1_RegisterFile_regfile_mem_0__13_), .B(datapath_1_Instr_16_bF_buf17_), .Y(_4267_) );
OAI21X1 OAI21X1_104 ( .A(datapath_1_RegisterFile_regfile_mem_1__13_), .B(_3588__bF_buf30), .C(_3566__bF_buf6), .Y(_4268_) );
NOR2X1 NOR2X1_49 ( .A(datapath_1_RegisterFile_regfile_mem_3__13_), .B(_3588__bF_buf30), .Y(_4269_) );
OAI21X1 OAI21X1_105 ( .A(datapath_1_RegisterFile_regfile_mem_2__13_), .B(datapath_1_Instr_16_bF_buf16_), .C(datapath_1_Instr_17_bF_buf18_), .Y(_4270_) );
OAI22X1 OAI22X1_41 ( .A(_4269_), .B(_4270_), .C(_4267_), .D(_4268_), .Y(_4271_) );
NOR2X1 NOR2X1_50 ( .A(datapath_1_Instr_18_bF_buf5_), .B(_4271_), .Y(_4272_) );
MUX2X1 MUX2X1_52 ( .A(datapath_1_RegisterFile_regfile_mem_5__13_), .B(datapath_1_RegisterFile_regfile_mem_4__13_), .S(datapath_1_Instr_16_bF_buf15_), .Y(_4273_) );
NOR2X1 NOR2X1_51 ( .A(datapath_1_RegisterFile_regfile_mem_7__13_), .B(_3588__bF_buf30), .Y(_4274_) );
OAI21X1 OAI21X1_106 ( .A(datapath_1_RegisterFile_regfile_mem_6__13_), .B(datapath_1_Instr_16_bF_buf14_), .C(datapath_1_Instr_17_bF_buf17_), .Y(_4275_) );
OAI22X1 OAI22X1_42 ( .A(_4275_), .B(_4274_), .C(datapath_1_Instr_17_bF_buf16_), .D(_4273_), .Y(_4276_) );
OAI21X1 OAI21X1_107 ( .A(_3567__bF_buf1), .B(_4276_), .C(_3571__bF_buf2), .Y(_4277_) );
OAI22X1 OAI22X1_43 ( .A(_3571__bF_buf2), .B(_4266_), .C(_4272_), .D(_4277_), .Y(_4278_) );
NAND2X1 NAND2X1_127 ( .A(_3570__bF_buf4), .B(_4278_), .Y(_4279_) );
INVX1 INVX1_31 ( .A(datapath_1_RegisterFile_regfile_mem_27__13_), .Y(_4280_) );
AOI21X1 AOI21X1_113 ( .A(datapath_1_RegisterFile_regfile_mem_31__13_), .B(datapath_1_Instr_18_bF_buf4_), .C(_3588__bF_buf41), .Y(_4281_) );
OAI21X1 OAI21X1_108 ( .A(_4280_), .B(datapath_1_Instr_18_bF_buf3_), .C(_4281_), .Y(_4282_) );
INVX1 INVX1_32 ( .A(datapath_1_RegisterFile_regfile_mem_26__13_), .Y(_4283_) );
AOI21X1 AOI21X1_114 ( .A(datapath_1_RegisterFile_regfile_mem_30__13_), .B(datapath_1_Instr_18_bF_buf2_), .C(datapath_1_Instr_16_bF_buf13_), .Y(_4284_) );
OAI21X1 OAI21X1_109 ( .A(_4283_), .B(datapath_1_Instr_18_bF_buf1_), .C(_4284_), .Y(_4285_) );
NAND3X1 NAND3X1_63 ( .A(datapath_1_Instr_17_bF_buf15_), .B(_4285_), .C(_4282_), .Y(_4286_) );
INVX1 INVX1_33 ( .A(datapath_1_RegisterFile_regfile_mem_25__13_), .Y(_4287_) );
AOI21X1 AOI21X1_115 ( .A(datapath_1_RegisterFile_regfile_mem_29__13_), .B(datapath_1_Instr_18_bF_buf0_), .C(_3588__bF_buf29), .Y(_4288_) );
OAI21X1 OAI21X1_110 ( .A(_4287_), .B(datapath_1_Instr_18_bF_buf44_), .C(_4288_), .Y(_4289_) );
INVX1 INVX1_34 ( .A(datapath_1_RegisterFile_regfile_mem_24__13_), .Y(_4290_) );
AOI21X1 AOI21X1_116 ( .A(datapath_1_RegisterFile_regfile_mem_28__13_), .B(datapath_1_Instr_18_bF_buf43_), .C(datapath_1_Instr_16_bF_buf12_), .Y(_4291_) );
OAI21X1 OAI21X1_111 ( .A(_4290_), .B(datapath_1_Instr_18_bF_buf42_), .C(_4291_), .Y(_4292_) );
NAND3X1 NAND3X1_64 ( .A(_3566__bF_buf4), .B(_4292_), .C(_4289_), .Y(_4293_) );
AOI21X1 AOI21X1_117 ( .A(_4286_), .B(_4293_), .C(_3571__bF_buf5), .Y(_4294_) );
MUX2X1 MUX2X1_53 ( .A(datapath_1_RegisterFile_regfile_mem_18__13_), .B(datapath_1_RegisterFile_regfile_mem_16__13_), .S(datapath_1_Instr_17_bF_buf14_), .Y(_4295_) );
NAND2X1 NAND2X1_128 ( .A(_3588__bF_buf32), .B(_4295_), .Y(_4296_) );
MUX2X1 MUX2X1_54 ( .A(datapath_1_RegisterFile_regfile_mem_19__13_), .B(datapath_1_RegisterFile_regfile_mem_17__13_), .S(datapath_1_Instr_17_bF_buf13_), .Y(_4297_) );
NAND2X1 NAND2X1_129 ( .A(datapath_1_Instr_16_bF_buf11_), .B(_4297_), .Y(_4298_) );
NAND3X1 NAND3X1_65 ( .A(_3567__bF_buf9), .B(_4296_), .C(_4298_), .Y(_4299_) );
MUX2X1 MUX2X1_55 ( .A(datapath_1_RegisterFile_regfile_mem_22__13_), .B(datapath_1_RegisterFile_regfile_mem_20__13_), .S(datapath_1_Instr_17_bF_buf12_), .Y(_4300_) );
NAND2X1 NAND2X1_130 ( .A(_3588__bF_buf27), .B(_4300_), .Y(_4301_) );
MUX2X1 MUX2X1_56 ( .A(datapath_1_RegisterFile_regfile_mem_23__13_), .B(datapath_1_RegisterFile_regfile_mem_21__13_), .S(datapath_1_Instr_17_bF_buf11_), .Y(_4302_) );
NAND2X1 NAND2X1_131 ( .A(datapath_1_Instr_16_bF_buf10_), .B(_4302_), .Y(_4303_) );
NAND3X1 NAND3X1_66 ( .A(datapath_1_Instr_18_bF_buf41_), .B(_4301_), .C(_4303_), .Y(_4304_) );
AOI21X1 AOI21X1_118 ( .A(_4299_), .B(_4304_), .C(datapath_1_Instr_19_bF_buf4_), .Y(_4305_) );
OAI21X1 OAI21X1_112 ( .A(_4294_), .B(_4305_), .C(datapath_1_Instr_20_bF_buf0_), .Y(_4306_) );
AOI22X1 AOI22X1_21 ( .A(_3565__bF_buf3), .B(_3569__bF_buf3), .C(_4306_), .D(_4279_), .Y(datapath_1_RD2_13_) );
NAND2X1 NAND2X1_132 ( .A(datapath_1_RegisterFile_regfile_mem_27__14_), .B(datapath_1_Instr_16_bF_buf9_), .Y(_4307_) );
NAND2X1 NAND2X1_133 ( .A(datapath_1_RegisterFile_regfile_mem_26__14_), .B(_3588__bF_buf38), .Y(_4308_) );
NAND3X1 NAND3X1_67 ( .A(datapath_1_Instr_17_bF_buf10_), .B(_4307_), .C(_4308_), .Y(_4309_) );
NAND2X1 NAND2X1_134 ( .A(datapath_1_RegisterFile_regfile_mem_25__14_), .B(datapath_1_Instr_16_bF_buf8_), .Y(_4310_) );
AOI21X1 AOI21X1_119 ( .A(_3588__bF_buf38), .B(datapath_1_RegisterFile_regfile_mem_24__14_), .C(datapath_1_Instr_17_bF_buf9_), .Y(_4311_) );
NAND2X1 NAND2X1_135 ( .A(_4310_), .B(_4311_), .Y(_4312_) );
NAND3X1 NAND3X1_68 ( .A(_3567__bF_buf9), .B(_4309_), .C(_4312_), .Y(_4313_) );
NAND2X1 NAND2X1_136 ( .A(datapath_1_RegisterFile_regfile_mem_31__14_), .B(datapath_1_Instr_16_bF_buf7_), .Y(_4314_) );
AOI21X1 AOI21X1_120 ( .A(_3588__bF_buf20), .B(datapath_1_RegisterFile_regfile_mem_30__14_), .C(_3566__bF_buf6), .Y(_4315_) );
NAND2X1 NAND2X1_137 ( .A(_4314_), .B(_4315_), .Y(_4316_) );
AOI21X1 AOI21X1_121 ( .A(datapath_1_RegisterFile_regfile_mem_29__14_), .B(datapath_1_Instr_16_bF_buf6_), .C(datapath_1_Instr_17_bF_buf8_), .Y(_4317_) );
OAI21X1 OAI21X1_113 ( .A(_2645_), .B(datapath_1_Instr_16_bF_buf5_), .C(_4317_), .Y(_4318_) );
NAND3X1 NAND3X1_69 ( .A(datapath_1_Instr_18_bF_buf40_), .B(_4318_), .C(_4316_), .Y(_4319_) );
AOI21X1 AOI21X1_122 ( .A(_4313_), .B(_4319_), .C(_3571__bF_buf2), .Y(_4320_) );
MUX2X1 MUX2X1_57 ( .A(datapath_1_RegisterFile_regfile_mem_17__14_), .B(datapath_1_RegisterFile_regfile_mem_16__14_), .S(datapath_1_Instr_16_bF_buf4_), .Y(_4321_) );
NOR2X1 NOR2X1_52 ( .A(datapath_1_RegisterFile_regfile_mem_19__14_), .B(_3588__bF_buf23), .Y(_4322_) );
OAI21X1 OAI21X1_114 ( .A(datapath_1_RegisterFile_regfile_mem_18__14_), .B(datapath_1_Instr_16_bF_buf3_), .C(datapath_1_Instr_17_bF_buf7_), .Y(_4323_) );
OAI22X1 OAI22X1_44 ( .A(_4323_), .B(_4322_), .C(datapath_1_Instr_17_bF_buf6_), .D(_4321_), .Y(_4324_) );
NAND2X1 NAND2X1_138 ( .A(_3567__bF_buf9), .B(_4324_), .Y(_4325_) );
MUX2X1 MUX2X1_58 ( .A(datapath_1_RegisterFile_regfile_mem_21__14_), .B(datapath_1_RegisterFile_regfile_mem_20__14_), .S(datapath_1_Instr_16_bF_buf2_), .Y(_4326_) );
NOR2X1 NOR2X1_53 ( .A(datapath_1_RegisterFile_regfile_mem_23__14_), .B(_3588__bF_buf32), .Y(_4327_) );
OAI21X1 OAI21X1_115 ( .A(datapath_1_RegisterFile_regfile_mem_22__14_), .B(datapath_1_Instr_16_bF_buf1_), .C(datapath_1_Instr_17_bF_buf5_), .Y(_4328_) );
OAI22X1 OAI22X1_45 ( .A(_4328_), .B(_4327_), .C(datapath_1_Instr_17_bF_buf4_), .D(_4326_), .Y(_4329_) );
NAND2X1 NAND2X1_139 ( .A(datapath_1_Instr_18_bF_buf39_), .B(_4329_), .Y(_4330_) );
AOI21X1 AOI21X1_123 ( .A(_4325_), .B(_4330_), .C(datapath_1_Instr_19_bF_buf3_), .Y(_4331_) );
OAI21X1 OAI21X1_116 ( .A(_4320_), .B(_4331_), .C(datapath_1_Instr_20_bF_buf5_), .Y(_4332_) );
NAND2X1 NAND2X1_140 ( .A(datapath_1_RegisterFile_regfile_mem_11__14_), .B(datapath_1_Instr_17_bF_buf3_), .Y(_4333_) );
NAND2X1 NAND2X1_141 ( .A(datapath_1_RegisterFile_regfile_mem_9__14_), .B(_3566__bF_buf5), .Y(_4334_) );
NAND3X1 NAND3X1_70 ( .A(datapath_1_Instr_16_bF_buf0_), .B(_4333_), .C(_4334_), .Y(_4335_) );
NAND2X1 NAND2X1_142 ( .A(datapath_1_RegisterFile_regfile_mem_10__14_), .B(datapath_1_Instr_17_bF_buf2_), .Y(_4336_) );
AOI21X1 AOI21X1_124 ( .A(_3566__bF_buf5), .B(datapath_1_RegisterFile_regfile_mem_8__14_), .C(datapath_1_Instr_16_bF_buf55_), .Y(_4337_) );
NAND2X1 NAND2X1_143 ( .A(_4336_), .B(_4337_), .Y(_4338_) );
NAND3X1 NAND3X1_71 ( .A(_3567__bF_buf8), .B(_4335_), .C(_4338_), .Y(_4339_) );
NAND2X1 NAND2X1_144 ( .A(datapath_1_RegisterFile_regfile_mem_15__14_), .B(datapath_1_Instr_17_bF_buf1_), .Y(_4340_) );
NAND2X1 NAND2X1_145 ( .A(datapath_1_RegisterFile_regfile_mem_13__14_), .B(_3566__bF_buf5), .Y(_4341_) );
NAND3X1 NAND3X1_72 ( .A(datapath_1_Instr_16_bF_buf54_), .B(_4340_), .C(_4341_), .Y(_4342_) );
NAND2X1 NAND2X1_146 ( .A(datapath_1_RegisterFile_regfile_mem_14__14_), .B(datapath_1_Instr_17_bF_buf0_), .Y(_4343_) );
AOI21X1 AOI21X1_125 ( .A(_3566__bF_buf5), .B(datapath_1_RegisterFile_regfile_mem_12__14_), .C(datapath_1_Instr_16_bF_buf53_), .Y(_4344_) );
NAND2X1 NAND2X1_147 ( .A(_4343_), .B(_4344_), .Y(_4345_) );
NAND3X1 NAND3X1_73 ( .A(datapath_1_Instr_18_bF_buf38_), .B(_4342_), .C(_4345_), .Y(_4346_) );
AOI21X1 AOI21X1_126 ( .A(_4339_), .B(_4346_), .C(_3571__bF_buf6), .Y(_4347_) );
INVX1 INVX1_35 ( .A(datapath_1_RegisterFile_regfile_mem_1__14_), .Y(_4348_) );
AOI21X1 AOI21X1_127 ( .A(datapath_1_RegisterFile_regfile_mem_5__14_), .B(datapath_1_Instr_18_bF_buf37_), .C(_3588__bF_buf7), .Y(_4349_) );
OAI21X1 OAI21X1_117 ( .A(_4348_), .B(datapath_1_Instr_18_bF_buf36_), .C(_4349_), .Y(_4350_) );
INVX1 INVX1_36 ( .A(datapath_1_RegisterFile_regfile_mem_0__14_), .Y(_4351_) );
AOI21X1 AOI21X1_128 ( .A(datapath_1_RegisterFile_regfile_mem_4__14_), .B(datapath_1_Instr_18_bF_buf35_), .C(datapath_1_Instr_16_bF_buf52_), .Y(_4352_) );
OAI21X1 OAI21X1_118 ( .A(_4351_), .B(datapath_1_Instr_18_bF_buf34_), .C(_4352_), .Y(_4353_) );
NAND3X1 NAND3X1_74 ( .A(_3566__bF_buf5), .B(_4353_), .C(_4350_), .Y(_4354_) );
INVX1 INVX1_37 ( .A(datapath_1_RegisterFile_regfile_mem_3__14_), .Y(_4355_) );
AOI21X1 AOI21X1_129 ( .A(datapath_1_RegisterFile_regfile_mem_7__14_), .B(datapath_1_Instr_18_bF_buf33_), .C(_3588__bF_buf3), .Y(_4356_) );
OAI21X1 OAI21X1_119 ( .A(_4355_), .B(datapath_1_Instr_18_bF_buf32_), .C(_4356_), .Y(_4357_) );
INVX1 INVX1_38 ( .A(datapath_1_RegisterFile_regfile_mem_2__14_), .Y(_4358_) );
AOI21X1 AOI21X1_130 ( .A(datapath_1_RegisterFile_regfile_mem_6__14_), .B(datapath_1_Instr_18_bF_buf31_), .C(datapath_1_Instr_16_bF_buf51_), .Y(_4359_) );
OAI21X1 OAI21X1_120 ( .A(_4358_), .B(datapath_1_Instr_18_bF_buf30_), .C(_4359_), .Y(_4360_) );
NAND3X1 NAND3X1_75 ( .A(datapath_1_Instr_17_bF_buf50_), .B(_4360_), .C(_4357_), .Y(_4361_) );
AOI21X1 AOI21X1_131 ( .A(_4354_), .B(_4361_), .C(datapath_1_Instr_19_bF_buf2_), .Y(_4362_) );
OAI21X1 OAI21X1_121 ( .A(_4362_), .B(_4347_), .C(_3570__bF_buf0), .Y(_4363_) );
AOI22X1 AOI22X1_22 ( .A(_3565__bF_buf3), .B(_3569__bF_buf3), .C(_4363_), .D(_4332_), .Y(datapath_1_RD2_14_) );
NAND2X1 NAND2X1_148 ( .A(datapath_1_RegisterFile_regfile_mem_27__15_), .B(datapath_1_Instr_16_bF_buf50_), .Y(_4364_) );
NAND2X1 NAND2X1_149 ( .A(datapath_1_RegisterFile_regfile_mem_26__15_), .B(_3588__bF_buf11), .Y(_4365_) );
NAND3X1 NAND3X1_76 ( .A(datapath_1_Instr_17_bF_buf49_), .B(_4364_), .C(_4365_), .Y(_4366_) );
NAND2X1 NAND2X1_150 ( .A(datapath_1_RegisterFile_regfile_mem_25__15_), .B(datapath_1_Instr_16_bF_buf49_), .Y(_4367_) );
AOI21X1 AOI21X1_132 ( .A(_3588__bF_buf11), .B(datapath_1_RegisterFile_regfile_mem_24__15_), .C(datapath_1_Instr_17_bF_buf48_), .Y(_4368_) );
NAND2X1 NAND2X1_151 ( .A(_4367_), .B(_4368_), .Y(_4369_) );
NAND3X1 NAND3X1_77 ( .A(_3567__bF_buf5), .B(_4366_), .C(_4369_), .Y(_4370_) );
NAND2X1 NAND2X1_152 ( .A(datapath_1_RegisterFile_regfile_mem_31__15_), .B(datapath_1_Instr_16_bF_buf48_), .Y(_4371_) );
AOI21X1 AOI21X1_133 ( .A(_3588__bF_buf26), .B(datapath_1_RegisterFile_regfile_mem_30__15_), .C(_3566__bF_buf9), .Y(_4372_) );
NAND2X1 NAND2X1_153 ( .A(_4371_), .B(_4372_), .Y(_4373_) );
AOI21X1 AOI21X1_134 ( .A(datapath_1_RegisterFile_regfile_mem_29__15_), .B(datapath_1_Instr_16_bF_buf47_), .C(datapath_1_Instr_17_bF_buf47_), .Y(_4374_) );
OAI21X1 OAI21X1_122 ( .A(_2696_), .B(datapath_1_Instr_16_bF_buf46_), .C(_4374_), .Y(_4375_) );
NAND3X1 NAND3X1_78 ( .A(datapath_1_Instr_18_bF_buf29_), .B(_4375_), .C(_4373_), .Y(_4376_) );
AOI21X1 AOI21X1_135 ( .A(_4370_), .B(_4376_), .C(_3571__bF_buf7), .Y(_4377_) );
MUX2X1 MUX2X1_59 ( .A(datapath_1_RegisterFile_regfile_mem_18__15_), .B(datapath_1_RegisterFile_regfile_mem_16__15_), .S(datapath_1_Instr_17_bF_buf46_), .Y(_4378_) );
NAND2X1 NAND2X1_154 ( .A(_3588__bF_buf19), .B(_4378_), .Y(_4379_) );
MUX2X1 MUX2X1_60 ( .A(datapath_1_RegisterFile_regfile_mem_19__15_), .B(datapath_1_RegisterFile_regfile_mem_17__15_), .S(datapath_1_Instr_17_bF_buf45_), .Y(_4380_) );
NAND2X1 NAND2X1_155 ( .A(datapath_1_Instr_16_bF_buf45_), .B(_4380_), .Y(_4381_) );
NAND3X1 NAND3X1_79 ( .A(_3567__bF_buf0), .B(_4379_), .C(_4381_), .Y(_4382_) );
MUX2X1 MUX2X1_61 ( .A(datapath_1_RegisterFile_regfile_mem_22__15_), .B(datapath_1_RegisterFile_regfile_mem_20__15_), .S(datapath_1_Instr_17_bF_buf44_), .Y(_4383_) );
NAND2X1 NAND2X1_156 ( .A(_3588__bF_buf14), .B(_4383_), .Y(_4384_) );
MUX2X1 MUX2X1_62 ( .A(datapath_1_RegisterFile_regfile_mem_23__15_), .B(datapath_1_RegisterFile_regfile_mem_21__15_), .S(datapath_1_Instr_17_bF_buf43_), .Y(_4385_) );
NAND2X1 NAND2X1_157 ( .A(datapath_1_Instr_16_bF_buf44_), .B(_4385_), .Y(_4386_) );
NAND3X1 NAND3X1_80 ( .A(datapath_1_Instr_18_bF_buf28_), .B(_4384_), .C(_4386_), .Y(_4387_) );
AOI21X1 AOI21X1_136 ( .A(_4382_), .B(_4387_), .C(datapath_1_Instr_19_bF_buf1_), .Y(_4388_) );
OAI21X1 OAI21X1_123 ( .A(_4388_), .B(_4377_), .C(datapath_1_Instr_20_bF_buf4_), .Y(_4389_) );
MUX2X1 MUX2X1_63 ( .A(datapath_1_RegisterFile_regfile_mem_9__15_), .B(datapath_1_RegisterFile_regfile_mem_8__15_), .S(datapath_1_Instr_16_bF_buf43_), .Y(_4390_) );
NOR2X1 NOR2X1_54 ( .A(datapath_1_RegisterFile_regfile_mem_11__15_), .B(_3588__bF_buf22), .Y(_4391_) );
OAI21X1 OAI21X1_124 ( .A(datapath_1_RegisterFile_regfile_mem_10__15_), .B(datapath_1_Instr_16_bF_buf42_), .C(datapath_1_Instr_17_bF_buf42_), .Y(_4392_) );
OAI22X1 OAI22X1_46 ( .A(_4392_), .B(_4391_), .C(datapath_1_Instr_17_bF_buf41_), .D(_4390_), .Y(_4393_) );
AOI21X1 AOI21X1_137 ( .A(_3588__bF_buf22), .B(datapath_1_RegisterFile_regfile_mem_14__15_), .C(_3566__bF_buf2), .Y(_4394_) );
OAI21X1 OAI21X1_125 ( .A(_2717_), .B(_3588__bF_buf22), .C(_4394_), .Y(_4395_) );
NAND2X1 NAND2X1_158 ( .A(datapath_1_RegisterFile_regfile_mem_12__15_), .B(_3588__bF_buf17), .Y(_4396_) );
AOI21X1 AOI21X1_138 ( .A(datapath_1_RegisterFile_regfile_mem_13__15_), .B(datapath_1_Instr_16_bF_buf41_), .C(datapath_1_Instr_17_bF_buf40_), .Y(_4397_) );
AOI21X1 AOI21X1_139 ( .A(_4396_), .B(_4397_), .C(_3567__bF_buf7), .Y(_4398_) );
AOI22X1 AOI22X1_23 ( .A(_4395_), .B(_4398_), .C(_3567__bF_buf7), .D(_4393_), .Y(_4399_) );
NOR2X1 NOR2X1_55 ( .A(datapath_1_RegisterFile_regfile_mem_0__15_), .B(datapath_1_Instr_16_bF_buf40_), .Y(_4400_) );
OAI21X1 OAI21X1_126 ( .A(datapath_1_RegisterFile_regfile_mem_1__15_), .B(_3588__bF_buf17), .C(_3566__bF_buf2), .Y(_4401_) );
NOR2X1 NOR2X1_56 ( .A(datapath_1_RegisterFile_regfile_mem_3__15_), .B(_3588__bF_buf34), .Y(_4402_) );
OAI21X1 OAI21X1_127 ( .A(datapath_1_RegisterFile_regfile_mem_2__15_), .B(datapath_1_Instr_16_bF_buf39_), .C(datapath_1_Instr_17_bF_buf39_), .Y(_4403_) );
OAI22X1 OAI22X1_47 ( .A(_4402_), .B(_4403_), .C(_4400_), .D(_4401_), .Y(_4404_) );
NOR2X1 NOR2X1_57 ( .A(datapath_1_Instr_18_bF_buf27_), .B(_4404_), .Y(_4405_) );
MUX2X1 MUX2X1_64 ( .A(datapath_1_RegisterFile_regfile_mem_5__15_), .B(datapath_1_RegisterFile_regfile_mem_4__15_), .S(datapath_1_Instr_16_bF_buf38_), .Y(_4406_) );
NOR2X1 NOR2X1_58 ( .A(datapath_1_RegisterFile_regfile_mem_7__15_), .B(_3588__bF_buf28), .Y(_4407_) );
OAI21X1 OAI21X1_128 ( .A(datapath_1_RegisterFile_regfile_mem_6__15_), .B(datapath_1_Instr_16_bF_buf37_), .C(datapath_1_Instr_17_bF_buf38_), .Y(_4408_) );
OAI22X1 OAI22X1_48 ( .A(_4408_), .B(_4407_), .C(datapath_1_Instr_17_bF_buf37_), .D(_4406_), .Y(_4409_) );
OAI21X1 OAI21X1_129 ( .A(_3567__bF_buf10), .B(_4409_), .C(_3571__bF_buf0), .Y(_4410_) );
OAI22X1 OAI22X1_49 ( .A(_3571__bF_buf0), .B(_4399_), .C(_4405_), .D(_4410_), .Y(_4411_) );
NAND2X1 NAND2X1_159 ( .A(_3570__bF_buf1), .B(_4411_), .Y(_4412_) );
AOI22X1 AOI22X1_24 ( .A(_3565__bF_buf0), .B(_3569__bF_buf0), .C(_4389_), .D(_4412_), .Y(datapath_1_RD2_15_) );
MUX2X1 MUX2X1_65 ( .A(datapath_1_RegisterFile_regfile_mem_9__16_), .B(datapath_1_RegisterFile_regfile_mem_8__16_), .S(datapath_1_Instr_16_bF_buf36_), .Y(_4413_) );
NOR2X1 NOR2X1_59 ( .A(datapath_1_RegisterFile_regfile_mem_11__16_), .B(_3588__bF_buf22), .Y(_4414_) );
OAI21X1 OAI21X1_130 ( .A(datapath_1_RegisterFile_regfile_mem_10__16_), .B(datapath_1_Instr_16_bF_buf35_), .C(datapath_1_Instr_17_bF_buf36_), .Y(_4415_) );
OAI22X1 OAI22X1_50 ( .A(_4415_), .B(_4414_), .C(datapath_1_Instr_17_bF_buf35_), .D(_4413_), .Y(_4416_) );
AOI21X1 AOI21X1_140 ( .A(_3588__bF_buf34), .B(datapath_1_RegisterFile_regfile_mem_14__16_), .C(_3566__bF_buf2), .Y(_4417_) );
OAI21X1 OAI21X1_131 ( .A(_2741_), .B(_3588__bF_buf34), .C(_4417_), .Y(_4418_) );
NAND2X1 NAND2X1_160 ( .A(datapath_1_RegisterFile_regfile_mem_12__16_), .B(_3588__bF_buf34), .Y(_4419_) );
AOI21X1 AOI21X1_141 ( .A(datapath_1_RegisterFile_regfile_mem_13__16_), .B(datapath_1_Instr_16_bF_buf34_), .C(datapath_1_Instr_17_bF_buf34_), .Y(_4420_) );
AOI21X1 AOI21X1_142 ( .A(_4419_), .B(_4420_), .C(_3567__bF_buf7), .Y(_4421_) );
AOI22X1 AOI22X1_25 ( .A(_4418_), .B(_4421_), .C(_3567__bF_buf7), .D(_4416_), .Y(_4422_) );
NOR2X1 NOR2X1_60 ( .A(datapath_1_RegisterFile_regfile_mem_0__16_), .B(datapath_1_Instr_16_bF_buf33_), .Y(_4423_) );
OAI21X1 OAI21X1_132 ( .A(datapath_1_RegisterFile_regfile_mem_1__16_), .B(_3588__bF_buf36), .C(_3566__bF_buf1), .Y(_4424_) );
NOR2X1 NOR2X1_61 ( .A(datapath_1_RegisterFile_regfile_mem_3__16_), .B(_3588__bF_buf36), .Y(_4425_) );
OAI21X1 OAI21X1_133 ( .A(datapath_1_RegisterFile_regfile_mem_2__16_), .B(datapath_1_Instr_16_bF_buf32_), .C(datapath_1_Instr_17_bF_buf33_), .Y(_4426_) );
OAI22X1 OAI22X1_51 ( .A(_4425_), .B(_4426_), .C(_4423_), .D(_4424_), .Y(_4427_) );
NOR2X1 NOR2X1_62 ( .A(datapath_1_Instr_18_bF_buf26_), .B(_4427_), .Y(_4428_) );
MUX2X1 MUX2X1_66 ( .A(datapath_1_RegisterFile_regfile_mem_5__16_), .B(datapath_1_RegisterFile_regfile_mem_4__16_), .S(datapath_1_Instr_16_bF_buf31_), .Y(_4429_) );
NOR2X1 NOR2X1_63 ( .A(datapath_1_RegisterFile_regfile_mem_7__16_), .B(_3588__bF_buf36), .Y(_4430_) );
OAI21X1 OAI21X1_134 ( .A(datapath_1_RegisterFile_regfile_mem_6__16_), .B(datapath_1_Instr_16_bF_buf30_), .C(datapath_1_Instr_17_bF_buf32_), .Y(_4431_) );
OAI22X1 OAI22X1_52 ( .A(_4431_), .B(_4430_), .C(datapath_1_Instr_17_bF_buf31_), .D(_4429_), .Y(_4432_) );
OAI21X1 OAI21X1_135 ( .A(_3567__bF_buf4), .B(_4432_), .C(_3571__bF_buf0), .Y(_4433_) );
OAI22X1 OAI22X1_53 ( .A(_3571__bF_buf1), .B(_4422_), .C(_4428_), .D(_4433_), .Y(_4434_) );
NAND2X1 NAND2X1_161 ( .A(_3570__bF_buf2), .B(_4434_), .Y(_4435_) );
INVX1 INVX1_39 ( .A(datapath_1_RegisterFile_regfile_mem_27__16_), .Y(_4436_) );
AOI21X1 AOI21X1_143 ( .A(datapath_1_RegisterFile_regfile_mem_31__16_), .B(datapath_1_Instr_18_bF_buf25_), .C(_3588__bF_buf31), .Y(_4437_) );
OAI21X1 OAI21X1_136 ( .A(_4436_), .B(datapath_1_Instr_18_bF_buf24_), .C(_4437_), .Y(_4438_) );
INVX1 INVX1_40 ( .A(datapath_1_RegisterFile_regfile_mem_26__16_), .Y(_4439_) );
AOI21X1 AOI21X1_144 ( .A(datapath_1_RegisterFile_regfile_mem_30__16_), .B(datapath_1_Instr_18_bF_buf23_), .C(datapath_1_Instr_16_bF_buf29_), .Y(_4440_) );
OAI21X1 OAI21X1_137 ( .A(_4439_), .B(datapath_1_Instr_18_bF_buf22_), .C(_4440_), .Y(_4441_) );
NAND3X1 NAND3X1_81 ( .A(datapath_1_Instr_17_bF_buf30_), .B(_4441_), .C(_4438_), .Y(_4442_) );
INVX1 INVX1_41 ( .A(datapath_1_RegisterFile_regfile_mem_25__16_), .Y(_4443_) );
AOI21X1 AOI21X1_145 ( .A(datapath_1_RegisterFile_regfile_mem_29__16_), .B(datapath_1_Instr_18_bF_buf21_), .C(_3588__bF_buf15), .Y(_4444_) );
OAI21X1 OAI21X1_138 ( .A(_4443_), .B(datapath_1_Instr_18_bF_buf20_), .C(_4444_), .Y(_4445_) );
INVX1 INVX1_42 ( .A(datapath_1_RegisterFile_regfile_mem_24__16_), .Y(_4446_) );
AOI21X1 AOI21X1_146 ( .A(datapath_1_RegisterFile_regfile_mem_28__16_), .B(datapath_1_Instr_18_bF_buf19_), .C(datapath_1_Instr_16_bF_buf28_), .Y(_4447_) );
OAI21X1 OAI21X1_139 ( .A(_4446_), .B(datapath_1_Instr_18_bF_buf18_), .C(_4447_), .Y(_4448_) );
NAND3X1 NAND3X1_82 ( .A(_3566__bF_buf9), .B(_4448_), .C(_4445_), .Y(_4449_) );
AOI21X1 AOI21X1_147 ( .A(_4442_), .B(_4449_), .C(_3571__bF_buf7), .Y(_4450_) );
MUX2X1 MUX2X1_67 ( .A(datapath_1_RegisterFile_regfile_mem_18__16_), .B(datapath_1_RegisterFile_regfile_mem_16__16_), .S(datapath_1_Instr_17_bF_buf29_), .Y(_4451_) );
NAND2X1 NAND2X1_162 ( .A(_3588__bF_buf39), .B(_4451_), .Y(_4452_) );
MUX2X1 MUX2X1_68 ( .A(datapath_1_RegisterFile_regfile_mem_19__16_), .B(datapath_1_RegisterFile_regfile_mem_17__16_), .S(datapath_1_Instr_17_bF_buf28_), .Y(_4453_) );
NAND2X1 NAND2X1_163 ( .A(datapath_1_Instr_16_bF_buf27_), .B(_4453_), .Y(_4454_) );
NAND3X1 NAND3X1_83 ( .A(_3567__bF_buf2), .B(_4452_), .C(_4454_), .Y(_4455_) );
MUX2X1 MUX2X1_69 ( .A(datapath_1_RegisterFile_regfile_mem_22__16_), .B(datapath_1_RegisterFile_regfile_mem_20__16_), .S(datapath_1_Instr_17_bF_buf27_), .Y(_4456_) );
NAND2X1 NAND2X1_164 ( .A(_3588__bF_buf39), .B(_4456_), .Y(_4457_) );
MUX2X1 MUX2X1_70 ( .A(datapath_1_RegisterFile_regfile_mem_23__16_), .B(datapath_1_RegisterFile_regfile_mem_21__16_), .S(datapath_1_Instr_17_bF_buf26_), .Y(_4458_) );
NAND2X1 NAND2X1_165 ( .A(datapath_1_Instr_16_bF_buf26_), .B(_4458_), .Y(_4459_) );
NAND3X1 NAND3X1_84 ( .A(datapath_1_Instr_18_bF_buf17_), .B(_4457_), .C(_4459_), .Y(_4460_) );
AOI21X1 AOI21X1_148 ( .A(_4455_), .B(_4460_), .C(datapath_1_Instr_19_bF_buf0_), .Y(_4461_) );
OAI21X1 OAI21X1_140 ( .A(_4450_), .B(_4461_), .C(datapath_1_Instr_20_bF_buf3_), .Y(_4462_) );
AOI22X1 AOI22X1_26 ( .A(_3565__bF_buf0), .B(_3569__bF_buf0), .C(_4462_), .D(_4435_), .Y(datapath_1_RD2_16_) );
NAND2X1 NAND2X1_166 ( .A(datapath_1_RegisterFile_regfile_mem_27__17_), .B(datapath_1_Instr_16_bF_buf25_), .Y(_4463_) );
NAND2X1 NAND2X1_167 ( .A(datapath_1_RegisterFile_regfile_mem_26__17_), .B(_3588__bF_buf16), .Y(_4464_) );
NAND3X1 NAND3X1_85 ( .A(datapath_1_Instr_17_bF_buf25_), .B(_4463_), .C(_4464_), .Y(_4465_) );
NAND2X1 NAND2X1_168 ( .A(datapath_1_RegisterFile_regfile_mem_25__17_), .B(datapath_1_Instr_16_bF_buf24_), .Y(_4466_) );
AOI21X1 AOI21X1_149 ( .A(_3588__bF_buf16), .B(datapath_1_RegisterFile_regfile_mem_24__17_), .C(datapath_1_Instr_17_bF_buf24_), .Y(_4467_) );
NAND2X1 NAND2X1_169 ( .A(_4466_), .B(_4467_), .Y(_4468_) );
NAND3X1 NAND3X1_86 ( .A(_3567__bF_buf3), .B(_4465_), .C(_4468_), .Y(_4469_) );
NAND2X1 NAND2X1_170 ( .A(datapath_1_RegisterFile_regfile_mem_31__17_), .B(datapath_1_Instr_16_bF_buf23_), .Y(_4470_) );
AOI21X1 AOI21X1_150 ( .A(_3588__bF_buf37), .B(datapath_1_RegisterFile_regfile_mem_30__17_), .C(_3566__bF_buf4), .Y(_4471_) );
NAND2X1 NAND2X1_171 ( .A(_4470_), .B(_4471_), .Y(_4472_) );
INVX1 INVX1_43 ( .A(datapath_1_RegisterFile_regfile_mem_28__17_), .Y(_4473_) );
AOI21X1 AOI21X1_151 ( .A(datapath_1_RegisterFile_regfile_mem_29__17_), .B(datapath_1_Instr_16_bF_buf22_), .C(datapath_1_Instr_17_bF_buf23_), .Y(_4474_) );
OAI21X1 OAI21X1_141 ( .A(_4473_), .B(datapath_1_Instr_16_bF_buf21_), .C(_4474_), .Y(_4475_) );
NAND3X1 NAND3X1_87 ( .A(datapath_1_Instr_18_bF_buf16_), .B(_4475_), .C(_4472_), .Y(_4476_) );
AOI21X1 AOI21X1_152 ( .A(_4469_), .B(_4476_), .C(_3571__bF_buf5), .Y(_4477_) );
MUX2X1 MUX2X1_71 ( .A(datapath_1_RegisterFile_regfile_mem_17__17_), .B(datapath_1_RegisterFile_regfile_mem_16__17_), .S(datapath_1_Instr_16_bF_buf20_), .Y(_4478_) );
NOR2X1 NOR2X1_64 ( .A(datapath_1_RegisterFile_regfile_mem_19__17_), .B(_3588__bF_buf16), .Y(_4479_) );
OAI21X1 OAI21X1_142 ( .A(datapath_1_RegisterFile_regfile_mem_18__17_), .B(datapath_1_Instr_16_bF_buf19_), .C(datapath_1_Instr_17_bF_buf22_), .Y(_4480_) );
OAI22X1 OAI22X1_54 ( .A(_4480_), .B(_4479_), .C(datapath_1_Instr_17_bF_buf21_), .D(_4478_), .Y(_4481_) );
NAND2X1 NAND2X1_172 ( .A(_3567__bF_buf3), .B(_4481_), .Y(_4482_) );
MUX2X1 MUX2X1_72 ( .A(datapath_1_RegisterFile_regfile_mem_21__17_), .B(datapath_1_RegisterFile_regfile_mem_20__17_), .S(datapath_1_Instr_16_bF_buf18_), .Y(_4483_) );
NOR2X1 NOR2X1_65 ( .A(datapath_1_RegisterFile_regfile_mem_23__17_), .B(_3588__bF_buf16), .Y(_4484_) );
OAI21X1 OAI21X1_143 ( .A(datapath_1_RegisterFile_regfile_mem_22__17_), .B(datapath_1_Instr_16_bF_buf17_), .C(datapath_1_Instr_17_bF_buf20_), .Y(_4485_) );
OAI22X1 OAI22X1_55 ( .A(_4485_), .B(_4484_), .C(datapath_1_Instr_17_bF_buf19_), .D(_4483_), .Y(_4486_) );
NAND2X1 NAND2X1_173 ( .A(datapath_1_Instr_18_bF_buf15_), .B(_4486_), .Y(_4487_) );
AOI21X1 AOI21X1_153 ( .A(_4482_), .B(_4487_), .C(datapath_1_Instr_19_bF_buf6_), .Y(_4488_) );
OAI21X1 OAI21X1_144 ( .A(_4477_), .B(_4488_), .C(datapath_1_Instr_20_bF_buf2_), .Y(_4489_) );
NAND2X1 NAND2X1_174 ( .A(datapath_1_RegisterFile_regfile_mem_11__17_), .B(datapath_1_Instr_17_bF_buf18_), .Y(_4490_) );
NAND2X1 NAND2X1_175 ( .A(datapath_1_RegisterFile_regfile_mem_9__17_), .B(_3566__bF_buf8), .Y(_4491_) );
NAND3X1 NAND3X1_88 ( .A(datapath_1_Instr_16_bF_buf16_), .B(_4490_), .C(_4491_), .Y(_4492_) );
NAND2X1 NAND2X1_176 ( .A(datapath_1_RegisterFile_regfile_mem_10__17_), .B(datapath_1_Instr_17_bF_buf17_), .Y(_4493_) );
AOI21X1 AOI21X1_154 ( .A(_3566__bF_buf8), .B(datapath_1_RegisterFile_regfile_mem_8__17_), .C(datapath_1_Instr_16_bF_buf15_), .Y(_4494_) );
NAND2X1 NAND2X1_177 ( .A(_4493_), .B(_4494_), .Y(_4495_) );
NAND3X1 NAND3X1_89 ( .A(_3567__bF_buf8), .B(_4492_), .C(_4495_), .Y(_4496_) );
NAND2X1 NAND2X1_178 ( .A(datapath_1_RegisterFile_regfile_mem_15__17_), .B(datapath_1_Instr_17_bF_buf16_), .Y(_4497_) );
NAND2X1 NAND2X1_179 ( .A(datapath_1_RegisterFile_regfile_mem_13__17_), .B(_3566__bF_buf8), .Y(_4498_) );
NAND3X1 NAND3X1_90 ( .A(datapath_1_Instr_16_bF_buf14_), .B(_4497_), .C(_4498_), .Y(_4499_) );
NAND2X1 NAND2X1_180 ( .A(datapath_1_RegisterFile_regfile_mem_14__17_), .B(datapath_1_Instr_17_bF_buf15_), .Y(_4500_) );
AOI21X1 AOI21X1_155 ( .A(_3566__bF_buf8), .B(datapath_1_RegisterFile_regfile_mem_12__17_), .C(datapath_1_Instr_16_bF_buf13_), .Y(_4501_) );
NAND2X1 NAND2X1_181 ( .A(_4500_), .B(_4501_), .Y(_4502_) );
NAND3X1 NAND3X1_91 ( .A(datapath_1_Instr_18_bF_buf14_), .B(_4499_), .C(_4502_), .Y(_4503_) );
AOI21X1 AOI21X1_156 ( .A(_4496_), .B(_4503_), .C(_3571__bF_buf3), .Y(_4504_) );
INVX1 INVX1_44 ( .A(datapath_1_RegisterFile_regfile_mem_1__17_), .Y(_4505_) );
AOI21X1 AOI21X1_157 ( .A(datapath_1_RegisterFile_regfile_mem_5__17_), .B(datapath_1_Instr_18_bF_buf13_), .C(_3588__bF_buf18), .Y(_4506_) );
OAI21X1 OAI21X1_145 ( .A(_4505_), .B(datapath_1_Instr_18_bF_buf12_), .C(_4506_), .Y(_4507_) );
INVX1 INVX1_45 ( .A(datapath_1_RegisterFile_regfile_mem_0__17_), .Y(_4508_) );
AOI21X1 AOI21X1_158 ( .A(datapath_1_RegisterFile_regfile_mem_4__17_), .B(datapath_1_Instr_18_bF_buf11_), .C(datapath_1_Instr_16_bF_buf12_), .Y(_4509_) );
OAI21X1 OAI21X1_146 ( .A(_4508_), .B(datapath_1_Instr_18_bF_buf10_), .C(_4509_), .Y(_4510_) );
NAND3X1 NAND3X1_92 ( .A(_3566__bF_buf4), .B(_4510_), .C(_4507_), .Y(_4511_) );
INVX1 INVX1_46 ( .A(datapath_1_RegisterFile_regfile_mem_3__17_), .Y(_4512_) );
AOI21X1 AOI21X1_159 ( .A(datapath_1_RegisterFile_regfile_mem_7__17_), .B(datapath_1_Instr_18_bF_buf9_), .C(_3588__bF_buf18), .Y(_4513_) );
OAI21X1 OAI21X1_147 ( .A(_4512_), .B(datapath_1_Instr_18_bF_buf8_), .C(_4513_), .Y(_4514_) );
INVX1 INVX1_47 ( .A(datapath_1_RegisterFile_regfile_mem_2__17_), .Y(_4515_) );
AOI21X1 AOI21X1_160 ( .A(datapath_1_RegisterFile_regfile_mem_6__17_), .B(datapath_1_Instr_18_bF_buf7_), .C(datapath_1_Instr_16_bF_buf11_), .Y(_4516_) );
OAI21X1 OAI21X1_148 ( .A(_4515_), .B(datapath_1_Instr_18_bF_buf6_), .C(_4516_), .Y(_4517_) );
NAND3X1 NAND3X1_93 ( .A(datapath_1_Instr_17_bF_buf14_), .B(_4517_), .C(_4514_), .Y(_4518_) );
AOI21X1 AOI21X1_161 ( .A(_4511_), .B(_4518_), .C(datapath_1_Instr_19_bF_buf5_), .Y(_4519_) );
OAI21X1 OAI21X1_149 ( .A(_4519_), .B(_4504_), .C(_3570__bF_buf0), .Y(_4520_) );
AOI22X1 AOI22X1_27 ( .A(_3565__bF_buf2), .B(_3569__bF_buf2), .C(_4520_), .D(_4489_), .Y(datapath_1_RD2_17_) );
MUX2X1 MUX2X1_73 ( .A(datapath_1_RegisterFile_regfile_mem_9__18_), .B(datapath_1_RegisterFile_regfile_mem_8__18_), .S(datapath_1_Instr_16_bF_buf10_), .Y(_4521_) );
NOR2X1 NOR2X1_66 ( .A(datapath_1_RegisterFile_regfile_mem_11__18_), .B(_3588__bF_buf4), .Y(_4522_) );
OAI21X1 OAI21X1_150 ( .A(datapath_1_RegisterFile_regfile_mem_10__18_), .B(datapath_1_Instr_16_bF_buf9_), .C(datapath_1_Instr_17_bF_buf13_), .Y(_4523_) );
OAI22X1 OAI22X1_56 ( .A(_4523_), .B(_4522_), .C(datapath_1_Instr_17_bF_buf12_), .D(_4521_), .Y(_4524_) );
INVX1 INVX1_48 ( .A(datapath_1_RegisterFile_regfile_mem_15__18_), .Y(_4525_) );
AOI21X1 AOI21X1_162 ( .A(_3588__bF_buf4), .B(datapath_1_RegisterFile_regfile_mem_14__18_), .C(_3566__bF_buf3), .Y(_4526_) );
OAI21X1 OAI21X1_151 ( .A(_4525_), .B(_3588__bF_buf4), .C(_4526_), .Y(_4527_) );
NAND2X1 NAND2X1_182 ( .A(datapath_1_RegisterFile_regfile_mem_12__18_), .B(_3588__bF_buf35), .Y(_4528_) );
AOI21X1 AOI21X1_163 ( .A(datapath_1_RegisterFile_regfile_mem_13__18_), .B(datapath_1_Instr_16_bF_buf8_), .C(datapath_1_Instr_17_bF_buf11_), .Y(_4529_) );
AOI21X1 AOI21X1_164 ( .A(_4528_), .B(_4529_), .C(_3567__bF_buf6), .Y(_4530_) );
AOI22X1 AOI22X1_28 ( .A(_4527_), .B(_4530_), .C(_3567__bF_buf6), .D(_4524_), .Y(_4531_) );
NOR2X1 NOR2X1_67 ( .A(datapath_1_RegisterFile_regfile_mem_0__18_), .B(datapath_1_Instr_16_bF_buf7_), .Y(_4532_) );
OAI21X1 OAI21X1_152 ( .A(datapath_1_RegisterFile_regfile_mem_1__18_), .B(_3588__bF_buf30), .C(_3566__bF_buf6), .Y(_4533_) );
NOR2X1 NOR2X1_68 ( .A(datapath_1_RegisterFile_regfile_mem_3__18_), .B(_3588__bF_buf30), .Y(_4534_) );
OAI21X1 OAI21X1_153 ( .A(datapath_1_RegisterFile_regfile_mem_2__18_), .B(datapath_1_Instr_16_bF_buf6_), .C(datapath_1_Instr_17_bF_buf10_), .Y(_4535_) );
OAI22X1 OAI22X1_57 ( .A(_4534_), .B(_4535_), .C(_4532_), .D(_4533_), .Y(_4536_) );
NOR2X1 NOR2X1_69 ( .A(datapath_1_Instr_18_bF_buf5_), .B(_4536_), .Y(_4537_) );
MUX2X1 MUX2X1_74 ( .A(datapath_1_RegisterFile_regfile_mem_5__18_), .B(datapath_1_RegisterFile_regfile_mem_4__18_), .S(datapath_1_Instr_16_bF_buf5_), .Y(_4538_) );
NOR2X1 NOR2X1_70 ( .A(datapath_1_RegisterFile_regfile_mem_7__18_), .B(_3588__bF_buf4), .Y(_4539_) );
OAI21X1 OAI21X1_154 ( .A(datapath_1_RegisterFile_regfile_mem_6__18_), .B(datapath_1_Instr_16_bF_buf4_), .C(datapath_1_Instr_17_bF_buf9_), .Y(_4540_) );
OAI22X1 OAI22X1_58 ( .A(_4540_), .B(_4539_), .C(datapath_1_Instr_17_bF_buf8_), .D(_4538_), .Y(_4541_) );
OAI21X1 OAI21X1_155 ( .A(_3567__bF_buf1), .B(_4541_), .C(_3571__bF_buf2), .Y(_4542_) );
OAI22X1 OAI22X1_59 ( .A(_3571__bF_buf2), .B(_4531_), .C(_4537_), .D(_4542_), .Y(_4543_) );
NAND2X1 NAND2X1_183 ( .A(_3570__bF_buf0), .B(_4543_), .Y(_4544_) );
INVX1 INVX1_49 ( .A(datapath_1_RegisterFile_regfile_mem_19__18_), .Y(_4545_) );
AOI21X1 AOI21X1_165 ( .A(datapath_1_RegisterFile_regfile_mem_23__18_), .B(datapath_1_Instr_18_bF_buf4_), .C(_3588__bF_buf27), .Y(_4546_) );
OAI21X1 OAI21X1_156 ( .A(_4545_), .B(datapath_1_Instr_18_bF_buf3_), .C(_4546_), .Y(_4547_) );
NAND2X1 NAND2X1_184 ( .A(datapath_1_RegisterFile_regfile_mem_18__18_), .B(_3567__bF_buf9), .Y(_4548_) );
AOI21X1 AOI21X1_166 ( .A(datapath_1_RegisterFile_regfile_mem_22__18_), .B(datapath_1_Instr_18_bF_buf2_), .C(datapath_1_Instr_16_bF_buf3_), .Y(_4549_) );
AOI21X1 AOI21X1_167 ( .A(_4548_), .B(_4549_), .C(_3566__bF_buf6), .Y(_4550_) );
INVX1 INVX1_50 ( .A(datapath_1_RegisterFile_regfile_mem_17__18_), .Y(_4551_) );
AOI21X1 AOI21X1_168 ( .A(datapath_1_RegisterFile_regfile_mem_21__18_), .B(datapath_1_Instr_18_bF_buf1_), .C(_3588__bF_buf32), .Y(_4552_) );
OAI21X1 OAI21X1_157 ( .A(_4551_), .B(datapath_1_Instr_18_bF_buf0_), .C(_4552_), .Y(_4553_) );
NAND2X1 NAND2X1_185 ( .A(datapath_1_RegisterFile_regfile_mem_16__18_), .B(_3567__bF_buf9), .Y(_4554_) );
AOI21X1 AOI21X1_169 ( .A(datapath_1_RegisterFile_regfile_mem_20__18_), .B(datapath_1_Instr_18_bF_buf44_), .C(datapath_1_Instr_16_bF_buf2_), .Y(_4555_) );
AOI21X1 AOI21X1_170 ( .A(_4554_), .B(_4555_), .C(datapath_1_Instr_17_bF_buf7_), .Y(_4556_) );
AOI22X1 AOI22X1_29 ( .A(_4550_), .B(_4547_), .C(_4553_), .D(_4556_), .Y(_4557_) );
NOR2X1 NOR2X1_71 ( .A(datapath_1_RegisterFile_regfile_mem_24__18_), .B(datapath_1_Instr_16_bF_buf1_), .Y(_4558_) );
OAI21X1 OAI21X1_158 ( .A(datapath_1_RegisterFile_regfile_mem_25__18_), .B(_3588__bF_buf23), .C(_3566__bF_buf6), .Y(_4559_) );
NOR2X1 NOR2X1_72 ( .A(datapath_1_RegisterFile_regfile_mem_27__18_), .B(_3588__bF_buf23), .Y(_4560_) );
OAI21X1 OAI21X1_159 ( .A(datapath_1_RegisterFile_regfile_mem_26__18_), .B(datapath_1_Instr_16_bF_buf0_), .C(datapath_1_Instr_17_bF_buf6_), .Y(_4561_) );
OAI22X1 OAI22X1_60 ( .A(_4560_), .B(_4561_), .C(_4558_), .D(_4559_), .Y(_4562_) );
NOR2X1 NOR2X1_73 ( .A(datapath_1_Instr_18_bF_buf43_), .B(_4562_), .Y(_4563_) );
MUX2X1 MUX2X1_75 ( .A(datapath_1_RegisterFile_regfile_mem_29__18_), .B(datapath_1_RegisterFile_regfile_mem_28__18_), .S(datapath_1_Instr_16_bF_buf55_), .Y(_4564_) );
NOR2X1 NOR2X1_74 ( .A(datapath_1_RegisterFile_regfile_mem_31__18_), .B(_3588__bF_buf20), .Y(_4565_) );
OAI21X1 OAI21X1_160 ( .A(datapath_1_RegisterFile_regfile_mem_30__18_), .B(datapath_1_Instr_16_bF_buf54_), .C(datapath_1_Instr_17_bF_buf5_), .Y(_4566_) );
OAI22X1 OAI22X1_61 ( .A(_4566_), .B(_4565_), .C(datapath_1_Instr_17_bF_buf4_), .D(_4564_), .Y(_4567_) );
OAI21X1 OAI21X1_161 ( .A(_3567__bF_buf9), .B(_4567_), .C(datapath_1_Instr_19_bF_buf4_), .Y(_4568_) );
OAI22X1 OAI22X1_62 ( .A(datapath_1_Instr_19_bF_buf3_), .B(_4557_), .C(_4563_), .D(_4568_), .Y(_4569_) );
NAND2X1 NAND2X1_186 ( .A(datapath_1_Instr_20_bF_buf1_), .B(_4569_), .Y(_4570_) );
AOI22X1 AOI22X1_30 ( .A(_3565__bF_buf2), .B(_3569__bF_buf2), .C(_4570_), .D(_4544_), .Y(datapath_1_RD2_18_) );
MUX2X1 MUX2X1_76 ( .A(datapath_1_RegisterFile_regfile_mem_2__19_), .B(datapath_1_RegisterFile_regfile_mem_0__19_), .S(datapath_1_Instr_17_bF_buf3_), .Y(_4571_) );
NAND2X1 NAND2X1_187 ( .A(_3588__bF_buf36), .B(_4571_), .Y(_4572_) );
MUX2X1 MUX2X1_77 ( .A(datapath_1_RegisterFile_regfile_mem_3__19_), .B(datapath_1_RegisterFile_regfile_mem_1__19_), .S(datapath_1_Instr_17_bF_buf2_), .Y(_4573_) );
NAND2X1 NAND2X1_188 ( .A(datapath_1_Instr_16_bF_buf53_), .B(_4573_), .Y(_4574_) );
NAND3X1 NAND3X1_94 ( .A(_3567__bF_buf7), .B(_4572_), .C(_4574_), .Y(_4575_) );
MUX2X1 MUX2X1_78 ( .A(datapath_1_RegisterFile_regfile_mem_6__19_), .B(datapath_1_RegisterFile_regfile_mem_4__19_), .S(datapath_1_Instr_17_bF_buf1_), .Y(_4576_) );
NAND2X1 NAND2X1_189 ( .A(_3588__bF_buf11), .B(_4576_), .Y(_4577_) );
MUX2X1 MUX2X1_79 ( .A(datapath_1_RegisterFile_regfile_mem_7__19_), .B(datapath_1_RegisterFile_regfile_mem_5__19_), .S(datapath_1_Instr_17_bF_buf0_), .Y(_4578_) );
NAND2X1 NAND2X1_190 ( .A(datapath_1_Instr_16_bF_buf52_), .B(_4578_), .Y(_4579_) );
NAND3X1 NAND3X1_95 ( .A(datapath_1_Instr_18_bF_buf42_), .B(_4577_), .C(_4579_), .Y(_4580_) );
AOI21X1 AOI21X1_171 ( .A(_4575_), .B(_4580_), .C(datapath_1_Instr_19_bF_buf2_), .Y(_4581_) );
INVX1 INVX1_51 ( .A(datapath_1_RegisterFile_regfile_mem_9__19_), .Y(_4582_) );
AOI21X1 AOI21X1_172 ( .A(datapath_1_RegisterFile_regfile_mem_13__19_), .B(datapath_1_Instr_18_bF_buf41_), .C(_3588__bF_buf13), .Y(_4583_) );
OAI21X1 OAI21X1_162 ( .A(_4582_), .B(datapath_1_Instr_18_bF_buf40_), .C(_4583_), .Y(_4584_) );
INVX1 INVX1_52 ( .A(datapath_1_RegisterFile_regfile_mem_8__19_), .Y(_4585_) );
AOI21X1 AOI21X1_173 ( .A(datapath_1_RegisterFile_regfile_mem_12__19_), .B(datapath_1_Instr_18_bF_buf39_), .C(datapath_1_Instr_16_bF_buf51_), .Y(_4586_) );
OAI21X1 OAI21X1_163 ( .A(_4585_), .B(datapath_1_Instr_18_bF_buf38_), .C(_4586_), .Y(_4587_) );
NAND3X1 NAND3X1_96 ( .A(_3566__bF_buf9), .B(_4587_), .C(_4584_), .Y(_4588_) );
INVX1 INVX1_53 ( .A(datapath_1_RegisterFile_regfile_mem_11__19_), .Y(_4589_) );
AOI21X1 AOI21X1_174 ( .A(datapath_1_RegisterFile_regfile_mem_15__19_), .B(datapath_1_Instr_18_bF_buf37_), .C(_3588__bF_buf36), .Y(_4590_) );
OAI21X1 OAI21X1_164 ( .A(_4589_), .B(datapath_1_Instr_18_bF_buf36_), .C(_4590_), .Y(_4591_) );
INVX1 INVX1_54 ( .A(datapath_1_RegisterFile_regfile_mem_10__19_), .Y(_4592_) );
AOI21X1 AOI21X1_175 ( .A(datapath_1_RegisterFile_regfile_mem_14__19_), .B(datapath_1_Instr_18_bF_buf35_), .C(datapath_1_Instr_16_bF_buf50_), .Y(_4593_) );
OAI21X1 OAI21X1_165 ( .A(_4592_), .B(datapath_1_Instr_18_bF_buf34_), .C(_4593_), .Y(_4594_) );
NAND3X1 NAND3X1_97 ( .A(datapath_1_Instr_17_bF_buf50_), .B(_4594_), .C(_4591_), .Y(_4595_) );
AOI21X1 AOI21X1_176 ( .A(_4588_), .B(_4595_), .C(_3571__bF_buf4), .Y(_4596_) );
OAI21X1 OAI21X1_166 ( .A(_4596_), .B(_4581_), .C(_3570__bF_buf2), .Y(_4597_) );
NOR2X1 NOR2X1_75 ( .A(datapath_1_RegisterFile_regfile_mem_24__19_), .B(datapath_1_Instr_16_bF_buf49_), .Y(_4598_) );
OAI21X1 OAI21X1_167 ( .A(datapath_1_RegisterFile_regfile_mem_25__19_), .B(_3588__bF_buf6), .C(_3566__bF_buf10), .Y(_4599_) );
NOR2X1 NOR2X1_76 ( .A(datapath_1_RegisterFile_regfile_mem_27__19_), .B(_3588__bF_buf33), .Y(_4600_) );
OAI21X1 OAI21X1_168 ( .A(datapath_1_RegisterFile_regfile_mem_26__19_), .B(datapath_1_Instr_16_bF_buf48_), .C(datapath_1_Instr_17_bF_buf49_), .Y(_4601_) );
OAI22X1 OAI22X1_63 ( .A(_4600_), .B(_4601_), .C(_4598_), .D(_4599_), .Y(_4602_) );
NOR2X1 NOR2X1_77 ( .A(datapath_1_Instr_18_bF_buf33_), .B(_4602_), .Y(_4603_) );
MUX2X1 MUX2X1_80 ( .A(datapath_1_RegisterFile_regfile_mem_29__19_), .B(datapath_1_RegisterFile_regfile_mem_28__19_), .S(datapath_1_Instr_16_bF_buf47_), .Y(_4604_) );
NOR2X1 NOR2X1_78 ( .A(datapath_1_RegisterFile_regfile_mem_31__19_), .B(_3588__bF_buf31), .Y(_4605_) );
OAI21X1 OAI21X1_169 ( .A(datapath_1_RegisterFile_regfile_mem_30__19_), .B(datapath_1_Instr_16_bF_buf46_), .C(datapath_1_Instr_17_bF_buf48_), .Y(_4606_) );
OAI22X1 OAI22X1_64 ( .A(_4606_), .B(_4605_), .C(datapath_1_Instr_17_bF_buf47_), .D(_4604_), .Y(_4607_) );
OAI21X1 OAI21X1_170 ( .A(_3567__bF_buf5), .B(_4607_), .C(datapath_1_Instr_19_bF_buf1_), .Y(_4608_) );
INVX1 INVX1_55 ( .A(datapath_1_RegisterFile_regfile_mem_19__19_), .Y(_4609_) );
AOI21X1 AOI21X1_177 ( .A(datapath_1_RegisterFile_regfile_mem_23__19_), .B(datapath_1_Instr_18_bF_buf32_), .C(_3588__bF_buf26), .Y(_4610_) );
OAI21X1 OAI21X1_171 ( .A(_4609_), .B(datapath_1_Instr_18_bF_buf31_), .C(_4610_), .Y(_4611_) );
NAND2X1 NAND2X1_191 ( .A(datapath_1_RegisterFile_regfile_mem_18__19_), .B(_3567__bF_buf0), .Y(_4612_) );
AOI21X1 AOI21X1_178 ( .A(datapath_1_RegisterFile_regfile_mem_22__19_), .B(datapath_1_Instr_18_bF_buf30_), .C(datapath_1_Instr_16_bF_buf45_), .Y(_4613_) );
AOI21X1 AOI21X1_179 ( .A(_4612_), .B(_4613_), .C(_3566__bF_buf9), .Y(_4614_) );
INVX1 INVX1_56 ( .A(datapath_1_RegisterFile_regfile_mem_17__19_), .Y(_4615_) );
AOI21X1 AOI21X1_180 ( .A(datapath_1_RegisterFile_regfile_mem_21__19_), .B(datapath_1_Instr_18_bF_buf29_), .C(_3588__bF_buf14), .Y(_4616_) );
OAI21X1 OAI21X1_172 ( .A(_4615_), .B(datapath_1_Instr_18_bF_buf28_), .C(_4616_), .Y(_4617_) );
NAND2X1 NAND2X1_192 ( .A(datapath_1_RegisterFile_regfile_mem_16__19_), .B(_3567__bF_buf5), .Y(_4618_) );
AOI21X1 AOI21X1_181 ( .A(datapath_1_RegisterFile_regfile_mem_20__19_), .B(datapath_1_Instr_18_bF_buf27_), .C(datapath_1_Instr_16_bF_buf44_), .Y(_4619_) );
AOI21X1 AOI21X1_182 ( .A(_4618_), .B(_4619_), .C(datapath_1_Instr_17_bF_buf46_), .Y(_4620_) );
AOI22X1 AOI22X1_31 ( .A(_4614_), .B(_4611_), .C(_4617_), .D(_4620_), .Y(_4621_) );
OAI22X1 OAI22X1_65 ( .A(datapath_1_Instr_19_bF_buf0_), .B(_4621_), .C(_4603_), .D(_4608_), .Y(_4622_) );
NAND2X1 NAND2X1_193 ( .A(datapath_1_Instr_20_bF_buf0_), .B(_4622_), .Y(_4623_) );
AOI22X1 AOI22X1_32 ( .A(_3565__bF_buf1), .B(_3569__bF_buf1), .C(_4597_), .D(_4623_), .Y(datapath_1_RD2_19_) );
NAND2X1 NAND2X1_194 ( .A(datapath_1_RegisterFile_regfile_mem_27__20_), .B(datapath_1_Instr_16_bF_buf43_), .Y(_4624_) );
NAND2X1 NAND2X1_195 ( .A(datapath_1_RegisterFile_regfile_mem_26__20_), .B(_3588__bF_buf0), .Y(_4625_) );
NAND3X1 NAND3X1_98 ( .A(datapath_1_Instr_17_bF_buf45_), .B(_4624_), .C(_4625_), .Y(_4626_) );
NAND2X1 NAND2X1_196 ( .A(datapath_1_RegisterFile_regfile_mem_25__20_), .B(datapath_1_Instr_16_bF_buf42_), .Y(_4627_) );
AOI21X1 AOI21X1_183 ( .A(_3588__bF_buf28), .B(datapath_1_RegisterFile_regfile_mem_24__20_), .C(datapath_1_Instr_17_bF_buf44_), .Y(_4628_) );
NAND2X1 NAND2X1_197 ( .A(_4627_), .B(_4628_), .Y(_4629_) );
NAND3X1 NAND3X1_99 ( .A(_3567__bF_buf10), .B(_4626_), .C(_4629_), .Y(_4630_) );
NAND2X1 NAND2X1_198 ( .A(datapath_1_RegisterFile_regfile_mem_31__20_), .B(datapath_1_Instr_16_bF_buf41_), .Y(_4631_) );
AOI21X1 AOI21X1_184 ( .A(_3588__bF_buf28), .B(datapath_1_RegisterFile_regfile_mem_30__20_), .C(_3566__bF_buf9), .Y(_4632_) );
NAND2X1 NAND2X1_199 ( .A(_4631_), .B(_4632_), .Y(_4633_) );
AOI21X1 AOI21X1_185 ( .A(datapath_1_RegisterFile_regfile_mem_29__20_), .B(datapath_1_Instr_16_bF_buf40_), .C(datapath_1_Instr_17_bF_buf43_), .Y(_4634_) );
OAI21X1 OAI21X1_173 ( .A(_2952_), .B(datapath_1_Instr_16_bF_buf39_), .C(_4634_), .Y(_4635_) );
NAND3X1 NAND3X1_100 ( .A(datapath_1_Instr_18_bF_buf26_), .B(_4635_), .C(_4633_), .Y(_4636_) );
AOI21X1 AOI21X1_186 ( .A(_4630_), .B(_4636_), .C(_3571__bF_buf4), .Y(_4637_) );
MUX2X1 MUX2X1_81 ( .A(datapath_1_RegisterFile_regfile_mem_18__20_), .B(datapath_1_RegisterFile_regfile_mem_16__20_), .S(datapath_1_Instr_17_bF_buf42_), .Y(_4638_) );
NAND2X1 NAND2X1_200 ( .A(_3588__bF_buf19), .B(_4638_), .Y(_4639_) );
MUX2X1 MUX2X1_82 ( .A(datapath_1_RegisterFile_regfile_mem_19__20_), .B(datapath_1_RegisterFile_regfile_mem_17__20_), .S(datapath_1_Instr_17_bF_buf41_), .Y(_4640_) );
NAND2X1 NAND2X1_201 ( .A(datapath_1_Instr_16_bF_buf38_), .B(_4640_), .Y(_4641_) );
NAND3X1 NAND3X1_101 ( .A(_3567__bF_buf5), .B(_4639_), .C(_4641_), .Y(_4642_) );
MUX2X1 MUX2X1_83 ( .A(datapath_1_RegisterFile_regfile_mem_22__20_), .B(datapath_1_RegisterFile_regfile_mem_20__20_), .S(datapath_1_Instr_17_bF_buf40_), .Y(_4643_) );
NAND2X1 NAND2X1_202 ( .A(_3588__bF_buf19), .B(_4643_), .Y(_4644_) );
MUX2X1 MUX2X1_84 ( .A(datapath_1_RegisterFile_regfile_mem_23__20_), .B(datapath_1_RegisterFile_regfile_mem_21__20_), .S(datapath_1_Instr_17_bF_buf39_), .Y(_4645_) );
NAND2X1 NAND2X1_203 ( .A(datapath_1_Instr_16_bF_buf37_), .B(_4645_), .Y(_4646_) );
NAND3X1 NAND3X1_102 ( .A(datapath_1_Instr_18_bF_buf25_), .B(_4644_), .C(_4646_), .Y(_4647_) );
AOI21X1 AOI21X1_187 ( .A(_4642_), .B(_4647_), .C(datapath_1_Instr_19_bF_buf6_), .Y(_4648_) );
OAI21X1 OAI21X1_174 ( .A(_4648_), .B(_4637_), .C(datapath_1_Instr_20_bF_buf5_), .Y(_4649_) );
MUX2X1 MUX2X1_85 ( .A(datapath_1_RegisterFile_regfile_mem_9__20_), .B(datapath_1_RegisterFile_regfile_mem_8__20_), .S(datapath_1_Instr_16_bF_buf36_), .Y(_4650_) );
NOR2X1 NOR2X1_79 ( .A(datapath_1_RegisterFile_regfile_mem_11__20_), .B(_3588__bF_buf40), .Y(_4651_) );
OAI21X1 OAI21X1_175 ( .A(datapath_1_RegisterFile_regfile_mem_10__20_), .B(datapath_1_Instr_16_bF_buf35_), .C(datapath_1_Instr_17_bF_buf38_), .Y(_4652_) );
OAI22X1 OAI22X1_66 ( .A(_4652_), .B(_4651_), .C(datapath_1_Instr_17_bF_buf37_), .D(_4650_), .Y(_4653_) );
AOI21X1 AOI21X1_188 ( .A(_3588__bF_buf40), .B(datapath_1_RegisterFile_regfile_mem_14__20_), .C(_3566__bF_buf1), .Y(_4654_) );
OAI21X1 OAI21X1_176 ( .A(_2973_), .B(_3588__bF_buf40), .C(_4654_), .Y(_4655_) );
NAND2X1 NAND2X1_204 ( .A(datapath_1_RegisterFile_regfile_mem_12__20_), .B(_3588__bF_buf40), .Y(_4656_) );
AOI21X1 AOI21X1_189 ( .A(datapath_1_RegisterFile_regfile_mem_13__20_), .B(datapath_1_Instr_16_bF_buf34_), .C(datapath_1_Instr_17_bF_buf36_), .Y(_4657_) );
AOI21X1 AOI21X1_190 ( .A(_4656_), .B(_4657_), .C(_3567__bF_buf7), .Y(_4658_) );
AOI22X1 AOI22X1_33 ( .A(_4655_), .B(_4658_), .C(_3567__bF_buf7), .D(_4653_), .Y(_4659_) );
NOR2X1 NOR2X1_80 ( .A(datapath_1_RegisterFile_regfile_mem_0__20_), .B(datapath_1_Instr_16_bF_buf33_), .Y(_4660_) );
OAI21X1 OAI21X1_177 ( .A(datapath_1_RegisterFile_regfile_mem_1__20_), .B(_3588__bF_buf36), .C(_3566__bF_buf1), .Y(_4661_) );
NOR2X1 NOR2X1_81 ( .A(datapath_1_RegisterFile_regfile_mem_3__20_), .B(_3588__bF_buf40), .Y(_4662_) );
OAI21X1 OAI21X1_178 ( .A(datapath_1_RegisterFile_regfile_mem_2__20_), .B(datapath_1_Instr_16_bF_buf32_), .C(datapath_1_Instr_17_bF_buf35_), .Y(_4663_) );
OAI22X1 OAI22X1_67 ( .A(_4662_), .B(_4663_), .C(_4660_), .D(_4661_), .Y(_4664_) );
NOR2X1 NOR2X1_82 ( .A(datapath_1_Instr_18_bF_buf24_), .B(_4664_), .Y(_4665_) );
MUX2X1 MUX2X1_86 ( .A(datapath_1_RegisterFile_regfile_mem_5__20_), .B(datapath_1_RegisterFile_regfile_mem_4__20_), .S(datapath_1_Instr_16_bF_buf31_), .Y(_4666_) );
NOR2X1 NOR2X1_83 ( .A(datapath_1_RegisterFile_regfile_mem_7__20_), .B(_3588__bF_buf42), .Y(_4667_) );
OAI21X1 OAI21X1_179 ( .A(datapath_1_RegisterFile_regfile_mem_6__20_), .B(datapath_1_Instr_16_bF_buf30_), .C(datapath_1_Instr_17_bF_buf34_), .Y(_4668_) );
OAI22X1 OAI22X1_68 ( .A(_4668_), .B(_4667_), .C(datapath_1_Instr_17_bF_buf33_), .D(_4666_), .Y(_4669_) );
OAI21X1 OAI21X1_180 ( .A(_3567__bF_buf4), .B(_4669_), .C(_3571__bF_buf0), .Y(_4670_) );
OAI22X1 OAI22X1_69 ( .A(_3571__bF_buf4), .B(_4659_), .C(_4665_), .D(_4670_), .Y(_4671_) );
NAND2X1 NAND2X1_205 ( .A(_3570__bF_buf2), .B(_4671_), .Y(_4672_) );
AOI22X1 AOI22X1_34 ( .A(_3565__bF_buf1), .B(_3569__bF_buf1), .C(_4649_), .D(_4672_), .Y(datapath_1_RD2_20_) );
INVX1 INVX1_57 ( .A(datapath_1_RegisterFile_regfile_mem_1__21_), .Y(_4673_) );
AOI21X1 AOI21X1_191 ( .A(datapath_1_RegisterFile_regfile_mem_5__21_), .B(datapath_1_Instr_18_bF_buf23_), .C(_3588__bF_buf5), .Y(_4674_) );
OAI21X1 OAI21X1_181 ( .A(_4673_), .B(datapath_1_Instr_18_bF_buf22_), .C(_4674_), .Y(_4675_) );
INVX1 INVX1_58 ( .A(datapath_1_RegisterFile_regfile_mem_0__21_), .Y(_4676_) );
AOI21X1 AOI21X1_192 ( .A(datapath_1_RegisterFile_regfile_mem_4__21_), .B(datapath_1_Instr_18_bF_buf21_), .C(datapath_1_Instr_16_bF_buf29_), .Y(_4677_) );
OAI21X1 OAI21X1_182 ( .A(_4676_), .B(datapath_1_Instr_18_bF_buf20_), .C(_4677_), .Y(_4678_) );
NAND3X1 NAND3X1_103 ( .A(_3566__bF_buf10), .B(_4678_), .C(_4675_), .Y(_4679_) );
INVX1 INVX1_59 ( .A(datapath_1_RegisterFile_regfile_mem_3__21_), .Y(_4680_) );
AOI21X1 AOI21X1_193 ( .A(datapath_1_RegisterFile_regfile_mem_7__21_), .B(datapath_1_Instr_18_bF_buf19_), .C(_3588__bF_buf9), .Y(_4681_) );
OAI21X1 OAI21X1_183 ( .A(_4680_), .B(datapath_1_Instr_18_bF_buf18_), .C(_4681_), .Y(_4682_) );
INVX1 INVX1_60 ( .A(datapath_1_RegisterFile_regfile_mem_2__21_), .Y(_4683_) );
AOI21X1 AOI21X1_194 ( .A(datapath_1_RegisterFile_regfile_mem_6__21_), .B(datapath_1_Instr_18_bF_buf17_), .C(datapath_1_Instr_16_bF_buf28_), .Y(_4684_) );
OAI21X1 OAI21X1_184 ( .A(_4683_), .B(datapath_1_Instr_18_bF_buf16_), .C(_4684_), .Y(_4685_) );
NAND3X1 NAND3X1_104 ( .A(datapath_1_Instr_17_bF_buf32_), .B(_4685_), .C(_4682_), .Y(_4686_) );
AOI21X1 AOI21X1_195 ( .A(_4679_), .B(_4686_), .C(datapath_1_Instr_19_bF_buf5_), .Y(_4687_) );
NAND2X1 NAND2X1_206 ( .A(datapath_1_RegisterFile_regfile_mem_11__21_), .B(datapath_1_Instr_17_bF_buf31_), .Y(_4688_) );
NAND2X1 NAND2X1_207 ( .A(datapath_1_RegisterFile_regfile_mem_9__21_), .B(_3566__bF_buf0), .Y(_4689_) );
NAND3X1 NAND3X1_105 ( .A(datapath_1_Instr_16_bF_buf27_), .B(_4688_), .C(_4689_), .Y(_4690_) );
NAND2X1 NAND2X1_208 ( .A(datapath_1_RegisterFile_regfile_mem_10__21_), .B(datapath_1_Instr_17_bF_buf30_), .Y(_4691_) );
AOI21X1 AOI21X1_196 ( .A(_3566__bF_buf0), .B(datapath_1_RegisterFile_regfile_mem_8__21_), .C(datapath_1_Instr_16_bF_buf26_), .Y(_4692_) );
NAND2X1 NAND2X1_209 ( .A(_4691_), .B(_4692_), .Y(_4693_) );
NAND3X1 NAND3X1_106 ( .A(_3567__bF_buf8), .B(_4690_), .C(_4693_), .Y(_4694_) );
NAND2X1 NAND2X1_210 ( .A(datapath_1_RegisterFile_regfile_mem_15__21_), .B(datapath_1_Instr_17_bF_buf29_), .Y(_4695_) );
NAND2X1 NAND2X1_211 ( .A(datapath_1_RegisterFile_regfile_mem_13__21_), .B(_3566__bF_buf0), .Y(_4696_) );
NAND3X1 NAND3X1_107 ( .A(datapath_1_Instr_16_bF_buf25_), .B(_4695_), .C(_4696_), .Y(_4697_) );
NAND2X1 NAND2X1_212 ( .A(datapath_1_RegisterFile_regfile_mem_14__21_), .B(datapath_1_Instr_17_bF_buf28_), .Y(_4698_) );
AOI21X1 AOI21X1_197 ( .A(_3566__bF_buf0), .B(datapath_1_RegisterFile_regfile_mem_12__21_), .C(datapath_1_Instr_16_bF_buf24_), .Y(_4699_) );
NAND2X1 NAND2X1_213 ( .A(_4698_), .B(_4699_), .Y(_4700_) );
NAND3X1 NAND3X1_108 ( .A(datapath_1_Instr_18_bF_buf15_), .B(_4697_), .C(_4700_), .Y(_4701_) );
AOI21X1 AOI21X1_198 ( .A(_4694_), .B(_4701_), .C(_3571__bF_buf3), .Y(_4702_) );
OAI21X1 OAI21X1_185 ( .A(_4687_), .B(_4702_), .C(_3570__bF_buf3), .Y(_4703_) );
MUX2X1 MUX2X1_87 ( .A(datapath_1_RegisterFile_regfile_mem_17__21_), .B(datapath_1_RegisterFile_regfile_mem_16__21_), .S(datapath_1_Instr_16_bF_buf23_), .Y(_4704_) );
NOR2X1 NOR2X1_84 ( .A(datapath_1_RegisterFile_regfile_mem_19__21_), .B(_3588__bF_buf24), .Y(_4705_) );
OAI21X1 OAI21X1_186 ( .A(datapath_1_RegisterFile_regfile_mem_18__21_), .B(datapath_1_Instr_16_bF_buf22_), .C(datapath_1_Instr_17_bF_buf27_), .Y(_4706_) );
OAI22X1 OAI22X1_70 ( .A(_4706_), .B(_4705_), .C(datapath_1_Instr_17_bF_buf26_), .D(_4704_), .Y(_4707_) );
NAND2X1 NAND2X1_214 ( .A(_3567__bF_buf2), .B(_4707_), .Y(_4708_) );
MUX2X1 MUX2X1_88 ( .A(datapath_1_RegisterFile_regfile_mem_21__21_), .B(datapath_1_RegisterFile_regfile_mem_20__21_), .S(datapath_1_Instr_16_bF_buf21_), .Y(_4709_) );
NOR2X1 NOR2X1_85 ( .A(datapath_1_RegisterFile_regfile_mem_23__21_), .B(_3588__bF_buf24), .Y(_4710_) );
OAI21X1 OAI21X1_187 ( .A(datapath_1_RegisterFile_regfile_mem_22__21_), .B(datapath_1_Instr_16_bF_buf20_), .C(datapath_1_Instr_17_bF_buf25_), .Y(_4711_) );
OAI22X1 OAI22X1_71 ( .A(_4711_), .B(_4710_), .C(datapath_1_Instr_17_bF_buf24_), .D(_4709_), .Y(_4712_) );
NAND2X1 NAND2X1_215 ( .A(datapath_1_Instr_18_bF_buf14_), .B(_4712_), .Y(_4713_) );
AOI21X1 AOI21X1_199 ( .A(_4708_), .B(_4713_), .C(datapath_1_Instr_19_bF_buf4_), .Y(_4714_) );
INVX1 INVX1_61 ( .A(datapath_1_RegisterFile_regfile_mem_27__21_), .Y(_4715_) );
AOI21X1 AOI21X1_200 ( .A(datapath_1_RegisterFile_regfile_mem_31__21_), .B(datapath_1_Instr_18_bF_buf13_), .C(_3588__bF_buf24), .Y(_4716_) );
OAI21X1 OAI21X1_188 ( .A(_4715_), .B(datapath_1_Instr_18_bF_buf12_), .C(_4716_), .Y(_4717_) );
INVX1 INVX1_62 ( .A(datapath_1_RegisterFile_regfile_mem_26__21_), .Y(_4718_) );
AOI21X1 AOI21X1_201 ( .A(datapath_1_RegisterFile_regfile_mem_30__21_), .B(datapath_1_Instr_18_bF_buf11_), .C(datapath_1_Instr_16_bF_buf19_), .Y(_4719_) );
OAI21X1 OAI21X1_189 ( .A(_4718_), .B(datapath_1_Instr_18_bF_buf10_), .C(_4719_), .Y(_4720_) );
NAND3X1 NAND3X1_109 ( .A(datapath_1_Instr_17_bF_buf23_), .B(_4720_), .C(_4717_), .Y(_4721_) );
INVX1 INVX1_63 ( .A(datapath_1_RegisterFile_regfile_mem_25__21_), .Y(_4722_) );
AOI21X1 AOI21X1_202 ( .A(datapath_1_RegisterFile_regfile_mem_29__21_), .B(datapath_1_Instr_18_bF_buf9_), .C(_3588__bF_buf5), .Y(_4723_) );
OAI21X1 OAI21X1_190 ( .A(_4722_), .B(datapath_1_Instr_18_bF_buf8_), .C(_4723_), .Y(_4724_) );
INVX1 INVX1_64 ( .A(datapath_1_RegisterFile_regfile_mem_24__21_), .Y(_4725_) );
AOI21X1 AOI21X1_203 ( .A(datapath_1_RegisterFile_regfile_mem_28__21_), .B(datapath_1_Instr_18_bF_buf7_), .C(datapath_1_Instr_16_bF_buf18_), .Y(_4726_) );
OAI21X1 OAI21X1_191 ( .A(_4725_), .B(datapath_1_Instr_18_bF_buf6_), .C(_4726_), .Y(_4727_) );
NAND3X1 NAND3X1_110 ( .A(_3566__bF_buf10), .B(_4727_), .C(_4724_), .Y(_4728_) );
AOI21X1 AOI21X1_204 ( .A(_4721_), .B(_4728_), .C(_3571__bF_buf5), .Y(_4729_) );
OAI21X1 OAI21X1_192 ( .A(_4729_), .B(_4714_), .C(datapath_1_Instr_20_bF_buf4_), .Y(_4730_) );
AOI22X1 AOI22X1_35 ( .A(_3565__bF_buf4), .B(_3569__bF_buf4), .C(_4703_), .D(_4730_), .Y(datapath_1_RD2_21_) );
NAND2X1 NAND2X1_216 ( .A(datapath_1_RegisterFile_regfile_mem_27__22_), .B(datapath_1_Instr_16_bF_buf17_), .Y(_4731_) );
NAND2X1 NAND2X1_217 ( .A(datapath_1_RegisterFile_regfile_mem_26__22_), .B(_3588__bF_buf27), .Y(_4732_) );
NAND3X1 NAND3X1_111 ( .A(datapath_1_Instr_17_bF_buf22_), .B(_4731_), .C(_4732_), .Y(_4733_) );
NAND2X1 NAND2X1_218 ( .A(datapath_1_RegisterFile_regfile_mem_25__22_), .B(datapath_1_Instr_16_bF_buf16_), .Y(_4734_) );
AOI21X1 AOI21X1_205 ( .A(_3588__bF_buf27), .B(datapath_1_RegisterFile_regfile_mem_24__22_), .C(datapath_1_Instr_17_bF_buf21_), .Y(_4735_) );
NAND2X1 NAND2X1_219 ( .A(_4734_), .B(_4735_), .Y(_4736_) );
NAND3X1 NAND3X1_112 ( .A(_3567__bF_buf9), .B(_4733_), .C(_4736_), .Y(_4737_) );
NAND2X1 NAND2X1_220 ( .A(datapath_1_RegisterFile_regfile_mem_31__22_), .B(datapath_1_Instr_16_bF_buf15_), .Y(_4738_) );
AOI21X1 AOI21X1_206 ( .A(_3588__bF_buf29), .B(datapath_1_RegisterFile_regfile_mem_30__22_), .C(_3566__bF_buf4), .Y(_4739_) );
NAND2X1 NAND2X1_221 ( .A(_4738_), .B(_4739_), .Y(_4740_) );
INVX1 INVX1_65 ( .A(datapath_1_RegisterFile_regfile_mem_28__22_), .Y(_4741_) );
AOI21X1 AOI21X1_207 ( .A(datapath_1_RegisterFile_regfile_mem_29__22_), .B(datapath_1_Instr_16_bF_buf14_), .C(datapath_1_Instr_17_bF_buf20_), .Y(_4742_) );
OAI21X1 OAI21X1_193 ( .A(_4741_), .B(datapath_1_Instr_16_bF_buf13_), .C(_4742_), .Y(_4743_) );
NAND3X1 NAND3X1_113 ( .A(datapath_1_Instr_18_bF_buf5_), .B(_4743_), .C(_4740_), .Y(_4744_) );
AOI21X1 AOI21X1_208 ( .A(_4737_), .B(_4744_), .C(_3571__bF_buf5), .Y(_4745_) );
MUX2X1 MUX2X1_89 ( .A(datapath_1_RegisterFile_regfile_mem_17__22_), .B(datapath_1_RegisterFile_regfile_mem_16__22_), .S(datapath_1_Instr_16_bF_buf12_), .Y(_4746_) );
NOR2X1 NOR2X1_86 ( .A(datapath_1_RegisterFile_regfile_mem_19__22_), .B(_3588__bF_buf41), .Y(_4747_) );
OAI21X1 OAI21X1_194 ( .A(datapath_1_RegisterFile_regfile_mem_18__22_), .B(datapath_1_Instr_16_bF_buf11_), .C(datapath_1_Instr_17_bF_buf19_), .Y(_4748_) );
OAI22X1 OAI22X1_72 ( .A(_4748_), .B(_4747_), .C(datapath_1_Instr_17_bF_buf18_), .D(_4746_), .Y(_4749_) );
NAND2X1 NAND2X1_222 ( .A(_3567__bF_buf3), .B(_4749_), .Y(_4750_) );
MUX2X1 MUX2X1_90 ( .A(datapath_1_RegisterFile_regfile_mem_21__22_), .B(datapath_1_RegisterFile_regfile_mem_20__22_), .S(datapath_1_Instr_16_bF_buf10_), .Y(_4751_) );
NOR2X1 NOR2X1_87 ( .A(datapath_1_RegisterFile_regfile_mem_23__22_), .B(_3588__bF_buf41), .Y(_4752_) );
OAI21X1 OAI21X1_195 ( .A(datapath_1_RegisterFile_regfile_mem_22__22_), .B(datapath_1_Instr_16_bF_buf9_), .C(datapath_1_Instr_17_bF_buf17_), .Y(_4753_) );
OAI22X1 OAI22X1_73 ( .A(_4753_), .B(_4752_), .C(datapath_1_Instr_17_bF_buf16_), .D(_4751_), .Y(_4754_) );
NAND2X1 NAND2X1_223 ( .A(datapath_1_Instr_18_bF_buf4_), .B(_4754_), .Y(_4755_) );
AOI21X1 AOI21X1_209 ( .A(_4750_), .B(_4755_), .C(datapath_1_Instr_19_bF_buf3_), .Y(_4756_) );
OAI21X1 OAI21X1_196 ( .A(_4745_), .B(_4756_), .C(datapath_1_Instr_20_bF_buf3_), .Y(_4757_) );
NAND2X1 NAND2X1_224 ( .A(datapath_1_RegisterFile_regfile_mem_11__22_), .B(datapath_1_Instr_17_bF_buf15_), .Y(_4758_) );
NAND2X1 NAND2X1_225 ( .A(datapath_1_RegisterFile_regfile_mem_9__22_), .B(_3566__bF_buf3), .Y(_4759_) );
NAND3X1 NAND3X1_114 ( .A(datapath_1_Instr_16_bF_buf8_), .B(_4758_), .C(_4759_), .Y(_4760_) );
NAND2X1 NAND2X1_226 ( .A(datapath_1_RegisterFile_regfile_mem_10__22_), .B(datapath_1_Instr_17_bF_buf14_), .Y(_4761_) );
AOI21X1 AOI21X1_210 ( .A(_3566__bF_buf3), .B(datapath_1_RegisterFile_regfile_mem_8__22_), .C(datapath_1_Instr_16_bF_buf7_), .Y(_4762_) );
NAND2X1 NAND2X1_227 ( .A(_4761_), .B(_4762_), .Y(_4763_) );
NAND3X1 NAND3X1_115 ( .A(_3567__bF_buf1), .B(_4760_), .C(_4763_), .Y(_4764_) );
NAND2X1 NAND2X1_228 ( .A(datapath_1_RegisterFile_regfile_mem_15__22_), .B(datapath_1_Instr_17_bF_buf13_), .Y(_4765_) );
NAND2X1 NAND2X1_229 ( .A(datapath_1_RegisterFile_regfile_mem_13__22_), .B(_3566__bF_buf3), .Y(_4766_) );
NAND3X1 NAND3X1_116 ( .A(datapath_1_Instr_16_bF_buf6_), .B(_4765_), .C(_4766_), .Y(_4767_) );
NAND2X1 NAND2X1_230 ( .A(datapath_1_RegisterFile_regfile_mem_14__22_), .B(datapath_1_Instr_17_bF_buf12_), .Y(_4768_) );
AOI21X1 AOI21X1_211 ( .A(_3566__bF_buf3), .B(datapath_1_RegisterFile_regfile_mem_12__22_), .C(datapath_1_Instr_16_bF_buf5_), .Y(_4769_) );
NAND2X1 NAND2X1_231 ( .A(_4768_), .B(_4769_), .Y(_4770_) );
NAND3X1 NAND3X1_117 ( .A(datapath_1_Instr_18_bF_buf3_), .B(_4767_), .C(_4770_), .Y(_4771_) );
AOI21X1 AOI21X1_212 ( .A(_4764_), .B(_4771_), .C(_3571__bF_buf6), .Y(_4772_) );
INVX1 INVX1_66 ( .A(datapath_1_RegisterFile_regfile_mem_1__22_), .Y(_4773_) );
AOI21X1 AOI21X1_213 ( .A(datapath_1_RegisterFile_regfile_mem_5__22_), .B(datapath_1_Instr_18_bF_buf2_), .C(_3588__bF_buf20), .Y(_4774_) );
OAI21X1 OAI21X1_197 ( .A(_4773_), .B(datapath_1_Instr_18_bF_buf1_), .C(_4774_), .Y(_4775_) );
INVX1 INVX1_67 ( .A(datapath_1_RegisterFile_regfile_mem_0__22_), .Y(_4776_) );
AOI21X1 AOI21X1_214 ( .A(datapath_1_RegisterFile_regfile_mem_4__22_), .B(datapath_1_Instr_18_bF_buf0_), .C(datapath_1_Instr_16_bF_buf4_), .Y(_4777_) );
OAI21X1 OAI21X1_198 ( .A(_4776_), .B(datapath_1_Instr_18_bF_buf44_), .C(_4777_), .Y(_4778_) );
NAND3X1 NAND3X1_118 ( .A(_3566__bF_buf6), .B(_4778_), .C(_4775_), .Y(_4779_) );
INVX1 INVX1_68 ( .A(datapath_1_RegisterFile_regfile_mem_3__22_), .Y(_4780_) );
AOI21X1 AOI21X1_215 ( .A(datapath_1_RegisterFile_regfile_mem_7__22_), .B(datapath_1_Instr_18_bF_buf43_), .C(_3588__bF_buf20), .Y(_4781_) );
OAI21X1 OAI21X1_199 ( .A(_4780_), .B(datapath_1_Instr_18_bF_buf42_), .C(_4781_), .Y(_4782_) );
INVX1 INVX1_69 ( .A(datapath_1_RegisterFile_regfile_mem_2__22_), .Y(_4783_) );
AOI21X1 AOI21X1_216 ( .A(datapath_1_RegisterFile_regfile_mem_6__22_), .B(datapath_1_Instr_18_bF_buf41_), .C(datapath_1_Instr_16_bF_buf3_), .Y(_4784_) );
OAI21X1 OAI21X1_200 ( .A(_4783_), .B(datapath_1_Instr_18_bF_buf40_), .C(_4784_), .Y(_4785_) );
NAND3X1 NAND3X1_119 ( .A(datapath_1_Instr_17_bF_buf11_), .B(_4785_), .C(_4782_), .Y(_4786_) );
AOI21X1 AOI21X1_217 ( .A(_4779_), .B(_4786_), .C(datapath_1_Instr_19_bF_buf2_), .Y(_4787_) );
OAI21X1 OAI21X1_201 ( .A(_4787_), .B(_4772_), .C(_3570__bF_buf4), .Y(_4788_) );
AOI22X1 AOI22X1_36 ( .A(_3565__bF_buf2), .B(_3569__bF_buf2), .C(_4788_), .D(_4757_), .Y(datapath_1_RD2_22_) );
MUX2X1 MUX2X1_91 ( .A(datapath_1_RegisterFile_regfile_mem_9__23_), .B(datapath_1_RegisterFile_regfile_mem_8__23_), .S(datapath_1_Instr_16_bF_buf2_), .Y(_4789_) );
NOR2X1 NOR2X1_88 ( .A(datapath_1_RegisterFile_regfile_mem_11__23_), .B(_3588__bF_buf3), .Y(_4790_) );
OAI21X1 OAI21X1_202 ( .A(datapath_1_RegisterFile_regfile_mem_10__23_), .B(datapath_1_Instr_16_bF_buf1_), .C(datapath_1_Instr_17_bF_buf10_), .Y(_4791_) );
OAI22X1 OAI22X1_74 ( .A(_4791_), .B(_4790_), .C(datapath_1_Instr_17_bF_buf9_), .D(_4789_), .Y(_4792_) );
INVX1 INVX1_70 ( .A(datapath_1_RegisterFile_regfile_mem_15__23_), .Y(_4793_) );
AOI21X1 AOI21X1_218 ( .A(_3588__bF_buf35), .B(datapath_1_RegisterFile_regfile_mem_14__23_), .C(_3566__bF_buf3), .Y(_4794_) );
OAI21X1 OAI21X1_203 ( .A(_4793_), .B(_3588__bF_buf35), .C(_4794_), .Y(_4795_) );
NAND2X1 NAND2X1_232 ( .A(datapath_1_RegisterFile_regfile_mem_12__23_), .B(_3588__bF_buf35), .Y(_4796_) );
AOI21X1 AOI21X1_219 ( .A(datapath_1_RegisterFile_regfile_mem_13__23_), .B(datapath_1_Instr_16_bF_buf0_), .C(datapath_1_Instr_17_bF_buf8_), .Y(_4797_) );
AOI21X1 AOI21X1_220 ( .A(_4796_), .B(_4797_), .C(_3567__bF_buf6), .Y(_4798_) );
AOI22X1 AOI22X1_37 ( .A(_4795_), .B(_4798_), .C(_3567__bF_buf6), .D(_4792_), .Y(_4799_) );
NOR2X1 NOR2X1_89 ( .A(datapath_1_RegisterFile_regfile_mem_0__23_), .B(datapath_1_Instr_16_bF_buf55_), .Y(_4800_) );
OAI21X1 OAI21X1_204 ( .A(datapath_1_RegisterFile_regfile_mem_1__23_), .B(_3588__bF_buf35), .C(_3566__bF_buf3), .Y(_4801_) );
NOR2X1 NOR2X1_90 ( .A(datapath_1_RegisterFile_regfile_mem_3__23_), .B(_3588__bF_buf35), .Y(_4802_) );
OAI21X1 OAI21X1_205 ( .A(datapath_1_RegisterFile_regfile_mem_2__23_), .B(datapath_1_Instr_16_bF_buf54_), .C(datapath_1_Instr_17_bF_buf7_), .Y(_4803_) );
OAI22X1 OAI22X1_75 ( .A(_4802_), .B(_4803_), .C(_4800_), .D(_4801_), .Y(_4804_) );
NOR2X1 NOR2X1_91 ( .A(datapath_1_Instr_18_bF_buf39_), .B(_4804_), .Y(_4805_) );
MUX2X1 MUX2X1_92 ( .A(datapath_1_RegisterFile_regfile_mem_5__23_), .B(datapath_1_RegisterFile_regfile_mem_4__23_), .S(datapath_1_Instr_16_bF_buf53_), .Y(_4806_) );
NOR2X1 NOR2X1_92 ( .A(datapath_1_RegisterFile_regfile_mem_7__23_), .B(_3588__bF_buf3), .Y(_4807_) );
OAI21X1 OAI21X1_206 ( .A(datapath_1_RegisterFile_regfile_mem_6__23_), .B(datapath_1_Instr_16_bF_buf52_), .C(datapath_1_Instr_17_bF_buf6_), .Y(_4808_) );
OAI22X1 OAI22X1_76 ( .A(_4808_), .B(_4807_), .C(datapath_1_Instr_17_bF_buf5_), .D(_4806_), .Y(_4809_) );
OAI21X1 OAI21X1_207 ( .A(_3567__bF_buf6), .B(_4809_), .C(_3571__bF_buf6), .Y(_4810_) );
OAI22X1 OAI22X1_77 ( .A(_3571__bF_buf6), .B(_4799_), .C(_4805_), .D(_4810_), .Y(_4811_) );
NAND2X1 NAND2X1_233 ( .A(_3570__bF_buf3), .B(_4811_), .Y(_4812_) );
AOI21X1 AOI21X1_221 ( .A(datapath_1_RegisterFile_regfile_mem_23__23_), .B(datapath_1_Instr_18_bF_buf38_), .C(_3588__bF_buf33), .Y(_4813_) );
OAI21X1 OAI21X1_208 ( .A(_3131_), .B(datapath_1_Instr_18_bF_buf37_), .C(_4813_), .Y(_4814_) );
NAND2X1 NAND2X1_234 ( .A(datapath_1_RegisterFile_regfile_mem_18__23_), .B(_3567__bF_buf2), .Y(_4815_) );
AOI21X1 AOI21X1_222 ( .A(datapath_1_RegisterFile_regfile_mem_22__23_), .B(datapath_1_Instr_18_bF_buf36_), .C(datapath_1_Instr_16_bF_buf51_), .Y(_4816_) );
AOI21X1 AOI21X1_223 ( .A(_4815_), .B(_4816_), .C(_3566__bF_buf10), .Y(_4817_) );
AOI21X1 AOI21X1_224 ( .A(datapath_1_RegisterFile_regfile_mem_21__23_), .B(datapath_1_Instr_18_bF_buf35_), .C(_3588__bF_buf33), .Y(_4818_) );
OAI21X1 OAI21X1_209 ( .A(_3137_), .B(datapath_1_Instr_18_bF_buf34_), .C(_4818_), .Y(_4819_) );
NAND2X1 NAND2X1_235 ( .A(datapath_1_RegisterFile_regfile_mem_16__23_), .B(_3567__bF_buf2), .Y(_4820_) );
AOI21X1 AOI21X1_225 ( .A(datapath_1_RegisterFile_regfile_mem_20__23_), .B(datapath_1_Instr_18_bF_buf33_), .C(datapath_1_Instr_16_bF_buf50_), .Y(_4821_) );
AOI21X1 AOI21X1_226 ( .A(_4820_), .B(_4821_), .C(datapath_1_Instr_17_bF_buf4_), .Y(_4822_) );
AOI22X1 AOI22X1_38 ( .A(_4817_), .B(_4814_), .C(_4819_), .D(_4822_), .Y(_4823_) );
NOR2X1 NOR2X1_93 ( .A(datapath_1_RegisterFile_regfile_mem_24__23_), .B(datapath_1_Instr_16_bF_buf49_), .Y(_4824_) );
OAI21X1 OAI21X1_210 ( .A(datapath_1_RegisterFile_regfile_mem_25__23_), .B(_3588__bF_buf5), .C(_3566__bF_buf10), .Y(_4825_) );
NOR2X1 NOR2X1_94 ( .A(datapath_1_RegisterFile_regfile_mem_27__23_), .B(_3588__bF_buf5), .Y(_4826_) );
OAI21X1 OAI21X1_211 ( .A(datapath_1_RegisterFile_regfile_mem_26__23_), .B(datapath_1_Instr_16_bF_buf48_), .C(datapath_1_Instr_17_bF_buf3_), .Y(_4827_) );
OAI22X1 OAI22X1_78 ( .A(_4826_), .B(_4827_), .C(_4824_), .D(_4825_), .Y(_4828_) );
NOR2X1 NOR2X1_95 ( .A(datapath_1_Instr_18_bF_buf32_), .B(_4828_), .Y(_4829_) );
MUX2X1 MUX2X1_93 ( .A(datapath_1_RegisterFile_regfile_mem_29__23_), .B(datapath_1_RegisterFile_regfile_mem_28__23_), .S(datapath_1_Instr_16_bF_buf47_), .Y(_4830_) );
NOR2X1 NOR2X1_96 ( .A(datapath_1_RegisterFile_regfile_mem_31__23_), .B(_3588__bF_buf33), .Y(_4831_) );
OAI21X1 OAI21X1_212 ( .A(datapath_1_RegisterFile_regfile_mem_30__23_), .B(datapath_1_Instr_16_bF_buf46_), .C(datapath_1_Instr_17_bF_buf2_), .Y(_4832_) );
OAI22X1 OAI22X1_79 ( .A(_4832_), .B(_4831_), .C(datapath_1_Instr_17_bF_buf1_), .D(_4830_), .Y(_4833_) );
OAI21X1 OAI21X1_213 ( .A(_3567__bF_buf2), .B(_4833_), .C(datapath_1_Instr_19_bF_buf1_), .Y(_4834_) );
OAI22X1 OAI22X1_80 ( .A(datapath_1_Instr_19_bF_buf0_), .B(_4823_), .C(_4829_), .D(_4834_), .Y(_4835_) );
NAND2X1 NAND2X1_236 ( .A(datapath_1_Instr_20_bF_buf2_), .B(_4835_), .Y(_4836_) );
AOI22X1 AOI22X1_39 ( .A(_3565__bF_buf4), .B(_3569__bF_buf4), .C(_4836_), .D(_4812_), .Y(datapath_1_RD2_23_) );
NAND2X1 NAND2X1_237 ( .A(datapath_1_RegisterFile_regfile_mem_11__24_), .B(datapath_1_Instr_17_bF_buf0_), .Y(_4837_) );
NAND2X1 NAND2X1_238 ( .A(datapath_1_RegisterFile_regfile_mem_9__24_), .B(_3566__bF_buf2), .Y(_4838_) );
NAND3X1 NAND3X1_120 ( .A(datapath_1_Instr_16_bF_buf45_), .B(_4837_), .C(_4838_), .Y(_4839_) );
NAND2X1 NAND2X1_239 ( .A(datapath_1_RegisterFile_regfile_mem_10__24_), .B(datapath_1_Instr_17_bF_buf50_), .Y(_4840_) );
AOI21X1 AOI21X1_227 ( .A(_3566__bF_buf2), .B(datapath_1_RegisterFile_regfile_mem_8__24_), .C(datapath_1_Instr_16_bF_buf44_), .Y(_4841_) );
NAND2X1 NAND2X1_240 ( .A(_4840_), .B(_4841_), .Y(_4842_) );
NAND3X1 NAND3X1_121 ( .A(_3567__bF_buf7), .B(_4839_), .C(_4842_), .Y(_4843_) );
NAND2X1 NAND2X1_241 ( .A(datapath_1_RegisterFile_regfile_mem_15__24_), .B(datapath_1_Instr_17_bF_buf49_), .Y(_4844_) );
NAND2X1 NAND2X1_242 ( .A(datapath_1_RegisterFile_regfile_mem_13__24_), .B(_3566__bF_buf2), .Y(_4845_) );
NAND3X1 NAND3X1_122 ( .A(datapath_1_Instr_16_bF_buf43_), .B(_4844_), .C(_4845_), .Y(_4846_) );
NAND2X1 NAND2X1_243 ( .A(datapath_1_RegisterFile_regfile_mem_14__24_), .B(datapath_1_Instr_17_bF_buf48_), .Y(_4847_) );
AOI21X1 AOI21X1_228 ( .A(_3566__bF_buf2), .B(datapath_1_RegisterFile_regfile_mem_12__24_), .C(datapath_1_Instr_16_bF_buf42_), .Y(_4848_) );
NAND2X1 NAND2X1_244 ( .A(_4847_), .B(_4848_), .Y(_4849_) );
NAND3X1 NAND3X1_123 ( .A(datapath_1_Instr_18_bF_buf31_), .B(_4846_), .C(_4849_), .Y(_4850_) );
AOI21X1 AOI21X1_229 ( .A(_4843_), .B(_4850_), .C(_3571__bF_buf0), .Y(_4851_) );
INVX1 INVX1_71 ( .A(datapath_1_RegisterFile_regfile_mem_1__24_), .Y(_4852_) );
AOI21X1 AOI21X1_230 ( .A(datapath_1_RegisterFile_regfile_mem_5__24_), .B(datapath_1_Instr_18_bF_buf30_), .C(_3588__bF_buf17), .Y(_4853_) );
OAI21X1 OAI21X1_214 ( .A(_4852_), .B(datapath_1_Instr_18_bF_buf29_), .C(_4853_), .Y(_4854_) );
INVX1 INVX1_72 ( .A(datapath_1_RegisterFile_regfile_mem_0__24_), .Y(_4855_) );
AOI21X1 AOI21X1_231 ( .A(datapath_1_RegisterFile_regfile_mem_4__24_), .B(datapath_1_Instr_18_bF_buf28_), .C(datapath_1_Instr_16_bF_buf41_), .Y(_4856_) );
OAI21X1 OAI21X1_215 ( .A(_4855_), .B(datapath_1_Instr_18_bF_buf27_), .C(_4856_), .Y(_4857_) );
NAND3X1 NAND3X1_124 ( .A(_3566__bF_buf2), .B(_4857_), .C(_4854_), .Y(_4858_) );
INVX1 INVX1_73 ( .A(datapath_1_RegisterFile_regfile_mem_3__24_), .Y(_4859_) );
AOI21X1 AOI21X1_232 ( .A(datapath_1_RegisterFile_regfile_mem_7__24_), .B(datapath_1_Instr_18_bF_buf26_), .C(_3588__bF_buf28), .Y(_4860_) );
OAI21X1 OAI21X1_216 ( .A(_4859_), .B(datapath_1_Instr_18_bF_buf25_), .C(_4860_), .Y(_4861_) );
INVX1 INVX1_74 ( .A(datapath_1_RegisterFile_regfile_mem_2__24_), .Y(_4862_) );
AOI21X1 AOI21X1_233 ( .A(datapath_1_RegisterFile_regfile_mem_6__24_), .B(datapath_1_Instr_18_bF_buf24_), .C(datapath_1_Instr_16_bF_buf40_), .Y(_4863_) );
OAI21X1 OAI21X1_217 ( .A(_4862_), .B(datapath_1_Instr_18_bF_buf23_), .C(_4863_), .Y(_4864_) );
NAND3X1 NAND3X1_125 ( .A(datapath_1_Instr_17_bF_buf47_), .B(_4864_), .C(_4861_), .Y(_4865_) );
AOI21X1 AOI21X1_234 ( .A(_4858_), .B(_4865_), .C(datapath_1_Instr_19_bF_buf6_), .Y(_4866_) );
OAI21X1 OAI21X1_218 ( .A(_4866_), .B(_4851_), .C(_3570__bF_buf1), .Y(_4867_) );
INVX1 INVX1_75 ( .A(datapath_1_RegisterFile_regfile_mem_19__24_), .Y(_4868_) );
AOI21X1 AOI21X1_235 ( .A(datapath_1_RegisterFile_regfile_mem_23__24_), .B(datapath_1_Instr_18_bF_buf22_), .C(_3588__bF_buf15), .Y(_4869_) );
OAI21X1 OAI21X1_219 ( .A(_4868_), .B(datapath_1_Instr_18_bF_buf21_), .C(_4869_), .Y(_4870_) );
NAND2X1 NAND2X1_245 ( .A(datapath_1_RegisterFile_regfile_mem_18__24_), .B(_3567__bF_buf0), .Y(_4871_) );
AOI21X1 AOI21X1_236 ( .A(datapath_1_RegisterFile_regfile_mem_22__24_), .B(datapath_1_Instr_18_bF_buf20_), .C(datapath_1_Instr_16_bF_buf39_), .Y(_4872_) );
AOI21X1 AOI21X1_237 ( .A(_4871_), .B(_4872_), .C(_3566__bF_buf9), .Y(_4873_) );
INVX1 INVX1_76 ( .A(datapath_1_RegisterFile_regfile_mem_17__24_), .Y(_4874_) );
AOI21X1 AOI21X1_238 ( .A(datapath_1_RegisterFile_regfile_mem_21__24_), .B(datapath_1_Instr_18_bF_buf19_), .C(_3588__bF_buf15), .Y(_4875_) );
OAI21X1 OAI21X1_220 ( .A(_4874_), .B(datapath_1_Instr_18_bF_buf18_), .C(_4875_), .Y(_4876_) );
NAND2X1 NAND2X1_246 ( .A(datapath_1_RegisterFile_regfile_mem_16__24_), .B(_3567__bF_buf0), .Y(_4877_) );
AOI21X1 AOI21X1_239 ( .A(datapath_1_RegisterFile_regfile_mem_20__24_), .B(datapath_1_Instr_18_bF_buf17_), .C(datapath_1_Instr_16_bF_buf38_), .Y(_4878_) );
AOI21X1 AOI21X1_240 ( .A(_4877_), .B(_4878_), .C(datapath_1_Instr_17_bF_buf46_), .Y(_4879_) );
AOI22X1 AOI22X1_40 ( .A(_4873_), .B(_4870_), .C(_4876_), .D(_4879_), .Y(_4880_) );
NOR2X1 NOR2X1_97 ( .A(datapath_1_RegisterFile_regfile_mem_24__24_), .B(datapath_1_Instr_16_bF_buf37_), .Y(_4881_) );
OAI21X1 OAI21X1_221 ( .A(datapath_1_RegisterFile_regfile_mem_25__24_), .B(_3588__bF_buf19), .C(_3566__bF_buf9), .Y(_4882_) );
NOR2X1 NOR2X1_98 ( .A(datapath_1_RegisterFile_regfile_mem_27__24_), .B(_3588__bF_buf19), .Y(_4883_) );
OAI21X1 OAI21X1_222 ( .A(datapath_1_RegisterFile_regfile_mem_26__24_), .B(datapath_1_Instr_16_bF_buf36_), .C(datapath_1_Instr_17_bF_buf45_), .Y(_4884_) );
OAI22X1 OAI22X1_81 ( .A(_4883_), .B(_4884_), .C(_4881_), .D(_4882_), .Y(_4885_) );
NOR2X1 NOR2X1_99 ( .A(datapath_1_Instr_18_bF_buf16_), .B(_4885_), .Y(_4886_) );
MUX2X1 MUX2X1_94 ( .A(datapath_1_RegisterFile_regfile_mem_29__24_), .B(datapath_1_RegisterFile_regfile_mem_28__24_), .S(datapath_1_Instr_16_bF_buf35_), .Y(_4887_) );
NOR2X1 NOR2X1_100 ( .A(datapath_1_RegisterFile_regfile_mem_31__24_), .B(_3588__bF_buf26), .Y(_4888_) );
OAI21X1 OAI21X1_223 ( .A(datapath_1_RegisterFile_regfile_mem_30__24_), .B(datapath_1_Instr_16_bF_buf34_), .C(datapath_1_Instr_17_bF_buf44_), .Y(_4889_) );
OAI22X1 OAI22X1_82 ( .A(_4889_), .B(_4888_), .C(datapath_1_Instr_17_bF_buf43_), .D(_4887_), .Y(_4890_) );
OAI21X1 OAI21X1_224 ( .A(_3567__bF_buf0), .B(_4890_), .C(datapath_1_Instr_19_bF_buf5_), .Y(_4891_) );
OAI22X1 OAI22X1_83 ( .A(datapath_1_Instr_19_bF_buf4_), .B(_4880_), .C(_4886_), .D(_4891_), .Y(_4892_) );
NAND2X1 NAND2X1_247 ( .A(datapath_1_Instr_20_bF_buf1_), .B(_4892_), .Y(_4893_) );
AOI22X1 AOI22X1_41 ( .A(_3565__bF_buf0), .B(_3569__bF_buf0), .C(_4867_), .D(_4893_), .Y(datapath_1_RD2_24_) );
NAND2X1 NAND2X1_248 ( .A(datapath_1_RegisterFile_regfile_mem_27__25_), .B(datapath_1_Instr_16_bF_buf33_), .Y(_4894_) );
NAND2X1 NAND2X1_249 ( .A(datapath_1_RegisterFile_regfile_mem_26__25_), .B(_3588__bF_buf39), .Y(_4895_) );
NAND3X1 NAND3X1_126 ( .A(datapath_1_Instr_17_bF_buf42_), .B(_4894_), .C(_4895_), .Y(_4896_) );
NAND2X1 NAND2X1_250 ( .A(datapath_1_RegisterFile_regfile_mem_25__25_), .B(datapath_1_Instr_16_bF_buf32_), .Y(_4897_) );
AOI21X1 AOI21X1_241 ( .A(_3588__bF_buf2), .B(datapath_1_RegisterFile_regfile_mem_24__25_), .C(datapath_1_Instr_17_bF_buf41_), .Y(_4898_) );
NAND2X1 NAND2X1_251 ( .A(_4897_), .B(_4898_), .Y(_4899_) );
NAND3X1 NAND3X1_127 ( .A(_3567__bF_buf2), .B(_4896_), .C(_4899_), .Y(_4900_) );
NAND2X1 NAND2X1_252 ( .A(datapath_1_RegisterFile_regfile_mem_31__25_), .B(datapath_1_Instr_16_bF_buf31_), .Y(_4901_) );
AOI21X1 AOI21X1_242 ( .A(_3588__bF_buf39), .B(datapath_1_RegisterFile_regfile_mem_30__25_), .C(_3566__bF_buf10), .Y(_4902_) );
NAND2X1 NAND2X1_253 ( .A(_4901_), .B(_4902_), .Y(_4903_) );
INVX1 INVX1_77 ( .A(datapath_1_RegisterFile_regfile_mem_28__25_), .Y(_4904_) );
AOI21X1 AOI21X1_243 ( .A(datapath_1_RegisterFile_regfile_mem_29__25_), .B(datapath_1_Instr_16_bF_buf30_), .C(datapath_1_Instr_17_bF_buf40_), .Y(_4905_) );
OAI21X1 OAI21X1_225 ( .A(_4904_), .B(datapath_1_Instr_16_bF_buf29_), .C(_4905_), .Y(_4906_) );
NAND3X1 NAND3X1_128 ( .A(datapath_1_Instr_18_bF_buf15_), .B(_4906_), .C(_4903_), .Y(_4907_) );
AOI21X1 AOI21X1_244 ( .A(_4900_), .B(_4907_), .C(_3571__bF_buf7), .Y(_4908_) );
MUX2X1 MUX2X1_95 ( .A(datapath_1_RegisterFile_regfile_mem_17__25_), .B(datapath_1_RegisterFile_regfile_mem_16__25_), .S(datapath_1_Instr_16_bF_buf28_), .Y(_4909_) );
NOR2X1 NOR2X1_101 ( .A(datapath_1_RegisterFile_regfile_mem_19__25_), .B(_3588__bF_buf15), .Y(_4910_) );
OAI21X1 OAI21X1_226 ( .A(datapath_1_RegisterFile_regfile_mem_18__25_), .B(datapath_1_Instr_16_bF_buf27_), .C(datapath_1_Instr_17_bF_buf39_), .Y(_4911_) );
OAI22X1 OAI22X1_84 ( .A(_4911_), .B(_4910_), .C(datapath_1_Instr_17_bF_buf38_), .D(_4909_), .Y(_4912_) );
NAND2X1 NAND2X1_254 ( .A(_3567__bF_buf0), .B(_4912_), .Y(_4913_) );
MUX2X1 MUX2X1_96 ( .A(datapath_1_RegisterFile_regfile_mem_21__25_), .B(datapath_1_RegisterFile_regfile_mem_20__25_), .S(datapath_1_Instr_16_bF_buf26_), .Y(_4914_) );
NOR2X1 NOR2X1_102 ( .A(datapath_1_RegisterFile_regfile_mem_23__25_), .B(_3588__bF_buf31), .Y(_4915_) );
OAI21X1 OAI21X1_227 ( .A(datapath_1_RegisterFile_regfile_mem_22__25_), .B(datapath_1_Instr_16_bF_buf25_), .C(datapath_1_Instr_17_bF_buf37_), .Y(_4916_) );
OAI22X1 OAI22X1_85 ( .A(_4916_), .B(_4915_), .C(datapath_1_Instr_17_bF_buf36_), .D(_4914_), .Y(_4917_) );
NAND2X1 NAND2X1_255 ( .A(datapath_1_Instr_18_bF_buf14_), .B(_4917_), .Y(_4918_) );
AOI21X1 AOI21X1_245 ( .A(_4913_), .B(_4918_), .C(datapath_1_Instr_19_bF_buf3_), .Y(_4919_) );
OAI21X1 OAI21X1_228 ( .A(_4908_), .B(_4919_), .C(datapath_1_Instr_20_bF_buf0_), .Y(_4920_) );
NAND2X1 NAND2X1_256 ( .A(datapath_1_RegisterFile_regfile_mem_11__25_), .B(datapath_1_Instr_17_bF_buf35_), .Y(_4921_) );
NAND2X1 NAND2X1_257 ( .A(datapath_1_RegisterFile_regfile_mem_9__25_), .B(_3566__bF_buf1), .Y(_4922_) );
NAND3X1 NAND3X1_129 ( .A(datapath_1_Instr_16_bF_buf24_), .B(_4921_), .C(_4922_), .Y(_4923_) );
NAND2X1 NAND2X1_258 ( .A(datapath_1_RegisterFile_regfile_mem_10__25_), .B(datapath_1_Instr_17_bF_buf34_), .Y(_4924_) );
AOI21X1 AOI21X1_246 ( .A(_3566__bF_buf1), .B(datapath_1_RegisterFile_regfile_mem_8__25_), .C(datapath_1_Instr_16_bF_buf23_), .Y(_4925_) );
NAND2X1 NAND2X1_259 ( .A(_4924_), .B(_4925_), .Y(_4926_) );
NAND3X1 NAND3X1_130 ( .A(_3567__bF_buf4), .B(_4923_), .C(_4926_), .Y(_4927_) );
NAND2X1 NAND2X1_260 ( .A(datapath_1_RegisterFile_regfile_mem_15__25_), .B(datapath_1_Instr_17_bF_buf33_), .Y(_4928_) );
NAND2X1 NAND2X1_261 ( .A(datapath_1_RegisterFile_regfile_mem_13__25_), .B(_3566__bF_buf7), .Y(_4929_) );
NAND3X1 NAND3X1_131 ( .A(datapath_1_Instr_16_bF_buf22_), .B(_4928_), .C(_4929_), .Y(_4930_) );
NAND2X1 NAND2X1_262 ( .A(datapath_1_RegisterFile_regfile_mem_14__25_), .B(datapath_1_Instr_17_bF_buf32_), .Y(_4931_) );
AOI21X1 AOI21X1_247 ( .A(_3566__bF_buf1), .B(datapath_1_RegisterFile_regfile_mem_12__25_), .C(datapath_1_Instr_16_bF_buf21_), .Y(_4932_) );
NAND2X1 NAND2X1_263 ( .A(_4931_), .B(_4932_), .Y(_4933_) );
NAND3X1 NAND3X1_132 ( .A(datapath_1_Instr_18_bF_buf13_), .B(_4930_), .C(_4933_), .Y(_4934_) );
AOI21X1 AOI21X1_248 ( .A(_4927_), .B(_4934_), .C(_3571__bF_buf1), .Y(_4935_) );
INVX1 INVX1_78 ( .A(datapath_1_RegisterFile_regfile_mem_1__25_), .Y(_4936_) );
AOI21X1 AOI21X1_249 ( .A(datapath_1_RegisterFile_regfile_mem_5__25_), .B(datapath_1_Instr_18_bF_buf12_), .C(_3588__bF_buf6), .Y(_4937_) );
OAI21X1 OAI21X1_229 ( .A(_4936_), .B(datapath_1_Instr_18_bF_buf11_), .C(_4937_), .Y(_4938_) );
INVX1 INVX1_79 ( .A(datapath_1_RegisterFile_regfile_mem_0__25_), .Y(_4939_) );
AOI21X1 AOI21X1_250 ( .A(datapath_1_RegisterFile_regfile_mem_4__25_), .B(datapath_1_Instr_18_bF_buf10_), .C(datapath_1_Instr_16_bF_buf20_), .Y(_4940_) );
OAI21X1 OAI21X1_230 ( .A(_4939_), .B(datapath_1_Instr_18_bF_buf9_), .C(_4940_), .Y(_4941_) );
NAND3X1 NAND3X1_133 ( .A(_3566__bF_buf7), .B(_4941_), .C(_4938_), .Y(_4942_) );
INVX1 INVX1_80 ( .A(datapath_1_RegisterFile_regfile_mem_3__25_), .Y(_4943_) );
AOI21X1 AOI21X1_251 ( .A(datapath_1_RegisterFile_regfile_mem_7__25_), .B(datapath_1_Instr_18_bF_buf8_), .C(_3588__bF_buf6), .Y(_4944_) );
OAI21X1 OAI21X1_231 ( .A(_4943_), .B(datapath_1_Instr_18_bF_buf7_), .C(_4944_), .Y(_4945_) );
INVX1 INVX1_81 ( .A(datapath_1_RegisterFile_regfile_mem_2__25_), .Y(_4946_) );
AOI21X1 AOI21X1_252 ( .A(datapath_1_RegisterFile_regfile_mem_6__25_), .B(datapath_1_Instr_18_bF_buf6_), .C(datapath_1_Instr_16_bF_buf19_), .Y(_4947_) );
OAI21X1 OAI21X1_232 ( .A(_4946_), .B(datapath_1_Instr_18_bF_buf5_), .C(_4947_), .Y(_4948_) );
NAND3X1 NAND3X1_134 ( .A(datapath_1_Instr_17_bF_buf31_), .B(_4948_), .C(_4945_), .Y(_4949_) );
AOI21X1 AOI21X1_253 ( .A(_4942_), .B(_4949_), .C(datapath_1_Instr_19_bF_buf2_), .Y(_4950_) );
OAI21X1 OAI21X1_233 ( .A(_4950_), .B(_4935_), .C(_3570__bF_buf2), .Y(_4951_) );
AOI22X1 AOI22X1_42 ( .A(_3565__bF_buf4), .B(_3569__bF_buf4), .C(_4951_), .D(_4920_), .Y(datapath_1_RD2_25_) );
MUX2X1 MUX2X1_97 ( .A(datapath_1_RegisterFile_regfile_mem_9__26_), .B(datapath_1_RegisterFile_regfile_mem_8__26_), .S(datapath_1_Instr_16_bF_buf18_), .Y(_4952_) );
NOR2X1 NOR2X1_103 ( .A(datapath_1_RegisterFile_regfile_mem_11__26_), .B(_3588__bF_buf44), .Y(_4953_) );
OAI21X1 OAI21X1_234 ( .A(datapath_1_RegisterFile_regfile_mem_10__26_), .B(datapath_1_Instr_16_bF_buf17_), .C(datapath_1_Instr_17_bF_buf30_), .Y(_4954_) );
OAI22X1 OAI22X1_86 ( .A(_4954_), .B(_4953_), .C(datapath_1_Instr_17_bF_buf29_), .D(_4952_), .Y(_4955_) );
INVX1 INVX1_82 ( .A(datapath_1_RegisterFile_regfile_mem_15__26_), .Y(_4956_) );
AOI21X1 AOI21X1_254 ( .A(_3588__bF_buf44), .B(datapath_1_RegisterFile_regfile_mem_14__26_), .C(_3566__bF_buf8), .Y(_4957_) );
OAI21X1 OAI21X1_235 ( .A(_4956_), .B(_3588__bF_buf44), .C(_4957_), .Y(_4958_) );
NAND2X1 NAND2X1_264 ( .A(datapath_1_RegisterFile_regfile_mem_12__26_), .B(_3588__bF_buf7), .Y(_4959_) );
AOI21X1 AOI21X1_255 ( .A(datapath_1_RegisterFile_regfile_mem_13__26_), .B(datapath_1_Instr_16_bF_buf16_), .C(datapath_1_Instr_17_bF_buf28_), .Y(_4960_) );
AOI21X1 AOI21X1_256 ( .A(_4959_), .B(_4960_), .C(_3567__bF_buf1), .Y(_4961_) );
AOI22X1 AOI22X1_43 ( .A(_4958_), .B(_4961_), .C(_3567__bF_buf1), .D(_4955_), .Y(_4962_) );
NOR2X1 NOR2X1_104 ( .A(datapath_1_RegisterFile_regfile_mem_0__26_), .B(datapath_1_Instr_16_bF_buf15_), .Y(_4963_) );
OAI21X1 OAI21X1_236 ( .A(datapath_1_RegisterFile_regfile_mem_1__26_), .B(_3588__bF_buf44), .C(_3566__bF_buf6), .Y(_4964_) );
NOR2X1 NOR2X1_105 ( .A(datapath_1_RegisterFile_regfile_mem_3__26_), .B(_3588__bF_buf44), .Y(_4965_) );
OAI21X1 OAI21X1_237 ( .A(datapath_1_RegisterFile_regfile_mem_2__26_), .B(datapath_1_Instr_16_bF_buf14_), .C(datapath_1_Instr_17_bF_buf27_), .Y(_4966_) );
OAI22X1 OAI22X1_87 ( .A(_4965_), .B(_4966_), .C(_4963_), .D(_4964_), .Y(_4967_) );
NOR2X1 NOR2X1_106 ( .A(datapath_1_Instr_18_bF_buf4_), .B(_4967_), .Y(_4968_) );
MUX2X1 MUX2X1_98 ( .A(datapath_1_RegisterFile_regfile_mem_5__26_), .B(datapath_1_RegisterFile_regfile_mem_4__26_), .S(datapath_1_Instr_16_bF_buf13_), .Y(_4969_) );
NOR2X1 NOR2X1_107 ( .A(datapath_1_RegisterFile_regfile_mem_7__26_), .B(_3588__bF_buf18), .Y(_4970_) );
OAI21X1 OAI21X1_238 ( .A(datapath_1_RegisterFile_regfile_mem_6__26_), .B(datapath_1_Instr_16_bF_buf12_), .C(datapath_1_Instr_17_bF_buf26_), .Y(_4971_) );
OAI22X1 OAI22X1_88 ( .A(_4971_), .B(_4970_), .C(datapath_1_Instr_17_bF_buf25_), .D(_4969_), .Y(_4972_) );
OAI21X1 OAI21X1_239 ( .A(_3567__bF_buf1), .B(_4972_), .C(_3571__bF_buf2), .Y(_4973_) );
OAI22X1 OAI22X1_89 ( .A(_3571__bF_buf2), .B(_4962_), .C(_4968_), .D(_4973_), .Y(_4974_) );
NAND2X1 NAND2X1_265 ( .A(_3570__bF_buf0), .B(_4974_), .Y(_4975_) );
INVX1 INVX1_83 ( .A(datapath_1_RegisterFile_regfile_mem_27__26_), .Y(_4976_) );
AOI21X1 AOI21X1_257 ( .A(datapath_1_RegisterFile_regfile_mem_31__26_), .B(datapath_1_Instr_18_bF_buf3_), .C(_3588__bF_buf41), .Y(_4977_) );
OAI21X1 OAI21X1_240 ( .A(_4976_), .B(datapath_1_Instr_18_bF_buf2_), .C(_4977_), .Y(_4978_) );
INVX1 INVX1_84 ( .A(datapath_1_RegisterFile_regfile_mem_26__26_), .Y(_4979_) );
AOI21X1 AOI21X1_258 ( .A(datapath_1_RegisterFile_regfile_mem_30__26_), .B(datapath_1_Instr_18_bF_buf1_), .C(datapath_1_Instr_16_bF_buf11_), .Y(_4980_) );
OAI21X1 OAI21X1_241 ( .A(_4979_), .B(datapath_1_Instr_18_bF_buf0_), .C(_4980_), .Y(_4981_) );
NAND3X1 NAND3X1_135 ( .A(datapath_1_Instr_17_bF_buf24_), .B(_4981_), .C(_4978_), .Y(_4982_) );
INVX1 INVX1_85 ( .A(datapath_1_RegisterFile_regfile_mem_25__26_), .Y(_4983_) );
AOI21X1 AOI21X1_259 ( .A(datapath_1_RegisterFile_regfile_mem_29__26_), .B(datapath_1_Instr_18_bF_buf44_), .C(_3588__bF_buf29), .Y(_4984_) );
OAI21X1 OAI21X1_242 ( .A(_4983_), .B(datapath_1_Instr_18_bF_buf43_), .C(_4984_), .Y(_4985_) );
INVX1 INVX1_86 ( .A(datapath_1_RegisterFile_regfile_mem_24__26_), .Y(_4986_) );
AOI21X1 AOI21X1_260 ( .A(datapath_1_RegisterFile_regfile_mem_28__26_), .B(datapath_1_Instr_18_bF_buf42_), .C(datapath_1_Instr_16_bF_buf10_), .Y(_4987_) );
OAI21X1 OAI21X1_243 ( .A(_4986_), .B(datapath_1_Instr_18_bF_buf41_), .C(_4987_), .Y(_4988_) );
NAND3X1 NAND3X1_136 ( .A(_3566__bF_buf4), .B(_4988_), .C(_4985_), .Y(_4989_) );
AOI21X1 AOI21X1_261 ( .A(_4982_), .B(_4989_), .C(_3571__bF_buf5), .Y(_4990_) );
MUX2X1 MUX2X1_99 ( .A(datapath_1_RegisterFile_regfile_mem_18__26_), .B(datapath_1_RegisterFile_regfile_mem_16__26_), .S(datapath_1_Instr_17_bF_buf23_), .Y(_4991_) );
NAND2X1 NAND2X1_266 ( .A(_3588__bF_buf41), .B(_4991_), .Y(_4992_) );
MUX2X1 MUX2X1_100 ( .A(datapath_1_RegisterFile_regfile_mem_19__26_), .B(datapath_1_RegisterFile_regfile_mem_17__26_), .S(datapath_1_Instr_17_bF_buf22_), .Y(_4993_) );
NAND2X1 NAND2X1_267 ( .A(datapath_1_Instr_16_bF_buf9_), .B(_4993_), .Y(_4994_) );
NAND3X1 NAND3X1_137 ( .A(_3567__bF_buf3), .B(_4992_), .C(_4994_), .Y(_4995_) );
MUX2X1 MUX2X1_101 ( .A(datapath_1_RegisterFile_regfile_mem_22__26_), .B(datapath_1_RegisterFile_regfile_mem_20__26_), .S(datapath_1_Instr_17_bF_buf21_), .Y(_4996_) );
NAND2X1 NAND2X1_268 ( .A(_3588__bF_buf29), .B(_4996_), .Y(_4997_) );
MUX2X1 MUX2X1_102 ( .A(datapath_1_RegisterFile_regfile_mem_23__26_), .B(datapath_1_RegisterFile_regfile_mem_21__26_), .S(datapath_1_Instr_17_bF_buf20_), .Y(_4998_) );
NAND2X1 NAND2X1_269 ( .A(datapath_1_Instr_16_bF_buf8_), .B(_4998_), .Y(_4999_) );
NAND3X1 NAND3X1_138 ( .A(datapath_1_Instr_18_bF_buf40_), .B(_4997_), .C(_4999_), .Y(_5000_) );
AOI21X1 AOI21X1_262 ( .A(_4995_), .B(_5000_), .C(datapath_1_Instr_19_bF_buf1_), .Y(_5001_) );
OAI21X1 OAI21X1_244 ( .A(_4990_), .B(_5001_), .C(datapath_1_Instr_20_bF_buf5_), .Y(_5002_) );
AOI22X1 AOI22X1_44 ( .A(_3565__bF_buf3), .B(_3569__bF_buf3), .C(_5002_), .D(_4975_), .Y(datapath_1_RD2_26_) );
NAND2X1 NAND2X1_270 ( .A(datapath_1_RegisterFile_regfile_mem_27__27_), .B(datapath_1_Instr_16_bF_buf7_), .Y(_5003_) );
NAND2X1 NAND2X1_271 ( .A(datapath_1_RegisterFile_regfile_mem_26__27_), .B(_3588__bF_buf38), .Y(_5004_) );
NAND3X1 NAND3X1_139 ( .A(datapath_1_Instr_17_bF_buf19_), .B(_5003_), .C(_5004_), .Y(_5005_) );
NAND2X1 NAND2X1_272 ( .A(datapath_1_RegisterFile_regfile_mem_25__27_), .B(datapath_1_Instr_16_bF_buf6_), .Y(_5006_) );
AOI21X1 AOI21X1_263 ( .A(_3588__bF_buf38), .B(datapath_1_RegisterFile_regfile_mem_24__27_), .C(datapath_1_Instr_17_bF_buf18_), .Y(_5007_) );
NAND2X1 NAND2X1_273 ( .A(_5006_), .B(_5007_), .Y(_5008_) );
NAND3X1 NAND3X1_140 ( .A(_3567__bF_buf1), .B(_5005_), .C(_5008_), .Y(_5009_) );
NAND2X1 NAND2X1_274 ( .A(datapath_1_RegisterFile_regfile_mem_31__27_), .B(datapath_1_Instr_16_bF_buf5_), .Y(_5010_) );
AOI21X1 AOI21X1_264 ( .A(_3588__bF_buf20), .B(datapath_1_RegisterFile_regfile_mem_30__27_), .C(_3566__bF_buf6), .Y(_5011_) );
NAND2X1 NAND2X1_275 ( .A(_5010_), .B(_5011_), .Y(_5012_) );
AOI21X1 AOI21X1_265 ( .A(datapath_1_RegisterFile_regfile_mem_29__27_), .B(datapath_1_Instr_16_bF_buf4_), .C(datapath_1_Instr_17_bF_buf17_), .Y(_5013_) );
OAI21X1 OAI21X1_245 ( .A(_3312_), .B(datapath_1_Instr_16_bF_buf3_), .C(_5013_), .Y(_5014_) );
NAND3X1 NAND3X1_141 ( .A(datapath_1_Instr_18_bF_buf39_), .B(_5014_), .C(_5012_), .Y(_5015_) );
AOI21X1 AOI21X1_266 ( .A(_5009_), .B(_5015_), .C(_3571__bF_buf2), .Y(_5016_) );
MUX2X1 MUX2X1_103 ( .A(datapath_1_RegisterFile_regfile_mem_18__27_), .B(datapath_1_RegisterFile_regfile_mem_16__27_), .S(datapath_1_Instr_17_bF_buf16_), .Y(_5017_) );
NAND2X1 NAND2X1_276 ( .A(_3588__bF_buf32), .B(_5017_), .Y(_5018_) );
MUX2X1 MUX2X1_104 ( .A(datapath_1_RegisterFile_regfile_mem_19__27_), .B(datapath_1_RegisterFile_regfile_mem_17__27_), .S(datapath_1_Instr_17_bF_buf15_), .Y(_5019_) );
NAND2X1 NAND2X1_277 ( .A(datapath_1_Instr_16_bF_buf2_), .B(_5019_), .Y(_5020_) );
NAND3X1 NAND3X1_142 ( .A(_3567__bF_buf9), .B(_5018_), .C(_5020_), .Y(_5021_) );
MUX2X1 MUX2X1_105 ( .A(datapath_1_RegisterFile_regfile_mem_22__27_), .B(datapath_1_RegisterFile_regfile_mem_20__27_), .S(datapath_1_Instr_17_bF_buf14_), .Y(_5022_) );
NAND2X1 NAND2X1_278 ( .A(_3588__bF_buf23), .B(_5022_), .Y(_5023_) );
MUX2X1 MUX2X1_106 ( .A(datapath_1_RegisterFile_regfile_mem_23__27_), .B(datapath_1_RegisterFile_regfile_mem_21__27_), .S(datapath_1_Instr_17_bF_buf13_), .Y(_5024_) );
NAND2X1 NAND2X1_279 ( .A(datapath_1_Instr_16_bF_buf1_), .B(_5024_), .Y(_5025_) );
NAND3X1 NAND3X1_143 ( .A(datapath_1_Instr_18_bF_buf38_), .B(_5023_), .C(_5025_), .Y(_5026_) );
AOI21X1 AOI21X1_267 ( .A(_5021_), .B(_5026_), .C(datapath_1_Instr_19_bF_buf0_), .Y(_5027_) );
OAI21X1 OAI21X1_246 ( .A(_5027_), .B(_5016_), .C(datapath_1_Instr_20_bF_buf4_), .Y(_5028_) );
INVX1 INVX1_87 ( .A(datapath_1_RegisterFile_regfile_mem_9__27_), .Y(_5029_) );
AOI21X1 AOI21X1_268 ( .A(datapath_1_RegisterFile_regfile_mem_13__27_), .B(datapath_1_Instr_18_bF_buf37_), .C(_3588__bF_buf7), .Y(_5030_) );
OAI21X1 OAI21X1_247 ( .A(_5029_), .B(datapath_1_Instr_18_bF_buf36_), .C(_5030_), .Y(_5031_) );
INVX1 INVX1_88 ( .A(datapath_1_RegisterFile_regfile_mem_8__27_), .Y(_5032_) );
AOI21X1 AOI21X1_269 ( .A(datapath_1_RegisterFile_regfile_mem_12__27_), .B(datapath_1_Instr_18_bF_buf35_), .C(datapath_1_Instr_16_bF_buf0_), .Y(_5033_) );
OAI21X1 OAI21X1_248 ( .A(_5032_), .B(datapath_1_Instr_18_bF_buf34_), .C(_5033_), .Y(_5034_) );
NAND3X1 NAND3X1_144 ( .A(_3566__bF_buf5), .B(_5034_), .C(_5031_), .Y(_5035_) );
INVX1 INVX1_89 ( .A(datapath_1_RegisterFile_regfile_mem_11__27_), .Y(_5036_) );
AOI21X1 AOI21X1_270 ( .A(datapath_1_RegisterFile_regfile_mem_15__27_), .B(datapath_1_Instr_18_bF_buf33_), .C(_3588__bF_buf3), .Y(_5037_) );
OAI21X1 OAI21X1_249 ( .A(_5036_), .B(datapath_1_Instr_18_bF_buf32_), .C(_5037_), .Y(_5038_) );
INVX1 INVX1_90 ( .A(datapath_1_RegisterFile_regfile_mem_10__27_), .Y(_5039_) );
AOI21X1 AOI21X1_271 ( .A(datapath_1_RegisterFile_regfile_mem_14__27_), .B(datapath_1_Instr_18_bF_buf31_), .C(datapath_1_Instr_16_bF_buf55_), .Y(_5040_) );
OAI21X1 OAI21X1_250 ( .A(_5039_), .B(datapath_1_Instr_18_bF_buf30_), .C(_5040_), .Y(_5041_) );
NAND3X1 NAND3X1_145 ( .A(datapath_1_Instr_17_bF_buf12_), .B(_5041_), .C(_5038_), .Y(_5042_) );
AOI21X1 AOI21X1_272 ( .A(_5035_), .B(_5042_), .C(_3571__bF_buf6), .Y(_5043_) );
MUX2X1 MUX2X1_107 ( .A(datapath_1_RegisterFile_regfile_mem_1__27_), .B(datapath_1_RegisterFile_regfile_mem_0__27_), .S(datapath_1_Instr_16_bF_buf54_), .Y(_5044_) );
NOR2X1 NOR2X1_108 ( .A(datapath_1_RegisterFile_regfile_mem_3__27_), .B(_3588__bF_buf3), .Y(_5045_) );
OAI21X1 OAI21X1_251 ( .A(datapath_1_RegisterFile_regfile_mem_2__27_), .B(datapath_1_Instr_16_bF_buf53_), .C(datapath_1_Instr_17_bF_buf11_), .Y(_5046_) );
OAI22X1 OAI22X1_90 ( .A(_5046_), .B(_5045_), .C(datapath_1_Instr_17_bF_buf10_), .D(_5044_), .Y(_5047_) );
NAND2X1 NAND2X1_280 ( .A(_3567__bF_buf6), .B(_5047_), .Y(_5048_) );
MUX2X1 MUX2X1_108 ( .A(datapath_1_RegisterFile_regfile_mem_5__27_), .B(datapath_1_RegisterFile_regfile_mem_4__27_), .S(datapath_1_Instr_16_bF_buf52_), .Y(_5049_) );
NOR2X1 NOR2X1_109 ( .A(datapath_1_RegisterFile_regfile_mem_7__27_), .B(_3588__bF_buf3), .Y(_5050_) );
OAI21X1 OAI21X1_252 ( .A(datapath_1_RegisterFile_regfile_mem_6__27_), .B(datapath_1_Instr_16_bF_buf51_), .C(datapath_1_Instr_17_bF_buf9_), .Y(_5051_) );
OAI22X1 OAI22X1_91 ( .A(_5051_), .B(_5050_), .C(datapath_1_Instr_17_bF_buf8_), .D(_5049_), .Y(_5052_) );
NAND2X1 NAND2X1_281 ( .A(datapath_1_Instr_18_bF_buf29_), .B(_5052_), .Y(_5053_) );
AOI21X1 AOI21X1_273 ( .A(_5048_), .B(_5053_), .C(datapath_1_Instr_19_bF_buf6_), .Y(_5054_) );
OAI21X1 OAI21X1_253 ( .A(_5043_), .B(_5054_), .C(_3570__bF_buf0), .Y(_5055_) );
AOI22X1 AOI22X1_45 ( .A(_3565__bF_buf3), .B(_3569__bF_buf3), .C(_5028_), .D(_5055_), .Y(datapath_1_RD2_27_) );
MUX2X1 MUX2X1_109 ( .A(datapath_1_RegisterFile_regfile_mem_9__28_), .B(datapath_1_RegisterFile_regfile_mem_8__28_), .S(datapath_1_Instr_16_bF_buf50_), .Y(_5056_) );
NOR2X1 NOR2X1_110 ( .A(datapath_1_RegisterFile_regfile_mem_11__28_), .B(_3588__bF_buf34), .Y(_5057_) );
OAI21X1 OAI21X1_254 ( .A(datapath_1_RegisterFile_regfile_mem_10__28_), .B(datapath_1_Instr_16_bF_buf49_), .C(datapath_1_Instr_17_bF_buf7_), .Y(_5058_) );
OAI22X1 OAI22X1_92 ( .A(_5058_), .B(_5057_), .C(datapath_1_Instr_17_bF_buf6_), .D(_5056_), .Y(_5059_) );
AOI21X1 AOI21X1_274 ( .A(_3588__bF_buf12), .B(datapath_1_RegisterFile_regfile_mem_14__28_), .C(_3566__bF_buf2), .Y(_5060_) );
OAI21X1 OAI21X1_255 ( .A(_3384_), .B(_3588__bF_buf12), .C(_5060_), .Y(_5061_) );
NAND2X1 NAND2X1_282 ( .A(datapath_1_RegisterFile_regfile_mem_12__28_), .B(_3588__bF_buf12), .Y(_5062_) );
AOI21X1 AOI21X1_275 ( .A(datapath_1_RegisterFile_regfile_mem_13__28_), .B(datapath_1_Instr_16_bF_buf48_), .C(datapath_1_Instr_17_bF_buf5_), .Y(_5063_) );
AOI21X1 AOI21X1_276 ( .A(_5062_), .B(_5063_), .C(_3567__bF_buf7), .Y(_5064_) );
AOI22X1 AOI22X1_46 ( .A(_5061_), .B(_5064_), .C(_3567__bF_buf7), .D(_5059_), .Y(_5065_) );
NOR2X1 NOR2X1_111 ( .A(datapath_1_RegisterFile_regfile_mem_0__28_), .B(datapath_1_Instr_16_bF_buf47_), .Y(_5066_) );
OAI21X1 OAI21X1_256 ( .A(datapath_1_RegisterFile_regfile_mem_1__28_), .B(_3588__bF_buf40), .C(_3566__bF_buf1), .Y(_5067_) );
NOR2X1 NOR2X1_112 ( .A(datapath_1_RegisterFile_regfile_mem_3__28_), .B(_3588__bF_buf40), .Y(_5068_) );
OAI21X1 OAI21X1_257 ( .A(datapath_1_RegisterFile_regfile_mem_2__28_), .B(datapath_1_Instr_16_bF_buf46_), .C(datapath_1_Instr_17_bF_buf4_), .Y(_5069_) );
OAI22X1 OAI22X1_93 ( .A(_5068_), .B(_5069_), .C(_5066_), .D(_5067_), .Y(_5070_) );
NOR2X1 NOR2X1_113 ( .A(datapath_1_Instr_18_bF_buf28_), .B(_5070_), .Y(_5071_) );
MUX2X1 MUX2X1_110 ( .A(datapath_1_RegisterFile_regfile_mem_5__28_), .B(datapath_1_RegisterFile_regfile_mem_4__28_), .S(datapath_1_Instr_16_bF_buf45_), .Y(_5072_) );
NOR2X1 NOR2X1_114 ( .A(datapath_1_RegisterFile_regfile_mem_7__28_), .B(_3588__bF_buf28), .Y(_5073_) );
OAI21X1 OAI21X1_258 ( .A(datapath_1_RegisterFile_regfile_mem_6__28_), .B(datapath_1_Instr_16_bF_buf44_), .C(datapath_1_Instr_17_bF_buf3_), .Y(_5074_) );
OAI22X1 OAI22X1_94 ( .A(_5074_), .B(_5073_), .C(datapath_1_Instr_17_bF_buf2_), .D(_5072_), .Y(_5075_) );
OAI21X1 OAI21X1_259 ( .A(_3567__bF_buf10), .B(_5075_), .C(_3571__bF_buf0), .Y(_5076_) );
OAI22X1 OAI22X1_95 ( .A(_3571__bF_buf0), .B(_5065_), .C(_5071_), .D(_5076_), .Y(_5077_) );
NAND2X1 NAND2X1_283 ( .A(_3570__bF_buf1), .B(_5077_), .Y(_5078_) );
INVX1 INVX1_91 ( .A(datapath_1_RegisterFile_regfile_mem_19__28_), .Y(_5079_) );
AOI21X1 AOI21X1_277 ( .A(datapath_1_RegisterFile_regfile_mem_23__28_), .B(datapath_1_Instr_18_bF_buf27_), .C(_3588__bF_buf26), .Y(_5080_) );
OAI21X1 OAI21X1_260 ( .A(_5079_), .B(datapath_1_Instr_18_bF_buf26_), .C(_5080_), .Y(_5081_) );
NAND2X1 NAND2X1_284 ( .A(datapath_1_RegisterFile_regfile_mem_18__28_), .B(_3567__bF_buf0), .Y(_5082_) );
AOI21X1 AOI21X1_278 ( .A(datapath_1_RegisterFile_regfile_mem_22__28_), .B(datapath_1_Instr_18_bF_buf25_), .C(datapath_1_Instr_16_bF_buf43_), .Y(_5083_) );
AOI21X1 AOI21X1_279 ( .A(_5082_), .B(_5083_), .C(_3566__bF_buf9), .Y(_5084_) );
INVX1 INVX1_92 ( .A(datapath_1_RegisterFile_regfile_mem_17__28_), .Y(_5085_) );
AOI21X1 AOI21X1_280 ( .A(datapath_1_RegisterFile_regfile_mem_21__28_), .B(datapath_1_Instr_18_bF_buf24_), .C(_3588__bF_buf26), .Y(_5086_) );
OAI21X1 OAI21X1_261 ( .A(_5085_), .B(datapath_1_Instr_18_bF_buf23_), .C(_5086_), .Y(_5087_) );
NAND2X1 NAND2X1_285 ( .A(datapath_1_RegisterFile_regfile_mem_16__28_), .B(_3567__bF_buf0), .Y(_5088_) );
AOI21X1 AOI21X1_281 ( .A(datapath_1_RegisterFile_regfile_mem_20__28_), .B(datapath_1_Instr_18_bF_buf22_), .C(datapath_1_Instr_16_bF_buf42_), .Y(_5089_) );
AOI21X1 AOI21X1_282 ( .A(_5088_), .B(_5089_), .C(datapath_1_Instr_17_bF_buf1_), .Y(_5090_) );
AOI22X1 AOI22X1_47 ( .A(_5084_), .B(_5081_), .C(_5087_), .D(_5090_), .Y(_5091_) );
NOR2X1 NOR2X1_115 ( .A(datapath_1_RegisterFile_regfile_mem_24__28_), .B(datapath_1_Instr_16_bF_buf41_), .Y(_5092_) );
OAI21X1 OAI21X1_262 ( .A(datapath_1_RegisterFile_regfile_mem_25__28_), .B(_3588__bF_buf0), .C(_3566__bF_buf9), .Y(_5093_) );
NOR2X1 NOR2X1_116 ( .A(datapath_1_RegisterFile_regfile_mem_27__28_), .B(_3588__bF_buf0), .Y(_5094_) );
OAI21X1 OAI21X1_263 ( .A(datapath_1_RegisterFile_regfile_mem_26__28_), .B(datapath_1_Instr_16_bF_buf40_), .C(datapath_1_Instr_17_bF_buf0_), .Y(_5095_) );
OAI22X1 OAI22X1_96 ( .A(_5094_), .B(_5095_), .C(_5092_), .D(_5093_), .Y(_5096_) );
NOR2X1 NOR2X1_117 ( .A(datapath_1_Instr_18_bF_buf21_), .B(_5096_), .Y(_5097_) );
MUX2X1 MUX2X1_111 ( .A(datapath_1_RegisterFile_regfile_mem_29__28_), .B(datapath_1_RegisterFile_regfile_mem_28__28_), .S(datapath_1_Instr_16_bF_buf39_), .Y(_5098_) );
NOR2X1 NOR2X1_118 ( .A(datapath_1_RegisterFile_regfile_mem_31__28_), .B(_3588__bF_buf14), .Y(_5099_) );
OAI21X1 OAI21X1_264 ( .A(datapath_1_RegisterFile_regfile_mem_30__28_), .B(datapath_1_Instr_16_bF_buf38_), .C(datapath_1_Instr_17_bF_buf50_), .Y(_5100_) );
OAI22X1 OAI22X1_97 ( .A(_5100_), .B(_5099_), .C(datapath_1_Instr_17_bF_buf49_), .D(_5098_), .Y(_5101_) );
OAI21X1 OAI21X1_265 ( .A(_3567__bF_buf5), .B(_5101_), .C(datapath_1_Instr_19_bF_buf5_), .Y(_5102_) );
OAI22X1 OAI22X1_98 ( .A(datapath_1_Instr_19_bF_buf4_), .B(_5091_), .C(_5097_), .D(_5102_), .Y(_5103_) );
NAND2X1 NAND2X1_286 ( .A(datapath_1_Instr_20_bF_buf3_), .B(_5103_), .Y(_5104_) );
AOI22X1 AOI22X1_48 ( .A(_3565__bF_buf0), .B(_3569__bF_buf0), .C(_5104_), .D(_5078_), .Y(datapath_1_RD2_28_) );
NAND2X1 NAND2X1_287 ( .A(datapath_1_RegisterFile_regfile_mem_27__29_), .B(datapath_1_Instr_16_bF_buf37_), .Y(_5105_) );
NAND2X1 NAND2X1_288 ( .A(datapath_1_RegisterFile_regfile_mem_26__29_), .B(_3588__bF_buf13), .Y(_5106_) );
NAND3X1 NAND3X1_146 ( .A(datapath_1_Instr_17_bF_buf48_), .B(_5105_), .C(_5106_), .Y(_5107_) );
NAND2X1 NAND2X1_289 ( .A(datapath_1_RegisterFile_regfile_mem_25__29_), .B(datapath_1_Instr_16_bF_buf36_), .Y(_5108_) );
AOI21X1 AOI21X1_283 ( .A(_3588__bF_buf13), .B(datapath_1_RegisterFile_regfile_mem_24__29_), .C(datapath_1_Instr_17_bF_buf47_), .Y(_5109_) );
NAND2X1 NAND2X1_290 ( .A(_5108_), .B(_5109_), .Y(_5110_) );
NAND3X1 NAND3X1_147 ( .A(_3567__bF_buf5), .B(_5107_), .C(_5110_), .Y(_5111_) );
NAND2X1 NAND2X1_291 ( .A(datapath_1_RegisterFile_regfile_mem_31__29_), .B(datapath_1_Instr_16_bF_buf35_), .Y(_5112_) );
AOI21X1 AOI21X1_284 ( .A(_3588__bF_buf39), .B(datapath_1_RegisterFile_regfile_mem_30__29_), .C(_3566__bF_buf10), .Y(_5113_) );
NAND2X1 NAND2X1_292 ( .A(_5112_), .B(_5113_), .Y(_5114_) );
INVX1 INVX1_93 ( .A(datapath_1_RegisterFile_regfile_mem_28__29_), .Y(_5115_) );
AOI21X1 AOI21X1_285 ( .A(datapath_1_RegisterFile_regfile_mem_29__29_), .B(datapath_1_Instr_16_bF_buf34_), .C(datapath_1_Instr_17_bF_buf46_), .Y(_5116_) );
OAI21X1 OAI21X1_266 ( .A(_5115_), .B(datapath_1_Instr_16_bF_buf33_), .C(_5116_), .Y(_5117_) );
NAND3X1 NAND3X1_148 ( .A(datapath_1_Instr_18_bF_buf20_), .B(_5117_), .C(_5114_), .Y(_5118_) );
AOI21X1 AOI21X1_286 ( .A(_5111_), .B(_5118_), .C(_3571__bF_buf7), .Y(_5119_) );
MUX2X1 MUX2X1_112 ( .A(datapath_1_RegisterFile_regfile_mem_18__29_), .B(datapath_1_RegisterFile_regfile_mem_16__29_), .S(datapath_1_Instr_17_bF_buf45_), .Y(_5120_) );
NAND2X1 NAND2X1_293 ( .A(_3588__bF_buf39), .B(_5120_), .Y(_5121_) );
MUX2X1 MUX2X1_113 ( .A(datapath_1_RegisterFile_regfile_mem_19__29_), .B(datapath_1_RegisterFile_regfile_mem_17__29_), .S(datapath_1_Instr_17_bF_buf44_), .Y(_5122_) );
NAND2X1 NAND2X1_294 ( .A(datapath_1_Instr_16_bF_buf32_), .B(_5122_), .Y(_5123_) );
NAND3X1 NAND3X1_149 ( .A(_3567__bF_buf2), .B(_5121_), .C(_5123_), .Y(_5124_) );
MUX2X1 MUX2X1_114 ( .A(datapath_1_RegisterFile_regfile_mem_22__29_), .B(datapath_1_RegisterFile_regfile_mem_20__29_), .S(datapath_1_Instr_17_bF_buf43_), .Y(_5125_) );
NAND2X1 NAND2X1_295 ( .A(_3588__bF_buf15), .B(_5125_), .Y(_5126_) );
MUX2X1 MUX2X1_115 ( .A(datapath_1_RegisterFile_regfile_mem_23__29_), .B(datapath_1_RegisterFile_regfile_mem_21__29_), .S(datapath_1_Instr_17_bF_buf42_), .Y(_5127_) );
NAND2X1 NAND2X1_296 ( .A(datapath_1_Instr_16_bF_buf31_), .B(_5127_), .Y(_5128_) );
NAND3X1 NAND3X1_150 ( .A(datapath_1_Instr_18_bF_buf19_), .B(_5126_), .C(_5128_), .Y(_5129_) );
AOI21X1 AOI21X1_287 ( .A(_5124_), .B(_5129_), .C(datapath_1_Instr_19_bF_buf3_), .Y(_5130_) );
OAI21X1 OAI21X1_267 ( .A(_5130_), .B(_5119_), .C(datapath_1_Instr_20_bF_buf2_), .Y(_5131_) );
MUX2X1 MUX2X1_116 ( .A(datapath_1_RegisterFile_regfile_mem_9__29_), .B(datapath_1_RegisterFile_regfile_mem_8__29_), .S(datapath_1_Instr_16_bF_buf30_), .Y(_5132_) );
NOR2X1 NOR2X1_119 ( .A(datapath_1_RegisterFile_regfile_mem_11__29_), .B(_3588__bF_buf12), .Y(_5133_) );
OAI21X1 OAI21X1_268 ( .A(datapath_1_RegisterFile_regfile_mem_10__29_), .B(datapath_1_Instr_16_bF_buf29_), .C(datapath_1_Instr_17_bF_buf41_), .Y(_5134_) );
OAI22X1 OAI22X1_99 ( .A(_5134_), .B(_5133_), .C(datapath_1_Instr_17_bF_buf40_), .D(_5132_), .Y(_5135_) );
INVX1 INVX1_94 ( .A(datapath_1_RegisterFile_regfile_mem_15__29_), .Y(_5136_) );
AOI21X1 AOI21X1_288 ( .A(_3588__bF_buf12), .B(datapath_1_RegisterFile_regfile_mem_14__29_), .C(_3566__bF_buf1), .Y(_5137_) );
OAI21X1 OAI21X1_269 ( .A(_5136_), .B(_3588__bF_buf12), .C(_5137_), .Y(_5138_) );
NAND2X1 NAND2X1_297 ( .A(datapath_1_RegisterFile_regfile_mem_12__29_), .B(_3588__bF_buf12), .Y(_5139_) );
AOI21X1 AOI21X1_289 ( .A(datapath_1_RegisterFile_regfile_mem_13__29_), .B(datapath_1_Instr_16_bF_buf28_), .C(datapath_1_Instr_17_bF_buf39_), .Y(_5140_) );
AOI21X1 AOI21X1_290 ( .A(_5139_), .B(_5140_), .C(_3567__bF_buf10), .Y(_5141_) );
AOI22X1 AOI22X1_49 ( .A(_5138_), .B(_5141_), .C(_3567__bF_buf10), .D(_5135_), .Y(_5142_) );
NOR2X1 NOR2X1_120 ( .A(datapath_1_RegisterFile_regfile_mem_0__29_), .B(datapath_1_Instr_16_bF_buf27_), .Y(_5143_) );
OAI21X1 OAI21X1_270 ( .A(datapath_1_RegisterFile_regfile_mem_1__29_), .B(_3588__bF_buf42), .C(_3566__bF_buf7), .Y(_5144_) );
NOR2X1 NOR2X1_121 ( .A(datapath_1_RegisterFile_regfile_mem_3__29_), .B(_3588__bF_buf42), .Y(_5145_) );
OAI21X1 OAI21X1_271 ( .A(datapath_1_RegisterFile_regfile_mem_2__29_), .B(datapath_1_Instr_16_bF_buf26_), .C(datapath_1_Instr_17_bF_buf38_), .Y(_5146_) );
OAI22X1 OAI22X1_100 ( .A(_5145_), .B(_5146_), .C(_5143_), .D(_5144_), .Y(_5147_) );
NOR2X1 NOR2X1_122 ( .A(datapath_1_Instr_18_bF_buf18_), .B(_5147_), .Y(_5148_) );
MUX2X1 MUX2X1_117 ( .A(datapath_1_RegisterFile_regfile_mem_5__29_), .B(datapath_1_RegisterFile_regfile_mem_4__29_), .S(datapath_1_Instr_16_bF_buf25_), .Y(_5149_) );
NOR2X1 NOR2X1_123 ( .A(datapath_1_RegisterFile_regfile_mem_7__29_), .B(_3588__bF_buf42), .Y(_5150_) );
OAI21X1 OAI21X1_272 ( .A(datapath_1_RegisterFile_regfile_mem_6__29_), .B(datapath_1_Instr_16_bF_buf24_), .C(datapath_1_Instr_17_bF_buf37_), .Y(_5151_) );
OAI22X1 OAI22X1_101 ( .A(_5151_), .B(_5150_), .C(datapath_1_Instr_17_bF_buf36_), .D(_5149_), .Y(_5152_) );
OAI21X1 OAI21X1_273 ( .A(_3567__bF_buf10), .B(_5152_), .C(_3571__bF_buf4), .Y(_5153_) );
OAI22X1 OAI22X1_102 ( .A(_3571__bF_buf4), .B(_5142_), .C(_5148_), .D(_5153_), .Y(_5154_) );
NAND2X1 NAND2X1_298 ( .A(_3570__bF_buf1), .B(_5154_), .Y(_5155_) );
AOI22X1 AOI22X1_50 ( .A(_3565__bF_buf0), .B(_3569__bF_buf0), .C(_5131_), .D(_5155_), .Y(datapath_1_RD2_29_) );
NAND2X1 NAND2X1_299 ( .A(datapath_1_RegisterFile_regfile_mem_27__30_), .B(datapath_1_Instr_16_bF_buf23_), .Y(_5156_) );
NAND2X1 NAND2X1_300 ( .A(datapath_1_RegisterFile_regfile_mem_26__30_), .B(_3588__bF_buf37), .Y(_5157_) );
NAND3X1 NAND3X1_151 ( .A(datapath_1_Instr_17_bF_buf35_), .B(_5156_), .C(_5157_), .Y(_5158_) );
NAND2X1 NAND2X1_301 ( .A(datapath_1_RegisterFile_regfile_mem_25__30_), .B(datapath_1_Instr_16_bF_buf22_), .Y(_5159_) );
AOI21X1 AOI21X1_291 ( .A(_3588__bF_buf5), .B(datapath_1_RegisterFile_regfile_mem_24__30_), .C(datapath_1_Instr_17_bF_buf34_), .Y(_5160_) );
NAND2X1 NAND2X1_302 ( .A(_5159_), .B(_5160_), .Y(_5161_) );
NAND3X1 NAND3X1_152 ( .A(_3567__bF_buf3), .B(_5158_), .C(_5161_), .Y(_5162_) );
NAND2X1 NAND2X1_303 ( .A(datapath_1_RegisterFile_regfile_mem_31__30_), .B(datapath_1_Instr_16_bF_buf21_), .Y(_5163_) );
AOI21X1 AOI21X1_292 ( .A(_3588__bF_buf16), .B(datapath_1_RegisterFile_regfile_mem_30__30_), .C(_3566__bF_buf4), .Y(_5164_) );
NAND2X1 NAND2X1_304 ( .A(_5163_), .B(_5164_), .Y(_5165_) );
INVX1 INVX1_95 ( .A(datapath_1_RegisterFile_regfile_mem_28__30_), .Y(_5166_) );
AOI21X1 AOI21X1_293 ( .A(datapath_1_RegisterFile_regfile_mem_29__30_), .B(datapath_1_Instr_16_bF_buf20_), .C(datapath_1_Instr_17_bF_buf33_), .Y(_5167_) );
OAI21X1 OAI21X1_274 ( .A(_5166_), .B(datapath_1_Instr_16_bF_buf19_), .C(_5167_), .Y(_5168_) );
NAND3X1 NAND3X1_153 ( .A(datapath_1_Instr_18_bF_buf17_), .B(_5168_), .C(_5165_), .Y(_5169_) );
AOI21X1 AOI21X1_294 ( .A(_5162_), .B(_5169_), .C(_3571__bF_buf5), .Y(_5170_) );
MUX2X1 MUX2X1_118 ( .A(datapath_1_RegisterFile_regfile_mem_17__30_), .B(datapath_1_RegisterFile_regfile_mem_16__30_), .S(datapath_1_Instr_16_bF_buf18_), .Y(_5171_) );
NOR2X1 NOR2X1_124 ( .A(datapath_1_RegisterFile_regfile_mem_19__30_), .B(_3588__bF_buf41), .Y(_5172_) );
OAI21X1 OAI21X1_275 ( .A(datapath_1_RegisterFile_regfile_mem_18__30_), .B(datapath_1_Instr_16_bF_buf17_), .C(datapath_1_Instr_17_bF_buf32_), .Y(_5173_) );
OAI22X1 OAI22X1_103 ( .A(_5173_), .B(_5172_), .C(datapath_1_Instr_17_bF_buf31_), .D(_5171_), .Y(_5174_) );
NAND2X1 NAND2X1_305 ( .A(_3567__bF_buf3), .B(_5174_), .Y(_5175_) );
MUX2X1 MUX2X1_119 ( .A(datapath_1_RegisterFile_regfile_mem_21__30_), .B(datapath_1_RegisterFile_regfile_mem_20__30_), .S(datapath_1_Instr_16_bF_buf16_), .Y(_5176_) );
NOR2X1 NOR2X1_125 ( .A(datapath_1_RegisterFile_regfile_mem_23__30_), .B(_3588__bF_buf41), .Y(_5177_) );
OAI21X1 OAI21X1_276 ( .A(datapath_1_RegisterFile_regfile_mem_22__30_), .B(datapath_1_Instr_16_bF_buf15_), .C(datapath_1_Instr_17_bF_buf30_), .Y(_5178_) );
OAI22X1 OAI22X1_104 ( .A(_5178_), .B(_5177_), .C(datapath_1_Instr_17_bF_buf29_), .D(_5176_), .Y(_5179_) );
NAND2X1 NAND2X1_306 ( .A(datapath_1_Instr_18_bF_buf16_), .B(_5179_), .Y(_5180_) );
AOI21X1 AOI21X1_295 ( .A(_5175_), .B(_5180_), .C(datapath_1_Instr_19_bF_buf2_), .Y(_5181_) );
OAI21X1 OAI21X1_277 ( .A(_5170_), .B(_5181_), .C(datapath_1_Instr_20_bF_buf1_), .Y(_5182_) );
NAND2X1 NAND2X1_307 ( .A(datapath_1_RegisterFile_regfile_mem_11__30_), .B(datapath_1_Instr_17_bF_buf28_), .Y(_5183_) );
NAND2X1 NAND2X1_308 ( .A(datapath_1_RegisterFile_regfile_mem_9__30_), .B(_3566__bF_buf5), .Y(_5184_) );
NAND3X1 NAND3X1_154 ( .A(datapath_1_Instr_16_bF_buf14_), .B(_5183_), .C(_5184_), .Y(_5185_) );
NAND2X1 NAND2X1_309 ( .A(datapath_1_RegisterFile_regfile_mem_10__30_), .B(datapath_1_Instr_17_bF_buf27_), .Y(_5186_) );
AOI21X1 AOI21X1_296 ( .A(_3566__bF_buf5), .B(datapath_1_RegisterFile_regfile_mem_8__30_), .C(datapath_1_Instr_16_bF_buf13_), .Y(_5187_) );
NAND2X1 NAND2X1_310 ( .A(_5186_), .B(_5187_), .Y(_5188_) );
NAND3X1 NAND3X1_155 ( .A(_3567__bF_buf8), .B(_5185_), .C(_5188_), .Y(_5189_) );
NAND2X1 NAND2X1_311 ( .A(datapath_1_RegisterFile_regfile_mem_15__30_), .B(datapath_1_Instr_17_bF_buf26_), .Y(_5190_) );
NAND2X1 NAND2X1_312 ( .A(datapath_1_RegisterFile_regfile_mem_13__30_), .B(_3566__bF_buf5), .Y(_5191_) );
NAND3X1 NAND3X1_156 ( .A(datapath_1_Instr_16_bF_buf12_), .B(_5190_), .C(_5191_), .Y(_5192_) );
NAND2X1 NAND2X1_313 ( .A(datapath_1_RegisterFile_regfile_mem_14__30_), .B(datapath_1_Instr_17_bF_buf25_), .Y(_5193_) );
AOI21X1 AOI21X1_297 ( .A(_3566__bF_buf5), .B(datapath_1_RegisterFile_regfile_mem_12__30_), .C(datapath_1_Instr_16_bF_buf11_), .Y(_5194_) );
NAND2X1 NAND2X1_314 ( .A(_5193_), .B(_5194_), .Y(_5195_) );
NAND3X1 NAND3X1_157 ( .A(datapath_1_Instr_18_bF_buf15_), .B(_5192_), .C(_5195_), .Y(_5196_) );
AOI21X1 AOI21X1_298 ( .A(_5189_), .B(_5196_), .C(_3571__bF_buf3), .Y(_5197_) );
INVX1 INVX1_96 ( .A(datapath_1_RegisterFile_regfile_mem_1__30_), .Y(_5198_) );
AOI21X1 AOI21X1_299 ( .A(datapath_1_RegisterFile_regfile_mem_5__30_), .B(datapath_1_Instr_18_bF_buf14_), .C(_3588__bF_buf37), .Y(_5199_) );
OAI21X1 OAI21X1_278 ( .A(_5198_), .B(datapath_1_Instr_18_bF_buf13_), .C(_5199_), .Y(_5200_) );
INVX1 INVX1_97 ( .A(datapath_1_RegisterFile_regfile_mem_0__30_), .Y(_5201_) );
AOI21X1 AOI21X1_300 ( .A(datapath_1_RegisterFile_regfile_mem_4__30_), .B(datapath_1_Instr_18_bF_buf12_), .C(datapath_1_Instr_16_bF_buf10_), .Y(_5202_) );
OAI21X1 OAI21X1_279 ( .A(_5201_), .B(datapath_1_Instr_18_bF_buf11_), .C(_5202_), .Y(_5203_) );
NAND3X1 NAND3X1_158 ( .A(_3566__bF_buf4), .B(_5203_), .C(_5200_), .Y(_5204_) );
INVX1 INVX1_98 ( .A(datapath_1_RegisterFile_regfile_mem_3__30_), .Y(_5205_) );
AOI21X1 AOI21X1_301 ( .A(datapath_1_RegisterFile_regfile_mem_7__30_), .B(datapath_1_Instr_18_bF_buf10_), .C(_3588__bF_buf18), .Y(_5206_) );
OAI21X1 OAI21X1_280 ( .A(_5205_), .B(datapath_1_Instr_18_bF_buf9_), .C(_5206_), .Y(_5207_) );
INVX1 INVX1_99 ( .A(datapath_1_RegisterFile_regfile_mem_2__30_), .Y(_5208_) );
AOI21X1 AOI21X1_302 ( .A(datapath_1_RegisterFile_regfile_mem_6__30_), .B(datapath_1_Instr_18_bF_buf8_), .C(datapath_1_Instr_16_bF_buf9_), .Y(_5209_) );
OAI21X1 OAI21X1_281 ( .A(_5208_), .B(datapath_1_Instr_18_bF_buf7_), .C(_5209_), .Y(_5210_) );
NAND3X1 NAND3X1_159 ( .A(datapath_1_Instr_17_bF_buf24_), .B(_5210_), .C(_5207_), .Y(_5211_) );
AOI21X1 AOI21X1_303 ( .A(_5204_), .B(_5211_), .C(datapath_1_Instr_19_bF_buf1_), .Y(_5212_) );
OAI21X1 OAI21X1_282 ( .A(_5212_), .B(_5197_), .C(_3570__bF_buf4), .Y(_5213_) );
AOI22X1 AOI22X1_51 ( .A(_3565__bF_buf2), .B(_3569__bF_buf2), .C(_5213_), .D(_5182_), .Y(datapath_1_RD2_30_) );
NAND2X1 NAND2X1_315 ( .A(datapath_1_RegisterFile_regfile_mem_27__31_), .B(datapath_1_Instr_16_bF_buf8_), .Y(_5214_) );
NAND2X1 NAND2X1_316 ( .A(datapath_1_RegisterFile_regfile_mem_26__31_), .B(_3588__bF_buf38), .Y(_5215_) );
NAND3X1 NAND3X1_160 ( .A(datapath_1_Instr_17_bF_buf23_), .B(_5214_), .C(_5215_), .Y(_5216_) );
NAND2X1 NAND2X1_317 ( .A(datapath_1_RegisterFile_regfile_mem_25__31_), .B(datapath_1_Instr_16_bF_buf7_), .Y(_5217_) );
AOI21X1 AOI21X1_304 ( .A(_3588__bF_buf20), .B(datapath_1_RegisterFile_regfile_mem_24__31_), .C(datapath_1_Instr_17_bF_buf22_), .Y(_5218_) );
NAND2X1 NAND2X1_318 ( .A(_5217_), .B(_5218_), .Y(_5219_) );
NAND3X1 NAND3X1_161 ( .A(_3567__bF_buf1), .B(_5216_), .C(_5219_), .Y(_5220_) );
NAND2X1 NAND2X1_319 ( .A(datapath_1_RegisterFile_regfile_mem_31__31_), .B(datapath_1_Instr_16_bF_buf6_), .Y(_5221_) );
AOI21X1 AOI21X1_305 ( .A(_3588__bF_buf38), .B(datapath_1_RegisterFile_regfile_mem_30__31_), .C(_3566__bF_buf6), .Y(_5222_) );
NAND2X1 NAND2X1_320 ( .A(_5221_), .B(_5222_), .Y(_5223_) );
AOI21X1 AOI21X1_306 ( .A(datapath_1_RegisterFile_regfile_mem_29__31_), .B(datapath_1_Instr_16_bF_buf5_), .C(datapath_1_Instr_17_bF_buf21_), .Y(_5224_) );
OAI21X1 OAI21X1_283 ( .A(_3521_), .B(datapath_1_Instr_16_bF_buf4_), .C(_5224_), .Y(_5225_) );
NAND3X1 NAND3X1_162 ( .A(datapath_1_Instr_18_bF_buf6_), .B(_5225_), .C(_5223_), .Y(_5226_) );
AOI21X1 AOI21X1_307 ( .A(_5220_), .B(_5226_), .C(_3571__bF_buf2), .Y(_5227_) );
MUX2X1 MUX2X1_120 ( .A(datapath_1_RegisterFile_regfile_mem_18__31_), .B(datapath_1_RegisterFile_regfile_mem_16__31_), .S(datapath_1_Instr_17_bF_buf20_), .Y(_5228_) );
NAND2X1 NAND2X1_321 ( .A(_3588__bF_buf32), .B(_5228_), .Y(_5229_) );
MUX2X1 MUX2X1_121 ( .A(datapath_1_RegisterFile_regfile_mem_19__31_), .B(datapath_1_RegisterFile_regfile_mem_17__31_), .S(datapath_1_Instr_17_bF_buf19_), .Y(_5230_) );
NAND2X1 NAND2X1_322 ( .A(datapath_1_Instr_16_bF_buf3_), .B(_5230_), .Y(_5231_) );
NAND3X1 NAND3X1_163 ( .A(_3567__bF_buf9), .B(_5229_), .C(_5231_), .Y(_5232_) );
MUX2X1 MUX2X1_122 ( .A(datapath_1_RegisterFile_regfile_mem_22__31_), .B(datapath_1_RegisterFile_regfile_mem_20__31_), .S(datapath_1_Instr_17_bF_buf18_), .Y(_5233_) );
NAND2X1 NAND2X1_323 ( .A(_3588__bF_buf32), .B(_5233_), .Y(_5234_) );
MUX2X1 MUX2X1_123 ( .A(datapath_1_RegisterFile_regfile_mem_23__31_), .B(datapath_1_RegisterFile_regfile_mem_21__31_), .S(datapath_1_Instr_17_bF_buf17_), .Y(_5235_) );
NAND2X1 NAND2X1_324 ( .A(datapath_1_Instr_16_bF_buf2_), .B(_5235_), .Y(_5236_) );
NAND3X1 NAND3X1_164 ( .A(datapath_1_Instr_18_bF_buf5_), .B(_5234_), .C(_5236_), .Y(_5237_) );
AOI21X1 AOI21X1_308 ( .A(_5232_), .B(_5237_), .C(datapath_1_Instr_19_bF_buf0_), .Y(_5238_) );
OAI21X1 OAI21X1_284 ( .A(_5238_), .B(_5227_), .C(datapath_1_Instr_20_bF_buf0_), .Y(_5239_) );
MUX2X1 MUX2X1_124 ( .A(datapath_1_RegisterFile_regfile_mem_9__31_), .B(datapath_1_RegisterFile_regfile_mem_8__31_), .S(datapath_1_Instr_16_bF_buf1_), .Y(_5240_) );
NOR2X1 NOR2X1_126 ( .A(datapath_1_RegisterFile_regfile_mem_11__31_), .B(_3588__bF_buf7), .Y(_5241_) );
OAI21X1 OAI21X1_285 ( .A(datapath_1_RegisterFile_regfile_mem_10__31_), .B(datapath_1_Instr_16_bF_buf0_), .C(datapath_1_Instr_17_bF_buf16_), .Y(_5242_) );
OAI22X1 OAI22X1_105 ( .A(_5242_), .B(_5241_), .C(datapath_1_Instr_17_bF_buf15_), .D(_5240_), .Y(_5243_) );
INVX1 INVX1_100 ( .A(datapath_1_RegisterFile_regfile_mem_15__31_), .Y(_5244_) );
AOI21X1 AOI21X1_309 ( .A(_3588__bF_buf7), .B(datapath_1_RegisterFile_regfile_mem_14__31_), .C(_3566__bF_buf8), .Y(_5245_) );
OAI21X1 OAI21X1_286 ( .A(_5244_), .B(_3588__bF_buf7), .C(_5245_), .Y(_5246_) );
NAND2X1 NAND2X1_325 ( .A(datapath_1_RegisterFile_regfile_mem_12__31_), .B(_3588__bF_buf7), .Y(_5247_) );
AOI21X1 AOI21X1_310 ( .A(datapath_1_RegisterFile_regfile_mem_13__31_), .B(datapath_1_Instr_16_bF_buf55_), .C(datapath_1_Instr_17_bF_buf14_), .Y(_5248_) );
AOI21X1 AOI21X1_311 ( .A(_5247_), .B(_5248_), .C(_3567__bF_buf6), .Y(_5249_) );
AOI22X1 AOI22X1_52 ( .A(_5246_), .B(_5249_), .C(_3567__bF_buf6), .D(_5243_), .Y(_5250_) );
NOR2X1 NOR2X1_127 ( .A(datapath_1_RegisterFile_regfile_mem_0__31_), .B(datapath_1_Instr_16_bF_buf54_), .Y(_5251_) );
OAI21X1 OAI21X1_287 ( .A(datapath_1_RegisterFile_regfile_mem_1__31_), .B(_3588__bF_buf30), .C(_3566__bF_buf6), .Y(_5252_) );
NOR2X1 NOR2X1_128 ( .A(datapath_1_RegisterFile_regfile_mem_3__31_), .B(_3588__bF_buf30), .Y(_5253_) );
OAI21X1 OAI21X1_288 ( .A(datapath_1_RegisterFile_regfile_mem_2__31_), .B(datapath_1_Instr_16_bF_buf53_), .C(datapath_1_Instr_17_bF_buf13_), .Y(_5254_) );
OAI22X1 OAI22X1_106 ( .A(_5253_), .B(_5254_), .C(_5251_), .D(_5252_), .Y(_5255_) );
NOR2X1 NOR2X1_129 ( .A(datapath_1_Instr_18_bF_buf4_), .B(_5255_), .Y(_5256_) );
MUX2X1 MUX2X1_125 ( .A(datapath_1_RegisterFile_regfile_mem_5__31_), .B(datapath_1_RegisterFile_regfile_mem_4__31_), .S(datapath_1_Instr_16_bF_buf52_), .Y(_5257_) );
NOR2X1 NOR2X1_130 ( .A(datapath_1_RegisterFile_regfile_mem_7__31_), .B(_3588__bF_buf35), .Y(_5258_) );
OAI21X1 OAI21X1_289 ( .A(datapath_1_RegisterFile_regfile_mem_6__31_), .B(datapath_1_Instr_16_bF_buf51_), .C(datapath_1_Instr_17_bF_buf12_), .Y(_5259_) );
OAI22X1 OAI22X1_107 ( .A(_5259_), .B(_5258_), .C(datapath_1_Instr_17_bF_buf11_), .D(_5257_), .Y(_5260_) );
OAI21X1 OAI21X1_290 ( .A(_3567__bF_buf6), .B(_5260_), .C(_3571__bF_buf6), .Y(_5261_) );
OAI22X1 OAI22X1_108 ( .A(_3571__bF_buf6), .B(_5250_), .C(_5256_), .D(_5261_), .Y(_5262_) );
NAND2X1 NAND2X1_326 ( .A(_3570__bF_buf4), .B(_5262_), .Y(_5263_) );
AOI22X1 AOI22X1_53 ( .A(_3565__bF_buf3), .B(_3569__bF_buf3), .C(_5239_), .D(_5263_), .Y(datapath_1_RD2_31_) );
INVX1 INVX1_101 ( .A(datapath_1_A3_3_), .Y(_5264_) );
INVX1 INVX1_102 ( .A(rst_bF_buf8), .Y(_5265_) );
NAND2X1 NAND2X1_327 ( .A(RegWrite), .B(_5265__bF_buf47), .Y(_5266_) );
NOR2X1 NOR2X1_131 ( .A(datapath_1_A3_4_), .B(_5266_), .Y(_5267_) );
NAND2X1 NAND2X1_328 ( .A(_5264_), .B(_5267_), .Y(_5268_) );
NOR2X1 NOR2X1_132 ( .A(datapath_1_A3_2_), .B(_5268_), .Y(_5269_) );
INVX1 INVX1_103 ( .A(datapath_1_A3_0_), .Y(_5270_) );
INVX1 INVX1_104 ( .A(datapath_1_A3_1_), .Y(_5271_) );
INVX1 INVX1_105 ( .A(_5266_), .Y(_5272_) );
NAND3X1 NAND3X1_165 ( .A(_5270_), .B(_5271_), .C(_5272__bF_buf2), .Y(_5273_) );
INVX1 INVX1_106 ( .A(_5273_), .Y(_5274_) );
NAND2X1 NAND2X1_329 ( .A(_5274_), .B(_5269_), .Y(_5275_) );
NAND2X1 NAND2X1_330 ( .A(datapath_1_RegisterFile_dataWrite_0_), .B(_5272__bF_buf5), .Y(_5276_) );
NAND3X1 NAND3X1_166 ( .A(datapath_1_RegisterFile_regfile_mem_0__0_), .B(_5265__bF_buf31), .C(_5275__bF_buf7), .Y(_5277_) );
OAI21X1 OAI21X1_291 ( .A(_5275__bF_buf7), .B(_5276__bF_buf3), .C(_5277_), .Y(_1861_) );
NAND2X1 NAND2X1_331 ( .A(datapath_1_RegisterFile_dataWrite_1_), .B(_5272__bF_buf5), .Y(_5278_) );
NAND3X1 NAND3X1_167 ( .A(datapath_1_RegisterFile_regfile_mem_0__1_), .B(_5265__bF_buf45), .C(_5275__bF_buf2), .Y(_5279_) );
OAI21X1 OAI21X1_292 ( .A(_5275__bF_buf2), .B(_5278__bF_buf2), .C(_5279_), .Y(_1862_) );
NAND2X1 NAND2X1_332 ( .A(datapath_1_RegisterFile_dataWrite_2_), .B(_5272__bF_buf5), .Y(_5280_) );
NAND3X1 NAND3X1_168 ( .A(datapath_1_RegisterFile_regfile_mem_0__2_), .B(_5265__bF_buf56), .C(_5275__bF_buf6), .Y(_5281_) );
OAI21X1 OAI21X1_293 ( .A(_5275__bF_buf6), .B(_5280__bF_buf2), .C(_5281_), .Y(_1863_) );
NAND2X1 NAND2X1_333 ( .A(datapath_1_RegisterFile_dataWrite_3_), .B(_5272__bF_buf4), .Y(_5282_) );
NAND3X1 NAND3X1_169 ( .A(datapath_1_RegisterFile_regfile_mem_0__3_), .B(_5265__bF_buf44), .C(_5275__bF_buf1), .Y(_5283_) );
OAI21X1 OAI21X1_294 ( .A(_5275__bF_buf1), .B(_5282__bF_buf4), .C(_5283_), .Y(_1864_) );
NAND2X1 NAND2X1_334 ( .A(datapath_1_RegisterFile_dataWrite_4_), .B(_5272__bF_buf4), .Y(_5284_) );
NAND3X1 NAND3X1_170 ( .A(datapath_1_RegisterFile_regfile_mem_0__4_), .B(_5265__bF_buf13), .C(_5275__bF_buf4), .Y(_5285_) );
OAI21X1 OAI21X1_295 ( .A(_5275__bF_buf4), .B(_5284__bF_buf4), .C(_5285_), .Y(_1865_) );
NAND2X1 NAND2X1_335 ( .A(datapath_1_RegisterFile_dataWrite_5_), .B(_5272__bF_buf1), .Y(_5286_) );
NAND3X1 NAND3X1_171 ( .A(datapath_1_RegisterFile_regfile_mem_0__5_), .B(_5265__bF_buf48), .C(_5275__bF_buf7), .Y(_5287_) );
OAI21X1 OAI21X1_296 ( .A(_5275__bF_buf7), .B(_5286__bF_buf4), .C(_5287_), .Y(_1866_) );
NAND2X1 NAND2X1_336 ( .A(datapath_1_RegisterFile_dataWrite_6_), .B(_5272__bF_buf0), .Y(_5288_) );
NAND3X1 NAND3X1_172 ( .A(datapath_1_RegisterFile_regfile_mem_0__6_), .B(_5265__bF_buf5), .C(_5275__bF_buf2), .Y(_5289_) );
OAI21X1 OAI21X1_297 ( .A(_5275__bF_buf2), .B(_5288__bF_buf4), .C(_5289_), .Y(_1867_) );
NAND2X1 NAND2X1_337 ( .A(datapath_1_RegisterFile_dataWrite_7_), .B(_5272__bF_buf0), .Y(_5290_) );
NAND3X1 NAND3X1_173 ( .A(datapath_1_RegisterFile_regfile_mem_0__7_), .B(_5265__bF_buf86), .C(_5275__bF_buf5), .Y(_5291_) );
OAI21X1 OAI21X1_298 ( .A(_5275__bF_buf5), .B(_5290__bF_buf4), .C(_5291_), .Y(_1868_) );
NAND2X1 NAND2X1_338 ( .A(datapath_1_RegisterFile_dataWrite_8_), .B(_5272__bF_buf1), .Y(_5292_) );
NAND3X1 NAND3X1_174 ( .A(datapath_1_RegisterFile_regfile_mem_0__8_), .B(_5265__bF_buf97), .C(_5275__bF_buf0), .Y(_5293_) );
OAI21X1 OAI21X1_299 ( .A(_5275__bF_buf0), .B(_5292__bF_buf4), .C(_5293_), .Y(_1869_) );
NAND2X1 NAND2X1_339 ( .A(datapath_1_RegisterFile_dataWrite_9_), .B(_5272__bF_buf3), .Y(_5294_) );
NAND3X1 NAND3X1_175 ( .A(datapath_1_RegisterFile_regfile_mem_0__9_), .B(_5265__bF_buf60), .C(_5275__bF_buf3), .Y(_5295_) );
OAI21X1 OAI21X1_300 ( .A(_5275__bF_buf3), .B(_5294__bF_buf2), .C(_5295_), .Y(_1870_) );
NAND2X1 NAND2X1_340 ( .A(datapath_1_RegisterFile_dataWrite_10_), .B(_5272__bF_buf1), .Y(_5296_) );
NAND3X1 NAND3X1_176 ( .A(datapath_1_RegisterFile_regfile_mem_0__10_), .B(_5265__bF_buf56), .C(_5275__bF_buf6), .Y(_5297_) );
OAI21X1 OAI21X1_301 ( .A(_5275__bF_buf6), .B(_5296__bF_buf4), .C(_5297_), .Y(_1871_) );
NAND2X1 NAND2X1_341 ( .A(datapath_1_RegisterFile_dataWrite_11_), .B(_5272__bF_buf4), .Y(_5298_) );
NAND3X1 NAND3X1_177 ( .A(datapath_1_RegisterFile_regfile_mem_0__11_), .B(_5265__bF_buf44), .C(_5275__bF_buf1), .Y(_5299_) );
OAI21X1 OAI21X1_302 ( .A(_5275__bF_buf1), .B(_5298__bF_buf2), .C(_5299_), .Y(_1872_) );
NAND2X1 NAND2X1_342 ( .A(datapath_1_RegisterFile_dataWrite_12_), .B(_5272__bF_buf4), .Y(_5300_) );
NAND3X1 NAND3X1_178 ( .A(datapath_1_RegisterFile_regfile_mem_0__12_), .B(_5265__bF_buf45), .C(_5275__bF_buf2), .Y(_5301_) );
OAI21X1 OAI21X1_303 ( .A(_5275__bF_buf2), .B(_5300__bF_buf4), .C(_5301_), .Y(_1873_) );
NAND2X1 NAND2X1_343 ( .A(datapath_1_RegisterFile_dataWrite_13_), .B(_5272__bF_buf1), .Y(_5302_) );
NAND3X1 NAND3X1_179 ( .A(datapath_1_RegisterFile_regfile_mem_0__13_), .B(_5265__bF_buf18), .C(_5275__bF_buf3), .Y(_5303_) );
OAI21X1 OAI21X1_304 ( .A(_5275__bF_buf3), .B(_5302__bF_buf0), .C(_5303_), .Y(_1874_) );
NAND2X1 NAND2X1_344 ( .A(datapath_1_RegisterFile_dataWrite_14_), .B(_5272__bF_buf3), .Y(_5304_) );
NAND3X1 NAND3X1_180 ( .A(datapath_1_RegisterFile_regfile_mem_0__14_), .B(_5265__bF_buf77), .C(_5275__bF_buf4), .Y(_5305_) );
OAI21X1 OAI21X1_305 ( .A(_5275__bF_buf4), .B(_5304__bF_buf3), .C(_5305_), .Y(_1875_) );
NAND2X1 NAND2X1_345 ( .A(datapath_1_RegisterFile_dataWrite_15_), .B(_5272__bF_buf0), .Y(_5306_) );
NAND3X1 NAND3X1_181 ( .A(datapath_1_RegisterFile_regfile_mem_0__15_), .B(_5265__bF_buf86), .C(_5275__bF_buf5), .Y(_5307_) );
OAI21X1 OAI21X1_306 ( .A(_5275__bF_buf5), .B(_5306__bF_buf1), .C(_5307_), .Y(_1876_) );
NAND2X1 NAND2X1_346 ( .A(datapath_1_RegisterFile_dataWrite_16_), .B(_5272__bF_buf4), .Y(_5308_) );
NAND3X1 NAND3X1_182 ( .A(datapath_1_RegisterFile_regfile_mem_0__16_), .B(_5265__bF_buf91), .C(_5275__bF_buf6), .Y(_5309_) );
OAI21X1 OAI21X1_307 ( .A(_5275__bF_buf6), .B(_5308__bF_buf2), .C(_5309_), .Y(_1877_) );
NAND2X1 NAND2X1_347 ( .A(datapath_1_RegisterFile_dataWrite_17_), .B(_5272__bF_buf0), .Y(_5310_) );
NAND3X1 NAND3X1_183 ( .A(datapath_1_RegisterFile_regfile_mem_0__17_), .B(_5265__bF_buf28), .C(_5275__bF_buf0), .Y(_5311_) );
OAI21X1 OAI21X1_308 ( .A(_5275__bF_buf0), .B(_5310__bF_buf2), .C(_5311_), .Y(_1878_) );
NAND2X1 NAND2X1_348 ( .A(datapath_1_RegisterFile_dataWrite_18_), .B(_5272__bF_buf3), .Y(_5312_) );
NAND3X1 NAND3X1_184 ( .A(datapath_1_RegisterFile_regfile_mem_0__18_), .B(_5265__bF_buf18), .C(_5275__bF_buf3), .Y(_5313_) );
OAI21X1 OAI21X1_309 ( .A(_5275__bF_buf3), .B(_5312__bF_buf3), .C(_5313_), .Y(_1879_) );
NAND2X1 NAND2X1_349 ( .A(datapath_1_RegisterFile_dataWrite_19_), .B(_5272__bF_buf4), .Y(_5314_) );
NAND3X1 NAND3X1_185 ( .A(datapath_1_RegisterFile_regfile_mem_0__19_), .B(_5265__bF_buf94), .C(_5275__bF_buf1), .Y(_5315_) );
OAI21X1 OAI21X1_310 ( .A(_5275__bF_buf1), .B(_5314__bF_buf3), .C(_5315_), .Y(_1880_) );
NAND2X1 NAND2X1_350 ( .A(datapath_1_RegisterFile_dataWrite_20_), .B(_5272__bF_buf0), .Y(_5316_) );
NAND3X1 NAND3X1_186 ( .A(datapath_1_RegisterFile_regfile_mem_0__20_), .B(_5265__bF_buf44), .C(_5275__bF_buf1), .Y(_5317_) );
OAI21X1 OAI21X1_311 ( .A(_5275__bF_buf1), .B(_5316__bF_buf2), .C(_5317_), .Y(_1881_) );
NAND2X1 NAND2X1_351 ( .A(datapath_1_RegisterFile_dataWrite_21_), .B(_5272__bF_buf5), .Y(_5318_) );
NAND3X1 NAND3X1_187 ( .A(datapath_1_RegisterFile_regfile_mem_0__21_), .B(_5265__bF_buf65), .C(_5275__bF_buf0), .Y(_5319_) );
OAI21X1 OAI21X1_312 ( .A(_5275__bF_buf0), .B(_5318__bF_buf2), .C(_5319_), .Y(_859_) );
NAND2X1 NAND2X1_352 ( .A(datapath_1_RegisterFile_dataWrite_22_), .B(_5272__bF_buf1), .Y(_5320_) );
NAND3X1 NAND3X1_188 ( .A(datapath_1_RegisterFile_regfile_mem_0__22_), .B(_5265__bF_buf22), .C(_5275__bF_buf7), .Y(_5321_) );
OAI21X1 OAI21X1_313 ( .A(_5275__bF_buf7), .B(_5320__bF_buf3), .C(_5321_), .Y(_860_) );
NAND2X1 NAND2X1_353 ( .A(datapath_1_RegisterFile_dataWrite_23_), .B(_5272__bF_buf1), .Y(_5322_) );
NAND3X1 NAND3X1_189 ( .A(datapath_1_RegisterFile_regfile_mem_0__23_), .B(_5265__bF_buf27), .C(_5275__bF_buf4), .Y(_5323_) );
OAI21X1 OAI21X1_314 ( .A(_5275__bF_buf4), .B(_5322__bF_buf1), .C(_5323_), .Y(_861_) );
NAND2X1 NAND2X1_354 ( .A(datapath_1_RegisterFile_dataWrite_24_), .B(_5272__bF_buf5), .Y(_5324_) );
NAND3X1 NAND3X1_190 ( .A(datapath_1_RegisterFile_regfile_mem_0__24_), .B(_5265__bF_buf85), .C(_5275__bF_buf5), .Y(_5325_) );
OAI21X1 OAI21X1_315 ( .A(_5275__bF_buf5), .B(_5324__bF_buf3), .C(_5325_), .Y(_862_) );
NAND2X1 NAND2X1_355 ( .A(datapath_1_RegisterFile_dataWrite_25_), .B(_5272__bF_buf5), .Y(_5326_) );
NAND3X1 NAND3X1_191 ( .A(datapath_1_RegisterFile_regfile_mem_0__25_), .B(_5265__bF_buf25), .C(_5275__bF_buf2), .Y(_5327_) );
OAI21X1 OAI21X1_316 ( .A(_5275__bF_buf2), .B(_5326__bF_buf2), .C(_5327_), .Y(_863_) );
NAND2X1 NAND2X1_356 ( .A(datapath_1_RegisterFile_dataWrite_26_), .B(_5272__bF_buf3), .Y(_5328_) );
NAND3X1 NAND3X1_192 ( .A(datapath_1_RegisterFile_regfile_mem_0__26_), .B(_5265__bF_buf64), .C(_5275__bF_buf7), .Y(_5329_) );
OAI21X1 OAI21X1_317 ( .A(_5275__bF_buf7), .B(_5328__bF_buf0), .C(_5329_), .Y(_1882_) );
NAND2X1 NAND2X1_357 ( .A(datapath_1_RegisterFile_dataWrite_27_), .B(_5272__bF_buf3), .Y(_5330_) );
NAND3X1 NAND3X1_193 ( .A(datapath_1_RegisterFile_regfile_mem_0__27_), .B(_5265__bF_buf27), .C(_5275__bF_buf4), .Y(_5331_) );
OAI21X1 OAI21X1_318 ( .A(_5275__bF_buf4), .B(_5330__bF_buf4), .C(_5331_), .Y(_864_) );
NAND2X1 NAND2X1_358 ( .A(datapath_1_RegisterFile_dataWrite_28_), .B(_5272__bF_buf5), .Y(_5332_) );
NAND3X1 NAND3X1_194 ( .A(datapath_1_RegisterFile_regfile_mem_0__28_), .B(_5265__bF_buf84), .C(_5275__bF_buf5), .Y(_5333_) );
OAI21X1 OAI21X1_319 ( .A(_5275__bF_buf5), .B(_5332__bF_buf4), .C(_5333_), .Y(_865_) );
NAND2X1 NAND2X1_359 ( .A(datapath_1_RegisterFile_dataWrite_29_), .B(_5272__bF_buf4), .Y(_5334_) );
NAND3X1 NAND3X1_195 ( .A(datapath_1_RegisterFile_regfile_mem_0__29_), .B(_5265__bF_buf35), .C(_5275__bF_buf6), .Y(_5335_) );
OAI21X1 OAI21X1_320 ( .A(_5275__bF_buf6), .B(_5334__bF_buf4), .C(_5335_), .Y(_866_) );
NAND2X1 NAND2X1_360 ( .A(datapath_1_RegisterFile_dataWrite_30_), .B(_5272__bF_buf0), .Y(_5336_) );
NAND3X1 NAND3X1_196 ( .A(datapath_1_RegisterFile_regfile_mem_0__30_), .B(_5265__bF_buf28), .C(_5275__bF_buf0), .Y(_5337_) );
OAI21X1 OAI21X1_321 ( .A(_5275__bF_buf0), .B(_5336__bF_buf0), .C(_5337_), .Y(_867_) );
NAND2X1 NAND2X1_361 ( .A(datapath_1_RegisterFile_dataWrite_31_), .B(_5272__bF_buf3), .Y(_5338_) );
NAND3X1 NAND3X1_197 ( .A(datapath_1_RegisterFile_regfile_mem_0__31_), .B(_5265__bF_buf73), .C(_5275__bF_buf3), .Y(_5339_) );
OAI21X1 OAI21X1_322 ( .A(_5275__bF_buf3), .B(_5338__bF_buf4), .C(_5339_), .Y(_868_) );
NAND2X1 NAND2X1_362 ( .A(_5271_), .B(_5272__bF_buf2), .Y(_5340_) );
NOR2X1 NOR2X1_133 ( .A(_5270_), .B(_5340_), .Y(_5341_) );
NAND2X1 NAND2X1_363 ( .A(_5341_), .B(_5269_), .Y(_5342_) );
NAND3X1 NAND3X1_198 ( .A(datapath_1_RegisterFile_regfile_mem_1__0_), .B(_5265__bF_buf31), .C(_5342__bF_buf0), .Y(_5343_) );
OAI21X1 OAI21X1_323 ( .A(_5276__bF_buf3), .B(_5342__bF_buf0), .C(_5343_), .Y(_1128_) );
NAND3X1 NAND3X1_199 ( .A(datapath_1_RegisterFile_regfile_mem_1__1_), .B(_5265__bF_buf45), .C(_5342__bF_buf3), .Y(_5344_) );
OAI21X1 OAI21X1_324 ( .A(_5278__bF_buf2), .B(_5342__bF_buf3), .C(_5344_), .Y(_1618_) );
NAND3X1 NAND3X1_200 ( .A(datapath_1_RegisterFile_regfile_mem_1__2_), .B(_5265__bF_buf56), .C(_5342__bF_buf3), .Y(_5345_) );
OAI21X1 OAI21X1_325 ( .A(_5280__bF_buf1), .B(_5342__bF_buf3), .C(_5345_), .Y(_1141_) );
NAND3X1 NAND3X1_201 ( .A(datapath_1_RegisterFile_regfile_mem_1__3_), .B(_5265__bF_buf45), .C(_5342__bF_buf3), .Y(_5346_) );
OAI21X1 OAI21X1_326 ( .A(_5282__bF_buf4), .B(_5342__bF_buf3), .C(_5346_), .Y(_1143_) );
NAND3X1 NAND3X1_202 ( .A(datapath_1_RegisterFile_regfile_mem_1__4_), .B(_5265__bF_buf97), .C(_5342__bF_buf2), .Y(_5347_) );
OAI21X1 OAI21X1_327 ( .A(_5284__bF_buf1), .B(_5342__bF_buf2), .C(_5347_), .Y(_1144_) );
NAND3X1 NAND3X1_203 ( .A(datapath_1_RegisterFile_regfile_mem_1__5_), .B(_5265__bF_buf77), .C(_5342__bF_buf4), .Y(_5348_) );
OAI21X1 OAI21X1_328 ( .A(_5286__bF_buf1), .B(_5342__bF_buf4), .C(_5348_), .Y(_1145_) );
NAND3X1 NAND3X1_204 ( .A(datapath_1_RegisterFile_regfile_mem_1__6_), .B(_5265__bF_buf92), .C(_5342__bF_buf2), .Y(_5349_) );
OAI21X1 OAI21X1_329 ( .A(_5288__bF_buf3), .B(_5342__bF_buf2), .C(_5349_), .Y(_1619_) );
NAND3X1 NAND3X1_205 ( .A(datapath_1_RegisterFile_regfile_mem_1__7_), .B(_5265__bF_buf86), .C(_5342__bF_buf1), .Y(_5350_) );
OAI21X1 OAI21X1_330 ( .A(_5290__bF_buf4), .B(_5342__bF_buf1), .C(_5350_), .Y(_1146_) );
NAND3X1 NAND3X1_206 ( .A(datapath_1_RegisterFile_regfile_mem_1__8_), .B(_5265__bF_buf97), .C(_5342__bF_buf2), .Y(_5351_) );
OAI21X1 OAI21X1_331 ( .A(_5292__bF_buf1), .B(_5342__bF_buf2), .C(_5351_), .Y(_1147_) );
NAND3X1 NAND3X1_207 ( .A(datapath_1_RegisterFile_regfile_mem_1__9_), .B(_5265__bF_buf27), .C(_5342__bF_buf4), .Y(_5352_) );
OAI21X1 OAI21X1_332 ( .A(_5294__bF_buf3), .B(_5342__bF_buf4), .C(_5352_), .Y(_1148_) );
NAND3X1 NAND3X1_208 ( .A(datapath_1_RegisterFile_regfile_mem_1__10_), .B(_5265__bF_buf65), .C(_5342__bF_buf6), .Y(_5353_) );
OAI21X1 OAI21X1_333 ( .A(_5296__bF_buf2), .B(_5342__bF_buf6), .C(_5353_), .Y(_1129_) );
NAND3X1 NAND3X1_209 ( .A(datapath_1_RegisterFile_regfile_mem_1__11_), .B(_5265__bF_buf93), .C(_5342__bF_buf6), .Y(_5354_) );
OAI21X1 OAI21X1_334 ( .A(_5298__bF_buf2), .B(_5342__bF_buf6), .C(_5354_), .Y(_1620_) );
NAND3X1 NAND3X1_210 ( .A(datapath_1_RegisterFile_regfile_mem_1__12_), .B(_5265__bF_buf50), .C(_5342__bF_buf3), .Y(_5355_) );
OAI21X1 OAI21X1_335 ( .A(_5300__bF_buf1), .B(_5342__bF_buf3), .C(_5355_), .Y(_1130_) );
NAND3X1 NAND3X1_211 ( .A(datapath_1_RegisterFile_regfile_mem_1__13_), .B(_5265__bF_buf48), .C(_5342__bF_buf7), .Y(_5356_) );
OAI21X1 OAI21X1_336 ( .A(_5302__bF_buf2), .B(_5342__bF_buf7), .C(_5356_), .Y(_1131_) );
NAND3X1 NAND3X1_212 ( .A(datapath_1_RegisterFile_regfile_mem_1__14_), .B(_5265__bF_buf27), .C(_5342__bF_buf4), .Y(_5357_) );
OAI21X1 OAI21X1_337 ( .A(_5304__bF_buf3), .B(_5342__bF_buf4), .C(_5357_), .Y(_1132_) );
NAND3X1 NAND3X1_213 ( .A(datapath_1_RegisterFile_regfile_mem_1__15_), .B(_5265__bF_buf85), .C(_5342__bF_buf1), .Y(_5358_) );
OAI21X1 OAI21X1_338 ( .A(_5306__bF_buf1), .B(_5342__bF_buf1), .C(_5358_), .Y(_1133_) );
NAND3X1 NAND3X1_214 ( .A(datapath_1_RegisterFile_regfile_mem_1__16_), .B(_5265__bF_buf35), .C(_5342__bF_buf5), .Y(_5359_) );
OAI21X1 OAI21X1_339 ( .A(_5308__bF_buf2), .B(_5342__bF_buf5), .C(_5359_), .Y(_1621_) );
NAND3X1 NAND3X1_215 ( .A(datapath_1_RegisterFile_regfile_mem_1__17_), .B(_5265__bF_buf38), .C(_5342__bF_buf0), .Y(_5360_) );
OAI21X1 OAI21X1_340 ( .A(_5310__bF_buf2), .B(_5342__bF_buf0), .C(_5360_), .Y(_1134_) );
NAND3X1 NAND3X1_216 ( .A(datapath_1_RegisterFile_regfile_mem_1__18_), .B(_5265__bF_buf18), .C(_5342__bF_buf7), .Y(_5361_) );
OAI21X1 OAI21X1_341 ( .A(_5312__bF_buf3), .B(_5342__bF_buf7), .C(_5361_), .Y(_1622_) );
NAND3X1 NAND3X1_217 ( .A(datapath_1_RegisterFile_regfile_mem_1__19_), .B(_5265__bF_buf35), .C(_5342__bF_buf5), .Y(_5362_) );
OAI21X1 OAI21X1_342 ( .A(_5314__bF_buf3), .B(_5342__bF_buf5), .C(_5362_), .Y(_1623_) );
NAND3X1 NAND3X1_218 ( .A(datapath_1_RegisterFile_regfile_mem_1__20_), .B(_5265__bF_buf35), .C(_5342__bF_buf5), .Y(_5363_) );
OAI21X1 OAI21X1_343 ( .A(_5316__bF_buf2), .B(_5342__bF_buf5), .C(_5363_), .Y(_1624_) );
NAND3X1 NAND3X1_219 ( .A(datapath_1_RegisterFile_regfile_mem_1__21_), .B(_5265__bF_buf65), .C(_5342__bF_buf6), .Y(_5364_) );
OAI21X1 OAI21X1_344 ( .A(_5318__bF_buf4), .B(_5342__bF_buf6), .C(_5364_), .Y(_1625_) );
NAND3X1 NAND3X1_220 ( .A(datapath_1_RegisterFile_regfile_mem_1__22_), .B(_5265__bF_buf22), .C(_5342__bF_buf7), .Y(_5365_) );
OAI21X1 OAI21X1_345 ( .A(_5320__bF_buf3), .B(_5342__bF_buf7), .C(_5365_), .Y(_1626_) );
NAND3X1 NAND3X1_221 ( .A(datapath_1_RegisterFile_regfile_mem_1__23_), .B(_5265__bF_buf21), .C(_5342__bF_buf0), .Y(_5366_) );
OAI21X1 OAI21X1_346 ( .A(_5322__bF_buf2), .B(_5342__bF_buf0), .C(_5366_), .Y(_1135_) );
NAND3X1 NAND3X1_222 ( .A(datapath_1_RegisterFile_regfile_mem_1__24_), .B(_5265__bF_buf86), .C(_5342__bF_buf1), .Y(_5367_) );
OAI21X1 OAI21X1_347 ( .A(_5324__bF_buf3), .B(_5342__bF_buf1), .C(_5367_), .Y(_1136_) );
NAND3X1 NAND3X1_223 ( .A(datapath_1_RegisterFile_regfile_mem_1__25_), .B(_5265__bF_buf25), .C(_5342__bF_buf6), .Y(_5368_) );
OAI21X1 OAI21X1_348 ( .A(_5326__bF_buf2), .B(_5342__bF_buf6), .C(_5368_), .Y(_1137_) );
NAND3X1 NAND3X1_224 ( .A(datapath_1_RegisterFile_regfile_mem_1__26_), .B(_5265__bF_buf64), .C(_5342__bF_buf0), .Y(_5369_) );
OAI21X1 OAI21X1_349 ( .A(_5328__bF_buf0), .B(_5342__bF_buf0), .C(_5369_), .Y(_1627_) );
NAND3X1 NAND3X1_225 ( .A(datapath_1_RegisterFile_regfile_mem_1__27_), .B(_5265__bF_buf27), .C(_5342__bF_buf4), .Y(_5370_) );
OAI21X1 OAI21X1_350 ( .A(_5330__bF_buf4), .B(_5342__bF_buf4), .C(_5370_), .Y(_1138_) );
NAND3X1 NAND3X1_226 ( .A(datapath_1_RegisterFile_regfile_mem_1__28_), .B(_5265__bF_buf84), .C(_5342__bF_buf1), .Y(_5371_) );
OAI21X1 OAI21X1_351 ( .A(_5332__bF_buf4), .B(_5342__bF_buf1), .C(_5371_), .Y(_1139_) );
NAND3X1 NAND3X1_227 ( .A(datapath_1_RegisterFile_regfile_mem_1__29_), .B(_5265__bF_buf35), .C(_5342__bF_buf5), .Y(_5372_) );
OAI21X1 OAI21X1_352 ( .A(_5334__bF_buf4), .B(_5342__bF_buf5), .C(_5372_), .Y(_1140_) );
NAND3X1 NAND3X1_228 ( .A(datapath_1_RegisterFile_regfile_mem_1__30_), .B(_5265__bF_buf28), .C(_5342__bF_buf2), .Y(_5373_) );
OAI21X1 OAI21X1_353 ( .A(_5336__bF_buf0), .B(_5342__bF_buf2), .C(_5373_), .Y(_1142_) );
NAND3X1 NAND3X1_229 ( .A(datapath_1_RegisterFile_regfile_mem_1__31_), .B(_5265__bF_buf73), .C(_5342__bF_buf7), .Y(_5374_) );
OAI21X1 OAI21X1_354 ( .A(_5338__bF_buf4), .B(_5342__bF_buf7), .C(_5374_), .Y(_1628_) );
NAND2X1 NAND2X1_364 ( .A(_5270_), .B(_5272__bF_buf2), .Y(_5375_) );
NOR2X1 NOR2X1_134 ( .A(_5271_), .B(_5375_), .Y(_5376_) );
NAND2X1 NAND2X1_365 ( .A(_5376_), .B(_5269_), .Y(_5377_) );
NAND3X1 NAND3X1_230 ( .A(datapath_1_RegisterFile_regfile_mem_2__0_), .B(_5265__bF_buf64), .C(_5377__bF_buf7), .Y(_5378_) );
OAI21X1 OAI21X1_355 ( .A(_5276__bF_buf0), .B(_5377__bF_buf7), .C(_5378_), .Y(_1367_) );
NAND3X1 NAND3X1_231 ( .A(datapath_1_RegisterFile_regfile_mem_2__1_), .B(_5265__bF_buf65), .C(_5377__bF_buf5), .Y(_5379_) );
OAI21X1 OAI21X1_356 ( .A(_5278__bF_buf4), .B(_5377__bF_buf5), .C(_5379_), .Y(_1377_) );
NAND3X1 NAND3X1_232 ( .A(datapath_1_RegisterFile_regfile_mem_2__2_), .B(_5265__bF_buf91), .C(_5377__bF_buf0), .Y(_5380_) );
OAI21X1 OAI21X1_357 ( .A(_5280__bF_buf2), .B(_5377__bF_buf0), .C(_5380_), .Y(_1387_) );
NAND3X1 NAND3X1_233 ( .A(datapath_1_RegisterFile_regfile_mem_2__3_), .B(_5265__bF_buf93), .C(_5377__bF_buf4), .Y(_5381_) );
OAI21X1 OAI21X1_358 ( .A(_5282__bF_buf4), .B(_5377__bF_buf4), .C(_5381_), .Y(_1390_) );
NAND3X1 NAND3X1_234 ( .A(datapath_1_RegisterFile_regfile_mem_2__4_), .B(_5265__bF_buf97), .C(_5377__bF_buf5), .Y(_5382_) );
OAI21X1 OAI21X1_359 ( .A(_5284__bF_buf2), .B(_5377__bF_buf5), .C(_5382_), .Y(_1391_) );
NAND3X1 NAND3X1_235 ( .A(datapath_1_RegisterFile_regfile_mem_2__5_), .B(_5265__bF_buf60), .C(_5377__bF_buf3), .Y(_5383_) );
OAI21X1 OAI21X1_360 ( .A(_5286__bF_buf0), .B(_5377__bF_buf3), .C(_5383_), .Y(_1392_) );
NAND3X1 NAND3X1_236 ( .A(datapath_1_RegisterFile_regfile_mem_2__6_), .B(_5265__bF_buf23), .C(_5377__bF_buf2), .Y(_5384_) );
OAI21X1 OAI21X1_361 ( .A(_5288__bF_buf3), .B(_5377__bF_buf2), .C(_5384_), .Y(_1629_) );
NAND3X1 NAND3X1_237 ( .A(datapath_1_RegisterFile_regfile_mem_2__7_), .B(_5265__bF_buf86), .C(_5377__bF_buf6), .Y(_5385_) );
OAI21X1 OAI21X1_362 ( .A(_5290__bF_buf4), .B(_5377__bF_buf6), .C(_5385_), .Y(_1393_) );
NAND3X1 NAND3X1_238 ( .A(datapath_1_RegisterFile_regfile_mem_2__8_), .B(_5265__bF_buf5), .C(_5377__bF_buf1), .Y(_5386_) );
OAI21X1 OAI21X1_363 ( .A(_5292__bF_buf1), .B(_5377__bF_buf1), .C(_5386_), .Y(_1394_) );
NAND3X1 NAND3X1_239 ( .A(datapath_1_RegisterFile_regfile_mem_2__9_), .B(_5265__bF_buf6), .C(_5377__bF_buf2), .Y(_5387_) );
OAI21X1 OAI21X1_364 ( .A(_5294__bF_buf3), .B(_5377__bF_buf2), .C(_5387_), .Y(_1395_) );
NAND3X1 NAND3X1_240 ( .A(datapath_1_RegisterFile_regfile_mem_2__10_), .B(_5265__bF_buf55), .C(_5377__bF_buf4), .Y(_5388_) );
OAI21X1 OAI21X1_365 ( .A(_5296__bF_buf2), .B(_5377__bF_buf4), .C(_5388_), .Y(_1368_) );
NAND3X1 NAND3X1_241 ( .A(datapath_1_RegisterFile_regfile_mem_2__11_), .B(_5265__bF_buf63), .C(_5377__bF_buf4), .Y(_5389_) );
OAI21X1 OAI21X1_366 ( .A(_5298__bF_buf2), .B(_5377__bF_buf4), .C(_5389_), .Y(_1369_) );
NAND3X1 NAND3X1_242 ( .A(datapath_1_RegisterFile_regfile_mem_2__12_), .B(_5265__bF_buf50), .C(_5377__bF_buf1), .Y(_5390_) );
OAI21X1 OAI21X1_367 ( .A(_5300__bF_buf1), .B(_5377__bF_buf1), .C(_5390_), .Y(_1370_) );
NAND3X1 NAND3X1_243 ( .A(datapath_1_RegisterFile_regfile_mem_2__13_), .B(_5265__bF_buf18), .C(_5377__bF_buf3), .Y(_5391_) );
OAI21X1 OAI21X1_368 ( .A(_5302__bF_buf0), .B(_5377__bF_buf3), .C(_5391_), .Y(_1371_) );
NAND3X1 NAND3X1_244 ( .A(datapath_1_RegisterFile_regfile_mem_2__14_), .B(_5265__bF_buf6), .C(_5377__bF_buf2), .Y(_5392_) );
OAI21X1 OAI21X1_369 ( .A(_5304__bF_buf0), .B(_5377__bF_buf2), .C(_5392_), .Y(_1372_) );
NAND3X1 NAND3X1_245 ( .A(datapath_1_RegisterFile_regfile_mem_2__15_), .B(_5265__bF_buf70), .C(_5377__bF_buf6), .Y(_5393_) );
OAI21X1 OAI21X1_370 ( .A(_5306__bF_buf1), .B(_5377__bF_buf6), .C(_5393_), .Y(_1373_) );
NAND3X1 NAND3X1_246 ( .A(datapath_1_RegisterFile_regfile_mem_2__16_), .B(_5265__bF_buf91), .C(_5377__bF_buf0), .Y(_5394_) );
OAI21X1 OAI21X1_371 ( .A(_5308__bF_buf2), .B(_5377__bF_buf0), .C(_5394_), .Y(_1630_) );
NAND3X1 NAND3X1_247 ( .A(datapath_1_RegisterFile_regfile_mem_2__17_), .B(_5265__bF_buf38), .C(_5377__bF_buf5), .Y(_5395_) );
OAI21X1 OAI21X1_372 ( .A(_5310__bF_buf1), .B(_5377__bF_buf5), .C(_5395_), .Y(_1374_) );
NAND3X1 NAND3X1_248 ( .A(datapath_1_RegisterFile_regfile_mem_2__18_), .B(_5265__bF_buf48), .C(_5377__bF_buf7), .Y(_5396_) );
OAI21X1 OAI21X1_373 ( .A(_5312__bF_buf3), .B(_5377__bF_buf7), .C(_5396_), .Y(_1375_) );
NAND3X1 NAND3X1_249 ( .A(datapath_1_RegisterFile_regfile_mem_2__19_), .B(_5265__bF_buf96), .C(_5377__bF_buf0), .Y(_5397_) );
OAI21X1 OAI21X1_374 ( .A(_5314__bF_buf3), .B(_5377__bF_buf0), .C(_5397_), .Y(_1376_) );
NAND3X1 NAND3X1_250 ( .A(datapath_1_RegisterFile_regfile_mem_2__20_), .B(_5265__bF_buf96), .C(_5377__bF_buf0), .Y(_5398_) );
OAI21X1 OAI21X1_375 ( .A(_5316__bF_buf3), .B(_5377__bF_buf0), .C(_5398_), .Y(_1378_) );
NAND3X1 NAND3X1_251 ( .A(datapath_1_RegisterFile_regfile_mem_2__21_), .B(_5265__bF_buf5), .C(_5377__bF_buf1), .Y(_5399_) );
OAI21X1 OAI21X1_376 ( .A(_5318__bF_buf4), .B(_5377__bF_buf1), .C(_5399_), .Y(_1379_) );
NAND3X1 NAND3X1_252 ( .A(datapath_1_RegisterFile_regfile_mem_2__22_), .B(_5265__bF_buf73), .C(_5377__bF_buf3), .Y(_5400_) );
OAI21X1 OAI21X1_377 ( .A(_5320__bF_buf4), .B(_5377__bF_buf3), .C(_5400_), .Y(_1380_) );
NAND3X1 NAND3X1_253 ( .A(datapath_1_RegisterFile_regfile_mem_2__23_), .B(_5265__bF_buf21), .C(_5377__bF_buf3), .Y(_5401_) );
OAI21X1 OAI21X1_378 ( .A(_5322__bF_buf2), .B(_5377__bF_buf3), .C(_5401_), .Y(_1381_) );
NAND3X1 NAND3X1_254 ( .A(datapath_1_RegisterFile_regfile_mem_2__24_), .B(_5265__bF_buf96), .C(_5377__bF_buf6), .Y(_5402_) );
OAI21X1 OAI21X1_379 ( .A(_5324__bF_buf3), .B(_5377__bF_buf6), .C(_5402_), .Y(_1382_) );
NAND3X1 NAND3X1_255 ( .A(datapath_1_RegisterFile_regfile_mem_2__25_), .B(_5265__bF_buf45), .C(_5377__bF_buf1), .Y(_5403_) );
OAI21X1 OAI21X1_380 ( .A(_5326__bF_buf2), .B(_5377__bF_buf1), .C(_5403_), .Y(_1383_) );
NAND3X1 NAND3X1_256 ( .A(datapath_1_RegisterFile_regfile_mem_2__26_), .B(_5265__bF_buf64), .C(_5377__bF_buf7), .Y(_5404_) );
OAI21X1 OAI21X1_381 ( .A(_5328__bF_buf3), .B(_5377__bF_buf7), .C(_5404_), .Y(_1631_) );
NAND3X1 NAND3X1_257 ( .A(datapath_1_RegisterFile_regfile_mem_2__27_), .B(_5265__bF_buf42), .C(_5377__bF_buf2), .Y(_5405_) );
OAI21X1 OAI21X1_382 ( .A(_5330__bF_buf3), .B(_5377__bF_buf2), .C(_5405_), .Y(_1384_) );
NAND3X1 NAND3X1_258 ( .A(datapath_1_RegisterFile_regfile_mem_2__28_), .B(_5265__bF_buf94), .C(_5377__bF_buf6), .Y(_5406_) );
OAI21X1 OAI21X1_383 ( .A(_5332__bF_buf1), .B(_5377__bF_buf6), .C(_5406_), .Y(_1385_) );
NAND3X1 NAND3X1_259 ( .A(datapath_1_RegisterFile_regfile_mem_2__29_), .B(_5265__bF_buf93), .C(_5377__bF_buf4), .Y(_5407_) );
OAI21X1 OAI21X1_384 ( .A(_5334__bF_buf1), .B(_5377__bF_buf4), .C(_5407_), .Y(_1386_) );
NAND3X1 NAND3X1_260 ( .A(datapath_1_RegisterFile_regfile_mem_2__30_), .B(_5265__bF_buf28), .C(_5377__bF_buf5), .Y(_5408_) );
OAI21X1 OAI21X1_385 ( .A(_5336__bF_buf2), .B(_5377__bF_buf5), .C(_5408_), .Y(_1388_) );
NAND3X1 NAND3X1_261 ( .A(datapath_1_RegisterFile_regfile_mem_2__31_), .B(_5265__bF_buf22), .C(_5377__bF_buf7), .Y(_5409_) );
OAI21X1 OAI21X1_386 ( .A(_5338__bF_buf4), .B(_5377__bF_buf7), .C(_5409_), .Y(_1389_) );
OAI21X1 OAI21X1_387 ( .A(_5270_), .B(_5271_), .C(_5272__bF_buf2), .Y(_5410_) );
NAND2X1 NAND2X1_366 ( .A(_5410_), .B(_5269_), .Y(_5411_) );
NAND3X1 NAND3X1_262 ( .A(datapath_1_RegisterFile_regfile_mem_3__0_), .B(_5265__bF_buf12), .C(_5411__bF_buf2), .Y(_5412_) );
OAI21X1 OAI21X1_388 ( .A(_5276__bF_buf3), .B(_5411__bF_buf2), .C(_5412_), .Y(_1447_) );
NAND3X1 NAND3X1_263 ( .A(datapath_1_RegisterFile_regfile_mem_3__1_), .B(_5265__bF_buf50), .C(_5411__bF_buf3), .Y(_5413_) );
OAI21X1 OAI21X1_389 ( .A(_5278__bF_buf2), .B(_5411__bF_buf3), .C(_5413_), .Y(_1457_) );
NAND3X1 NAND3X1_264 ( .A(datapath_1_RegisterFile_regfile_mem_3__2_), .B(_5265__bF_buf56), .C(_5411__bF_buf0), .Y(_5414_) );
OAI21X1 OAI21X1_390 ( .A(_5280__bF_buf1), .B(_5411__bF_buf0), .C(_5414_), .Y(_1467_) );
NAND3X1 NAND3X1_265 ( .A(datapath_1_RegisterFile_regfile_mem_3__3_), .B(_5265__bF_buf93), .C(_5411__bF_buf5), .Y(_5415_) );
OAI21X1 OAI21X1_391 ( .A(_5282__bF_buf2), .B(_5411__bF_buf5), .C(_5415_), .Y(_1470_) );
NAND3X1 NAND3X1_266 ( .A(datapath_1_RegisterFile_regfile_mem_3__4_), .B(_5265__bF_buf5), .C(_5411__bF_buf3), .Y(_5416_) );
OAI21X1 OAI21X1_392 ( .A(_5284__bF_buf1), .B(_5411__bF_buf3), .C(_5416_), .Y(_1471_) );
NAND3X1 NAND3X1_267 ( .A(datapath_1_RegisterFile_regfile_mem_3__5_), .B(_5265__bF_buf60), .C(_5411__bF_buf4), .Y(_5417_) );
OAI21X1 OAI21X1_393 ( .A(_5286__bF_buf0), .B(_5411__bF_buf4), .C(_5417_), .Y(_1472_) );
NAND3X1 NAND3X1_268 ( .A(datapath_1_RegisterFile_regfile_mem_3__6_), .B(_5265__bF_buf5), .C(_5411__bF_buf3), .Y(_5418_) );
OAI21X1 OAI21X1_394 ( .A(_5288__bF_buf2), .B(_5411__bF_buf3), .C(_5418_), .Y(_1473_) );
NAND3X1 NAND3X1_269 ( .A(datapath_1_RegisterFile_regfile_mem_3__7_), .B(_5265__bF_buf85), .C(_5411__bF_buf6), .Y(_5419_) );
OAI21X1 OAI21X1_395 ( .A(_5290__bF_buf4), .B(_5411__bF_buf6), .C(_5419_), .Y(_1474_) );
NAND3X1 NAND3X1_270 ( .A(datapath_1_RegisterFile_regfile_mem_3__8_), .B(_5265__bF_buf65), .C(_5411__bF_buf1), .Y(_5420_) );
OAI21X1 OAI21X1_396 ( .A(_5292__bF_buf4), .B(_5411__bF_buf1), .C(_5420_), .Y(_1475_) );
NAND3X1 NAND3X1_271 ( .A(datapath_1_RegisterFile_regfile_mem_3__9_), .B(_5265__bF_buf38), .C(_5411__bF_buf2), .Y(_5421_) );
OAI21X1 OAI21X1_397 ( .A(_5294__bF_buf4), .B(_5411__bF_buf2), .C(_5421_), .Y(_1632_) );
NAND3X1 NAND3X1_272 ( .A(datapath_1_RegisterFile_regfile_mem_3__10_), .B(_5265__bF_buf65), .C(_5411__bF_buf1), .Y(_5422_) );
OAI21X1 OAI21X1_398 ( .A(_5296__bF_buf2), .B(_5411__bF_buf1), .C(_5422_), .Y(_1448_) );
NAND3X1 NAND3X1_273 ( .A(datapath_1_RegisterFile_regfile_mem_3__11_), .B(_5265__bF_buf63), .C(_5411__bF_buf5), .Y(_5423_) );
OAI21X1 OAI21X1_399 ( .A(_5298__bF_buf2), .B(_5411__bF_buf5), .C(_5423_), .Y(_1449_) );
NAND3X1 NAND3X1_274 ( .A(datapath_1_RegisterFile_regfile_mem_3__12_), .B(_5265__bF_buf56), .C(_5411__bF_buf3), .Y(_5424_) );
OAI21X1 OAI21X1_400 ( .A(_5300__bF_buf1), .B(_5411__bF_buf3), .C(_5424_), .Y(_1450_) );
NAND3X1 NAND3X1_275 ( .A(datapath_1_RegisterFile_regfile_mem_3__13_), .B(_5265__bF_buf18), .C(_5411__bF_buf4), .Y(_5425_) );
OAI21X1 OAI21X1_401 ( .A(_5302__bF_buf0), .B(_5411__bF_buf4), .C(_5425_), .Y(_1451_) );
NAND3X1 NAND3X1_276 ( .A(datapath_1_RegisterFile_regfile_mem_3__14_), .B(_5265__bF_buf77), .C(_5411__bF_buf7), .Y(_5426_) );
OAI21X1 OAI21X1_402 ( .A(_5304__bF_buf3), .B(_5411__bF_buf7), .C(_5426_), .Y(_1452_) );
NAND3X1 NAND3X1_277 ( .A(datapath_1_RegisterFile_regfile_mem_3__15_), .B(_5265__bF_buf85), .C(_5411__bF_buf6), .Y(_5427_) );
OAI21X1 OAI21X1_403 ( .A(_5306__bF_buf1), .B(_5411__bF_buf6), .C(_5427_), .Y(_1453_) );
NAND3X1 NAND3X1_278 ( .A(datapath_1_RegisterFile_regfile_mem_3__16_), .B(_5265__bF_buf35), .C(_5411__bF_buf0), .Y(_5428_) );
OAI21X1 OAI21X1_404 ( .A(_5308__bF_buf2), .B(_5411__bF_buf0), .C(_5428_), .Y(_1454_) );
NAND3X1 NAND3X1_279 ( .A(datapath_1_RegisterFile_regfile_mem_3__17_), .B(_5265__bF_buf12), .C(_5411__bF_buf2), .Y(_5429_) );
OAI21X1 OAI21X1_405 ( .A(_5310__bF_buf2), .B(_5411__bF_buf2), .C(_5429_), .Y(_1455_) );
NAND3X1 NAND3X1_280 ( .A(datapath_1_RegisterFile_regfile_mem_3__18_), .B(_5265__bF_buf52), .C(_5411__bF_buf4), .Y(_5430_) );
OAI21X1 OAI21X1_406 ( .A(_5312__bF_buf1), .B(_5411__bF_buf4), .C(_5430_), .Y(_1456_) );
NAND3X1 NAND3X1_281 ( .A(datapath_1_RegisterFile_regfile_mem_3__19_), .B(_5265__bF_buf35), .C(_5411__bF_buf0), .Y(_5431_) );
OAI21X1 OAI21X1_407 ( .A(_5314__bF_buf3), .B(_5411__bF_buf0), .C(_5431_), .Y(_1633_) );
NAND3X1 NAND3X1_282 ( .A(datapath_1_RegisterFile_regfile_mem_3__20_), .B(_5265__bF_buf96), .C(_5411__bF_buf0), .Y(_5432_) );
OAI21X1 OAI21X1_408 ( .A(_5316__bF_buf2), .B(_5411__bF_buf0), .C(_5432_), .Y(_1458_) );
NAND3X1 NAND3X1_283 ( .A(datapath_1_RegisterFile_regfile_mem_3__21_), .B(_5265__bF_buf65), .C(_5411__bF_buf1), .Y(_5433_) );
OAI21X1 OAI21X1_409 ( .A(_5318__bF_buf4), .B(_5411__bF_buf1), .C(_5433_), .Y(_1459_) );
NAND3X1 NAND3X1_284 ( .A(datapath_1_RegisterFile_regfile_mem_3__22_), .B(_5265__bF_buf31), .C(_5411__bF_buf2), .Y(_5434_) );
OAI21X1 OAI21X1_410 ( .A(_5320__bF_buf3), .B(_5411__bF_buf2), .C(_5434_), .Y(_1460_) );
NAND3X1 NAND3X1_285 ( .A(datapath_1_RegisterFile_regfile_mem_3__23_), .B(_5265__bF_buf68), .C(_5411__bF_buf7), .Y(_5435_) );
OAI21X1 OAI21X1_411 ( .A(_5322__bF_buf1), .B(_5411__bF_buf7), .C(_5435_), .Y(_1461_) );
NAND3X1 NAND3X1_286 ( .A(datapath_1_RegisterFile_regfile_mem_3__24_), .B(_5265__bF_buf85), .C(_5411__bF_buf6), .Y(_5436_) );
OAI21X1 OAI21X1_412 ( .A(_5324__bF_buf3), .B(_5411__bF_buf6), .C(_5436_), .Y(_1462_) );
NAND3X1 NAND3X1_287 ( .A(datapath_1_RegisterFile_regfile_mem_3__25_), .B(_5265__bF_buf63), .C(_5411__bF_buf5), .Y(_5437_) );
OAI21X1 OAI21X1_413 ( .A(_5326__bF_buf0), .B(_5411__bF_buf5), .C(_5437_), .Y(_1463_) );
NAND3X1 NAND3X1_288 ( .A(datapath_1_RegisterFile_regfile_mem_3__26_), .B(_5265__bF_buf64), .C(_5411__bF_buf4), .Y(_5438_) );
OAI21X1 OAI21X1_414 ( .A(_5328__bF_buf3), .B(_5411__bF_buf4), .C(_5438_), .Y(_1464_) );
NAND3X1 NAND3X1_289 ( .A(datapath_1_RegisterFile_regfile_mem_3__27_), .B(_5265__bF_buf77), .C(_5411__bF_buf7), .Y(_5439_) );
OAI21X1 OAI21X1_415 ( .A(_5330__bF_buf4), .B(_5411__bF_buf7), .C(_5439_), .Y(_1465_) );
NAND3X1 NAND3X1_290 ( .A(datapath_1_RegisterFile_regfile_mem_3__28_), .B(_5265__bF_buf84), .C(_5411__bF_buf6), .Y(_5440_) );
OAI21X1 OAI21X1_416 ( .A(_5332__bF_buf4), .B(_5411__bF_buf6), .C(_5440_), .Y(_1466_) );
NAND3X1 NAND3X1_291 ( .A(datapath_1_RegisterFile_regfile_mem_3__29_), .B(_5265__bF_buf63), .C(_5411__bF_buf5), .Y(_5441_) );
OAI21X1 OAI21X1_417 ( .A(_5334__bF_buf2), .B(_5411__bF_buf5), .C(_5441_), .Y(_1634_) );
NAND3X1 NAND3X1_292 ( .A(datapath_1_RegisterFile_regfile_mem_3__30_), .B(_5265__bF_buf97), .C(_5411__bF_buf1), .Y(_5442_) );
OAI21X1 OAI21X1_418 ( .A(_5336__bF_buf0), .B(_5411__bF_buf1), .C(_5442_), .Y(_1468_) );
NAND3X1 NAND3X1_293 ( .A(datapath_1_RegisterFile_regfile_mem_3__31_), .B(_5265__bF_buf77), .C(_5411__bF_buf7), .Y(_5443_) );
OAI21X1 OAI21X1_419 ( .A(_5338__bF_buf0), .B(_5411__bF_buf7), .C(_5443_), .Y(_1469_) );
INVX1 INVX1_107 ( .A(datapath_1_A3_2_), .Y(_5444_) );
NOR2X1 NOR2X1_135 ( .A(_5444_), .B(_5268_), .Y(_5445_) );
NAND2X1 NAND2X1_367 ( .A(_5274_), .B(_5445_), .Y(_5446_) );
NAND3X1 NAND3X1_294 ( .A(datapath_1_RegisterFile_regfile_mem_4__0_), .B(_5265__bF_buf38), .C(_5446__bF_buf4), .Y(_5447_) );
OAI21X1 OAI21X1_420 ( .A(_5276__bF_buf0), .B(_5446__bF_buf4), .C(_5447_), .Y(_1476_) );
NAND3X1 NAND3X1_295 ( .A(datapath_1_RegisterFile_regfile_mem_4__1_), .B(_5265__bF_buf25), .C(_5446__bF_buf5), .Y(_5448_) );
OAI21X1 OAI21X1_421 ( .A(_5278__bF_buf4), .B(_5446__bF_buf5), .C(_5448_), .Y(_1486_) );
NAND3X1 NAND3X1_296 ( .A(datapath_1_RegisterFile_regfile_mem_4__2_), .B(_5265__bF_buf93), .C(_5446__bF_buf3), .Y(_5449_) );
OAI21X1 OAI21X1_422 ( .A(_5280__bF_buf0), .B(_5446__bF_buf3), .C(_5449_), .Y(_1635_) );
NAND3X1 NAND3X1_297 ( .A(datapath_1_RegisterFile_regfile_mem_4__3_), .B(_5265__bF_buf44), .C(_5446__bF_buf0), .Y(_5450_) );
OAI21X1 OAI21X1_423 ( .A(_5282__bF_buf2), .B(_5446__bF_buf0), .C(_5450_), .Y(_1498_) );
NAND3X1 NAND3X1_298 ( .A(datapath_1_RegisterFile_regfile_mem_4__4_), .B(_5265__bF_buf97), .C(_5446__bF_buf5), .Y(_5451_) );
OAI21X1 OAI21X1_424 ( .A(_5284__bF_buf2), .B(_5446__bF_buf5), .C(_5451_), .Y(_1499_) );
NAND3X1 NAND3X1_299 ( .A(datapath_1_RegisterFile_regfile_mem_4__5_), .B(_5265__bF_buf18), .C(_5446__bF_buf2), .Y(_5452_) );
OAI21X1 OAI21X1_425 ( .A(_5286__bF_buf4), .B(_5446__bF_buf2), .C(_5452_), .Y(_1500_) );
NAND3X1 NAND3X1_300 ( .A(datapath_1_RegisterFile_regfile_mem_4__6_), .B(_5265__bF_buf5), .C(_5446__bF_buf6), .Y(_5453_) );
OAI21X1 OAI21X1_426 ( .A(_5288__bF_buf4), .B(_5446__bF_buf6), .C(_5453_), .Y(_1501_) );
NAND3X1 NAND3X1_301 ( .A(datapath_1_RegisterFile_regfile_mem_4__7_), .B(_5265__bF_buf62), .C(_5446__bF_buf7), .Y(_5454_) );
OAI21X1 OAI21X1_427 ( .A(_5290__bF_buf0), .B(_5446__bF_buf7), .C(_5454_), .Y(_1502_) );
NAND3X1 NAND3X1_302 ( .A(datapath_1_RegisterFile_regfile_mem_4__8_), .B(_5265__bF_buf5), .C(_5446__bF_buf6), .Y(_5455_) );
OAI21X1 OAI21X1_428 ( .A(_5292__bF_buf1), .B(_5446__bF_buf6), .C(_5455_), .Y(_1503_) );
NAND3X1 NAND3X1_303 ( .A(datapath_1_RegisterFile_regfile_mem_4__9_), .B(_5265__bF_buf48), .C(_5446__bF_buf2), .Y(_5456_) );
OAI21X1 OAI21X1_429 ( .A(_5294__bF_buf4), .B(_5446__bF_buf2), .C(_5456_), .Y(_1504_) );
NAND3X1 NAND3X1_304 ( .A(datapath_1_RegisterFile_regfile_mem_4__10_), .B(_5265__bF_buf25), .C(_5446__bF_buf5), .Y(_5457_) );
OAI21X1 OAI21X1_430 ( .A(_5296__bF_buf4), .B(_5446__bF_buf5), .C(_5457_), .Y(_1477_) );
NAND3X1 NAND3X1_305 ( .A(datapath_1_RegisterFile_regfile_mem_4__11_), .B(_5265__bF_buf63), .C(_5446__bF_buf3), .Y(_5458_) );
OAI21X1 OAI21X1_431 ( .A(_5298__bF_buf2), .B(_5446__bF_buf3), .C(_5458_), .Y(_1478_) );
NAND3X1 NAND3X1_306 ( .A(datapath_1_RegisterFile_regfile_mem_4__12_), .B(_5265__bF_buf50), .C(_5446__bF_buf6), .Y(_5459_) );
OAI21X1 OAI21X1_432 ( .A(_5300__bF_buf1), .B(_5446__bF_buf6), .C(_5459_), .Y(_1636_) );
NAND3X1 NAND3X1_307 ( .A(datapath_1_RegisterFile_regfile_mem_4__13_), .B(_5265__bF_buf18), .C(_5446__bF_buf2), .Y(_5460_) );
OAI21X1 OAI21X1_433 ( .A(_5302__bF_buf0), .B(_5446__bF_buf2), .C(_5460_), .Y(_1479_) );
NAND3X1 NAND3X1_308 ( .A(datapath_1_RegisterFile_regfile_mem_4__14_), .B(_5265__bF_buf23), .C(_5446__bF_buf6), .Y(_5461_) );
OAI21X1 OAI21X1_434 ( .A(_5304__bF_buf0), .B(_5446__bF_buf6), .C(_5461_), .Y(_1480_) );
NAND3X1 NAND3X1_309 ( .A(datapath_1_RegisterFile_regfile_mem_4__15_), .B(_5265__bF_buf70), .C(_5446__bF_buf7), .Y(_5462_) );
OAI21X1 OAI21X1_435 ( .A(_5306__bF_buf3), .B(_5446__bF_buf7), .C(_5462_), .Y(_1481_) );
NAND3X1 NAND3X1_310 ( .A(datapath_1_RegisterFile_regfile_mem_4__16_), .B(_5265__bF_buf44), .C(_5446__bF_buf0), .Y(_5463_) );
OAI21X1 OAI21X1_436 ( .A(_5308__bF_buf3), .B(_5446__bF_buf0), .C(_5463_), .Y(_1482_) );
NAND3X1 NAND3X1_311 ( .A(datapath_1_RegisterFile_regfile_mem_4__17_), .B(_5265__bF_buf38), .C(_5446__bF_buf4), .Y(_5464_) );
OAI21X1 OAI21X1_437 ( .A(_5310__bF_buf1), .B(_5446__bF_buf4), .C(_5464_), .Y(_1483_) );
NAND3X1 NAND3X1_312 ( .A(datapath_1_RegisterFile_regfile_mem_4__18_), .B(_5265__bF_buf52), .C(_5446__bF_buf1), .Y(_5465_) );
OAI21X1 OAI21X1_438 ( .A(_5312__bF_buf0), .B(_5446__bF_buf1), .C(_5465_), .Y(_1484_) );
NAND3X1 NAND3X1_313 ( .A(datapath_1_RegisterFile_regfile_mem_4__19_), .B(_5265__bF_buf39), .C(_5446__bF_buf0), .Y(_5466_) );
OAI21X1 OAI21X1_439 ( .A(_5314__bF_buf1), .B(_5446__bF_buf0), .C(_5466_), .Y(_1485_) );
NAND3X1 NAND3X1_314 ( .A(datapath_1_RegisterFile_regfile_mem_4__20_), .B(_5265__bF_buf39), .C(_5446__bF_buf0), .Y(_5467_) );
OAI21X1 OAI21X1_440 ( .A(_5316__bF_buf1), .B(_5446__bF_buf0), .C(_5467_), .Y(_1487_) );
NAND3X1 NAND3X1_315 ( .A(datapath_1_RegisterFile_regfile_mem_4__21_), .B(_5265__bF_buf65), .C(_5446__bF_buf5), .Y(_5468_) );
OAI21X1 OAI21X1_441 ( .A(_5318__bF_buf4), .B(_5446__bF_buf5), .C(_5468_), .Y(_1488_) );
NAND3X1 NAND3X1_316 ( .A(datapath_1_RegisterFile_regfile_mem_4__22_), .B(_5265__bF_buf18), .C(_5446__bF_buf2), .Y(_5469_) );
OAI21X1 OAI21X1_442 ( .A(_5320__bF_buf4), .B(_5446__bF_buf2), .C(_5469_), .Y(_1637_) );
NAND3X1 NAND3X1_317 ( .A(datapath_1_RegisterFile_regfile_mem_4__23_), .B(_5265__bF_buf7), .C(_5446__bF_buf1), .Y(_5470_) );
OAI21X1 OAI21X1_443 ( .A(_5322__bF_buf3), .B(_5446__bF_buf1), .C(_5470_), .Y(_1489_) );
NAND3X1 NAND3X1_318 ( .A(datapath_1_RegisterFile_regfile_mem_4__24_), .B(_5265__bF_buf62), .C(_5446__bF_buf7), .Y(_5471_) );
OAI21X1 OAI21X1_444 ( .A(_5324__bF_buf4), .B(_5446__bF_buf7), .C(_5471_), .Y(_1490_) );
NAND3X1 NAND3X1_319 ( .A(datapath_1_RegisterFile_regfile_mem_4__25_), .B(_5265__bF_buf93), .C(_5446__bF_buf3), .Y(_5472_) );
OAI21X1 OAI21X1_445 ( .A(_5326__bF_buf0), .B(_5446__bF_buf3), .C(_5472_), .Y(_1491_) );
NAND3X1 NAND3X1_320 ( .A(datapath_1_RegisterFile_regfile_mem_4__26_), .B(_5265__bF_buf38), .C(_5446__bF_buf4), .Y(_5473_) );
OAI21X1 OAI21X1_446 ( .A(_5328__bF_buf2), .B(_5446__bF_buf4), .C(_5473_), .Y(_1492_) );
NAND3X1 NAND3X1_321 ( .A(datapath_1_RegisterFile_regfile_mem_4__27_), .B(_5265__bF_buf52), .C(_5446__bF_buf1), .Y(_5474_) );
OAI21X1 OAI21X1_447 ( .A(_5330__bF_buf0), .B(_5446__bF_buf1), .C(_5474_), .Y(_1493_) );
NAND3X1 NAND3X1_322 ( .A(datapath_1_RegisterFile_regfile_mem_4__28_), .B(_5265__bF_buf62), .C(_5446__bF_buf7), .Y(_5475_) );
OAI21X1 OAI21X1_448 ( .A(_5332__bF_buf0), .B(_5446__bF_buf7), .C(_5475_), .Y(_1494_) );
NAND3X1 NAND3X1_323 ( .A(datapath_1_RegisterFile_regfile_mem_4__29_), .B(_5265__bF_buf89), .C(_5446__bF_buf3), .Y(_5476_) );
OAI21X1 OAI21X1_449 ( .A(_5334__bF_buf2), .B(_5446__bF_buf3), .C(_5476_), .Y(_1495_) );
NAND3X1 NAND3X1_324 ( .A(datapath_1_RegisterFile_regfile_mem_4__30_), .B(_5265__bF_buf38), .C(_5446__bF_buf4), .Y(_5477_) );
OAI21X1 OAI21X1_450 ( .A(_5336__bF_buf2), .B(_5446__bF_buf4), .C(_5477_), .Y(_1496_) );
NAND3X1 NAND3X1_325 ( .A(datapath_1_RegisterFile_regfile_mem_4__31_), .B(_5265__bF_buf77), .C(_5446__bF_buf1), .Y(_5478_) );
OAI21X1 OAI21X1_451 ( .A(_5338__bF_buf0), .B(_5446__bF_buf1), .C(_5478_), .Y(_1497_) );
NAND2X1 NAND2X1_368 ( .A(_5341_), .B(_5445_), .Y(_5479_) );
NAND3X1 NAND3X1_326 ( .A(datapath_1_RegisterFile_regfile_mem_5__0_), .B(_5265__bF_buf31), .C(_5479__bF_buf5), .Y(_5480_) );
OAI21X1 OAI21X1_452 ( .A(_5276__bF_buf3), .B(_5479__bF_buf5), .C(_5480_), .Y(_1505_) );
NAND3X1 NAND3X1_327 ( .A(datapath_1_RegisterFile_regfile_mem_5__1_), .B(_5265__bF_buf45), .C(_5479__bF_buf1), .Y(_5481_) );
OAI21X1 OAI21X1_453 ( .A(_5278__bF_buf2), .B(_5479__bF_buf1), .C(_5481_), .Y(_1515_) );
NAND3X1 NAND3X1_328 ( .A(datapath_1_RegisterFile_regfile_mem_5__2_), .B(_5265__bF_buf93), .C(_5479__bF_buf7), .Y(_5482_) );
OAI21X1 OAI21X1_454 ( .A(_5280__bF_buf0), .B(_5479__bF_buf7), .C(_5482_), .Y(_1525_) );
NAND3X1 NAND3X1_329 ( .A(datapath_1_RegisterFile_regfile_mem_5__3_), .B(_5265__bF_buf44), .C(_5479__bF_buf1), .Y(_5483_) );
OAI21X1 OAI21X1_455 ( .A(_5282__bF_buf4), .B(_5479__bF_buf1), .C(_5483_), .Y(_1528_) );
NAND3X1 NAND3X1_330 ( .A(datapath_1_RegisterFile_regfile_mem_5__4_), .B(_5265__bF_buf92), .C(_5479__bF_buf6), .Y(_5484_) );
OAI21X1 OAI21X1_456 ( .A(_5284__bF_buf4), .B(_5479__bF_buf6), .C(_5484_), .Y(_1529_) );
NAND3X1 NAND3X1_331 ( .A(datapath_1_RegisterFile_regfile_mem_5__5_), .B(_5265__bF_buf18), .C(_5479__bF_buf5), .Y(_5485_) );
OAI21X1 OAI21X1_457 ( .A(_5286__bF_buf4), .B(_5479__bF_buf5), .C(_5485_), .Y(_1638_) );
NAND3X1 NAND3X1_332 ( .A(datapath_1_RegisterFile_regfile_mem_5__6_), .B(_5265__bF_buf5), .C(_5479__bF_buf6), .Y(_5486_) );
OAI21X1 OAI21X1_458 ( .A(_5288__bF_buf3), .B(_5479__bF_buf6), .C(_5486_), .Y(_1530_) );
NAND3X1 NAND3X1_333 ( .A(datapath_1_RegisterFile_regfile_mem_5__7_), .B(_5265__bF_buf62), .C(_5479__bF_buf2), .Y(_5487_) );
OAI21X1 OAI21X1_459 ( .A(_5290__bF_buf1), .B(_5479__bF_buf2), .C(_5487_), .Y(_1531_) );
NAND3X1 NAND3X1_334 ( .A(datapath_1_RegisterFile_regfile_mem_5__8_), .B(_5265__bF_buf72), .C(_5479__bF_buf3), .Y(_5488_) );
OAI21X1 OAI21X1_460 ( .A(_5292__bF_buf1), .B(_5479__bF_buf3), .C(_5488_), .Y(_1532_) );
NAND3X1 NAND3X1_335 ( .A(datapath_1_RegisterFile_regfile_mem_5__9_), .B(_5265__bF_buf48), .C(_5479__bF_buf0), .Y(_5489_) );
OAI21X1 OAI21X1_461 ( .A(_5294__bF_buf2), .B(_5479__bF_buf0), .C(_5489_), .Y(_1533_) );
NAND3X1 NAND3X1_336 ( .A(datapath_1_RegisterFile_regfile_mem_5__10_), .B(_5265__bF_buf55), .C(_5479__bF_buf7), .Y(_5490_) );
OAI21X1 OAI21X1_462 ( .A(_5296__bF_buf2), .B(_5479__bF_buf7), .C(_5490_), .Y(_1506_) );
NAND3X1 NAND3X1_337 ( .A(datapath_1_RegisterFile_regfile_mem_5__11_), .B(_5265__bF_buf89), .C(_5479__bF_buf4), .Y(_5491_) );
OAI21X1 OAI21X1_463 ( .A(_5298__bF_buf2), .B(_5479__bF_buf4), .C(_5491_), .Y(_1507_) );
NAND3X1 NAND3X1_338 ( .A(datapath_1_RegisterFile_regfile_mem_5__12_), .B(_5265__bF_buf50), .C(_5479__bF_buf1), .Y(_5492_) );
OAI21X1 OAI21X1_464 ( .A(_5300__bF_buf1), .B(_5479__bF_buf1), .C(_5492_), .Y(_1508_) );
NAND3X1 NAND3X1_339 ( .A(datapath_1_RegisterFile_regfile_mem_5__13_), .B(_5265__bF_buf18), .C(_5479__bF_buf5), .Y(_5493_) );
OAI21X1 OAI21X1_465 ( .A(_5302__bF_buf0), .B(_5479__bF_buf5), .C(_5493_), .Y(_1509_) );
NAND3X1 NAND3X1_340 ( .A(datapath_1_RegisterFile_regfile_mem_5__14_), .B(_5265__bF_buf6), .C(_5479__bF_buf6), .Y(_5494_) );
OAI21X1 OAI21X1_466 ( .A(_5304__bF_buf1), .B(_5479__bF_buf6), .C(_5494_), .Y(_1510_) );
NAND3X1 NAND3X1_341 ( .A(datapath_1_RegisterFile_regfile_mem_5__15_), .B(_5265__bF_buf70), .C(_5479__bF_buf2), .Y(_5495_) );
OAI21X1 OAI21X1_467 ( .A(_5306__bF_buf3), .B(_5479__bF_buf2), .C(_5495_), .Y(_1639_) );
NAND3X1 NAND3X1_342 ( .A(datapath_1_RegisterFile_regfile_mem_5__16_), .B(_5265__bF_buf26), .C(_5479__bF_buf1), .Y(_5496_) );
OAI21X1 OAI21X1_468 ( .A(_5308__bF_buf2), .B(_5479__bF_buf1), .C(_5496_), .Y(_1511_) );
NAND3X1 NAND3X1_343 ( .A(datapath_1_RegisterFile_regfile_mem_5__17_), .B(_5265__bF_buf97), .C(_5479__bF_buf3), .Y(_5497_) );
OAI21X1 OAI21X1_469 ( .A(_5310__bF_buf1), .B(_5479__bF_buf3), .C(_5497_), .Y(_1512_) );
NAND3X1 NAND3X1_344 ( .A(datapath_1_RegisterFile_regfile_mem_5__18_), .B(_5265__bF_buf7), .C(_5479__bF_buf0), .Y(_5498_) );
OAI21X1 OAI21X1_470 ( .A(_5312__bF_buf1), .B(_5479__bF_buf0), .C(_5498_), .Y(_1513_) );
NAND3X1 NAND3X1_345 ( .A(datapath_1_RegisterFile_regfile_mem_5__19_), .B(_5265__bF_buf89), .C(_5479__bF_buf4), .Y(_5499_) );
OAI21X1 OAI21X1_471 ( .A(_5314__bF_buf2), .B(_5479__bF_buf4), .C(_5499_), .Y(_1514_) );
NAND3X1 NAND3X1_346 ( .A(datapath_1_RegisterFile_regfile_mem_5__20_), .B(_5265__bF_buf44), .C(_5479__bF_buf4), .Y(_5500_) );
OAI21X1 OAI21X1_472 ( .A(_5316__bF_buf1), .B(_5479__bF_buf4), .C(_5500_), .Y(_1516_) );
NAND3X1 NAND3X1_347 ( .A(datapath_1_RegisterFile_regfile_mem_5__21_), .B(_5265__bF_buf65), .C(_5479__bF_buf7), .Y(_5501_) );
OAI21X1 OAI21X1_473 ( .A(_5318__bF_buf2), .B(_5479__bF_buf7), .C(_5501_), .Y(_1517_) );
NAND3X1 NAND3X1_348 ( .A(datapath_1_RegisterFile_regfile_mem_5__22_), .B(_5265__bF_buf73), .C(_5479__bF_buf5), .Y(_5502_) );
OAI21X1 OAI21X1_474 ( .A(_5320__bF_buf4), .B(_5479__bF_buf5), .C(_5502_), .Y(_1518_) );
NAND3X1 NAND3X1_349 ( .A(datapath_1_RegisterFile_regfile_mem_5__23_), .B(_5265__bF_buf7), .C(_5479__bF_buf0), .Y(_5503_) );
OAI21X1 OAI21X1_475 ( .A(_5322__bF_buf3), .B(_5479__bF_buf0), .C(_5503_), .Y(_1519_) );
NAND3X1 NAND3X1_350 ( .A(datapath_1_RegisterFile_regfile_mem_5__24_), .B(_5265__bF_buf70), .C(_5479__bF_buf2), .Y(_5504_) );
OAI21X1 OAI21X1_476 ( .A(_5324__bF_buf0), .B(_5479__bF_buf2), .C(_5504_), .Y(_1520_) );
NAND3X1 NAND3X1_351 ( .A(datapath_1_RegisterFile_regfile_mem_5__25_), .B(_5265__bF_buf55), .C(_5479__bF_buf7), .Y(_5505_) );
OAI21X1 OAI21X1_477 ( .A(_5326__bF_buf0), .B(_5479__bF_buf7), .C(_5505_), .Y(_1640_) );
NAND3X1 NAND3X1_352 ( .A(datapath_1_RegisterFile_regfile_mem_5__26_), .B(_5265__bF_buf38), .C(_5479__bF_buf3), .Y(_5506_) );
OAI21X1 OAI21X1_478 ( .A(_5328__bF_buf0), .B(_5479__bF_buf3), .C(_5506_), .Y(_1521_) );
NAND3X1 NAND3X1_353 ( .A(datapath_1_RegisterFile_regfile_mem_5__27_), .B(_5265__bF_buf68), .C(_5479__bF_buf6), .Y(_5507_) );
OAI21X1 OAI21X1_479 ( .A(_5330__bF_buf4), .B(_5479__bF_buf6), .C(_5507_), .Y(_1522_) );
NAND3X1 NAND3X1_354 ( .A(datapath_1_RegisterFile_regfile_mem_5__28_), .B(_5265__bF_buf62), .C(_5479__bF_buf2), .Y(_5508_) );
OAI21X1 OAI21X1_480 ( .A(_5332__bF_buf0), .B(_5479__bF_buf2), .C(_5508_), .Y(_1523_) );
NAND3X1 NAND3X1_355 ( .A(datapath_1_RegisterFile_regfile_mem_5__29_), .B(_5265__bF_buf44), .C(_5479__bF_buf4), .Y(_5509_) );
OAI21X1 OAI21X1_481 ( .A(_5334__bF_buf1), .B(_5479__bF_buf4), .C(_5509_), .Y(_1524_) );
NAND3X1 NAND3X1_356 ( .A(datapath_1_RegisterFile_regfile_mem_5__30_), .B(_5265__bF_buf28), .C(_5479__bF_buf3), .Y(_5510_) );
OAI21X1 OAI21X1_482 ( .A(_5336__bF_buf2), .B(_5479__bF_buf3), .C(_5510_), .Y(_1526_) );
NAND3X1 NAND3X1_357 ( .A(datapath_1_RegisterFile_regfile_mem_5__31_), .B(_5265__bF_buf7), .C(_5479__bF_buf0), .Y(_5511_) );
OAI21X1 OAI21X1_483 ( .A(_5338__bF_buf0), .B(_5479__bF_buf0), .C(_5511_), .Y(_1527_) );
NAND2X1 NAND2X1_369 ( .A(_5376_), .B(_5445_), .Y(_5512_) );
NAND3X1 NAND3X1_358 ( .A(datapath_1_RegisterFile_regfile_mem_6__0_), .B(_5265__bF_buf38), .C(_5512__bF_buf1), .Y(_5513_) );
OAI21X1 OAI21X1_484 ( .A(_5276__bF_buf0), .B(_5512__bF_buf1), .C(_5513_), .Y(_1534_) );
NAND3X1 NAND3X1_359 ( .A(datapath_1_RegisterFile_regfile_mem_6__1_), .B(_5265__bF_buf25), .C(_5512__bF_buf7), .Y(_5514_) );
OAI21X1 OAI21X1_485 ( .A(_5278__bF_buf4), .B(_5512__bF_buf7), .C(_5514_), .Y(_1544_) );
NAND3X1 NAND3X1_360 ( .A(datapath_1_RegisterFile_regfile_mem_6__2_), .B(_5265__bF_buf45), .C(_5512__bF_buf2), .Y(_5515_) );
OAI21X1 OAI21X1_486 ( .A(_5280__bF_buf0), .B(_5512__bF_buf2), .C(_5515_), .Y(_1554_) );
NAND3X1 NAND3X1_361 ( .A(datapath_1_RegisterFile_regfile_mem_6__3_), .B(_5265__bF_buf93), .C(_5512__bF_buf2), .Y(_5516_) );
OAI21X1 OAI21X1_487 ( .A(_5282__bF_buf4), .B(_5512__bF_buf2), .C(_5516_), .Y(_1557_) );
NAND3X1 NAND3X1_362 ( .A(datapath_1_RegisterFile_regfile_mem_6__4_), .B(_5265__bF_buf97), .C(_5512__bF_buf3), .Y(_5517_) );
OAI21X1 OAI21X1_488 ( .A(_5284__bF_buf1), .B(_5512__bF_buf3), .C(_5517_), .Y(_1558_) );
NAND3X1 NAND3X1_363 ( .A(datapath_1_RegisterFile_regfile_mem_6__5_), .B(_5265__bF_buf48), .C(_5512__bF_buf4), .Y(_5518_) );
OAI21X1 OAI21X1_489 ( .A(_5286__bF_buf4), .B(_5512__bF_buf4), .C(_5518_), .Y(_1559_) );
NAND3X1 NAND3X1_364 ( .A(datapath_1_RegisterFile_regfile_mem_6__6_), .B(_5265__bF_buf5), .C(_5512__bF_buf3), .Y(_5519_) );
OAI21X1 OAI21X1_490 ( .A(_5288__bF_buf4), .B(_5512__bF_buf3), .C(_5519_), .Y(_1560_) );
NAND3X1 NAND3X1_365 ( .A(datapath_1_RegisterFile_regfile_mem_6__7_), .B(_5265__bF_buf62), .C(_5512__bF_buf6), .Y(_5520_) );
OAI21X1 OAI21X1_491 ( .A(_5290__bF_buf0), .B(_5512__bF_buf6), .C(_5520_), .Y(_1561_) );
NAND3X1 NAND3X1_366 ( .A(datapath_1_RegisterFile_regfile_mem_6__8_), .B(_5265__bF_buf25), .C(_5512__bF_buf7), .Y(_5521_) );
OAI21X1 OAI21X1_492 ( .A(_5292__bF_buf4), .B(_5512__bF_buf7), .C(_5521_), .Y(_1641_) );
NAND3X1 NAND3X1_367 ( .A(datapath_1_RegisterFile_regfile_mem_6__9_), .B(_5265__bF_buf64), .C(_5512__bF_buf4), .Y(_5522_) );
OAI21X1 OAI21X1_493 ( .A(_5294__bF_buf4), .B(_5512__bF_buf4), .C(_5522_), .Y(_1562_) );
NAND3X1 NAND3X1_368 ( .A(datapath_1_RegisterFile_regfile_mem_6__10_), .B(_5265__bF_buf25), .C(_5512__bF_buf7), .Y(_5523_) );
OAI21X1 OAI21X1_494 ( .A(_5296__bF_buf2), .B(_5512__bF_buf7), .C(_5523_), .Y(_1535_) );
NAND3X1 NAND3X1_369 ( .A(datapath_1_RegisterFile_regfile_mem_6__11_), .B(_5265__bF_buf89), .C(_5512__bF_buf5), .Y(_5524_) );
OAI21X1 OAI21X1_495 ( .A(_5298__bF_buf0), .B(_5512__bF_buf5), .C(_5524_), .Y(_1536_) );
NAND3X1 NAND3X1_370 ( .A(datapath_1_RegisterFile_regfile_mem_6__12_), .B(_5265__bF_buf45), .C(_5512__bF_buf2), .Y(_5525_) );
OAI21X1 OAI21X1_496 ( .A(_5300__bF_buf4), .B(_5512__bF_buf2), .C(_5525_), .Y(_1537_) );
NAND3X1 NAND3X1_371 ( .A(datapath_1_RegisterFile_regfile_mem_6__13_), .B(_5265__bF_buf77), .C(_5512__bF_buf0), .Y(_5526_) );
OAI21X1 OAI21X1_497 ( .A(_5302__bF_buf4), .B(_5512__bF_buf0), .C(_5526_), .Y(_1538_) );
NAND3X1 NAND3X1_372 ( .A(datapath_1_RegisterFile_regfile_mem_6__14_), .B(_5265__bF_buf23), .C(_5512__bF_buf3), .Y(_5527_) );
OAI21X1 OAI21X1_498 ( .A(_5304__bF_buf0), .B(_5512__bF_buf3), .C(_5527_), .Y(_1539_) );
NAND3X1 NAND3X1_373 ( .A(datapath_1_RegisterFile_regfile_mem_6__15_), .B(_5265__bF_buf30), .C(_5512__bF_buf6), .Y(_5528_) );
OAI21X1 OAI21X1_499 ( .A(_5306__bF_buf4), .B(_5512__bF_buf6), .C(_5528_), .Y(_1540_) );
NAND3X1 NAND3X1_374 ( .A(datapath_1_RegisterFile_regfile_mem_6__16_), .B(_5265__bF_buf89), .C(_5512__bF_buf5), .Y(_5529_) );
OAI21X1 OAI21X1_500 ( .A(_5308__bF_buf3), .B(_5512__bF_buf5), .C(_5529_), .Y(_1541_) );
NAND3X1 NAND3X1_375 ( .A(datapath_1_RegisterFile_regfile_mem_6__17_), .B(_5265__bF_buf38), .C(_5512__bF_buf1), .Y(_5530_) );
OAI21X1 OAI21X1_501 ( .A(_5310__bF_buf1), .B(_5512__bF_buf1), .C(_5530_), .Y(_1542_) );
NAND3X1 NAND3X1_376 ( .A(datapath_1_RegisterFile_regfile_mem_6__18_), .B(_5265__bF_buf52), .C(_5512__bF_buf0), .Y(_5531_) );
OAI21X1 OAI21X1_502 ( .A(_5312__bF_buf0), .B(_5512__bF_buf0), .C(_5531_), .Y(_1642_) );
NAND3X1 NAND3X1_377 ( .A(datapath_1_RegisterFile_regfile_mem_6__19_), .B(_5265__bF_buf89), .C(_5512__bF_buf5), .Y(_5532_) );
OAI21X1 OAI21X1_503 ( .A(_5314__bF_buf2), .B(_5512__bF_buf5), .C(_5532_), .Y(_1543_) );
NAND3X1 NAND3X1_378 ( .A(datapath_1_RegisterFile_regfile_mem_6__20_), .B(_5265__bF_buf45), .C(_5512__bF_buf2), .Y(_5533_) );
OAI21X1 OAI21X1_504 ( .A(_5316__bF_buf2), .B(_5512__bF_buf2), .C(_5533_), .Y(_1545_) );
NAND3X1 NAND3X1_379 ( .A(datapath_1_RegisterFile_regfile_mem_6__21_), .B(_5265__bF_buf72), .C(_5512__bF_buf3), .Y(_5534_) );
OAI21X1 OAI21X1_505 ( .A(_5318__bF_buf4), .B(_5512__bF_buf3), .C(_5534_), .Y(_1546_) );
NAND3X1 NAND3X1_380 ( .A(datapath_1_RegisterFile_regfile_mem_6__22_), .B(_5265__bF_buf73), .C(_5512__bF_buf4), .Y(_5535_) );
OAI21X1 OAI21X1_506 ( .A(_5320__bF_buf4), .B(_5512__bF_buf4), .C(_5535_), .Y(_1547_) );
NAND3X1 NAND3X1_381 ( .A(datapath_1_RegisterFile_regfile_mem_6__23_), .B(_5265__bF_buf7), .C(_5512__bF_buf0), .Y(_5536_) );
OAI21X1 OAI21X1_507 ( .A(_5322__bF_buf3), .B(_5512__bF_buf0), .C(_5536_), .Y(_1548_) );
NAND3X1 NAND3X1_382 ( .A(datapath_1_RegisterFile_regfile_mem_6__24_), .B(_5265__bF_buf39), .C(_5512__bF_buf6), .Y(_5537_) );
OAI21X1 OAI21X1_508 ( .A(_5324__bF_buf4), .B(_5512__bF_buf6), .C(_5537_), .Y(_1549_) );
NAND3X1 NAND3X1_383 ( .A(datapath_1_RegisterFile_regfile_mem_6__25_), .B(_5265__bF_buf25), .C(_5512__bF_buf7), .Y(_5538_) );
OAI21X1 OAI21X1_509 ( .A(_5326__bF_buf2), .B(_5512__bF_buf7), .C(_5538_), .Y(_1550_) );
NAND3X1 NAND3X1_384 ( .A(datapath_1_RegisterFile_regfile_mem_6__26_), .B(_5265__bF_buf64), .C(_5512__bF_buf1), .Y(_5539_) );
OAI21X1 OAI21X1_510 ( .A(_5328__bF_buf2), .B(_5512__bF_buf1), .C(_5539_), .Y(_1551_) );
NAND3X1 NAND3X1_385 ( .A(datapath_1_RegisterFile_regfile_mem_6__27_), .B(_5265__bF_buf98), .C(_5512__bF_buf0), .Y(_5540_) );
OAI21X1 OAI21X1_511 ( .A(_5330__bF_buf0), .B(_5512__bF_buf0), .C(_5540_), .Y(_1552_) );
NAND3X1 NAND3X1_386 ( .A(datapath_1_RegisterFile_regfile_mem_6__28_), .B(_5265__bF_buf62), .C(_5512__bF_buf6), .Y(_5541_) );
OAI21X1 OAI21X1_512 ( .A(_5332__bF_buf1), .B(_5512__bF_buf6), .C(_5541_), .Y(_1643_) );
NAND3X1 NAND3X1_387 ( .A(datapath_1_RegisterFile_regfile_mem_6__29_), .B(_5265__bF_buf89), .C(_5512__bF_buf5), .Y(_5542_) );
OAI21X1 OAI21X1_513 ( .A(_5334__bF_buf2), .B(_5512__bF_buf5), .C(_5542_), .Y(_1553_) );
NAND3X1 NAND3X1_388 ( .A(datapath_1_RegisterFile_regfile_mem_6__30_), .B(_5265__bF_buf72), .C(_5512__bF_buf1), .Y(_5543_) );
OAI21X1 OAI21X1_514 ( .A(_5336__bF_buf2), .B(_5512__bF_buf1), .C(_5543_), .Y(_1555_) );
NAND3X1 NAND3X1_389 ( .A(datapath_1_RegisterFile_regfile_mem_6__31_), .B(_5265__bF_buf64), .C(_5512__bF_buf4), .Y(_5544_) );
OAI21X1 OAI21X1_515 ( .A(_5338__bF_buf3), .B(_5512__bF_buf4), .C(_5544_), .Y(_1556_) );
NAND2X1 NAND2X1_370 ( .A(_5410_), .B(_5445_), .Y(_5545_) );
NAND3X1 NAND3X1_390 ( .A(datapath_1_RegisterFile_regfile_mem_7__0_), .B(_5265__bF_buf87), .C(_5545__bF_buf0), .Y(_5546_) );
OAI21X1 OAI21X1_516 ( .A(_5276__bF_buf2), .B(_5545__bF_buf0), .C(_5546_), .Y(_1563_) );
NAND3X1 NAND3X1_391 ( .A(datapath_1_RegisterFile_regfile_mem_7__1_), .B(_5265__bF_buf25), .C(_5545__bF_buf2), .Y(_5547_) );
OAI21X1 OAI21X1_517 ( .A(_5278__bF_buf4), .B(_5545__bF_buf2), .C(_5547_), .Y(_1644_) );
NAND3X1 NAND3X1_392 ( .A(datapath_1_RegisterFile_regfile_mem_7__2_), .B(_5265__bF_buf25), .C(_5545__bF_buf3), .Y(_5548_) );
OAI21X1 OAI21X1_518 ( .A(_5280__bF_buf0), .B(_5545__bF_buf3), .C(_5548_), .Y(_1567_) );
NAND3X1 NAND3X1_393 ( .A(datapath_1_RegisterFile_regfile_mem_7__3_), .B(_5265__bF_buf93), .C(_5545__bF_buf3), .Y(_5549_) );
OAI21X1 OAI21X1_519 ( .A(_5282__bF_buf2), .B(_5545__bF_buf3), .C(_5549_), .Y(_1568_) );
NAND3X1 NAND3X1_394 ( .A(datapath_1_RegisterFile_regfile_mem_7__4_), .B(_5265__bF_buf97), .C(_5545__bF_buf5), .Y(_5550_) );
OAI21X1 OAI21X1_520 ( .A(_5284__bF_buf2), .B(_5545__bF_buf5), .C(_5550_), .Y(_1569_) );
NAND3X1 NAND3X1_395 ( .A(datapath_1_RegisterFile_regfile_mem_7__5_), .B(_5265__bF_buf52), .C(_5545__bF_buf6), .Y(_5551_) );
OAI21X1 OAI21X1_521 ( .A(_5286__bF_buf1), .B(_5545__bF_buf6), .C(_5551_), .Y(_1570_) );
NAND3X1 NAND3X1_396 ( .A(datapath_1_RegisterFile_regfile_mem_7__6_), .B(_5265__bF_buf23), .C(_5545__bF_buf0), .Y(_5552_) );
OAI21X1 OAI21X1_522 ( .A(_5288__bF_buf3), .B(_5545__bF_buf0), .C(_5552_), .Y(_1571_) );
NAND3X1 NAND3X1_397 ( .A(datapath_1_RegisterFile_regfile_mem_7__7_), .B(_5265__bF_buf62), .C(_5545__bF_buf4), .Y(_5553_) );
OAI21X1 OAI21X1_523 ( .A(_5290__bF_buf0), .B(_5545__bF_buf4), .C(_5553_), .Y(_1572_) );
NAND3X1 NAND3X1_398 ( .A(datapath_1_RegisterFile_regfile_mem_7__8_), .B(_5265__bF_buf5), .C(_5545__bF_buf5), .Y(_5554_) );
OAI21X1 OAI21X1_524 ( .A(_5292__bF_buf1), .B(_5545__bF_buf5), .C(_5554_), .Y(_1573_) );
NAND3X1 NAND3X1_399 ( .A(datapath_1_RegisterFile_regfile_mem_7__9_), .B(_5265__bF_buf6), .C(_5545__bF_buf0), .Y(_5555_) );
OAI21X1 OAI21X1_525 ( .A(_5294__bF_buf3), .B(_5545__bF_buf0), .C(_5555_), .Y(_1574_) );
NAND3X1 NAND3X1_400 ( .A(datapath_1_RegisterFile_regfile_mem_7__10_), .B(_5265__bF_buf55), .C(_5545__bF_buf2), .Y(_5556_) );
OAI21X1 OAI21X1_526 ( .A(_5296__bF_buf2), .B(_5545__bF_buf2), .C(_5556_), .Y(_1564_) );
NAND3X1 NAND3X1_401 ( .A(datapath_1_RegisterFile_regfile_mem_7__11_), .B(_5265__bF_buf36), .C(_5545__bF_buf1), .Y(_5557_) );
OAI21X1 OAI21X1_527 ( .A(_5298__bF_buf0), .B(_5545__bF_buf1), .C(_5557_), .Y(_1645_) );
NAND3X1 NAND3X1_402 ( .A(datapath_1_RegisterFile_regfile_mem_7__12_), .B(_5265__bF_buf45), .C(_5545__bF_buf3), .Y(_5558_) );
OAI21X1 OAI21X1_528 ( .A(_5300__bF_buf4), .B(_5545__bF_buf3), .C(_5558_), .Y(_1565_) );
NAND3X1 NAND3X1_403 ( .A(datapath_1_RegisterFile_regfile_mem_7__13_), .B(_5265__bF_buf73), .C(_5545__bF_buf7), .Y(_5559_) );
OAI21X1 OAI21X1_529 ( .A(_5302__bF_buf0), .B(_5545__bF_buf7), .C(_5559_), .Y(_1566_) );
NAND3X1 NAND3X1_404 ( .A(datapath_1_RegisterFile_regfile_mem_7__14_), .B(_5265__bF_buf6), .C(_5545__bF_buf0), .Y(_5560_) );
OAI21X1 OAI21X1_530 ( .A(_5304__bF_buf0), .B(_5545__bF_buf0), .C(_5560_), .Y(_1646_) );
NAND3X1 NAND3X1_405 ( .A(datapath_1_RegisterFile_regfile_mem_7__15_), .B(_5265__bF_buf39), .C(_5545__bF_buf1), .Y(_5561_) );
OAI21X1 OAI21X1_531 ( .A(_5306__bF_buf4), .B(_5545__bF_buf1), .C(_5561_), .Y(_1647_) );
NAND3X1 NAND3X1_406 ( .A(datapath_1_RegisterFile_regfile_mem_7__16_), .B(_5265__bF_buf62), .C(_5545__bF_buf4), .Y(_5562_) );
OAI21X1 OAI21X1_532 ( .A(_5308__bF_buf3), .B(_5545__bF_buf4), .C(_5562_), .Y(_1648_) );
NAND3X1 NAND3X1_407 ( .A(datapath_1_RegisterFile_regfile_mem_7__17_), .B(_5265__bF_buf97), .C(_5545__bF_buf5), .Y(_5563_) );
OAI21X1 OAI21X1_533 ( .A(_5310__bF_buf1), .B(_5545__bF_buf5), .C(_5563_), .Y(_1649_) );
NAND3X1 NAND3X1_408 ( .A(datapath_1_RegisterFile_regfile_mem_7__18_), .B(_5265__bF_buf60), .C(_5545__bF_buf7), .Y(_5564_) );
OAI21X1 OAI21X1_534 ( .A(_5312__bF_buf3), .B(_5545__bF_buf7), .C(_5564_), .Y(_1650_) );
NAND3X1 NAND3X1_409 ( .A(datapath_1_RegisterFile_regfile_mem_7__19_), .B(_5265__bF_buf89), .C(_5545__bF_buf1), .Y(_5565_) );
OAI21X1 OAI21X1_535 ( .A(_5314__bF_buf1), .B(_5545__bF_buf1), .C(_5565_), .Y(_1651_) );
NAND3X1 NAND3X1_410 ( .A(datapath_1_RegisterFile_regfile_mem_7__20_), .B(_5265__bF_buf39), .C(_5545__bF_buf1), .Y(_5566_) );
OAI21X1 OAI21X1_536 ( .A(_5316__bF_buf1), .B(_5545__bF_buf1), .C(_5566_), .Y(_1652_) );
NAND3X1 NAND3X1_411 ( .A(datapath_1_RegisterFile_regfile_mem_7__21_), .B(_5265__bF_buf65), .C(_5545__bF_buf2), .Y(_5567_) );
OAI21X1 OAI21X1_537 ( .A(_5318__bF_buf2), .B(_5545__bF_buf2), .C(_5567_), .Y(_1653_) );
NAND3X1 NAND3X1_412 ( .A(datapath_1_RegisterFile_regfile_mem_7__22_), .B(_5265__bF_buf73), .C(_5545__bF_buf7), .Y(_5568_) );
OAI21X1 OAI21X1_538 ( .A(_5320__bF_buf4), .B(_5545__bF_buf7), .C(_5568_), .Y(_1654_) );
NAND3X1 NAND3X1_413 ( .A(datapath_1_RegisterFile_regfile_mem_7__23_), .B(_5265__bF_buf77), .C(_5545__bF_buf6), .Y(_5569_) );
OAI21X1 OAI21X1_539 ( .A(_5322__bF_buf1), .B(_5545__bF_buf6), .C(_5569_), .Y(_1655_) );
NAND3X1 NAND3X1_414 ( .A(datapath_1_RegisterFile_regfile_mem_7__24_), .B(_5265__bF_buf30), .C(_5545__bF_buf4), .Y(_5570_) );
OAI21X1 OAI21X1_540 ( .A(_5324__bF_buf4), .B(_5545__bF_buf4), .C(_5570_), .Y(_1656_) );
NAND3X1 NAND3X1_415 ( .A(datapath_1_RegisterFile_regfile_mem_7__25_), .B(_5265__bF_buf55), .C(_5545__bF_buf2), .Y(_5571_) );
OAI21X1 OAI21X1_541 ( .A(_5326__bF_buf0), .B(_5545__bF_buf2), .C(_5571_), .Y(_1657_) );
NAND3X1 NAND3X1_416 ( .A(datapath_1_RegisterFile_regfile_mem_7__26_), .B(_5265__bF_buf64), .C(_5545__bF_buf7), .Y(_5572_) );
OAI21X1 OAI21X1_542 ( .A(_5328__bF_buf3), .B(_5545__bF_buf7), .C(_5572_), .Y(_1658_) );
NAND3X1 NAND3X1_417 ( .A(datapath_1_RegisterFile_regfile_mem_7__27_), .B(_5265__bF_buf68), .C(_5545__bF_buf6), .Y(_5573_) );
OAI21X1 OAI21X1_543 ( .A(_5330__bF_buf4), .B(_5545__bF_buf6), .C(_5573_), .Y(_1659_) );
NAND3X1 NAND3X1_418 ( .A(datapath_1_RegisterFile_regfile_mem_7__28_), .B(_5265__bF_buf30), .C(_5545__bF_buf4), .Y(_5574_) );
OAI21X1 OAI21X1_544 ( .A(_5332__bF_buf0), .B(_5545__bF_buf4), .C(_5574_), .Y(_1660_) );
NAND3X1 NAND3X1_419 ( .A(datapath_1_RegisterFile_regfile_mem_7__29_), .B(_5265__bF_buf93), .C(_5545__bF_buf3), .Y(_5575_) );
OAI21X1 OAI21X1_545 ( .A(_5334__bF_buf1), .B(_5545__bF_buf3), .C(_5575_), .Y(_1661_) );
NAND3X1 NAND3X1_420 ( .A(datapath_1_RegisterFile_regfile_mem_7__30_), .B(_5265__bF_buf97), .C(_5545__bF_buf5), .Y(_5576_) );
OAI21X1 OAI21X1_546 ( .A(_5336__bF_buf2), .B(_5545__bF_buf5), .C(_5576_), .Y(_1662_) );
NAND3X1 NAND3X1_421 ( .A(datapath_1_RegisterFile_regfile_mem_7__31_), .B(_5265__bF_buf77), .C(_5545__bF_buf6), .Y(_5577_) );
OAI21X1 OAI21X1_547 ( .A(_5338__bF_buf0), .B(_5545__bF_buf6), .C(_5577_), .Y(_1663_) );
NAND2X1 NAND2X1_371 ( .A(datapath_1_A3_3_), .B(_5267_), .Y(_5578_) );
NOR2X1 NOR2X1_136 ( .A(datapath_1_A3_2_), .B(_5578_), .Y(_5579_) );
NAND2X1 NAND2X1_372 ( .A(_5274_), .B(_5579_), .Y(_5580_) );
NAND3X1 NAND3X1_422 ( .A(datapath_1_RegisterFile_regfile_mem_8__0_), .B(_5265__bF_buf23), .C(_5580__bF_buf4), .Y(_5581_) );
OAI21X1 OAI21X1_548 ( .A(_5276__bF_buf0), .B(_5580__bF_buf4), .C(_5581_), .Y(_1664_) );
NAND3X1 NAND3X1_423 ( .A(datapath_1_RegisterFile_regfile_mem_8__1_), .B(_5265__bF_buf56), .C(_5580__bF_buf5), .Y(_5582_) );
OAI21X1 OAI21X1_549 ( .A(_5278__bF_buf0), .B(_5580__bF_buf5), .C(_5582_), .Y(_1665_) );
NAND3X1 NAND3X1_424 ( .A(datapath_1_RegisterFile_regfile_mem_8__2_), .B(_5265__bF_buf43), .C(_5580__bF_buf0), .Y(_5583_) );
OAI21X1 OAI21X1_550 ( .A(_5280__bF_buf2), .B(_5580__bF_buf0), .C(_5583_), .Y(_1666_) );
NAND3X1 NAND3X1_425 ( .A(datapath_1_RegisterFile_regfile_mem_8__3_), .B(_5265__bF_buf56), .C(_5580__bF_buf5), .Y(_5584_) );
OAI21X1 OAI21X1_551 ( .A(_5282__bF_buf0), .B(_5580__bF_buf5), .C(_5584_), .Y(_1667_) );
NAND3X1 NAND3X1_426 ( .A(datapath_1_RegisterFile_regfile_mem_8__4_), .B(_5265__bF_buf43), .C(_5580__bF_buf0), .Y(_5585_) );
OAI21X1 OAI21X1_552 ( .A(_5284__bF_buf4), .B(_5580__bF_buf0), .C(_5585_), .Y(_1668_) );
NAND3X1 NAND3X1_427 ( .A(datapath_1_RegisterFile_regfile_mem_8__5_), .B(_5265__bF_buf98), .C(_5580__bF_buf2), .Y(_5586_) );
OAI21X1 OAI21X1_553 ( .A(_5286__bF_buf0), .B(_5580__bF_buf2), .C(_5586_), .Y(_1669_) );
NAND3X1 NAND3X1_428 ( .A(datapath_1_RegisterFile_regfile_mem_8__6_), .B(_5265__bF_buf74), .C(_5580__bF_buf1), .Y(_5587_) );
OAI21X1 OAI21X1_554 ( .A(_5288__bF_buf3), .B(_5580__bF_buf1), .C(_5587_), .Y(_1670_) );
NAND3X1 NAND3X1_429 ( .A(datapath_1_RegisterFile_regfile_mem_8__7_), .B(_5265__bF_buf70), .C(_5580__bF_buf7), .Y(_5588_) );
OAI21X1 OAI21X1_555 ( .A(_5290__bF_buf1), .B(_5580__bF_buf7), .C(_5588_), .Y(_1671_) );
NAND3X1 NAND3X1_430 ( .A(datapath_1_RegisterFile_regfile_mem_8__8_), .B(_5265__bF_buf74), .C(_5580__bF_buf0), .Y(_5589_) );
OAI21X1 OAI21X1_556 ( .A(_5292__bF_buf3), .B(_5580__bF_buf0), .C(_5589_), .Y(_1672_) );
NAND3X1 NAND3X1_431 ( .A(datapath_1_RegisterFile_regfile_mem_8__9_), .B(_5265__bF_buf42), .C(_5580__bF_buf3), .Y(_5590_) );
OAI21X1 OAI21X1_557 ( .A(_5294__bF_buf3), .B(_5580__bF_buf3), .C(_5590_), .Y(_1673_) );
NAND3X1 NAND3X1_432 ( .A(datapath_1_RegisterFile_regfile_mem_8__10_), .B(_5265__bF_buf83), .C(_5580__bF_buf1), .Y(_5591_) );
OAI21X1 OAI21X1_558 ( .A(_5296__bF_buf3), .B(_5580__bF_buf1), .C(_5591_), .Y(_1674_) );
NAND3X1 NAND3X1_433 ( .A(datapath_1_RegisterFile_regfile_mem_8__11_), .B(_5265__bF_buf30), .C(_5580__bF_buf7), .Y(_5592_) );
OAI21X1 OAI21X1_559 ( .A(_5298__bF_buf3), .B(_5580__bF_buf7), .C(_5592_), .Y(_1675_) );
NAND3X1 NAND3X1_434 ( .A(datapath_1_RegisterFile_regfile_mem_8__12_), .B(_5265__bF_buf43), .C(_5580__bF_buf0), .Y(_5593_) );
OAI21X1 OAI21X1_560 ( .A(_5300__bF_buf1), .B(_5580__bF_buf0), .C(_5593_), .Y(_1676_) );
NAND3X1 NAND3X1_435 ( .A(datapath_1_RegisterFile_regfile_mem_8__13_), .B(_5265__bF_buf52), .C(_5580__bF_buf2), .Y(_5594_) );
OAI21X1 OAI21X1_561 ( .A(_5302__bF_buf4), .B(_5580__bF_buf2), .C(_5594_), .Y(_1677_) );
NAND3X1 NAND3X1_436 ( .A(datapath_1_RegisterFile_regfile_mem_8__14_), .B(_5265__bF_buf42), .C(_5580__bF_buf3), .Y(_5595_) );
OAI21X1 OAI21X1_562 ( .A(_5304__bF_buf3), .B(_5580__bF_buf3), .C(_5595_), .Y(_1678_) );
NAND3X1 NAND3X1_437 ( .A(datapath_1_RegisterFile_regfile_mem_8__15_), .B(_5265__bF_buf57), .C(_5580__bF_buf6), .Y(_5596_) );
OAI21X1 OAI21X1_563 ( .A(_5306__bF_buf3), .B(_5580__bF_buf6), .C(_5596_), .Y(_1679_) );
NAND3X1 NAND3X1_438 ( .A(datapath_1_RegisterFile_regfile_mem_8__16_), .B(_5265__bF_buf86), .C(_5580__bF_buf6), .Y(_5597_) );
OAI21X1 OAI21X1_564 ( .A(_5308__bF_buf0), .B(_5580__bF_buf6), .C(_5597_), .Y(_1680_) );
NAND3X1 NAND3X1_439 ( .A(datapath_1_RegisterFile_regfile_mem_8__17_), .B(_5265__bF_buf72), .C(_5580__bF_buf4), .Y(_5598_) );
OAI21X1 OAI21X1_565 ( .A(_5310__bF_buf4), .B(_5580__bF_buf4), .C(_5598_), .Y(_1575_) );
NAND3X1 NAND3X1_440 ( .A(datapath_1_RegisterFile_regfile_mem_8__18_), .B(_5265__bF_buf52), .C(_5580__bF_buf2), .Y(_5599_) );
OAI21X1 OAI21X1_566 ( .A(_5312__bF_buf0), .B(_5580__bF_buf2), .C(_5599_), .Y(_1576_) );
NAND3X1 NAND3X1_441 ( .A(datapath_1_RegisterFile_regfile_mem_8__19_), .B(_5265__bF_buf39), .C(_5580__bF_buf7), .Y(_5600_) );
OAI21X1 OAI21X1_567 ( .A(_5314__bF_buf1), .B(_5580__bF_buf7), .C(_5600_), .Y(_1577_) );
NAND3X1 NAND3X1_442 ( .A(datapath_1_RegisterFile_regfile_mem_8__20_), .B(_5265__bF_buf94), .C(_5580__bF_buf5), .Y(_5601_) );
OAI21X1 OAI21X1_568 ( .A(_5316__bF_buf3), .B(_5580__bF_buf5), .C(_5601_), .Y(_1578_) );
NAND3X1 NAND3X1_443 ( .A(datapath_1_RegisterFile_regfile_mem_8__21_), .B(_5265__bF_buf74), .C(_5580__bF_buf1), .Y(_5602_) );
OAI21X1 OAI21X1_569 ( .A(_5318__bF_buf0), .B(_5580__bF_buf1), .C(_5602_), .Y(_1579_) );
NAND3X1 NAND3X1_444 ( .A(datapath_1_RegisterFile_regfile_mem_8__22_), .B(_5265__bF_buf98), .C(_5580__bF_buf2), .Y(_5603_) );
OAI21X1 OAI21X1_570 ( .A(_5320__bF_buf2), .B(_5580__bF_buf2), .C(_5603_), .Y(_1580_) );
NAND3X1 NAND3X1_445 ( .A(datapath_1_RegisterFile_regfile_mem_8__23_), .B(_5265__bF_buf7), .C(_5580__bF_buf3), .Y(_5604_) );
OAI21X1 OAI21X1_571 ( .A(_5322__bF_buf3), .B(_5580__bF_buf3), .C(_5604_), .Y(_1581_) );
NAND3X1 NAND3X1_446 ( .A(datapath_1_RegisterFile_regfile_mem_8__24_), .B(_5265__bF_buf70), .C(_5580__bF_buf6), .Y(_5605_) );
OAI21X1 OAI21X1_572 ( .A(_5324__bF_buf0), .B(_5580__bF_buf6), .C(_5605_), .Y(_1681_) );
NAND3X1 NAND3X1_447 ( .A(datapath_1_RegisterFile_regfile_mem_8__25_), .B(_5265__bF_buf26), .C(_5580__bF_buf5), .Y(_5606_) );
OAI21X1 OAI21X1_573 ( .A(_5326__bF_buf1), .B(_5580__bF_buf5), .C(_5606_), .Y(_1582_) );
NAND3X1 NAND3X1_448 ( .A(datapath_1_RegisterFile_regfile_mem_8__26_), .B(_5265__bF_buf51), .C(_5580__bF_buf4), .Y(_5607_) );
OAI21X1 OAI21X1_574 ( .A(_5328__bF_buf2), .B(_5580__bF_buf4), .C(_5607_), .Y(_1583_) );
NAND3X1 NAND3X1_449 ( .A(datapath_1_RegisterFile_regfile_mem_8__27_), .B(_5265__bF_buf6), .C(_5580__bF_buf4), .Y(_5608_) );
OAI21X1 OAI21X1_575 ( .A(_5330__bF_buf3), .B(_5580__bF_buf4), .C(_5608_), .Y(_1584_) );
NAND3X1 NAND3X1_450 ( .A(datapath_1_RegisterFile_regfile_mem_8__28_), .B(_5265__bF_buf94), .C(_5580__bF_buf6), .Y(_5609_) );
OAI21X1 OAI21X1_576 ( .A(_5332__bF_buf1), .B(_5580__bF_buf6), .C(_5609_), .Y(_1585_) );
NAND3X1 NAND3X1_451 ( .A(datapath_1_RegisterFile_regfile_mem_8__29_), .B(_5265__bF_buf39), .C(_5580__bF_buf7), .Y(_5610_) );
OAI21X1 OAI21X1_577 ( .A(_5334__bF_buf1), .B(_5580__bF_buf7), .C(_5610_), .Y(_1586_) );
NAND3X1 NAND3X1_452 ( .A(datapath_1_RegisterFile_regfile_mem_8__30_), .B(_5265__bF_buf23), .C(_5580__bF_buf1), .Y(_5611_) );
OAI21X1 OAI21X1_578 ( .A(_5336__bF_buf4), .B(_5580__bF_buf1), .C(_5611_), .Y(_1587_) );
NAND3X1 NAND3X1_453 ( .A(datapath_1_RegisterFile_regfile_mem_8__31_), .B(_5265__bF_buf68), .C(_5580__bF_buf3), .Y(_5612_) );
OAI21X1 OAI21X1_579 ( .A(_5338__bF_buf0), .B(_5580__bF_buf3), .C(_5612_), .Y(_1588_) );
NAND2X1 NAND2X1_373 ( .A(_5341_), .B(_5579_), .Y(_5613_) );
NAND3X1 NAND3X1_454 ( .A(datapath_1_RegisterFile_regfile_mem_9__0_), .B(_5265__bF_buf83), .C(_5613__bF_buf1), .Y(_5614_) );
OAI21X1 OAI21X1_580 ( .A(_5276__bF_buf2), .B(_5613__bF_buf1), .C(_5614_), .Y(_1589_) );
NAND3X1 NAND3X1_455 ( .A(datapath_1_RegisterFile_regfile_mem_9__1_), .B(_5265__bF_buf91), .C(_5613__bF_buf6), .Y(_5615_) );
OAI21X1 OAI21X1_581 ( .A(_5278__bF_buf0), .B(_5613__bF_buf6), .C(_5615_), .Y(_1599_) );
NAND3X1 NAND3X1_456 ( .A(datapath_1_RegisterFile_regfile_mem_9__2_), .B(_5265__bF_buf26), .C(_5613__bF_buf4), .Y(_5616_) );
OAI21X1 OAI21X1_582 ( .A(_5280__bF_buf1), .B(_5613__bF_buf4), .C(_5616_), .Y(_1609_) );
NAND3X1 NAND3X1_457 ( .A(datapath_1_RegisterFile_regfile_mem_9__3_), .B(_5265__bF_buf35), .C(_5613__bF_buf4), .Y(_5617_) );
OAI21X1 OAI21X1_583 ( .A(_5282__bF_buf0), .B(_5613__bF_buf4), .C(_5617_), .Y(_1612_) );
NAND3X1 NAND3X1_458 ( .A(datapath_1_RegisterFile_regfile_mem_9__4_), .B(_5265__bF_buf83), .C(_5613__bF_buf1), .Y(_5618_) );
OAI21X1 OAI21X1_584 ( .A(_5284__bF_buf4), .B(_5613__bF_buf1), .C(_5618_), .Y(_1613_) );
NAND3X1 NAND3X1_459 ( .A(datapath_1_RegisterFile_regfile_mem_9__5_), .B(_5265__bF_buf21), .C(_5613__bF_buf3), .Y(_5619_) );
OAI21X1 OAI21X1_585 ( .A(_5286__bF_buf1), .B(_5613__bF_buf3), .C(_5619_), .Y(_1614_) );
NAND3X1 NAND3X1_460 ( .A(datapath_1_RegisterFile_regfile_mem_9__6_), .B(_5265__bF_buf0), .C(_5613__bF_buf6), .Y(_5620_) );
OAI21X1 OAI21X1_586 ( .A(_5288__bF_buf2), .B(_5613__bF_buf6), .C(_5620_), .Y(_1615_) );
NAND3X1 NAND3X1_461 ( .A(datapath_1_RegisterFile_regfile_mem_9__7_), .B(_5265__bF_buf76), .C(_5613__bF_buf5), .Y(_5621_) );
OAI21X1 OAI21X1_587 ( .A(_5290__bF_buf1), .B(_5613__bF_buf5), .C(_5621_), .Y(_1682_) );
NAND3X1 NAND3X1_462 ( .A(datapath_1_RegisterFile_regfile_mem_9__8_), .B(_5265__bF_buf0), .C(_5613__bF_buf6), .Y(_5622_) );
OAI21X1 OAI21X1_588 ( .A(_5292__bF_buf3), .B(_5613__bF_buf6), .C(_5622_), .Y(_1616_) );
NAND3X1 NAND3X1_463 ( .A(datapath_1_RegisterFile_regfile_mem_9__9_), .B(_5265__bF_buf98), .C(_5613__bF_buf7), .Y(_5623_) );
OAI21X1 OAI21X1_589 ( .A(_5294__bF_buf2), .B(_5613__bF_buf7), .C(_5623_), .Y(_1617_) );
NAND3X1 NAND3X1_464 ( .A(datapath_1_RegisterFile_regfile_mem_9__10_), .B(_5265__bF_buf83), .C(_5613__bF_buf0), .Y(_5624_) );
OAI21X1 OAI21X1_590 ( .A(_5296__bF_buf3), .B(_5613__bF_buf0), .C(_5624_), .Y(_1590_) );
NAND3X1 NAND3X1_465 ( .A(datapath_1_RegisterFile_regfile_mem_9__11_), .B(_5265__bF_buf30), .C(_5613__bF_buf5), .Y(_5625_) );
OAI21X1 OAI21X1_591 ( .A(_5298__bF_buf3), .B(_5613__bF_buf5), .C(_5625_), .Y(_1591_) );
NAND3X1 NAND3X1_466 ( .A(datapath_1_RegisterFile_regfile_mem_9__12_), .B(_5265__bF_buf43), .C(_5613__bF_buf6), .Y(_5626_) );
OAI21X1 OAI21X1_592 ( .A(_5300__bF_buf3), .B(_5613__bF_buf6), .C(_5626_), .Y(_1592_) );
NAND3X1 NAND3X1_467 ( .A(datapath_1_RegisterFile_regfile_mem_9__13_), .B(_5265__bF_buf21), .C(_5613__bF_buf7), .Y(_5627_) );
OAI21X1 OAI21X1_593 ( .A(_5302__bF_buf4), .B(_5613__bF_buf7), .C(_5627_), .Y(_1593_) );
NAND3X1 NAND3X1_468 ( .A(datapath_1_RegisterFile_regfile_mem_9__14_), .B(_5265__bF_buf87), .C(_5613__bF_buf0), .Y(_5628_) );
OAI21X1 OAI21X1_594 ( .A(_5304__bF_buf1), .B(_5613__bF_buf0), .C(_5628_), .Y(_1594_) );
NAND3X1 NAND3X1_469 ( .A(datapath_1_RegisterFile_regfile_mem_9__15_), .B(_5265__bF_buf70), .C(_5613__bF_buf2), .Y(_5629_) );
OAI21X1 OAI21X1_595 ( .A(_5306__bF_buf1), .B(_5613__bF_buf2), .C(_5629_), .Y(_1595_) );
NAND3X1 NAND3X1_470 ( .A(datapath_1_RegisterFile_regfile_mem_9__16_), .B(_5265__bF_buf86), .C(_5613__bF_buf2), .Y(_5630_) );
OAI21X1 OAI21X1_596 ( .A(_5308__bF_buf0), .B(_5613__bF_buf2), .C(_5630_), .Y(_1596_) );
NAND3X1 NAND3X1_471 ( .A(datapath_1_RegisterFile_regfile_mem_9__17_), .B(_5265__bF_buf83), .C(_5613__bF_buf0), .Y(_5631_) );
OAI21X1 OAI21X1_597 ( .A(_5310__bF_buf4), .B(_5613__bF_buf0), .C(_5631_), .Y(_1683_) );
NAND3X1 NAND3X1_472 ( .A(datapath_1_RegisterFile_regfile_mem_9__18_), .B(_5265__bF_buf52), .C(_5613__bF_buf7), .Y(_5632_) );
OAI21X1 OAI21X1_598 ( .A(_5312__bF_buf0), .B(_5613__bF_buf7), .C(_5632_), .Y(_1597_) );
NAND3X1 NAND3X1_473 ( .A(datapath_1_RegisterFile_regfile_mem_9__19_), .B(_5265__bF_buf39), .C(_5613__bF_buf5), .Y(_5633_) );
OAI21X1 OAI21X1_599 ( .A(_5314__bF_buf1), .B(_5613__bF_buf5), .C(_5633_), .Y(_1598_) );
NAND3X1 NAND3X1_474 ( .A(datapath_1_RegisterFile_regfile_mem_9__20_), .B(_5265__bF_buf96), .C(_5613__bF_buf4), .Y(_5634_) );
OAI21X1 OAI21X1_600 ( .A(_5316__bF_buf3), .B(_5613__bF_buf4), .C(_5634_), .Y(_1600_) );
NAND3X1 NAND3X1_475 ( .A(datapath_1_RegisterFile_regfile_mem_9__21_), .B(_5265__bF_buf83), .C(_5613__bF_buf1), .Y(_5635_) );
OAI21X1 OAI21X1_601 ( .A(_5318__bF_buf0), .B(_5613__bF_buf1), .C(_5635_), .Y(_1601_) );
NAND3X1 NAND3X1_476 ( .A(datapath_1_RegisterFile_regfile_mem_9__22_), .B(_5265__bF_buf98), .C(_5613__bF_buf7), .Y(_5636_) );
OAI21X1 OAI21X1_602 ( .A(_5320__bF_buf2), .B(_5613__bF_buf7), .C(_5636_), .Y(_1602_) );
NAND3X1 NAND3X1_477 ( .A(datapath_1_RegisterFile_regfile_mem_9__23_), .B(_5265__bF_buf21), .C(_5613__bF_buf3), .Y(_5637_) );
OAI21X1 OAI21X1_603 ( .A(_5322__bF_buf2), .B(_5613__bF_buf3), .C(_5637_), .Y(_1603_) );
NAND3X1 NAND3X1_478 ( .A(datapath_1_RegisterFile_regfile_mem_9__24_), .B(_5265__bF_buf76), .C(_5613__bF_buf5), .Y(_5638_) );
OAI21X1 OAI21X1_604 ( .A(_5324__bF_buf0), .B(_5613__bF_buf5), .C(_5638_), .Y(_1604_) );
NAND3X1 NAND3X1_479 ( .A(datapath_1_RegisterFile_regfile_mem_9__25_), .B(_5265__bF_buf26), .C(_5613__bF_buf4), .Y(_5639_) );
OAI21X1 OAI21X1_605 ( .A(_5326__bF_buf1), .B(_5613__bF_buf4), .C(_5639_), .Y(_1605_) );
NAND3X1 NAND3X1_480 ( .A(datapath_1_RegisterFile_regfile_mem_9__26_), .B(_5265__bF_buf51), .C(_5613__bF_buf3), .Y(_5640_) );
OAI21X1 OAI21X1_606 ( .A(_5328__bF_buf3), .B(_5613__bF_buf3), .C(_5640_), .Y(_1606_) );
NAND3X1 NAND3X1_481 ( .A(datapath_1_RegisterFile_regfile_mem_9__27_), .B(_5265__bF_buf42), .C(_5613__bF_buf0), .Y(_5641_) );
OAI21X1 OAI21X1_607 ( .A(_5330__bF_buf3), .B(_5613__bF_buf0), .C(_5641_), .Y(_1684_) );
NAND3X1 NAND3X1_482 ( .A(datapath_1_RegisterFile_regfile_mem_9__28_), .B(_5265__bF_buf94), .C(_5613__bF_buf2), .Y(_5642_) );
OAI21X1 OAI21X1_608 ( .A(_5332__bF_buf1), .B(_5613__bF_buf2), .C(_5642_), .Y(_1607_) );
NAND3X1 NAND3X1_483 ( .A(datapath_1_RegisterFile_regfile_mem_9__29_), .B(_5265__bF_buf96), .C(_5613__bF_buf2), .Y(_5643_) );
OAI21X1 OAI21X1_609 ( .A(_5334__bF_buf4), .B(_5613__bF_buf2), .C(_5643_), .Y(_1608_) );
NAND3X1 NAND3X1_484 ( .A(datapath_1_RegisterFile_regfile_mem_9__30_), .B(_5265__bF_buf83), .C(_5613__bF_buf1), .Y(_5644_) );
OAI21X1 OAI21X1_610 ( .A(_5336__bF_buf4), .B(_5613__bF_buf1), .C(_5644_), .Y(_1610_) );
NAND3X1 NAND3X1_485 ( .A(datapath_1_RegisterFile_regfile_mem_9__31_), .B(_5265__bF_buf7), .C(_5613__bF_buf3), .Y(_5645_) );
OAI21X1 OAI21X1_611 ( .A(_5338__bF_buf3), .B(_5613__bF_buf3), .C(_5645_), .Y(_1611_) );
NAND2X1 NAND2X1_374 ( .A(_5376_), .B(_5579_), .Y(_5646_) );
NAND3X1 NAND3X1_486 ( .A(datapath_1_RegisterFile_regfile_mem_10__0_), .B(_5265__bF_buf83), .C(_5646__bF_buf2), .Y(_5647_) );
OAI21X1 OAI21X1_612 ( .A(_5276__bF_buf2), .B(_5646__bF_buf2), .C(_5647_), .Y(_869_) );
NAND3X1 NAND3X1_487 ( .A(datapath_1_RegisterFile_regfile_mem_10__1_), .B(_5265__bF_buf91), .C(_5646__bF_buf7), .Y(_5648_) );
OAI21X1 OAI21X1_613 ( .A(_5278__bF_buf0), .B(_5646__bF_buf7), .C(_5648_), .Y(_879_) );
NAND3X1 NAND3X1_488 ( .A(datapath_1_RegisterFile_regfile_mem_10__2_), .B(_5265__bF_buf50), .C(_5646__bF_buf6), .Y(_5649_) );
OAI21X1 OAI21X1_614 ( .A(_5280__bF_buf1), .B(_5646__bF_buf6), .C(_5649_), .Y(_1685_) );
NAND3X1 NAND3X1_489 ( .A(datapath_1_RegisterFile_regfile_mem_10__3_), .B(_5265__bF_buf56), .C(_5646__bF_buf6), .Y(_5650_) );
OAI21X1 OAI21X1_615 ( .A(_5282__bF_buf0), .B(_5646__bF_buf6), .C(_5650_), .Y(_884_) );
NAND3X1 NAND3X1_490 ( .A(datapath_1_RegisterFile_regfile_mem_10__4_), .B(_5265__bF_buf92), .C(_5646__bF_buf3), .Y(_5651_) );
OAI21X1 OAI21X1_616 ( .A(_5284__bF_buf4), .B(_5646__bF_buf3), .C(_5651_), .Y(_885_) );
NAND3X1 NAND3X1_491 ( .A(datapath_1_RegisterFile_regfile_mem_10__5_), .B(_5265__bF_buf60), .C(_5646__bF_buf0), .Y(_5652_) );
OAI21X1 OAI21X1_617 ( .A(_5286__bF_buf0), .B(_5646__bF_buf0), .C(_5652_), .Y(_886_) );
NAND3X1 NAND3X1_492 ( .A(datapath_1_RegisterFile_regfile_mem_10__6_), .B(_5265__bF_buf92), .C(_5646__bF_buf3), .Y(_5653_) );
OAI21X1 OAI21X1_618 ( .A(_5288__bF_buf3), .B(_5646__bF_buf3), .C(_5653_), .Y(_887_) );
NAND3X1 NAND3X1_493 ( .A(datapath_1_RegisterFile_regfile_mem_10__7_), .B(_5265__bF_buf76), .C(_5646__bF_buf1), .Y(_5654_) );
OAI21X1 OAI21X1_619 ( .A(_5290__bF_buf1), .B(_5646__bF_buf1), .C(_5654_), .Y(_888_) );
NAND3X1 NAND3X1_494 ( .A(datapath_1_RegisterFile_regfile_mem_10__8_), .B(_5265__bF_buf43), .C(_5646__bF_buf7), .Y(_5655_) );
OAI21X1 OAI21X1_620 ( .A(_5292__bF_buf3), .B(_5646__bF_buf7), .C(_5655_), .Y(_889_) );
NAND3X1 NAND3X1_495 ( .A(datapath_1_RegisterFile_regfile_mem_10__9_), .B(_5265__bF_buf60), .C(_5646__bF_buf0), .Y(_5656_) );
OAI21X1 OAI21X1_621 ( .A(_5294__bF_buf2), .B(_5646__bF_buf0), .C(_5656_), .Y(_890_) );
NAND3X1 NAND3X1_496 ( .A(datapath_1_RegisterFile_regfile_mem_10__10_), .B(_5265__bF_buf0), .C(_5646__bF_buf7), .Y(_5657_) );
OAI21X1 OAI21X1_622 ( .A(_5296__bF_buf4), .B(_5646__bF_buf7), .C(_5657_), .Y(_870_) );
NAND3X1 NAND3X1_497 ( .A(datapath_1_RegisterFile_regfile_mem_10__11_), .B(_5265__bF_buf85), .C(_5646__bF_buf5), .Y(_5658_) );
OAI21X1 OAI21X1_623 ( .A(_5298__bF_buf3), .B(_5646__bF_buf5), .C(_5658_), .Y(_871_) );
NAND3X1 NAND3X1_498 ( .A(datapath_1_RegisterFile_regfile_mem_10__12_), .B(_5265__bF_buf43), .C(_5646__bF_buf7), .Y(_5659_) );
OAI21X1 OAI21X1_624 ( .A(_5300__bF_buf3), .B(_5646__bF_buf7), .C(_5659_), .Y(_1686_) );
NAND3X1 NAND3X1_499 ( .A(datapath_1_RegisterFile_regfile_mem_10__13_), .B(_5265__bF_buf48), .C(_5646__bF_buf0), .Y(_5660_) );
OAI21X1 OAI21X1_625 ( .A(_5302__bF_buf2), .B(_5646__bF_buf0), .C(_5660_), .Y(_872_) );
NAND3X1 NAND3X1_500 ( .A(datapath_1_RegisterFile_regfile_mem_10__14_), .B(_5265__bF_buf6), .C(_5646__bF_buf2), .Y(_5661_) );
OAI21X1 OAI21X1_626 ( .A(_5304__bF_buf0), .B(_5646__bF_buf2), .C(_5661_), .Y(_873_) );
NAND3X1 NAND3X1_501 ( .A(datapath_1_RegisterFile_regfile_mem_10__15_), .B(_5265__bF_buf57), .C(_5646__bF_buf5), .Y(_5662_) );
OAI21X1 OAI21X1_627 ( .A(_5306__bF_buf1), .B(_5646__bF_buf5), .C(_5662_), .Y(_874_) );
NAND3X1 NAND3X1_502 ( .A(datapath_1_RegisterFile_regfile_mem_10__16_), .B(_5265__bF_buf57), .C(_5646__bF_buf5), .Y(_5663_) );
OAI21X1 OAI21X1_628 ( .A(_5308__bF_buf0), .B(_5646__bF_buf5), .C(_5663_), .Y(_875_) );
NAND3X1 NAND3X1_503 ( .A(datapath_1_RegisterFile_regfile_mem_10__17_), .B(_5265__bF_buf23), .C(_5646__bF_buf3), .Y(_5664_) );
OAI21X1 OAI21X1_629 ( .A(_5310__bF_buf4), .B(_5646__bF_buf3), .C(_5664_), .Y(_876_) );
NAND3X1 NAND3X1_504 ( .A(datapath_1_RegisterFile_regfile_mem_10__18_), .B(_5265__bF_buf52), .C(_5646__bF_buf4), .Y(_5665_) );
OAI21X1 OAI21X1_630 ( .A(_5312__bF_buf1), .B(_5646__bF_buf4), .C(_5665_), .Y(_877_) );
NAND3X1 NAND3X1_505 ( .A(datapath_1_RegisterFile_regfile_mem_10__19_), .B(_5265__bF_buf44), .C(_5646__bF_buf6), .Y(_5666_) );
OAI21X1 OAI21X1_631 ( .A(_5314__bF_buf1), .B(_5646__bF_buf6), .C(_5666_), .Y(_878_) );
NAND3X1 NAND3X1_506 ( .A(datapath_1_RegisterFile_regfile_mem_10__20_), .B(_5265__bF_buf96), .C(_5646__bF_buf1), .Y(_5667_) );
OAI21X1 OAI21X1_632 ( .A(_5316__bF_buf3), .B(_5646__bF_buf1), .C(_5667_), .Y(_880_) );
NAND3X1 NAND3X1_507 ( .A(datapath_1_RegisterFile_regfile_mem_10__21_), .B(_5265__bF_buf92), .C(_5646__bF_buf3), .Y(_5668_) );
OAI21X1 OAI21X1_633 ( .A(_5318__bF_buf4), .B(_5646__bF_buf3), .C(_5668_), .Y(_881_) );
NAND3X1 NAND3X1_508 ( .A(datapath_1_RegisterFile_regfile_mem_10__22_), .B(_5265__bF_buf60), .C(_5646__bF_buf0), .Y(_5669_) );
OAI21X1 OAI21X1_634 ( .A(_5320__bF_buf4), .B(_5646__bF_buf0), .C(_5669_), .Y(_1687_) );
NAND3X1 NAND3X1_509 ( .A(datapath_1_RegisterFile_regfile_mem_10__23_), .B(_5265__bF_buf7), .C(_5646__bF_buf4), .Y(_5670_) );
OAI21X1 OAI21X1_635 ( .A(_5322__bF_buf3), .B(_5646__bF_buf4), .C(_5670_), .Y(_882_) );
NAND3X1 NAND3X1_510 ( .A(datapath_1_RegisterFile_regfile_mem_10__24_), .B(_5265__bF_buf70), .C(_5646__bF_buf1), .Y(_5671_) );
OAI21X1 OAI21X1_636 ( .A(_5324__bF_buf3), .B(_5646__bF_buf1), .C(_5671_), .Y(_883_) );
NAND3X1 NAND3X1_511 ( .A(datapath_1_RegisterFile_regfile_mem_10__25_), .B(_5265__bF_buf96), .C(_5646__bF_buf1), .Y(_5672_) );
OAI21X1 OAI21X1_637 ( .A(_5326__bF_buf1), .B(_5646__bF_buf1), .C(_5672_), .Y(_1688_) );
NAND3X1 NAND3X1_512 ( .A(datapath_1_RegisterFile_regfile_mem_10__26_), .B(_5265__bF_buf51), .C(_5646__bF_buf2), .Y(_5673_) );
OAI21X1 OAI21X1_638 ( .A(_5328__bF_buf2), .B(_5646__bF_buf2), .C(_5673_), .Y(_1689_) );
NAND3X1 NAND3X1_513 ( .A(datapath_1_RegisterFile_regfile_mem_10__27_), .B(_5265__bF_buf7), .C(_5646__bF_buf4), .Y(_5674_) );
OAI21X1 OAI21X1_639 ( .A(_5330__bF_buf3), .B(_5646__bF_buf4), .C(_5674_), .Y(_1690_) );
NAND3X1 NAND3X1_514 ( .A(datapath_1_RegisterFile_regfile_mem_10__28_), .B(_5265__bF_buf85), .C(_5646__bF_buf5), .Y(_5675_) );
OAI21X1 OAI21X1_640 ( .A(_5332__bF_buf4), .B(_5646__bF_buf5), .C(_5675_), .Y(_1691_) );
NAND3X1 NAND3X1_515 ( .A(datapath_1_RegisterFile_regfile_mem_10__29_), .B(_5265__bF_buf44), .C(_5646__bF_buf6), .Y(_5676_) );
OAI21X1 OAI21X1_641 ( .A(_5334__bF_buf1), .B(_5646__bF_buf6), .C(_5676_), .Y(_1692_) );
NAND3X1 NAND3X1_516 ( .A(datapath_1_RegisterFile_regfile_mem_10__30_), .B(_5265__bF_buf13), .C(_5646__bF_buf2), .Y(_5677_) );
OAI21X1 OAI21X1_642 ( .A(_5336__bF_buf4), .B(_5646__bF_buf2), .C(_5677_), .Y(_1693_) );
NAND3X1 NAND3X1_517 ( .A(datapath_1_RegisterFile_regfile_mem_10__31_), .B(_5265__bF_buf42), .C(_5646__bF_buf4), .Y(_5678_) );
OAI21X1 OAI21X1_643 ( .A(_5338__bF_buf0), .B(_5646__bF_buf4), .C(_5678_), .Y(_1694_) );
NAND2X1 NAND2X1_375 ( .A(_5410_), .B(_5579_), .Y(_5679_) );
NAND3X1 NAND3X1_518 ( .A(datapath_1_RegisterFile_regfile_mem_11__0_), .B(_5265__bF_buf23), .C(_5679__bF_buf1), .Y(_5680_) );
OAI21X1 OAI21X1_644 ( .A(_5276__bF_buf2), .B(_5679__bF_buf1), .C(_5680_), .Y(_891_) );
NAND3X1 NAND3X1_519 ( .A(datapath_1_RegisterFile_regfile_mem_11__1_), .B(_5265__bF_buf91), .C(_5679__bF_buf0), .Y(_5681_) );
OAI21X1 OAI21X1_645 ( .A(_5278__bF_buf0), .B(_5679__bF_buf0), .C(_5681_), .Y(_901_) );
NAND3X1 NAND3X1_520 ( .A(datapath_1_RegisterFile_regfile_mem_11__2_), .B(_5265__bF_buf0), .C(_5679__bF_buf3), .Y(_5682_) );
OAI21X1 OAI21X1_646 ( .A(_5280__bF_buf2), .B(_5679__bF_buf3), .C(_5682_), .Y(_911_) );
NAND3X1 NAND3X1_521 ( .A(datapath_1_RegisterFile_regfile_mem_11__3_), .B(_5265__bF_buf91), .C(_5679__bF_buf0), .Y(_5683_) );
OAI21X1 OAI21X1_647 ( .A(_5282__bF_buf0), .B(_5679__bF_buf0), .C(_5683_), .Y(_914_) );
NAND3X1 NAND3X1_522 ( .A(datapath_1_RegisterFile_regfile_mem_11__4_), .B(_5265__bF_buf72), .C(_5679__bF_buf5), .Y(_5684_) );
OAI21X1 OAI21X1_648 ( .A(_5284__bF_buf1), .B(_5679__bF_buf5), .C(_5684_), .Y(_915_) );
NAND3X1 NAND3X1_523 ( .A(datapath_1_RegisterFile_regfile_mem_11__5_), .B(_5265__bF_buf21), .C(_5679__bF_buf7), .Y(_5685_) );
OAI21X1 OAI21X1_649 ( .A(_5286__bF_buf1), .B(_5679__bF_buf7), .C(_5685_), .Y(_916_) );
NAND3X1 NAND3X1_524 ( .A(datapath_1_RegisterFile_regfile_mem_11__6_), .B(_5265__bF_buf92), .C(_5679__bF_buf5), .Y(_5686_) );
OAI21X1 OAI21X1_650 ( .A(_5288__bF_buf3), .B(_5679__bF_buf5), .C(_5686_), .Y(_917_) );
NAND3X1 NAND3X1_525 ( .A(datapath_1_RegisterFile_regfile_mem_11__7_), .B(_5265__bF_buf57), .C(_5679__bF_buf2), .Y(_5687_) );
OAI21X1 OAI21X1_651 ( .A(_5290__bF_buf4), .B(_5679__bF_buf2), .C(_5687_), .Y(_1695_) );
NAND3X1 NAND3X1_526 ( .A(datapath_1_RegisterFile_regfile_mem_11__8_), .B(_5265__bF_buf0), .C(_5679__bF_buf3), .Y(_5688_) );
OAI21X1 OAI21X1_652 ( .A(_5292__bF_buf3), .B(_5679__bF_buf3), .C(_5688_), .Y(_918_) );
NAND3X1 NAND3X1_527 ( .A(datapath_1_RegisterFile_regfile_mem_11__9_), .B(_5265__bF_buf21), .C(_5679__bF_buf4), .Y(_5689_) );
OAI21X1 OAI21X1_653 ( .A(_5294__bF_buf2), .B(_5679__bF_buf4), .C(_5689_), .Y(_919_) );
NAND3X1 NAND3X1_528 ( .A(datapath_1_RegisterFile_regfile_mem_11__10_), .B(_5265__bF_buf43), .C(_5679__bF_buf3), .Y(_5690_) );
OAI21X1 OAI21X1_654 ( .A(_5296__bF_buf4), .B(_5679__bF_buf3), .C(_5690_), .Y(_892_) );
NAND3X1 NAND3X1_529 ( .A(datapath_1_RegisterFile_regfile_mem_11__11_), .B(_5265__bF_buf70), .C(_5679__bF_buf6), .Y(_5691_) );
OAI21X1 OAI21X1_655 ( .A(_5298__bF_buf3), .B(_5679__bF_buf6), .C(_5691_), .Y(_893_) );
NAND3X1 NAND3X1_530 ( .A(datapath_1_RegisterFile_regfile_mem_11__12_), .B(_5265__bF_buf0), .C(_5679__bF_buf3), .Y(_5692_) );
OAI21X1 OAI21X1_656 ( .A(_5300__bF_buf3), .B(_5679__bF_buf3), .C(_5692_), .Y(_894_) );
NAND3X1 NAND3X1_531 ( .A(datapath_1_RegisterFile_regfile_mem_11__13_), .B(_5265__bF_buf52), .C(_5679__bF_buf4), .Y(_5693_) );
OAI21X1 OAI21X1_657 ( .A(_5302__bF_buf4), .B(_5679__bF_buf4), .C(_5693_), .Y(_895_) );
NAND3X1 NAND3X1_532 ( .A(datapath_1_RegisterFile_regfile_mem_11__14_), .B(_5265__bF_buf87), .C(_5679__bF_buf1), .Y(_5694_) );
OAI21X1 OAI21X1_658 ( .A(_5304__bF_buf1), .B(_5679__bF_buf1), .C(_5694_), .Y(_896_) );
NAND3X1 NAND3X1_533 ( .A(datapath_1_RegisterFile_regfile_mem_11__15_), .B(_5265__bF_buf76), .C(_5679__bF_buf2), .Y(_5695_) );
OAI21X1 OAI21X1_659 ( .A(_5306__bF_buf3), .B(_5679__bF_buf2), .C(_5695_), .Y(_897_) );
NAND3X1 NAND3X1_534 ( .A(datapath_1_RegisterFile_regfile_mem_11__16_), .B(_5265__bF_buf57), .C(_5679__bF_buf2), .Y(_5696_) );
OAI21X1 OAI21X1_660 ( .A(_5308__bF_buf0), .B(_5679__bF_buf2), .C(_5696_), .Y(_898_) );
NAND3X1 NAND3X1_535 ( .A(datapath_1_RegisterFile_regfile_mem_11__17_), .B(_5265__bF_buf72), .C(_5679__bF_buf5), .Y(_5697_) );
OAI21X1 OAI21X1_661 ( .A(_5310__bF_buf1), .B(_5679__bF_buf5), .C(_5697_), .Y(_1696_) );
NAND3X1 NAND3X1_536 ( .A(datapath_1_RegisterFile_regfile_mem_11__18_), .B(_5265__bF_buf98), .C(_5679__bF_buf4), .Y(_5698_) );
OAI21X1 OAI21X1_662 ( .A(_5312__bF_buf0), .B(_5679__bF_buf4), .C(_5698_), .Y(_899_) );
NAND3X1 NAND3X1_537 ( .A(datapath_1_RegisterFile_regfile_mem_11__19_), .B(_5265__bF_buf84), .C(_5679__bF_buf0), .Y(_5699_) );
OAI21X1 OAI21X1_663 ( .A(_5314__bF_buf3), .B(_5679__bF_buf0), .C(_5699_), .Y(_900_) );
NAND3X1 NAND3X1_538 ( .A(datapath_1_RegisterFile_regfile_mem_11__20_), .B(_5265__bF_buf84), .C(_5679__bF_buf0), .Y(_5700_) );
OAI21X1 OAI21X1_664 ( .A(_5316__bF_buf3), .B(_5679__bF_buf0), .C(_5700_), .Y(_902_) );
NAND3X1 NAND3X1_539 ( .A(datapath_1_RegisterFile_regfile_mem_11__21_), .B(_5265__bF_buf92), .C(_5679__bF_buf5), .Y(_5701_) );
OAI21X1 OAI21X1_665 ( .A(_5318__bF_buf0), .B(_5679__bF_buf5), .C(_5701_), .Y(_903_) );
NAND3X1 NAND3X1_540 ( .A(datapath_1_RegisterFile_regfile_mem_11__22_), .B(_5265__bF_buf98), .C(_5679__bF_buf4), .Y(_5702_) );
OAI21X1 OAI21X1_666 ( .A(_5320__bF_buf2), .B(_5679__bF_buf4), .C(_5702_), .Y(_904_) );
NAND3X1 NAND3X1_541 ( .A(datapath_1_RegisterFile_regfile_mem_11__23_), .B(_5265__bF_buf7), .C(_5679__bF_buf7), .Y(_5703_) );
OAI21X1 OAI21X1_667 ( .A(_5322__bF_buf3), .B(_5679__bF_buf7), .C(_5703_), .Y(_905_) );
NAND3X1 NAND3X1_542 ( .A(datapath_1_RegisterFile_regfile_mem_11__24_), .B(_5265__bF_buf86), .C(_5679__bF_buf2), .Y(_5704_) );
OAI21X1 OAI21X1_668 ( .A(_5324__bF_buf3), .B(_5679__bF_buf2), .C(_5704_), .Y(_906_) );
NAND3X1 NAND3X1_543 ( .A(datapath_1_RegisterFile_regfile_mem_11__25_), .B(_5265__bF_buf94), .C(_5679__bF_buf6), .Y(_5705_) );
OAI21X1 OAI21X1_669 ( .A(_5326__bF_buf1), .B(_5679__bF_buf6), .C(_5705_), .Y(_907_) );
NAND3X1 NAND3X1_544 ( .A(datapath_1_RegisterFile_regfile_mem_11__26_), .B(_5265__bF_buf51), .C(_5679__bF_buf7), .Y(_5706_) );
OAI21X1 OAI21X1_670 ( .A(_5328__bF_buf3), .B(_5679__bF_buf7), .C(_5706_), .Y(_908_) );
NAND3X1 NAND3X1_545 ( .A(datapath_1_RegisterFile_regfile_mem_11__27_), .B(_5265__bF_buf42), .C(_5679__bF_buf7), .Y(_5707_) );
OAI21X1 OAI21X1_671 ( .A(_5330__bF_buf3), .B(_5679__bF_buf7), .C(_5707_), .Y(_1697_) );
NAND3X1 NAND3X1_546 ( .A(datapath_1_RegisterFile_regfile_mem_11__28_), .B(_5265__bF_buf94), .C(_5679__bF_buf6), .Y(_5708_) );
OAI21X1 OAI21X1_672 ( .A(_5332__bF_buf1), .B(_5679__bF_buf6), .C(_5708_), .Y(_909_) );
NAND3X1 NAND3X1_547 ( .A(datapath_1_RegisterFile_regfile_mem_11__29_), .B(_5265__bF_buf94), .C(_5679__bF_buf6), .Y(_5709_) );
OAI21X1 OAI21X1_673 ( .A(_5334__bF_buf4), .B(_5679__bF_buf6), .C(_5709_), .Y(_910_) );
NAND3X1 NAND3X1_548 ( .A(datapath_1_RegisterFile_regfile_mem_11__30_), .B(_5265__bF_buf13), .C(_5679__bF_buf1), .Y(_5710_) );
OAI21X1 OAI21X1_674 ( .A(_5336__bF_buf4), .B(_5679__bF_buf1), .C(_5710_), .Y(_912_) );
NAND3X1 NAND3X1_549 ( .A(datapath_1_RegisterFile_regfile_mem_11__31_), .B(_5265__bF_buf6), .C(_5679__bF_buf1), .Y(_5711_) );
OAI21X1 OAI21X1_675 ( .A(_5338__bF_buf3), .B(_5679__bF_buf1), .C(_5711_), .Y(_913_) );
NOR2X1 NOR2X1_137 ( .A(_5444_), .B(_5578_), .Y(_5712_) );
NAND2X1 NAND2X1_376 ( .A(_5274_), .B(_5712_), .Y(_5713_) );
NAND3X1 NAND3X1_550 ( .A(datapath_1_RegisterFile_regfile_mem_12__0_), .B(_5265__bF_buf72), .C(_5713__bF_buf5), .Y(_5714_) );
OAI21X1 OAI21X1_676 ( .A(_5276__bF_buf0), .B(_5713__bF_buf5), .C(_5714_), .Y(_1698_) );
NAND3X1 NAND3X1_551 ( .A(datapath_1_RegisterFile_regfile_mem_12__1_), .B(_5265__bF_buf50), .C(_5713__bF_buf4), .Y(_5715_) );
OAI21X1 OAI21X1_677 ( .A(_5278__bF_buf2), .B(_5713__bF_buf4), .C(_5715_), .Y(_1699_) );
NAND3X1 NAND3X1_552 ( .A(datapath_1_RegisterFile_regfile_mem_12__2_), .B(_5265__bF_buf50), .C(_5713__bF_buf6), .Y(_5716_) );
OAI21X1 OAI21X1_678 ( .A(_5280__bF_buf1), .B(_5713__bF_buf6), .C(_5716_), .Y(_1700_) );
NAND3X1 NAND3X1_553 ( .A(datapath_1_RegisterFile_regfile_mem_12__3_), .B(_5265__bF_buf26), .C(_5713__bF_buf6), .Y(_5717_) );
OAI21X1 OAI21X1_679 ( .A(_5282__bF_buf4), .B(_5713__bF_buf6), .C(_5717_), .Y(_1701_) );
NAND3X1 NAND3X1_554 ( .A(datapath_1_RegisterFile_regfile_mem_12__4_), .B(_5265__bF_buf72), .C(_5713__bF_buf5), .Y(_5718_) );
OAI21X1 OAI21X1_680 ( .A(_5284__bF_buf1), .B(_5713__bF_buf5), .C(_5718_), .Y(_1702_) );
NAND3X1 NAND3X1_555 ( .A(datapath_1_RegisterFile_regfile_mem_12__5_), .B(_5265__bF_buf98), .C(_5713__bF_buf0), .Y(_5719_) );
OAI21X1 OAI21X1_681 ( .A(_5286__bF_buf0), .B(_5713__bF_buf0), .C(_5719_), .Y(_940_) );
NAND3X1 NAND3X1_556 ( .A(datapath_1_RegisterFile_regfile_mem_12__6_), .B(_5265__bF_buf50), .C(_5713__bF_buf4), .Y(_5720_) );
OAI21X1 OAI21X1_682 ( .A(_5288__bF_buf2), .B(_5713__bF_buf4), .C(_5720_), .Y(_941_) );
NAND3X1 NAND3X1_557 ( .A(datapath_1_RegisterFile_regfile_mem_12__7_), .B(_5265__bF_buf57), .C(_5713__bF_buf7), .Y(_5721_) );
OAI21X1 OAI21X1_683 ( .A(_5290__bF_buf4), .B(_5713__bF_buf7), .C(_5721_), .Y(_942_) );
NAND3X1 NAND3X1_558 ( .A(datapath_1_RegisterFile_regfile_mem_12__8_), .B(_5265__bF_buf13), .C(_5713__bF_buf2), .Y(_5722_) );
OAI21X1 OAI21X1_684 ( .A(_5292__bF_buf3), .B(_5713__bF_buf2), .C(_5722_), .Y(_943_) );
NAND3X1 NAND3X1_559 ( .A(datapath_1_RegisterFile_regfile_mem_12__9_), .B(_5265__bF_buf68), .C(_5713__bF_buf3), .Y(_5723_) );
OAI21X1 OAI21X1_685 ( .A(_5294__bF_buf3), .B(_5713__bF_buf3), .C(_5723_), .Y(_944_) );
NAND3X1 NAND3X1_560 ( .A(datapath_1_RegisterFile_regfile_mem_12__10_), .B(_5265__bF_buf74), .C(_5713__bF_buf4), .Y(_5724_) );
OAI21X1 OAI21X1_686 ( .A(_5296__bF_buf4), .B(_5713__bF_buf4), .C(_5724_), .Y(_920_) );
NAND3X1 NAND3X1_561 ( .A(datapath_1_RegisterFile_regfile_mem_12__11_), .B(_5265__bF_buf30), .C(_5713__bF_buf1), .Y(_5725_) );
OAI21X1 OAI21X1_687 ( .A(_5298__bF_buf0), .B(_5713__bF_buf1), .C(_5725_), .Y(_921_) );
NAND3X1 NAND3X1_562 ( .A(datapath_1_RegisterFile_regfile_mem_12__12_), .B(_5265__bF_buf74), .C(_5713__bF_buf4), .Y(_5726_) );
OAI21X1 OAI21X1_688 ( .A(_5300__bF_buf3), .B(_5713__bF_buf4), .C(_5726_), .Y(_1703_) );
NAND3X1 NAND3X1_563 ( .A(datapath_1_RegisterFile_regfile_mem_12__13_), .B(_5265__bF_buf98), .C(_5713__bF_buf0), .Y(_5727_) );
OAI21X1 OAI21X1_689 ( .A(_5302__bF_buf4), .B(_5713__bF_buf0), .C(_5727_), .Y(_922_) );
NAND3X1 NAND3X1_564 ( .A(datapath_1_RegisterFile_regfile_mem_12__14_), .B(_5265__bF_buf87), .C(_5713__bF_buf2), .Y(_5728_) );
OAI21X1 OAI21X1_690 ( .A(_5304__bF_buf1), .B(_5713__bF_buf2), .C(_5728_), .Y(_923_) );
NAND3X1 NAND3X1_565 ( .A(datapath_1_RegisterFile_regfile_mem_12__15_), .B(_5265__bF_buf30), .C(_5713__bF_buf1), .Y(_5729_) );
OAI21X1 OAI21X1_691 ( .A(_5306__bF_buf4), .B(_5713__bF_buf1), .C(_5729_), .Y(_924_) );
NAND3X1 NAND3X1_566 ( .A(datapath_1_RegisterFile_regfile_mem_12__16_), .B(_5265__bF_buf57), .C(_5713__bF_buf7), .Y(_5730_) );
OAI21X1 OAI21X1_692 ( .A(_5308__bF_buf0), .B(_5713__bF_buf7), .C(_5730_), .Y(_925_) );
NAND3X1 NAND3X1_567 ( .A(datapath_1_RegisterFile_regfile_mem_12__17_), .B(_5265__bF_buf51), .C(_5713__bF_buf5), .Y(_5731_) );
OAI21X1 OAI21X1_693 ( .A(_5310__bF_buf4), .B(_5713__bF_buf5), .C(_5731_), .Y(_926_) );
NAND3X1 NAND3X1_568 ( .A(datapath_1_RegisterFile_regfile_mem_12__18_), .B(_5265__bF_buf68), .C(_5713__bF_buf3), .Y(_5732_) );
OAI21X1 OAI21X1_694 ( .A(_5312__bF_buf1), .B(_5713__bF_buf3), .C(_5732_), .Y(_927_) );
NAND3X1 NAND3X1_569 ( .A(datapath_1_RegisterFile_regfile_mem_12__19_), .B(_5265__bF_buf39), .C(_5713__bF_buf1), .Y(_5733_) );
OAI21X1 OAI21X1_695 ( .A(_5314__bF_buf1), .B(_5713__bF_buf1), .C(_5733_), .Y(_928_) );
NAND3X1 NAND3X1_570 ( .A(datapath_1_RegisterFile_regfile_mem_12__20_), .B(_5265__bF_buf26), .C(_5713__bF_buf6), .Y(_5734_) );
OAI21X1 OAI21X1_696 ( .A(_5316__bF_buf2), .B(_5713__bF_buf6), .C(_5734_), .Y(_929_) );
NAND3X1 NAND3X1_571 ( .A(datapath_1_RegisterFile_regfile_mem_12__21_), .B(_5265__bF_buf13), .C(_5713__bF_buf2), .Y(_5735_) );
OAI21X1 OAI21X1_697 ( .A(_5318__bF_buf0), .B(_5713__bF_buf2), .C(_5735_), .Y(_930_) );
NAND3X1 NAND3X1_572 ( .A(datapath_1_RegisterFile_regfile_mem_12__22_), .B(_5265__bF_buf60), .C(_5713__bF_buf0), .Y(_5736_) );
OAI21X1 OAI21X1_698 ( .A(_5320__bF_buf2), .B(_5713__bF_buf0), .C(_5736_), .Y(_1704_) );
NAND3X1 NAND3X1_573 ( .A(datapath_1_RegisterFile_regfile_mem_12__23_), .B(_5265__bF_buf27), .C(_5713__bF_buf3), .Y(_5737_) );
OAI21X1 OAI21X1_699 ( .A(_5322__bF_buf1), .B(_5713__bF_buf3), .C(_5737_), .Y(_931_) );
NAND3X1 NAND3X1_574 ( .A(datapath_1_RegisterFile_regfile_mem_12__24_), .B(_5265__bF_buf76), .C(_5713__bF_buf7), .Y(_5738_) );
OAI21X1 OAI21X1_700 ( .A(_5324__bF_buf0), .B(_5713__bF_buf7), .C(_5738_), .Y(_932_) );
NAND3X1 NAND3X1_575 ( .A(datapath_1_RegisterFile_regfile_mem_12__25_), .B(_5265__bF_buf26), .C(_5713__bF_buf6), .Y(_5739_) );
OAI21X1 OAI21X1_701 ( .A(_5326__bF_buf2), .B(_5713__bF_buf6), .C(_5739_), .Y(_933_) );
NAND3X1 NAND3X1_576 ( .A(datapath_1_RegisterFile_regfile_mem_12__26_), .B(_5265__bF_buf21), .C(_5713__bF_buf0), .Y(_5740_) );
OAI21X1 OAI21X1_702 ( .A(_5328__bF_buf3), .B(_5713__bF_buf0), .C(_5740_), .Y(_934_) );
NAND3X1 NAND3X1_577 ( .A(datapath_1_RegisterFile_regfile_mem_12__27_), .B(_5265__bF_buf42), .C(_5713__bF_buf2), .Y(_5741_) );
OAI21X1 OAI21X1_703 ( .A(_5330__bF_buf3), .B(_5713__bF_buf2), .C(_5741_), .Y(_935_) );
NAND3X1 NAND3X1_578 ( .A(datapath_1_RegisterFile_regfile_mem_12__28_), .B(_5265__bF_buf96), .C(_5713__bF_buf7), .Y(_5742_) );
OAI21X1 OAI21X1_704 ( .A(_5332__bF_buf4), .B(_5713__bF_buf7), .C(_5742_), .Y(_936_) );
NAND3X1 NAND3X1_579 ( .A(datapath_1_RegisterFile_regfile_mem_12__29_), .B(_5265__bF_buf39), .C(_5713__bF_buf1), .Y(_5743_) );
OAI21X1 OAI21X1_705 ( .A(_5334__bF_buf1), .B(_5713__bF_buf1), .C(_5743_), .Y(_937_) );
NAND3X1 NAND3X1_580 ( .A(datapath_1_RegisterFile_regfile_mem_12__30_), .B(_5265__bF_buf72), .C(_5713__bF_buf5), .Y(_5744_) );
OAI21X1 OAI21X1_706 ( .A(_5336__bF_buf2), .B(_5713__bF_buf5), .C(_5744_), .Y(_938_) );
NAND3X1 NAND3X1_581 ( .A(datapath_1_RegisterFile_regfile_mem_12__31_), .B(_5265__bF_buf27), .C(_5713__bF_buf3), .Y(_5745_) );
OAI21X1 OAI21X1_707 ( .A(_5338__bF_buf3), .B(_5713__bF_buf3), .C(_5745_), .Y(_939_) );
NAND2X1 NAND2X1_377 ( .A(_5341_), .B(_5712_), .Y(_5746_) );
NAND3X1 NAND3X1_582 ( .A(datapath_1_RegisterFile_regfile_mem_13__0_), .B(_5265__bF_buf51), .C(_5746__bF_buf7), .Y(_5747_) );
OAI21X1 OAI21X1_708 ( .A(_5276__bF_buf0), .B(_5746__bF_buf7), .C(_5747_), .Y(_945_) );
NAND3X1 NAND3X1_583 ( .A(datapath_1_RegisterFile_regfile_mem_13__1_), .B(_5265__bF_buf74), .C(_5746__bF_buf2), .Y(_5748_) );
OAI21X1 OAI21X1_709 ( .A(_5278__bF_buf2), .B(_5746__bF_buf2), .C(_5748_), .Y(_955_) );
NAND3X1 NAND3X1_584 ( .A(datapath_1_RegisterFile_regfile_mem_13__2_), .B(_5265__bF_buf43), .C(_5746__bF_buf2), .Y(_5749_) );
OAI21X1 OAI21X1_710 ( .A(_5280__bF_buf2), .B(_5746__bF_buf2), .C(_5749_), .Y(_965_) );
NAND3X1 NAND3X1_585 ( .A(datapath_1_RegisterFile_regfile_mem_13__3_), .B(_5265__bF_buf26), .C(_5746__bF_buf1), .Y(_5750_) );
OAI21X1 OAI21X1_711 ( .A(_5282__bF_buf4), .B(_5746__bF_buf1), .C(_5750_), .Y(_966_) );
NAND3X1 NAND3X1_586 ( .A(datapath_1_RegisterFile_regfile_mem_13__4_), .B(_5265__bF_buf74), .C(_5746__bF_buf4), .Y(_5751_) );
OAI21X1 OAI21X1_712 ( .A(_5284__bF_buf4), .B(_5746__bF_buf4), .C(_5751_), .Y(_967_) );
NAND3X1 NAND3X1_587 ( .A(datapath_1_RegisterFile_regfile_mem_13__5_), .B(_5265__bF_buf68), .C(_5746__bF_buf5), .Y(_5752_) );
OAI21X1 OAI21X1_713 ( .A(_5286__bF_buf1), .B(_5746__bF_buf5), .C(_5752_), .Y(_968_) );
NAND3X1 NAND3X1_588 ( .A(datapath_1_RegisterFile_regfile_mem_13__6_), .B(_5265__bF_buf50), .C(_5746__bF_buf1), .Y(_5753_) );
OAI21X1 OAI21X1_714 ( .A(_5288__bF_buf2), .B(_5746__bF_buf1), .C(_5753_), .Y(_969_) );
NAND3X1 NAND3X1_589 ( .A(datapath_1_RegisterFile_regfile_mem_13__7_), .B(_5265__bF_buf62), .C(_5746__bF_buf6), .Y(_5754_) );
OAI21X1 OAI21X1_715 ( .A(_5290__bF_buf1), .B(_5746__bF_buf6), .C(_5754_), .Y(_1705_) );
NAND3X1 NAND3X1_590 ( .A(datapath_1_RegisterFile_regfile_mem_13__8_), .B(_5265__bF_buf92), .C(_5746__bF_buf4), .Y(_5755_) );
OAI21X1 OAI21X1_716 ( .A(_5292__bF_buf1), .B(_5746__bF_buf4), .C(_5755_), .Y(_970_) );
NAND3X1 NAND3X1_591 ( .A(datapath_1_RegisterFile_regfile_mem_13__9_), .B(_5265__bF_buf42), .C(_5746__bF_buf5), .Y(_5756_) );
OAI21X1 OAI21X1_717 ( .A(_5294__bF_buf3), .B(_5746__bF_buf5), .C(_5756_), .Y(_971_) );
NAND3X1 NAND3X1_592 ( .A(datapath_1_RegisterFile_regfile_mem_13__10_), .B(_5265__bF_buf74), .C(_5746__bF_buf2), .Y(_5757_) );
OAI21X1 OAI21X1_718 ( .A(_5296__bF_buf4), .B(_5746__bF_buf2), .C(_5757_), .Y(_946_) );
NAND3X1 NAND3X1_593 ( .A(datapath_1_RegisterFile_regfile_mem_13__11_), .B(_5265__bF_buf30), .C(_5746__bF_buf6), .Y(_5758_) );
OAI21X1 OAI21X1_719 ( .A(_5298__bF_buf3), .B(_5746__bF_buf6), .C(_5758_), .Y(_947_) );
NAND3X1 NAND3X1_594 ( .A(datapath_1_RegisterFile_regfile_mem_13__12_), .B(_5265__bF_buf43), .C(_5746__bF_buf2), .Y(_5759_) );
OAI21X1 OAI21X1_720 ( .A(_5300__bF_buf3), .B(_5746__bF_buf2), .C(_5759_), .Y(_948_) );
NAND3X1 NAND3X1_595 ( .A(datapath_1_RegisterFile_regfile_mem_13__13_), .B(_5265__bF_buf48), .C(_5746__bF_buf3), .Y(_5760_) );
OAI21X1 OAI21X1_721 ( .A(_5302__bF_buf2), .B(_5746__bF_buf3), .C(_5760_), .Y(_949_) );
NAND3X1 NAND3X1_596 ( .A(datapath_1_RegisterFile_regfile_mem_13__14_), .B(_5265__bF_buf6), .C(_5746__bF_buf7), .Y(_5761_) );
OAI21X1 OAI21X1_722 ( .A(_5304__bF_buf0), .B(_5746__bF_buf7), .C(_5761_), .Y(_950_) );
NAND3X1 NAND3X1_597 ( .A(datapath_1_RegisterFile_regfile_mem_13__15_), .B(_5265__bF_buf70), .C(_5746__bF_buf6), .Y(_5762_) );
OAI21X1 OAI21X1_723 ( .A(_5306__bF_buf3), .B(_5746__bF_buf6), .C(_5762_), .Y(_951_) );
NAND3X1 NAND3X1_598 ( .A(datapath_1_RegisterFile_regfile_mem_13__16_), .B(_5265__bF_buf94), .C(_5746__bF_buf0), .Y(_5763_) );
OAI21X1 OAI21X1_724 ( .A(_5308__bF_buf3), .B(_5746__bF_buf0), .C(_5763_), .Y(_952_) );
NAND3X1 NAND3X1_599 ( .A(datapath_1_RegisterFile_regfile_mem_13__17_), .B(_5265__bF_buf51), .C(_5746__bF_buf7), .Y(_5764_) );
OAI21X1 OAI21X1_725 ( .A(_5310__bF_buf4), .B(_5746__bF_buf7), .C(_5764_), .Y(_1706_) );
NAND3X1 NAND3X1_600 ( .A(datapath_1_RegisterFile_regfile_mem_13__18_), .B(_5265__bF_buf68), .C(_5746__bF_buf5), .Y(_5765_) );
OAI21X1 OAI21X1_726 ( .A(_5312__bF_buf1), .B(_5746__bF_buf5), .C(_5765_), .Y(_953_) );
NAND3X1 NAND3X1_601 ( .A(datapath_1_RegisterFile_regfile_mem_13__19_), .B(_5265__bF_buf89), .C(_5746__bF_buf6), .Y(_5766_) );
OAI21X1 OAI21X1_727 ( .A(_5314__bF_buf2), .B(_5746__bF_buf6), .C(_5766_), .Y(_954_) );
NAND3X1 NAND3X1_602 ( .A(datapath_1_RegisterFile_regfile_mem_13__20_), .B(_5265__bF_buf26), .C(_5746__bF_buf1), .Y(_5767_) );
OAI21X1 OAI21X1_728 ( .A(_5316__bF_buf2), .B(_5746__bF_buf1), .C(_5767_), .Y(_956_) );
NAND3X1 NAND3X1_603 ( .A(datapath_1_RegisterFile_regfile_mem_13__21_), .B(_5265__bF_buf92), .C(_5746__bF_buf4), .Y(_5768_) );
OAI21X1 OAI21X1_729 ( .A(_5318__bF_buf4), .B(_5746__bF_buf4), .C(_5768_), .Y(_957_) );
NAND3X1 NAND3X1_604 ( .A(datapath_1_RegisterFile_regfile_mem_13__22_), .B(_5265__bF_buf48), .C(_5746__bF_buf3), .Y(_5769_) );
OAI21X1 OAI21X1_730 ( .A(_5320__bF_buf4), .B(_5746__bF_buf3), .C(_5769_), .Y(_958_) );
NAND3X1 NAND3X1_605 ( .A(datapath_1_RegisterFile_regfile_mem_13__23_), .B(_5265__bF_buf68), .C(_5746__bF_buf5), .Y(_5770_) );
OAI21X1 OAI21X1_731 ( .A(_5322__bF_buf3), .B(_5746__bF_buf5), .C(_5770_), .Y(_959_) );
NAND3X1 NAND3X1_606 ( .A(datapath_1_RegisterFile_regfile_mem_13__24_), .B(_5265__bF_buf86), .C(_5746__bF_buf0), .Y(_5771_) );
OAI21X1 OAI21X1_732 ( .A(_5324__bF_buf3), .B(_5746__bF_buf0), .C(_5771_), .Y(_960_) );
NAND3X1 NAND3X1_607 ( .A(datapath_1_RegisterFile_regfile_mem_13__25_), .B(_5265__bF_buf26), .C(_5746__bF_buf1), .Y(_5772_) );
OAI21X1 OAI21X1_733 ( .A(_5326__bF_buf2), .B(_5746__bF_buf1), .C(_5772_), .Y(_961_) );
NAND3X1 NAND3X1_608 ( .A(datapath_1_RegisterFile_regfile_mem_13__26_), .B(_5265__bF_buf51), .C(_5746__bF_buf3), .Y(_5773_) );
OAI21X1 OAI21X1_734 ( .A(_5328__bF_buf2), .B(_5746__bF_buf3), .C(_5773_), .Y(_962_) );
NAND3X1 NAND3X1_609 ( .A(datapath_1_RegisterFile_regfile_mem_13__27_), .B(_5265__bF_buf6), .C(_5746__bF_buf7), .Y(_5774_) );
OAI21X1 OAI21X1_735 ( .A(_5330__bF_buf3), .B(_5746__bF_buf7), .C(_5774_), .Y(_1707_) );
NAND3X1 NAND3X1_610 ( .A(datapath_1_RegisterFile_regfile_mem_13__28_), .B(_5265__bF_buf86), .C(_5746__bF_buf0), .Y(_5775_) );
OAI21X1 OAI21X1_736 ( .A(_5332__bF_buf1), .B(_5746__bF_buf0), .C(_5775_), .Y(_963_) );
NAND3X1 NAND3X1_611 ( .A(datapath_1_RegisterFile_regfile_mem_13__29_), .B(_5265__bF_buf94), .C(_5746__bF_buf0), .Y(_5776_) );
OAI21X1 OAI21X1_737 ( .A(_5334__bF_buf4), .B(_5746__bF_buf0), .C(_5776_), .Y(_964_) );
NAND3X1 NAND3X1_612 ( .A(datapath_1_RegisterFile_regfile_mem_13__30_), .B(_5265__bF_buf92), .C(_5746__bF_buf4), .Y(_5777_) );
OAI21X1 OAI21X1_738 ( .A(_5336__bF_buf4), .B(_5746__bF_buf4), .C(_5777_), .Y(_1708_) );
NAND3X1 NAND3X1_613 ( .A(datapath_1_RegisterFile_regfile_mem_13__31_), .B(_5265__bF_buf51), .C(_5746__bF_buf3), .Y(_5778_) );
OAI21X1 OAI21X1_739 ( .A(_5338__bF_buf3), .B(_5746__bF_buf3), .C(_5778_), .Y(_1709_) );
NAND2X1 NAND2X1_378 ( .A(_5376_), .B(_5712_), .Y(_5779_) );
NAND3X1 NAND3X1_614 ( .A(datapath_1_RegisterFile_regfile_mem_14__0_), .B(_5265__bF_buf23), .C(_5779__bF_buf2), .Y(_5780_) );
OAI21X1 OAI21X1_740 ( .A(_5276__bF_buf2), .B(_5779__bF_buf2), .C(_5780_), .Y(_972_) );
NAND3X1 NAND3X1_615 ( .A(datapath_1_RegisterFile_regfile_mem_14__1_), .B(_5265__bF_buf91), .C(_5779__bF_buf3), .Y(_5781_) );
OAI21X1 OAI21X1_741 ( .A(_5278__bF_buf0), .B(_5779__bF_buf3), .C(_5781_), .Y(_982_) );
NAND3X1 NAND3X1_616 ( .A(datapath_1_RegisterFile_regfile_mem_14__2_), .B(_5265__bF_buf56), .C(_5779__bF_buf0), .Y(_5782_) );
OAI21X1 OAI21X1_742 ( .A(_5280__bF_buf1), .B(_5779__bF_buf0), .C(_5782_), .Y(_1710_) );
NAND3X1 NAND3X1_617 ( .A(datapath_1_RegisterFile_regfile_mem_14__3_), .B(_5265__bF_buf91), .C(_5779__bF_buf3), .Y(_5783_) );
OAI21X1 OAI21X1_743 ( .A(_5282__bF_buf0), .B(_5779__bF_buf3), .C(_5783_), .Y(_994_) );
NAND3X1 NAND3X1_618 ( .A(datapath_1_RegisterFile_regfile_mem_14__4_), .B(_5265__bF_buf72), .C(_5779__bF_buf7), .Y(_5784_) );
OAI21X1 OAI21X1_744 ( .A(_5284__bF_buf1), .B(_5779__bF_buf7), .C(_5784_), .Y(_995_) );
NAND3X1 NAND3X1_619 ( .A(datapath_1_RegisterFile_regfile_mem_14__5_), .B(_5265__bF_buf48), .C(_5779__bF_buf1), .Y(_5785_) );
OAI21X1 OAI21X1_745 ( .A(_5286__bF_buf0), .B(_5779__bF_buf1), .C(_5785_), .Y(_996_) );
NAND3X1 NAND3X1_620 ( .A(datapath_1_RegisterFile_regfile_mem_14__6_), .B(_5265__bF_buf43), .C(_5779__bF_buf0), .Y(_5786_) );
OAI21X1 OAI21X1_746 ( .A(_5288__bF_buf2), .B(_5779__bF_buf0), .C(_5786_), .Y(_997_) );
NAND3X1 NAND3X1_621 ( .A(datapath_1_RegisterFile_regfile_mem_14__7_), .B(_5265__bF_buf57), .C(_5779__bF_buf4), .Y(_5787_) );
OAI21X1 OAI21X1_747 ( .A(_5290__bF_buf4), .B(_5779__bF_buf4), .C(_5787_), .Y(_998_) );
NAND3X1 NAND3X1_622 ( .A(datapath_1_RegisterFile_regfile_mem_14__8_), .B(_5265__bF_buf74), .C(_5779__bF_buf0), .Y(_5788_) );
OAI21X1 OAI21X1_748 ( .A(_5292__bF_buf3), .B(_5779__bF_buf0), .C(_5788_), .Y(_999_) );
NAND3X1 NAND3X1_623 ( .A(datapath_1_RegisterFile_regfile_mem_14__9_), .B(_5265__bF_buf60), .C(_5779__bF_buf1), .Y(_5789_) );
OAI21X1 OAI21X1_749 ( .A(_5294__bF_buf2), .B(_5779__bF_buf1), .C(_5789_), .Y(_1000_) );
NAND3X1 NAND3X1_624 ( .A(datapath_1_RegisterFile_regfile_mem_14__10_), .B(_5265__bF_buf83), .C(_5779__bF_buf2), .Y(_5790_) );
OAI21X1 OAI21X1_750 ( .A(_5296__bF_buf3), .B(_5779__bF_buf2), .C(_5790_), .Y(_973_) );
NAND3X1 NAND3X1_625 ( .A(datapath_1_RegisterFile_regfile_mem_14__11_), .B(_5265__bF_buf85), .C(_5779__bF_buf6), .Y(_5791_) );
OAI21X1 OAI21X1_751 ( .A(_5298__bF_buf3), .B(_5779__bF_buf6), .C(_5791_), .Y(_974_) );
NAND3X1 NAND3X1_626 ( .A(datapath_1_RegisterFile_regfile_mem_14__12_), .B(_5265__bF_buf74), .C(_5779__bF_buf0), .Y(_5792_) );
OAI21X1 OAI21X1_752 ( .A(_5300__bF_buf3), .B(_5779__bF_buf0), .C(_5792_), .Y(_1711_) );
NAND3X1 NAND3X1_627 ( .A(datapath_1_RegisterFile_regfile_mem_14__13_), .B(_5265__bF_buf77), .C(_5779__bF_buf5), .Y(_5793_) );
OAI21X1 OAI21X1_753 ( .A(_5302__bF_buf4), .B(_5779__bF_buf5), .C(_5793_), .Y(_975_) );
NAND3X1 NAND3X1_628 ( .A(datapath_1_RegisterFile_regfile_mem_14__14_), .B(_5265__bF_buf87), .C(_5779__bF_buf5), .Y(_5794_) );
OAI21X1 OAI21X1_754 ( .A(_5304__bF_buf1), .B(_5779__bF_buf5), .C(_5794_), .Y(_976_) );
NAND3X1 NAND3X1_629 ( .A(datapath_1_RegisterFile_regfile_mem_14__15_), .B(_5265__bF_buf76), .C(_5779__bF_buf4), .Y(_5795_) );
OAI21X1 OAI21X1_755 ( .A(_5306__bF_buf3), .B(_5779__bF_buf4), .C(_5795_), .Y(_977_) );
NAND3X1 NAND3X1_630 ( .A(datapath_1_RegisterFile_regfile_mem_14__16_), .B(_5265__bF_buf76), .C(_5779__bF_buf4), .Y(_5796_) );
OAI21X1 OAI21X1_756 ( .A(_5308__bF_buf0), .B(_5779__bF_buf4), .C(_5796_), .Y(_978_) );
NAND3X1 NAND3X1_631 ( .A(datapath_1_RegisterFile_regfile_mem_14__17_), .B(_5265__bF_buf87), .C(_5779__bF_buf7), .Y(_5797_) );
OAI21X1 OAI21X1_757 ( .A(_5310__bF_buf4), .B(_5779__bF_buf7), .C(_5797_), .Y(_979_) );
NAND3X1 NAND3X1_632 ( .A(datapath_1_RegisterFile_regfile_mem_14__18_), .B(_5265__bF_buf21), .C(_5779__bF_buf1), .Y(_5798_) );
OAI21X1 OAI21X1_758 ( .A(_5312__bF_buf1), .B(_5779__bF_buf1), .C(_5798_), .Y(_980_) );
NAND3X1 NAND3X1_633 ( .A(datapath_1_RegisterFile_regfile_mem_14__19_), .B(_5265__bF_buf84), .C(_5779__bF_buf3), .Y(_5799_) );
OAI21X1 OAI21X1_759 ( .A(_5314__bF_buf3), .B(_5779__bF_buf3), .C(_5799_), .Y(_981_) );
NAND3X1 NAND3X1_634 ( .A(datapath_1_RegisterFile_regfile_mem_14__20_), .B(_5265__bF_buf84), .C(_5779__bF_buf3), .Y(_5800_) );
OAI21X1 OAI21X1_760 ( .A(_5316__bF_buf3), .B(_5779__bF_buf3), .C(_5800_), .Y(_983_) );
NAND3X1 NAND3X1_635 ( .A(datapath_1_RegisterFile_regfile_mem_14__21_), .B(_5265__bF_buf83), .C(_5779__bF_buf2), .Y(_5801_) );
OAI21X1 OAI21X1_761 ( .A(_5318__bF_buf0), .B(_5779__bF_buf2), .C(_5801_), .Y(_984_) );
NAND3X1 NAND3X1_636 ( .A(datapath_1_RegisterFile_regfile_mem_14__22_), .B(_5265__bF_buf60), .C(_5779__bF_buf1), .Y(_5802_) );
OAI21X1 OAI21X1_762 ( .A(_5320__bF_buf2), .B(_5779__bF_buf1), .C(_5802_), .Y(_1712_) );
NAND3X1 NAND3X1_637 ( .A(datapath_1_RegisterFile_regfile_mem_14__23_), .B(_5265__bF_buf27), .C(_5779__bF_buf5), .Y(_5803_) );
OAI21X1 OAI21X1_763 ( .A(_5322__bF_buf1), .B(_5779__bF_buf5), .C(_5803_), .Y(_985_) );
NAND3X1 NAND3X1_638 ( .A(datapath_1_RegisterFile_regfile_mem_14__24_), .B(_5265__bF_buf57), .C(_5779__bF_buf4), .Y(_5804_) );
OAI21X1 OAI21X1_764 ( .A(_5324__bF_buf0), .B(_5779__bF_buf4), .C(_5804_), .Y(_986_) );
NAND3X1 NAND3X1_639 ( .A(datapath_1_RegisterFile_regfile_mem_14__25_), .B(_5265__bF_buf96), .C(_5779__bF_buf6), .Y(_5805_) );
OAI21X1 OAI21X1_765 ( .A(_5326__bF_buf1), .B(_5779__bF_buf6), .C(_5805_), .Y(_987_) );
NAND3X1 NAND3X1_640 ( .A(datapath_1_RegisterFile_regfile_mem_14__26_), .B(_5265__bF_buf64), .C(_5779__bF_buf7), .Y(_5806_) );
OAI21X1 OAI21X1_766 ( .A(_5328__bF_buf2), .B(_5779__bF_buf7), .C(_5806_), .Y(_988_) );
NAND3X1 NAND3X1_641 ( .A(datapath_1_RegisterFile_regfile_mem_14__27_), .B(_5265__bF_buf42), .C(_5779__bF_buf7), .Y(_5807_) );
OAI21X1 OAI21X1_767 ( .A(_5330__bF_buf4), .B(_5779__bF_buf7), .C(_5807_), .Y(_989_) );
NAND3X1 NAND3X1_642 ( .A(datapath_1_RegisterFile_regfile_mem_14__28_), .B(_5265__bF_buf96), .C(_5779__bF_buf6), .Y(_5808_) );
OAI21X1 OAI21X1_768 ( .A(_5332__bF_buf4), .B(_5779__bF_buf6), .C(_5808_), .Y(_990_) );
NAND3X1 NAND3X1_643 ( .A(datapath_1_RegisterFile_regfile_mem_14__29_), .B(_5265__bF_buf84), .C(_5779__bF_buf6), .Y(_5809_) );
OAI21X1 OAI21X1_769 ( .A(_5334__bF_buf4), .B(_5779__bF_buf6), .C(_5809_), .Y(_991_) );
NAND3X1 NAND3X1_644 ( .A(datapath_1_RegisterFile_regfile_mem_14__30_), .B(_5265__bF_buf23), .C(_5779__bF_buf2), .Y(_5810_) );
OAI21X1 OAI21X1_770 ( .A(_5336__bF_buf4), .B(_5779__bF_buf2), .C(_5810_), .Y(_992_) );
NAND3X1 NAND3X1_645 ( .A(datapath_1_RegisterFile_regfile_mem_14__31_), .B(_5265__bF_buf87), .C(_5779__bF_buf5), .Y(_5811_) );
OAI21X1 OAI21X1_771 ( .A(_5338__bF_buf3), .B(_5779__bF_buf5), .C(_5811_), .Y(_993_) );
NAND2X1 NAND2X1_379 ( .A(_5410_), .B(_5712_), .Y(_5812_) );
NAND3X1 NAND3X1_646 ( .A(datapath_1_RegisterFile_regfile_mem_15__0_), .B(_5265__bF_buf13), .C(_5812__bF_buf3), .Y(_5813_) );
OAI21X1 OAI21X1_772 ( .A(_5276__bF_buf2), .B(_5812__bF_buf3), .C(_5813_), .Y(_1713_) );
NAND3X1 NAND3X1_647 ( .A(datapath_1_RegisterFile_regfile_mem_15__1_), .B(_5265__bF_buf56), .C(_5812__bF_buf1), .Y(_5814_) );
OAI21X1 OAI21X1_773 ( .A(_5278__bF_buf0), .B(_5812__bF_buf1), .C(_5814_), .Y(_1714_) );
NAND3X1 NAND3X1_648 ( .A(datapath_1_RegisterFile_regfile_mem_15__2_), .B(_5265__bF_buf0), .C(_5812__bF_buf4), .Y(_5815_) );
OAI21X1 OAI21X1_774 ( .A(_5280__bF_buf2), .B(_5812__bF_buf4), .C(_5815_), .Y(_1715_) );
NAND3X1 NAND3X1_649 ( .A(datapath_1_RegisterFile_regfile_mem_15__3_), .B(_5265__bF_buf91), .C(_5812__bF_buf1), .Y(_5816_) );
OAI21X1 OAI21X1_775 ( .A(_5282__bF_buf0), .B(_5812__bF_buf1), .C(_5816_), .Y(_1716_) );
NAND3X1 NAND3X1_650 ( .A(datapath_1_RegisterFile_regfile_mem_15__4_), .B(_5265__bF_buf13), .C(_5812__bF_buf7), .Y(_5817_) );
OAI21X1 OAI21X1_776 ( .A(_5284__bF_buf4), .B(_5812__bF_buf7), .C(_5817_), .Y(_1717_) );
NAND3X1 NAND3X1_651 ( .A(datapath_1_RegisterFile_regfile_mem_15__5_), .B(_5265__bF_buf27), .C(_5812__bF_buf6), .Y(_5818_) );
OAI21X1 OAI21X1_777 ( .A(_5286__bF_buf1), .B(_5812__bF_buf6), .C(_5818_), .Y(_1718_) );
NAND3X1 NAND3X1_652 ( .A(datapath_1_RegisterFile_regfile_mem_15__6_), .B(_5265__bF_buf0), .C(_5812__bF_buf4), .Y(_5819_) );
OAI21X1 OAI21X1_778 ( .A(_5288__bF_buf2), .B(_5812__bF_buf4), .C(_5819_), .Y(_1719_) );
NAND3X1 NAND3X1_653 ( .A(datapath_1_RegisterFile_regfile_mem_15__7_), .B(_5265__bF_buf76), .C(_5812__bF_buf0), .Y(_5820_) );
OAI21X1 OAI21X1_779 ( .A(_5290__bF_buf1), .B(_5812__bF_buf0), .C(_5820_), .Y(_1720_) );
NAND3X1 NAND3X1_654 ( .A(datapath_1_RegisterFile_regfile_mem_15__8_), .B(_5265__bF_buf0), .C(_5812__bF_buf4), .Y(_5821_) );
OAI21X1 OAI21X1_780 ( .A(_5292__bF_buf3), .B(_5812__bF_buf4), .C(_5821_), .Y(_1721_) );
NAND3X1 NAND3X1_655 ( .A(datapath_1_RegisterFile_regfile_mem_15__9_), .B(_5265__bF_buf27), .C(_5812__bF_buf6), .Y(_5822_) );
OAI21X1 OAI21X1_781 ( .A(_5294__bF_buf3), .B(_5812__bF_buf6), .C(_5822_), .Y(_1722_) );
NAND3X1 NAND3X1_656 ( .A(datapath_1_RegisterFile_regfile_mem_15__10_), .B(_5265__bF_buf13), .C(_5812__bF_buf7), .Y(_5823_) );
OAI21X1 OAI21X1_782 ( .A(_5296__bF_buf4), .B(_5812__bF_buf7), .C(_5823_), .Y(_1001_) );
NAND3X1 NAND3X1_657 ( .A(datapath_1_RegisterFile_regfile_mem_15__11_), .B(_5265__bF_buf76), .C(_5812__bF_buf0), .Y(_5824_) );
OAI21X1 OAI21X1_783 ( .A(_5298__bF_buf3), .B(_5812__bF_buf0), .C(_5824_), .Y(_1002_) );
NAND3X1 NAND3X1_658 ( .A(datapath_1_RegisterFile_regfile_mem_15__12_), .B(_5265__bF_buf0), .C(_5812__bF_buf4), .Y(_5825_) );
OAI21X1 OAI21X1_784 ( .A(_5300__bF_buf3), .B(_5812__bF_buf4), .C(_5825_), .Y(_1003_) );
NAND3X1 NAND3X1_659 ( .A(datapath_1_RegisterFile_regfile_mem_15__13_), .B(_5265__bF_buf21), .C(_5812__bF_buf2), .Y(_5826_) );
OAI21X1 OAI21X1_785 ( .A(_5302__bF_buf4), .B(_5812__bF_buf2), .C(_5826_), .Y(_1004_) );
NAND3X1 NAND3X1_660 ( .A(datapath_1_RegisterFile_regfile_mem_15__14_), .B(_5265__bF_buf87), .C(_5812__bF_buf3), .Y(_5827_) );
OAI21X1 OAI21X1_786 ( .A(_5304__bF_buf1), .B(_5812__bF_buf3), .C(_5827_), .Y(_1005_) );
NAND3X1 NAND3X1_661 ( .A(datapath_1_RegisterFile_regfile_mem_15__15_), .B(_5265__bF_buf57), .C(_5812__bF_buf0), .Y(_5828_) );
OAI21X1 OAI21X1_787 ( .A(_5306__bF_buf3), .B(_5812__bF_buf0), .C(_5828_), .Y(_1006_) );
NAND3X1 NAND3X1_662 ( .A(datapath_1_RegisterFile_regfile_mem_15__16_), .B(_5265__bF_buf84), .C(_5812__bF_buf5), .Y(_5829_) );
OAI21X1 OAI21X1_788 ( .A(_5308__bF_buf2), .B(_5812__bF_buf5), .C(_5829_), .Y(_1007_) );
NAND3X1 NAND3X1_663 ( .A(datapath_1_RegisterFile_regfile_mem_15__17_), .B(_5265__bF_buf87), .C(_5812__bF_buf3), .Y(_5830_) );
OAI21X1 OAI21X1_789 ( .A(_5310__bF_buf4), .B(_5812__bF_buf3), .C(_5830_), .Y(_1723_) );
NAND3X1 NAND3X1_664 ( .A(datapath_1_RegisterFile_regfile_mem_15__18_), .B(_5265__bF_buf98), .C(_5812__bF_buf2), .Y(_5831_) );
OAI21X1 OAI21X1_790 ( .A(_5312__bF_buf0), .B(_5812__bF_buf2), .C(_5831_), .Y(_1008_) );
NAND3X1 NAND3X1_665 ( .A(datapath_1_RegisterFile_regfile_mem_15__19_), .B(_5265__bF_buf35), .C(_5812__bF_buf1), .Y(_5832_) );
OAI21X1 OAI21X1_791 ( .A(_5314__bF_buf3), .B(_5812__bF_buf1), .C(_5832_), .Y(_1009_) );
NAND3X1 NAND3X1_666 ( .A(datapath_1_RegisterFile_regfile_mem_15__20_), .B(_5265__bF_buf84), .C(_5812__bF_buf5), .Y(_5833_) );
OAI21X1 OAI21X1_792 ( .A(_5316__bF_buf3), .B(_5812__bF_buf5), .C(_5833_), .Y(_1010_) );
NAND3X1 NAND3X1_667 ( .A(datapath_1_RegisterFile_regfile_mem_15__21_), .B(_5265__bF_buf13), .C(_5812__bF_buf7), .Y(_5834_) );
OAI21X1 OAI21X1_793 ( .A(_5318__bF_buf0), .B(_5812__bF_buf7), .C(_5834_), .Y(_1011_) );
NAND3X1 NAND3X1_668 ( .A(datapath_1_RegisterFile_regfile_mem_15__22_), .B(_5265__bF_buf98), .C(_5812__bF_buf2), .Y(_5835_) );
OAI21X1 OAI21X1_794 ( .A(_5320__bF_buf2), .B(_5812__bF_buf2), .C(_5835_), .Y(_1012_) );
NAND3X1 NAND3X1_669 ( .A(datapath_1_RegisterFile_regfile_mem_15__23_), .B(_5265__bF_buf68), .C(_5812__bF_buf6), .Y(_5836_) );
OAI21X1 OAI21X1_795 ( .A(_5322__bF_buf1), .B(_5812__bF_buf6), .C(_5836_), .Y(_1013_) );
NAND3X1 NAND3X1_670 ( .A(datapath_1_RegisterFile_regfile_mem_15__24_), .B(_5265__bF_buf76), .C(_5812__bF_buf0), .Y(_5837_) );
OAI21X1 OAI21X1_796 ( .A(_5324__bF_buf0), .B(_5812__bF_buf0), .C(_5837_), .Y(_1014_) );
NAND3X1 NAND3X1_671 ( .A(datapath_1_RegisterFile_regfile_mem_15__25_), .B(_5265__bF_buf35), .C(_5812__bF_buf1), .Y(_5838_) );
OAI21X1 OAI21X1_797 ( .A(_5326__bF_buf1), .B(_5812__bF_buf1), .C(_5838_), .Y(_1015_) );
NAND3X1 NAND3X1_672 ( .A(datapath_1_RegisterFile_regfile_mem_15__26_), .B(_5265__bF_buf51), .C(_5812__bF_buf2), .Y(_5839_) );
OAI21X1 OAI21X1_798 ( .A(_5328__bF_buf3), .B(_5812__bF_buf2), .C(_5839_), .Y(_1016_) );
NAND3X1 NAND3X1_673 ( .A(datapath_1_RegisterFile_regfile_mem_15__27_), .B(_5265__bF_buf42), .C(_5812__bF_buf6), .Y(_5840_) );
OAI21X1 OAI21X1_799 ( .A(_5330__bF_buf4), .B(_5812__bF_buf6), .C(_5840_), .Y(_1724_) );
NAND3X1 NAND3X1_674 ( .A(datapath_1_RegisterFile_regfile_mem_15__28_), .B(_5265__bF_buf85), .C(_5812__bF_buf5), .Y(_5841_) );
OAI21X1 OAI21X1_800 ( .A(_5332__bF_buf4), .B(_5812__bF_buf5), .C(_5841_), .Y(_1017_) );
NAND3X1 NAND3X1_675 ( .A(datapath_1_RegisterFile_regfile_mem_15__29_), .B(_5265__bF_buf85), .C(_5812__bF_buf5), .Y(_5842_) );
OAI21X1 OAI21X1_801 ( .A(_5334__bF_buf4), .B(_5812__bF_buf5), .C(_5842_), .Y(_1018_) );
NAND3X1 NAND3X1_676 ( .A(datapath_1_RegisterFile_regfile_mem_15__30_), .B(_5265__bF_buf13), .C(_5812__bF_buf7), .Y(_5843_) );
OAI21X1 OAI21X1_802 ( .A(_5336__bF_buf4), .B(_5812__bF_buf7), .C(_5843_), .Y(_1019_) );
NAND3X1 NAND3X1_677 ( .A(datapath_1_RegisterFile_regfile_mem_15__31_), .B(_5265__bF_buf87), .C(_5812__bF_buf3), .Y(_5844_) );
OAI21X1 OAI21X1_803 ( .A(_5338__bF_buf3), .B(_5812__bF_buf3), .C(_5844_), .Y(_1020_) );
NAND3X1 NAND3X1_678 ( .A(_5264_), .B(datapath_1_A3_4_), .C(_5272__bF_buf2), .Y(_5845_) );
NOR2X1 NOR2X1_138 ( .A(datapath_1_A3_2_), .B(_5845_), .Y(_5846_) );
NAND2X1 NAND2X1_380 ( .A(_5274_), .B(_5846_), .Y(_5847_) );
NAND3X1 NAND3X1_679 ( .A(datapath_1_RegisterFile_regfile_mem_16__0_), .B(_5265__bF_buf47), .C(_5847__bF_buf0), .Y(_5848_) );
OAI21X1 OAI21X1_804 ( .A(_5276__bF_buf4), .B(_5847__bF_buf0), .C(_5848_), .Y(_1021_) );
NAND3X1 NAND3X1_680 ( .A(datapath_1_RegisterFile_regfile_mem_16__1_), .B(_5265__bF_buf34), .C(_5847__bF_buf3), .Y(_5849_) );
OAI21X1 OAI21X1_805 ( .A(_5278__bF_buf1), .B(_5847__bF_buf3), .C(_5849_), .Y(_1031_) );
NAND3X1 NAND3X1_681 ( .A(datapath_1_RegisterFile_regfile_mem_16__2_), .B(_5265__bF_buf34), .C(_5847__bF_buf3), .Y(_5850_) );
OAI21X1 OAI21X1_806 ( .A(_5280__bF_buf3), .B(_5847__bF_buf1), .C(_5850_), .Y(_1725_) );
NAND3X1 NAND3X1_682 ( .A(datapath_1_RegisterFile_regfile_mem_16__3_), .B(_5265__bF_buf69), .C(_5847__bF_buf1), .Y(_5851_) );
OAI21X1 OAI21X1_807 ( .A(_5282__bF_buf1), .B(_5847__bF_buf1), .C(_5851_), .Y(_1043_) );
NAND3X1 NAND3X1_683 ( .A(datapath_1_RegisterFile_regfile_mem_16__4_), .B(_5265__bF_buf8), .C(_5847__bF_buf7), .Y(_5852_) );
OAI21X1 OAI21X1_808 ( .A(_5284__bF_buf2), .B(_5847__bF_buf7), .C(_5852_), .Y(_1044_) );
NAND3X1 NAND3X1_684 ( .A(datapath_1_RegisterFile_regfile_mem_16__5_), .B(_5265__bF_buf79), .C(_5847__bF_buf2), .Y(_5853_) );
OAI21X1 OAI21X1_809 ( .A(_5286__bF_buf2), .B(_5847__bF_buf2), .C(_5853_), .Y(_1045_) );
NAND3X1 NAND3X1_685 ( .A(datapath_1_RegisterFile_regfile_mem_16__6_), .B(_5265__bF_buf53), .C(_5847__bF_buf4), .Y(_5854_) );
OAI21X1 OAI21X1_810 ( .A(_5288__bF_buf1), .B(_5847__bF_buf4), .C(_5854_), .Y(_1046_) );
NAND3X1 NAND3X1_686 ( .A(datapath_1_RegisterFile_regfile_mem_16__7_), .B(_5265__bF_buf78), .C(_5847__bF_buf1), .Y(_5855_) );
OAI21X1 OAI21X1_811 ( .A(_5290__bF_buf2), .B(_5847__bF_buf5), .C(_5855_), .Y(_1047_) );
NAND3X1 NAND3X1_687 ( .A(datapath_1_RegisterFile_regfile_mem_16__8_), .B(_5265__bF_buf46), .C(_5847__bF_buf7), .Y(_5856_) );
OAI21X1 OAI21X1_812 ( .A(_5292__bF_buf2), .B(_5847__bF_buf7), .C(_5856_), .Y(_1048_) );
NAND3X1 NAND3X1_688 ( .A(datapath_1_RegisterFile_regfile_mem_16__9_), .B(_5265__bF_buf29), .C(_5847__bF_buf6), .Y(_5857_) );
OAI21X1 OAI21X1_813 ( .A(_5294__bF_buf1), .B(_5847__bF_buf6), .C(_5857_), .Y(_1049_) );
NAND3X1 NAND3X1_689 ( .A(datapath_1_RegisterFile_regfile_mem_16__10_), .B(_5265__bF_buf79), .C(_5847__bF_buf2), .Y(_5858_) );
OAI21X1 OAI21X1_814 ( .A(_5296__bF_buf0), .B(_5847__bF_buf2), .C(_5858_), .Y(_1022_) );
NAND3X1 NAND3X1_690 ( .A(datapath_1_RegisterFile_regfile_mem_16__11_), .B(_5265__bF_buf71), .C(_5847__bF_buf5), .Y(_5859_) );
OAI21X1 OAI21X1_815 ( .A(_5298__bF_buf1), .B(_5847__bF_buf5), .C(_5859_), .Y(_1023_) );
NAND3X1 NAND3X1_691 ( .A(datapath_1_RegisterFile_regfile_mem_16__12_), .B(_5265__bF_buf20), .C(_5847__bF_buf1), .Y(_5860_) );
OAI21X1 OAI21X1_816 ( .A(_5300__bF_buf0), .B(_5847__bF_buf1), .C(_5860_), .Y(_1726_) );
NAND3X1 NAND3X1_692 ( .A(datapath_1_RegisterFile_regfile_mem_16__13_), .B(_5265__bF_buf79), .C(_5847__bF_buf2), .Y(_5861_) );
OAI21X1 OAI21X1_817 ( .A(_5302__bF_buf1), .B(_5847__bF_buf2), .C(_5861_), .Y(_1024_) );
NAND3X1 NAND3X1_693 ( .A(datapath_1_RegisterFile_regfile_mem_16__14_), .B(_5265__bF_buf81), .C(_5847__bF_buf6), .Y(_5862_) );
OAI21X1 OAI21X1_818 ( .A(_5304__bF_buf2), .B(_5847__bF_buf6), .C(_5862_), .Y(_1025_) );
NAND3X1 NAND3X1_694 ( .A(datapath_1_RegisterFile_regfile_mem_16__15_), .B(_5265__bF_buf32), .C(_5847__bF_buf5), .Y(_5863_) );
OAI21X1 OAI21X1_819 ( .A(_5306__bF_buf2), .B(_5847__bF_buf5), .C(_5863_), .Y(_1026_) );
NAND3X1 NAND3X1_695 ( .A(datapath_1_RegisterFile_regfile_mem_16__16_), .B(_5265__bF_buf24), .C(_5847__bF_buf4), .Y(_5864_) );
OAI21X1 OAI21X1_820 ( .A(_5308__bF_buf1), .B(_5847__bF_buf4), .C(_5864_), .Y(_1027_) );
NAND3X1 NAND3X1_696 ( .A(datapath_1_RegisterFile_regfile_mem_16__17_), .B(_5265__bF_buf8), .C(_5847__bF_buf7), .Y(_5865_) );
OAI21X1 OAI21X1_821 ( .A(_5310__bF_buf3), .B(_5847__bF_buf7), .C(_5865_), .Y(_1028_) );
NAND3X1 NAND3X1_697 ( .A(datapath_1_RegisterFile_regfile_mem_16__18_), .B(_5265__bF_buf58), .C(_5847__bF_buf2), .Y(_5866_) );
OAI21X1 OAI21X1_822 ( .A(_5312__bF_buf4), .B(_5847__bF_buf2), .C(_5866_), .Y(_1029_) );
NAND3X1 NAND3X1_698 ( .A(datapath_1_RegisterFile_regfile_mem_16__19_), .B(_5265__bF_buf71), .C(_5847__bF_buf5), .Y(_5867_) );
OAI21X1 OAI21X1_823 ( .A(_5314__bF_buf4), .B(_5847__bF_buf5), .C(_5867_), .Y(_1030_) );
NAND3X1 NAND3X1_699 ( .A(datapath_1_RegisterFile_regfile_mem_16__20_), .B(_5265__bF_buf88), .C(_5847__bF_buf1), .Y(_5868_) );
OAI21X1 OAI21X1_824 ( .A(_5316__bF_buf4), .B(_5847__bF_buf1), .C(_5868_), .Y(_1032_) );
NAND3X1 NAND3X1_700 ( .A(datapath_1_RegisterFile_regfile_mem_16__21_), .B(_5265__bF_buf46), .C(_5847__bF_buf7), .Y(_5869_) );
OAI21X1 OAI21X1_825 ( .A(_5318__bF_buf1), .B(_5847__bF_buf7), .C(_5869_), .Y(_1033_) );
NAND3X1 NAND3X1_701 ( .A(datapath_1_RegisterFile_regfile_mem_16__22_), .B(_5265__bF_buf66), .C(_5847__bF_buf0), .Y(_5870_) );
OAI21X1 OAI21X1_826 ( .A(_5320__bF_buf1), .B(_5847__bF_buf0), .C(_5870_), .Y(_1727_) );
NAND3X1 NAND3X1_702 ( .A(datapath_1_RegisterFile_regfile_mem_16__23_), .B(_5265__bF_buf53), .C(_5847__bF_buf4), .Y(_5871_) );
OAI21X1 OAI21X1_827 ( .A(_5322__bF_buf4), .B(_5847__bF_buf4), .C(_5871_), .Y(_1034_) );
NAND3X1 NAND3X1_703 ( .A(datapath_1_RegisterFile_regfile_mem_16__24_), .B(_5265__bF_buf32), .C(_5847__bF_buf3), .Y(_5872_) );
OAI21X1 OAI21X1_828 ( .A(_5324__bF_buf2), .B(_5847__bF_buf3), .C(_5872_), .Y(_1035_) );
NAND3X1 NAND3X1_704 ( .A(datapath_1_RegisterFile_regfile_mem_16__25_), .B(_5265__bF_buf34), .C(_5847__bF_buf3), .Y(_5873_) );
OAI21X1 OAI21X1_829 ( .A(_5326__bF_buf4), .B(_5847__bF_buf3), .C(_5873_), .Y(_1036_) );
NAND3X1 NAND3X1_705 ( .A(datapath_1_RegisterFile_regfile_mem_16__26_), .B(_5265__bF_buf47), .C(_5847__bF_buf0), .Y(_5874_) );
OAI21X1 OAI21X1_830 ( .A(_5328__bF_buf1), .B(_5847__bF_buf0), .C(_5874_), .Y(_1037_) );
NAND3X1 NAND3X1_706 ( .A(datapath_1_RegisterFile_regfile_mem_16__27_), .B(_5265__bF_buf29), .C(_5847__bF_buf6), .Y(_5875_) );
OAI21X1 OAI21X1_831 ( .A(_5330__bF_buf2), .B(_5847__bF_buf6), .C(_5875_), .Y(_1038_) );
NAND3X1 NAND3X1_707 ( .A(datapath_1_RegisterFile_regfile_mem_16__28_), .B(_5265__bF_buf11), .C(_5847__bF_buf5), .Y(_5876_) );
OAI21X1 OAI21X1_832 ( .A(_5332__bF_buf2), .B(_5847__bF_buf3), .C(_5876_), .Y(_1039_) );
NAND3X1 NAND3X1_708 ( .A(datapath_1_RegisterFile_regfile_mem_16__29_), .B(_5265__bF_buf80), .C(_5847__bF_buf4), .Y(_5877_) );
OAI21X1 OAI21X1_833 ( .A(_5334__bF_buf0), .B(_5847__bF_buf4), .C(_5877_), .Y(_1040_) );
NAND3X1 NAND3X1_709 ( .A(datapath_1_RegisterFile_regfile_mem_16__30_), .B(_5265__bF_buf66), .C(_5847__bF_buf0), .Y(_5878_) );
OAI21X1 OAI21X1_834 ( .A(_5336__bF_buf3), .B(_5847__bF_buf0), .C(_5878_), .Y(_1041_) );
NAND3X1 NAND3X1_710 ( .A(datapath_1_RegisterFile_regfile_mem_16__31_), .B(_5265__bF_buf81), .C(_5847__bF_buf6), .Y(_5879_) );
OAI21X1 OAI21X1_835 ( .A(_5338__bF_buf2), .B(_5847__bF_buf6), .C(_5879_), .Y(_1042_) );
NAND2X1 NAND2X1_381 ( .A(_5341_), .B(_5846_), .Y(_5880_) );
NAND3X1 NAND3X1_711 ( .A(datapath_1_RegisterFile_regfile_mem_17__0_), .B(_5265__bF_buf47), .C(_5880__bF_buf5), .Y(_5881_) );
OAI21X1 OAI21X1_836 ( .A(_5276__bF_buf4), .B(_5880__bF_buf5), .C(_5881_), .Y(_1050_) );
NAND3X1 NAND3X1_712 ( .A(datapath_1_RegisterFile_regfile_mem_17__1_), .B(_5265__bF_buf16), .C(_5880__bF_buf1), .Y(_5882_) );
OAI21X1 OAI21X1_837 ( .A(_5278__bF_buf1), .B(_5880__bF_buf1), .C(_5882_), .Y(_1060_) );
NAND3X1 NAND3X1_713 ( .A(datapath_1_RegisterFile_regfile_mem_17__2_), .B(_5265__bF_buf16), .C(_5880__bF_buf1), .Y(_5883_) );
OAI21X1 OAI21X1_838 ( .A(_5280__bF_buf3), .B(_5880__bF_buf1), .C(_5883_), .Y(_1070_) );
NAND3X1 NAND3X1_714 ( .A(datapath_1_RegisterFile_regfile_mem_17__3_), .B(_5265__bF_buf14), .C(_5880__bF_buf2), .Y(_5884_) );
OAI21X1 OAI21X1_839 ( .A(_5282__bF_buf1), .B(_5880__bF_buf2), .C(_5884_), .Y(_1073_) );
NAND3X1 NAND3X1_715 ( .A(datapath_1_RegisterFile_regfile_mem_17__4_), .B(_5265__bF_buf49), .C(_5880__bF_buf0), .Y(_5885_) );
OAI21X1 OAI21X1_840 ( .A(_5284__bF_buf0), .B(_5880__bF_buf0), .C(_5885_), .Y(_1074_) );
NAND3X1 NAND3X1_716 ( .A(datapath_1_RegisterFile_regfile_mem_17__5_), .B(_5265__bF_buf29), .C(_5880__bF_buf3), .Y(_5886_) );
OAI21X1 OAI21X1_841 ( .A(_5286__bF_buf3), .B(_5880__bF_buf3), .C(_5886_), .Y(_1075_) );
NAND3X1 NAND3X1_717 ( .A(datapath_1_RegisterFile_regfile_mem_17__6_), .B(_5265__bF_buf67), .C(_5880__bF_buf4), .Y(_5887_) );
OAI21X1 OAI21X1_842 ( .A(_5288__bF_buf1), .B(_5880__bF_buf4), .C(_5887_), .Y(_1076_) );
NAND3X1 NAND3X1_718 ( .A(datapath_1_RegisterFile_regfile_mem_17__7_), .B(_5265__bF_buf11), .C(_5880__bF_buf7), .Y(_5888_) );
OAI21X1 OAI21X1_843 ( .A(_5290__bF_buf2), .B(_5880__bF_buf7), .C(_5888_), .Y(_1728_) );
NAND3X1 NAND3X1_719 ( .A(datapath_1_RegisterFile_regfile_mem_17__8_), .B(_5265__bF_buf67), .C(_5880__bF_buf0), .Y(_5889_) );
OAI21X1 OAI21X1_844 ( .A(_5292__bF_buf0), .B(_5880__bF_buf0), .C(_5889_), .Y(_1077_) );
NAND3X1 NAND3X1_720 ( .A(datapath_1_RegisterFile_regfile_mem_17__9_), .B(_5265__bF_buf81), .C(_5880__bF_buf6), .Y(_5890_) );
OAI21X1 OAI21X1_845 ( .A(_5294__bF_buf1), .B(_5880__bF_buf6), .C(_5890_), .Y(_1078_) );
NAND3X1 NAND3X1_721 ( .A(datapath_1_RegisterFile_regfile_mem_17__10_), .B(_5265__bF_buf79), .C(_5880__bF_buf3), .Y(_5891_) );
OAI21X1 OAI21X1_846 ( .A(_5296__bF_buf0), .B(_5880__bF_buf3), .C(_5891_), .Y(_1051_) );
NAND3X1 NAND3X1_722 ( .A(datapath_1_RegisterFile_regfile_mem_17__11_), .B(_5265__bF_buf78), .C(_5880__bF_buf2), .Y(_5892_) );
OAI21X1 OAI21X1_847 ( .A(_5298__bF_buf1), .B(_5880__bF_buf2), .C(_5892_), .Y(_1052_) );
NAND3X1 NAND3X1_723 ( .A(datapath_1_RegisterFile_regfile_mem_17__12_), .B(_5265__bF_buf40), .C(_5880__bF_buf4), .Y(_5893_) );
OAI21X1 OAI21X1_848 ( .A(_5300__bF_buf2), .B(_5880__bF_buf4), .C(_5893_), .Y(_1053_) );
NAND3X1 NAND3X1_724 ( .A(datapath_1_RegisterFile_regfile_mem_17__13_), .B(_5265__bF_buf29), .C(_5880__bF_buf3), .Y(_5894_) );
OAI21X1 OAI21X1_849 ( .A(_5302__bF_buf1), .B(_5880__bF_buf3), .C(_5894_), .Y(_1054_) );
NAND3X1 NAND3X1_725 ( .A(datapath_1_RegisterFile_regfile_mem_17__14_), .B(_5265__bF_buf81), .C(_5880__bF_buf6), .Y(_5895_) );
OAI21X1 OAI21X1_850 ( .A(_5304__bF_buf2), .B(_5880__bF_buf6), .C(_5895_), .Y(_1055_) );
NAND3X1 NAND3X1_726 ( .A(datapath_1_RegisterFile_regfile_mem_17__15_), .B(_5265__bF_buf32), .C(_5880__bF_buf7), .Y(_5896_) );
OAI21X1 OAI21X1_851 ( .A(_5306__bF_buf2), .B(_5880__bF_buf7), .C(_5896_), .Y(_1056_) );
NAND3X1 NAND3X1_727 ( .A(datapath_1_RegisterFile_regfile_mem_17__16_), .B(_5265__bF_buf24), .C(_5880__bF_buf4), .Y(_5897_) );
OAI21X1 OAI21X1_852 ( .A(_5308__bF_buf1), .B(_5880__bF_buf4), .C(_5897_), .Y(_1057_) );
NAND3X1 NAND3X1_728 ( .A(datapath_1_RegisterFile_regfile_mem_17__17_), .B(_5265__bF_buf8), .C(_5880__bF_buf0), .Y(_5898_) );
OAI21X1 OAI21X1_853 ( .A(_5310__bF_buf0), .B(_5880__bF_buf0), .C(_5898_), .Y(_1729_) );
NAND3X1 NAND3X1_729 ( .A(datapath_1_RegisterFile_regfile_mem_17__18_), .B(_5265__bF_buf58), .C(_5880__bF_buf3), .Y(_5899_) );
OAI21X1 OAI21X1_854 ( .A(_5312__bF_buf2), .B(_5880__bF_buf3), .C(_5899_), .Y(_1058_) );
NAND3X1 NAND3X1_730 ( .A(datapath_1_RegisterFile_regfile_mem_17__19_), .B(_5265__bF_buf78), .C(_5880__bF_buf2), .Y(_5900_) );
OAI21X1 OAI21X1_855 ( .A(_5314__bF_buf4), .B(_5880__bF_buf2), .C(_5900_), .Y(_1059_) );
NAND3X1 NAND3X1_731 ( .A(datapath_1_RegisterFile_regfile_mem_17__20_), .B(_5265__bF_buf88), .C(_5880__bF_buf2), .Y(_5901_) );
OAI21X1 OAI21X1_856 ( .A(_5316__bF_buf4), .B(_5880__bF_buf2), .C(_5901_), .Y(_1061_) );
NAND3X1 NAND3X1_732 ( .A(datapath_1_RegisterFile_regfile_mem_17__21_), .B(_5265__bF_buf54), .C(_5880__bF_buf0), .Y(_5902_) );
OAI21X1 OAI21X1_857 ( .A(_5318__bF_buf1), .B(_5880__bF_buf0), .C(_5902_), .Y(_1062_) );
NAND3X1 NAND3X1_733 ( .A(datapath_1_RegisterFile_regfile_mem_17__22_), .B(_5265__bF_buf66), .C(_5880__bF_buf5), .Y(_5903_) );
OAI21X1 OAI21X1_858 ( .A(_5320__bF_buf1), .B(_5880__bF_buf5), .C(_5903_), .Y(_1063_) );
NAND3X1 NAND3X1_734 ( .A(datapath_1_RegisterFile_regfile_mem_17__23_), .B(_5265__bF_buf95), .C(_5880__bF_buf4), .Y(_5904_) );
OAI21X1 OAI21X1_859 ( .A(_5322__bF_buf4), .B(_5880__bF_buf4), .C(_5904_), .Y(_1064_) );
NAND3X1 NAND3X1_735 ( .A(datapath_1_RegisterFile_regfile_mem_17__24_), .B(_5265__bF_buf16), .C(_5880__bF_buf1), .Y(_5905_) );
OAI21X1 OAI21X1_860 ( .A(_5324__bF_buf2), .B(_5880__bF_buf1), .C(_5905_), .Y(_1065_) );
NAND3X1 NAND3X1_736 ( .A(datapath_1_RegisterFile_regfile_mem_17__25_), .B(_5265__bF_buf34), .C(_5880__bF_buf7), .Y(_5906_) );
OAI21X1 OAI21X1_861 ( .A(_5326__bF_buf4), .B(_5880__bF_buf7), .C(_5906_), .Y(_1066_) );
NAND3X1 NAND3X1_737 ( .A(datapath_1_RegisterFile_regfile_mem_17__26_), .B(_5265__bF_buf47), .C(_5880__bF_buf5), .Y(_5907_) );
OAI21X1 OAI21X1_862 ( .A(_5328__bF_buf1), .B(_5880__bF_buf5), .C(_5907_), .Y(_1067_) );
NAND3X1 NAND3X1_738 ( .A(datapath_1_RegisterFile_regfile_mem_17__27_), .B(_5265__bF_buf81), .C(_5880__bF_buf6), .Y(_5908_) );
OAI21X1 OAI21X1_863 ( .A(_5330__bF_buf2), .B(_5880__bF_buf6), .C(_5908_), .Y(_1730_) );
NAND3X1 NAND3X1_739 ( .A(datapath_1_RegisterFile_regfile_mem_17__28_), .B(_5265__bF_buf11), .C(_5880__bF_buf7), .Y(_5909_) );
OAI21X1 OAI21X1_864 ( .A(_5332__bF_buf2), .B(_5880__bF_buf7), .C(_5909_), .Y(_1068_) );
NAND3X1 NAND3X1_740 ( .A(datapath_1_RegisterFile_regfile_mem_17__29_), .B(_5265__bF_buf16), .C(_5880__bF_buf1), .Y(_5910_) );
OAI21X1 OAI21X1_865 ( .A(_5334__bF_buf3), .B(_5880__bF_buf1), .C(_5910_), .Y(_1069_) );
NAND3X1 NAND3X1_741 ( .A(datapath_1_RegisterFile_regfile_mem_17__30_), .B(_5265__bF_buf66), .C(_5880__bF_buf5), .Y(_5911_) );
OAI21X1 OAI21X1_866 ( .A(_5336__bF_buf3), .B(_5880__bF_buf5), .C(_5911_), .Y(_1071_) );
NAND3X1 NAND3X1_742 ( .A(datapath_1_RegisterFile_regfile_mem_17__31_), .B(_5265__bF_buf81), .C(_5880__bF_buf6), .Y(_5912_) );
OAI21X1 OAI21X1_867 ( .A(_5338__bF_buf2), .B(_5880__bF_buf6), .C(_5912_), .Y(_1072_) );
NAND2X1 NAND2X1_382 ( .A(_5376_), .B(_5846_), .Y(_5913_) );
NAND3X1 NAND3X1_743 ( .A(datapath_1_RegisterFile_regfile_mem_18__0_), .B(_5265__bF_buf1), .C(_5913__bF_buf7), .Y(_5914_) );
OAI21X1 OAI21X1_868 ( .A(_5276__bF_buf4), .B(_5913__bF_buf7), .C(_5914_), .Y(_1079_) );
NAND3X1 NAND3X1_744 ( .A(datapath_1_RegisterFile_regfile_mem_18__1_), .B(_5265__bF_buf32), .C(_5913__bF_buf1), .Y(_5915_) );
OAI21X1 OAI21X1_869 ( .A(_5278__bF_buf1), .B(_5913__bF_buf1), .C(_5915_), .Y(_1085_) );
NAND3X1 NAND3X1_745 ( .A(datapath_1_RegisterFile_regfile_mem_18__2_), .B(_5265__bF_buf32), .C(_5913__bF_buf1), .Y(_5916_) );
OAI21X1 OAI21X1_870 ( .A(_5280__bF_buf3), .B(_5913__bF_buf1), .C(_5916_), .Y(_1731_) );
NAND3X1 NAND3X1_746 ( .A(datapath_1_RegisterFile_regfile_mem_18__3_), .B(_5265__bF_buf14), .C(_5913__bF_buf5), .Y(_5917_) );
OAI21X1 OAI21X1_871 ( .A(_5282__bF_buf1), .B(_5913__bF_buf5), .C(_5917_), .Y(_1097_) );
NAND3X1 NAND3X1_747 ( .A(datapath_1_RegisterFile_regfile_mem_18__4_), .B(_5265__bF_buf49), .C(_5913__bF_buf4), .Y(_5918_) );
OAI21X1 OAI21X1_872 ( .A(_5284__bF_buf0), .B(_5913__bF_buf4), .C(_5918_), .Y(_1098_) );
NAND3X1 NAND3X1_748 ( .A(datapath_1_RegisterFile_regfile_mem_18__5_), .B(_5265__bF_buf37), .C(_5913__bF_buf3), .Y(_5919_) );
OAI21X1 OAI21X1_873 ( .A(_5286__bF_buf3), .B(_5913__bF_buf3), .C(_5919_), .Y(_1732_) );
NAND3X1 NAND3X1_749 ( .A(datapath_1_RegisterFile_regfile_mem_18__6_), .B(_5265__bF_buf95), .C(_5913__bF_buf6), .Y(_5920_) );
OAI21X1 OAI21X1_874 ( .A(_5288__bF_buf1), .B(_5913__bF_buf6), .C(_5920_), .Y(_1733_) );
NAND3X1 NAND3X1_750 ( .A(datapath_1_RegisterFile_regfile_mem_18__7_), .B(_5265__bF_buf88), .C(_5913__bF_buf5), .Y(_5921_) );
OAI21X1 OAI21X1_875 ( .A(_5290__bF_buf2), .B(_5913__bF_buf5), .C(_5921_), .Y(_1734_) );
NAND3X1 NAND3X1_751 ( .A(datapath_1_RegisterFile_regfile_mem_18__8_), .B(_5265__bF_buf54), .C(_5913__bF_buf4), .Y(_5922_) );
OAI21X1 OAI21X1_876 ( .A(_5292__bF_buf0), .B(_5913__bF_buf4), .C(_5922_), .Y(_1735_) );
NAND3X1 NAND3X1_752 ( .A(datapath_1_RegisterFile_regfile_mem_18__9_), .B(_5265__bF_buf29), .C(_5913__bF_buf3), .Y(_5923_) );
OAI21X1 OAI21X1_877 ( .A(_5294__bF_buf1), .B(_5913__bF_buf3), .C(_5923_), .Y(_1736_) );
NAND3X1 NAND3X1_753 ( .A(datapath_1_RegisterFile_regfile_mem_18__10_), .B(_5265__bF_buf15), .C(_5913__bF_buf2), .Y(_5924_) );
OAI21X1 OAI21X1_878 ( .A(_5296__bF_buf0), .B(_5913__bF_buf2), .C(_5924_), .Y(_1737_) );
NAND3X1 NAND3X1_754 ( .A(datapath_1_RegisterFile_regfile_mem_18__11_), .B(_5265__bF_buf71), .C(_5913__bF_buf0), .Y(_5925_) );
OAI21X1 OAI21X1_879 ( .A(_5298__bF_buf1), .B(_5913__bF_buf0), .C(_5925_), .Y(_1738_) );
NAND3X1 NAND3X1_755 ( .A(datapath_1_RegisterFile_regfile_mem_18__12_), .B(_5265__bF_buf20), .C(_5913__bF_buf5), .Y(_5926_) );
OAI21X1 OAI21X1_880 ( .A(_5300__bF_buf0), .B(_5913__bF_buf5), .C(_5926_), .Y(_1739_) );
NAND3X1 NAND3X1_756 ( .A(datapath_1_RegisterFile_regfile_mem_18__13_), .B(_5265__bF_buf17), .C(_5913__bF_buf2), .Y(_5927_) );
OAI21X1 OAI21X1_881 ( .A(_5302__bF_buf1), .B(_5913__bF_buf2), .C(_5927_), .Y(_1740_) );
NAND3X1 NAND3X1_757 ( .A(datapath_1_RegisterFile_regfile_mem_18__14_), .B(_5265__bF_buf81), .C(_5913__bF_buf2), .Y(_5928_) );
OAI21X1 OAI21X1_882 ( .A(_5304__bF_buf2), .B(_5913__bF_buf2), .C(_5928_), .Y(_1741_) );
NAND3X1 NAND3X1_758 ( .A(datapath_1_RegisterFile_regfile_mem_18__15_), .B(_5265__bF_buf32), .C(_5913__bF_buf1), .Y(_5929_) );
OAI21X1 OAI21X1_883 ( .A(_5306__bF_buf2), .B(_5913__bF_buf1), .C(_5929_), .Y(_1080_) );
NAND3X1 NAND3X1_759 ( .A(datapath_1_RegisterFile_regfile_mem_18__16_), .B(_5265__bF_buf80), .C(_5913__bF_buf6), .Y(_5930_) );
OAI21X1 OAI21X1_884 ( .A(_5308__bF_buf4), .B(_5913__bF_buf6), .C(_5930_), .Y(_1081_) );
NAND3X1 NAND3X1_760 ( .A(datapath_1_RegisterFile_regfile_mem_18__17_), .B(_5265__bF_buf8), .C(_5913__bF_buf4), .Y(_5931_) );
OAI21X1 OAI21X1_885 ( .A(_5310__bF_buf0), .B(_5913__bF_buf4), .C(_5931_), .Y(_1082_) );
NAND3X1 NAND3X1_761 ( .A(datapath_1_RegisterFile_regfile_mem_18__18_), .B(_5265__bF_buf37), .C(_5913__bF_buf3), .Y(_5932_) );
OAI21X1 OAI21X1_886 ( .A(_5312__bF_buf4), .B(_5913__bF_buf3), .C(_5932_), .Y(_1083_) );
NAND3X1 NAND3X1_762 ( .A(datapath_1_RegisterFile_regfile_mem_18__19_), .B(_5265__bF_buf78), .C(_5913__bF_buf0), .Y(_5933_) );
OAI21X1 OAI21X1_887 ( .A(_5314__bF_buf4), .B(_5913__bF_buf0), .C(_5933_), .Y(_1084_) );
NAND3X1 NAND3X1_763 ( .A(datapath_1_RegisterFile_regfile_mem_18__20_), .B(_5265__bF_buf88), .C(_5913__bF_buf5), .Y(_5934_) );
OAI21X1 OAI21X1_888 ( .A(_5316__bF_buf4), .B(_5913__bF_buf5), .C(_5934_), .Y(_1086_) );
NAND3X1 NAND3X1_764 ( .A(datapath_1_RegisterFile_regfile_mem_18__21_), .B(_5265__bF_buf54), .C(_5913__bF_buf4), .Y(_5935_) );
OAI21X1 OAI21X1_889 ( .A(_5318__bF_buf1), .B(_5913__bF_buf4), .C(_5935_), .Y(_1087_) );
NAND3X1 NAND3X1_765 ( .A(datapath_1_RegisterFile_regfile_mem_18__22_), .B(_5265__bF_buf82), .C(_5913__bF_buf7), .Y(_5936_) );
OAI21X1 OAI21X1_890 ( .A(_5320__bF_buf1), .B(_5913__bF_buf7), .C(_5936_), .Y(_1742_) );
NAND3X1 NAND3X1_766 ( .A(datapath_1_RegisterFile_regfile_mem_18__23_), .B(_5265__bF_buf95), .C(_5913__bF_buf6), .Y(_5937_) );
OAI21X1 OAI21X1_891 ( .A(_5322__bF_buf4), .B(_5913__bF_buf6), .C(_5937_), .Y(_1088_) );
NAND3X1 NAND3X1_767 ( .A(datapath_1_RegisterFile_regfile_mem_18__24_), .B(_5265__bF_buf32), .C(_5913__bF_buf1), .Y(_5938_) );
OAI21X1 OAI21X1_892 ( .A(_5324__bF_buf2), .B(_5913__bF_buf1), .C(_5938_), .Y(_1089_) );
NAND3X1 NAND3X1_768 ( .A(datapath_1_RegisterFile_regfile_mem_18__25_), .B(_5265__bF_buf32), .C(_5913__bF_buf0), .Y(_5939_) );
OAI21X1 OAI21X1_893 ( .A(_5326__bF_buf4), .B(_5913__bF_buf0), .C(_5939_), .Y(_1090_) );
NAND3X1 NAND3X1_769 ( .A(datapath_1_RegisterFile_regfile_mem_18__26_), .B(_5265__bF_buf1), .C(_5913__bF_buf7), .Y(_5940_) );
OAI21X1 OAI21X1_894 ( .A(_5328__bF_buf4), .B(_5913__bF_buf7), .C(_5940_), .Y(_1091_) );
NAND3X1 NAND3X1_770 ( .A(datapath_1_RegisterFile_regfile_mem_18__27_), .B(_5265__bF_buf29), .C(_5913__bF_buf3), .Y(_5941_) );
OAI21X1 OAI21X1_895 ( .A(_5330__bF_buf2), .B(_5913__bF_buf3), .C(_5941_), .Y(_1092_) );
NAND3X1 NAND3X1_771 ( .A(datapath_1_RegisterFile_regfile_mem_18__28_), .B(_5265__bF_buf32), .C(_5913__bF_buf0), .Y(_5942_) );
OAI21X1 OAI21X1_896 ( .A(_5332__bF_buf2), .B(_5913__bF_buf0), .C(_5942_), .Y(_1093_) );
NAND3X1 NAND3X1_772 ( .A(datapath_1_RegisterFile_regfile_mem_18__29_), .B(_5265__bF_buf80), .C(_5913__bF_buf6), .Y(_5943_) );
OAI21X1 OAI21X1_897 ( .A(_5334__bF_buf0), .B(_5913__bF_buf6), .C(_5943_), .Y(_1094_) );
NAND3X1 NAND3X1_773 ( .A(datapath_1_RegisterFile_regfile_mem_18__30_), .B(_5265__bF_buf82), .C(_5913__bF_buf7), .Y(_5944_) );
OAI21X1 OAI21X1_898 ( .A(_5336__bF_buf1), .B(_5913__bF_buf7), .C(_5944_), .Y(_1095_) );
NAND3X1 NAND3X1_774 ( .A(datapath_1_RegisterFile_regfile_mem_18__31_), .B(_5265__bF_buf17), .C(_5913__bF_buf2), .Y(_5945_) );
OAI21X1 OAI21X1_899 ( .A(_5338__bF_buf2), .B(_5913__bF_buf2), .C(_5945_), .Y(_1096_) );
NAND2X1 NAND2X1_383 ( .A(_5410_), .B(_5846_), .Y(_5946_) );
NAND3X1 NAND3X1_775 ( .A(datapath_1_RegisterFile_regfile_mem_19__0_), .B(_5265__bF_buf47), .C(_5946__bF_buf7), .Y(_5947_) );
OAI21X1 OAI21X1_900 ( .A(_5276__bF_buf4), .B(_5946__bF_buf7), .C(_5947_), .Y(_1099_) );
NAND3X1 NAND3X1_776 ( .A(datapath_1_RegisterFile_regfile_mem_19__1_), .B(_5265__bF_buf34), .C(_5946__bF_buf0), .Y(_5948_) );
OAI21X1 OAI21X1_901 ( .A(_5278__bF_buf1), .B(_5946__bF_buf0), .C(_5948_), .Y(_1109_) );
NAND3X1 NAND3X1_777 ( .A(datapath_1_RegisterFile_regfile_mem_19__2_), .B(_5265__bF_buf71), .C(_5946__bF_buf5), .Y(_5949_) );
OAI21X1 OAI21X1_902 ( .A(_5280__bF_buf3), .B(_5946__bF_buf5), .C(_5949_), .Y(_1119_) );
NAND3X1 NAND3X1_778 ( .A(datapath_1_RegisterFile_regfile_mem_19__3_), .B(_5265__bF_buf14), .C(_5946__bF_buf3), .Y(_5950_) );
OAI21X1 OAI21X1_903 ( .A(_5282__bF_buf1), .B(_5946__bF_buf3), .C(_5950_), .Y(_1122_) );
NAND3X1 NAND3X1_779 ( .A(datapath_1_RegisterFile_regfile_mem_19__4_), .B(_5265__bF_buf49), .C(_5946__bF_buf6), .Y(_5951_) );
OAI21X1 OAI21X1_904 ( .A(_5284__bF_buf0), .B(_5946__bF_buf6), .C(_5951_), .Y(_1123_) );
NAND3X1 NAND3X1_780 ( .A(datapath_1_RegisterFile_regfile_mem_19__5_), .B(_5265__bF_buf15), .C(_5946__bF_buf1), .Y(_5952_) );
OAI21X1 OAI21X1_905 ( .A(_5286__bF_buf2), .B(_5946__bF_buf1), .C(_5952_), .Y(_1124_) );
NAND3X1 NAND3X1_781 ( .A(datapath_1_RegisterFile_regfile_mem_19__6_), .B(_5265__bF_buf67), .C(_5946__bF_buf2), .Y(_5953_) );
OAI21X1 OAI21X1_906 ( .A(_5288__bF_buf1), .B(_5946__bF_buf2), .C(_5953_), .Y(_1125_) );
NAND3X1 NAND3X1_782 ( .A(datapath_1_RegisterFile_regfile_mem_19__7_), .B(_5265__bF_buf71), .C(_5946__bF_buf3), .Y(_5954_) );
OAI21X1 OAI21X1_907 ( .A(_5290__bF_buf2), .B(_5946__bF_buf3), .C(_5954_), .Y(_1743_) );
NAND3X1 NAND3X1_783 ( .A(datapath_1_RegisterFile_regfile_mem_19__8_), .B(_5265__bF_buf54), .C(_5946__bF_buf6), .Y(_5955_) );
OAI21X1 OAI21X1_908 ( .A(_5292__bF_buf0), .B(_5946__bF_buf6), .C(_5955_), .Y(_1126_) );
NAND3X1 NAND3X1_784 ( .A(datapath_1_RegisterFile_regfile_mem_19__9_), .B(_5265__bF_buf17), .C(_5946__bF_buf1), .Y(_5956_) );
OAI21X1 OAI21X1_909 ( .A(_5294__bF_buf1), .B(_5946__bF_buf1), .C(_5956_), .Y(_1127_) );
NAND3X1 NAND3X1_785 ( .A(datapath_1_RegisterFile_regfile_mem_19__10_), .B(_5265__bF_buf79), .C(_5946__bF_buf4), .Y(_5957_) );
OAI21X1 OAI21X1_910 ( .A(_5296__bF_buf0), .B(_5946__bF_buf4), .C(_5957_), .Y(_1100_) );
NAND3X1 NAND3X1_786 ( .A(datapath_1_RegisterFile_regfile_mem_19__11_), .B(_5265__bF_buf71), .C(_5946__bF_buf5), .Y(_5958_) );
OAI21X1 OAI21X1_911 ( .A(_5298__bF_buf1), .B(_5946__bF_buf5), .C(_5958_), .Y(_1101_) );
NAND3X1 NAND3X1_787 ( .A(datapath_1_RegisterFile_regfile_mem_19__12_), .B(_5265__bF_buf40), .C(_5946__bF_buf2), .Y(_5959_) );
OAI21X1 OAI21X1_912 ( .A(_5300__bF_buf2), .B(_5946__bF_buf2), .C(_5959_), .Y(_1102_) );
NAND3X1 NAND3X1_788 ( .A(datapath_1_RegisterFile_regfile_mem_19__13_), .B(_5265__bF_buf58), .C(_5946__bF_buf4), .Y(_5960_) );
OAI21X1 OAI21X1_913 ( .A(_5302__bF_buf1), .B(_5946__bF_buf4), .C(_5960_), .Y(_1103_) );
NAND3X1 NAND3X1_789 ( .A(datapath_1_RegisterFile_regfile_mem_19__14_), .B(_5265__bF_buf17), .C(_5946__bF_buf1), .Y(_5961_) );
OAI21X1 OAI21X1_914 ( .A(_5304__bF_buf2), .B(_5946__bF_buf1), .C(_5961_), .Y(_1104_) );
NAND3X1 NAND3X1_790 ( .A(datapath_1_RegisterFile_regfile_mem_19__15_), .B(_5265__bF_buf71), .C(_5946__bF_buf5), .Y(_5962_) );
OAI21X1 OAI21X1_915 ( .A(_5306__bF_buf2), .B(_5946__bF_buf5), .C(_5962_), .Y(_1105_) );
NAND3X1 NAND3X1_791 ( .A(datapath_1_RegisterFile_regfile_mem_19__16_), .B(_5265__bF_buf80), .C(_5946__bF_buf2), .Y(_5963_) );
OAI21X1 OAI21X1_916 ( .A(_5308__bF_buf4), .B(_5946__bF_buf2), .C(_5963_), .Y(_1106_) );
NAND3X1 NAND3X1_792 ( .A(datapath_1_RegisterFile_regfile_mem_19__17_), .B(_5265__bF_buf49), .C(_5946__bF_buf6), .Y(_5964_) );
OAI21X1 OAI21X1_917 ( .A(_5310__bF_buf0), .B(_5946__bF_buf6), .C(_5964_), .Y(_1744_) );
NAND3X1 NAND3X1_793 ( .A(datapath_1_RegisterFile_regfile_mem_19__18_), .B(_5265__bF_buf58), .C(_5946__bF_buf4), .Y(_5965_) );
OAI21X1 OAI21X1_918 ( .A(_5312__bF_buf2), .B(_5946__bF_buf4), .C(_5965_), .Y(_1107_) );
NAND3X1 NAND3X1_794 ( .A(datapath_1_RegisterFile_regfile_mem_19__19_), .B(_5265__bF_buf71), .C(_5946__bF_buf5), .Y(_5966_) );
OAI21X1 OAI21X1_919 ( .A(_5314__bF_buf4), .B(_5946__bF_buf5), .C(_5966_), .Y(_1108_) );
NAND3X1 NAND3X1_795 ( .A(datapath_1_RegisterFile_regfile_mem_19__20_), .B(_5265__bF_buf88), .C(_5946__bF_buf3), .Y(_5967_) );
OAI21X1 OAI21X1_920 ( .A(_5316__bF_buf4), .B(_5946__bF_buf3), .C(_5967_), .Y(_1110_) );
NAND3X1 NAND3X1_796 ( .A(datapath_1_RegisterFile_regfile_mem_19__21_), .B(_5265__bF_buf54), .C(_5946__bF_buf6), .Y(_5968_) );
OAI21X1 OAI21X1_921 ( .A(_5318__bF_buf1), .B(_5946__bF_buf6), .C(_5968_), .Y(_1111_) );
NAND3X1 NAND3X1_797 ( .A(datapath_1_RegisterFile_regfile_mem_19__22_), .B(_5265__bF_buf66), .C(_5946__bF_buf7), .Y(_5969_) );
OAI21X1 OAI21X1_922 ( .A(_5320__bF_buf1), .B(_5946__bF_buf7), .C(_5969_), .Y(_1112_) );
NAND3X1 NAND3X1_798 ( .A(datapath_1_RegisterFile_regfile_mem_19__23_), .B(_5265__bF_buf46), .C(_5946__bF_buf2), .Y(_5970_) );
OAI21X1 OAI21X1_923 ( .A(_5322__bF_buf4), .B(_5946__bF_buf2), .C(_5970_), .Y(_1113_) );
NAND3X1 NAND3X1_799 ( .A(datapath_1_RegisterFile_regfile_mem_19__24_), .B(_5265__bF_buf32), .C(_5946__bF_buf0), .Y(_5971_) );
OAI21X1 OAI21X1_924 ( .A(_5324__bF_buf2), .B(_5946__bF_buf0), .C(_5971_), .Y(_1114_) );
NAND3X1 NAND3X1_800 ( .A(datapath_1_RegisterFile_regfile_mem_19__25_), .B(_5265__bF_buf34), .C(_5946__bF_buf0), .Y(_5972_) );
OAI21X1 OAI21X1_925 ( .A(_5326__bF_buf4), .B(_5946__bF_buf0), .C(_5972_), .Y(_1115_) );
NAND3X1 NAND3X1_801 ( .A(datapath_1_RegisterFile_regfile_mem_19__26_), .B(_5265__bF_buf47), .C(_5946__bF_buf7), .Y(_5973_) );
OAI21X1 OAI21X1_926 ( .A(_5328__bF_buf4), .B(_5946__bF_buf7), .C(_5973_), .Y(_1116_) );
NAND3X1 NAND3X1_802 ( .A(datapath_1_RegisterFile_regfile_mem_19__27_), .B(_5265__bF_buf29), .C(_5946__bF_buf4), .Y(_5974_) );
OAI21X1 OAI21X1_927 ( .A(_5330__bF_buf2), .B(_5946__bF_buf4), .C(_5974_), .Y(_1745_) );
NAND3X1 NAND3X1_803 ( .A(datapath_1_RegisterFile_regfile_mem_19__28_), .B(_5265__bF_buf78), .C(_5946__bF_buf3), .Y(_5975_) );
OAI21X1 OAI21X1_928 ( .A(_5332__bF_buf3), .B(_5946__bF_buf3), .C(_5975_), .Y(_1117_) );
NAND3X1 NAND3X1_804 ( .A(datapath_1_RegisterFile_regfile_mem_19__29_), .B(_5265__bF_buf34), .C(_5946__bF_buf0), .Y(_5976_) );
OAI21X1 OAI21X1_929 ( .A(_5334__bF_buf3), .B(_5946__bF_buf0), .C(_5976_), .Y(_1118_) );
NAND3X1 NAND3X1_805 ( .A(datapath_1_RegisterFile_regfile_mem_19__30_), .B(_5265__bF_buf82), .C(_5946__bF_buf7), .Y(_5977_) );
OAI21X1 OAI21X1_930 ( .A(_5336__bF_buf3), .B(_5946__bF_buf7), .C(_5977_), .Y(_1120_) );
NAND3X1 NAND3X1_806 ( .A(datapath_1_RegisterFile_regfile_mem_19__31_), .B(_5265__bF_buf81), .C(_5946__bF_buf1), .Y(_5978_) );
OAI21X1 OAI21X1_931 ( .A(_5338__bF_buf2), .B(_5946__bF_buf1), .C(_5978_), .Y(_1121_) );
NOR2X1 NOR2X1_139 ( .A(_5444_), .B(_5845_), .Y(_5979_) );
NAND2X1 NAND2X1_384 ( .A(_5274_), .B(_5979_), .Y(_5980_) );
NAND3X1 NAND3X1_807 ( .A(datapath_1_RegisterFile_regfile_mem_20__0_), .B(_5265__bF_buf1), .C(_5980__bF_buf0), .Y(_5981_) );
OAI21X1 OAI21X1_932 ( .A(_5276__bF_buf4), .B(_5980__bF_buf0), .C(_5981_), .Y(_1149_) );
NAND3X1 NAND3X1_808 ( .A(datapath_1_RegisterFile_regfile_mem_20__1_), .B(_5265__bF_buf67), .C(_5980__bF_buf1), .Y(_5982_) );
OAI21X1 OAI21X1_933 ( .A(_5278__bF_buf3), .B(_5980__bF_buf1), .C(_5982_), .Y(_1159_) );
NAND3X1 NAND3X1_809 ( .A(datapath_1_RegisterFile_regfile_mem_20__2_), .B(_5265__bF_buf34), .C(_5980__bF_buf6), .Y(_5983_) );
OAI21X1 OAI21X1_934 ( .A(_5280__bF_buf3), .B(_5980__bF_buf6), .C(_5983_), .Y(_1746_) );
NAND3X1 NAND3X1_810 ( .A(datapath_1_RegisterFile_regfile_mem_20__3_), .B(_5265__bF_buf69), .C(_5980__bF_buf4), .Y(_5984_) );
OAI21X1 OAI21X1_935 ( .A(_5282__bF_buf1), .B(_5980__bF_buf4), .C(_5984_), .Y(_1171_) );
NAND3X1 NAND3X1_811 ( .A(datapath_1_RegisterFile_regfile_mem_20__4_), .B(_5265__bF_buf46), .C(_5980__bF_buf5), .Y(_5985_) );
OAI21X1 OAI21X1_936 ( .A(_5284__bF_buf3), .B(_5980__bF_buf5), .C(_5985_), .Y(_1172_) );
NAND3X1 NAND3X1_812 ( .A(datapath_1_RegisterFile_regfile_mem_20__5_), .B(_5265__bF_buf79), .C(_5980__bF_buf7), .Y(_5986_) );
OAI21X1 OAI21X1_937 ( .A(_5286__bF_buf2), .B(_5980__bF_buf7), .C(_5986_), .Y(_1173_) );
NAND3X1 NAND3X1_813 ( .A(datapath_1_RegisterFile_regfile_mem_20__6_), .B(_5265__bF_buf95), .C(_5980__bF_buf2), .Y(_5987_) );
OAI21X1 OAI21X1_938 ( .A(_5288__bF_buf0), .B(_5980__bF_buf2), .C(_5987_), .Y(_1174_) );
NAND3X1 NAND3X1_814 ( .A(datapath_1_RegisterFile_regfile_mem_20__7_), .B(_5265__bF_buf14), .C(_5980__bF_buf4), .Y(_5988_) );
OAI21X1 OAI21X1_939 ( .A(_5290__bF_buf3), .B(_5980__bF_buf4), .C(_5988_), .Y(_1175_) );
NAND3X1 NAND3X1_815 ( .A(datapath_1_RegisterFile_regfile_mem_20__8_), .B(_5265__bF_buf46), .C(_5980__bF_buf5), .Y(_5989_) );
OAI21X1 OAI21X1_940 ( .A(_5292__bF_buf2), .B(_5980__bF_buf5), .C(_5989_), .Y(_1176_) );
NAND3X1 NAND3X1_816 ( .A(datapath_1_RegisterFile_regfile_mem_20__9_), .B(_5265__bF_buf37), .C(_5980__bF_buf7), .Y(_5990_) );
OAI21X1 OAI21X1_941 ( .A(_5294__bF_buf4), .B(_5980__bF_buf7), .C(_5990_), .Y(_1177_) );
NAND3X1 NAND3X1_817 ( .A(datapath_1_RegisterFile_regfile_mem_20__10_), .B(_5265__bF_buf90), .C(_5980__bF_buf0), .Y(_5991_) );
OAI21X1 OAI21X1_942 ( .A(_5296__bF_buf3), .B(_5980__bF_buf0), .C(_5991_), .Y(_1150_) );
NAND3X1 NAND3X1_818 ( .A(datapath_1_RegisterFile_regfile_mem_20__11_), .B(_5265__bF_buf11), .C(_5980__bF_buf6), .Y(_5992_) );
OAI21X1 OAI21X1_943 ( .A(_5298__bF_buf1), .B(_5980__bF_buf6), .C(_5992_), .Y(_1151_) );
NAND3X1 NAND3X1_819 ( .A(datapath_1_RegisterFile_regfile_mem_20__12_), .B(_5265__bF_buf19), .C(_5980__bF_buf2), .Y(_5993_) );
OAI21X1 OAI21X1_944 ( .A(_5300__bF_buf2), .B(_5980__bF_buf2), .C(_5993_), .Y(_1747_) );
NAND3X1 NAND3X1_820 ( .A(datapath_1_RegisterFile_regfile_mem_20__13_), .B(_5265__bF_buf17), .C(_5980__bF_buf3), .Y(_5994_) );
OAI21X1 OAI21X1_945 ( .A(_5302__bF_buf1), .B(_5980__bF_buf3), .C(_5994_), .Y(_1152_) );
NAND3X1 NAND3X1_821 ( .A(datapath_1_RegisterFile_regfile_mem_20__14_), .B(_5265__bF_buf17), .C(_5980__bF_buf3), .Y(_5995_) );
OAI21X1 OAI21X1_946 ( .A(_5304__bF_buf2), .B(_5980__bF_buf3), .C(_5995_), .Y(_1153_) );
NAND3X1 NAND3X1_822 ( .A(datapath_1_RegisterFile_regfile_mem_20__15_), .B(_5265__bF_buf10), .C(_5980__bF_buf4), .Y(_5996_) );
OAI21X1 OAI21X1_947 ( .A(_5306__bF_buf0), .B(_5980__bF_buf4), .C(_5996_), .Y(_1154_) );
NAND3X1 NAND3X1_823 ( .A(datapath_1_RegisterFile_regfile_mem_20__16_), .B(_5265__bF_buf41), .C(_5980__bF_buf1), .Y(_5997_) );
OAI21X1 OAI21X1_948 ( .A(_5308__bF_buf4), .B(_5980__bF_buf1), .C(_5997_), .Y(_1155_) );
NAND3X1 NAND3X1_824 ( .A(datapath_1_RegisterFile_regfile_mem_20__17_), .B(_5265__bF_buf8), .C(_5980__bF_buf5), .Y(_5998_) );
OAI21X1 OAI21X1_949 ( .A(_5310__bF_buf3), .B(_5980__bF_buf5), .C(_5998_), .Y(_1156_) );
NAND3X1 NAND3X1_825 ( .A(datapath_1_RegisterFile_regfile_mem_20__18_), .B(_5265__bF_buf17), .C(_5980__bF_buf3), .Y(_5999_) );
OAI21X1 OAI21X1_950 ( .A(_5312__bF_buf2), .B(_5980__bF_buf3), .C(_5999_), .Y(_1157_) );
NAND3X1 NAND3X1_826 ( .A(datapath_1_RegisterFile_regfile_mem_20__19_), .B(_5265__bF_buf11), .C(_5980__bF_buf6), .Y(_6000_) );
OAI21X1 OAI21X1_951 ( .A(_5314__bF_buf4), .B(_5980__bF_buf6), .C(_6000_), .Y(_1158_) );
NAND3X1 NAND3X1_827 ( .A(datapath_1_RegisterFile_regfile_mem_20__20_), .B(_5265__bF_buf14), .C(_5980__bF_buf4), .Y(_6001_) );
OAI21X1 OAI21X1_952 ( .A(_5316__bF_buf4), .B(_5980__bF_buf4), .C(_6001_), .Y(_1160_) );
NAND3X1 NAND3X1_828 ( .A(datapath_1_RegisterFile_regfile_mem_20__21_), .B(_5265__bF_buf49), .C(_5980__bF_buf5), .Y(_6002_) );
OAI21X1 OAI21X1_953 ( .A(_5318__bF_buf3), .B(_5980__bF_buf5), .C(_6002_), .Y(_1161_) );
NAND3X1 NAND3X1_829 ( .A(datapath_1_RegisterFile_regfile_mem_20__22_), .B(_5265__bF_buf82), .C(_5980__bF_buf0), .Y(_6003_) );
OAI21X1 OAI21X1_954 ( .A(_5320__bF_buf1), .B(_5980__bF_buf0), .C(_6003_), .Y(_1748_) );
NAND3X1 NAND3X1_830 ( .A(datapath_1_RegisterFile_regfile_mem_20__23_), .B(_5265__bF_buf4), .C(_5980__bF_buf2), .Y(_6004_) );
OAI21X1 OAI21X1_955 ( .A(_5322__bF_buf0), .B(_5980__bF_buf2), .C(_6004_), .Y(_1162_) );
NAND3X1 NAND3X1_831 ( .A(datapath_1_RegisterFile_regfile_mem_20__24_), .B(_5265__bF_buf11), .C(_5980__bF_buf6), .Y(_6005_) );
OAI21X1 OAI21X1_956 ( .A(_5324__bF_buf1), .B(_5980__bF_buf6), .C(_6005_), .Y(_1163_) );
NAND3X1 NAND3X1_832 ( .A(datapath_1_RegisterFile_regfile_mem_20__25_), .B(_5265__bF_buf80), .C(_5980__bF_buf2), .Y(_6006_) );
OAI21X1 OAI21X1_957 ( .A(_5326__bF_buf3), .B(_5980__bF_buf2), .C(_6006_), .Y(_1164_) );
NAND3X1 NAND3X1_833 ( .A(datapath_1_RegisterFile_regfile_mem_20__26_), .B(_5265__bF_buf15), .C(_5980__bF_buf3), .Y(_6007_) );
OAI21X1 OAI21X1_958 ( .A(_5328__bF_buf1), .B(_5980__bF_buf3), .C(_6007_), .Y(_1165_) );
NAND3X1 NAND3X1_834 ( .A(datapath_1_RegisterFile_regfile_mem_20__27_), .B(_5265__bF_buf37), .C(_5980__bF_buf7), .Y(_6008_) );
OAI21X1 OAI21X1_959 ( .A(_5330__bF_buf1), .B(_5980__bF_buf7), .C(_6008_), .Y(_1166_) );
NAND3X1 NAND3X1_835 ( .A(datapath_1_RegisterFile_regfile_mem_20__28_), .B(_5265__bF_buf41), .C(_5980__bF_buf1), .Y(_6009_) );
OAI21X1 OAI21X1_960 ( .A(_5332__bF_buf2), .B(_5980__bF_buf1), .C(_6009_), .Y(_1167_) );
NAND3X1 NAND3X1_836 ( .A(datapath_1_RegisterFile_regfile_mem_20__29_), .B(_5265__bF_buf24), .C(_5980__bF_buf1), .Y(_6010_) );
OAI21X1 OAI21X1_961 ( .A(_5334__bF_buf3), .B(_5980__bF_buf1), .C(_6010_), .Y(_1168_) );
NAND3X1 NAND3X1_837 ( .A(datapath_1_RegisterFile_regfile_mem_20__30_), .B(_5265__bF_buf82), .C(_5980__bF_buf0), .Y(_6011_) );
OAI21X1 OAI21X1_962 ( .A(_5336__bF_buf1), .B(_5980__bF_buf0), .C(_6011_), .Y(_1169_) );
NAND3X1 NAND3X1_838 ( .A(datapath_1_RegisterFile_regfile_mem_20__31_), .B(_5265__bF_buf37), .C(_5980__bF_buf7), .Y(_6012_) );
OAI21X1 OAI21X1_963 ( .A(_5338__bF_buf1), .B(_5980__bF_buf7), .C(_6012_), .Y(_1170_) );
NAND2X1 NAND2X1_385 ( .A(_5341_), .B(_5979_), .Y(_6013_) );
NAND3X1 NAND3X1_839 ( .A(datapath_1_RegisterFile_regfile_mem_21__0_), .B(_5265__bF_buf47), .C(_6013__bF_buf6), .Y(_6014_) );
OAI21X1 OAI21X1_964 ( .A(_5276__bF_buf4), .B(_6013__bF_buf6), .C(_6014_), .Y(_1178_) );
NAND3X1 NAND3X1_840 ( .A(datapath_1_RegisterFile_regfile_mem_21__1_), .B(_5265__bF_buf24), .C(_6013__bF_buf5), .Y(_6015_) );
OAI21X1 OAI21X1_965 ( .A(_5278__bF_buf3), .B(_6013__bF_buf5), .C(_6015_), .Y(_1179_) );
NAND3X1 NAND3X1_841 ( .A(datapath_1_RegisterFile_regfile_mem_21__2_), .B(_5265__bF_buf80), .C(_6013__bF_buf3), .Y(_6016_) );
OAI21X1 OAI21X1_966 ( .A(_5280__bF_buf4), .B(_6013__bF_buf3), .C(_6016_), .Y(_1189_) );
NAND3X1 NAND3X1_842 ( .A(datapath_1_RegisterFile_regfile_mem_21__3_), .B(_5265__bF_buf10), .C(_6013__bF_buf4), .Y(_6017_) );
OAI21X1 OAI21X1_967 ( .A(_5282__bF_buf3), .B(_6013__bF_buf4), .C(_6017_), .Y(_1192_) );
NAND3X1 NAND3X1_843 ( .A(datapath_1_RegisterFile_regfile_mem_21__4_), .B(_5265__bF_buf49), .C(_6013__bF_buf7), .Y(_6018_) );
OAI21X1 OAI21X1_968 ( .A(_5284__bF_buf0), .B(_6013__bF_buf7), .C(_6018_), .Y(_1193_) );
NAND3X1 NAND3X1_844 ( .A(datapath_1_RegisterFile_regfile_mem_21__5_), .B(_5265__bF_buf15), .C(_6013__bF_buf0), .Y(_6019_) );
OAI21X1 OAI21X1_969 ( .A(_5286__bF_buf2), .B(_6013__bF_buf0), .C(_6019_), .Y(_1194_) );
NAND3X1 NAND3X1_845 ( .A(datapath_1_RegisterFile_regfile_mem_21__6_), .B(_5265__bF_buf95), .C(_6013__bF_buf3), .Y(_6020_) );
OAI21X1 OAI21X1_970 ( .A(_5288__bF_buf0), .B(_6013__bF_buf3), .C(_6020_), .Y(_1195_) );
NAND3X1 NAND3X1_846 ( .A(datapath_1_RegisterFile_regfile_mem_21__7_), .B(_5265__bF_buf78), .C(_6013__bF_buf1), .Y(_6021_) );
OAI21X1 OAI21X1_971 ( .A(_5290__bF_buf2), .B(_6013__bF_buf1), .C(_6021_), .Y(_1749_) );
NAND3X1 NAND3X1_847 ( .A(datapath_1_RegisterFile_regfile_mem_21__8_), .B(_5265__bF_buf54), .C(_6013__bF_buf7), .Y(_6022_) );
OAI21X1 OAI21X1_972 ( .A(_5292__bF_buf2), .B(_6013__bF_buf7), .C(_6022_), .Y(_1196_) );
NAND3X1 NAND3X1_848 ( .A(datapath_1_RegisterFile_regfile_mem_21__9_), .B(_5265__bF_buf29), .C(_6013__bF_buf2), .Y(_6023_) );
OAI21X1 OAI21X1_973 ( .A(_5294__bF_buf1), .B(_6013__bF_buf2), .C(_6023_), .Y(_1197_) );
NAND3X1 NAND3X1_849 ( .A(datapath_1_RegisterFile_regfile_mem_21__10_), .B(_5265__bF_buf1), .C(_6013__bF_buf6), .Y(_6024_) );
OAI21X1 OAI21X1_974 ( .A(_5296__bF_buf0), .B(_6013__bF_buf6), .C(_6024_), .Y(_1750_) );
NAND3X1 NAND3X1_850 ( .A(datapath_1_RegisterFile_regfile_mem_21__11_), .B(_5265__bF_buf78), .C(_6013__bF_buf1), .Y(_6025_) );
OAI21X1 OAI21X1_975 ( .A(_5298__bF_buf4), .B(_6013__bF_buf1), .C(_6025_), .Y(_1751_) );
NAND3X1 NAND3X1_851 ( .A(datapath_1_RegisterFile_regfile_mem_21__12_), .B(_5265__bF_buf40), .C(_6013__bF_buf1), .Y(_6026_) );
OAI21X1 OAI21X1_976 ( .A(_5300__bF_buf2), .B(_6013__bF_buf1), .C(_6026_), .Y(_1752_) );
NAND3X1 NAND3X1_852 ( .A(datapath_1_RegisterFile_regfile_mem_21__13_), .B(_5265__bF_buf15), .C(_6013__bF_buf0), .Y(_6027_) );
OAI21X1 OAI21X1_977 ( .A(_5302__bF_buf3), .B(_6013__bF_buf0), .C(_6027_), .Y(_1753_) );
NAND3X1 NAND3X1_853 ( .A(datapath_1_RegisterFile_regfile_mem_21__14_), .B(_5265__bF_buf81), .C(_6013__bF_buf2), .Y(_6028_) );
OAI21X1 OAI21X1_978 ( .A(_5304__bF_buf2), .B(_6013__bF_buf2), .C(_6028_), .Y(_1754_) );
NAND3X1 NAND3X1_854 ( .A(datapath_1_RegisterFile_regfile_mem_21__15_), .B(_5265__bF_buf10), .C(_6013__bF_buf4), .Y(_6029_) );
OAI21X1 OAI21X1_979 ( .A(_5306__bF_buf0), .B(_6013__bF_buf4), .C(_6029_), .Y(_1755_) );
NAND3X1 NAND3X1_855 ( .A(datapath_1_RegisterFile_regfile_mem_21__16_), .B(_5265__bF_buf24), .C(_6013__bF_buf5), .Y(_6030_) );
OAI21X1 OAI21X1_980 ( .A(_5308__bF_buf1), .B(_6013__bF_buf5), .C(_6030_), .Y(_1756_) );
NAND3X1 NAND3X1_856 ( .A(datapath_1_RegisterFile_regfile_mem_21__17_), .B(_5265__bF_buf49), .C(_6013__bF_buf7), .Y(_6031_) );
OAI21X1 OAI21X1_981 ( .A(_5310__bF_buf0), .B(_6013__bF_buf7), .C(_6031_), .Y(_1757_) );
NAND3X1 NAND3X1_857 ( .A(datapath_1_RegisterFile_regfile_mem_21__18_), .B(_5265__bF_buf17), .C(_6013__bF_buf0), .Y(_6032_) );
OAI21X1 OAI21X1_982 ( .A(_5312__bF_buf2), .B(_6013__bF_buf0), .C(_6032_), .Y(_1758_) );
NAND3X1 NAND3X1_858 ( .A(datapath_1_RegisterFile_regfile_mem_21__19_), .B(_5265__bF_buf14), .C(_6013__bF_buf4), .Y(_6033_) );
OAI21X1 OAI21X1_983 ( .A(_5314__bF_buf2), .B(_6013__bF_buf4), .C(_6033_), .Y(_1759_) );
NAND3X1 NAND3X1_859 ( .A(datapath_1_RegisterFile_regfile_mem_21__20_), .B(_5265__bF_buf88), .C(_6013__bF_buf4), .Y(_6034_) );
OAI21X1 OAI21X1_984 ( .A(_5316__bF_buf4), .B(_6013__bF_buf4), .C(_6034_), .Y(_1180_) );
NAND3X1 NAND3X1_860 ( .A(datapath_1_RegisterFile_regfile_mem_21__21_), .B(_5265__bF_buf46), .C(_6013__bF_buf7), .Y(_6035_) );
OAI21X1 OAI21X1_985 ( .A(_5318__bF_buf1), .B(_6013__bF_buf7), .C(_6035_), .Y(_1181_) );
NAND3X1 NAND3X1_861 ( .A(datapath_1_RegisterFile_regfile_mem_21__22_), .B(_5265__bF_buf82), .C(_6013__bF_buf6), .Y(_6036_) );
OAI21X1 OAI21X1_986 ( .A(_5320__bF_buf0), .B(_6013__bF_buf6), .C(_6036_), .Y(_1182_) );
NAND3X1 NAND3X1_862 ( .A(datapath_1_RegisterFile_regfile_mem_21__23_), .B(_5265__bF_buf4), .C(_6013__bF_buf3), .Y(_6037_) );
OAI21X1 OAI21X1_987 ( .A(_5322__bF_buf0), .B(_6013__bF_buf3), .C(_6037_), .Y(_1183_) );
NAND3X1 NAND3X1_863 ( .A(datapath_1_RegisterFile_regfile_mem_21__24_), .B(_5265__bF_buf16), .C(_6013__bF_buf5), .Y(_6038_) );
OAI21X1 OAI21X1_988 ( .A(_5324__bF_buf2), .B(_6013__bF_buf5), .C(_6038_), .Y(_1184_) );
NAND3X1 NAND3X1_864 ( .A(datapath_1_RegisterFile_regfile_mem_21__25_), .B(_5265__bF_buf19), .C(_6013__bF_buf3), .Y(_6039_) );
OAI21X1 OAI21X1_989 ( .A(_5326__bF_buf0), .B(_6013__bF_buf3), .C(_6039_), .Y(_1185_) );
NAND3X1 NAND3X1_865 ( .A(datapath_1_RegisterFile_regfile_mem_21__26_), .B(_5265__bF_buf15), .C(_6013__bF_buf0), .Y(_6040_) );
OAI21X1 OAI21X1_990 ( .A(_5328__bF_buf1), .B(_6013__bF_buf0), .C(_6040_), .Y(_1186_) );
NAND3X1 NAND3X1_866 ( .A(datapath_1_RegisterFile_regfile_mem_21__27_), .B(_5265__bF_buf81), .C(_6013__bF_buf2), .Y(_6041_) );
OAI21X1 OAI21X1_991 ( .A(_5330__bF_buf2), .B(_6013__bF_buf2), .C(_6041_), .Y(_1760_) );
NAND3X1 NAND3X1_867 ( .A(datapath_1_RegisterFile_regfile_mem_21__28_), .B(_5265__bF_buf88), .C(_6013__bF_buf1), .Y(_6042_) );
OAI21X1 OAI21X1_992 ( .A(_5332__bF_buf3), .B(_6013__bF_buf1), .C(_6042_), .Y(_1187_) );
NAND3X1 NAND3X1_868 ( .A(datapath_1_RegisterFile_regfile_mem_21__29_), .B(_5265__bF_buf41), .C(_6013__bF_buf5), .Y(_6043_) );
OAI21X1 OAI21X1_993 ( .A(_5334__bF_buf3), .B(_6013__bF_buf5), .C(_6043_), .Y(_1188_) );
NAND3X1 NAND3X1_869 ( .A(datapath_1_RegisterFile_regfile_mem_21__30_), .B(_5265__bF_buf66), .C(_6013__bF_buf6), .Y(_6044_) );
OAI21X1 OAI21X1_994 ( .A(_5336__bF_buf3), .B(_6013__bF_buf6), .C(_6044_), .Y(_1190_) );
NAND3X1 NAND3X1_870 ( .A(datapath_1_RegisterFile_regfile_mem_21__31_), .B(_5265__bF_buf17), .C(_6013__bF_buf2), .Y(_6045_) );
OAI21X1 OAI21X1_995 ( .A(_5338__bF_buf2), .B(_6013__bF_buf2), .C(_6045_), .Y(_1191_) );
NAND2X1 NAND2X1_386 ( .A(_5376_), .B(_5979_), .Y(_6046_) );
NAND3X1 NAND3X1_871 ( .A(datapath_1_RegisterFile_regfile_mem_22__0_), .B(_5265__bF_buf1), .C(_6046__bF_buf6), .Y(_6047_) );
OAI21X1 OAI21X1_996 ( .A(_5276__bF_buf4), .B(_6046__bF_buf6), .C(_6047_), .Y(_1761_) );
NAND3X1 NAND3X1_872 ( .A(datapath_1_RegisterFile_regfile_mem_22__1_), .B(_5265__bF_buf24), .C(_6046__bF_buf2), .Y(_6048_) );
OAI21X1 OAI21X1_997 ( .A(_5278__bF_buf1), .B(_6046__bF_buf2), .C(_6048_), .Y(_1762_) );
NAND3X1 NAND3X1_873 ( .A(datapath_1_RegisterFile_regfile_mem_22__2_), .B(_5265__bF_buf40), .C(_6046__bF_buf1), .Y(_6049_) );
OAI21X1 OAI21X1_998 ( .A(_5280__bF_buf4), .B(_6046__bF_buf1), .C(_6049_), .Y(_1763_) );
NAND3X1 NAND3X1_874 ( .A(datapath_1_RegisterFile_regfile_mem_22__3_), .B(_5265__bF_buf69), .C(_6046__bF_buf4), .Y(_6050_) );
OAI21X1 OAI21X1_999 ( .A(_5282__bF_buf3), .B(_6046__bF_buf4), .C(_6050_), .Y(_1764_) );
NAND3X1 NAND3X1_875 ( .A(datapath_1_RegisterFile_regfile_mem_22__4_), .B(_5265__bF_buf8), .C(_6046__bF_buf5), .Y(_6051_) );
OAI21X1 OAI21X1_1000 ( .A(_5284__bF_buf0), .B(_6046__bF_buf5), .C(_6051_), .Y(_1765_) );
NAND3X1 NAND3X1_876 ( .A(datapath_1_RegisterFile_regfile_mem_22__5_), .B(_5265__bF_buf79), .C(_6046__bF_buf3), .Y(_6052_) );
OAI21X1 OAI21X1_1001 ( .A(_5286__bF_buf2), .B(_6046__bF_buf3), .C(_6052_), .Y(_1766_) );
NAND3X1 NAND3X1_877 ( .A(datapath_1_RegisterFile_regfile_mem_22__6_), .B(_5265__bF_buf54), .C(_6046__bF_buf5), .Y(_6053_) );
OAI21X1 OAI21X1_1002 ( .A(_5288__bF_buf1), .B(_6046__bF_buf5), .C(_6053_), .Y(_1767_) );
NAND3X1 NAND3X1_878 ( .A(datapath_1_RegisterFile_regfile_mem_22__7_), .B(_5265__bF_buf69), .C(_6046__bF_buf4), .Y(_6054_) );
OAI21X1 OAI21X1_1003 ( .A(_5290__bF_buf3), .B(_6046__bF_buf4), .C(_6054_), .Y(_1768_) );
NAND3X1 NAND3X1_879 ( .A(datapath_1_RegisterFile_regfile_mem_22__8_), .B(_5265__bF_buf54), .C(_6046__bF_buf5), .Y(_6055_) );
OAI21X1 OAI21X1_1004 ( .A(_5292__bF_buf2), .B(_6046__bF_buf5), .C(_6055_), .Y(_1769_) );
NAND3X1 NAND3X1_880 ( .A(datapath_1_RegisterFile_regfile_mem_22__9_), .B(_5265__bF_buf29), .C(_6046__bF_buf0), .Y(_6056_) );
OAI21X1 OAI21X1_1005 ( .A(_5294__bF_buf1), .B(_6046__bF_buf0), .C(_6056_), .Y(_1770_) );
NAND3X1 NAND3X1_881 ( .A(datapath_1_RegisterFile_regfile_mem_22__10_), .B(_5265__bF_buf90), .C(_6046__bF_buf6), .Y(_6057_) );
OAI21X1 OAI21X1_1006 ( .A(_5296__bF_buf1), .B(_6046__bF_buf6), .C(_6057_), .Y(_1771_) );
NAND3X1 NAND3X1_882 ( .A(datapath_1_RegisterFile_regfile_mem_22__11_), .B(_5265__bF_buf78), .C(_6046__bF_buf1), .Y(_6058_) );
OAI21X1 OAI21X1_1007 ( .A(_5298__bF_buf1), .B(_6046__bF_buf1), .C(_6058_), .Y(_1772_) );
NAND3X1 NAND3X1_883 ( .A(datapath_1_RegisterFile_regfile_mem_22__12_), .B(_5265__bF_buf19), .C(_6046__bF_buf7), .Y(_6059_) );
OAI21X1 OAI21X1_1008 ( .A(_5300__bF_buf2), .B(_6046__bF_buf7), .C(_6059_), .Y(_1773_) );
NAND3X1 NAND3X1_884 ( .A(datapath_1_RegisterFile_regfile_mem_22__13_), .B(_5265__bF_buf79), .C(_6046__bF_buf3), .Y(_6060_) );
OAI21X1 OAI21X1_1009 ( .A(_5302__bF_buf1), .B(_6046__bF_buf3), .C(_6060_), .Y(_1774_) );
NAND3X1 NAND3X1_885 ( .A(datapath_1_RegisterFile_regfile_mem_22__14_), .B(_5265__bF_buf37), .C(_6046__bF_buf0), .Y(_6061_) );
OAI21X1 OAI21X1_1010 ( .A(_5304__bF_buf4), .B(_6046__bF_buf0), .C(_6061_), .Y(_1775_) );
NAND3X1 NAND3X1_886 ( .A(datapath_1_RegisterFile_regfile_mem_22__15_), .B(_5265__bF_buf69), .C(_6046__bF_buf4), .Y(_6062_) );
OAI21X1 OAI21X1_1011 ( .A(_5306__bF_buf0), .B(_6046__bF_buf4), .C(_6062_), .Y(_1776_) );
NAND3X1 NAND3X1_887 ( .A(datapath_1_RegisterFile_regfile_mem_22__16_), .B(_5265__bF_buf24), .C(_6046__bF_buf2), .Y(_6063_) );
OAI21X1 OAI21X1_1012 ( .A(_5308__bF_buf1), .B(_6046__bF_buf2), .C(_6063_), .Y(_1777_) );
NAND3X1 NAND3X1_888 ( .A(datapath_1_RegisterFile_regfile_mem_22__17_), .B(_5265__bF_buf8), .C(_6046__bF_buf5), .Y(_6064_) );
OAI21X1 OAI21X1_1013 ( .A(_5310__bF_buf3), .B(_6046__bF_buf5), .C(_6064_), .Y(_1778_) );
NAND3X1 NAND3X1_889 ( .A(datapath_1_RegisterFile_regfile_mem_22__18_), .B(_5265__bF_buf58), .C(_6046__bF_buf3), .Y(_6065_) );
OAI21X1 OAI21X1_1014 ( .A(_5312__bF_buf2), .B(_6046__bF_buf3), .C(_6065_), .Y(_1779_) );
NAND3X1 NAND3X1_890 ( .A(datapath_1_RegisterFile_regfile_mem_22__19_), .B(_5265__bF_buf78), .C(_6046__bF_buf1), .Y(_6066_) );
OAI21X1 OAI21X1_1015 ( .A(_5314__bF_buf4), .B(_6046__bF_buf1), .C(_6066_), .Y(_1780_) );
NAND3X1 NAND3X1_891 ( .A(datapath_1_RegisterFile_regfile_mem_22__20_), .B(_5265__bF_buf10), .C(_6046__bF_buf4), .Y(_6067_) );
OAI21X1 OAI21X1_1016 ( .A(_5316__bF_buf0), .B(_6046__bF_buf4), .C(_6067_), .Y(_1781_) );
NAND3X1 NAND3X1_892 ( .A(datapath_1_RegisterFile_regfile_mem_22__21_), .B(_5265__bF_buf4), .C(_6046__bF_buf7), .Y(_6068_) );
OAI21X1 OAI21X1_1017 ( .A(_5318__bF_buf2), .B(_6046__bF_buf7), .C(_6068_), .Y(_1782_) );
NAND3X1 NAND3X1_893 ( .A(datapath_1_RegisterFile_regfile_mem_22__22_), .B(_5265__bF_buf82), .C(_6046__bF_buf6), .Y(_6069_) );
OAI21X1 OAI21X1_1018 ( .A(_5320__bF_buf0), .B(_6046__bF_buf6), .C(_6069_), .Y(_1783_) );
NAND3X1 NAND3X1_894 ( .A(datapath_1_RegisterFile_regfile_mem_22__23_), .B(_5265__bF_buf4), .C(_6046__bF_buf7), .Y(_6070_) );
OAI21X1 OAI21X1_1019 ( .A(_5322__bF_buf0), .B(_6046__bF_buf7), .C(_6070_), .Y(_1784_) );
NAND3X1 NAND3X1_895 ( .A(datapath_1_RegisterFile_regfile_mem_22__24_), .B(_5265__bF_buf11), .C(_6046__bF_buf1), .Y(_6071_) );
OAI21X1 OAI21X1_1020 ( .A(_5324__bF_buf1), .B(_6046__bF_buf1), .C(_6071_), .Y(_1785_) );
NAND3X1 NAND3X1_896 ( .A(datapath_1_RegisterFile_regfile_mem_22__25_), .B(_5265__bF_buf19), .C(_6046__bF_buf7), .Y(_6072_) );
OAI21X1 OAI21X1_1021 ( .A(_5326__bF_buf0), .B(_6046__bF_buf7), .C(_6072_), .Y(_1786_) );
NAND3X1 NAND3X1_897 ( .A(datapath_1_RegisterFile_regfile_mem_22__26_), .B(_5265__bF_buf1), .C(_6046__bF_buf3), .Y(_6073_) );
OAI21X1 OAI21X1_1022 ( .A(_5328__bF_buf4), .B(_6046__bF_buf3), .C(_6073_), .Y(_1787_) );
NAND3X1 NAND3X1_898 ( .A(datapath_1_RegisterFile_regfile_mem_22__27_), .B(_5265__bF_buf29), .C(_6046__bF_buf0), .Y(_6074_) );
OAI21X1 OAI21X1_1023 ( .A(_5330__bF_buf2), .B(_6046__bF_buf0), .C(_6074_), .Y(_1788_) );
NAND3X1 NAND3X1_899 ( .A(datapath_1_RegisterFile_regfile_mem_22__28_), .B(_5265__bF_buf16), .C(_6046__bF_buf2), .Y(_6075_) );
OAI21X1 OAI21X1_1024 ( .A(_5332__bF_buf2), .B(_6046__bF_buf2), .C(_6075_), .Y(_1789_) );
NAND3X1 NAND3X1_900 ( .A(datapath_1_RegisterFile_regfile_mem_22__29_), .B(_5265__bF_buf41), .C(_6046__bF_buf2), .Y(_6076_) );
OAI21X1 OAI21X1_1025 ( .A(_5334__bF_buf3), .B(_6046__bF_buf2), .C(_6076_), .Y(_1790_) );
NAND3X1 NAND3X1_901 ( .A(datapath_1_RegisterFile_regfile_mem_22__30_), .B(_5265__bF_buf82), .C(_6046__bF_buf6), .Y(_6077_) );
OAI21X1 OAI21X1_1026 ( .A(_5336__bF_buf1), .B(_6046__bF_buf6), .C(_6077_), .Y(_1791_) );
NAND3X1 NAND3X1_902 ( .A(datapath_1_RegisterFile_regfile_mem_22__31_), .B(_5265__bF_buf37), .C(_6046__bF_buf0), .Y(_6078_) );
OAI21X1 OAI21X1_1027 ( .A(_5338__bF_buf1), .B(_6046__bF_buf0), .C(_6078_), .Y(_1792_) );
NAND2X1 NAND2X1_387 ( .A(_5410_), .B(_5979_), .Y(_6079_) );
NAND3X1 NAND3X1_903 ( .A(datapath_1_RegisterFile_regfile_mem_23__0_), .B(_5265__bF_buf33), .C(_6079__bF_buf3), .Y(_6080_) );
OAI21X1 OAI21X1_1028 ( .A(_5276__bF_buf3), .B(_6079__bF_buf3), .C(_6080_), .Y(_1198_) );
NAND3X1 NAND3X1_904 ( .A(datapath_1_RegisterFile_regfile_mem_23__1_), .B(_5265__bF_buf53), .C(_6079__bF_buf7), .Y(_6081_) );
OAI21X1 OAI21X1_1029 ( .A(_5278__bF_buf3), .B(_6079__bF_buf7), .C(_6081_), .Y(_1204_) );
NAND3X1 NAND3X1_905 ( .A(datapath_1_RegisterFile_regfile_mem_23__2_), .B(_5265__bF_buf34), .C(_6079__bF_buf4), .Y(_6082_) );
OAI21X1 OAI21X1_1030 ( .A(_5280__bF_buf3), .B(_6079__bF_buf4), .C(_6082_), .Y(_1209_) );
NAND3X1 NAND3X1_906 ( .A(datapath_1_RegisterFile_regfile_mem_23__3_), .B(_5265__bF_buf10), .C(_6079__bF_buf1), .Y(_6083_) );
OAI21X1 OAI21X1_1031 ( .A(_5282__bF_buf3), .B(_6079__bF_buf1), .C(_6083_), .Y(_1793_) );
NAND3X1 NAND3X1_907 ( .A(datapath_1_RegisterFile_regfile_mem_23__4_), .B(_5265__bF_buf61), .C(_6079__bF_buf5), .Y(_6084_) );
OAI21X1 OAI21X1_1032 ( .A(_5284__bF_buf2), .B(_6079__bF_buf5), .C(_6084_), .Y(_1212_) );
NAND3X1 NAND3X1_908 ( .A(datapath_1_RegisterFile_regfile_mem_23__5_), .B(_5265__bF_buf15), .C(_6079__bF_buf0), .Y(_6085_) );
OAI21X1 OAI21X1_1033 ( .A(_5286__bF_buf2), .B(_6079__bF_buf0), .C(_6085_), .Y(_1213_) );
NAND3X1 NAND3X1_909 ( .A(datapath_1_RegisterFile_regfile_mem_23__6_), .B(_5265__bF_buf53), .C(_6079__bF_buf7), .Y(_6086_) );
OAI21X1 OAI21X1_1034 ( .A(_5288__bF_buf1), .B(_6079__bF_buf7), .C(_6086_), .Y(_1214_) );
NAND3X1 NAND3X1_910 ( .A(datapath_1_RegisterFile_regfile_mem_23__7_), .B(_5265__bF_buf71), .C(_6079__bF_buf6), .Y(_6087_) );
OAI21X1 OAI21X1_1035 ( .A(_5290__bF_buf2), .B(_6079__bF_buf6), .C(_6087_), .Y(_1215_) );
NAND3X1 NAND3X1_911 ( .A(datapath_1_RegisterFile_regfile_mem_23__8_), .B(_5265__bF_buf53), .C(_6079__bF_buf7), .Y(_6088_) );
OAI21X1 OAI21X1_1036 ( .A(_5292__bF_buf0), .B(_6079__bF_buf7), .C(_6088_), .Y(_1216_) );
NAND3X1 NAND3X1_912 ( .A(datapath_1_RegisterFile_regfile_mem_23__9_), .B(_5265__bF_buf37), .C(_6079__bF_buf3), .Y(_6089_) );
OAI21X1 OAI21X1_1037 ( .A(_5294__bF_buf4), .B(_6079__bF_buf3), .C(_6089_), .Y(_1217_) );
NAND3X1 NAND3X1_913 ( .A(datapath_1_RegisterFile_regfile_mem_23__10_), .B(_5265__bF_buf15), .C(_6079__bF_buf0), .Y(_6090_) );
OAI21X1 OAI21X1_1038 ( .A(_5296__bF_buf0), .B(_6079__bF_buf0), .C(_6090_), .Y(_1199_) );
NAND3X1 NAND3X1_914 ( .A(datapath_1_RegisterFile_regfile_mem_23__11_), .B(_5265__bF_buf88), .C(_6079__bF_buf1), .Y(_6091_) );
OAI21X1 OAI21X1_1039 ( .A(_5298__bF_buf4), .B(_6079__bF_buf1), .C(_6091_), .Y(_1200_) );
NAND3X1 NAND3X1_915 ( .A(datapath_1_RegisterFile_regfile_mem_23__12_), .B(_5265__bF_buf41), .C(_6079__bF_buf4), .Y(_6092_) );
OAI21X1 OAI21X1_1040 ( .A(_5300__bF_buf2), .B(_6079__bF_buf4), .C(_6092_), .Y(_1201_) );
NAND3X1 NAND3X1_916 ( .A(datapath_1_RegisterFile_regfile_mem_23__13_), .B(_5265__bF_buf15), .C(_6079__bF_buf2), .Y(_6093_) );
OAI21X1 OAI21X1_1041 ( .A(_5302__bF_buf3), .B(_6079__bF_buf2), .C(_6093_), .Y(_1794_) );
NAND3X1 NAND3X1_917 ( .A(datapath_1_RegisterFile_regfile_mem_23__14_), .B(_5265__bF_buf37), .C(_6079__bF_buf3), .Y(_6094_) );
OAI21X1 OAI21X1_1042 ( .A(_5304__bF_buf4), .B(_6079__bF_buf3), .C(_6094_), .Y(_1202_) );
NAND3X1 NAND3X1_918 ( .A(datapath_1_RegisterFile_regfile_mem_23__15_), .B(_5265__bF_buf69), .C(_6079__bF_buf1), .Y(_6095_) );
OAI21X1 OAI21X1_1043 ( .A(_5306__bF_buf0), .B(_6079__bF_buf1), .C(_6095_), .Y(_1203_) );
NAND3X1 NAND3X1_919 ( .A(datapath_1_RegisterFile_regfile_mem_23__16_), .B(_5265__bF_buf24), .C(_6079__bF_buf7), .Y(_6096_) );
OAI21X1 OAI21X1_1044 ( .A(_5308__bF_buf1), .B(_6079__bF_buf7), .C(_6096_), .Y(_1795_) );
NAND3X1 NAND3X1_920 ( .A(datapath_1_RegisterFile_regfile_mem_23__17_), .B(_5265__bF_buf61), .C(_6079__bF_buf5), .Y(_6097_) );
OAI21X1 OAI21X1_1045 ( .A(_5310__bF_buf3), .B(_6079__bF_buf5), .C(_6097_), .Y(_1796_) );
NAND3X1 NAND3X1_921 ( .A(datapath_1_RegisterFile_regfile_mem_23__18_), .B(_5265__bF_buf15), .C(_6079__bF_buf0), .Y(_6098_) );
OAI21X1 OAI21X1_1046 ( .A(_5312__bF_buf2), .B(_6079__bF_buf0), .C(_6098_), .Y(_1797_) );
NAND3X1 NAND3X1_922 ( .A(datapath_1_RegisterFile_regfile_mem_23__19_), .B(_5265__bF_buf11), .C(_6079__bF_buf6), .Y(_6099_) );
OAI21X1 OAI21X1_1047 ( .A(_5314__bF_buf4), .B(_6079__bF_buf6), .C(_6099_), .Y(_1798_) );
NAND3X1 NAND3X1_923 ( .A(datapath_1_RegisterFile_regfile_mem_23__20_), .B(_5265__bF_buf88), .C(_6079__bF_buf1), .Y(_6100_) );
OAI21X1 OAI21X1_1048 ( .A(_5316__bF_buf4), .B(_6079__bF_buf1), .C(_6100_), .Y(_1799_) );
NAND3X1 NAND3X1_924 ( .A(datapath_1_RegisterFile_regfile_mem_23__21_), .B(_5265__bF_buf61), .C(_6079__bF_buf5), .Y(_6101_) );
OAI21X1 OAI21X1_1049 ( .A(_5318__bF_buf3), .B(_6079__bF_buf5), .C(_6101_), .Y(_1800_) );
NAND3X1 NAND3X1_925 ( .A(datapath_1_RegisterFile_regfile_mem_23__22_), .B(_5265__bF_buf1), .C(_6079__bF_buf2), .Y(_6102_) );
OAI21X1 OAI21X1_1050 ( .A(_5320__bF_buf0), .B(_6079__bF_buf2), .C(_6102_), .Y(_1801_) );
NAND3X1 NAND3X1_926 ( .A(datapath_1_RegisterFile_regfile_mem_23__23_), .B(_5265__bF_buf4), .C(_6079__bF_buf5), .Y(_6103_) );
OAI21X1 OAI21X1_1051 ( .A(_5322__bF_buf4), .B(_6079__bF_buf5), .C(_6103_), .Y(_1802_) );
NAND3X1 NAND3X1_927 ( .A(datapath_1_RegisterFile_regfile_mem_23__24_), .B(_5265__bF_buf11), .C(_6079__bF_buf6), .Y(_6104_) );
OAI21X1 OAI21X1_1052 ( .A(_5324__bF_buf1), .B(_6079__bF_buf6), .C(_6104_), .Y(_1803_) );
NAND3X1 NAND3X1_928 ( .A(datapath_1_RegisterFile_regfile_mem_23__25_), .B(_5265__bF_buf41), .C(_6079__bF_buf4), .Y(_6105_) );
OAI21X1 OAI21X1_1053 ( .A(_5326__bF_buf4), .B(_6079__bF_buf4), .C(_6105_), .Y(_1804_) );
NAND3X1 NAND3X1_929 ( .A(datapath_1_RegisterFile_regfile_mem_23__26_), .B(_5265__bF_buf47), .C(_6079__bF_buf2), .Y(_6106_) );
OAI21X1 OAI21X1_1054 ( .A(_5328__bF_buf1), .B(_6079__bF_buf2), .C(_6106_), .Y(_1205_) );
NAND3X1 NAND3X1_930 ( .A(datapath_1_RegisterFile_regfile_mem_23__27_), .B(_5265__bF_buf37), .C(_6079__bF_buf3), .Y(_6107_) );
OAI21X1 OAI21X1_1055 ( .A(_5330__bF_buf1), .B(_6079__bF_buf3), .C(_6107_), .Y(_1206_) );
NAND3X1 NAND3X1_931 ( .A(datapath_1_RegisterFile_regfile_mem_23__28_), .B(_5265__bF_buf11), .C(_6079__bF_buf6), .Y(_6108_) );
OAI21X1 OAI21X1_1056 ( .A(_5332__bF_buf2), .B(_6079__bF_buf6), .C(_6108_), .Y(_1207_) );
NAND3X1 NAND3X1_932 ( .A(datapath_1_RegisterFile_regfile_mem_23__29_), .B(_5265__bF_buf16), .C(_6079__bF_buf4), .Y(_6109_) );
OAI21X1 OAI21X1_1057 ( .A(_5334__bF_buf3), .B(_6079__bF_buf4), .C(_6109_), .Y(_1208_) );
NAND3X1 NAND3X1_933 ( .A(datapath_1_RegisterFile_regfile_mem_23__30_), .B(_5265__bF_buf66), .C(_6079__bF_buf2), .Y(_6110_) );
OAI21X1 OAI21X1_1058 ( .A(_5336__bF_buf3), .B(_6079__bF_buf2), .C(_6110_), .Y(_1210_) );
NAND3X1 NAND3X1_934 ( .A(datapath_1_RegisterFile_regfile_mem_23__31_), .B(_5265__bF_buf17), .C(_6079__bF_buf0), .Y(_6111_) );
OAI21X1 OAI21X1_1059 ( .A(_5338__bF_buf2), .B(_6079__bF_buf0), .C(_6111_), .Y(_1211_) );
NOR2X1 NOR2X1_140 ( .A(datapath_1_A3_2_), .B(_5266_), .Y(_6112_) );
INVX1 INVX1_108 ( .A(datapath_1_A3_4_), .Y(_6113_) );
OAI21X1 OAI21X1_1060 ( .A(_5264_), .B(_6113_), .C(_5272__bF_buf2), .Y(_6114_) );
NAND2X1 NAND2X1_388 ( .A(_6112_), .B(_6114_), .Y(_6115_) );
OR2X2 OR2X2_1 ( .A(_6115_), .B(_5273_), .Y(_6116_) );
NAND3X1 NAND3X1_935 ( .A(datapath_1_RegisterFile_regfile_mem_24__0_), .B(_5265__bF_buf28), .C(_6116__bF_buf3), .Y(_6117_) );
OAI21X1 OAI21X1_1061 ( .A(_5276__bF_buf1), .B(_6116__bF_buf3), .C(_6117_), .Y(_1218_) );
NAND3X1 NAND3X1_936 ( .A(datapath_1_RegisterFile_regfile_mem_24__1_), .B(_5265__bF_buf67), .C(_6116__bF_buf5), .Y(_6118_) );
OAI21X1 OAI21X1_1062 ( .A(_5278__bF_buf3), .B(_6116__bF_buf5), .C(_6118_), .Y(_1227_) );
NAND3X1 NAND3X1_937 ( .A(datapath_1_RegisterFile_regfile_mem_24__2_), .B(_5265__bF_buf19), .C(_6116__bF_buf4), .Y(_6119_) );
OAI21X1 OAI21X1_1063 ( .A(_5280__bF_buf4), .B(_6116__bF_buf4), .C(_6119_), .Y(_1229_) );
NAND3X1 NAND3X1_938 ( .A(datapath_1_RegisterFile_regfile_mem_24__3_), .B(_5265__bF_buf9), .C(_6116__bF_buf6), .Y(_6120_) );
OAI21X1 OAI21X1_1064 ( .A(_5282__bF_buf3), .B(_6116__bF_buf6), .C(_6120_), .Y(_1232_) );
NAND3X1 NAND3X1_939 ( .A(datapath_1_RegisterFile_regfile_mem_24__4_), .B(_5265__bF_buf67), .C(_6116__bF_buf5), .Y(_6121_) );
OAI21X1 OAI21X1_1065 ( .A(_5284__bF_buf3), .B(_6116__bF_buf5), .C(_6121_), .Y(_1233_) );
NAND3X1 NAND3X1_940 ( .A(datapath_1_RegisterFile_regfile_mem_24__5_), .B(_5265__bF_buf2), .C(_6116__bF_buf2), .Y(_6122_) );
OAI21X1 OAI21X1_1066 ( .A(_5286__bF_buf3), .B(_6116__bF_buf2), .C(_6122_), .Y(_1234_) );
NAND3X1 NAND3X1_941 ( .A(datapath_1_RegisterFile_regfile_mem_24__6_), .B(_5265__bF_buf75), .C(_6116__bF_buf0), .Y(_6123_) );
OAI21X1 OAI21X1_1067 ( .A(_5288__bF_buf4), .B(_6116__bF_buf0), .C(_6123_), .Y(_1805_) );
NAND3X1 NAND3X1_942 ( .A(datapath_1_RegisterFile_regfile_mem_24__7_), .B(_5265__bF_buf36), .C(_6116__bF_buf6), .Y(_6124_) );
OAI21X1 OAI21X1_1068 ( .A(_5290__bF_buf0), .B(_6116__bF_buf6), .C(_6124_), .Y(_1235_) );
NAND3X1 NAND3X1_943 ( .A(datapath_1_RegisterFile_regfile_mem_24__8_), .B(_5265__bF_buf67), .C(_6116__bF_buf5), .Y(_6125_) );
OAI21X1 OAI21X1_1069 ( .A(_5292__bF_buf0), .B(_6116__bF_buf5), .C(_6125_), .Y(_1236_) );
NAND3X1 NAND3X1_944 ( .A(datapath_1_RegisterFile_regfile_mem_24__9_), .B(_5265__bF_buf31), .C(_6116__bF_buf1), .Y(_6126_) );
OAI21X1 OAI21X1_1070 ( .A(_5294__bF_buf4), .B(_6116__bF_buf1), .C(_6126_), .Y(_1237_) );
NAND3X1 NAND3X1_945 ( .A(datapath_1_RegisterFile_regfile_mem_24__10_), .B(_5265__bF_buf90), .C(_6116__bF_buf3), .Y(_6127_) );
OAI21X1 OAI21X1_1071 ( .A(_5296__bF_buf1), .B(_6116__bF_buf3), .C(_6127_), .Y(_1219_) );
NAND3X1 NAND3X1_946 ( .A(datapath_1_RegisterFile_regfile_mem_24__11_), .B(_5265__bF_buf10), .C(_6116__bF_buf7), .Y(_6128_) );
OAI21X1 OAI21X1_1072 ( .A(_5298__bF_buf4), .B(_6116__bF_buf7), .C(_6128_), .Y(_1220_) );
NAND3X1 NAND3X1_947 ( .A(datapath_1_RegisterFile_regfile_mem_24__12_), .B(_5265__bF_buf63), .C(_6116__bF_buf4), .Y(_6129_) );
OAI21X1 OAI21X1_1073 ( .A(_5300__bF_buf4), .B(_6116__bF_buf4), .C(_6129_), .Y(_1221_) );
NAND3X1 NAND3X1_948 ( .A(datapath_1_RegisterFile_regfile_mem_24__13_), .B(_5265__bF_buf33), .C(_6116__bF_buf2), .Y(_6130_) );
OAI21X1 OAI21X1_1074 ( .A(_5302__bF_buf2), .B(_6116__bF_buf2), .C(_6130_), .Y(_1222_) );
NAND3X1 NAND3X1_949 ( .A(datapath_1_RegisterFile_regfile_mem_24__14_), .B(_5265__bF_buf59), .C(_6116__bF_buf1), .Y(_6131_) );
OAI21X1 OAI21X1_1075 ( .A(_5304__bF_buf4), .B(_6116__bF_buf1), .C(_6131_), .Y(_1223_) );
NAND3X1 NAND3X1_950 ( .A(datapath_1_RegisterFile_regfile_mem_24__15_), .B(_5265__bF_buf10), .C(_6116__bF_buf7), .Y(_6132_) );
OAI21X1 OAI21X1_1076 ( .A(_5306__bF_buf0), .B(_6116__bF_buf7), .C(_6132_), .Y(_1224_) );
NAND3X1 NAND3X1_951 ( .A(datapath_1_RegisterFile_regfile_mem_24__16_), .B(_5265__bF_buf14), .C(_6116__bF_buf7), .Y(_6133_) );
OAI21X1 OAI21X1_1077 ( .A(_5308__bF_buf3), .B(_6116__bF_buf7), .C(_6133_), .Y(_1806_) );
NAND3X1 NAND3X1_952 ( .A(datapath_1_RegisterFile_regfile_mem_24__17_), .B(_5265__bF_buf28), .C(_6116__bF_buf3), .Y(_6134_) );
OAI21X1 OAI21X1_1078 ( .A(_5310__bF_buf2), .B(_6116__bF_buf3), .C(_6134_), .Y(_1225_) );
NAND3X1 NAND3X1_953 ( .A(datapath_1_RegisterFile_regfile_mem_24__18_), .B(_5265__bF_buf2), .C(_6116__bF_buf2), .Y(_6135_) );
OAI21X1 OAI21X1_1079 ( .A(_5312__bF_buf4), .B(_6116__bF_buf2), .C(_6135_), .Y(_1226_) );
NAND3X1 NAND3X1_954 ( .A(datapath_1_RegisterFile_regfile_mem_24__19_), .B(_5265__bF_buf19), .C(_6116__bF_buf4), .Y(_6136_) );
OAI21X1 OAI21X1_1080 ( .A(_5314__bF_buf0), .B(_6116__bF_buf4), .C(_6136_), .Y(_1807_) );
NAND3X1 NAND3X1_955 ( .A(datapath_1_RegisterFile_regfile_mem_24__20_), .B(_5265__bF_buf9), .C(_6116__bF_buf6), .Y(_6137_) );
OAI21X1 OAI21X1_1081 ( .A(_5316__bF_buf1), .B(_6116__bF_buf6), .C(_6137_), .Y(_1808_) );
NAND3X1 NAND3X1_956 ( .A(datapath_1_RegisterFile_regfile_mem_24__21_), .B(_5265__bF_buf75), .C(_6116__bF_buf0), .Y(_6138_) );
OAI21X1 OAI21X1_1082 ( .A(_5318__bF_buf2), .B(_6116__bF_buf0), .C(_6138_), .Y(_1809_) );
NAND3X1 NAND3X1_957 ( .A(datapath_1_RegisterFile_regfile_mem_24__22_), .B(_5265__bF_buf33), .C(_6116__bF_buf2), .Y(_6139_) );
OAI21X1 OAI21X1_1083 ( .A(_5320__bF_buf0), .B(_6116__bF_buf2), .C(_6139_), .Y(_1810_) );
NAND3X1 NAND3X1_958 ( .A(datapath_1_RegisterFile_regfile_mem_24__23_), .B(_5265__bF_buf75), .C(_6116__bF_buf0), .Y(_6140_) );
OAI21X1 OAI21X1_1084 ( .A(_5322__bF_buf2), .B(_6116__bF_buf0), .C(_6140_), .Y(_1811_) );
NAND3X1 NAND3X1_959 ( .A(datapath_1_RegisterFile_regfile_mem_24__24_), .B(_5265__bF_buf14), .C(_6116__bF_buf7), .Y(_6141_) );
OAI21X1 OAI21X1_1085 ( .A(_5324__bF_buf4), .B(_6116__bF_buf7), .C(_6141_), .Y(_1812_) );
NAND3X1 NAND3X1_960 ( .A(datapath_1_RegisterFile_regfile_mem_24__25_), .B(_5265__bF_buf67), .C(_6116__bF_buf5), .Y(_6142_) );
OAI21X1 OAI21X1_1086 ( .A(_5326__bF_buf3), .B(_6116__bF_buf5), .C(_6142_), .Y(_1813_) );
NAND3X1 NAND3X1_961 ( .A(datapath_1_RegisterFile_regfile_mem_24__26_), .B(_5265__bF_buf12), .C(_6116__bF_buf3), .Y(_6143_) );
OAI21X1 OAI21X1_1087 ( .A(_5328__bF_buf0), .B(_6116__bF_buf3), .C(_6143_), .Y(_1814_) );
NAND3X1 NAND3X1_962 ( .A(datapath_1_RegisterFile_regfile_mem_24__27_), .B(_5265__bF_buf59), .C(_6116__bF_buf1), .Y(_6144_) );
OAI21X1 OAI21X1_1088 ( .A(_5330__bF_buf1), .B(_6116__bF_buf1), .C(_6144_), .Y(_1815_) );
NAND3X1 NAND3X1_963 ( .A(datapath_1_RegisterFile_regfile_mem_24__28_), .B(_5265__bF_buf9), .C(_6116__bF_buf6), .Y(_6145_) );
OAI21X1 OAI21X1_1089 ( .A(_5332__bF_buf0), .B(_6116__bF_buf6), .C(_6145_), .Y(_1816_) );
NAND3X1 NAND3X1_964 ( .A(datapath_1_RegisterFile_regfile_mem_24__29_), .B(_5265__bF_buf63), .C(_6116__bF_buf4), .Y(_6146_) );
OAI21X1 OAI21X1_1090 ( .A(_5334__bF_buf2), .B(_6116__bF_buf4), .C(_6146_), .Y(_1228_) );
NAND3X1 NAND3X1_965 ( .A(datapath_1_RegisterFile_regfile_mem_24__30_), .B(_5265__bF_buf75), .C(_6116__bF_buf0), .Y(_6147_) );
OAI21X1 OAI21X1_1091 ( .A(_5336__bF_buf0), .B(_6116__bF_buf0), .C(_6147_), .Y(_1230_) );
NAND3X1 NAND3X1_966 ( .A(datapath_1_RegisterFile_regfile_mem_24__31_), .B(_5265__bF_buf59), .C(_6116__bF_buf1), .Y(_6148_) );
OAI21X1 OAI21X1_1092 ( .A(_5338__bF_buf1), .B(_6116__bF_buf1), .C(_6148_), .Y(_1231_) );
NAND3X1 NAND3X1_967 ( .A(_6112_), .B(_6114_), .C(_5341_), .Y(_6149_) );
NAND3X1 NAND3X1_968 ( .A(datapath_1_RegisterFile_regfile_mem_25__0_), .B(_5265__bF_buf28), .C(_6149__bF_buf3), .Y(_6150_) );
OAI21X1 OAI21X1_1093 ( .A(_5276__bF_buf1), .B(_6149__bF_buf3), .C(_6150_), .Y(_1238_) );
NAND3X1 NAND3X1_969 ( .A(datapath_1_RegisterFile_regfile_mem_25__1_), .B(_5265__bF_buf53), .C(_6149__bF_buf6), .Y(_6151_) );
OAI21X1 OAI21X1_1094 ( .A(_5278__bF_buf3), .B(_6149__bF_buf6), .C(_6151_), .Y(_1248_) );
NAND3X1 NAND3X1_970 ( .A(datapath_1_RegisterFile_regfile_mem_25__2_), .B(_5265__bF_buf16), .C(_6149__bF_buf4), .Y(_6152_) );
OAI21X1 OAI21X1_1095 ( .A(_5280__bF_buf3), .B(_6149__bF_buf4), .C(_6152_), .Y(_1251_) );
NAND3X1 NAND3X1_971 ( .A(datapath_1_RegisterFile_regfile_mem_25__3_), .B(_5265__bF_buf36), .C(_6149__bF_buf1), .Y(_6153_) );
OAI21X1 OAI21X1_1096 ( .A(_5282__bF_buf2), .B(_6149__bF_buf1), .C(_6153_), .Y(_1252_) );
NAND3X1 NAND3X1_972 ( .A(datapath_1_RegisterFile_regfile_mem_25__4_), .B(_5265__bF_buf53), .C(_6149__bF_buf6), .Y(_6154_) );
OAI21X1 OAI21X1_1097 ( .A(_5284__bF_buf3), .B(_6149__bF_buf6), .C(_6154_), .Y(_1253_) );
NAND3X1 NAND3X1_973 ( .A(datapath_1_RegisterFile_regfile_mem_25__5_), .B(_5265__bF_buf2), .C(_6149__bF_buf2), .Y(_6155_) );
OAI21X1 OAI21X1_1098 ( .A(_5286__bF_buf3), .B(_6149__bF_buf2), .C(_6155_), .Y(_1254_) );
NAND3X1 NAND3X1_974 ( .A(datapath_1_RegisterFile_regfile_mem_25__6_), .B(_5265__bF_buf61), .C(_6149__bF_buf5), .Y(_6156_) );
OAI21X1 OAI21X1_1099 ( .A(_5288__bF_buf0), .B(_6149__bF_buf5), .C(_6156_), .Y(_1255_) );
NAND3X1 NAND3X1_975 ( .A(datapath_1_RegisterFile_regfile_mem_25__7_), .B(_5265__bF_buf36), .C(_6149__bF_buf1), .Y(_6157_) );
OAI21X1 OAI21X1_1100 ( .A(_5290__bF_buf0), .B(_6149__bF_buf1), .C(_6157_), .Y(_1256_) );
NAND3X1 NAND3X1_976 ( .A(datapath_1_RegisterFile_regfile_mem_25__8_), .B(_5265__bF_buf95), .C(_6149__bF_buf6), .Y(_6158_) );
OAI21X1 OAI21X1_1101 ( .A(_5292__bF_buf4), .B(_6149__bF_buf6), .C(_6158_), .Y(_1257_) );
NAND3X1 NAND3X1_977 ( .A(datapath_1_RegisterFile_regfile_mem_25__9_), .B(_5265__bF_buf12), .C(_6149__bF_buf7), .Y(_6159_) );
OAI21X1 OAI21X1_1102 ( .A(_5294__bF_buf0), .B(_6149__bF_buf7), .C(_6159_), .Y(_1817_) );
NAND3X1 NAND3X1_978 ( .A(datapath_1_RegisterFile_regfile_mem_25__10_), .B(_5265__bF_buf31), .C(_6149__bF_buf7), .Y(_6160_) );
OAI21X1 OAI21X1_1103 ( .A(_5296__bF_buf1), .B(_6149__bF_buf7), .C(_6160_), .Y(_1239_) );
NAND3X1 NAND3X1_979 ( .A(datapath_1_RegisterFile_regfile_mem_25__11_), .B(_5265__bF_buf3), .C(_6149__bF_buf0), .Y(_6161_) );
OAI21X1 OAI21X1_1104 ( .A(_5298__bF_buf0), .B(_6149__bF_buf0), .C(_6161_), .Y(_1240_) );
NAND3X1 NAND3X1_980 ( .A(datapath_1_RegisterFile_regfile_mem_25__12_), .B(_5265__bF_buf63), .C(_6149__bF_buf0), .Y(_6162_) );
OAI21X1 OAI21X1_1105 ( .A(_5300__bF_buf0), .B(_6149__bF_buf0), .C(_6162_), .Y(_1241_) );
NAND3X1 NAND3X1_981 ( .A(datapath_1_RegisterFile_regfile_mem_25__13_), .B(_5265__bF_buf33), .C(_6149__bF_buf5), .Y(_6163_) );
OAI21X1 OAI21X1_1106 ( .A(_5302__bF_buf3), .B(_6149__bF_buf5), .C(_6163_), .Y(_1242_) );
NAND3X1 NAND3X1_982 ( .A(datapath_1_RegisterFile_regfile_mem_25__14_), .B(_5265__bF_buf2), .C(_6149__bF_buf2), .Y(_6164_) );
OAI21X1 OAI21X1_1107 ( .A(_5304__bF_buf4), .B(_6149__bF_buf2), .C(_6164_), .Y(_1243_) );
NAND3X1 NAND3X1_983 ( .A(datapath_1_RegisterFile_regfile_mem_25__15_), .B(_5265__bF_buf3), .C(_6149__bF_buf0), .Y(_6165_) );
OAI21X1 OAI21X1_1108 ( .A(_5306__bF_buf4), .B(_6149__bF_buf0), .C(_6165_), .Y(_1244_) );
NAND3X1 NAND3X1_984 ( .A(datapath_1_RegisterFile_regfile_mem_25__16_), .B(_5265__bF_buf41), .C(_6149__bF_buf4), .Y(_6166_) );
OAI21X1 OAI21X1_1109 ( .A(_5308__bF_buf4), .B(_6149__bF_buf4), .C(_6166_), .Y(_1245_) );
NAND3X1 NAND3X1_985 ( .A(datapath_1_RegisterFile_regfile_mem_25__17_), .B(_5265__bF_buf8), .C(_6149__bF_buf5), .Y(_6167_) );
OAI21X1 OAI21X1_1110 ( .A(_5310__bF_buf3), .B(_6149__bF_buf5), .C(_6167_), .Y(_1246_) );
NAND3X1 NAND3X1_986 ( .A(datapath_1_RegisterFile_regfile_mem_25__18_), .B(_5265__bF_buf2), .C(_6149__bF_buf2), .Y(_6168_) );
OAI21X1 OAI21X1_1111 ( .A(_5312__bF_buf4), .B(_6149__bF_buf2), .C(_6168_), .Y(_1247_) );
NAND3X1 NAND3X1_987 ( .A(datapath_1_RegisterFile_regfile_mem_25__19_), .B(_5265__bF_buf63), .C(_6149__bF_buf0), .Y(_6169_) );
OAI21X1 OAI21X1_1112 ( .A(_5314__bF_buf0), .B(_6149__bF_buf0), .C(_6169_), .Y(_1818_) );
NAND3X1 NAND3X1_988 ( .A(datapath_1_RegisterFile_regfile_mem_25__20_), .B(_5265__bF_buf30), .C(_6149__bF_buf1), .Y(_6170_) );
OAI21X1 OAI21X1_1113 ( .A(_5316__bF_buf1), .B(_6149__bF_buf1), .C(_6170_), .Y(_1249_) );
NAND3X1 NAND3X1_989 ( .A(datapath_1_RegisterFile_regfile_mem_25__21_), .B(_5265__bF_buf75), .C(_6149__bF_buf3), .Y(_6171_) );
OAI21X1 OAI21X1_1114 ( .A(_5318__bF_buf3), .B(_6149__bF_buf3), .C(_6171_), .Y(_1250_) );
NAND3X1 NAND3X1_990 ( .A(datapath_1_RegisterFile_regfile_mem_25__22_), .B(_5265__bF_buf33), .C(_6149__bF_buf7), .Y(_6172_) );
OAI21X1 OAI21X1_1115 ( .A(_5320__bF_buf3), .B(_6149__bF_buf7), .C(_6172_), .Y(_1819_) );
NAND3X1 NAND3X1_991 ( .A(datapath_1_RegisterFile_regfile_mem_25__23_), .B(_5265__bF_buf75), .C(_6149__bF_buf3), .Y(_6173_) );
OAI21X1 OAI21X1_1116 ( .A(_5322__bF_buf2), .B(_6149__bF_buf3), .C(_6173_), .Y(_1820_) );
NAND3X1 NAND3X1_992 ( .A(datapath_1_RegisterFile_regfile_mem_25__24_), .B(_5265__bF_buf34), .C(_6149__bF_buf4), .Y(_6174_) );
OAI21X1 OAI21X1_1117 ( .A(_5324__bF_buf2), .B(_6149__bF_buf4), .C(_6174_), .Y(_1821_) );
NAND3X1 NAND3X1_993 ( .A(datapath_1_RegisterFile_regfile_mem_25__25_), .B(_5265__bF_buf95), .C(_6149__bF_buf6), .Y(_6175_) );
OAI21X1 OAI21X1_1118 ( .A(_5326__bF_buf3), .B(_6149__bF_buf6), .C(_6175_), .Y(_1822_) );
NAND3X1 NAND3X1_994 ( .A(datapath_1_RegisterFile_regfile_mem_25__26_), .B(_5265__bF_buf33), .C(_6149__bF_buf5), .Y(_6176_) );
OAI21X1 OAI21X1_1119 ( .A(_5328__bF_buf4), .B(_6149__bF_buf5), .C(_6176_), .Y(_1823_) );
NAND3X1 NAND3X1_995 ( .A(datapath_1_RegisterFile_regfile_mem_25__27_), .B(_5265__bF_buf2), .C(_6149__bF_buf2), .Y(_6177_) );
OAI21X1 OAI21X1_1120 ( .A(_5330__bF_buf1), .B(_6149__bF_buf2), .C(_6177_), .Y(_1824_) );
NAND3X1 NAND3X1_996 ( .A(datapath_1_RegisterFile_regfile_mem_25__28_), .B(_5265__bF_buf36), .C(_6149__bF_buf1), .Y(_6178_) );
OAI21X1 OAI21X1_1121 ( .A(_5332__bF_buf0), .B(_6149__bF_buf1), .C(_6178_), .Y(_1825_) );
NAND3X1 NAND3X1_997 ( .A(datapath_1_RegisterFile_regfile_mem_25__29_), .B(_5265__bF_buf24), .C(_6149__bF_buf4), .Y(_6179_) );
OAI21X1 OAI21X1_1122 ( .A(_5334__bF_buf3), .B(_6149__bF_buf4), .C(_6179_), .Y(_1826_) );
NAND3X1 NAND3X1_998 ( .A(datapath_1_RegisterFile_regfile_mem_25__30_), .B(_5265__bF_buf28), .C(_6149__bF_buf3), .Y(_6180_) );
OAI21X1 OAI21X1_1123 ( .A(_5336__bF_buf0), .B(_6149__bF_buf3), .C(_6180_), .Y(_1827_) );
NAND3X1 NAND3X1_999 ( .A(datapath_1_RegisterFile_regfile_mem_25__31_), .B(_5265__bF_buf22), .C(_6149__bF_buf7), .Y(_6181_) );
OAI21X1 OAI21X1_1124 ( .A(_5338__bF_buf4), .B(_6149__bF_buf7), .C(_6181_), .Y(_1828_) );
NAND3X1 NAND3X1_1000 ( .A(_6112_), .B(_6114_), .C(_5376_), .Y(_6182_) );
NAND3X1 NAND3X1_1001 ( .A(datapath_1_RegisterFile_regfile_mem_26__0_), .B(_5265__bF_buf75), .C(_6182__bF_buf7), .Y(_6183_) );
OAI21X1 OAI21X1_1125 ( .A(_5276__bF_buf1), .B(_6182__bF_buf7), .C(_6183_), .Y(_1258_) );
NAND3X1 NAND3X1_1002 ( .A(datapath_1_RegisterFile_regfile_mem_26__1_), .B(_5265__bF_buf53), .C(_6182__bF_buf1), .Y(_6184_) );
OAI21X1 OAI21X1_1126 ( .A(_5278__bF_buf3), .B(_6182__bF_buf1), .C(_6184_), .Y(_1268_) );
NAND3X1 NAND3X1_1003 ( .A(datapath_1_RegisterFile_regfile_mem_26__2_), .B(_5265__bF_buf20), .C(_6182__bF_buf6), .Y(_6185_) );
OAI21X1 OAI21X1_1127 ( .A(_5280__bF_buf4), .B(_6182__bF_buf6), .C(_6185_), .Y(_1278_) );
NAND3X1 NAND3X1_1004 ( .A(datapath_1_RegisterFile_regfile_mem_26__3_), .B(_5265__bF_buf10), .C(_6182__bF_buf5), .Y(_6186_) );
OAI21X1 OAI21X1_1128 ( .A(_5282__bF_buf3), .B(_6182__bF_buf5), .C(_6186_), .Y(_1281_) );
NAND3X1 NAND3X1_1005 ( .A(datapath_1_RegisterFile_regfile_mem_26__4_), .B(_5265__bF_buf54), .C(_6182__bF_buf2), .Y(_6187_) );
OAI21X1 OAI21X1_1129 ( .A(_5284__bF_buf0), .B(_6182__bF_buf2), .C(_6187_), .Y(_1829_) );
NAND3X1 NAND3X1_1006 ( .A(datapath_1_RegisterFile_regfile_mem_26__5_), .B(_5265__bF_buf2), .C(_6182__bF_buf4), .Y(_6188_) );
OAI21X1 OAI21X1_1130 ( .A(_5286__bF_buf3), .B(_6182__bF_buf4), .C(_6188_), .Y(_1282_) );
NAND3X1 NAND3X1_1007 ( .A(datapath_1_RegisterFile_regfile_mem_26__6_), .B(_5265__bF_buf4), .C(_6182__bF_buf1), .Y(_6189_) );
OAI21X1 OAI21X1_1131 ( .A(_5288__bF_buf0), .B(_6182__bF_buf1), .C(_6189_), .Y(_1283_) );
NAND3X1 NAND3X1_1008 ( .A(datapath_1_RegisterFile_regfile_mem_26__7_), .B(_5265__bF_buf89), .C(_6182__bF_buf3), .Y(_6190_) );
OAI21X1 OAI21X1_1132 ( .A(_5290__bF_buf3), .B(_6182__bF_buf3), .C(_6190_), .Y(_1284_) );
NAND3X1 NAND3X1_1009 ( .A(datapath_1_RegisterFile_regfile_mem_26__8_), .B(_5265__bF_buf95), .C(_6182__bF_buf1), .Y(_6191_) );
OAI21X1 OAI21X1_1133 ( .A(_5292__bF_buf4), .B(_6182__bF_buf1), .C(_6191_), .Y(_1285_) );
NAND3X1 NAND3X1_1010 ( .A(datapath_1_RegisterFile_regfile_mem_26__9_), .B(_5265__bF_buf12), .C(_6182__bF_buf7), .Y(_6192_) );
OAI21X1 OAI21X1_1134 ( .A(_5294__bF_buf0), .B(_6182__bF_buf7), .C(_6192_), .Y(_1286_) );
NAND3X1 NAND3X1_1011 ( .A(datapath_1_RegisterFile_regfile_mem_26__10_), .B(_5265__bF_buf12), .C(_6182__bF_buf7), .Y(_6193_) );
OAI21X1 OAI21X1_1135 ( .A(_5296__bF_buf3), .B(_6182__bF_buf7), .C(_6193_), .Y(_1259_) );
NAND3X1 NAND3X1_1012 ( .A(datapath_1_RegisterFile_regfile_mem_26__11_), .B(_5265__bF_buf3), .C(_6182__bF_buf5), .Y(_6194_) );
OAI21X1 OAI21X1_1136 ( .A(_5298__bF_buf4), .B(_6182__bF_buf5), .C(_6194_), .Y(_1260_) );
NAND3X1 NAND3X1_1013 ( .A(datapath_1_RegisterFile_regfile_mem_26__12_), .B(_5265__bF_buf3), .C(_6182__bF_buf3), .Y(_6195_) );
OAI21X1 OAI21X1_1137 ( .A(_5300__bF_buf0), .B(_6182__bF_buf3), .C(_6195_), .Y(_1261_) );
NAND3X1 NAND3X1_1014 ( .A(datapath_1_RegisterFile_regfile_mem_26__13_), .B(_5265__bF_buf1), .C(_6182__bF_buf0), .Y(_6196_) );
OAI21X1 OAI21X1_1138 ( .A(_5302__bF_buf3), .B(_6182__bF_buf0), .C(_6196_), .Y(_1262_) );
NAND3X1 NAND3X1_1015 ( .A(datapath_1_RegisterFile_regfile_mem_26__14_), .B(_5265__bF_buf59), .C(_6182__bF_buf4), .Y(_6197_) );
OAI21X1 OAI21X1_1139 ( .A(_5304__bF_buf4), .B(_6182__bF_buf4), .C(_6197_), .Y(_1830_) );
NAND3X1 NAND3X1_1016 ( .A(datapath_1_RegisterFile_regfile_mem_26__15_), .B(_5265__bF_buf20), .C(_6182__bF_buf3), .Y(_6198_) );
OAI21X1 OAI21X1_1140 ( .A(_5306__bF_buf4), .B(_6182__bF_buf3), .C(_6198_), .Y(_1263_) );
NAND3X1 NAND3X1_1017 ( .A(datapath_1_RegisterFile_regfile_mem_26__16_), .B(_5265__bF_buf40), .C(_6182__bF_buf6), .Y(_6199_) );
OAI21X1 OAI21X1_1141 ( .A(_5308__bF_buf3), .B(_6182__bF_buf6), .C(_6199_), .Y(_1264_) );
NAND3X1 NAND3X1_1018 ( .A(datapath_1_RegisterFile_regfile_mem_26__17_), .B(_5265__bF_buf49), .C(_6182__bF_buf2), .Y(_6200_) );
OAI21X1 OAI21X1_1142 ( .A(_5310__bF_buf0), .B(_6182__bF_buf2), .C(_6200_), .Y(_1265_) );
NAND3X1 NAND3X1_1019 ( .A(datapath_1_RegisterFile_regfile_mem_26__18_), .B(_5265__bF_buf58), .C(_6182__bF_buf0), .Y(_6201_) );
OAI21X1 OAI21X1_1143 ( .A(_5312__bF_buf4), .B(_6182__bF_buf0), .C(_6201_), .Y(_1266_) );
NAND3X1 NAND3X1_1020 ( .A(datapath_1_RegisterFile_regfile_mem_26__19_), .B(_5265__bF_buf20), .C(_6182__bF_buf6), .Y(_6202_) );
OAI21X1 OAI21X1_1144 ( .A(_5314__bF_buf2), .B(_6182__bF_buf6), .C(_6202_), .Y(_1267_) );
NAND3X1 NAND3X1_1021 ( .A(datapath_1_RegisterFile_regfile_mem_26__20_), .B(_5265__bF_buf9), .C(_6182__bF_buf5), .Y(_6203_) );
OAI21X1 OAI21X1_1145 ( .A(_5316__bF_buf0), .B(_6182__bF_buf5), .C(_6203_), .Y(_1269_) );
NAND3X1 NAND3X1_1022 ( .A(datapath_1_RegisterFile_regfile_mem_26__21_), .B(_5265__bF_buf8), .C(_6182__bF_buf2), .Y(_6204_) );
OAI21X1 OAI21X1_1146 ( .A(_5318__bF_buf3), .B(_6182__bF_buf2), .C(_6204_), .Y(_1270_) );
NAND3X1 NAND3X1_1023 ( .A(datapath_1_RegisterFile_regfile_mem_26__22_), .B(_5265__bF_buf79), .C(_6182__bF_buf0), .Y(_6205_) );
OAI21X1 OAI21X1_1147 ( .A(_5320__bF_buf0), .B(_6182__bF_buf0), .C(_6205_), .Y(_1271_) );
NAND3X1 NAND3X1_1024 ( .A(datapath_1_RegisterFile_regfile_mem_26__23_), .B(_5265__bF_buf12), .C(_6182__bF_buf7), .Y(_6206_) );
OAI21X1 OAI21X1_1148 ( .A(_5322__bF_buf2), .B(_6182__bF_buf7), .C(_6206_), .Y(_1272_) );
NAND3X1 NAND3X1_1025 ( .A(datapath_1_RegisterFile_regfile_mem_26__24_), .B(_5265__bF_buf78), .C(_6182__bF_buf6), .Y(_6207_) );
OAI21X1 OAI21X1_1149 ( .A(_5324__bF_buf4), .B(_6182__bF_buf6), .C(_6207_), .Y(_1831_) );
NAND3X1 NAND3X1_1026 ( .A(datapath_1_RegisterFile_regfile_mem_26__25_), .B(_5265__bF_buf80), .C(_6182__bF_buf1), .Y(_6208_) );
OAI21X1 OAI21X1_1150 ( .A(_5326__bF_buf3), .B(_6182__bF_buf1), .C(_6208_), .Y(_1273_) );
NAND3X1 NAND3X1_1027 ( .A(datapath_1_RegisterFile_regfile_mem_26__26_), .B(_5265__bF_buf79), .C(_6182__bF_buf0), .Y(_6209_) );
OAI21X1 OAI21X1_1151 ( .A(_5328__bF_buf4), .B(_6182__bF_buf0), .C(_6209_), .Y(_1274_) );
NAND3X1 NAND3X1_1028 ( .A(datapath_1_RegisterFile_regfile_mem_26__27_), .B(_5265__bF_buf2), .C(_6182__bF_buf4), .Y(_6210_) );
OAI21X1 OAI21X1_1152 ( .A(_5330__bF_buf1), .B(_6182__bF_buf4), .C(_6210_), .Y(_1275_) );
NAND3X1 NAND3X1_1029 ( .A(datapath_1_RegisterFile_regfile_mem_26__28_), .B(_5265__bF_buf9), .C(_6182__bF_buf5), .Y(_6211_) );
OAI21X1 OAI21X1_1153 ( .A(_5332__bF_buf0), .B(_6182__bF_buf5), .C(_6211_), .Y(_1276_) );
NAND3X1 NAND3X1_1030 ( .A(datapath_1_RegisterFile_regfile_mem_26__29_), .B(_5265__bF_buf20), .C(_6182__bF_buf3), .Y(_6212_) );
OAI21X1 OAI21X1_1154 ( .A(_5334__bF_buf2), .B(_6182__bF_buf3), .C(_6212_), .Y(_1277_) );
NAND3X1 NAND3X1_1031 ( .A(datapath_1_RegisterFile_regfile_mem_26__30_), .B(_5265__bF_buf49), .C(_6182__bF_buf2), .Y(_6213_) );
OAI21X1 OAI21X1_1155 ( .A(_5336__bF_buf3), .B(_6182__bF_buf2), .C(_6213_), .Y(_1279_) );
NAND3X1 NAND3X1_1032 ( .A(datapath_1_RegisterFile_regfile_mem_26__31_), .B(_5265__bF_buf59), .C(_6182__bF_buf4), .Y(_6214_) );
OAI21X1 OAI21X1_1156 ( .A(_5338__bF_buf1), .B(_6182__bF_buf4), .C(_6214_), .Y(_1280_) );
NAND3X1 NAND3X1_1033 ( .A(_6112_), .B(_5410_), .C(_6114_), .Y(_6215_) );
NAND3X1 NAND3X1_1034 ( .A(datapath_1_RegisterFile_regfile_mem_27__0_), .B(_5265__bF_buf75), .C(_6215__bF_buf5), .Y(_6216_) );
OAI21X1 OAI21X1_1157 ( .A(_5276__bF_buf1), .B(_6215__bF_buf5), .C(_6216_), .Y(_1832_) );
NAND3X1 NAND3X1_1035 ( .A(datapath_1_RegisterFile_regfile_mem_27__1_), .B(_5265__bF_buf53), .C(_6215__bF_buf2), .Y(_6217_) );
OAI21X1 OAI21X1_1158 ( .A(_5278__bF_buf3), .B(_6215__bF_buf2), .C(_6217_), .Y(_1833_) );
NAND3X1 NAND3X1_1036 ( .A(datapath_1_RegisterFile_regfile_mem_27__2_), .B(_5265__bF_buf20), .C(_6215__bF_buf7), .Y(_6218_) );
OAI21X1 OAI21X1_1159 ( .A(_5280__bF_buf4), .B(_6215__bF_buf7), .C(_6218_), .Y(_1305_) );
NAND3X1 NAND3X1_1037 ( .A(datapath_1_RegisterFile_regfile_mem_27__3_), .B(_5265__bF_buf10), .C(_6215__bF_buf3), .Y(_6219_) );
OAI21X1 OAI21X1_1160 ( .A(_5282__bF_buf3), .B(_6215__bF_buf3), .C(_6219_), .Y(_1308_) );
NAND3X1 NAND3X1_1038 ( .A(datapath_1_RegisterFile_regfile_mem_27__4_), .B(_5265__bF_buf46), .C(_6215__bF_buf2), .Y(_6220_) );
OAI21X1 OAI21X1_1161 ( .A(_5284__bF_buf3), .B(_6215__bF_buf2), .C(_6220_), .Y(_1309_) );
NAND3X1 NAND3X1_1039 ( .A(datapath_1_RegisterFile_regfile_mem_27__5_), .B(_5265__bF_buf2), .C(_6215__bF_buf0), .Y(_6221_) );
OAI21X1 OAI21X1_1162 ( .A(_5286__bF_buf3), .B(_6215__bF_buf0), .C(_6221_), .Y(_1310_) );
NAND3X1 NAND3X1_1040 ( .A(datapath_1_RegisterFile_regfile_mem_27__6_), .B(_5265__bF_buf4), .C(_6215__bF_buf5), .Y(_6222_) );
OAI21X1 OAI21X1_1163 ( .A(_5288__bF_buf4), .B(_6215__bF_buf5), .C(_6222_), .Y(_1311_) );
NAND3X1 NAND3X1_1041 ( .A(datapath_1_RegisterFile_regfile_mem_27__7_), .B(_5265__bF_buf9), .C(_6215__bF_buf3), .Y(_6223_) );
OAI21X1 OAI21X1_1164 ( .A(_5290__bF_buf0), .B(_6215__bF_buf3), .C(_6223_), .Y(_1312_) );
NAND3X1 NAND3X1_1042 ( .A(datapath_1_RegisterFile_regfile_mem_27__8_), .B(_5265__bF_buf67), .C(_6215__bF_buf2), .Y(_6224_) );
OAI21X1 OAI21X1_1165 ( .A(_5292__bF_buf0), .B(_6215__bF_buf2), .C(_6224_), .Y(_1313_) );
NAND3X1 NAND3X1_1043 ( .A(datapath_1_RegisterFile_regfile_mem_27__9_), .B(_5265__bF_buf90), .C(_6215__bF_buf1), .Y(_6225_) );
OAI21X1 OAI21X1_1166 ( .A(_5294__bF_buf4), .B(_6215__bF_buf1), .C(_6225_), .Y(_1834_) );
NAND3X1 NAND3X1_1044 ( .A(datapath_1_RegisterFile_regfile_mem_27__10_), .B(_5265__bF_buf31), .C(_6215__bF_buf1), .Y(_6226_) );
OAI21X1 OAI21X1_1167 ( .A(_5296__bF_buf1), .B(_6215__bF_buf1), .C(_6226_), .Y(_1287_) );
NAND3X1 NAND3X1_1045 ( .A(datapath_1_RegisterFile_regfile_mem_27__11_), .B(_5265__bF_buf69), .C(_6215__bF_buf6), .Y(_6227_) );
OAI21X1 OAI21X1_1168 ( .A(_5298__bF_buf4), .B(_6215__bF_buf6), .C(_6227_), .Y(_1288_) );
NAND3X1 NAND3X1_1046 ( .A(datapath_1_RegisterFile_regfile_mem_27__12_), .B(_5265__bF_buf3), .C(_6215__bF_buf7), .Y(_6228_) );
OAI21X1 OAI21X1_1169 ( .A(_5300__bF_buf0), .B(_6215__bF_buf7), .C(_6228_), .Y(_1289_) );
NAND3X1 NAND3X1_1047 ( .A(datapath_1_RegisterFile_regfile_mem_27__13_), .B(_5265__bF_buf47), .C(_6215__bF_buf4), .Y(_6229_) );
OAI21X1 OAI21X1_1170 ( .A(_5302__bF_buf3), .B(_6215__bF_buf4), .C(_6229_), .Y(_1290_) );
NAND3X1 NAND3X1_1048 ( .A(datapath_1_RegisterFile_regfile_mem_27__14_), .B(_5265__bF_buf22), .C(_6215__bF_buf1), .Y(_6230_) );
OAI21X1 OAI21X1_1171 ( .A(_5304__bF_buf4), .B(_6215__bF_buf1), .C(_6230_), .Y(_1291_) );
NAND3X1 NAND3X1_1049 ( .A(datapath_1_RegisterFile_regfile_mem_27__15_), .B(_5265__bF_buf3), .C(_6215__bF_buf7), .Y(_6231_) );
OAI21X1 OAI21X1_1172 ( .A(_5306__bF_buf4), .B(_6215__bF_buf7), .C(_6231_), .Y(_1292_) );
NAND3X1 NAND3X1_1050 ( .A(datapath_1_RegisterFile_regfile_mem_27__16_), .B(_5265__bF_buf40), .C(_6215__bF_buf6), .Y(_6232_) );
OAI21X1 OAI21X1_1173 ( .A(_5308__bF_buf3), .B(_6215__bF_buf6), .C(_6232_), .Y(_1293_) );
NAND3X1 NAND3X1_1051 ( .A(datapath_1_RegisterFile_regfile_mem_27__17_), .B(_5265__bF_buf66), .C(_6215__bF_buf4), .Y(_6233_) );
OAI21X1 OAI21X1_1174 ( .A(_5310__bF_buf0), .B(_6215__bF_buf4), .C(_6233_), .Y(_1294_) );
NAND3X1 NAND3X1_1052 ( .A(datapath_1_RegisterFile_regfile_mem_27__18_), .B(_5265__bF_buf2), .C(_6215__bF_buf0), .Y(_6234_) );
OAI21X1 OAI21X1_1175 ( .A(_5312__bF_buf4), .B(_6215__bF_buf0), .C(_6234_), .Y(_1295_) );
NAND3X1 NAND3X1_1053 ( .A(datapath_1_RegisterFile_regfile_mem_27__19_), .B(_5265__bF_buf55), .C(_6215__bF_buf5), .Y(_6235_) );
OAI21X1 OAI21X1_1176 ( .A(_5314__bF_buf0), .B(_6215__bF_buf5), .C(_6235_), .Y(_1835_) );
NAND3X1 NAND3X1_1054 ( .A(datapath_1_RegisterFile_regfile_mem_27__20_), .B(_5265__bF_buf9), .C(_6215__bF_buf3), .Y(_6236_) );
OAI21X1 OAI21X1_1177 ( .A(_5316__bF_buf0), .B(_6215__bF_buf3), .C(_6236_), .Y(_1296_) );
NAND3X1 NAND3X1_1055 ( .A(datapath_1_RegisterFile_regfile_mem_27__21_), .B(_5265__bF_buf54), .C(_6215__bF_buf2), .Y(_6237_) );
OAI21X1 OAI21X1_1178 ( .A(_5318__bF_buf1), .B(_6215__bF_buf2), .C(_6237_), .Y(_1297_) );
NAND3X1 NAND3X1_1056 ( .A(datapath_1_RegisterFile_regfile_mem_27__22_), .B(_5265__bF_buf58), .C(_6215__bF_buf0), .Y(_6238_) );
OAI21X1 OAI21X1_1179 ( .A(_5320__bF_buf3), .B(_6215__bF_buf0), .C(_6238_), .Y(_1298_) );
NAND3X1 NAND3X1_1057 ( .A(datapath_1_RegisterFile_regfile_mem_27__23_), .B(_5265__bF_buf4), .C(_6215__bF_buf5), .Y(_6239_) );
OAI21X1 OAI21X1_1180 ( .A(_5322__bF_buf0), .B(_6215__bF_buf5), .C(_6239_), .Y(_1299_) );
NAND3X1 NAND3X1_1058 ( .A(datapath_1_RegisterFile_regfile_mem_27__24_), .B(_5265__bF_buf71), .C(_6215__bF_buf6), .Y(_6240_) );
OAI21X1 OAI21X1_1181 ( .A(_5324__bF_buf1), .B(_6215__bF_buf6), .C(_6240_), .Y(_1300_) );
NAND3X1 NAND3X1_1059 ( .A(datapath_1_RegisterFile_regfile_mem_27__25_), .B(_5265__bF_buf41), .C(_6215__bF_buf6), .Y(_6241_) );
OAI21X1 OAI21X1_1182 ( .A(_5326__bF_buf4), .B(_6215__bF_buf6), .C(_6241_), .Y(_1301_) );
NAND3X1 NAND3X1_1060 ( .A(datapath_1_RegisterFile_regfile_mem_27__26_), .B(_5265__bF_buf66), .C(_6215__bF_buf4), .Y(_6242_) );
OAI21X1 OAI21X1_1183 ( .A(_5328__bF_buf1), .B(_6215__bF_buf4), .C(_6242_), .Y(_1302_) );
NAND3X1 NAND3X1_1061 ( .A(datapath_1_RegisterFile_regfile_mem_27__27_), .B(_5265__bF_buf59), .C(_6215__bF_buf0), .Y(_6243_) );
OAI21X1 OAI21X1_1184 ( .A(_5330__bF_buf1), .B(_6215__bF_buf0), .C(_6243_), .Y(_1303_) );
NAND3X1 NAND3X1_1062 ( .A(datapath_1_RegisterFile_regfile_mem_27__28_), .B(_5265__bF_buf9), .C(_6215__bF_buf3), .Y(_6244_) );
OAI21X1 OAI21X1_1185 ( .A(_5332__bF_buf3), .B(_6215__bF_buf3), .C(_6244_), .Y(_1304_) );
NAND3X1 NAND3X1_1063 ( .A(datapath_1_RegisterFile_regfile_mem_27__29_), .B(_5265__bF_buf3), .C(_6215__bF_buf7), .Y(_6245_) );
OAI21X1 OAI21X1_1186 ( .A(_5334__bF_buf2), .B(_6215__bF_buf7), .C(_6245_), .Y(_1836_) );
NAND3X1 NAND3X1_1064 ( .A(datapath_1_RegisterFile_regfile_mem_27__30_), .B(_5265__bF_buf66), .C(_6215__bF_buf4), .Y(_6246_) );
OAI21X1 OAI21X1_1187 ( .A(_5336__bF_buf3), .B(_6215__bF_buf4), .C(_6246_), .Y(_1306_) );
NAND3X1 NAND3X1_1065 ( .A(datapath_1_RegisterFile_regfile_mem_27__31_), .B(_5265__bF_buf22), .C(_6215__bF_buf1), .Y(_6247_) );
OAI21X1 OAI21X1_1188 ( .A(_5338__bF_buf1), .B(_6215__bF_buf1), .C(_6247_), .Y(_1307_) );
AOI21X1 AOI21X1_312 ( .A(datapath_1_A3_3_), .B(datapath_1_A3_4_), .C(_5266_), .Y(_6248_) );
NOR2X1 NOR2X1_141 ( .A(_6248_), .B(_6112_), .Y(_6249_) );
NAND2X1 NAND2X1_389 ( .A(_6249_), .B(_5274_), .Y(_6250_) );
NAND3X1 NAND3X1_1066 ( .A(datapath_1_RegisterFile_regfile_mem_28__0_), .B(_5265__bF_buf90), .C(_6250__bF_buf2), .Y(_6251_) );
OAI21X1 OAI21X1_1189 ( .A(_5276__bF_buf3), .B(_6250__bF_buf2), .C(_6251_), .Y(_1314_) );
NAND3X1 NAND3X1_1067 ( .A(datapath_1_RegisterFile_regfile_mem_28__1_), .B(_5265__bF_buf95), .C(_6250__bF_buf0), .Y(_6252_) );
OAI21X1 OAI21X1_1190 ( .A(_5278__bF_buf4), .B(_6250__bF_buf0), .C(_6252_), .Y(_1324_) );
NAND3X1 NAND3X1_1068 ( .A(datapath_1_RegisterFile_regfile_mem_28__2_), .B(_5265__bF_buf20), .C(_6250__bF_buf1), .Y(_6253_) );
OAI21X1 OAI21X1_1191 ( .A(_5280__bF_buf4), .B(_6250__bF_buf1), .C(_6253_), .Y(_1331_) );
NAND3X1 NAND3X1_1069 ( .A(datapath_1_RegisterFile_regfile_mem_28__3_), .B(_5265__bF_buf10), .C(_6250__bF_buf4), .Y(_6254_) );
OAI21X1 OAI21X1_1192 ( .A(_5282__bF_buf3), .B(_6250__bF_buf4), .C(_6254_), .Y(_1332_) );
NAND3X1 NAND3X1_1070 ( .A(datapath_1_RegisterFile_regfile_mem_28__4_), .B(_5265__bF_buf53), .C(_6250__bF_buf0), .Y(_6255_) );
OAI21X1 OAI21X1_1193 ( .A(_5284__bF_buf3), .B(_6250__bF_buf0), .C(_6255_), .Y(_1837_) );
NAND3X1 NAND3X1_1071 ( .A(datapath_1_RegisterFile_regfile_mem_28__5_), .B(_5265__bF_buf22), .C(_6250__bF_buf6), .Y(_6256_) );
OAI21X1 OAI21X1_1194 ( .A(_5286__bF_buf4), .B(_6250__bF_buf6), .C(_6256_), .Y(_1333_) );
NAND3X1 NAND3X1_1072 ( .A(datapath_1_RegisterFile_regfile_mem_28__6_), .B(_5265__bF_buf61), .C(_6250__bF_buf3), .Y(_6257_) );
OAI21X1 OAI21X1_1195 ( .A(_5288__bF_buf0), .B(_6250__bF_buf3), .C(_6257_), .Y(_1334_) );
NAND3X1 NAND3X1_1073 ( .A(datapath_1_RegisterFile_regfile_mem_28__7_), .B(_5265__bF_buf36), .C(_6250__bF_buf5), .Y(_6258_) );
OAI21X1 OAI21X1_1196 ( .A(_5290__bF_buf3), .B(_6250__bF_buf5), .C(_6258_), .Y(_1335_) );
NAND3X1 NAND3X1_1074 ( .A(datapath_1_RegisterFile_regfile_mem_28__8_), .B(_5265__bF_buf49), .C(_6250__bF_buf3), .Y(_6259_) );
OAI21X1 OAI21X1_1197 ( .A(_5292__bF_buf2), .B(_6250__bF_buf3), .C(_6259_), .Y(_1336_) );
NAND3X1 NAND3X1_1075 ( .A(datapath_1_RegisterFile_regfile_mem_28__9_), .B(_5265__bF_buf12), .C(_6250__bF_buf2), .Y(_6260_) );
OAI21X1 OAI21X1_1198 ( .A(_5294__bF_buf0), .B(_6250__bF_buf2), .C(_6260_), .Y(_1337_) );
NAND3X1 NAND3X1_1076 ( .A(datapath_1_RegisterFile_regfile_mem_28__10_), .B(_5265__bF_buf90), .C(_6250__bF_buf2), .Y(_6261_) );
OAI21X1 OAI21X1_1199 ( .A(_5296__bF_buf3), .B(_6250__bF_buf2), .C(_6261_), .Y(_1315_) );
NAND3X1 NAND3X1_1077 ( .A(datapath_1_RegisterFile_regfile_mem_28__11_), .B(_5265__bF_buf9), .C(_6250__bF_buf5), .Y(_6262_) );
OAI21X1 OAI21X1_1200 ( .A(_5298__bF_buf4), .B(_6250__bF_buf5), .C(_6262_), .Y(_1316_) );
NAND3X1 NAND3X1_1078 ( .A(datapath_1_RegisterFile_regfile_mem_28__12_), .B(_5265__bF_buf3), .C(_6250__bF_buf5), .Y(_6263_) );
OAI21X1 OAI21X1_1201 ( .A(_5300__bF_buf0), .B(_6250__bF_buf5), .C(_6263_), .Y(_1317_) );
NAND3X1 NAND3X1_1079 ( .A(datapath_1_RegisterFile_regfile_mem_28__13_), .B(_5265__bF_buf33), .C(_6250__bF_buf6), .Y(_6264_) );
OAI21X1 OAI21X1_1202 ( .A(_5302__bF_buf2), .B(_6250__bF_buf6), .C(_6264_), .Y(_1318_) );
NAND3X1 NAND3X1_1080 ( .A(datapath_1_RegisterFile_regfile_mem_28__14_), .B(_5265__bF_buf59), .C(_6250__bF_buf7), .Y(_6265_) );
OAI21X1 OAI21X1_1203 ( .A(_5304__bF_buf4), .B(_6250__bF_buf7), .C(_6265_), .Y(_1838_) );
NAND3X1 NAND3X1_1081 ( .A(datapath_1_RegisterFile_regfile_mem_28__15_), .B(_5265__bF_buf69), .C(_6250__bF_buf4), .Y(_6266_) );
OAI21X1 OAI21X1_1204 ( .A(_5306__bF_buf0), .B(_6250__bF_buf4), .C(_6266_), .Y(_1319_) );
NAND3X1 NAND3X1_1082 ( .A(datapath_1_RegisterFile_regfile_mem_28__16_), .B(_5265__bF_buf40), .C(_6250__bF_buf1), .Y(_6267_) );
OAI21X1 OAI21X1_1205 ( .A(_5308__bF_buf4), .B(_6250__bF_buf1), .C(_6267_), .Y(_1320_) );
NAND3X1 NAND3X1_1083 ( .A(datapath_1_RegisterFile_regfile_mem_28__17_), .B(_5265__bF_buf90), .C(_6250__bF_buf2), .Y(_6268_) );
OAI21X1 OAI21X1_1206 ( .A(_5310__bF_buf2), .B(_6250__bF_buf2), .C(_6268_), .Y(_1321_) );
NAND3X1 NAND3X1_1084 ( .A(datapath_1_RegisterFile_regfile_mem_28__18_), .B(_5265__bF_buf59), .C(_6250__bF_buf7), .Y(_6269_) );
OAI21X1 OAI21X1_1207 ( .A(_5312__bF_buf3), .B(_6250__bF_buf7), .C(_6269_), .Y(_1322_) );
NAND3X1 NAND3X1_1085 ( .A(datapath_1_RegisterFile_regfile_mem_28__19_), .B(_5265__bF_buf20), .C(_6250__bF_buf1), .Y(_6270_) );
OAI21X1 OAI21X1_1208 ( .A(_5314__bF_buf2), .B(_6250__bF_buf1), .C(_6270_), .Y(_1323_) );
NAND3X1 NAND3X1_1086 ( .A(datapath_1_RegisterFile_regfile_mem_28__20_), .B(_5265__bF_buf9), .C(_6250__bF_buf5), .Y(_6271_) );
OAI21X1 OAI21X1_1209 ( .A(_5316__bF_buf0), .B(_6250__bF_buf5), .C(_6271_), .Y(_1325_) );
NAND3X1 NAND3X1_1087 ( .A(datapath_1_RegisterFile_regfile_mem_28__21_), .B(_5265__bF_buf61), .C(_6250__bF_buf3), .Y(_6272_) );
OAI21X1 OAI21X1_1210 ( .A(_5318__bF_buf3), .B(_6250__bF_buf3), .C(_6272_), .Y(_1326_) );
NAND3X1 NAND3X1_1088 ( .A(datapath_1_RegisterFile_regfile_mem_28__22_), .B(_5265__bF_buf33), .C(_6250__bF_buf6), .Y(_6273_) );
OAI21X1 OAI21X1_1211 ( .A(_5320__bF_buf3), .B(_6250__bF_buf6), .C(_6273_), .Y(_1327_) );
NAND3X1 NAND3X1_1089 ( .A(datapath_1_RegisterFile_regfile_mem_28__23_), .B(_5265__bF_buf95), .C(_6250__bF_buf0), .Y(_6274_) );
OAI21X1 OAI21X1_1212 ( .A(_5322__bF_buf4), .B(_6250__bF_buf0), .C(_6274_), .Y(_1328_) );
NAND3X1 NAND3X1_1090 ( .A(datapath_1_RegisterFile_regfile_mem_28__24_), .B(_5265__bF_buf88), .C(_6250__bF_buf4), .Y(_6275_) );
OAI21X1 OAI21X1_1213 ( .A(_5324__bF_buf4), .B(_6250__bF_buf4), .C(_6275_), .Y(_1839_) );
NAND3X1 NAND3X1_1091 ( .A(datapath_1_RegisterFile_regfile_mem_28__25_), .B(_5265__bF_buf80), .C(_6250__bF_buf0), .Y(_6276_) );
OAI21X1 OAI21X1_1214 ( .A(_5326__bF_buf3), .B(_6250__bF_buf0), .C(_6276_), .Y(_1329_) );
NAND3X1 NAND3X1_1092 ( .A(datapath_1_RegisterFile_regfile_mem_28__26_), .B(_5265__bF_buf90), .C(_6250__bF_buf6), .Y(_6277_) );
OAI21X1 OAI21X1_1215 ( .A(_5328__bF_buf0), .B(_6250__bF_buf6), .C(_6277_), .Y(_1330_) );
NAND3X1 NAND3X1_1093 ( .A(datapath_1_RegisterFile_regfile_mem_28__27_), .B(_5265__bF_buf73), .C(_6250__bF_buf7), .Y(_6278_) );
OAI21X1 OAI21X1_1216 ( .A(_5330__bF_buf0), .B(_6250__bF_buf7), .C(_6278_), .Y(_1840_) );
NAND3X1 NAND3X1_1094 ( .A(datapath_1_RegisterFile_regfile_mem_28__28_), .B(_5265__bF_buf69), .C(_6250__bF_buf4), .Y(_6279_) );
OAI21X1 OAI21X1_1217 ( .A(_5332__bF_buf3), .B(_6250__bF_buf4), .C(_6279_), .Y(_1841_) );
NAND3X1 NAND3X1_1095 ( .A(datapath_1_RegisterFile_regfile_mem_28__29_), .B(_5265__bF_buf40), .C(_6250__bF_buf1), .Y(_6280_) );
OAI21X1 OAI21X1_1218 ( .A(_5334__bF_buf0), .B(_6250__bF_buf1), .C(_6280_), .Y(_1842_) );
NAND3X1 NAND3X1_1096 ( .A(datapath_1_RegisterFile_regfile_mem_28__30_), .B(_5265__bF_buf8), .C(_6250__bF_buf3), .Y(_6281_) );
OAI21X1 OAI21X1_1219 ( .A(_5336__bF_buf1), .B(_6250__bF_buf3), .C(_6281_), .Y(_1843_) );
NAND3X1 NAND3X1_1097 ( .A(datapath_1_RegisterFile_regfile_mem_28__31_), .B(_5265__bF_buf59), .C(_6250__bF_buf7), .Y(_6282_) );
OAI21X1 OAI21X1_1220 ( .A(_5338__bF_buf1), .B(_6250__bF_buf7), .C(_6282_), .Y(_1844_) );
NAND2X1 NAND2X1_390 ( .A(_6249_), .B(_5341_), .Y(_6283_) );
NAND3X1 NAND3X1_1098 ( .A(datapath_1_RegisterFile_regfile_mem_29__0_), .B(_5265__bF_buf90), .C(_6283__bF_buf7), .Y(_6284_) );
OAI21X1 OAI21X1_1221 ( .A(_5276__bF_buf3), .B(_6283__bF_buf7), .C(_6284_), .Y(_1338_) );
NAND3X1 NAND3X1_1099 ( .A(datapath_1_RegisterFile_regfile_mem_29__1_), .B(_5265__bF_buf19), .C(_6283__bF_buf3), .Y(_6285_) );
OAI21X1 OAI21X1_1222 ( .A(_5278__bF_buf4), .B(_6283__bF_buf3), .C(_6285_), .Y(_1348_) );
NAND3X1 NAND3X1_1100 ( .A(datapath_1_RegisterFile_regfile_mem_29__2_), .B(_5265__bF_buf19), .C(_6283__bF_buf6), .Y(_6286_) );
OAI21X1 OAI21X1_1223 ( .A(_5280__bF_buf0), .B(_6283__bF_buf6), .C(_6286_), .Y(_1358_) );
NAND3X1 NAND3X1_1101 ( .A(datapath_1_RegisterFile_regfile_mem_29__3_), .B(_5265__bF_buf3), .C(_6283__bF_buf6), .Y(_6287_) );
OAI21X1 OAI21X1_1224 ( .A(_5282__bF_buf2), .B(_6283__bF_buf6), .C(_6287_), .Y(_1361_) );
NAND3X1 NAND3X1_1102 ( .A(datapath_1_RegisterFile_regfile_mem_29__4_), .B(_5265__bF_buf46), .C(_6283__bF_buf0), .Y(_6288_) );
OAI21X1 OAI21X1_1225 ( .A(_5284__bF_buf3), .B(_6283__bF_buf0), .C(_6288_), .Y(_1362_) );
NAND3X1 NAND3X1_1103 ( .A(datapath_1_RegisterFile_regfile_mem_29__5_), .B(_5265__bF_buf58), .C(_6283__bF_buf5), .Y(_6289_) );
OAI21X1 OAI21X1_1226 ( .A(_5286__bF_buf3), .B(_6283__bF_buf5), .C(_6289_), .Y(_1363_) );
NAND3X1 NAND3X1_1104 ( .A(datapath_1_RegisterFile_regfile_mem_29__6_), .B(_5265__bF_buf61), .C(_6283__bF_buf0), .Y(_6290_) );
OAI21X1 OAI21X1_1227 ( .A(_5288__bF_buf0), .B(_6283__bF_buf0), .C(_6290_), .Y(_1364_) );
NAND3X1 NAND3X1_1105 ( .A(datapath_1_RegisterFile_regfile_mem_29__7_), .B(_5265__bF_buf36), .C(_6283__bF_buf1), .Y(_6291_) );
OAI21X1 OAI21X1_1228 ( .A(_5290__bF_buf3), .B(_6283__bF_buf1), .C(_6291_), .Y(_1365_) );
NAND3X1 NAND3X1_1106 ( .A(datapath_1_RegisterFile_regfile_mem_29__8_), .B(_5265__bF_buf46), .C(_6283__bF_buf0), .Y(_6292_) );
OAI21X1 OAI21X1_1229 ( .A(_5292__bF_buf2), .B(_6283__bF_buf0), .C(_6292_), .Y(_1366_) );
NAND3X1 NAND3X1_1107 ( .A(datapath_1_RegisterFile_regfile_mem_29__9_), .B(_5265__bF_buf12), .C(_6283__bF_buf7), .Y(_6293_) );
OAI21X1 OAI21X1_1230 ( .A(_5294__bF_buf0), .B(_6283__bF_buf7), .C(_6293_), .Y(_1845_) );
NAND3X1 NAND3X1_1108 ( .A(datapath_1_RegisterFile_regfile_mem_29__10_), .B(_5265__bF_buf12), .C(_6283__bF_buf7), .Y(_6294_) );
OAI21X1 OAI21X1_1231 ( .A(_5296__bF_buf3), .B(_6283__bF_buf7), .C(_6294_), .Y(_1339_) );
NAND3X1 NAND3X1_1109 ( .A(datapath_1_RegisterFile_regfile_mem_29__11_), .B(_5265__bF_buf36), .C(_6283__bF_buf1), .Y(_6295_) );
OAI21X1 OAI21X1_1232 ( .A(_5298__bF_buf4), .B(_6283__bF_buf1), .C(_6295_), .Y(_1340_) );
NAND3X1 NAND3X1_1110 ( .A(datapath_1_RegisterFile_regfile_mem_29__12_), .B(_5265__bF_buf63), .C(_6283__bF_buf6), .Y(_6296_) );
OAI21X1 OAI21X1_1233 ( .A(_5300__bF_buf4), .B(_6283__bF_buf6), .C(_6296_), .Y(_1341_) );
NAND3X1 NAND3X1_1111 ( .A(datapath_1_RegisterFile_regfile_mem_29__13_), .B(_5265__bF_buf33), .C(_6283__bF_buf5), .Y(_6297_) );
OAI21X1 OAI21X1_1234 ( .A(_5302__bF_buf2), .B(_6283__bF_buf5), .C(_6297_), .Y(_1342_) );
NAND3X1 NAND3X1_1112 ( .A(datapath_1_RegisterFile_regfile_mem_29__14_), .B(_5265__bF_buf22), .C(_6283__bF_buf4), .Y(_6298_) );
OAI21X1 OAI21X1_1235 ( .A(_5304__bF_buf3), .B(_6283__bF_buf4), .C(_6298_), .Y(_1343_) );
NAND3X1 NAND3X1_1113 ( .A(datapath_1_RegisterFile_regfile_mem_29__15_), .B(_5265__bF_buf20), .C(_6283__bF_buf6), .Y(_6299_) );
OAI21X1 OAI21X1_1236 ( .A(_5306__bF_buf4), .B(_6283__bF_buf6), .C(_6299_), .Y(_1344_) );
NAND3X1 NAND3X1_1114 ( .A(datapath_1_RegisterFile_regfile_mem_29__16_), .B(_5265__bF_buf41), .C(_6283__bF_buf2), .Y(_6300_) );
OAI21X1 OAI21X1_1237 ( .A(_5308__bF_buf4), .B(_6283__bF_buf2), .C(_6300_), .Y(_1345_) );
NAND3X1 NAND3X1_1115 ( .A(datapath_1_RegisterFile_regfile_mem_29__17_), .B(_5265__bF_buf28), .C(_6283__bF_buf7), .Y(_6301_) );
OAI21X1 OAI21X1_1238 ( .A(_5310__bF_buf2), .B(_6283__bF_buf7), .C(_6301_), .Y(_1346_) );
NAND3X1 NAND3X1_1116 ( .A(datapath_1_RegisterFile_regfile_mem_29__18_), .B(_5265__bF_buf58), .C(_6283__bF_buf5), .Y(_6302_) );
OAI21X1 OAI21X1_1239 ( .A(_5312__bF_buf4), .B(_6283__bF_buf5), .C(_6302_), .Y(_1347_) );
NAND3X1 NAND3X1_1117 ( .A(datapath_1_RegisterFile_regfile_mem_29__19_), .B(_5265__bF_buf19), .C(_6283__bF_buf3), .Y(_6303_) );
OAI21X1 OAI21X1_1240 ( .A(_5314__bF_buf0), .B(_6283__bF_buf3), .C(_6303_), .Y(_1846_) );
NAND3X1 NAND3X1_1118 ( .A(datapath_1_RegisterFile_regfile_mem_29__20_), .B(_5265__bF_buf30), .C(_6283__bF_buf1), .Y(_6304_) );
OAI21X1 OAI21X1_1241 ( .A(_5316__bF_buf1), .B(_6283__bF_buf1), .C(_6304_), .Y(_1349_) );
NAND3X1 NAND3X1_1119 ( .A(datapath_1_RegisterFile_regfile_mem_29__21_), .B(_5265__bF_buf4), .C(_6283__bF_buf3), .Y(_6305_) );
OAI21X1 OAI21X1_1242 ( .A(_5318__bF_buf2), .B(_6283__bF_buf3), .C(_6305_), .Y(_1350_) );
NAND3X1 NAND3X1_1120 ( .A(datapath_1_RegisterFile_regfile_mem_29__22_), .B(_5265__bF_buf33), .C(_6283__bF_buf5), .Y(_6306_) );
OAI21X1 OAI21X1_1243 ( .A(_5320__bF_buf3), .B(_6283__bF_buf5), .C(_6306_), .Y(_1351_) );
NAND3X1 NAND3X1_1121 ( .A(datapath_1_RegisterFile_regfile_mem_29__23_), .B(_5265__bF_buf4), .C(_6283__bF_buf3), .Y(_6307_) );
OAI21X1 OAI21X1_1244 ( .A(_5322__bF_buf0), .B(_6283__bF_buf3), .C(_6307_), .Y(_1352_) );
NAND3X1 NAND3X1_1122 ( .A(datapath_1_RegisterFile_regfile_mem_29__24_), .B(_5265__bF_buf40), .C(_6283__bF_buf2), .Y(_6308_) );
OAI21X1 OAI21X1_1245 ( .A(_5324__bF_buf1), .B(_6283__bF_buf2), .C(_6308_), .Y(_1353_) );
NAND3X1 NAND3X1_1123 ( .A(datapath_1_RegisterFile_regfile_mem_29__25_), .B(_5265__bF_buf80), .C(_6283__bF_buf2), .Y(_6309_) );
OAI21X1 OAI21X1_1246 ( .A(_5326__bF_buf3), .B(_6283__bF_buf2), .C(_6309_), .Y(_1354_) );
NAND3X1 NAND3X1_1124 ( .A(datapath_1_RegisterFile_regfile_mem_29__26_), .B(_5265__bF_buf31), .C(_6283__bF_buf4), .Y(_6310_) );
OAI21X1 OAI21X1_1247 ( .A(_5328__bF_buf0), .B(_6283__bF_buf4), .C(_6310_), .Y(_1355_) );
NAND3X1 NAND3X1_1125 ( .A(datapath_1_RegisterFile_regfile_mem_29__27_), .B(_5265__bF_buf22), .C(_6283__bF_buf4), .Y(_6311_) );
OAI21X1 OAI21X1_1248 ( .A(_5330__bF_buf0), .B(_6283__bF_buf4), .C(_6311_), .Y(_1356_) );
NAND3X1 NAND3X1_1126 ( .A(datapath_1_RegisterFile_regfile_mem_29__28_), .B(_5265__bF_buf69), .C(_6283__bF_buf1), .Y(_6312_) );
OAI21X1 OAI21X1_1249 ( .A(_5332__bF_buf3), .B(_6283__bF_buf1), .C(_6312_), .Y(_1357_) );
NAND3X1 NAND3X1_1127 ( .A(datapath_1_RegisterFile_regfile_mem_29__29_), .B(_5265__bF_buf41), .C(_6283__bF_buf2), .Y(_6313_) );
OAI21X1 OAI21X1_1250 ( .A(_5334__bF_buf0), .B(_6283__bF_buf2), .C(_6313_), .Y(_1847_) );
NAND3X1 NAND3X1_1128 ( .A(datapath_1_RegisterFile_regfile_mem_29__30_), .B(_5265__bF_buf61), .C(_6283__bF_buf0), .Y(_6314_) );
OAI21X1 OAI21X1_1251 ( .A(_5336__bF_buf0), .B(_6283__bF_buf0), .C(_6314_), .Y(_1359_) );
NAND3X1 NAND3X1_1129 ( .A(datapath_1_RegisterFile_regfile_mem_29__31_), .B(_5265__bF_buf31), .C(_6283__bF_buf4), .Y(_6315_) );
OAI21X1 OAI21X1_1252 ( .A(_5338__bF_buf4), .B(_6283__bF_buf4), .C(_6315_), .Y(_1360_) );
NAND2X1 NAND2X1_391 ( .A(_6249_), .B(_5376_), .Y(_6316_) );
NAND3X1 NAND3X1_1130 ( .A(datapath_1_RegisterFile_regfile_mem_30__0_), .B(_5265__bF_buf75), .C(_6316__bF_buf7), .Y(_6317_) );
OAI21X1 OAI21X1_1253 ( .A(_5276__bF_buf1), .B(_6316__bF_buf7), .C(_6317_), .Y(_1848_) );
NAND3X1 NAND3X1_1131 ( .A(datapath_1_RegisterFile_regfile_mem_30__1_), .B(_5265__bF_buf16), .C(_6316__bF_buf0), .Y(_6318_) );
OAI21X1 OAI21X1_1254 ( .A(_5278__bF_buf1), .B(_6316__bF_buf0), .C(_6318_), .Y(_1849_) );
NAND3X1 NAND3X1_1132 ( .A(datapath_1_RegisterFile_regfile_mem_30__2_), .B(_5265__bF_buf19), .C(_6316__bF_buf5), .Y(_6319_) );
OAI21X1 OAI21X1_1255 ( .A(_5280__bF_buf4), .B(_6316__bF_buf5), .C(_6319_), .Y(_1850_) );
NAND3X1 NAND3X1_1133 ( .A(datapath_1_RegisterFile_regfile_mem_30__3_), .B(_5265__bF_buf14), .C(_6316__bF_buf5), .Y(_6320_) );
OAI21X1 OAI21X1_1256 ( .A(_5282__bF_buf1), .B(_6316__bF_buf5), .C(_6320_), .Y(_1851_) );
NAND3X1 NAND3X1_1134 ( .A(datapath_1_RegisterFile_regfile_mem_30__4_), .B(_5265__bF_buf61), .C(_6316__bF_buf1), .Y(_6321_) );
OAI21X1 OAI21X1_1257 ( .A(_5284__bF_buf2), .B(_6316__bF_buf1), .C(_6321_), .Y(_1852_) );
NAND3X1 NAND3X1_1135 ( .A(datapath_1_RegisterFile_regfile_mem_30__5_), .B(_5265__bF_buf58), .C(_6316__bF_buf3), .Y(_6322_) );
OAI21X1 OAI21X1_1258 ( .A(_5286__bF_buf4), .B(_6316__bF_buf3), .C(_6322_), .Y(_1853_) );
NAND3X1 NAND3X1_1136 ( .A(datapath_1_RegisterFile_regfile_mem_30__6_), .B(_5265__bF_buf55), .C(_6316__bF_buf6), .Y(_6323_) );
OAI21X1 OAI21X1_1259 ( .A(_5288__bF_buf4), .B(_6316__bF_buf6), .C(_6323_), .Y(_1854_) );
NAND3X1 NAND3X1_1137 ( .A(datapath_1_RegisterFile_regfile_mem_30__7_), .B(_5265__bF_buf3), .C(_6316__bF_buf4), .Y(_6324_) );
OAI21X1 OAI21X1_1260 ( .A(_5290__bF_buf3), .B(_6316__bF_buf4), .C(_6324_), .Y(_1416_) );
NAND3X1 NAND3X1_1138 ( .A(datapath_1_RegisterFile_regfile_mem_30__8_), .B(_5265__bF_buf46), .C(_6316__bF_buf1), .Y(_6325_) );
OAI21X1 OAI21X1_1261 ( .A(_5292__bF_buf4), .B(_6316__bF_buf1), .C(_6325_), .Y(_1417_) );
NAND3X1 NAND3X1_1139 ( .A(datapath_1_RegisterFile_regfile_mem_30__9_), .B(_5265__bF_buf90), .C(_6316__bF_buf7), .Y(_6326_) );
OAI21X1 OAI21X1_1262 ( .A(_5294__bF_buf0), .B(_6316__bF_buf7), .C(_6326_), .Y(_1418_) );
NAND3X1 NAND3X1_1140 ( .A(datapath_1_RegisterFile_regfile_mem_30__10_), .B(_5265__bF_buf31), .C(_6316__bF_buf3), .Y(_6327_) );
OAI21X1 OAI21X1_1263 ( .A(_5296__bF_buf1), .B(_6316__bF_buf3), .C(_6327_), .Y(_1396_) );
NAND3X1 NAND3X1_1141 ( .A(datapath_1_RegisterFile_regfile_mem_30__11_), .B(_5265__bF_buf36), .C(_6316__bF_buf4), .Y(_6328_) );
OAI21X1 OAI21X1_1264 ( .A(_5298__bF_buf0), .B(_6316__bF_buf4), .C(_6328_), .Y(_1397_) );
NAND3X1 NAND3X1_1142 ( .A(datapath_1_RegisterFile_regfile_mem_30__12_), .B(_5265__bF_buf55), .C(_6316__bF_buf6), .Y(_6329_) );
OAI21X1 OAI21X1_1265 ( .A(_5300__bF_buf4), .B(_6316__bF_buf6), .C(_6329_), .Y(_1398_) );
NAND3X1 NAND3X1_1143 ( .A(datapath_1_RegisterFile_regfile_mem_30__13_), .B(_5265__bF_buf1), .C(_6316__bF_buf3), .Y(_6330_) );
OAI21X1 OAI21X1_1266 ( .A(_5302__bF_buf3), .B(_6316__bF_buf3), .C(_6330_), .Y(_1399_) );
NAND3X1 NAND3X1_1144 ( .A(datapath_1_RegisterFile_regfile_mem_30__14_), .B(_5265__bF_buf22), .C(_6316__bF_buf2), .Y(_6331_) );
OAI21X1 OAI21X1_1267 ( .A(_5304__bF_buf3), .B(_6316__bF_buf2), .C(_6331_), .Y(_1855_) );
NAND3X1 NAND3X1_1145 ( .A(datapath_1_RegisterFile_regfile_mem_30__15_), .B(_5265__bF_buf16), .C(_6316__bF_buf0), .Y(_6332_) );
OAI21X1 OAI21X1_1268 ( .A(_5306__bF_buf2), .B(_6316__bF_buf0), .C(_6332_), .Y(_1400_) );
NAND3X1 NAND3X1_1146 ( .A(datapath_1_RegisterFile_regfile_mem_30__16_), .B(_5265__bF_buf24), .C(_6316__bF_buf0), .Y(_6333_) );
OAI21X1 OAI21X1_1269 ( .A(_5308__bF_buf1), .B(_6316__bF_buf0), .C(_6333_), .Y(_1401_) );
NAND3X1 NAND3X1_1147 ( .A(datapath_1_RegisterFile_regfile_mem_30__17_), .B(_5265__bF_buf61), .C(_6316__bF_buf7), .Y(_6334_) );
OAI21X1 OAI21X1_1270 ( .A(_5310__bF_buf3), .B(_6316__bF_buf7), .C(_6334_), .Y(_1402_) );
NAND3X1 NAND3X1_1148 ( .A(datapath_1_RegisterFile_regfile_mem_30__18_), .B(_5265__bF_buf73), .C(_6316__bF_buf2), .Y(_6335_) );
OAI21X1 OAI21X1_1271 ( .A(_5312__bF_buf3), .B(_6316__bF_buf2), .C(_6335_), .Y(_1403_) );
NAND3X1 NAND3X1_1149 ( .A(datapath_1_RegisterFile_regfile_mem_30__19_), .B(_5265__bF_buf55), .C(_6316__bF_buf6), .Y(_6336_) );
OAI21X1 OAI21X1_1272 ( .A(_5314__bF_buf0), .B(_6316__bF_buf6), .C(_6336_), .Y(_1404_) );
NAND3X1 NAND3X1_1150 ( .A(datapath_1_RegisterFile_regfile_mem_30__20_), .B(_5265__bF_buf36), .C(_6316__bF_buf4), .Y(_6337_) );
OAI21X1 OAI21X1_1273 ( .A(_5316__bF_buf0), .B(_6316__bF_buf4), .C(_6337_), .Y(_1405_) );
NAND3X1 NAND3X1_1151 ( .A(datapath_1_RegisterFile_regfile_mem_30__21_), .B(_5265__bF_buf75), .C(_6316__bF_buf7), .Y(_6338_) );
OAI21X1 OAI21X1_1274 ( .A(_5318__bF_buf3), .B(_6316__bF_buf7), .C(_6338_), .Y(_1406_) );
NAND3X1 NAND3X1_1152 ( .A(datapath_1_RegisterFile_regfile_mem_30__22_), .B(_5265__bF_buf1), .C(_6316__bF_buf3), .Y(_6339_) );
OAI21X1 OAI21X1_1275 ( .A(_5320__bF_buf0), .B(_6316__bF_buf3), .C(_6339_), .Y(_1407_) );
NAND3X1 NAND3X1_1153 ( .A(datapath_1_RegisterFile_regfile_mem_30__23_), .B(_5265__bF_buf55), .C(_6316__bF_buf6), .Y(_6340_) );
OAI21X1 OAI21X1_1276 ( .A(_5322__bF_buf0), .B(_6316__bF_buf6), .C(_6340_), .Y(_1408_) );
NAND3X1 NAND3X1_1154 ( .A(datapath_1_RegisterFile_regfile_mem_30__24_), .B(_5265__bF_buf40), .C(_6316__bF_buf5), .Y(_6341_) );
OAI21X1 OAI21X1_1277 ( .A(_5324__bF_buf1), .B(_6316__bF_buf5), .C(_6341_), .Y(_1856_) );
NAND3X1 NAND3X1_1155 ( .A(datapath_1_RegisterFile_regfile_mem_30__25_), .B(_5265__bF_buf67), .C(_6316__bF_buf0), .Y(_6342_) );
OAI21X1 OAI21X1_1278 ( .A(_5326__bF_buf4), .B(_6316__bF_buf0), .C(_6342_), .Y(_1409_) );
NAND3X1 NAND3X1_1156 ( .A(datapath_1_RegisterFile_regfile_mem_30__26_), .B(_5265__bF_buf82), .C(_6316__bF_buf1), .Y(_6343_) );
OAI21X1 OAI21X1_1279 ( .A(_5328__bF_buf4), .B(_6316__bF_buf1), .C(_6343_), .Y(_1410_) );
NAND3X1 NAND3X1_1157 ( .A(datapath_1_RegisterFile_regfile_mem_30__27_), .B(_5265__bF_buf73), .C(_6316__bF_buf2), .Y(_6344_) );
OAI21X1 OAI21X1_1280 ( .A(_5330__bF_buf0), .B(_6316__bF_buf2), .C(_6344_), .Y(_1411_) );
NAND3X1 NAND3X1_1158 ( .A(datapath_1_RegisterFile_regfile_mem_30__28_), .B(_5265__bF_buf14), .C(_6316__bF_buf4), .Y(_6345_) );
OAI21X1 OAI21X1_1281 ( .A(_5332__bF_buf3), .B(_6316__bF_buf4), .C(_6345_), .Y(_1412_) );
NAND3X1 NAND3X1_1159 ( .A(datapath_1_RegisterFile_regfile_mem_30__29_), .B(_5265__bF_buf80), .C(_6316__bF_buf5), .Y(_6346_) );
OAI21X1 OAI21X1_1282 ( .A(_5334__bF_buf0), .B(_6316__bF_buf5), .C(_6346_), .Y(_1413_) );
NAND3X1 NAND3X1_1160 ( .A(datapath_1_RegisterFile_regfile_mem_30__30_), .B(_5265__bF_buf82), .C(_6316__bF_buf1), .Y(_6347_) );
OAI21X1 OAI21X1_1283 ( .A(_5336__bF_buf1), .B(_6316__bF_buf1), .C(_6347_), .Y(_1414_) );
NAND3X1 NAND3X1_1161 ( .A(datapath_1_RegisterFile_regfile_mem_30__31_), .B(_5265__bF_buf59), .C(_6316__bF_buf2), .Y(_6348_) );
OAI21X1 OAI21X1_1284 ( .A(_5338__bF_buf4), .B(_6316__bF_buf2), .C(_6348_), .Y(_1415_) );
OR2X2 OR2X2_2 ( .A(rst_bF_buf2), .B(RegWrite), .Y(_6349_) );
NAND3X1 NAND3X1_1162 ( .A(_5410_), .B(_6349_), .C(_6249_), .Y(_6350_) );
NAND2X1 NAND2X1_392 ( .A(datapath_1_RegisterFile_regfile_mem_31__0_), .B(_6350__bF_buf1), .Y(_6351_) );
OAI21X1 OAI21X1_1285 ( .A(_5276__bF_buf1), .B(_6350__bF_buf1), .C(_6351_), .Y(_1419_) );
NAND2X1 NAND2X1_393 ( .A(datapath_1_RegisterFile_regfile_mem_31__1_), .B(_6350__bF_buf4), .Y(_6352_) );
OAI21X1 OAI21X1_1286 ( .A(_5278__bF_buf4), .B(_6350__bF_buf4), .C(_6352_), .Y(_1857_) );
NAND2X1 NAND2X1_394 ( .A(datapath_1_RegisterFile_regfile_mem_31__2_), .B(_6350__bF_buf4), .Y(_6353_) );
OAI21X1 OAI21X1_1287 ( .A(_5280__bF_buf0), .B(_6350__bF_buf4), .C(_6353_), .Y(_1438_) );
NAND2X1 NAND2X1_395 ( .A(datapath_1_RegisterFile_regfile_mem_31__3_), .B(_6350__bF_buf5), .Y(_6354_) );
OAI21X1 OAI21X1_1288 ( .A(_5282__bF_buf2), .B(_6350__bF_buf5), .C(_6354_), .Y(_1440_) );
NAND2X1 NAND2X1_396 ( .A(datapath_1_RegisterFile_regfile_mem_31__4_), .B(_6350__bF_buf7), .Y(_6355_) );
OAI21X1 OAI21X1_1289 ( .A(_5284__bF_buf3), .B(_6350__bF_buf7), .C(_6355_), .Y(_1441_) );
NAND2X1 NAND2X1_397 ( .A(datapath_1_RegisterFile_regfile_mem_31__5_), .B(_6350__bF_buf6), .Y(_6356_) );
OAI21X1 OAI21X1_1290 ( .A(_5286__bF_buf4), .B(_6350__bF_buf6), .C(_6356_), .Y(_1442_) );
NAND2X1 NAND2X1_398 ( .A(datapath_1_RegisterFile_regfile_mem_31__6_), .B(_6350__bF_buf1), .Y(_6357_) );
OAI21X1 OAI21X1_1291 ( .A(_5288__bF_buf4), .B(_6350__bF_buf1), .C(_6357_), .Y(_1443_) );
NAND2X1 NAND2X1_399 ( .A(datapath_1_RegisterFile_regfile_mem_31__7_), .B(_6350__bF_buf5), .Y(_6358_) );
OAI21X1 OAI21X1_1292 ( .A(_5290__bF_buf3), .B(_6350__bF_buf5), .C(_6358_), .Y(_1444_) );
NAND2X1 NAND2X1_400 ( .A(datapath_1_RegisterFile_regfile_mem_31__8_), .B(_6350__bF_buf1), .Y(_6359_) );
OAI21X1 OAI21X1_1293 ( .A(_5292__bF_buf4), .B(_6350__bF_buf1), .C(_6359_), .Y(_1445_) );
NAND2X1 NAND2X1_401 ( .A(datapath_1_RegisterFile_regfile_mem_31__9_), .B(_6350__bF_buf6), .Y(_6360_) );
OAI21X1 OAI21X1_1294 ( .A(_5294__bF_buf0), .B(_6350__bF_buf6), .C(_6360_), .Y(_1446_) );
NAND2X1 NAND2X1_402 ( .A(datapath_1_RegisterFile_regfile_mem_31__10_), .B(_6350__bF_buf6), .Y(_6361_) );
OAI21X1 OAI21X1_1295 ( .A(_5296__bF_buf1), .B(_6350__bF_buf6), .C(_6361_), .Y(_1420_) );
NAND2X1 NAND2X1_403 ( .A(datapath_1_RegisterFile_regfile_mem_31__11_), .B(_6350__bF_buf5), .Y(_6362_) );
OAI21X1 OAI21X1_1296 ( .A(_5298__bF_buf0), .B(_6350__bF_buf5), .C(_6362_), .Y(_1858_) );
NAND2X1 NAND2X1_404 ( .A(datapath_1_RegisterFile_regfile_mem_31__12_), .B(_6350__bF_buf4), .Y(_6363_) );
OAI21X1 OAI21X1_1297 ( .A(_5300__bF_buf4), .B(_6350__bF_buf4), .C(_6363_), .Y(_1421_) );
NAND2X1 NAND2X1_405 ( .A(datapath_1_RegisterFile_regfile_mem_31__13_), .B(_6350__bF_buf2), .Y(_6364_) );
OAI21X1 OAI21X1_1298 ( .A(_5302__bF_buf3), .B(_6350__bF_buf2), .C(_6364_), .Y(_1422_) );
NAND2X1 NAND2X1_406 ( .A(datapath_1_RegisterFile_regfile_mem_31__14_), .B(_6350__bF_buf3), .Y(_6365_) );
OAI21X1 OAI21X1_1299 ( .A(_5304__bF_buf3), .B(_6350__bF_buf3), .C(_6365_), .Y(_1423_) );
NAND2X1 NAND2X1_407 ( .A(datapath_1_RegisterFile_regfile_mem_31__15_), .B(_6350__bF_buf0), .Y(_6366_) );
OAI21X1 OAI21X1_1300 ( .A(_5306__bF_buf2), .B(_6350__bF_buf0), .C(_6366_), .Y(_1424_) );
NAND2X1 NAND2X1_408 ( .A(datapath_1_RegisterFile_regfile_mem_31__16_), .B(_6350__bF_buf0), .Y(_6367_) );
OAI21X1 OAI21X1_1301 ( .A(_5308__bF_buf4), .B(_6350__bF_buf0), .C(_6367_), .Y(_1425_) );
NAND2X1 NAND2X1_409 ( .A(datapath_1_RegisterFile_regfile_mem_31__17_), .B(_6350__bF_buf6), .Y(_6368_) );
OAI21X1 OAI21X1_1302 ( .A(_5310__bF_buf3), .B(_6350__bF_buf6), .C(_6368_), .Y(_1426_) );
NAND2X1 NAND2X1_410 ( .A(datapath_1_RegisterFile_regfile_mem_31__18_), .B(_6350__bF_buf3), .Y(_6369_) );
OAI21X1 OAI21X1_1303 ( .A(_5312__bF_buf3), .B(_6350__bF_buf3), .C(_6369_), .Y(_1427_) );
NAND2X1 NAND2X1_411 ( .A(datapath_1_RegisterFile_regfile_mem_31__19_), .B(_6350__bF_buf4), .Y(_6370_) );
OAI21X1 OAI21X1_1304 ( .A(_5314__bF_buf0), .B(_6350__bF_buf4), .C(_6370_), .Y(_1428_) );
NAND2X1 NAND2X1_412 ( .A(datapath_1_RegisterFile_regfile_mem_31__20_), .B(_6350__bF_buf5), .Y(_6371_) );
OAI21X1 OAI21X1_1305 ( .A(_5316__bF_buf0), .B(_6350__bF_buf5), .C(_6371_), .Y(_1429_) );
NAND2X1 NAND2X1_413 ( .A(datapath_1_RegisterFile_regfile_mem_31__21_), .B(_6350__bF_buf1), .Y(_6372_) );
OAI21X1 OAI21X1_1306 ( .A(_5318__bF_buf3), .B(_6350__bF_buf1), .C(_6372_), .Y(_1859_) );
NAND2X1 NAND2X1_414 ( .A(datapath_1_RegisterFile_regfile_mem_31__22_), .B(_6350__bF_buf2), .Y(_6373_) );
OAI21X1 OAI21X1_1307 ( .A(_5320__bF_buf1), .B(_6350__bF_buf2), .C(_6373_), .Y(_1430_) );
NAND2X1 NAND2X1_415 ( .A(datapath_1_RegisterFile_regfile_mem_31__23_), .B(_6350__bF_buf7), .Y(_6374_) );
OAI21X1 OAI21X1_1308 ( .A(_5322__bF_buf4), .B(_6350__bF_buf7), .C(_6374_), .Y(_1431_) );
NAND2X1 NAND2X1_416 ( .A(datapath_1_RegisterFile_regfile_mem_31__24_), .B(_6350__bF_buf0), .Y(_6375_) );
OAI21X1 OAI21X1_1309 ( .A(_5324__bF_buf4), .B(_6350__bF_buf0), .C(_6375_), .Y(_1432_) );
NAND2X1 NAND2X1_417 ( .A(datapath_1_RegisterFile_regfile_mem_31__25_), .B(_6350__bF_buf7), .Y(_6376_) );
OAI21X1 OAI21X1_1310 ( .A(_5326__bF_buf3), .B(_6350__bF_buf7), .C(_6376_), .Y(_1433_) );
NAND2X1 NAND2X1_418 ( .A(datapath_1_RegisterFile_regfile_mem_31__26_), .B(_6350__bF_buf2), .Y(_6377_) );
OAI21X1 OAI21X1_1311 ( .A(_5328__bF_buf4), .B(_6350__bF_buf2), .C(_6377_), .Y(_1434_) );
NAND2X1 NAND2X1_419 ( .A(datapath_1_RegisterFile_regfile_mem_31__27_), .B(_6350__bF_buf3), .Y(_6378_) );
OAI21X1 OAI21X1_1312 ( .A(_5330__bF_buf0), .B(_6350__bF_buf3), .C(_6378_), .Y(_1435_) );
NAND2X1 NAND2X1_420 ( .A(datapath_1_RegisterFile_regfile_mem_31__28_), .B(_6350__bF_buf0), .Y(_6379_) );
OAI21X1 OAI21X1_1313 ( .A(_5332__bF_buf3), .B(_6350__bF_buf0), .C(_6379_), .Y(_1436_) );
NAND2X1 NAND2X1_421 ( .A(datapath_1_RegisterFile_regfile_mem_31__29_), .B(_6350__bF_buf7), .Y(_6380_) );
OAI21X1 OAI21X1_1314 ( .A(_5334__bF_buf0), .B(_6350__bF_buf7), .C(_6380_), .Y(_1437_) );
NAND2X1 NAND2X1_422 ( .A(datapath_1_RegisterFile_regfile_mem_31__30_), .B(_6350__bF_buf2), .Y(_6381_) );
OAI21X1 OAI21X1_1315 ( .A(_5336__bF_buf1), .B(_6350__bF_buf2), .C(_6381_), .Y(_1439_) );
NAND2X1 NAND2X1_423 ( .A(datapath_1_RegisterFile_regfile_mem_31__31_), .B(_6350__bF_buf3), .Y(_6382_) );
OAI21X1 OAI21X1_1316 ( .A(_5338__bF_buf4), .B(_6350__bF_buf3), .C(_6382_), .Y(_1860_) );
DFFPOSX1 DFFPOSX1_1 ( .CLK(clk_bF_buf111), .D(_1698_), .Q(datapath_1_RegisterFile_regfile_mem_12__0_) );
DFFPOSX1 DFFPOSX1_2 ( .CLK(clk_bF_buf107), .D(_1699_), .Q(datapath_1_RegisterFile_regfile_mem_12__1_) );
DFFPOSX1 DFFPOSX1_3 ( .CLK(clk_bF_buf33), .D(_1700_), .Q(datapath_1_RegisterFile_regfile_mem_12__2_) );
DFFPOSX1 DFFPOSX1_4 ( .CLK(clk_bF_buf62), .D(_1701_), .Q(datapath_1_RegisterFile_regfile_mem_12__3_) );
DFFPOSX1 DFFPOSX1_5 ( .CLK(clk_bF_buf111), .D(_1702_), .Q(datapath_1_RegisterFile_regfile_mem_12__4_) );
DFFPOSX1 DFFPOSX1_6 ( .CLK(clk_bF_buf102), .D(_940_), .Q(datapath_1_RegisterFile_regfile_mem_12__5_) );
DFFPOSX1 DFFPOSX1_7 ( .CLK(clk_bF_buf107), .D(_941_), .Q(datapath_1_RegisterFile_regfile_mem_12__6_) );
DFFPOSX1 DFFPOSX1_8 ( .CLK(clk_bF_buf64), .D(_942_), .Q(datapath_1_RegisterFile_regfile_mem_12__7_) );
DFFPOSX1 DFFPOSX1_9 ( .CLK(clk_bF_buf94), .D(_943_), .Q(datapath_1_RegisterFile_regfile_mem_12__8_) );
DFFPOSX1 DFFPOSX1_10 ( .CLK(clk_bF_buf20), .D(_944_), .Q(datapath_1_RegisterFile_regfile_mem_12__9_) );
DFFPOSX1 DFFPOSX1_11 ( .CLK(clk_bF_buf92), .D(_920_), .Q(datapath_1_RegisterFile_regfile_mem_12__10_) );
DFFPOSX1 DFFPOSX1_12 ( .CLK(clk_bF_buf54), .D(_921_), .Q(datapath_1_RegisterFile_regfile_mem_12__11_) );
DFFPOSX1 DFFPOSX1_13 ( .CLK(clk_bF_buf92), .D(_1703_), .Q(datapath_1_RegisterFile_regfile_mem_12__12_) );
DFFPOSX1 DFFPOSX1_14 ( .CLK(clk_bF_buf102), .D(_922_), .Q(datapath_1_RegisterFile_regfile_mem_12__13_) );
DFFPOSX1 DFFPOSX1_15 ( .CLK(clk_bF_buf15), .D(_923_), .Q(datapath_1_RegisterFile_regfile_mem_12__14_) );
DFFPOSX1 DFFPOSX1_16 ( .CLK(clk_bF_buf54), .D(_924_), .Q(datapath_1_RegisterFile_regfile_mem_12__15_) );
DFFPOSX1 DFFPOSX1_17 ( .CLK(clk_bF_buf55), .D(_925_), .Q(datapath_1_RegisterFile_regfile_mem_12__16_) );
DFFPOSX1 DFFPOSX1_18 ( .CLK(clk_bF_buf53), .D(_926_), .Q(datapath_1_RegisterFile_regfile_mem_12__17_) );
DFFPOSX1 DFFPOSX1_19 ( .CLK(clk_bF_buf16), .D(_927_), .Q(datapath_1_RegisterFile_regfile_mem_12__18_) );
DFFPOSX1 DFFPOSX1_20 ( .CLK(clk_bF_buf54), .D(_928_), .Q(datapath_1_RegisterFile_regfile_mem_12__19_) );
DFFPOSX1 DFFPOSX1_21 ( .CLK(clk_bF_buf62), .D(_929_), .Q(datapath_1_RegisterFile_regfile_mem_12__20_) );
DFFPOSX1 DFFPOSX1_22 ( .CLK(clk_bF_buf37), .D(_930_), .Q(datapath_1_RegisterFile_regfile_mem_12__21_) );
DFFPOSX1 DFFPOSX1_23 ( .CLK(clk_bF_buf45), .D(_1704_), .Q(datapath_1_RegisterFile_regfile_mem_12__22_) );
DFFPOSX1 DFFPOSX1_24 ( .CLK(clk_bF_buf20), .D(_931_), .Q(datapath_1_RegisterFile_regfile_mem_12__23_) );
DFFPOSX1 DFFPOSX1_25 ( .CLK(clk_bF_buf64), .D(_932_), .Q(datapath_1_RegisterFile_regfile_mem_12__24_) );
DFFPOSX1 DFFPOSX1_26 ( .CLK(clk_bF_buf33), .D(_933_), .Q(datapath_1_RegisterFile_regfile_mem_12__25_) );
DFFPOSX1 DFFPOSX1_27 ( .CLK(clk_bF_buf112), .D(_934_), .Q(datapath_1_RegisterFile_regfile_mem_12__26_) );
DFFPOSX1 DFFPOSX1_28 ( .CLK(clk_bF_buf15), .D(_935_), .Q(datapath_1_RegisterFile_regfile_mem_12__27_) );
DFFPOSX1 DFFPOSX1_29 ( .CLK(clk_bF_buf35), .D(_936_), .Q(datapath_1_RegisterFile_regfile_mem_12__28_) );
DFFPOSX1 DFFPOSX1_30 ( .CLK(clk_bF_buf101), .D(_937_), .Q(datapath_1_RegisterFile_regfile_mem_12__29_) );
DFFPOSX1 DFFPOSX1_31 ( .CLK(clk_bF_buf111), .D(_938_), .Q(datapath_1_RegisterFile_regfile_mem_12__30_) );
DFFPOSX1 DFFPOSX1_32 ( .CLK(clk_bF_buf20), .D(_939_), .Q(datapath_1_RegisterFile_regfile_mem_12__31_) );
DFFPOSX1 DFFPOSX1_33 ( .CLK(clk_bF_buf106), .D(_1218_), .Q(datapath_1_RegisterFile_regfile_mem_24__0_) );
DFFPOSX1 DFFPOSX1_34 ( .CLK(clk_bF_buf65), .D(_1227_), .Q(datapath_1_RegisterFile_regfile_mem_24__1_) );
DFFPOSX1 DFFPOSX1_35 ( .CLK(clk_bF_buf2), .D(_1229_), .Q(datapath_1_RegisterFile_regfile_mem_24__2_) );
DFFPOSX1 DFFPOSX1_36 ( .CLK(clk_bF_buf89), .D(_1232_), .Q(datapath_1_RegisterFile_regfile_mem_24__3_) );
DFFPOSX1 DFFPOSX1_37 ( .CLK(clk_bF_buf96), .D(_1233_), .Q(datapath_1_RegisterFile_regfile_mem_24__4_) );
DFFPOSX1 DFFPOSX1_38 ( .CLK(clk_bF_buf56), .D(_1234_), .Q(datapath_1_RegisterFile_regfile_mem_24__5_) );
DFFPOSX1 DFFPOSX1_39 ( .CLK(clk_bF_buf1), .D(_1805_), .Q(datapath_1_RegisterFile_regfile_mem_24__6_) );
DFFPOSX1 DFFPOSX1_40 ( .CLK(clk_bF_buf49), .D(_1235_), .Q(datapath_1_RegisterFile_regfile_mem_24__7_) );
DFFPOSX1 DFFPOSX1_41 ( .CLK(clk_bF_buf96), .D(_1236_), .Q(datapath_1_RegisterFile_regfile_mem_24__8_) );
DFFPOSX1 DFFPOSX1_42 ( .CLK(clk_bF_buf100), .D(_1237_), .Q(datapath_1_RegisterFile_regfile_mem_24__9_) );
DFFPOSX1 DFFPOSX1_43 ( .CLK(clk_bF_buf23), .D(_1219_), .Q(datapath_1_RegisterFile_regfile_mem_24__10_) );
DFFPOSX1 DFFPOSX1_44 ( .CLK(clk_bF_buf63), .D(_1220_), .Q(datapath_1_RegisterFile_regfile_mem_24__11_) );
DFFPOSX1 DFFPOSX1_45 ( .CLK(clk_bF_buf2), .D(_1221_), .Q(datapath_1_RegisterFile_regfile_mem_24__12_) );
DFFPOSX1 DFFPOSX1_46 ( .CLK(clk_bF_buf13), .D(_1222_), .Q(datapath_1_RegisterFile_regfile_mem_24__13_) );
DFFPOSX1 DFFPOSX1_47 ( .CLK(clk_bF_buf48), .D(_1223_), .Q(datapath_1_RegisterFile_regfile_mem_24__14_) );
DFFPOSX1 DFFPOSX1_48 ( .CLK(clk_bF_buf63), .D(_1224_), .Q(datapath_1_RegisterFile_regfile_mem_24__15_) );
DFFPOSX1 DFFPOSX1_49 ( .CLK(clk_bF_buf42), .D(_1806_), .Q(datapath_1_RegisterFile_regfile_mem_24__16_) );
DFFPOSX1 DFFPOSX1_50 ( .CLK(clk_bF_buf106), .D(_1225_), .Q(datapath_1_RegisterFile_regfile_mem_24__17_) );
DFFPOSX1 DFFPOSX1_51 ( .CLK(clk_bF_buf56), .D(_1226_), .Q(datapath_1_RegisterFile_regfile_mem_24__18_) );
DFFPOSX1 DFFPOSX1_52 ( .CLK(clk_bF_buf2), .D(_1807_), .Q(datapath_1_RegisterFile_regfile_mem_24__19_) );
DFFPOSX1 DFFPOSX1_53 ( .CLK(clk_bF_buf70), .D(_1808_), .Q(datapath_1_RegisterFile_regfile_mem_24__20_) );
DFFPOSX1 DFFPOSX1_54 ( .CLK(clk_bF_buf67), .D(_1809_), .Q(datapath_1_RegisterFile_regfile_mem_24__21_) );
DFFPOSX1 DFFPOSX1_55 ( .CLK(clk_bF_buf34), .D(_1810_), .Q(datapath_1_RegisterFile_regfile_mem_24__22_) );
DFFPOSX1 DFFPOSX1_56 ( .CLK(clk_bF_buf67), .D(_1811_), .Q(datapath_1_RegisterFile_regfile_mem_24__23_) );
DFFPOSX1 DFFPOSX1_57 ( .CLK(clk_bF_buf42), .D(_1812_), .Q(datapath_1_RegisterFile_regfile_mem_24__24_) );
DFFPOSX1 DFFPOSX1_58 ( .CLK(clk_bF_buf65), .D(_1813_), .Q(datapath_1_RegisterFile_regfile_mem_24__25_) );
DFFPOSX1 DFFPOSX1_59 ( .CLK(clk_bF_buf79), .D(_1814_), .Q(datapath_1_RegisterFile_regfile_mem_24__26_) );
DFFPOSX1 DFFPOSX1_60 ( .CLK(clk_bF_buf48), .D(_1815_), .Q(datapath_1_RegisterFile_regfile_mem_24__27_) );
DFFPOSX1 DFFPOSX1_61 ( .CLK(clk_bF_buf49), .D(_1816_), .Q(datapath_1_RegisterFile_regfile_mem_24__28_) );
DFFPOSX1 DFFPOSX1_62 ( .CLK(clk_bF_buf2), .D(_1228_), .Q(datapath_1_RegisterFile_regfile_mem_24__29_) );
DFFPOSX1 DFFPOSX1_63 ( .CLK(clk_bF_buf1), .D(_1230_), .Q(datapath_1_RegisterFile_regfile_mem_24__30_) );
DFFPOSX1 DFFPOSX1_64 ( .CLK(clk_bF_buf48), .D(_1231_), .Q(datapath_1_RegisterFile_regfile_mem_24__31_) );
DFFPOSX1 DFFPOSX1_65 ( .CLK(clk_bF_buf34), .D(_1761_), .Q(datapath_1_RegisterFile_regfile_mem_22__0_) );
DFFPOSX1 DFFPOSX1_66 ( .CLK(clk_bF_buf31), .D(_1762_), .Q(datapath_1_RegisterFile_regfile_mem_22__1_) );
DFFPOSX1 DFFPOSX1_67 ( .CLK(clk_bF_buf3), .D(_1763_), .Q(datapath_1_RegisterFile_regfile_mem_22__2_) );
DFFPOSX1 DFFPOSX1_68 ( .CLK(clk_bF_buf89), .D(_1764_), .Q(datapath_1_RegisterFile_regfile_mem_22__3_) );
DFFPOSX1 DFFPOSX1_69 ( .CLK(clk_bF_buf88), .D(_1765_), .Q(datapath_1_RegisterFile_regfile_mem_22__4_) );
DFFPOSX1 DFFPOSX1_70 ( .CLK(clk_bF_buf105), .D(_1766_), .Q(datapath_1_RegisterFile_regfile_mem_22__5_) );
DFFPOSX1 DFFPOSX1_71 ( .CLK(clk_bF_buf96), .D(_1767_), .Q(datapath_1_RegisterFile_regfile_mem_22__6_) );
DFFPOSX1 DFFPOSX1_72 ( .CLK(clk_bF_buf42), .D(_1768_), .Q(datapath_1_RegisterFile_regfile_mem_22__7_) );
DFFPOSX1 DFFPOSX1_73 ( .CLK(clk_bF_buf57), .D(_1769_), .Q(datapath_1_RegisterFile_regfile_mem_22__8_) );
DFFPOSX1 DFFPOSX1_74 ( .CLK(clk_bF_buf22), .D(_1770_), .Q(datapath_1_RegisterFile_regfile_mem_22__9_) );
DFFPOSX1 DFFPOSX1_75 ( .CLK(clk_bF_buf79), .D(_1771_), .Q(datapath_1_RegisterFile_regfile_mem_22__10_) );
DFFPOSX1 DFFPOSX1_76 ( .CLK(clk_bF_buf25), .D(_1772_), .Q(datapath_1_RegisterFile_regfile_mem_22__11_) );
DFFPOSX1 DFFPOSX1_77 ( .CLK(clk_bF_buf2), .D(_1773_), .Q(datapath_1_RegisterFile_regfile_mem_22__12_) );
DFFPOSX1 DFFPOSX1_78 ( .CLK(clk_bF_buf22), .D(_1774_), .Q(datapath_1_RegisterFile_regfile_mem_22__13_) );
DFFPOSX1 DFFPOSX1_79 ( .CLK(clk_bF_buf90), .D(_1775_), .Q(datapath_1_RegisterFile_regfile_mem_22__14_) );
DFFPOSX1 DFFPOSX1_80 ( .CLK(clk_bF_buf63), .D(_1776_), .Q(datapath_1_RegisterFile_regfile_mem_22__15_) );
DFFPOSX1 DFFPOSX1_81 ( .CLK(clk_bF_buf78), .D(_1777_), .Q(datapath_1_RegisterFile_regfile_mem_22__16_) );
DFFPOSX1 DFFPOSX1_82 ( .CLK(clk_bF_buf60), .D(_1778_), .Q(datapath_1_RegisterFile_regfile_mem_22__17_) );
DFFPOSX1 DFFPOSX1_83 ( .CLK(clk_bF_buf44), .D(_1779_), .Q(datapath_1_RegisterFile_regfile_mem_22__18_) );
DFFPOSX1 DFFPOSX1_84 ( .CLK(clk_bF_buf85), .D(_1780_), .Q(datapath_1_RegisterFile_regfile_mem_22__19_) );
DFFPOSX1 DFFPOSX1_85 ( .CLK(clk_bF_buf63), .D(_1781_), .Q(datapath_1_RegisterFile_regfile_mem_22__20_) );
DFFPOSX1 DFFPOSX1_86 ( .CLK(clk_bF_buf67), .D(_1782_), .Q(datapath_1_RegisterFile_regfile_mem_22__21_) );
DFFPOSX1 DFFPOSX1_87 ( .CLK(clk_bF_buf34), .D(_1783_), .Q(datapath_1_RegisterFile_regfile_mem_22__22_) );
DFFPOSX1 DFFPOSX1_88 ( .CLK(clk_bF_buf21), .D(_1784_), .Q(datapath_1_RegisterFile_regfile_mem_22__23_) );
DFFPOSX1 DFFPOSX1_89 ( .CLK(clk_bF_buf85), .D(_1785_), .Q(datapath_1_RegisterFile_regfile_mem_22__24_) );
DFFPOSX1 DFFPOSX1_90 ( .CLK(clk_bF_buf21), .D(_1786_), .Q(datapath_1_RegisterFile_regfile_mem_22__25_) );
DFFPOSX1 DFFPOSX1_91 ( .CLK(clk_bF_buf105), .D(_1787_), .Q(datapath_1_RegisterFile_regfile_mem_22__26_) );
DFFPOSX1 DFFPOSX1_92 ( .CLK(clk_bF_buf90), .D(_1788_), .Q(datapath_1_RegisterFile_regfile_mem_22__27_) );
DFFPOSX1 DFFPOSX1_93 ( .CLK(clk_bF_buf95), .D(_1789_), .Q(datapath_1_RegisterFile_regfile_mem_22__28_) );
DFFPOSX1 DFFPOSX1_94 ( .CLK(clk_bF_buf59), .D(_1790_), .Q(datapath_1_RegisterFile_regfile_mem_22__29_) );
DFFPOSX1 DFFPOSX1_95 ( .CLK(clk_bF_buf60), .D(_1791_), .Q(datapath_1_RegisterFile_regfile_mem_22__30_) );
DFFPOSX1 DFFPOSX1_96 ( .CLK(clk_bF_buf22), .D(_1792_), .Q(datapath_1_RegisterFile_regfile_mem_22__31_) );
DFFPOSX1 DFFPOSX1_97 ( .CLK(clk_bF_buf105), .D(_1178_), .Q(datapath_1_RegisterFile_regfile_mem_21__0_) );
DFFPOSX1 DFFPOSX1_98 ( .CLK(clk_bF_buf83), .D(_1179_), .Q(datapath_1_RegisterFile_regfile_mem_21__1_) );
DFFPOSX1 DFFPOSX1_99 ( .CLK(clk_bF_buf31), .D(_1189_), .Q(datapath_1_RegisterFile_regfile_mem_21__2_) );
DFFPOSX1 DFFPOSX1_100 ( .CLK(clk_bF_buf63), .D(_1192_), .Q(datapath_1_RegisterFile_regfile_mem_21__3_) );
DFFPOSX1 DFFPOSX1_101 ( .CLK(clk_bF_buf26), .D(_1193_), .Q(datapath_1_RegisterFile_regfile_mem_21__4_) );
DFFPOSX1 DFFPOSX1_102 ( .CLK(clk_bF_buf105), .D(_1194_), .Q(datapath_1_RegisterFile_regfile_mem_21__5_) );
DFFPOSX1 DFFPOSX1_103 ( .CLK(clk_bF_buf113), .D(_1195_), .Q(datapath_1_RegisterFile_regfile_mem_21__6_) );
DFFPOSX1 DFFPOSX1_104 ( .CLK(clk_bF_buf3), .D(_1749_), .Q(datapath_1_RegisterFile_regfile_mem_21__7_) );
DFFPOSX1 DFFPOSX1_105 ( .CLK(clk_bF_buf57), .D(_1196_), .Q(datapath_1_RegisterFile_regfile_mem_21__8_) );
DFFPOSX1 DFFPOSX1_106 ( .CLK(clk_bF_buf69), .D(_1197_), .Q(datapath_1_RegisterFile_regfile_mem_21__9_) );
DFFPOSX1 DFFPOSX1_107 ( .CLK(clk_bF_buf34), .D(_1750_), .Q(datapath_1_RegisterFile_regfile_mem_21__10_) );
DFFPOSX1 DFFPOSX1_108 ( .CLK(clk_bF_buf25), .D(_1751_), .Q(datapath_1_RegisterFile_regfile_mem_21__11_) );
DFFPOSX1 DFFPOSX1_109 ( .CLK(clk_bF_buf31), .D(_1752_), .Q(datapath_1_RegisterFile_regfile_mem_21__12_) );
DFFPOSX1 DFFPOSX1_110 ( .CLK(clk_bF_buf80), .D(_1753_), .Q(datapath_1_RegisterFile_regfile_mem_21__13_) );
DFFPOSX1 DFFPOSX1_111 ( .CLK(clk_bF_buf69), .D(_1754_), .Q(datapath_1_RegisterFile_regfile_mem_21__14_) );
DFFPOSX1 DFFPOSX1_112 ( .CLK(clk_bF_buf42), .D(_1755_), .Q(datapath_1_RegisterFile_regfile_mem_21__15_) );
DFFPOSX1 DFFPOSX1_113 ( .CLK(clk_bF_buf83), .D(_1756_), .Q(datapath_1_RegisterFile_regfile_mem_21__16_) );
DFFPOSX1 DFFPOSX1_114 ( .CLK(clk_bF_buf26), .D(_1757_), .Q(datapath_1_RegisterFile_regfile_mem_21__17_) );
DFFPOSX1 DFFPOSX1_115 ( .CLK(clk_bF_buf44), .D(_1758_), .Q(datapath_1_RegisterFile_regfile_mem_21__18_) );
DFFPOSX1 DFFPOSX1_116 ( .CLK(clk_bF_buf3), .D(_1759_), .Q(datapath_1_RegisterFile_regfile_mem_21__19_) );
DFFPOSX1 DFFPOSX1_117 ( .CLK(clk_bF_buf42), .D(_1180_), .Q(datapath_1_RegisterFile_regfile_mem_21__20_) );
DFFPOSX1 DFFPOSX1_118 ( .CLK(clk_bF_buf113), .D(_1181_), .Q(datapath_1_RegisterFile_regfile_mem_21__21_) );
DFFPOSX1 DFFPOSX1_119 ( .CLK(clk_bF_buf66), .D(_1182_), .Q(datapath_1_RegisterFile_regfile_mem_21__22_) );
DFFPOSX1 DFFPOSX1_120 ( .CLK(clk_bF_buf21), .D(_1183_), .Q(datapath_1_RegisterFile_regfile_mem_21__23_) );
DFFPOSX1 DFFPOSX1_121 ( .CLK(clk_bF_buf14), .D(_1184_), .Q(datapath_1_RegisterFile_regfile_mem_21__24_) );
DFFPOSX1 DFFPOSX1_122 ( .CLK(clk_bF_buf21), .D(_1185_), .Q(datapath_1_RegisterFile_regfile_mem_21__25_) );
DFFPOSX1 DFFPOSX1_123 ( .CLK(clk_bF_buf80), .D(_1186_), .Q(datapath_1_RegisterFile_regfile_mem_21__26_) );
DFFPOSX1 DFFPOSX1_124 ( .CLK(clk_bF_buf69), .D(_1760_), .Q(datapath_1_RegisterFile_regfile_mem_21__27_) );
DFFPOSX1 DFFPOSX1_125 ( .CLK(clk_bF_buf6), .D(_1187_), .Q(datapath_1_RegisterFile_regfile_mem_21__28_) );
DFFPOSX1 DFFPOSX1_126 ( .CLK(clk_bF_buf95), .D(_1188_), .Q(datapath_1_RegisterFile_regfile_mem_21__29_) );
DFFPOSX1 DFFPOSX1_127 ( .CLK(clk_bF_buf60), .D(_1190_), .Q(datapath_1_RegisterFile_regfile_mem_21__30_) );
DFFPOSX1 DFFPOSX1_128 ( .CLK(clk_bF_buf44), .D(_1191_), .Q(datapath_1_RegisterFile_regfile_mem_21__31_) );
DFFPOSX1 DFFPOSX1_129 ( .CLK(clk_bF_buf34), .D(_1149_), .Q(datapath_1_RegisterFile_regfile_mem_20__0_) );
DFFPOSX1 DFFPOSX1_130 ( .CLK(clk_bF_buf78), .D(_1159_), .Q(datapath_1_RegisterFile_regfile_mem_20__1_) );
DFFPOSX1 DFFPOSX1_131 ( .CLK(clk_bF_buf38), .D(_1746_), .Q(datapath_1_RegisterFile_regfile_mem_20__2_) );
DFFPOSX1 DFFPOSX1_132 ( .CLK(clk_bF_buf63), .D(_1171_), .Q(datapath_1_RegisterFile_regfile_mem_20__3_) );
DFFPOSX1 DFFPOSX1_133 ( .CLK(clk_bF_buf76), .D(_1172_), .Q(datapath_1_RegisterFile_regfile_mem_20__4_) );
DFFPOSX1 DFFPOSX1_134 ( .CLK(clk_bF_buf80), .D(_1173_), .Q(datapath_1_RegisterFile_regfile_mem_20__5_) );
DFFPOSX1 DFFPOSX1_135 ( .CLK(clk_bF_buf113), .D(_1174_), .Q(datapath_1_RegisterFile_regfile_mem_20__6_) );
DFFPOSX1 DFFPOSX1_136 ( .CLK(clk_bF_buf63), .D(_1175_), .Q(datapath_1_RegisterFile_regfile_mem_20__7_) );
DFFPOSX1 DFFPOSX1_137 ( .CLK(clk_bF_buf26), .D(_1176_), .Q(datapath_1_RegisterFile_regfile_mem_20__8_) );
DFFPOSX1 DFFPOSX1_138 ( .CLK(clk_bF_buf90), .D(_1177_), .Q(datapath_1_RegisterFile_regfile_mem_20__9_) );
DFFPOSX1 DFFPOSX1_139 ( .CLK(clk_bF_buf13), .D(_1150_), .Q(datapath_1_RegisterFile_regfile_mem_20__10_) );
DFFPOSX1 DFFPOSX1_140 ( .CLK(clk_bF_buf85), .D(_1151_), .Q(datapath_1_RegisterFile_regfile_mem_20__11_) );
DFFPOSX1 DFFPOSX1_141 ( .CLK(clk_bF_buf21), .D(_1747_), .Q(datapath_1_RegisterFile_regfile_mem_20__12_) );
DFFPOSX1 DFFPOSX1_142 ( .CLK(clk_bF_buf44), .D(_1152_), .Q(datapath_1_RegisterFile_regfile_mem_20__13_) );
DFFPOSX1 DFFPOSX1_143 ( .CLK(clk_bF_buf44), .D(_1153_), .Q(datapath_1_RegisterFile_regfile_mem_20__14_) );
DFFPOSX1 DFFPOSX1_144 ( .CLK(clk_bF_buf63), .D(_1154_), .Q(datapath_1_RegisterFile_regfile_mem_20__15_) );
DFFPOSX1 DFFPOSX1_145 ( .CLK(clk_bF_buf78), .D(_1155_), .Q(datapath_1_RegisterFile_regfile_mem_20__16_) );
DFFPOSX1 DFFPOSX1_146 ( .CLK(clk_bF_buf76), .D(_1156_), .Q(datapath_1_RegisterFile_regfile_mem_20__17_) );
DFFPOSX1 DFFPOSX1_147 ( .CLK(clk_bF_buf4), .D(_1157_), .Q(datapath_1_RegisterFile_regfile_mem_20__18_) );
DFFPOSX1 DFFPOSX1_148 ( .CLK(clk_bF_buf85), .D(_1158_), .Q(datapath_1_RegisterFile_regfile_mem_20__19_) );
DFFPOSX1 DFFPOSX1_149 ( .CLK(clk_bF_buf42), .D(_1160_), .Q(datapath_1_RegisterFile_regfile_mem_20__20_) );
DFFPOSX1 DFFPOSX1_150 ( .CLK(clk_bF_buf26), .D(_1161_), .Q(datapath_1_RegisterFile_regfile_mem_20__21_) );
DFFPOSX1 DFFPOSX1_151 ( .CLK(clk_bF_buf66), .D(_1748_), .Q(datapath_1_RegisterFile_regfile_mem_20__22_) );
DFFPOSX1 DFFPOSX1_152 ( .CLK(clk_bF_buf67), .D(_1162_), .Q(datapath_1_RegisterFile_regfile_mem_20__23_) );
DFFPOSX1 DFFPOSX1_153 ( .CLK(clk_bF_buf85), .D(_1163_), .Q(datapath_1_RegisterFile_regfile_mem_20__24_) );
DFFPOSX1 DFFPOSX1_154 ( .CLK(clk_bF_buf21), .D(_1164_), .Q(datapath_1_RegisterFile_regfile_mem_20__25_) );
DFFPOSX1 DFFPOSX1_155 ( .CLK(clk_bF_buf105), .D(_1165_), .Q(datapath_1_RegisterFile_regfile_mem_20__26_) );
DFFPOSX1 DFFPOSX1_156 ( .CLK(clk_bF_buf90), .D(_1166_), .Q(datapath_1_RegisterFile_regfile_mem_20__27_) );
DFFPOSX1 DFFPOSX1_157 ( .CLK(clk_bF_buf59), .D(_1167_), .Q(datapath_1_RegisterFile_regfile_mem_20__28_) );
DFFPOSX1 DFFPOSX1_158 ( .CLK(clk_bF_buf95), .D(_1168_), .Q(datapath_1_RegisterFile_regfile_mem_20__29_) );
DFFPOSX1 DFFPOSX1_159 ( .CLK(clk_bF_buf60), .D(_1169_), .Q(datapath_1_RegisterFile_regfile_mem_20__30_) );
DFFPOSX1 DFFPOSX1_160 ( .CLK(clk_bF_buf22), .D(_1170_), .Q(datapath_1_RegisterFile_regfile_mem_20__31_) );
DFFPOSX1 DFFPOSX1_161 ( .CLK(clk_bF_buf105), .D(_1099_), .Q(datapath_1_RegisterFile_regfile_mem_19__0_) );
DFFPOSX1 DFFPOSX1_162 ( .CLK(clk_bF_buf14), .D(_1109_), .Q(datapath_1_RegisterFile_regfile_mem_19__1_) );
DFFPOSX1 DFFPOSX1_163 ( .CLK(clk_bF_buf85), .D(_1119_), .Q(datapath_1_RegisterFile_regfile_mem_19__2_) );
DFFPOSX1 DFFPOSX1_164 ( .CLK(clk_bF_buf6), .D(_1122_), .Q(datapath_1_RegisterFile_regfile_mem_19__3_) );
DFFPOSX1 DFFPOSX1_165 ( .CLK(clk_bF_buf26), .D(_1123_), .Q(datapath_1_RegisterFile_regfile_mem_19__4_) );
DFFPOSX1 DFFPOSX1_166 ( .CLK(clk_bF_buf80), .D(_1124_), .Q(datapath_1_RegisterFile_regfile_mem_19__5_) );
DFFPOSX1 DFFPOSX1_167 ( .CLK(clk_bF_buf65), .D(_1125_), .Q(datapath_1_RegisterFile_regfile_mem_19__6_) );
DFFPOSX1 DFFPOSX1_168 ( .CLK(clk_bF_buf25), .D(_1743_), .Q(datapath_1_RegisterFile_regfile_mem_19__7_) );
DFFPOSX1 DFFPOSX1_169 ( .CLK(clk_bF_buf96), .D(_1126_), .Q(datapath_1_RegisterFile_regfile_mem_19__8_) );
DFFPOSX1 DFFPOSX1_170 ( .CLK(clk_bF_buf69), .D(_1127_), .Q(datapath_1_RegisterFile_regfile_mem_19__9_) );
DFFPOSX1 DFFPOSX1_171 ( .CLK(clk_bF_buf80), .D(_1100_), .Q(datapath_1_RegisterFile_regfile_mem_19__10_) );
DFFPOSX1 DFFPOSX1_172 ( .CLK(clk_bF_buf85), .D(_1101_), .Q(datapath_1_RegisterFile_regfile_mem_19__11_) );
DFFPOSX1 DFFPOSX1_173 ( .CLK(clk_bF_buf31), .D(_1102_), .Q(datapath_1_RegisterFile_regfile_mem_19__12_) );
DFFPOSX1 DFFPOSX1_174 ( .CLK(clk_bF_buf44), .D(_1103_), .Q(datapath_1_RegisterFile_regfile_mem_19__13_) );
DFFPOSX1 DFFPOSX1_175 ( .CLK(clk_bF_buf44), .D(_1104_), .Q(datapath_1_RegisterFile_regfile_mem_19__14_) );
DFFPOSX1 DFFPOSX1_176 ( .CLK(clk_bF_buf75), .D(_1105_), .Q(datapath_1_RegisterFile_regfile_mem_19__15_) );
DFFPOSX1 DFFPOSX1_177 ( .CLK(clk_bF_buf59), .D(_1106_), .Q(datapath_1_RegisterFile_regfile_mem_19__16_) );
DFFPOSX1 DFFPOSX1_178 ( .CLK(clk_bF_buf88), .D(_1744_), .Q(datapath_1_RegisterFile_regfile_mem_19__17_) );
DFFPOSX1 DFFPOSX1_179 ( .CLK(clk_bF_buf80), .D(_1107_), .Q(datapath_1_RegisterFile_regfile_mem_19__18_) );
DFFPOSX1 DFFPOSX1_180 ( .CLK(clk_bF_buf75), .D(_1108_), .Q(datapath_1_RegisterFile_regfile_mem_19__19_) );
DFFPOSX1 DFFPOSX1_181 ( .CLK(clk_bF_buf6), .D(_1110_), .Q(datapath_1_RegisterFile_regfile_mem_19__20_) );
DFFPOSX1 DFFPOSX1_182 ( .CLK(clk_bF_buf57), .D(_1111_), .Q(datapath_1_RegisterFile_regfile_mem_19__21_) );
DFFPOSX1 DFFPOSX1_183 ( .CLK(clk_bF_buf66), .D(_1112_), .Q(datapath_1_RegisterFile_regfile_mem_19__22_) );
DFFPOSX1 DFFPOSX1_184 ( .CLK(clk_bF_buf113), .D(_1113_), .Q(datapath_1_RegisterFile_regfile_mem_19__23_) );
DFFPOSX1 DFFPOSX1_185 ( .CLK(clk_bF_buf75), .D(_1114_), .Q(datapath_1_RegisterFile_regfile_mem_19__24_) );
DFFPOSX1 DFFPOSX1_186 ( .CLK(clk_bF_buf14), .D(_1115_), .Q(datapath_1_RegisterFile_regfile_mem_19__25_) );
DFFPOSX1 DFFPOSX1_187 ( .CLK(clk_bF_buf105), .D(_1116_), .Q(datapath_1_RegisterFile_regfile_mem_19__26_) );
DFFPOSX1 DFFPOSX1_188 ( .CLK(clk_bF_buf22), .D(_1745_), .Q(datapath_1_RegisterFile_regfile_mem_19__27_) );
DFFPOSX1 DFFPOSX1_189 ( .CLK(clk_bF_buf6), .D(_1117_), .Q(datapath_1_RegisterFile_regfile_mem_19__28_) );
DFFPOSX1 DFFPOSX1_190 ( .CLK(clk_bF_buf38), .D(_1118_), .Q(datapath_1_RegisterFile_regfile_mem_19__29_) );
DFFPOSX1 DFFPOSX1_191 ( .CLK(clk_bF_buf60), .D(_1120_), .Q(datapath_1_RegisterFile_regfile_mem_19__30_) );
DFFPOSX1 DFFPOSX1_192 ( .CLK(clk_bF_buf69), .D(_1121_), .Q(datapath_1_RegisterFile_regfile_mem_19__31_) );
DFFPOSX1 DFFPOSX1_193 ( .CLK(clk_bF_buf66), .D(_1079_), .Q(datapath_1_RegisterFile_regfile_mem_18__0_) );
DFFPOSX1 DFFPOSX1_194 ( .CLK(clk_bF_buf14), .D(_1085_), .Q(datapath_1_RegisterFile_regfile_mem_18__1_) );
DFFPOSX1 DFFPOSX1_195 ( .CLK(clk_bF_buf75), .D(_1731_), .Q(datapath_1_RegisterFile_regfile_mem_18__2_) );
DFFPOSX1 DFFPOSX1_196 ( .CLK(clk_bF_buf42), .D(_1097_), .Q(datapath_1_RegisterFile_regfile_mem_18__3_) );
DFFPOSX1 DFFPOSX1_197 ( .CLK(clk_bF_buf88), .D(_1098_), .Q(datapath_1_RegisterFile_regfile_mem_18__4_) );
DFFPOSX1 DFFPOSX1_198 ( .CLK(clk_bF_buf90), .D(_1732_), .Q(datapath_1_RegisterFile_regfile_mem_18__5_) );
DFFPOSX1 DFFPOSX1_199 ( .CLK(clk_bF_buf58), .D(_1733_), .Q(datapath_1_RegisterFile_regfile_mem_18__6_) );
DFFPOSX1 DFFPOSX1_200 ( .CLK(clk_bF_buf6), .D(_1734_), .Q(datapath_1_RegisterFile_regfile_mem_18__7_) );
DFFPOSX1 DFFPOSX1_201 ( .CLK(clk_bF_buf57), .D(_1735_), .Q(datapath_1_RegisterFile_regfile_mem_18__8_) );
DFFPOSX1 DFFPOSX1_202 ( .CLK(clk_bF_buf22), .D(_1736_), .Q(datapath_1_RegisterFile_regfile_mem_18__9_) );
DFFPOSX1 DFFPOSX1_203 ( .CLK(clk_bF_buf44), .D(_1737_), .Q(datapath_1_RegisterFile_regfile_mem_18__10_) );
DFFPOSX1 DFFPOSX1_204 ( .CLK(clk_bF_buf25), .D(_1738_), .Q(datapath_1_RegisterFile_regfile_mem_18__11_) );
DFFPOSX1 DFFPOSX1_205 ( .CLK(clk_bF_buf41), .D(_1739_), .Q(datapath_1_RegisterFile_regfile_mem_18__12_) );
DFFPOSX1 DFFPOSX1_206 ( .CLK(clk_bF_buf44), .D(_1740_), .Q(datapath_1_RegisterFile_regfile_mem_18__13_) );
DFFPOSX1 DFFPOSX1_207 ( .CLK(clk_bF_buf9), .D(_1741_), .Q(datapath_1_RegisterFile_regfile_mem_18__14_) );
DFFPOSX1 DFFPOSX1_208 ( .CLK(clk_bF_buf75), .D(_1080_), .Q(datapath_1_RegisterFile_regfile_mem_18__15_) );
DFFPOSX1 DFFPOSX1_209 ( .CLK(clk_bF_buf78), .D(_1081_), .Q(datapath_1_RegisterFile_regfile_mem_18__16_) );
DFFPOSX1 DFFPOSX1_210 ( .CLK(clk_bF_buf60), .D(_1082_), .Q(datapath_1_RegisterFile_regfile_mem_18__17_) );
DFFPOSX1 DFFPOSX1_211 ( .CLK(clk_bF_buf90), .D(_1083_), .Q(datapath_1_RegisterFile_regfile_mem_18__18_) );
DFFPOSX1 DFFPOSX1_212 ( .CLK(clk_bF_buf3), .D(_1084_), .Q(datapath_1_RegisterFile_regfile_mem_18__19_) );
DFFPOSX1 DFFPOSX1_213 ( .CLK(clk_bF_buf6), .D(_1086_), .Q(datapath_1_RegisterFile_regfile_mem_18__20_) );
DFFPOSX1 DFFPOSX1_214 ( .CLK(clk_bF_buf57), .D(_1087_), .Q(datapath_1_RegisterFile_regfile_mem_18__21_) );
DFFPOSX1 DFFPOSX1_215 ( .CLK(clk_bF_buf66), .D(_1742_), .Q(datapath_1_RegisterFile_regfile_mem_18__22_) );
DFFPOSX1 DFFPOSX1_216 ( .CLK(clk_bF_buf21), .D(_1088_), .Q(datapath_1_RegisterFile_regfile_mem_18__23_) );
DFFPOSX1 DFFPOSX1_217 ( .CLK(clk_bF_buf14), .D(_1089_), .Q(datapath_1_RegisterFile_regfile_mem_18__24_) );
DFFPOSX1 DFFPOSX1_218 ( .CLK(clk_bF_buf38), .D(_1090_), .Q(datapath_1_RegisterFile_regfile_mem_18__25_) );
DFFPOSX1 DFFPOSX1_219 ( .CLK(clk_bF_buf47), .D(_1091_), .Q(datapath_1_RegisterFile_regfile_mem_18__26_) );
DFFPOSX1 DFFPOSX1_220 ( .CLK(clk_bF_buf22), .D(_1092_), .Q(datapath_1_RegisterFile_regfile_mem_18__27_) );
DFFPOSX1 DFFPOSX1_221 ( .CLK(clk_bF_buf75), .D(_1093_), .Q(datapath_1_RegisterFile_regfile_mem_18__28_) );
DFFPOSX1 DFFPOSX1_222 ( .CLK(clk_bF_buf78), .D(_1094_), .Q(datapath_1_RegisterFile_regfile_mem_18__29_) );
DFFPOSX1 DFFPOSX1_223 ( .CLK(clk_bF_buf60), .D(_1095_), .Q(datapath_1_RegisterFile_regfile_mem_18__30_) );
DFFPOSX1 DFFPOSX1_224 ( .CLK(clk_bF_buf9), .D(_1096_), .Q(datapath_1_RegisterFile_regfile_mem_18__31_) );
DFFPOSX1 DFFPOSX1_225 ( .CLK(clk_bF_buf47), .D(_1050_), .Q(datapath_1_RegisterFile_regfile_mem_17__0_) );
DFFPOSX1 DFFPOSX1_226 ( .CLK(clk_bF_buf14), .D(_1060_), .Q(datapath_1_RegisterFile_regfile_mem_17__1_) );
DFFPOSX1 DFFPOSX1_227 ( .CLK(clk_bF_buf14), .D(_1070_), .Q(datapath_1_RegisterFile_regfile_mem_17__2_) );
DFFPOSX1 DFFPOSX1_228 ( .CLK(clk_bF_buf42), .D(_1073_), .Q(datapath_1_RegisterFile_regfile_mem_17__3_) );
DFFPOSX1 DFFPOSX1_229 ( .CLK(clk_bF_buf26), .D(_1074_), .Q(datapath_1_RegisterFile_regfile_mem_17__4_) );
DFFPOSX1 DFFPOSX1_230 ( .CLK(clk_bF_buf22), .D(_1075_), .Q(datapath_1_RegisterFile_regfile_mem_17__5_) );
DFFPOSX1 DFFPOSX1_231 ( .CLK(clk_bF_buf65), .D(_1076_), .Q(datapath_1_RegisterFile_regfile_mem_17__6_) );
DFFPOSX1 DFFPOSX1_232 ( .CLK(clk_bF_buf75), .D(_1728_), .Q(datapath_1_RegisterFile_regfile_mem_17__7_) );
DFFPOSX1 DFFPOSX1_233 ( .CLK(clk_bF_buf96), .D(_1077_), .Q(datapath_1_RegisterFile_regfile_mem_17__8_) );
DFFPOSX1 DFFPOSX1_234 ( .CLK(clk_bF_buf9), .D(_1078_), .Q(datapath_1_RegisterFile_regfile_mem_17__9_) );
DFFPOSX1 DFFPOSX1_235 ( .CLK(clk_bF_buf80), .D(_1051_), .Q(datapath_1_RegisterFile_regfile_mem_17__10_) );
DFFPOSX1 DFFPOSX1_236 ( .CLK(clk_bF_buf25), .D(_1052_), .Q(datapath_1_RegisterFile_regfile_mem_17__11_) );
DFFPOSX1 DFFPOSX1_237 ( .CLK(clk_bF_buf59), .D(_1053_), .Q(datapath_1_RegisterFile_regfile_mem_17__12_) );
DFFPOSX1 DFFPOSX1_238 ( .CLK(clk_bF_buf69), .D(_1054_), .Q(datapath_1_RegisterFile_regfile_mem_17__13_) );
DFFPOSX1 DFFPOSX1_239 ( .CLK(clk_bF_buf69), .D(_1055_), .Q(datapath_1_RegisterFile_regfile_mem_17__14_) );
DFFPOSX1 DFFPOSX1_240 ( .CLK(clk_bF_buf75), .D(_1056_), .Q(datapath_1_RegisterFile_regfile_mem_17__15_) );
DFFPOSX1 DFFPOSX1_241 ( .CLK(clk_bF_buf95), .D(_1057_), .Q(datapath_1_RegisterFile_regfile_mem_17__16_) );
DFFPOSX1 DFFPOSX1_242 ( .CLK(clk_bF_buf88), .D(_1729_), .Q(datapath_1_RegisterFile_regfile_mem_17__17_) );
DFFPOSX1 DFFPOSX1_243 ( .CLK(clk_bF_buf22), .D(_1058_), .Q(datapath_1_RegisterFile_regfile_mem_17__18_) );
DFFPOSX1 DFFPOSX1_244 ( .CLK(clk_bF_buf25), .D(_1059_), .Q(datapath_1_RegisterFile_regfile_mem_17__19_) );
DFFPOSX1 DFFPOSX1_245 ( .CLK(clk_bF_buf6), .D(_1061_), .Q(datapath_1_RegisterFile_regfile_mem_17__20_) );
DFFPOSX1 DFFPOSX1_246 ( .CLK(clk_bF_buf57), .D(_1062_), .Q(datapath_1_RegisterFile_regfile_mem_17__21_) );
DFFPOSX1 DFFPOSX1_247 ( .CLK(clk_bF_buf66), .D(_1063_), .Q(datapath_1_RegisterFile_regfile_mem_17__22_) );
DFFPOSX1 DFFPOSX1_248 ( .CLK(clk_bF_buf58), .D(_1064_), .Q(datapath_1_RegisterFile_regfile_mem_17__23_) );
DFFPOSX1 DFFPOSX1_249 ( .CLK(clk_bF_buf38), .D(_1065_), .Q(datapath_1_RegisterFile_regfile_mem_17__24_) );
DFFPOSX1 DFFPOSX1_250 ( .CLK(clk_bF_buf85), .D(_1066_), .Q(datapath_1_RegisterFile_regfile_mem_17__25_) );
DFFPOSX1 DFFPOSX1_251 ( .CLK(clk_bF_buf47), .D(_1067_), .Q(datapath_1_RegisterFile_regfile_mem_17__26_) );
DFFPOSX1 DFFPOSX1_252 ( .CLK(clk_bF_buf9), .D(_1730_), .Q(datapath_1_RegisterFile_regfile_mem_17__27_) );
DFFPOSX1 DFFPOSX1_253 ( .CLK(clk_bF_buf38), .D(_1068_), .Q(datapath_1_RegisterFile_regfile_mem_17__28_) );
DFFPOSX1 DFFPOSX1_254 ( .CLK(clk_bF_buf14), .D(_1069_), .Q(datapath_1_RegisterFile_regfile_mem_17__29_) );
DFFPOSX1 DFFPOSX1_255 ( .CLK(clk_bF_buf88), .D(_1071_), .Q(datapath_1_RegisterFile_regfile_mem_17__30_) );
DFFPOSX1 DFFPOSX1_256 ( .CLK(clk_bF_buf9), .D(_1072_), .Q(datapath_1_RegisterFile_regfile_mem_17__31_) );
DFFPOSX1 DFFPOSX1_257 ( .CLK(clk_bF_buf47), .D(_1021_), .Q(datapath_1_RegisterFile_regfile_mem_16__0_) );
DFFPOSX1 DFFPOSX1_258 ( .CLK(clk_bF_buf38), .D(_1031_), .Q(datapath_1_RegisterFile_regfile_mem_16__1_) );
DFFPOSX1 DFFPOSX1_259 ( .CLK(clk_bF_buf59), .D(_1725_), .Q(datapath_1_RegisterFile_regfile_mem_16__2_) );
DFFPOSX1 DFFPOSX1_260 ( .CLK(clk_bF_buf42), .D(_1043_), .Q(datapath_1_RegisterFile_regfile_mem_16__3_) );
DFFPOSX1 DFFPOSX1_261 ( .CLK(clk_bF_buf76), .D(_1044_), .Q(datapath_1_RegisterFile_regfile_mem_16__4_) );
DFFPOSX1 DFFPOSX1_262 ( .CLK(clk_bF_buf105), .D(_1045_), .Q(datapath_1_RegisterFile_regfile_mem_16__5_) );
DFFPOSX1 DFFPOSX1_263 ( .CLK(clk_bF_buf58), .D(_1046_), .Q(datapath_1_RegisterFile_regfile_mem_16__6_) );
DFFPOSX1 DFFPOSX1_264 ( .CLK(clk_bF_buf25), .D(_1047_), .Q(datapath_1_RegisterFile_regfile_mem_16__7_) );
DFFPOSX1 DFFPOSX1_265 ( .CLK(clk_bF_buf113), .D(_1048_), .Q(datapath_1_RegisterFile_regfile_mem_16__8_) );
DFFPOSX1 DFFPOSX1_266 ( .CLK(clk_bF_buf69), .D(_1049_), .Q(datapath_1_RegisterFile_regfile_mem_16__9_) );
DFFPOSX1 DFFPOSX1_267 ( .CLK(clk_bF_buf44), .D(_1022_), .Q(datapath_1_RegisterFile_regfile_mem_16__10_) );
DFFPOSX1 DFFPOSX1_268 ( .CLK(clk_bF_buf25), .D(_1023_), .Q(datapath_1_RegisterFile_regfile_mem_16__11_) );
DFFPOSX1 DFFPOSX1_269 ( .CLK(clk_bF_buf40), .D(_1726_), .Q(datapath_1_RegisterFile_regfile_mem_16__12_) );
DFFPOSX1 DFFPOSX1_270 ( .CLK(clk_bF_buf22), .D(_1024_), .Q(datapath_1_RegisterFile_regfile_mem_16__13_) );
DFFPOSX1 DFFPOSX1_271 ( .CLK(clk_bF_buf69), .D(_1025_), .Q(datapath_1_RegisterFile_regfile_mem_16__14_) );
DFFPOSX1 DFFPOSX1_272 ( .CLK(clk_bF_buf75), .D(_1026_), .Q(datapath_1_RegisterFile_regfile_mem_16__15_) );
DFFPOSX1 DFFPOSX1_273 ( .CLK(clk_bF_buf78), .D(_1027_), .Q(datapath_1_RegisterFile_regfile_mem_16__16_) );
DFFPOSX1 DFFPOSX1_274 ( .CLK(clk_bF_buf60), .D(_1028_), .Q(datapath_1_RegisterFile_regfile_mem_16__17_) );
DFFPOSX1 DFFPOSX1_275 ( .CLK(clk_bF_buf90), .D(_1029_), .Q(datapath_1_RegisterFile_regfile_mem_16__18_) );
DFFPOSX1 DFFPOSX1_276 ( .CLK(clk_bF_buf25), .D(_1030_), .Q(datapath_1_RegisterFile_regfile_mem_16__19_) );
DFFPOSX1 DFFPOSX1_277 ( .CLK(clk_bF_buf6), .D(_1032_), .Q(datapath_1_RegisterFile_regfile_mem_16__20_) );
DFFPOSX1 DFFPOSX1_278 ( .CLK(clk_bF_buf113), .D(_1033_), .Q(datapath_1_RegisterFile_regfile_mem_16__21_) );
DFFPOSX1 DFFPOSX1_279 ( .CLK(clk_bF_buf66), .D(_1727_), .Q(datapath_1_RegisterFile_regfile_mem_16__22_) );
DFFPOSX1 DFFPOSX1_280 ( .CLK(clk_bF_buf96), .D(_1034_), .Q(datapath_1_RegisterFile_regfile_mem_16__23_) );
DFFPOSX1 DFFPOSX1_281 ( .CLK(clk_bF_buf38), .D(_1035_), .Q(datapath_1_RegisterFile_regfile_mem_16__24_) );
DFFPOSX1 DFFPOSX1_282 ( .CLK(clk_bF_buf38), .D(_1036_), .Q(datapath_1_RegisterFile_regfile_mem_16__25_) );
DFFPOSX1 DFFPOSX1_283 ( .CLK(clk_bF_buf47), .D(_1037_), .Q(datapath_1_RegisterFile_regfile_mem_16__26_) );
DFFPOSX1 DFFPOSX1_284 ( .CLK(clk_bF_buf69), .D(_1038_), .Q(datapath_1_RegisterFile_regfile_mem_16__27_) );
DFFPOSX1 DFFPOSX1_285 ( .CLK(clk_bF_buf85), .D(_1039_), .Q(datapath_1_RegisterFile_regfile_mem_16__28_) );
DFFPOSX1 DFFPOSX1_286 ( .CLK(clk_bF_buf31), .D(_1040_), .Q(datapath_1_RegisterFile_regfile_mem_16__29_) );
DFFPOSX1 DFFPOSX1_287 ( .CLK(clk_bF_buf88), .D(_1041_), .Q(datapath_1_RegisterFile_regfile_mem_16__30_) );
DFFPOSX1 DFFPOSX1_288 ( .CLK(clk_bF_buf69), .D(_1042_), .Q(datapath_1_RegisterFile_regfile_mem_16__31_) );
DFFPOSX1 DFFPOSX1_289 ( .CLK(clk_bF_buf15), .D(_1713_), .Q(datapath_1_RegisterFile_regfile_mem_15__0_) );
DFFPOSX1 DFFPOSX1_290 ( .CLK(clk_bF_buf39), .D(_1714_), .Q(datapath_1_RegisterFile_regfile_mem_15__1_) );
DFFPOSX1 DFFPOSX1_291 ( .CLK(clk_bF_buf93), .D(_1715_), .Q(datapath_1_RegisterFile_regfile_mem_15__2_) );
DFFPOSX1 DFFPOSX1_292 ( .CLK(clk_bF_buf39), .D(_1716_), .Q(datapath_1_RegisterFile_regfile_mem_15__3_) );
DFFPOSX1 DFFPOSX1_293 ( .CLK(clk_bF_buf37), .D(_1717_), .Q(datapath_1_RegisterFile_regfile_mem_15__4_) );
DFFPOSX1 DFFPOSX1_294 ( .CLK(clk_bF_buf11), .D(_1718_), .Q(datapath_1_RegisterFile_regfile_mem_15__5_) );
DFFPOSX1 DFFPOSX1_295 ( .CLK(clk_bF_buf93), .D(_1719_), .Q(datapath_1_RegisterFile_regfile_mem_15__6_) );
DFFPOSX1 DFFPOSX1_296 ( .CLK(clk_bF_buf55), .D(_1720_), .Q(datapath_1_RegisterFile_regfile_mem_15__7_) );
DFFPOSX1 DFFPOSX1_297 ( .CLK(clk_bF_buf94), .D(_1721_), .Q(datapath_1_RegisterFile_regfile_mem_15__8_) );
DFFPOSX1 DFFPOSX1_298 ( .CLK(clk_bF_buf72), .D(_1722_), .Q(datapath_1_RegisterFile_regfile_mem_15__9_) );
DFFPOSX1 DFFPOSX1_299 ( .CLK(clk_bF_buf94), .D(_1001_), .Q(datapath_1_RegisterFile_regfile_mem_15__10_) );
DFFPOSX1 DFFPOSX1_300 ( .CLK(clk_bF_buf55), .D(_1002_), .Q(datapath_1_RegisterFile_regfile_mem_15__11_) );
DFFPOSX1 DFFPOSX1_301 ( .CLK(clk_bF_buf94), .D(_1003_), .Q(datapath_1_RegisterFile_regfile_mem_15__12_) );
DFFPOSX1 DFFPOSX1_302 ( .CLK(clk_bF_buf16), .D(_1004_), .Q(datapath_1_RegisterFile_regfile_mem_15__13_) );
DFFPOSX1 DFFPOSX1_303 ( .CLK(clk_bF_buf15), .D(_1005_), .Q(datapath_1_RegisterFile_regfile_mem_15__14_) );
DFFPOSX1 DFFPOSX1_304 ( .CLK(clk_bF_buf64), .D(_1006_), .Q(datapath_1_RegisterFile_regfile_mem_15__15_) );
DFFPOSX1 DFFPOSX1_305 ( .CLK(clk_bF_buf35), .D(_1007_), .Q(datapath_1_RegisterFile_regfile_mem_15__16_) );
DFFPOSX1 DFFPOSX1_306 ( .CLK(clk_bF_buf15), .D(_1723_), .Q(datapath_1_RegisterFile_regfile_mem_15__17_) );
DFFPOSX1 DFFPOSX1_307 ( .CLK(clk_bF_buf102), .D(_1008_), .Q(datapath_1_RegisterFile_regfile_mem_15__18_) );
DFFPOSX1 DFFPOSX1_308 ( .CLK(clk_bF_buf84), .D(_1009_), .Q(datapath_1_RegisterFile_regfile_mem_15__19_) );
DFFPOSX1 DFFPOSX1_309 ( .CLK(clk_bF_buf84), .D(_1010_), .Q(datapath_1_RegisterFile_regfile_mem_15__20_) );
DFFPOSX1 DFFPOSX1_310 ( .CLK(clk_bF_buf37), .D(_1011_), .Q(datapath_1_RegisterFile_regfile_mem_15__21_) );
DFFPOSX1 DFFPOSX1_311 ( .CLK(clk_bF_buf102), .D(_1012_), .Q(datapath_1_RegisterFile_regfile_mem_15__22_) );
DFFPOSX1 DFFPOSX1_312 ( .CLK(clk_bF_buf20), .D(_1013_), .Q(datapath_1_RegisterFile_regfile_mem_15__23_) );
DFFPOSX1 DFFPOSX1_313 ( .CLK(clk_bF_buf64), .D(_1014_), .Q(datapath_1_RegisterFile_regfile_mem_15__24_) );
DFFPOSX1 DFFPOSX1_314 ( .CLK(clk_bF_buf62), .D(_1015_), .Q(datapath_1_RegisterFile_regfile_mem_15__25_) );
DFFPOSX1 DFFPOSX1_315 ( .CLK(clk_bF_buf36), .D(_1016_), .Q(datapath_1_RegisterFile_regfile_mem_15__26_) );
DFFPOSX1 DFFPOSX1_316 ( .CLK(clk_bF_buf72), .D(_1724_), .Q(datapath_1_RegisterFile_regfile_mem_15__27_) );
DFFPOSX1 DFFPOSX1_317 ( .CLK(clk_bF_buf61), .D(_1017_), .Q(datapath_1_RegisterFile_regfile_mem_15__28_) );
DFFPOSX1 DFFPOSX1_318 ( .CLK(clk_bF_buf61), .D(_1018_), .Q(datapath_1_RegisterFile_regfile_mem_15__29_) );
DFFPOSX1 DFFPOSX1_319 ( .CLK(clk_bF_buf37), .D(_1019_), .Q(datapath_1_RegisterFile_regfile_mem_15__30_) );
DFFPOSX1 DFFPOSX1_320 ( .CLK(clk_bF_buf15), .D(_1020_), .Q(datapath_1_RegisterFile_regfile_mem_15__31_) );
DFFPOSX1 DFFPOSX1_321 ( .CLK(clk_bF_buf37), .D(_972_), .Q(datapath_1_RegisterFile_regfile_mem_14__0_) );
DFFPOSX1 DFFPOSX1_322 ( .CLK(clk_bF_buf39), .D(_982_), .Q(datapath_1_RegisterFile_regfile_mem_14__1_) );
DFFPOSX1 DFFPOSX1_323 ( .CLK(clk_bF_buf33), .D(_1710_), .Q(datapath_1_RegisterFile_regfile_mem_14__2_) );
DFFPOSX1 DFFPOSX1_324 ( .CLK(clk_bF_buf39), .D(_994_), .Q(datapath_1_RegisterFile_regfile_mem_14__3_) );
DFFPOSX1 DFFPOSX1_325 ( .CLK(clk_bF_buf111), .D(_995_), .Q(datapath_1_RegisterFile_regfile_mem_14__4_) );
DFFPOSX1 DFFPOSX1_326 ( .CLK(clk_bF_buf45), .D(_996_), .Q(datapath_1_RegisterFile_regfile_mem_14__5_) );
DFFPOSX1 DFFPOSX1_327 ( .CLK(clk_bF_buf107), .D(_997_), .Q(datapath_1_RegisterFile_regfile_mem_14__6_) );
DFFPOSX1 DFFPOSX1_328 ( .CLK(clk_bF_buf61), .D(_998_), .Q(datapath_1_RegisterFile_regfile_mem_14__7_) );
DFFPOSX1 DFFPOSX1_329 ( .CLK(clk_bF_buf92), .D(_999_), .Q(datapath_1_RegisterFile_regfile_mem_14__8_) );
DFFPOSX1 DFFPOSX1_330 ( .CLK(clk_bF_buf45), .D(_1000_), .Q(datapath_1_RegisterFile_regfile_mem_14__9_) );
DFFPOSX1 DFFPOSX1_331 ( .CLK(clk_bF_buf30), .D(_973_), .Q(datapath_1_RegisterFile_regfile_mem_14__10_) );
DFFPOSX1 DFFPOSX1_332 ( .CLK(clk_bF_buf61), .D(_974_), .Q(datapath_1_RegisterFile_regfile_mem_14__11_) );
DFFPOSX1 DFFPOSX1_333 ( .CLK(clk_bF_buf92), .D(_1711_), .Q(datapath_1_RegisterFile_regfile_mem_14__12_) );
DFFPOSX1 DFFPOSX1_334 ( .CLK(clk_bF_buf11), .D(_975_), .Q(datapath_1_RegisterFile_regfile_mem_14__13_) );
DFFPOSX1 DFFPOSX1_335 ( .CLK(clk_bF_buf72), .D(_976_), .Q(datapath_1_RegisterFile_regfile_mem_14__14_) );
DFFPOSX1 DFFPOSX1_336 ( .CLK(clk_bF_buf64), .D(_977_), .Q(datapath_1_RegisterFile_regfile_mem_14__15_) );
DFFPOSX1 DFFPOSX1_337 ( .CLK(clk_bF_buf55), .D(_978_), .Q(datapath_1_RegisterFile_regfile_mem_14__16_) );
DFFPOSX1 DFFPOSX1_338 ( .CLK(clk_bF_buf15), .D(_979_), .Q(datapath_1_RegisterFile_regfile_mem_14__17_) );
DFFPOSX1 DFFPOSX1_339 ( .CLK(clk_bF_buf45), .D(_980_), .Q(datapath_1_RegisterFile_regfile_mem_14__18_) );
DFFPOSX1 DFFPOSX1_340 ( .CLK(clk_bF_buf39), .D(_981_), .Q(datapath_1_RegisterFile_regfile_mem_14__19_) );
DFFPOSX1 DFFPOSX1_341 ( .CLK(clk_bF_buf84), .D(_983_), .Q(datapath_1_RegisterFile_regfile_mem_14__20_) );
DFFPOSX1 DFFPOSX1_342 ( .CLK(clk_bF_buf37), .D(_984_), .Q(datapath_1_RegisterFile_regfile_mem_14__21_) );
DFFPOSX1 DFFPOSX1_343 ( .CLK(clk_bF_buf45), .D(_1712_), .Q(datapath_1_RegisterFile_regfile_mem_14__22_) );
DFFPOSX1 DFFPOSX1_344 ( .CLK(clk_bF_buf20), .D(_985_), .Q(datapath_1_RegisterFile_regfile_mem_14__23_) );
DFFPOSX1 DFFPOSX1_345 ( .CLK(clk_bF_buf64), .D(_986_), .Q(datapath_1_RegisterFile_regfile_mem_14__24_) );
DFFPOSX1 DFFPOSX1_346 ( .CLK(clk_bF_buf99), .D(_987_), .Q(datapath_1_RegisterFile_regfile_mem_14__25_) );
DFFPOSX1 DFFPOSX1_347 ( .CLK(clk_bF_buf36), .D(_988_), .Q(datapath_1_RegisterFile_regfile_mem_14__26_) );
DFFPOSX1 DFFPOSX1_348 ( .CLK(clk_bF_buf72), .D(_989_), .Q(datapath_1_RegisterFile_regfile_mem_14__27_) );
DFFPOSX1 DFFPOSX1_349 ( .CLK(clk_bF_buf35), .D(_990_), .Q(datapath_1_RegisterFile_regfile_mem_14__28_) );
DFFPOSX1 DFFPOSX1_350 ( .CLK(clk_bF_buf61), .D(_991_), .Q(datapath_1_RegisterFile_regfile_mem_14__29_) );
DFFPOSX1 DFFPOSX1_351 ( .CLK(clk_bF_buf37), .D(_992_), .Q(datapath_1_RegisterFile_regfile_mem_14__30_) );
DFFPOSX1 DFFPOSX1_352 ( .CLK(clk_bF_buf72), .D(_993_), .Q(datapath_1_RegisterFile_regfile_mem_14__31_) );
DFFPOSX1 DFFPOSX1_353 ( .CLK(clk_bF_buf53), .D(_945_), .Q(datapath_1_RegisterFile_regfile_mem_13__0_) );
DFFPOSX1 DFFPOSX1_354 ( .CLK(clk_bF_buf107), .D(_955_), .Q(datapath_1_RegisterFile_regfile_mem_13__1_) );
DFFPOSX1 DFFPOSX1_355 ( .CLK(clk_bF_buf92), .D(_965_), .Q(datapath_1_RegisterFile_regfile_mem_13__2_) );
DFFPOSX1 DFFPOSX1_356 ( .CLK(clk_bF_buf62), .D(_966_), .Q(datapath_1_RegisterFile_regfile_mem_13__3_) );
DFFPOSX1 DFFPOSX1_357 ( .CLK(clk_bF_buf37), .D(_967_), .Q(datapath_1_RegisterFile_regfile_mem_13__4_) );
DFFPOSX1 DFFPOSX1_358 ( .CLK(clk_bF_buf46), .D(_968_), .Q(datapath_1_RegisterFile_regfile_mem_13__5_) );
DFFPOSX1 DFFPOSX1_359 ( .CLK(clk_bF_buf107), .D(_969_), .Q(datapath_1_RegisterFile_regfile_mem_13__6_) );
DFFPOSX1 DFFPOSX1_360 ( .CLK(clk_bF_buf32), .D(_1705_), .Q(datapath_1_RegisterFile_regfile_mem_13__7_) );
DFFPOSX1 DFFPOSX1_361 ( .CLK(clk_bF_buf19), .D(_970_), .Q(datapath_1_RegisterFile_regfile_mem_13__8_) );
DFFPOSX1 DFFPOSX1_362 ( .CLK(clk_bF_buf46), .D(_971_), .Q(datapath_1_RegisterFile_regfile_mem_13__9_) );
DFFPOSX1 DFFPOSX1_363 ( .CLK(clk_bF_buf92), .D(_946_), .Q(datapath_1_RegisterFile_regfile_mem_13__10_) );
DFFPOSX1 DFFPOSX1_364 ( .CLK(clk_bF_buf70), .D(_947_), .Q(datapath_1_RegisterFile_regfile_mem_13__11_) );
DFFPOSX1 DFFPOSX1_365 ( .CLK(clk_bF_buf94), .D(_948_), .Q(datapath_1_RegisterFile_regfile_mem_13__12_) );
DFFPOSX1 DFFPOSX1_366 ( .CLK(clk_bF_buf45), .D(_949_), .Q(datapath_1_RegisterFile_regfile_mem_13__13_) );
DFFPOSX1 DFFPOSX1_367 ( .CLK(clk_bF_buf74), .D(_950_), .Q(datapath_1_RegisterFile_regfile_mem_13__14_) );
DFFPOSX1 DFFPOSX1_368 ( .CLK(clk_bF_buf101), .D(_951_), .Q(datapath_1_RegisterFile_regfile_mem_13__15_) );
DFFPOSX1 DFFPOSX1_369 ( .CLK(clk_bF_buf101), .D(_952_), .Q(datapath_1_RegisterFile_regfile_mem_13__16_) );
DFFPOSX1 DFFPOSX1_370 ( .CLK(clk_bF_buf53), .D(_1706_), .Q(datapath_1_RegisterFile_regfile_mem_13__17_) );
DFFPOSX1 DFFPOSX1_371 ( .CLK(clk_bF_buf20), .D(_953_), .Q(datapath_1_RegisterFile_regfile_mem_13__18_) );
DFFPOSX1 DFFPOSX1_372 ( .CLK(clk_bF_buf98), .D(_954_), .Q(datapath_1_RegisterFile_regfile_mem_13__19_) );
DFFPOSX1 DFFPOSX1_373 ( .CLK(clk_bF_buf99), .D(_956_), .Q(datapath_1_RegisterFile_regfile_mem_13__20_) );
DFFPOSX1 DFFPOSX1_374 ( .CLK(clk_bF_buf5), .D(_957_), .Q(datapath_1_RegisterFile_regfile_mem_13__21_) );
DFFPOSX1 DFFPOSX1_375 ( .CLK(clk_bF_buf109), .D(_958_), .Q(datapath_1_RegisterFile_regfile_mem_13__22_) );
DFFPOSX1 DFFPOSX1_376 ( .CLK(clk_bF_buf46), .D(_959_), .Q(datapath_1_RegisterFile_regfile_mem_13__23_) );
DFFPOSX1 DFFPOSX1_377 ( .CLK(clk_bF_buf73), .D(_960_), .Q(datapath_1_RegisterFile_regfile_mem_13__24_) );
DFFPOSX1 DFFPOSX1_378 ( .CLK(clk_bF_buf33), .D(_961_), .Q(datapath_1_RegisterFile_regfile_mem_13__25_) );
DFFPOSX1 DFFPOSX1_379 ( .CLK(clk_bF_buf53), .D(_962_), .Q(datapath_1_RegisterFile_regfile_mem_13__26_) );
DFFPOSX1 DFFPOSX1_380 ( .CLK(clk_bF_buf74), .D(_1707_), .Q(datapath_1_RegisterFile_regfile_mem_13__27_) );
DFFPOSX1 DFFPOSX1_381 ( .CLK(clk_bF_buf73), .D(_963_), .Q(datapath_1_RegisterFile_regfile_mem_13__28_) );
DFFPOSX1 DFFPOSX1_382 ( .CLK(clk_bF_buf35), .D(_964_), .Q(datapath_1_RegisterFile_regfile_mem_13__29_) );
DFFPOSX1 DFFPOSX1_383 ( .CLK(clk_bF_buf111), .D(_1708_), .Q(datapath_1_RegisterFile_regfile_mem_13__30_) );
DFFPOSX1 DFFPOSX1_384 ( .CLK(clk_bF_buf112), .D(_1709_), .Q(datapath_1_RegisterFile_regfile_mem_13__31_) );
DFFPOSX1 DFFPOSX1_385 ( .CLK(clk_bF_buf72), .D(_1563_), .Q(datapath_1_RegisterFile_regfile_mem_7__0_) );
DFFPOSX1 DFFPOSX1_386 ( .CLK(clk_bF_buf81), .D(_1644_), .Q(datapath_1_RegisterFile_regfile_mem_7__1_) );
DFFPOSX1 DFFPOSX1_387 ( .CLK(clk_bF_buf81), .D(_1567_), .Q(datapath_1_RegisterFile_regfile_mem_7__2_) );
DFFPOSX1 DFFPOSX1_388 ( .CLK(clk_bF_buf17), .D(_1568_), .Q(datapath_1_RegisterFile_regfile_mem_7__3_) );
DFFPOSX1 DFFPOSX1_389 ( .CLK(clk_bF_buf82), .D(_1569_), .Q(datapath_1_RegisterFile_regfile_mem_7__4_) );
DFFPOSX1 DFFPOSX1_390 ( .CLK(clk_bF_buf7), .D(_1570_), .Q(datapath_1_RegisterFile_regfile_mem_7__5_) );
DFFPOSX1 DFFPOSX1_391 ( .CLK(clk_bF_buf5), .D(_1571_), .Q(datapath_1_RegisterFile_regfile_mem_7__6_) );
DFFPOSX1 DFFPOSX1_392 ( .CLK(clk_bF_buf32), .D(_1572_), .Q(datapath_1_RegisterFile_regfile_mem_7__7_) );
DFFPOSX1 DFFPOSX1_393 ( .CLK(clk_bF_buf82), .D(_1573_), .Q(datapath_1_RegisterFile_regfile_mem_7__8_) );
DFFPOSX1 DFFPOSX1_394 ( .CLK(clk_bF_buf15), .D(_1574_), .Q(datapath_1_RegisterFile_regfile_mem_7__9_) );
DFFPOSX1 DFFPOSX1_395 ( .CLK(clk_bF_buf51), .D(_1564_), .Q(datapath_1_RegisterFile_regfile_mem_7__10_) );
DFFPOSX1 DFFPOSX1_396 ( .CLK(clk_bF_buf98), .D(_1645_), .Q(datapath_1_RegisterFile_regfile_mem_7__11_) );
DFFPOSX1 DFFPOSX1_397 ( .CLK(clk_bF_buf81), .D(_1565_), .Q(datapath_1_RegisterFile_regfile_mem_7__12_) );
DFFPOSX1 DFFPOSX1_398 ( .CLK(clk_bF_buf87), .D(_1566_), .Q(datapath_1_RegisterFile_regfile_mem_7__13_) );
DFFPOSX1 DFFPOSX1_399 ( .CLK(clk_bF_buf30), .D(_1646_), .Q(datapath_1_RegisterFile_regfile_mem_7__14_) );
DFFPOSX1 DFFPOSX1_400 ( .CLK(clk_bF_buf54), .D(_1647_), .Q(datapath_1_RegisterFile_regfile_mem_7__15_) );
DFFPOSX1 DFFPOSX1_401 ( .CLK(clk_bF_buf32), .D(_1648_), .Q(datapath_1_RegisterFile_regfile_mem_7__16_) );
DFFPOSX1 DFFPOSX1_402 ( .CLK(clk_bF_buf82), .D(_1649_), .Q(datapath_1_RegisterFile_regfile_mem_7__17_) );
DFFPOSX1 DFFPOSX1_403 ( .CLK(clk_bF_buf109), .D(_1650_), .Q(datapath_1_RegisterFile_regfile_mem_7__18_) );
DFFPOSX1 DFFPOSX1_404 ( .CLK(clk_bF_buf98), .D(_1651_), .Q(datapath_1_RegisterFile_regfile_mem_7__19_) );
DFFPOSX1 DFFPOSX1_405 ( .CLK(clk_bF_buf101), .D(_1652_), .Q(datapath_1_RegisterFile_regfile_mem_7__20_) );
DFFPOSX1 DFFPOSX1_406 ( .CLK(clk_bF_buf103), .D(_1653_), .Q(datapath_1_RegisterFile_regfile_mem_7__21_) );
DFFPOSX1 DFFPOSX1_407 ( .CLK(clk_bF_buf87), .D(_1654_), .Q(datapath_1_RegisterFile_regfile_mem_7__22_) );
DFFPOSX1 DFFPOSX1_408 ( .CLK(clk_bF_buf11), .D(_1655_), .Q(datapath_1_RegisterFile_regfile_mem_7__23_) );
DFFPOSX1 DFFPOSX1_409 ( .CLK(clk_bF_buf70), .D(_1656_), .Q(datapath_1_RegisterFile_regfile_mem_7__24_) );
DFFPOSX1 DFFPOSX1_410 ( .CLK(clk_bF_buf51), .D(_1657_), .Q(datapath_1_RegisterFile_regfile_mem_7__25_) );
DFFPOSX1 DFFPOSX1_411 ( .CLK(clk_bF_buf36), .D(_1658_), .Q(datapath_1_RegisterFile_regfile_mem_7__26_) );
DFFPOSX1 DFFPOSX1_412 ( .CLK(clk_bF_buf20), .D(_1659_), .Q(datapath_1_RegisterFile_regfile_mem_7__27_) );
DFFPOSX1 DFFPOSX1_413 ( .CLK(clk_bF_buf32), .D(_1660_), .Q(datapath_1_RegisterFile_regfile_mem_7__28_) );
DFFPOSX1 DFFPOSX1_414 ( .CLK(clk_bF_buf12), .D(_1661_), .Q(datapath_1_RegisterFile_regfile_mem_7__29_) );
DFFPOSX1 DFFPOSX1_415 ( .CLK(clk_bF_buf82), .D(_1662_), .Q(datapath_1_RegisterFile_regfile_mem_7__30_) );
DFFPOSX1 DFFPOSX1_416 ( .CLK(clk_bF_buf7), .D(_1663_), .Q(datapath_1_RegisterFile_regfile_mem_7__31_) );
DFFPOSX1 DFFPOSX1_417 ( .CLK(clk_bF_buf100), .D(_1861_), .Q(datapath_1_RegisterFile_regfile_mem_0__0_) );
DFFPOSX1 DFFPOSX1_418 ( .CLK(clk_bF_buf28), .D(_1862_), .Q(datapath_1_RegisterFile_regfile_mem_0__1_) );
DFFPOSX1 DFFPOSX1_419 ( .CLK(clk_bF_buf93), .D(_1863_), .Q(datapath_1_RegisterFile_regfile_mem_0__2_) );
DFFPOSX1 DFFPOSX1_420 ( .CLK(clk_bF_buf12), .D(_1864_), .Q(datapath_1_RegisterFile_regfile_mem_0__3_) );
DFFPOSX1 DFFPOSX1_421 ( .CLK(clk_bF_buf30), .D(_1865_), .Q(datapath_1_RegisterFile_regfile_mem_0__4_) );
DFFPOSX1 DFFPOSX1_422 ( .CLK(clk_bF_buf36), .D(_1866_), .Q(datapath_1_RegisterFile_regfile_mem_0__5_) );
DFFPOSX1 DFFPOSX1_423 ( .CLK(clk_bF_buf19), .D(_1867_), .Q(datapath_1_RegisterFile_regfile_mem_0__6_) );
DFFPOSX1 DFFPOSX1_424 ( .CLK(clk_bF_buf73), .D(_1868_), .Q(datapath_1_RegisterFile_regfile_mem_0__7_) );
DFFPOSX1 DFFPOSX1_425 ( .CLK(clk_bF_buf82), .D(_1869_), .Q(datapath_1_RegisterFile_regfile_mem_0__8_) );
DFFPOSX1 DFFPOSX1_426 ( .CLK(clk_bF_buf109), .D(_1870_), .Q(datapath_1_RegisterFile_regfile_mem_0__9_) );
DFFPOSX1 DFFPOSX1_427 ( .CLK(clk_bF_buf93), .D(_1871_), .Q(datapath_1_RegisterFile_regfile_mem_0__10_) );
DFFPOSX1 DFFPOSX1_428 ( .CLK(clk_bF_buf12), .D(_1872_), .Q(datapath_1_RegisterFile_regfile_mem_0__11_) );
DFFPOSX1 DFFPOSX1_429 ( .CLK(clk_bF_buf28), .D(_1873_), .Q(datapath_1_RegisterFile_regfile_mem_0__12_) );
DFFPOSX1 DFFPOSX1_430 ( .CLK(clk_bF_buf87), .D(_1874_), .Q(datapath_1_RegisterFile_regfile_mem_0__13_) );
DFFPOSX1 DFFPOSX1_431 ( .CLK(clk_bF_buf11), .D(_1875_), .Q(datapath_1_RegisterFile_regfile_mem_0__14_) );
DFFPOSX1 DFFPOSX1_432 ( .CLK(clk_bF_buf73), .D(_1876_), .Q(datapath_1_RegisterFile_regfile_mem_0__15_) );
DFFPOSX1 DFFPOSX1_433 ( .CLK(clk_bF_buf62), .D(_1877_), .Q(datapath_1_RegisterFile_regfile_mem_0__16_) );
DFFPOSX1 DFFPOSX1_434 ( .CLK(clk_bF_buf106), .D(_1878_), .Q(datapath_1_RegisterFile_regfile_mem_0__17_) );
DFFPOSX1 DFFPOSX1_435 ( .CLK(clk_bF_buf109), .D(_1879_), .Q(datapath_1_RegisterFile_regfile_mem_0__18_) );
DFFPOSX1 DFFPOSX1_436 ( .CLK(clk_bF_buf99), .D(_1880_), .Q(datapath_1_RegisterFile_regfile_mem_0__19_) );
DFFPOSX1 DFFPOSX1_437 ( .CLK(clk_bF_buf12), .D(_1881_), .Q(datapath_1_RegisterFile_regfile_mem_0__20_) );
DFFPOSX1 DFFPOSX1_438 ( .CLK(clk_bF_buf103), .D(_859_), .Q(datapath_1_RegisterFile_regfile_mem_0__21_) );
DFFPOSX1 DFFPOSX1_439 ( .CLK(clk_bF_buf100), .D(_860_), .Q(datapath_1_RegisterFile_regfile_mem_0__22_) );
DFFPOSX1 DFFPOSX1_440 ( .CLK(clk_bF_buf11), .D(_861_), .Q(datapath_1_RegisterFile_regfile_mem_0__23_) );
DFFPOSX1 DFFPOSX1_441 ( .CLK(clk_bF_buf61), .D(_862_), .Q(datapath_1_RegisterFile_regfile_mem_0__24_) );
DFFPOSX1 DFFPOSX1_442 ( .CLK(clk_bF_buf81), .D(_863_), .Q(datapath_1_RegisterFile_regfile_mem_0__25_) );
DFFPOSX1 DFFPOSX1_443 ( .CLK(clk_bF_buf100), .D(_1882_), .Q(datapath_1_RegisterFile_regfile_mem_0__26_) );
DFFPOSX1 DFFPOSX1_444 ( .CLK(clk_bF_buf72), .D(_864_), .Q(datapath_1_RegisterFile_regfile_mem_0__27_) );
DFFPOSX1 DFFPOSX1_445 ( .CLK(clk_bF_buf84), .D(_865_), .Q(datapath_1_RegisterFile_regfile_mem_0__28_) );
DFFPOSX1 DFFPOSX1_446 ( .CLK(clk_bF_buf62), .D(_866_), .Q(datapath_1_RegisterFile_regfile_mem_0__29_) );
DFFPOSX1 DFFPOSX1_447 ( .CLK(clk_bF_buf106), .D(_867_), .Q(datapath_1_RegisterFile_regfile_mem_0__30_) );
DFFPOSX1 DFFPOSX1_448 ( .CLK(clk_bF_buf87), .D(_868_), .Q(datapath_1_RegisterFile_regfile_mem_0__31_) );
DFFPOSX1 DFFPOSX1_449 ( .CLK(clk_bF_buf100), .D(_1128_), .Q(datapath_1_RegisterFile_regfile_mem_1__0_) );
DFFPOSX1 DFFPOSX1_450 ( .CLK(clk_bF_buf28), .D(_1618_), .Q(datapath_1_RegisterFile_regfile_mem_1__1_) );
DFFPOSX1 DFFPOSX1_451 ( .CLK(clk_bF_buf33), .D(_1141_), .Q(datapath_1_RegisterFile_regfile_mem_1__2_) );
DFFPOSX1 DFFPOSX1_452 ( .CLK(clk_bF_buf12), .D(_1143_), .Q(datapath_1_RegisterFile_regfile_mem_1__3_) );
DFFPOSX1 DFFPOSX1_453 ( .CLK(clk_bF_buf82), .D(_1144_), .Q(datapath_1_RegisterFile_regfile_mem_1__4_) );
DFFPOSX1 DFFPOSX1_454 ( .CLK(clk_bF_buf11), .D(_1145_), .Q(datapath_1_RegisterFile_regfile_mem_1__5_) );
DFFPOSX1 DFFPOSX1_455 ( .CLK(clk_bF_buf19), .D(_1619_), .Q(datapath_1_RegisterFile_regfile_mem_1__6_) );
DFFPOSX1 DFFPOSX1_456 ( .CLK(clk_bF_buf73), .D(_1146_), .Q(datapath_1_RegisterFile_regfile_mem_1__7_) );
DFFPOSX1 DFFPOSX1_457 ( .CLK(clk_bF_buf82), .D(_1147_), .Q(datapath_1_RegisterFile_regfile_mem_1__8_) );
DFFPOSX1 DFFPOSX1_458 ( .CLK(clk_bF_buf20), .D(_1148_), .Q(datapath_1_RegisterFile_regfile_mem_1__9_) );
DFFPOSX1 DFFPOSX1_459 ( .CLK(clk_bF_buf103), .D(_1129_), .Q(datapath_1_RegisterFile_regfile_mem_1__10_) );
DFFPOSX1 DFFPOSX1_460 ( .CLK(clk_bF_buf17), .D(_1620_), .Q(datapath_1_RegisterFile_regfile_mem_1__11_) );
DFFPOSX1 DFFPOSX1_461 ( .CLK(clk_bF_buf33), .D(_1130_), .Q(datapath_1_RegisterFile_regfile_mem_1__12_) );
DFFPOSX1 DFFPOSX1_462 ( .CLK(clk_bF_buf109), .D(_1131_), .Q(datapath_1_RegisterFile_regfile_mem_1__13_) );
DFFPOSX1 DFFPOSX1_463 ( .CLK(clk_bF_buf72), .D(_1132_), .Q(datapath_1_RegisterFile_regfile_mem_1__14_) );
DFFPOSX1 DFFPOSX1_464 ( .CLK(clk_bF_buf61), .D(_1133_), .Q(datapath_1_RegisterFile_regfile_mem_1__15_) );
DFFPOSX1 DFFPOSX1_465 ( .CLK(clk_bF_buf39), .D(_1621_), .Q(datapath_1_RegisterFile_regfile_mem_1__16_) );
DFFPOSX1 DFFPOSX1_466 ( .CLK(clk_bF_buf23), .D(_1134_), .Q(datapath_1_RegisterFile_regfile_mem_1__17_) );
DFFPOSX1 DFFPOSX1_467 ( .CLK(clk_bF_buf109), .D(_1622_), .Q(datapath_1_RegisterFile_regfile_mem_1__18_) );
DFFPOSX1 DFFPOSX1_468 ( .CLK(clk_bF_buf84), .D(_1623_), .Q(datapath_1_RegisterFile_regfile_mem_1__19_) );
DFFPOSX1 DFFPOSX1_469 ( .CLK(clk_bF_buf84), .D(_1624_), .Q(datapath_1_RegisterFile_regfile_mem_1__20_) );
DFFPOSX1 DFFPOSX1_470 ( .CLK(clk_bF_buf103), .D(_1625_), .Q(datapath_1_RegisterFile_regfile_mem_1__21_) );
DFFPOSX1 DFFPOSX1_471 ( .CLK(clk_bF_buf100), .D(_1626_), .Q(datapath_1_RegisterFile_regfile_mem_1__22_) );
DFFPOSX1 DFFPOSX1_472 ( .CLK(clk_bF_buf112), .D(_1135_), .Q(datapath_1_RegisterFile_regfile_mem_1__23_) );
DFFPOSX1 DFFPOSX1_473 ( .CLK(clk_bF_buf73), .D(_1136_), .Q(datapath_1_RegisterFile_regfile_mem_1__24_) );
DFFPOSX1 DFFPOSX1_474 ( .CLK(clk_bF_buf17), .D(_1137_), .Q(datapath_1_RegisterFile_regfile_mem_1__25_) );
DFFPOSX1 DFFPOSX1_475 ( .CLK(clk_bF_buf36), .D(_1627_), .Q(datapath_1_RegisterFile_regfile_mem_1__26_) );
DFFPOSX1 DFFPOSX1_476 ( .CLK(clk_bF_buf11), .D(_1138_), .Q(datapath_1_RegisterFile_regfile_mem_1__27_) );
DFFPOSX1 DFFPOSX1_477 ( .CLK(clk_bF_buf99), .D(_1139_), .Q(datapath_1_RegisterFile_regfile_mem_1__28_) );
DFFPOSX1 DFFPOSX1_478 ( .CLK(clk_bF_buf39), .D(_1140_), .Q(datapath_1_RegisterFile_regfile_mem_1__29_) );
DFFPOSX1 DFFPOSX1_479 ( .CLK(clk_bF_buf106), .D(_1142_), .Q(datapath_1_RegisterFile_regfile_mem_1__30_) );
DFFPOSX1 DFFPOSX1_480 ( .CLK(clk_bF_buf86), .D(_1628_), .Q(datapath_1_RegisterFile_regfile_mem_1__31_) );
DFFPOSX1 DFFPOSX1_481 ( .CLK(clk_bF_buf53), .D(_1534_), .Q(datapath_1_RegisterFile_regfile_mem_6__0_) );
DFFPOSX1 DFFPOSX1_482 ( .CLK(clk_bF_buf81), .D(_1544_), .Q(datapath_1_RegisterFile_regfile_mem_6__1_) );
DFFPOSX1 DFFPOSX1_483 ( .CLK(clk_bF_buf17), .D(_1554_), .Q(datapath_1_RegisterFile_regfile_mem_6__2_) );
DFFPOSX1 DFFPOSX1_484 ( .CLK(clk_bF_buf17), .D(_1557_), .Q(datapath_1_RegisterFile_regfile_mem_6__3_) );
DFFPOSX1 DFFPOSX1_485 ( .CLK(clk_bF_buf111), .D(_1558_), .Q(datapath_1_RegisterFile_regfile_mem_6__4_) );
DFFPOSX1 DFFPOSX1_486 ( .CLK(clk_bF_buf109), .D(_1559_), .Q(datapath_1_RegisterFile_regfile_mem_6__5_) );
DFFPOSX1 DFFPOSX1_487 ( .CLK(clk_bF_buf28), .D(_1560_), .Q(datapath_1_RegisterFile_regfile_mem_6__6_) );
DFFPOSX1 DFFPOSX1_488 ( .CLK(clk_bF_buf32), .D(_1561_), .Q(datapath_1_RegisterFile_regfile_mem_6__7_) );
DFFPOSX1 DFFPOSX1_489 ( .CLK(clk_bF_buf81), .D(_1641_), .Q(datapath_1_RegisterFile_regfile_mem_6__8_) );
DFFPOSX1 DFFPOSX1_490 ( .CLK(clk_bF_buf36), .D(_1562_), .Q(datapath_1_RegisterFile_regfile_mem_6__9_) );
DFFPOSX1 DFFPOSX1_491 ( .CLK(clk_bF_buf103), .D(_1535_), .Q(datapath_1_RegisterFile_regfile_mem_6__10_) );
DFFPOSX1 DFFPOSX1_492 ( .CLK(clk_bF_buf98), .D(_1536_), .Q(datapath_1_RegisterFile_regfile_mem_6__11_) );
DFFPOSX1 DFFPOSX1_493 ( .CLK(clk_bF_buf81), .D(_1537_), .Q(datapath_1_RegisterFile_regfile_mem_6__12_) );
DFFPOSX1 DFFPOSX1_494 ( .CLK(clk_bF_buf7), .D(_1538_), .Q(datapath_1_RegisterFile_regfile_mem_6__13_) );
DFFPOSX1 DFFPOSX1_495 ( .CLK(clk_bF_buf5), .D(_1539_), .Q(datapath_1_RegisterFile_regfile_mem_6__14_) );
DFFPOSX1 DFFPOSX1_496 ( .CLK(clk_bF_buf54), .D(_1540_), .Q(datapath_1_RegisterFile_regfile_mem_6__15_) );
DFFPOSX1 DFFPOSX1_497 ( .CLK(clk_bF_buf110), .D(_1541_), .Q(datapath_1_RegisterFile_regfile_mem_6__16_) );
DFFPOSX1 DFFPOSX1_498 ( .CLK(clk_bF_buf111), .D(_1542_), .Q(datapath_1_RegisterFile_regfile_mem_6__17_) );
DFFPOSX1 DFFPOSX1_499 ( .CLK(clk_bF_buf7), .D(_1642_), .Q(datapath_1_RegisterFile_regfile_mem_6__18_) );
DFFPOSX1 DFFPOSX1_500 ( .CLK(clk_bF_buf98), .D(_1543_), .Q(datapath_1_RegisterFile_regfile_mem_6__19_) );
DFFPOSX1 DFFPOSX1_501 ( .CLK(clk_bF_buf12), .D(_1545_), .Q(datapath_1_RegisterFile_regfile_mem_6__20_) );
DFFPOSX1 DFFPOSX1_502 ( .CLK(clk_bF_buf82), .D(_1546_), .Q(datapath_1_RegisterFile_regfile_mem_6__21_) );
DFFPOSX1 DFFPOSX1_503 ( .CLK(clk_bF_buf87), .D(_1547_), .Q(datapath_1_RegisterFile_regfile_mem_6__22_) );
DFFPOSX1 DFFPOSX1_504 ( .CLK(clk_bF_buf46), .D(_1548_), .Q(datapath_1_RegisterFile_regfile_mem_6__23_) );
DFFPOSX1 DFFPOSX1_505 ( .CLK(clk_bF_buf54), .D(_1549_), .Q(datapath_1_RegisterFile_regfile_mem_6__24_) );
DFFPOSX1 DFFPOSX1_506 ( .CLK(clk_bF_buf81), .D(_1550_), .Q(datapath_1_RegisterFile_regfile_mem_6__25_) );
DFFPOSX1 DFFPOSX1_507 ( .CLK(clk_bF_buf53), .D(_1551_), .Q(datapath_1_RegisterFile_regfile_mem_6__26_) );
DFFPOSX1 DFFPOSX1_508 ( .CLK(clk_bF_buf16), .D(_1552_), .Q(datapath_1_RegisterFile_regfile_mem_6__27_) );
DFFPOSX1 DFFPOSX1_509 ( .CLK(clk_bF_buf32), .D(_1643_), .Q(datapath_1_RegisterFile_regfile_mem_6__28_) );
DFFPOSX1 DFFPOSX1_510 ( .CLK(clk_bF_buf110), .D(_1553_), .Q(datapath_1_RegisterFile_regfile_mem_6__29_) );
DFFPOSX1 DFFPOSX1_511 ( .CLK(clk_bF_buf111), .D(_1555_), .Q(datapath_1_RegisterFile_regfile_mem_6__30_) );
DFFPOSX1 DFFPOSX1_512 ( .CLK(clk_bF_buf36), .D(_1556_), .Q(datapath_1_RegisterFile_regfile_mem_6__31_) );
DFFPOSX1 DFFPOSX1_513 ( .CLK(clk_bF_buf74), .D(_891_), .Q(datapath_1_RegisterFile_regfile_mem_11__0_) );
DFFPOSX1 DFFPOSX1_514 ( .CLK(clk_bF_buf39), .D(_901_), .Q(datapath_1_RegisterFile_regfile_mem_11__1_) );
DFFPOSX1 DFFPOSX1_515 ( .CLK(clk_bF_buf93), .D(_911_), .Q(datapath_1_RegisterFile_regfile_mem_11__2_) );
DFFPOSX1 DFFPOSX1_516 ( .CLK(clk_bF_buf39), .D(_914_), .Q(datapath_1_RegisterFile_regfile_mem_11__3_) );
DFFPOSX1 DFFPOSX1_517 ( .CLK(clk_bF_buf82), .D(_915_), .Q(datapath_1_RegisterFile_regfile_mem_11__4_) );
DFFPOSX1 DFFPOSX1_518 ( .CLK(clk_bF_buf16), .D(_916_), .Q(datapath_1_RegisterFile_regfile_mem_11__5_) );
DFFPOSX1 DFFPOSX1_519 ( .CLK(clk_bF_buf5), .D(_917_), .Q(datapath_1_RegisterFile_regfile_mem_11__6_) );
DFFPOSX1 DFFPOSX1_520 ( .CLK(clk_bF_buf64), .D(_1695_), .Q(datapath_1_RegisterFile_regfile_mem_11__7_) );
DFFPOSX1 DFFPOSX1_521 ( .CLK(clk_bF_buf94), .D(_918_), .Q(datapath_1_RegisterFile_regfile_mem_11__8_) );
DFFPOSX1 DFFPOSX1_522 ( .CLK(clk_bF_buf16), .D(_919_), .Q(datapath_1_RegisterFile_regfile_mem_11__9_) );
DFFPOSX1 DFFPOSX1_523 ( .CLK(clk_bF_buf94), .D(_892_), .Q(datapath_1_RegisterFile_regfile_mem_11__10_) );
DFFPOSX1 DFFPOSX1_524 ( .CLK(clk_bF_buf73), .D(_893_), .Q(datapath_1_RegisterFile_regfile_mem_11__11_) );
DFFPOSX1 DFFPOSX1_525 ( .CLK(clk_bF_buf107), .D(_894_), .Q(datapath_1_RegisterFile_regfile_mem_11__12_) );
DFFPOSX1 DFFPOSX1_526 ( .CLK(clk_bF_buf16), .D(_895_), .Q(datapath_1_RegisterFile_regfile_mem_11__13_) );
DFFPOSX1 DFFPOSX1_527 ( .CLK(clk_bF_buf15), .D(_896_), .Q(datapath_1_RegisterFile_regfile_mem_11__14_) );
DFFPOSX1 DFFPOSX1_528 ( .CLK(clk_bF_buf64), .D(_897_), .Q(datapath_1_RegisterFile_regfile_mem_11__15_) );
DFFPOSX1 DFFPOSX1_529 ( .CLK(clk_bF_buf64), .D(_898_), .Q(datapath_1_RegisterFile_regfile_mem_11__16_) );
DFFPOSX1 DFFPOSX1_530 ( .CLK(clk_bF_buf111), .D(_1696_), .Q(datapath_1_RegisterFile_regfile_mem_11__17_) );
DFFPOSX1 DFFPOSX1_531 ( .CLK(clk_bF_buf102), .D(_899_), .Q(datapath_1_RegisterFile_regfile_mem_11__18_) );
DFFPOSX1 DFFPOSX1_532 ( .CLK(clk_bF_buf84), .D(_900_), .Q(datapath_1_RegisterFile_regfile_mem_11__19_) );
DFFPOSX1 DFFPOSX1_533 ( .CLK(clk_bF_buf84), .D(_902_), .Q(datapath_1_RegisterFile_regfile_mem_11__20_) );
DFFPOSX1 DFFPOSX1_534 ( .CLK(clk_bF_buf5), .D(_903_), .Q(datapath_1_RegisterFile_regfile_mem_11__21_) );
DFFPOSX1 DFFPOSX1_535 ( .CLK(clk_bF_buf102), .D(_904_), .Q(datapath_1_RegisterFile_regfile_mem_11__22_) );
DFFPOSX1 DFFPOSX1_536 ( .CLK(clk_bF_buf46), .D(_905_), .Q(datapath_1_RegisterFile_regfile_mem_11__23_) );
DFFPOSX1 DFFPOSX1_537 ( .CLK(clk_bF_buf55), .D(_906_), .Q(datapath_1_RegisterFile_regfile_mem_11__24_) );
DFFPOSX1 DFFPOSX1_538 ( .CLK(clk_bF_buf101), .D(_907_), .Q(datapath_1_RegisterFile_regfile_mem_11__25_) );
DFFPOSX1 DFFPOSX1_539 ( .CLK(clk_bF_buf112), .D(_908_), .Q(datapath_1_RegisterFile_regfile_mem_11__26_) );
DFFPOSX1 DFFPOSX1_540 ( .CLK(clk_bF_buf74), .D(_1697_), .Q(datapath_1_RegisterFile_regfile_mem_11__27_) );
DFFPOSX1 DFFPOSX1_541 ( .CLK(clk_bF_buf35), .D(_909_), .Q(datapath_1_RegisterFile_regfile_mem_11__28_) );
DFFPOSX1 DFFPOSX1_542 ( .CLK(clk_bF_buf99), .D(_910_), .Q(datapath_1_RegisterFile_regfile_mem_11__29_) );
DFFPOSX1 DFFPOSX1_543 ( .CLK(clk_bF_buf37), .D(_912_), .Q(datapath_1_RegisterFile_regfile_mem_11__30_) );
DFFPOSX1 DFFPOSX1_544 ( .CLK(clk_bF_buf74), .D(_913_), .Q(datapath_1_RegisterFile_regfile_mem_11__31_) );
DFFPOSX1 DFFPOSX1_545 ( .CLK(clk_bF_buf77), .D(_1314_), .Q(datapath_1_RegisterFile_regfile_mem_28__0_) );
DFFPOSX1 DFFPOSX1_546 ( .CLK(clk_bF_buf21), .D(_1324_), .Q(datapath_1_RegisterFile_regfile_mem_28__1_) );
DFFPOSX1 DFFPOSX1_547 ( .CLK(clk_bF_buf40), .D(_1331_), .Q(datapath_1_RegisterFile_regfile_mem_28__2_) );
DFFPOSX1 DFFPOSX1_548 ( .CLK(clk_bF_buf63), .D(_1332_), .Q(datapath_1_RegisterFile_regfile_mem_28__3_) );
DFFPOSX1 DFFPOSX1_549 ( .CLK(clk_bF_buf96), .D(_1837_), .Q(datapath_1_RegisterFile_regfile_mem_28__4_) );
DFFPOSX1 DFFPOSX1_550 ( .CLK(clk_bF_buf29), .D(_1333_), .Q(datapath_1_RegisterFile_regfile_mem_28__5_) );
DFFPOSX1 DFFPOSX1_551 ( .CLK(clk_bF_buf76), .D(_1334_), .Q(datapath_1_RegisterFile_regfile_mem_28__6_) );
DFFPOSX1 DFFPOSX1_552 ( .CLK(clk_bF_buf98), .D(_1335_), .Q(datapath_1_RegisterFile_regfile_mem_28__7_) );
DFFPOSX1 DFFPOSX1_553 ( .CLK(clk_bF_buf26), .D(_1336_), .Q(datapath_1_RegisterFile_regfile_mem_28__8_) );
DFFPOSX1 DFFPOSX1_554 ( .CLK(clk_bF_buf79), .D(_1337_), .Q(datapath_1_RegisterFile_regfile_mem_28__9_) );
DFFPOSX1 DFFPOSX1_555 ( .CLK(clk_bF_buf13), .D(_1315_), .Q(datapath_1_RegisterFile_regfile_mem_28__10_) );
DFFPOSX1 DFFPOSX1_556 ( .CLK(clk_bF_buf89), .D(_1316_), .Q(datapath_1_RegisterFile_regfile_mem_28__11_) );
DFFPOSX1 DFFPOSX1_557 ( .CLK(clk_bF_buf41), .D(_1317_), .Q(datapath_1_RegisterFile_regfile_mem_28__12_) );
DFFPOSX1 DFFPOSX1_558 ( .CLK(clk_bF_buf13), .D(_1318_), .Q(datapath_1_RegisterFile_regfile_mem_28__13_) );
DFFPOSX1 DFFPOSX1_559 ( .CLK(clk_bF_buf48), .D(_1838_), .Q(datapath_1_RegisterFile_regfile_mem_28__14_) );
DFFPOSX1 DFFPOSX1_560 ( .CLK(clk_bF_buf42), .D(_1319_), .Q(datapath_1_RegisterFile_regfile_mem_28__15_) );
DFFPOSX1 DFFPOSX1_561 ( .CLK(clk_bF_buf31), .D(_1320_), .Q(datapath_1_RegisterFile_regfile_mem_28__16_) );
DFFPOSX1 DFFPOSX1_562 ( .CLK(clk_bF_buf77), .D(_1321_), .Q(datapath_1_RegisterFile_regfile_mem_28__17_) );
DFFPOSX1 DFFPOSX1_563 ( .CLK(clk_bF_buf86), .D(_1322_), .Q(datapath_1_RegisterFile_regfile_mem_28__18_) );
DFFPOSX1 DFFPOSX1_564 ( .CLK(clk_bF_buf40), .D(_1323_), .Q(datapath_1_RegisterFile_regfile_mem_28__19_) );
DFFPOSX1 DFFPOSX1_565 ( .CLK(clk_bF_buf49), .D(_1325_), .Q(datapath_1_RegisterFile_regfile_mem_28__20_) );
DFFPOSX1 DFFPOSX1_566 ( .CLK(clk_bF_buf1), .D(_1326_), .Q(datapath_1_RegisterFile_regfile_mem_28__21_) );
DFFPOSX1 DFFPOSX1_567 ( .CLK(clk_bF_buf29), .D(_1327_), .Q(datapath_1_RegisterFile_regfile_mem_28__22_) );
DFFPOSX1 DFFPOSX1_568 ( .CLK(clk_bF_buf113), .D(_1328_), .Q(datapath_1_RegisterFile_regfile_mem_28__23_) );
DFFPOSX1 DFFPOSX1_569 ( .CLK(clk_bF_buf6), .D(_1839_), .Q(datapath_1_RegisterFile_regfile_mem_28__24_) );
DFFPOSX1 DFFPOSX1_570 ( .CLK(clk_bF_buf65), .D(_1329_), .Q(datapath_1_RegisterFile_regfile_mem_28__25_) );
DFFPOSX1 DFFPOSX1_571 ( .CLK(clk_bF_buf13), .D(_1330_), .Q(datapath_1_RegisterFile_regfile_mem_28__26_) );
DFFPOSX1 DFFPOSX1_572 ( .CLK(clk_bF_buf86), .D(_1840_), .Q(datapath_1_RegisterFile_regfile_mem_28__27_) );
DFFPOSX1 DFFPOSX1_573 ( .CLK(clk_bF_buf63), .D(_1841_), .Q(datapath_1_RegisterFile_regfile_mem_28__28_) );
DFFPOSX1 DFFPOSX1_574 ( .CLK(clk_bF_buf31), .D(_1842_), .Q(datapath_1_RegisterFile_regfile_mem_28__29_) );
DFFPOSX1 DFFPOSX1_575 ( .CLK(clk_bF_buf60), .D(_1843_), .Q(datapath_1_RegisterFile_regfile_mem_28__30_) );
DFFPOSX1 DFFPOSX1_576 ( .CLK(clk_bF_buf48), .D(_1844_), .Q(datapath_1_RegisterFile_regfile_mem_28__31_) );
DFFPOSX1 DFFPOSX1_577 ( .CLK(clk_bF_buf23), .D(_1447_), .Q(datapath_1_RegisterFile_regfile_mem_3__0_) );
DFFPOSX1 DFFPOSX1_578 ( .CLK(clk_bF_buf107), .D(_1457_), .Q(datapath_1_RegisterFile_regfile_mem_3__1_) );
DFFPOSX1 DFFPOSX1_579 ( .CLK(clk_bF_buf93), .D(_1467_), .Q(datapath_1_RegisterFile_regfile_mem_3__2_) );
DFFPOSX1 DFFPOSX1_580 ( .CLK(clk_bF_buf110), .D(_1470_), .Q(datapath_1_RegisterFile_regfile_mem_3__3_) );
DFFPOSX1 DFFPOSX1_581 ( .CLK(clk_bF_buf19), .D(_1471_), .Q(datapath_1_RegisterFile_regfile_mem_3__4_) );
DFFPOSX1 DFFPOSX1_582 ( .CLK(clk_bF_buf45), .D(_1472_), .Q(datapath_1_RegisterFile_regfile_mem_3__5_) );
DFFPOSX1 DFFPOSX1_583 ( .CLK(clk_bF_buf28), .D(_1473_), .Q(datapath_1_RegisterFile_regfile_mem_3__6_) );
DFFPOSX1 DFFPOSX1_584 ( .CLK(clk_bF_buf61), .D(_1474_), .Q(datapath_1_RegisterFile_regfile_mem_3__7_) );
DFFPOSX1 DFFPOSX1_585 ( .CLK(clk_bF_buf103), .D(_1475_), .Q(datapath_1_RegisterFile_regfile_mem_3__8_) );
DFFPOSX1 DFFPOSX1_586 ( .CLK(clk_bF_buf23), .D(_1632_), .Q(datapath_1_RegisterFile_regfile_mem_3__9_) );
DFFPOSX1 DFFPOSX1_587 ( .CLK(clk_bF_buf103), .D(_1448_), .Q(datapath_1_RegisterFile_regfile_mem_3__10_) );
DFFPOSX1 DFFPOSX1_588 ( .CLK(clk_bF_buf110), .D(_1449_), .Q(datapath_1_RegisterFile_regfile_mem_3__11_) );
DFFPOSX1 DFFPOSX1_589 ( .CLK(clk_bF_buf33), .D(_1450_), .Q(datapath_1_RegisterFile_regfile_mem_3__12_) );
DFFPOSX1 DFFPOSX1_590 ( .CLK(clk_bF_buf109), .D(_1451_), .Q(datapath_1_RegisterFile_regfile_mem_3__13_) );
DFFPOSX1 DFFPOSX1_591 ( .CLK(clk_bF_buf7), .D(_1452_), .Q(datapath_1_RegisterFile_regfile_mem_3__14_) );
DFFPOSX1 DFFPOSX1_592 ( .CLK(clk_bF_buf73), .D(_1453_), .Q(datapath_1_RegisterFile_regfile_mem_3__15_) );
DFFPOSX1 DFFPOSX1_593 ( .CLK(clk_bF_buf84), .D(_1454_), .Q(datapath_1_RegisterFile_regfile_mem_3__16_) );
DFFPOSX1 DFFPOSX1_594 ( .CLK(clk_bF_buf23), .D(_1455_), .Q(datapath_1_RegisterFile_regfile_mem_3__17_) );
DFFPOSX1 DFFPOSX1_595 ( .CLK(clk_bF_buf46), .D(_1456_), .Q(datapath_1_RegisterFile_regfile_mem_3__18_) );
DFFPOSX1 DFFPOSX1_596 ( .CLK(clk_bF_buf84), .D(_1633_), .Q(datapath_1_RegisterFile_regfile_mem_3__19_) );
DFFPOSX1 DFFPOSX1_597 ( .CLK(clk_bF_buf99), .D(_1458_), .Q(datapath_1_RegisterFile_regfile_mem_3__20_) );
DFFPOSX1 DFFPOSX1_598 ( .CLK(clk_bF_buf103), .D(_1459_), .Q(datapath_1_RegisterFile_regfile_mem_3__21_) );
DFFPOSX1 DFFPOSX1_599 ( .CLK(clk_bF_buf23), .D(_1460_), .Q(datapath_1_RegisterFile_regfile_mem_3__22_) );
DFFPOSX1 DFFPOSX1_600 ( .CLK(clk_bF_buf11), .D(_1461_), .Q(datapath_1_RegisterFile_regfile_mem_3__23_) );
DFFPOSX1 DFFPOSX1_601 ( .CLK(clk_bF_buf35), .D(_1462_), .Q(datapath_1_RegisterFile_regfile_mem_3__24_) );
DFFPOSX1 DFFPOSX1_602 ( .CLK(clk_bF_buf17), .D(_1463_), .Q(datapath_1_RegisterFile_regfile_mem_3__25_) );
DFFPOSX1 DFFPOSX1_603 ( .CLK(clk_bF_buf36), .D(_1464_), .Q(datapath_1_RegisterFile_regfile_mem_3__26_) );
DFFPOSX1 DFFPOSX1_604 ( .CLK(clk_bF_buf7), .D(_1465_), .Q(datapath_1_RegisterFile_regfile_mem_3__27_) );
DFFPOSX1 DFFPOSX1_605 ( .CLK(clk_bF_buf99), .D(_1466_), .Q(datapath_1_RegisterFile_regfile_mem_3__28_) );
DFFPOSX1 DFFPOSX1_606 ( .CLK(clk_bF_buf110), .D(_1634_), .Q(datapath_1_RegisterFile_regfile_mem_3__29_) );
DFFPOSX1 DFFPOSX1_607 ( .CLK(clk_bF_buf106), .D(_1468_), .Q(datapath_1_RegisterFile_regfile_mem_3__30_) );
DFFPOSX1 DFFPOSX1_608 ( .CLK(clk_bF_buf11), .D(_1469_), .Q(datapath_1_RegisterFile_regfile_mem_3__31_) );
DFFPOSX1 DFFPOSX1_609 ( .CLK(clk_bF_buf23), .D(_1367_), .Q(datapath_1_RegisterFile_regfile_mem_2__0_) );
DFFPOSX1 DFFPOSX1_610 ( .CLK(clk_bF_buf103), .D(_1377_), .Q(datapath_1_RegisterFile_regfile_mem_2__1_) );
DFFPOSX1 DFFPOSX1_611 ( .CLK(clk_bF_buf93), .D(_1387_), .Q(datapath_1_RegisterFile_regfile_mem_2__2_) );
DFFPOSX1 DFFPOSX1_612 ( .CLK(clk_bF_buf17), .D(_1390_), .Q(datapath_1_RegisterFile_regfile_mem_2__3_) );
DFFPOSX1 DFFPOSX1_613 ( .CLK(clk_bF_buf106), .D(_1391_), .Q(datapath_1_RegisterFile_regfile_mem_2__4_) );
DFFPOSX1 DFFPOSX1_614 ( .CLK(clk_bF_buf45), .D(_1392_), .Q(datapath_1_RegisterFile_regfile_mem_2__5_) );
DFFPOSX1 DFFPOSX1_615 ( .CLK(clk_bF_buf5), .D(_1629_), .Q(datapath_1_RegisterFile_regfile_mem_2__6_) );
DFFPOSX1 DFFPOSX1_616 ( .CLK(clk_bF_buf73), .D(_1393_), .Q(datapath_1_RegisterFile_regfile_mem_2__7_) );
DFFPOSX1 DFFPOSX1_617 ( .CLK(clk_bF_buf19), .D(_1394_), .Q(datapath_1_RegisterFile_regfile_mem_2__8_) );
DFFPOSX1 DFFPOSX1_618 ( .CLK(clk_bF_buf74), .D(_1395_), .Q(datapath_1_RegisterFile_regfile_mem_2__9_) );
DFFPOSX1 DFFPOSX1_619 ( .CLK(clk_bF_buf51), .D(_1368_), .Q(datapath_1_RegisterFile_regfile_mem_2__10_) );
DFFPOSX1 DFFPOSX1_620 ( .CLK(clk_bF_buf110), .D(_1369_), .Q(datapath_1_RegisterFile_regfile_mem_2__11_) );
DFFPOSX1 DFFPOSX1_621 ( .CLK(clk_bF_buf107), .D(_1370_), .Q(datapath_1_RegisterFile_regfile_mem_2__12_) );
DFFPOSX1 DFFPOSX1_622 ( .CLK(clk_bF_buf109), .D(_1371_), .Q(datapath_1_RegisterFile_regfile_mem_2__13_) );
DFFPOSX1 DFFPOSX1_623 ( .CLK(clk_bF_buf74), .D(_1372_), .Q(datapath_1_RegisterFile_regfile_mem_2__14_) );
DFFPOSX1 DFFPOSX1_624 ( .CLK(clk_bF_buf73), .D(_1373_), .Q(datapath_1_RegisterFile_regfile_mem_2__15_) );
DFFPOSX1 DFFPOSX1_625 ( .CLK(clk_bF_buf39), .D(_1630_), .Q(datapath_1_RegisterFile_regfile_mem_2__16_) );
DFFPOSX1 DFFPOSX1_626 ( .CLK(clk_bF_buf53), .D(_1374_), .Q(datapath_1_RegisterFile_regfile_mem_2__17_) );
DFFPOSX1 DFFPOSX1_627 ( .CLK(clk_bF_buf87), .D(_1375_), .Q(datapath_1_RegisterFile_regfile_mem_2__18_) );
DFFPOSX1 DFFPOSX1_628 ( .CLK(clk_bF_buf99), .D(_1376_), .Q(datapath_1_RegisterFile_regfile_mem_2__19_) );
DFFPOSX1 DFFPOSX1_629 ( .CLK(clk_bF_buf84), .D(_1378_), .Q(datapath_1_RegisterFile_regfile_mem_2__20_) );
DFFPOSX1 DFFPOSX1_630 ( .CLK(clk_bF_buf28), .D(_1379_), .Q(datapath_1_RegisterFile_regfile_mem_2__21_) );
DFFPOSX1 DFFPOSX1_631 ( .CLK(clk_bF_buf87), .D(_1380_), .Q(datapath_1_RegisterFile_regfile_mem_2__22_) );
DFFPOSX1 DFFPOSX1_632 ( .CLK(clk_bF_buf112), .D(_1381_), .Q(datapath_1_RegisterFile_regfile_mem_2__23_) );
DFFPOSX1 DFFPOSX1_633 ( .CLK(clk_bF_buf35), .D(_1382_), .Q(datapath_1_RegisterFile_regfile_mem_2__24_) );
DFFPOSX1 DFFPOSX1_634 ( .CLK(clk_bF_buf28), .D(_1383_), .Q(datapath_1_RegisterFile_regfile_mem_2__25_) );
DFFPOSX1 DFFPOSX1_635 ( .CLK(clk_bF_buf36), .D(_1631_), .Q(datapath_1_RegisterFile_regfile_mem_2__26_) );
DFFPOSX1 DFFPOSX1_636 ( .CLK(clk_bF_buf74), .D(_1384_), .Q(datapath_1_RegisterFile_regfile_mem_2__27_) );
DFFPOSX1 DFFPOSX1_637 ( .CLK(clk_bF_buf35), .D(_1385_), .Q(datapath_1_RegisterFile_regfile_mem_2__28_) );
DFFPOSX1 DFFPOSX1_638 ( .CLK(clk_bF_buf110), .D(_1386_), .Q(datapath_1_RegisterFile_regfile_mem_2__29_) );
DFFPOSX1 DFFPOSX1_639 ( .CLK(clk_bF_buf106), .D(_1388_), .Q(datapath_1_RegisterFile_regfile_mem_2__30_) );
DFFPOSX1 DFFPOSX1_640 ( .CLK(clk_bF_buf100), .D(_1389_), .Q(datapath_1_RegisterFile_regfile_mem_2__31_) );
DFFPOSX1 DFFPOSX1_641 ( .CLK(clk_bF_buf23), .D(_1476_), .Q(datapath_1_RegisterFile_regfile_mem_4__0_) );
DFFPOSX1 DFFPOSX1_642 ( .CLK(clk_bF_buf81), .D(_1486_), .Q(datapath_1_RegisterFile_regfile_mem_4__1_) );
DFFPOSX1 DFFPOSX1_643 ( .CLK(clk_bF_buf17), .D(_1635_), .Q(datapath_1_RegisterFile_regfile_mem_4__2_) );
DFFPOSX1 DFFPOSX1_644 ( .CLK(clk_bF_buf12), .D(_1498_), .Q(datapath_1_RegisterFile_regfile_mem_4__3_) );
DFFPOSX1 DFFPOSX1_645 ( .CLK(clk_bF_buf82), .D(_1499_), .Q(datapath_1_RegisterFile_regfile_mem_4__4_) );
DFFPOSX1 DFFPOSX1_646 ( .CLK(clk_bF_buf109), .D(_1500_), .Q(datapath_1_RegisterFile_regfile_mem_4__5_) );
DFFPOSX1 DFFPOSX1_647 ( .CLK(clk_bF_buf28), .D(_1501_), .Q(datapath_1_RegisterFile_regfile_mem_4__6_) );
DFFPOSX1 DFFPOSX1_648 ( .CLK(clk_bF_buf32), .D(_1502_), .Q(datapath_1_RegisterFile_regfile_mem_4__7_) );
DFFPOSX1 DFFPOSX1_649 ( .CLK(clk_bF_buf19), .D(_1503_), .Q(datapath_1_RegisterFile_regfile_mem_4__8_) );
DFFPOSX1 DFFPOSX1_650 ( .CLK(clk_bF_buf100), .D(_1504_), .Q(datapath_1_RegisterFile_regfile_mem_4__9_) );
DFFPOSX1 DFFPOSX1_651 ( .CLK(clk_bF_buf81), .D(_1477_), .Q(datapath_1_RegisterFile_regfile_mem_4__10_) );
DFFPOSX1 DFFPOSX1_652 ( .CLK(clk_bF_buf110), .D(_1478_), .Q(datapath_1_RegisterFile_regfile_mem_4__11_) );
DFFPOSX1 DFFPOSX1_653 ( .CLK(clk_bF_buf107), .D(_1636_), .Q(datapath_1_RegisterFile_regfile_mem_4__12_) );
DFFPOSX1 DFFPOSX1_654 ( .CLK(clk_bF_buf87), .D(_1479_), .Q(datapath_1_RegisterFile_regfile_mem_4__13_) );
DFFPOSX1 DFFPOSX1_655 ( .CLK(clk_bF_buf111), .D(_1480_), .Q(datapath_1_RegisterFile_regfile_mem_4__14_) );
DFFPOSX1 DFFPOSX1_656 ( .CLK(clk_bF_buf101), .D(_1481_), .Q(datapath_1_RegisterFile_regfile_mem_4__15_) );
DFFPOSX1 DFFPOSX1_657 ( .CLK(clk_bF_buf101), .D(_1482_), .Q(datapath_1_RegisterFile_regfile_mem_4__16_) );
DFFPOSX1 DFFPOSX1_658 ( .CLK(clk_bF_buf23), .D(_1483_), .Q(datapath_1_RegisterFile_regfile_mem_4__17_) );
DFFPOSX1 DFFPOSX1_659 ( .CLK(clk_bF_buf16), .D(_1484_), .Q(datapath_1_RegisterFile_regfile_mem_4__18_) );
DFFPOSX1 DFFPOSX1_660 ( .CLK(clk_bF_buf54), .D(_1485_), .Q(datapath_1_RegisterFile_regfile_mem_4__19_) );
DFFPOSX1 DFFPOSX1_661 ( .CLK(clk_bF_buf54), .D(_1487_), .Q(datapath_1_RegisterFile_regfile_mem_4__20_) );
DFFPOSX1 DFFPOSX1_662 ( .CLK(clk_bF_buf103), .D(_1488_), .Q(datapath_1_RegisterFile_regfile_mem_4__21_) );
DFFPOSX1 DFFPOSX1_663 ( .CLK(clk_bF_buf87), .D(_1637_), .Q(datapath_1_RegisterFile_regfile_mem_4__22_) );
DFFPOSX1 DFFPOSX1_664 ( .CLK(clk_bF_buf7), .D(_1489_), .Q(datapath_1_RegisterFile_regfile_mem_4__23_) );
DFFPOSX1 DFFPOSX1_665 ( .CLK(clk_bF_buf70), .D(_1490_), .Q(datapath_1_RegisterFile_regfile_mem_4__24_) );
DFFPOSX1 DFFPOSX1_666 ( .CLK(clk_bF_buf17), .D(_1491_), .Q(datapath_1_RegisterFile_regfile_mem_4__25_) );
DFFPOSX1 DFFPOSX1_667 ( .CLK(clk_bF_buf53), .D(_1492_), .Q(datapath_1_RegisterFile_regfile_mem_4__26_) );
DFFPOSX1 DFFPOSX1_668 ( .CLK(clk_bF_buf7), .D(_1493_), .Q(datapath_1_RegisterFile_regfile_mem_4__27_) );
DFFPOSX1 DFFPOSX1_669 ( .CLK(clk_bF_buf32), .D(_1494_), .Q(datapath_1_RegisterFile_regfile_mem_4__28_) );
DFFPOSX1 DFFPOSX1_670 ( .CLK(clk_bF_buf110), .D(_1495_), .Q(datapath_1_RegisterFile_regfile_mem_4__29_) );
DFFPOSX1 DFFPOSX1_671 ( .CLK(clk_bF_buf53), .D(_1496_), .Q(datapath_1_RegisterFile_regfile_mem_4__30_) );
DFFPOSX1 DFFPOSX1_672 ( .CLK(clk_bF_buf11), .D(_1497_), .Q(datapath_1_RegisterFile_regfile_mem_4__31_) );
DFFPOSX1 DFFPOSX1_673 ( .CLK(clk_bF_buf30), .D(_869_), .Q(datapath_1_RegisterFile_regfile_mem_10__0_) );
DFFPOSX1 DFFPOSX1_674 ( .CLK(clk_bF_buf93), .D(_879_), .Q(datapath_1_RegisterFile_regfile_mem_10__1_) );
DFFPOSX1 DFFPOSX1_675 ( .CLK(clk_bF_buf33), .D(_1685_), .Q(datapath_1_RegisterFile_regfile_mem_10__2_) );
DFFPOSX1 DFFPOSX1_676 ( .CLK(clk_bF_buf39), .D(_884_), .Q(datapath_1_RegisterFile_regfile_mem_10__3_) );
DFFPOSX1 DFFPOSX1_677 ( .CLK(clk_bF_buf19), .D(_885_), .Q(datapath_1_RegisterFile_regfile_mem_10__4_) );
DFFPOSX1 DFFPOSX1_678 ( .CLK(clk_bF_buf45), .D(_886_), .Q(datapath_1_RegisterFile_regfile_mem_10__5_) );
DFFPOSX1 DFFPOSX1_679 ( .CLK(clk_bF_buf5), .D(_887_), .Q(datapath_1_RegisterFile_regfile_mem_10__6_) );
DFFPOSX1 DFFPOSX1_680 ( .CLK(clk_bF_buf55), .D(_888_), .Q(datapath_1_RegisterFile_regfile_mem_10__7_) );
DFFPOSX1 DFFPOSX1_681 ( .CLK(clk_bF_buf92), .D(_889_), .Q(datapath_1_RegisterFile_regfile_mem_10__8_) );
DFFPOSX1 DFFPOSX1_682 ( .CLK(clk_bF_buf45), .D(_890_), .Q(datapath_1_RegisterFile_regfile_mem_10__9_) );
DFFPOSX1 DFFPOSX1_683 ( .CLK(clk_bF_buf94), .D(_870_), .Q(datapath_1_RegisterFile_regfile_mem_10__10_) );
DFFPOSX1 DFFPOSX1_684 ( .CLK(clk_bF_buf61), .D(_871_), .Q(datapath_1_RegisterFile_regfile_mem_10__11_) );
DFFPOSX1 DFFPOSX1_685 ( .CLK(clk_bF_buf107), .D(_1686_), .Q(datapath_1_RegisterFile_regfile_mem_10__12_) );
DFFPOSX1 DFFPOSX1_686 ( .CLK(clk_bF_buf36), .D(_872_), .Q(datapath_1_RegisterFile_regfile_mem_10__13_) );
DFFPOSX1 DFFPOSX1_687 ( .CLK(clk_bF_buf74), .D(_873_), .Q(datapath_1_RegisterFile_regfile_mem_10__14_) );
DFFPOSX1 DFFPOSX1_688 ( .CLK(clk_bF_buf64), .D(_874_), .Q(datapath_1_RegisterFile_regfile_mem_10__15_) );
DFFPOSX1 DFFPOSX1_689 ( .CLK(clk_bF_buf73), .D(_875_), .Q(datapath_1_RegisterFile_regfile_mem_10__16_) );
DFFPOSX1 DFFPOSX1_690 ( .CLK(clk_bF_buf5), .D(_876_), .Q(datapath_1_RegisterFile_regfile_mem_10__17_) );
DFFPOSX1 DFFPOSX1_691 ( .CLK(clk_bF_buf7), .D(_877_), .Q(datapath_1_RegisterFile_regfile_mem_10__18_) );
DFFPOSX1 DFFPOSX1_692 ( .CLK(clk_bF_buf12), .D(_878_), .Q(datapath_1_RegisterFile_regfile_mem_10__19_) );
DFFPOSX1 DFFPOSX1_693 ( .CLK(clk_bF_buf99), .D(_880_), .Q(datapath_1_RegisterFile_regfile_mem_10__20_) );
DFFPOSX1 DFFPOSX1_694 ( .CLK(clk_bF_buf19), .D(_881_), .Q(datapath_1_RegisterFile_regfile_mem_10__21_) );
DFFPOSX1 DFFPOSX1_695 ( .CLK(clk_bF_buf45), .D(_1687_), .Q(datapath_1_RegisterFile_regfile_mem_10__22_) );
DFFPOSX1 DFFPOSX1_696 ( .CLK(clk_bF_buf46), .D(_882_), .Q(datapath_1_RegisterFile_regfile_mem_10__23_) );
DFFPOSX1 DFFPOSX1_697 ( .CLK(clk_bF_buf55), .D(_883_), .Q(datapath_1_RegisterFile_regfile_mem_10__24_) );
DFFPOSX1 DFFPOSX1_698 ( .CLK(clk_bF_buf99), .D(_1688_), .Q(datapath_1_RegisterFile_regfile_mem_10__25_) );
DFFPOSX1 DFFPOSX1_699 ( .CLK(clk_bF_buf53), .D(_1689_), .Q(datapath_1_RegisterFile_regfile_mem_10__26_) );
DFFPOSX1 DFFPOSX1_700 ( .CLK(clk_bF_buf46), .D(_1690_), .Q(datapath_1_RegisterFile_regfile_mem_10__27_) );
DFFPOSX1 DFFPOSX1_701 ( .CLK(clk_bF_buf61), .D(_1691_), .Q(datapath_1_RegisterFile_regfile_mem_10__28_) );
DFFPOSX1 DFFPOSX1_702 ( .CLK(clk_bF_buf12), .D(_1692_), .Q(datapath_1_RegisterFile_regfile_mem_10__29_) );
DFFPOSX1 DFFPOSX1_703 ( .CLK(clk_bF_buf30), .D(_1693_), .Q(datapath_1_RegisterFile_regfile_mem_10__30_) );
DFFPOSX1 DFFPOSX1_704 ( .CLK(clk_bF_buf72), .D(_1694_), .Q(datapath_1_RegisterFile_regfile_mem_10__31_) );
DFFPOSX1 DFFPOSX1_705 ( .CLK(clk_bF_buf36), .D(_1505_), .Q(datapath_1_RegisterFile_regfile_mem_5__0_) );
DFFPOSX1 DFFPOSX1_706 ( .CLK(clk_bF_buf28), .D(_1515_), .Q(datapath_1_RegisterFile_regfile_mem_5__1_) );
DFFPOSX1 DFFPOSX1_707 ( .CLK(clk_bF_buf81), .D(_1525_), .Q(datapath_1_RegisterFile_regfile_mem_5__2_) );
DFFPOSX1 DFFPOSX1_708 ( .CLK(clk_bF_buf62), .D(_1528_), .Q(datapath_1_RegisterFile_regfile_mem_5__3_) );
DFFPOSX1 DFFPOSX1_709 ( .CLK(clk_bF_buf19), .D(_1529_), .Q(datapath_1_RegisterFile_regfile_mem_5__4_) );
DFFPOSX1 DFFPOSX1_710 ( .CLK(clk_bF_buf87), .D(_1638_), .Q(datapath_1_RegisterFile_regfile_mem_5__5_) );
DFFPOSX1 DFFPOSX1_711 ( .CLK(clk_bF_buf19), .D(_1530_), .Q(datapath_1_RegisterFile_regfile_mem_5__6_) );
DFFPOSX1 DFFPOSX1_712 ( .CLK(clk_bF_buf32), .D(_1531_), .Q(datapath_1_RegisterFile_regfile_mem_5__7_) );
DFFPOSX1 DFFPOSX1_713 ( .CLK(clk_bF_buf82), .D(_1532_), .Q(datapath_1_RegisterFile_regfile_mem_5__8_) );
DFFPOSX1 DFFPOSX1_714 ( .CLK(clk_bF_buf112), .D(_1533_), .Q(datapath_1_RegisterFile_regfile_mem_5__9_) );
DFFPOSX1 DFFPOSX1_715 ( .CLK(clk_bF_buf51), .D(_1506_), .Q(datapath_1_RegisterFile_regfile_mem_5__10_) );
DFFPOSX1 DFFPOSX1_716 ( .CLK(clk_bF_buf110), .D(_1507_), .Q(datapath_1_RegisterFile_regfile_mem_5__11_) );
DFFPOSX1 DFFPOSX1_717 ( .CLK(clk_bF_buf28), .D(_1508_), .Q(datapath_1_RegisterFile_regfile_mem_5__12_) );
DFFPOSX1 DFFPOSX1_718 ( .CLK(clk_bF_buf109), .D(_1509_), .Q(datapath_1_RegisterFile_regfile_mem_5__13_) );
DFFPOSX1 DFFPOSX1_719 ( .CLK(clk_bF_buf30), .D(_1510_), .Q(datapath_1_RegisterFile_regfile_mem_5__14_) );
DFFPOSX1 DFFPOSX1_720 ( .CLK(clk_bF_buf101), .D(_1639_), .Q(datapath_1_RegisterFile_regfile_mem_5__15_) );
DFFPOSX1 DFFPOSX1_721 ( .CLK(clk_bF_buf62), .D(_1511_), .Q(datapath_1_RegisterFile_regfile_mem_5__16_) );
DFFPOSX1 DFFPOSX1_722 ( .CLK(clk_bF_buf106), .D(_1512_), .Q(datapath_1_RegisterFile_regfile_mem_5__17_) );
DFFPOSX1 DFFPOSX1_723 ( .CLK(clk_bF_buf16), .D(_1513_), .Q(datapath_1_RegisterFile_regfile_mem_5__18_) );
DFFPOSX1 DFFPOSX1_724 ( .CLK(clk_bF_buf98), .D(_1514_), .Q(datapath_1_RegisterFile_regfile_mem_5__19_) );
DFFPOSX1 DFFPOSX1_725 ( .CLK(clk_bF_buf110), .D(_1516_), .Q(datapath_1_RegisterFile_regfile_mem_5__20_) );
DFFPOSX1 DFFPOSX1_726 ( .CLK(clk_bF_buf103), .D(_1517_), .Q(datapath_1_RegisterFile_regfile_mem_5__21_) );
DFFPOSX1 DFFPOSX1_727 ( .CLK(clk_bF_buf87), .D(_1518_), .Q(datapath_1_RegisterFile_regfile_mem_5__22_) );
DFFPOSX1 DFFPOSX1_728 ( .CLK(clk_bF_buf46), .D(_1519_), .Q(datapath_1_RegisterFile_regfile_mem_5__23_) );
DFFPOSX1 DFFPOSX1_729 ( .CLK(clk_bF_buf101), .D(_1520_), .Q(datapath_1_RegisterFile_regfile_mem_5__24_) );
DFFPOSX1 DFFPOSX1_730 ( .CLK(clk_bF_buf17), .D(_1640_), .Q(datapath_1_RegisterFile_regfile_mem_5__25_) );
DFFPOSX1 DFFPOSX1_731 ( .CLK(clk_bF_buf23), .D(_1521_), .Q(datapath_1_RegisterFile_regfile_mem_5__26_) );
DFFPOSX1 DFFPOSX1_732 ( .CLK(clk_bF_buf20), .D(_1522_), .Q(datapath_1_RegisterFile_regfile_mem_5__27_) );
DFFPOSX1 DFFPOSX1_733 ( .CLK(clk_bF_buf70), .D(_1523_), .Q(datapath_1_RegisterFile_regfile_mem_5__28_) );
DFFPOSX1 DFFPOSX1_734 ( .CLK(clk_bF_buf12), .D(_1524_), .Q(datapath_1_RegisterFile_regfile_mem_5__29_) );
DFFPOSX1 DFFPOSX1_735 ( .CLK(clk_bF_buf106), .D(_1526_), .Q(datapath_1_RegisterFile_regfile_mem_5__30_) );
DFFPOSX1 DFFPOSX1_736 ( .CLK(clk_bF_buf112), .D(_1527_), .Q(datapath_1_RegisterFile_regfile_mem_5__31_) );
DFFPOSX1 DFFPOSX1_737 ( .CLK(clk_bF_buf30), .D(_1589_), .Q(datapath_1_RegisterFile_regfile_mem_9__0_) );
DFFPOSX1 DFFPOSX1_738 ( .CLK(clk_bF_buf93), .D(_1599_), .Q(datapath_1_RegisterFile_regfile_mem_9__1_) );
DFFPOSX1 DFFPOSX1_739 ( .CLK(clk_bF_buf33), .D(_1609_), .Q(datapath_1_RegisterFile_regfile_mem_9__2_) );
DFFPOSX1 DFFPOSX1_740 ( .CLK(clk_bF_buf62), .D(_1612_), .Q(datapath_1_RegisterFile_regfile_mem_9__3_) );
DFFPOSX1 DFFPOSX1_741 ( .CLK(clk_bF_buf92), .D(_1613_), .Q(datapath_1_RegisterFile_regfile_mem_9__4_) );
DFFPOSX1 DFFPOSX1_742 ( .CLK(clk_bF_buf112), .D(_1614_), .Q(datapath_1_RegisterFile_regfile_mem_9__5_) );
DFFPOSX1 DFFPOSX1_743 ( .CLK(clk_bF_buf94), .D(_1615_), .Q(datapath_1_RegisterFile_regfile_mem_9__6_) );
DFFPOSX1 DFFPOSX1_744 ( .CLK(clk_bF_buf101), .D(_1682_), .Q(datapath_1_RegisterFile_regfile_mem_9__7_) );
DFFPOSX1 DFFPOSX1_745 ( .CLK(clk_bF_buf94), .D(_1616_), .Q(datapath_1_RegisterFile_regfile_mem_9__8_) );
DFFPOSX1 DFFPOSX1_746 ( .CLK(clk_bF_buf102), .D(_1617_), .Q(datapath_1_RegisterFile_regfile_mem_9__9_) );
DFFPOSX1 DFFPOSX1_747 ( .CLK(clk_bF_buf30), .D(_1590_), .Q(datapath_1_RegisterFile_regfile_mem_9__10_) );
DFFPOSX1 DFFPOSX1_748 ( .CLK(clk_bF_buf70), .D(_1591_), .Q(datapath_1_RegisterFile_regfile_mem_9__11_) );
DFFPOSX1 DFFPOSX1_749 ( .CLK(clk_bF_buf94), .D(_1592_), .Q(datapath_1_RegisterFile_regfile_mem_9__12_) );
DFFPOSX1 DFFPOSX1_750 ( .CLK(clk_bF_buf102), .D(_1593_), .Q(datapath_1_RegisterFile_regfile_mem_9__13_) );
DFFPOSX1 DFFPOSX1_751 ( .CLK(clk_bF_buf15), .D(_1594_), .Q(datapath_1_RegisterFile_regfile_mem_9__14_) );
DFFPOSX1 DFFPOSX1_752 ( .CLK(clk_bF_buf55), .D(_1595_), .Q(datapath_1_RegisterFile_regfile_mem_9__15_) );
DFFPOSX1 DFFPOSX1_753 ( .CLK(clk_bF_buf55), .D(_1596_), .Q(datapath_1_RegisterFile_regfile_mem_9__16_) );
DFFPOSX1 DFFPOSX1_754 ( .CLK(clk_bF_buf30), .D(_1683_), .Q(datapath_1_RegisterFile_regfile_mem_9__17_) );
DFFPOSX1 DFFPOSX1_755 ( .CLK(clk_bF_buf16), .D(_1597_), .Q(datapath_1_RegisterFile_regfile_mem_9__18_) );
DFFPOSX1 DFFPOSX1_756 ( .CLK(clk_bF_buf54), .D(_1598_), .Q(datapath_1_RegisterFile_regfile_mem_9__19_) );
DFFPOSX1 DFFPOSX1_757 ( .CLK(clk_bF_buf61), .D(_1600_), .Q(datapath_1_RegisterFile_regfile_mem_9__20_) );
DFFPOSX1 DFFPOSX1_758 ( .CLK(clk_bF_buf37), .D(_1601_), .Q(datapath_1_RegisterFile_regfile_mem_9__21_) );
DFFPOSX1 DFFPOSX1_759 ( .CLK(clk_bF_buf102), .D(_1602_), .Q(datapath_1_RegisterFile_regfile_mem_9__22_) );
DFFPOSX1 DFFPOSX1_760 ( .CLK(clk_bF_buf112), .D(_1603_), .Q(datapath_1_RegisterFile_regfile_mem_9__23_) );
DFFPOSX1 DFFPOSX1_761 ( .CLK(clk_bF_buf101), .D(_1604_), .Q(datapath_1_RegisterFile_regfile_mem_9__24_) );
DFFPOSX1 DFFPOSX1_762 ( .CLK(clk_bF_buf62), .D(_1605_), .Q(datapath_1_RegisterFile_regfile_mem_9__25_) );
DFFPOSX1 DFFPOSX1_763 ( .CLK(clk_bF_buf112), .D(_1606_), .Q(datapath_1_RegisterFile_regfile_mem_9__26_) );
DFFPOSX1 DFFPOSX1_764 ( .CLK(clk_bF_buf72), .D(_1684_), .Q(datapath_1_RegisterFile_regfile_mem_9__27_) );
DFFPOSX1 DFFPOSX1_765 ( .CLK(clk_bF_buf35), .D(_1607_), .Q(datapath_1_RegisterFile_regfile_mem_9__28_) );
DFFPOSX1 DFFPOSX1_766 ( .CLK(clk_bF_buf35), .D(_1608_), .Q(datapath_1_RegisterFile_regfile_mem_9__29_) );
DFFPOSX1 DFFPOSX1_767 ( .CLK(clk_bF_buf30), .D(_1610_), .Q(datapath_1_RegisterFile_regfile_mem_9__30_) );
DFFPOSX1 DFFPOSX1_768 ( .CLK(clk_bF_buf112), .D(_1611_), .Q(datapath_1_RegisterFile_regfile_mem_9__31_) );
DFFPOSX1 DFFPOSX1_769 ( .CLK(clk_bF_buf5), .D(_1664_), .Q(datapath_1_RegisterFile_regfile_mem_8__0_) );
DFFPOSX1 DFFPOSX1_770 ( .CLK(clk_bF_buf93), .D(_1665_), .Q(datapath_1_RegisterFile_regfile_mem_8__1_) );
DFFPOSX1 DFFPOSX1_771 ( .CLK(clk_bF_buf93), .D(_1666_), .Q(datapath_1_RegisterFile_regfile_mem_8__2_) );
DFFPOSX1 DFFPOSX1_772 ( .CLK(clk_bF_buf33), .D(_1667_), .Q(datapath_1_RegisterFile_regfile_mem_8__3_) );
DFFPOSX1 DFFPOSX1_773 ( .CLK(clk_bF_buf92), .D(_1668_), .Q(datapath_1_RegisterFile_regfile_mem_8__4_) );
DFFPOSX1 DFFPOSX1_774 ( .CLK(clk_bF_buf102), .D(_1669_), .Q(datapath_1_RegisterFile_regfile_mem_8__5_) );
DFFPOSX1 DFFPOSX1_775 ( .CLK(clk_bF_buf5), .D(_1670_), .Q(datapath_1_RegisterFile_regfile_mem_8__6_) );
DFFPOSX1 DFFPOSX1_776 ( .CLK(clk_bF_buf32), .D(_1671_), .Q(datapath_1_RegisterFile_regfile_mem_8__7_) );
DFFPOSX1 DFFPOSX1_777 ( .CLK(clk_bF_buf92), .D(_1672_), .Q(datapath_1_RegisterFile_regfile_mem_8__8_) );
DFFPOSX1 DFFPOSX1_778 ( .CLK(clk_bF_buf72), .D(_1673_), .Q(datapath_1_RegisterFile_regfile_mem_8__9_) );
DFFPOSX1 DFFPOSX1_779 ( .CLK(clk_bF_buf37), .D(_1674_), .Q(datapath_1_RegisterFile_regfile_mem_8__10_) );
DFFPOSX1 DFFPOSX1_780 ( .CLK(clk_bF_buf70), .D(_1675_), .Q(datapath_1_RegisterFile_regfile_mem_8__11_) );
DFFPOSX1 DFFPOSX1_781 ( .CLK(clk_bF_buf107), .D(_1676_), .Q(datapath_1_RegisterFile_regfile_mem_8__12_) );
DFFPOSX1 DFFPOSX1_782 ( .CLK(clk_bF_buf16), .D(_1677_), .Q(datapath_1_RegisterFile_regfile_mem_8__13_) );
DFFPOSX1 DFFPOSX1_783 ( .CLK(clk_bF_buf46), .D(_1678_), .Q(datapath_1_RegisterFile_regfile_mem_8__14_) );
DFFPOSX1 DFFPOSX1_784 ( .CLK(clk_bF_buf64), .D(_1679_), .Q(datapath_1_RegisterFile_regfile_mem_8__15_) );
DFFPOSX1 DFFPOSX1_785 ( .CLK(clk_bF_buf55), .D(_1680_), .Q(datapath_1_RegisterFile_regfile_mem_8__16_) );
DFFPOSX1 DFFPOSX1_786 ( .CLK(clk_bF_buf111), .D(_1575_), .Q(datapath_1_RegisterFile_regfile_mem_8__17_) );
DFFPOSX1 DFFPOSX1_787 ( .CLK(clk_bF_buf7), .D(_1576_), .Q(datapath_1_RegisterFile_regfile_mem_8__18_) );
DFFPOSX1 DFFPOSX1_788 ( .CLK(clk_bF_buf54), .D(_1577_), .Q(datapath_1_RegisterFile_regfile_mem_8__19_) );
DFFPOSX1 DFFPOSX1_789 ( .CLK(clk_bF_buf99), .D(_1578_), .Q(datapath_1_RegisterFile_regfile_mem_8__20_) );
DFFPOSX1 DFFPOSX1_790 ( .CLK(clk_bF_buf92), .D(_1579_), .Q(datapath_1_RegisterFile_regfile_mem_8__21_) );
DFFPOSX1 DFFPOSX1_791 ( .CLK(clk_bF_buf102), .D(_1580_), .Q(datapath_1_RegisterFile_regfile_mem_8__22_) );
DFFPOSX1 DFFPOSX1_792 ( .CLK(clk_bF_buf46), .D(_1581_), .Q(datapath_1_RegisterFile_regfile_mem_8__23_) );
DFFPOSX1 DFFPOSX1_793 ( .CLK(clk_bF_buf55), .D(_1681_), .Q(datapath_1_RegisterFile_regfile_mem_8__24_) );
DFFPOSX1 DFFPOSX1_794 ( .CLK(clk_bF_buf62), .D(_1582_), .Q(datapath_1_RegisterFile_regfile_mem_8__25_) );
DFFPOSX1 DFFPOSX1_795 ( .CLK(clk_bF_buf53), .D(_1583_), .Q(datapath_1_RegisterFile_regfile_mem_8__26_) );
DFFPOSX1 DFFPOSX1_796 ( .CLK(clk_bF_buf74), .D(_1584_), .Q(datapath_1_RegisterFile_regfile_mem_8__27_) );
DFFPOSX1 DFFPOSX1_797 ( .CLK(clk_bF_buf35), .D(_1585_), .Q(datapath_1_RegisterFile_regfile_mem_8__28_) );
DFFPOSX1 DFFPOSX1_798 ( .CLK(clk_bF_buf54), .D(_1586_), .Q(datapath_1_RegisterFile_regfile_mem_8__29_) );
DFFPOSX1 DFFPOSX1_799 ( .CLK(clk_bF_buf74), .D(_1587_), .Q(datapath_1_RegisterFile_regfile_mem_8__30_) );
DFFPOSX1 DFFPOSX1_800 ( .CLK(clk_bF_buf20), .D(_1588_), .Q(datapath_1_RegisterFile_regfile_mem_8__31_) );
DFFPOSX1 DFFPOSX1_801 ( .CLK(clk_bF_buf106), .D(_1258_), .Q(datapath_1_RegisterFile_regfile_mem_26__0_) );
DFFPOSX1 DFFPOSX1_802 ( .CLK(clk_bF_buf58), .D(_1268_), .Q(datapath_1_RegisterFile_regfile_mem_26__1_) );
DFFPOSX1 DFFPOSX1_803 ( .CLK(clk_bF_buf3), .D(_1278_), .Q(datapath_1_RegisterFile_regfile_mem_26__2_) );
DFFPOSX1 DFFPOSX1_804 ( .CLK(clk_bF_buf89), .D(_1281_), .Q(datapath_1_RegisterFile_regfile_mem_26__3_) );
DFFPOSX1 DFFPOSX1_805 ( .CLK(clk_bF_buf26), .D(_1829_), .Q(datapath_1_RegisterFile_regfile_mem_26__4_) );
DFFPOSX1 DFFPOSX1_806 ( .CLK(clk_bF_buf56), .D(_1282_), .Q(datapath_1_RegisterFile_regfile_mem_26__5_) );
DFFPOSX1 DFFPOSX1_807 ( .CLK(clk_bF_buf113), .D(_1283_), .Q(datapath_1_RegisterFile_regfile_mem_26__6_) );
DFFPOSX1 DFFPOSX1_808 ( .CLK(clk_bF_buf98), .D(_1284_), .Q(datapath_1_RegisterFile_regfile_mem_26__7_) );
DFFPOSX1 DFFPOSX1_809 ( .CLK(clk_bF_buf96), .D(_1285_), .Q(datapath_1_RegisterFile_regfile_mem_26__8_) );
DFFPOSX1 DFFPOSX1_810 ( .CLK(clk_bF_buf79), .D(_1286_), .Q(datapath_1_RegisterFile_regfile_mem_26__9_) );
DFFPOSX1 DFFPOSX1_811 ( .CLK(clk_bF_buf79), .D(_1259_), .Q(datapath_1_RegisterFile_regfile_mem_26__10_) );
DFFPOSX1 DFFPOSX1_812 ( .CLK(clk_bF_buf40), .D(_1260_), .Q(datapath_1_RegisterFile_regfile_mem_26__11_) );
DFFPOSX1 DFFPOSX1_813 ( .CLK(clk_bF_buf41), .D(_1261_), .Q(datapath_1_RegisterFile_regfile_mem_26__12_) );
DFFPOSX1 DFFPOSX1_814 ( .CLK(clk_bF_buf34), .D(_1262_), .Q(datapath_1_RegisterFile_regfile_mem_26__13_) );
DFFPOSX1 DFFPOSX1_815 ( .CLK(clk_bF_buf48), .D(_1830_), .Q(datapath_1_RegisterFile_regfile_mem_26__14_) );
DFFPOSX1 DFFPOSX1_816 ( .CLK(clk_bF_buf40), .D(_1263_), .Q(datapath_1_RegisterFile_regfile_mem_26__15_) );
DFFPOSX1 DFFPOSX1_817 ( .CLK(clk_bF_buf40), .D(_1264_), .Q(datapath_1_RegisterFile_regfile_mem_26__16_) );
DFFPOSX1 DFFPOSX1_818 ( .CLK(clk_bF_buf26), .D(_1265_), .Q(datapath_1_RegisterFile_regfile_mem_26__17_) );
DFFPOSX1 DFFPOSX1_819 ( .CLK(clk_bF_buf90), .D(_1266_), .Q(datapath_1_RegisterFile_regfile_mem_26__18_) );
DFFPOSX1 DFFPOSX1_820 ( .CLK(clk_bF_buf3), .D(_1267_), .Q(datapath_1_RegisterFile_regfile_mem_26__19_) );
DFFPOSX1 DFFPOSX1_821 ( .CLK(clk_bF_buf49), .D(_1269_), .Q(datapath_1_RegisterFile_regfile_mem_26__20_) );
DFFPOSX1 DFFPOSX1_822 ( .CLK(clk_bF_buf76), .D(_1270_), .Q(datapath_1_RegisterFile_regfile_mem_26__21_) );
DFFPOSX1 DFFPOSX1_823 ( .CLK(clk_bF_buf105), .D(_1271_), .Q(datapath_1_RegisterFile_regfile_mem_26__22_) );
DFFPOSX1 DFFPOSX1_824 ( .CLK(clk_bF_buf79), .D(_1272_), .Q(datapath_1_RegisterFile_regfile_mem_26__23_) );
DFFPOSX1 DFFPOSX1_825 ( .CLK(clk_bF_buf3), .D(_1831_), .Q(datapath_1_RegisterFile_regfile_mem_26__24_) );
DFFPOSX1 DFFPOSX1_826 ( .CLK(clk_bF_buf58), .D(_1273_), .Q(datapath_1_RegisterFile_regfile_mem_26__25_) );
DFFPOSX1 DFFPOSX1_827 ( .CLK(clk_bF_buf105), .D(_1274_), .Q(datapath_1_RegisterFile_regfile_mem_26__26_) );
DFFPOSX1 DFFPOSX1_828 ( .CLK(clk_bF_buf56), .D(_1275_), .Q(datapath_1_RegisterFile_regfile_mem_26__27_) );
DFFPOSX1 DFFPOSX1_829 ( .CLK(clk_bF_buf70), .D(_1276_), .Q(datapath_1_RegisterFile_regfile_mem_26__28_) );
DFFPOSX1 DFFPOSX1_830 ( .CLK(clk_bF_buf41), .D(_1277_), .Q(datapath_1_RegisterFile_regfile_mem_26__29_) );
DFFPOSX1 DFFPOSX1_831 ( .CLK(clk_bF_buf88), .D(_1279_), .Q(datapath_1_RegisterFile_regfile_mem_26__30_) );
DFFPOSX1 DFFPOSX1_832 ( .CLK(clk_bF_buf48), .D(_1280_), .Q(datapath_1_RegisterFile_regfile_mem_26__31_) );
DFFPOSX1 DFFPOSX1_833 ( .CLK(clk_bF_buf77), .D(_1238_), .Q(datapath_1_RegisterFile_regfile_mem_25__0_) );
DFFPOSX1 DFFPOSX1_834 ( .CLK(clk_bF_buf58), .D(_1248_), .Q(datapath_1_RegisterFile_regfile_mem_25__1_) );
DFFPOSX1 DFFPOSX1_835 ( .CLK(clk_bF_buf95), .D(_1251_), .Q(datapath_1_RegisterFile_regfile_mem_25__2_) );
DFFPOSX1 DFFPOSX1_836 ( .CLK(clk_bF_buf49), .D(_1252_), .Q(datapath_1_RegisterFile_regfile_mem_25__3_) );
DFFPOSX1 DFFPOSX1_837 ( .CLK(clk_bF_buf96), .D(_1253_), .Q(datapath_1_RegisterFile_regfile_mem_25__4_) );
DFFPOSX1 DFFPOSX1_838 ( .CLK(clk_bF_buf56), .D(_1254_), .Q(datapath_1_RegisterFile_regfile_mem_25__5_) );
DFFPOSX1 DFFPOSX1_839 ( .CLK(clk_bF_buf1), .D(_1255_), .Q(datapath_1_RegisterFile_regfile_mem_25__6_) );
DFFPOSX1 DFFPOSX1_840 ( .CLK(clk_bF_buf89), .D(_1256_), .Q(datapath_1_RegisterFile_regfile_mem_25__7_) );
DFFPOSX1 DFFPOSX1_841 ( .CLK(clk_bF_buf58), .D(_1257_), .Q(datapath_1_RegisterFile_regfile_mem_25__8_) );
DFFPOSX1 DFFPOSX1_842 ( .CLK(clk_bF_buf79), .D(_1817_), .Q(datapath_1_RegisterFile_regfile_mem_25__9_) );
DFFPOSX1 DFFPOSX1_843 ( .CLK(clk_bF_buf100), .D(_1239_), .Q(datapath_1_RegisterFile_regfile_mem_25__10_) );
DFFPOSX1 DFFPOSX1_844 ( .CLK(clk_bF_buf40), .D(_1240_), .Q(datapath_1_RegisterFile_regfile_mem_25__11_) );
DFFPOSX1 DFFPOSX1_845 ( .CLK(clk_bF_buf41), .D(_1241_), .Q(datapath_1_RegisterFile_regfile_mem_25__12_) );
DFFPOSX1 DFFPOSX1_846 ( .CLK(clk_bF_buf77), .D(_1242_), .Q(datapath_1_RegisterFile_regfile_mem_25__13_) );
DFFPOSX1 DFFPOSX1_847 ( .CLK(clk_bF_buf56), .D(_1243_), .Q(datapath_1_RegisterFile_regfile_mem_25__14_) );
DFFPOSX1 DFFPOSX1_848 ( .CLK(clk_bF_buf41), .D(_1244_), .Q(datapath_1_RegisterFile_regfile_mem_25__15_) );
DFFPOSX1 DFFPOSX1_849 ( .CLK(clk_bF_buf59), .D(_1245_), .Q(datapath_1_RegisterFile_regfile_mem_25__16_) );
DFFPOSX1 DFFPOSX1_850 ( .CLK(clk_bF_buf60), .D(_1246_), .Q(datapath_1_RegisterFile_regfile_mem_25__17_) );
DFFPOSX1 DFFPOSX1_851 ( .CLK(clk_bF_buf56), .D(_1247_), .Q(datapath_1_RegisterFile_regfile_mem_25__18_) );
DFFPOSX1 DFFPOSX1_852 ( .CLK(clk_bF_buf2), .D(_1818_), .Q(datapath_1_RegisterFile_regfile_mem_25__19_) );
DFFPOSX1 DFFPOSX1_853 ( .CLK(clk_bF_buf70), .D(_1249_), .Q(datapath_1_RegisterFile_regfile_mem_25__20_) );
DFFPOSX1 DFFPOSX1_854 ( .CLK(clk_bF_buf1), .D(_1250_), .Q(datapath_1_RegisterFile_regfile_mem_25__21_) );
DFFPOSX1 DFFPOSX1_855 ( .CLK(clk_bF_buf29), .D(_1819_), .Q(datapath_1_RegisterFile_regfile_mem_25__22_) );
DFFPOSX1 DFFPOSX1_856 ( .CLK(clk_bF_buf67), .D(_1820_), .Q(datapath_1_RegisterFile_regfile_mem_25__23_) );
DFFPOSX1 DFFPOSX1_857 ( .CLK(clk_bF_buf38), .D(_1821_), .Q(datapath_1_RegisterFile_regfile_mem_25__24_) );
DFFPOSX1 DFFPOSX1_858 ( .CLK(clk_bF_buf58), .D(_1822_), .Q(datapath_1_RegisterFile_regfile_mem_25__25_) );
DFFPOSX1 DFFPOSX1_859 ( .CLK(clk_bF_buf34), .D(_1823_), .Q(datapath_1_RegisterFile_regfile_mem_25__26_) );
DFFPOSX1 DFFPOSX1_860 ( .CLK(clk_bF_buf56), .D(_1824_), .Q(datapath_1_RegisterFile_regfile_mem_25__27_) );
DFFPOSX1 DFFPOSX1_861 ( .CLK(clk_bF_buf70), .D(_1825_), .Q(datapath_1_RegisterFile_regfile_mem_25__28_) );
DFFPOSX1 DFFPOSX1_862 ( .CLK(clk_bF_buf95), .D(_1826_), .Q(datapath_1_RegisterFile_regfile_mem_25__29_) );
DFFPOSX1 DFFPOSX1_863 ( .CLK(clk_bF_buf77), .D(_1827_), .Q(datapath_1_RegisterFile_regfile_mem_25__30_) );
DFFPOSX1 DFFPOSX1_864 ( .CLK(clk_bF_buf29), .D(_1828_), .Q(datapath_1_RegisterFile_regfile_mem_25__31_) );
DFFPOSX1 DFFPOSX1_865 ( .CLK(clk_bF_buf29), .D(_1198_), .Q(datapath_1_RegisterFile_regfile_mem_23__0_) );
DFFPOSX1 DFFPOSX1_866 ( .CLK(clk_bF_buf65), .D(_1204_), .Q(datapath_1_RegisterFile_regfile_mem_23__1_) );
DFFPOSX1 DFFPOSX1_867 ( .CLK(clk_bF_buf38), .D(_1209_), .Q(datapath_1_RegisterFile_regfile_mem_23__2_) );
DFFPOSX1 DFFPOSX1_868 ( .CLK(clk_bF_buf89), .D(_1793_), .Q(datapath_1_RegisterFile_regfile_mem_23__3_) );
DFFPOSX1 DFFPOSX1_869 ( .CLK(clk_bF_buf26), .D(_1212_), .Q(datapath_1_RegisterFile_regfile_mem_23__4_) );
DFFPOSX1 DFFPOSX1_870 ( .CLK(clk_bF_buf4), .D(_1213_), .Q(datapath_1_RegisterFile_regfile_mem_23__5_) );
DFFPOSX1 DFFPOSX1_871 ( .CLK(clk_bF_buf65), .D(_1214_), .Q(datapath_1_RegisterFile_regfile_mem_23__6_) );
DFFPOSX1 DFFPOSX1_872 ( .CLK(clk_bF_buf75), .D(_1215_), .Q(datapath_1_RegisterFile_regfile_mem_23__7_) );
DFFPOSX1 DFFPOSX1_873 ( .CLK(clk_bF_buf96), .D(_1216_), .Q(datapath_1_RegisterFile_regfile_mem_23__8_) );
DFFPOSX1 DFFPOSX1_874 ( .CLK(clk_bF_buf29), .D(_1217_), .Q(datapath_1_RegisterFile_regfile_mem_23__9_) );
DFFPOSX1 DFFPOSX1_875 ( .CLK(clk_bF_buf80), .D(_1199_), .Q(datapath_1_RegisterFile_regfile_mem_23__10_) );
DFFPOSX1 DFFPOSX1_876 ( .CLK(clk_bF_buf25), .D(_1200_), .Q(datapath_1_RegisterFile_regfile_mem_23__11_) );
DFFPOSX1 DFFPOSX1_877 ( .CLK(clk_bF_buf59), .D(_1201_), .Q(datapath_1_RegisterFile_regfile_mem_23__12_) );
DFFPOSX1 DFFPOSX1_878 ( .CLK(clk_bF_buf47), .D(_1794_), .Q(datapath_1_RegisterFile_regfile_mem_23__13_) );
DFFPOSX1 DFFPOSX1_879 ( .CLK(clk_bF_buf90), .D(_1202_), .Q(datapath_1_RegisterFile_regfile_mem_23__14_) );
DFFPOSX1 DFFPOSX1_880 ( .CLK(clk_bF_buf42), .D(_1203_), .Q(datapath_1_RegisterFile_regfile_mem_23__15_) );
DFFPOSX1 DFFPOSX1_881 ( .CLK(clk_bF_buf78), .D(_1795_), .Q(datapath_1_RegisterFile_regfile_mem_23__16_) );
DFFPOSX1 DFFPOSX1_882 ( .CLK(clk_bF_buf76), .D(_1796_), .Q(datapath_1_RegisterFile_regfile_mem_23__17_) );
DFFPOSX1 DFFPOSX1_883 ( .CLK(clk_bF_buf80), .D(_1797_), .Q(datapath_1_RegisterFile_regfile_mem_23__18_) );
DFFPOSX1 DFFPOSX1_884 ( .CLK(clk_bF_buf75), .D(_1798_), .Q(datapath_1_RegisterFile_regfile_mem_23__19_) );
DFFPOSX1 DFFPOSX1_885 ( .CLK(clk_bF_buf6), .D(_1799_), .Q(datapath_1_RegisterFile_regfile_mem_23__20_) );
DFFPOSX1 DFFPOSX1_886 ( .CLK(clk_bF_buf76), .D(_1800_), .Q(datapath_1_RegisterFile_regfile_mem_23__21_) );
DFFPOSX1 DFFPOSX1_887 ( .CLK(clk_bF_buf105), .D(_1801_), .Q(datapath_1_RegisterFile_regfile_mem_23__22_) );
DFFPOSX1 DFFPOSX1_888 ( .CLK(clk_bF_buf113), .D(_1802_), .Q(datapath_1_RegisterFile_regfile_mem_23__23_) );
DFFPOSX1 DFFPOSX1_889 ( .CLK(clk_bF_buf85), .D(_1803_), .Q(datapath_1_RegisterFile_regfile_mem_23__24_) );
DFFPOSX1 DFFPOSX1_890 ( .CLK(clk_bF_buf59), .D(_1804_), .Q(datapath_1_RegisterFile_regfile_mem_23__25_) );
DFFPOSX1 DFFPOSX1_891 ( .CLK(clk_bF_buf47), .D(_1205_), .Q(datapath_1_RegisterFile_regfile_mem_23__26_) );
DFFPOSX1 DFFPOSX1_892 ( .CLK(clk_bF_buf90), .D(_1206_), .Q(datapath_1_RegisterFile_regfile_mem_23__27_) );
DFFPOSX1 DFFPOSX1_893 ( .CLK(clk_bF_buf38), .D(_1207_), .Q(datapath_1_RegisterFile_regfile_mem_23__28_) );
DFFPOSX1 DFFPOSX1_894 ( .CLK(clk_bF_buf95), .D(_1208_), .Q(datapath_1_RegisterFile_regfile_mem_23__29_) );
DFFPOSX1 DFFPOSX1_895 ( .CLK(clk_bF_buf66), .D(_1210_), .Q(datapath_1_RegisterFile_regfile_mem_23__30_) );
DFFPOSX1 DFFPOSX1_896 ( .CLK(clk_bF_buf44), .D(_1211_), .Q(datapath_1_RegisterFile_regfile_mem_23__31_) );
DFFPOSX1 DFFPOSX1_897 ( .CLK(clk_bF_buf1), .D(_1832_), .Q(datapath_1_RegisterFile_regfile_mem_27__0_) );
DFFPOSX1 DFFPOSX1_898 ( .CLK(clk_bF_buf65), .D(_1833_), .Q(datapath_1_RegisterFile_regfile_mem_27__1_) );
DFFPOSX1 DFFPOSX1_899 ( .CLK(clk_bF_buf40), .D(_1305_), .Q(datapath_1_RegisterFile_regfile_mem_27__2_) );
DFFPOSX1 DFFPOSX1_900 ( .CLK(clk_bF_buf89), .D(_1308_), .Q(datapath_1_RegisterFile_regfile_mem_27__3_) );
DFFPOSX1 DFFPOSX1_901 ( .CLK(clk_bF_buf57), .D(_1309_), .Q(datapath_1_RegisterFile_regfile_mem_27__4_) );
DFFPOSX1 DFFPOSX1_902 ( .CLK(clk_bF_buf56), .D(_1310_), .Q(datapath_1_RegisterFile_regfile_mem_27__5_) );
DFFPOSX1 DFFPOSX1_903 ( .CLK(clk_bF_buf67), .D(_1311_), .Q(datapath_1_RegisterFile_regfile_mem_27__6_) );
DFFPOSX1 DFFPOSX1_904 ( .CLK(clk_bF_buf49), .D(_1312_), .Q(datapath_1_RegisterFile_regfile_mem_27__7_) );
DFFPOSX1 DFFPOSX1_905 ( .CLK(clk_bF_buf65), .D(_1313_), .Q(datapath_1_RegisterFile_regfile_mem_27__8_) );
DFFPOSX1 DFFPOSX1_906 ( .CLK(clk_bF_buf79), .D(_1834_), .Q(datapath_1_RegisterFile_regfile_mem_27__9_) );
DFFPOSX1 DFFPOSX1_907 ( .CLK(clk_bF_buf29), .D(_1287_), .Q(datapath_1_RegisterFile_regfile_mem_27__10_) );
DFFPOSX1 DFFPOSX1_908 ( .CLK(clk_bF_buf63), .D(_1288_), .Q(datapath_1_RegisterFile_regfile_mem_27__11_) );
DFFPOSX1 DFFPOSX1_909 ( .CLK(clk_bF_buf41), .D(_1289_), .Q(datapath_1_RegisterFile_regfile_mem_27__12_) );
DFFPOSX1 DFFPOSX1_910 ( .CLK(clk_bF_buf47), .D(_1290_), .Q(datapath_1_RegisterFile_regfile_mem_27__13_) );
DFFPOSX1 DFFPOSX1_911 ( .CLK(clk_bF_buf48), .D(_1291_), .Q(datapath_1_RegisterFile_regfile_mem_27__14_) );
DFFPOSX1 DFFPOSX1_912 ( .CLK(clk_bF_buf41), .D(_1292_), .Q(datapath_1_RegisterFile_regfile_mem_27__15_) );
DFFPOSX1 DFFPOSX1_913 ( .CLK(clk_bF_buf3), .D(_1293_), .Q(datapath_1_RegisterFile_regfile_mem_27__16_) );
DFFPOSX1 DFFPOSX1_914 ( .CLK(clk_bF_buf88), .D(_1294_), .Q(datapath_1_RegisterFile_regfile_mem_27__17_) );
DFFPOSX1 DFFPOSX1_915 ( .CLK(clk_bF_buf90), .D(_1295_), .Q(datapath_1_RegisterFile_regfile_mem_27__18_) );
DFFPOSX1 DFFPOSX1_916 ( .CLK(clk_bF_buf51), .D(_1835_), .Q(datapath_1_RegisterFile_regfile_mem_27__19_) );
DFFPOSX1 DFFPOSX1_917 ( .CLK(clk_bF_buf49), .D(_1296_), .Q(datapath_1_RegisterFile_regfile_mem_27__20_) );
DFFPOSX1 DFFPOSX1_918 ( .CLK(clk_bF_buf57), .D(_1297_), .Q(datapath_1_RegisterFile_regfile_mem_27__21_) );
DFFPOSX1 DFFPOSX1_919 ( .CLK(clk_bF_buf29), .D(_1298_), .Q(datapath_1_RegisterFile_regfile_mem_27__22_) );
DFFPOSX1 DFFPOSX1_920 ( .CLK(clk_bF_buf67), .D(_1299_), .Q(datapath_1_RegisterFile_regfile_mem_27__23_) );
DFFPOSX1 DFFPOSX1_921 ( .CLK(clk_bF_buf85), .D(_1300_), .Q(datapath_1_RegisterFile_regfile_mem_27__24_) );
DFFPOSX1 DFFPOSX1_922 ( .CLK(clk_bF_buf59), .D(_1301_), .Q(datapath_1_RegisterFile_regfile_mem_27__25_) );
DFFPOSX1 DFFPOSX1_923 ( .CLK(clk_bF_buf66), .D(_1302_), .Q(datapath_1_RegisterFile_regfile_mem_27__26_) );
DFFPOSX1 DFFPOSX1_924 ( .CLK(clk_bF_buf48), .D(_1303_), .Q(datapath_1_RegisterFile_regfile_mem_27__27_) );
DFFPOSX1 DFFPOSX1_925 ( .CLK(clk_bF_buf49), .D(_1304_), .Q(datapath_1_RegisterFile_regfile_mem_27__28_) );
DFFPOSX1 DFFPOSX1_926 ( .CLK(clk_bF_buf41), .D(_1836_), .Q(datapath_1_RegisterFile_regfile_mem_27__29_) );
DFFPOSX1 DFFPOSX1_927 ( .CLK(clk_bF_buf88), .D(_1306_), .Q(datapath_1_RegisterFile_regfile_mem_27__30_) );
DFFPOSX1 DFFPOSX1_928 ( .CLK(clk_bF_buf48), .D(_1307_), .Q(datapath_1_RegisterFile_regfile_mem_27__31_) );
DFFPOSX1 DFFPOSX1_929 ( .CLK(clk_bF_buf77), .D(_1338_), .Q(datapath_1_RegisterFile_regfile_mem_29__0_) );
DFFPOSX1 DFFPOSX1_930 ( .CLK(clk_bF_buf21), .D(_1348_), .Q(datapath_1_RegisterFile_regfile_mem_29__1_) );
DFFPOSX1 DFFPOSX1_931 ( .CLK(clk_bF_buf2), .D(_1358_), .Q(datapath_1_RegisterFile_regfile_mem_29__2_) );
DFFPOSX1 DFFPOSX1_932 ( .CLK(clk_bF_buf41), .D(_1361_), .Q(datapath_1_RegisterFile_regfile_mem_29__3_) );
DFFPOSX1 DFFPOSX1_933 ( .CLK(clk_bF_buf96), .D(_1362_), .Q(datapath_1_RegisterFile_regfile_mem_29__4_) );
DFFPOSX1 DFFPOSX1_934 ( .CLK(clk_bF_buf56), .D(_1363_), .Q(datapath_1_RegisterFile_regfile_mem_29__5_) );
DFFPOSX1 DFFPOSX1_935 ( .CLK(clk_bF_buf1), .D(_1364_), .Q(datapath_1_RegisterFile_regfile_mem_29__6_) );
DFFPOSX1 DFFPOSX1_936 ( .CLK(clk_bF_buf89), .D(_1365_), .Q(datapath_1_RegisterFile_regfile_mem_29__7_) );
DFFPOSX1 DFFPOSX1_937 ( .CLK(clk_bF_buf113), .D(_1366_), .Q(datapath_1_RegisterFile_regfile_mem_29__8_) );
DFFPOSX1 DFFPOSX1_938 ( .CLK(clk_bF_buf79), .D(_1845_), .Q(datapath_1_RegisterFile_regfile_mem_29__9_) );
DFFPOSX1 DFFPOSX1_939 ( .CLK(clk_bF_buf79), .D(_1339_), .Q(datapath_1_RegisterFile_regfile_mem_29__10_) );
DFFPOSX1 DFFPOSX1_940 ( .CLK(clk_bF_buf89), .D(_1340_), .Q(datapath_1_RegisterFile_regfile_mem_29__11_) );
DFFPOSX1 DFFPOSX1_941 ( .CLK(clk_bF_buf2), .D(_1341_), .Q(datapath_1_RegisterFile_regfile_mem_29__12_) );
DFFPOSX1 DFFPOSX1_942 ( .CLK(clk_bF_buf13), .D(_1342_), .Q(datapath_1_RegisterFile_regfile_mem_29__13_) );
DFFPOSX1 DFFPOSX1_943 ( .CLK(clk_bF_buf100), .D(_1343_), .Q(datapath_1_RegisterFile_regfile_mem_29__14_) );
DFFPOSX1 DFFPOSX1_944 ( .CLK(clk_bF_buf41), .D(_1344_), .Q(datapath_1_RegisterFile_regfile_mem_29__15_) );
DFFPOSX1 DFFPOSX1_945 ( .CLK(clk_bF_buf59), .D(_1345_), .Q(datapath_1_RegisterFile_regfile_mem_29__16_) );
DFFPOSX1 DFFPOSX1_946 ( .CLK(clk_bF_buf77), .D(_1346_), .Q(datapath_1_RegisterFile_regfile_mem_29__17_) );
DFFPOSX1 DFFPOSX1_947 ( .CLK(clk_bF_buf56), .D(_1347_), .Q(datapath_1_RegisterFile_regfile_mem_29__18_) );
DFFPOSX1 DFFPOSX1_948 ( .CLK(clk_bF_buf51), .D(_1846_), .Q(datapath_1_RegisterFile_regfile_mem_29__19_) );
DFFPOSX1 DFFPOSX1_949 ( .CLK(clk_bF_buf70), .D(_1349_), .Q(datapath_1_RegisterFile_regfile_mem_29__20_) );
DFFPOSX1 DFFPOSX1_950 ( .CLK(clk_bF_buf67), .D(_1350_), .Q(datapath_1_RegisterFile_regfile_mem_29__21_) );
DFFPOSX1 DFFPOSX1_951 ( .CLK(clk_bF_buf13), .D(_1351_), .Q(datapath_1_RegisterFile_regfile_mem_29__22_) );
DFFPOSX1 DFFPOSX1_952 ( .CLK(clk_bF_buf51), .D(_1352_), .Q(datapath_1_RegisterFile_regfile_mem_29__23_) );
DFFPOSX1 DFFPOSX1_953 ( .CLK(clk_bF_buf59), .D(_1353_), .Q(datapath_1_RegisterFile_regfile_mem_29__24_) );
DFFPOSX1 DFFPOSX1_954 ( .CLK(clk_bF_buf78), .D(_1354_), .Q(datapath_1_RegisterFile_regfile_mem_29__25_) );
DFFPOSX1 DFFPOSX1_955 ( .CLK(clk_bF_buf13), .D(_1355_), .Q(datapath_1_RegisterFile_regfile_mem_29__26_) );
DFFPOSX1 DFFPOSX1_956 ( .CLK(clk_bF_buf86), .D(_1356_), .Q(datapath_1_RegisterFile_regfile_mem_29__27_) );
DFFPOSX1 DFFPOSX1_957 ( .CLK(clk_bF_buf89), .D(_1357_), .Q(datapath_1_RegisterFile_regfile_mem_29__28_) );
DFFPOSX1 DFFPOSX1_958 ( .CLK(clk_bF_buf31), .D(_1847_), .Q(datapath_1_RegisterFile_regfile_mem_29__29_) );
DFFPOSX1 DFFPOSX1_959 ( .CLK(clk_bF_buf76), .D(_1359_), .Q(datapath_1_RegisterFile_regfile_mem_29__30_) );
DFFPOSX1 DFFPOSX1_960 ( .CLK(clk_bF_buf100), .D(_1360_), .Q(datapath_1_RegisterFile_regfile_mem_29__31_) );
DFFPOSX1 DFFPOSX1_961 ( .CLK(clk_bF_buf1), .D(_1848_), .Q(datapath_1_RegisterFile_regfile_mem_30__0_) );
DFFPOSX1 DFFPOSX1_962 ( .CLK(clk_bF_buf14), .D(_1849_), .Q(datapath_1_RegisterFile_regfile_mem_30__1_) );
DFFPOSX1 DFFPOSX1_963 ( .CLK(clk_bF_buf2), .D(_1850_), .Q(datapath_1_RegisterFile_regfile_mem_30__2_) );
DFFPOSX1 DFFPOSX1_964 ( .CLK(clk_bF_buf40), .D(_1851_), .Q(datapath_1_RegisterFile_regfile_mem_30__3_) );
DFFPOSX1 DFFPOSX1_965 ( .CLK(clk_bF_buf76), .D(_1852_), .Q(datapath_1_RegisterFile_regfile_mem_30__4_) );
DFFPOSX1 DFFPOSX1_966 ( .CLK(clk_bF_buf29), .D(_1853_), .Q(datapath_1_RegisterFile_regfile_mem_30__5_) );
DFFPOSX1 DFFPOSX1_967 ( .CLK(clk_bF_buf67), .D(_1854_), .Q(datapath_1_RegisterFile_regfile_mem_30__6_) );
DFFPOSX1 DFFPOSX1_968 ( .CLK(clk_bF_buf98), .D(_1416_), .Q(datapath_1_RegisterFile_regfile_mem_30__7_) );
DFFPOSX1 DFFPOSX1_969 ( .CLK(clk_bF_buf76), .D(_1417_), .Q(datapath_1_RegisterFile_regfile_mem_30__8_) );
DFFPOSX1 DFFPOSX1_970 ( .CLK(clk_bF_buf79), .D(_1418_), .Q(datapath_1_RegisterFile_regfile_mem_30__9_) );
DFFPOSX1 DFFPOSX1_971 ( .CLK(clk_bF_buf29), .D(_1396_), .Q(datapath_1_RegisterFile_regfile_mem_30__10_) );
DFFPOSX1 DFFPOSX1_972 ( .CLK(clk_bF_buf49), .D(_1397_), .Q(datapath_1_RegisterFile_regfile_mem_30__11_) );
DFFPOSX1 DFFPOSX1_973 ( .CLK(clk_bF_buf51), .D(_1398_), .Q(datapath_1_RegisterFile_regfile_mem_30__12_) );
DFFPOSX1 DFFPOSX1_974 ( .CLK(clk_bF_buf34), .D(_1399_), .Q(datapath_1_RegisterFile_regfile_mem_30__13_) );
DFFPOSX1 DFFPOSX1_975 ( .CLK(clk_bF_buf86), .D(_1855_), .Q(datapath_1_RegisterFile_regfile_mem_30__14_) );
DFFPOSX1 DFFPOSX1_976 ( .CLK(clk_bF_buf14), .D(_1400_), .Q(datapath_1_RegisterFile_regfile_mem_30__15_) );
DFFPOSX1 DFFPOSX1_977 ( .CLK(clk_bF_buf95), .D(_1401_), .Q(datapath_1_RegisterFile_regfile_mem_30__16_) );
DFFPOSX1 DFFPOSX1_978 ( .CLK(clk_bF_buf77), .D(_1402_), .Q(datapath_1_RegisterFile_regfile_mem_30__17_) );
DFFPOSX1 DFFPOSX1_979 ( .CLK(clk_bF_buf86), .D(_1403_), .Q(datapath_1_RegisterFile_regfile_mem_30__18_) );
DFFPOSX1 DFFPOSX1_980 ( .CLK(clk_bF_buf51), .D(_1404_), .Q(datapath_1_RegisterFile_regfile_mem_30__19_) );
DFFPOSX1 DFFPOSX1_981 ( .CLK(clk_bF_buf49), .D(_1405_), .Q(datapath_1_RegisterFile_regfile_mem_30__20_) );
DFFPOSX1 DFFPOSX1_982 ( .CLK(clk_bF_buf1), .D(_1406_), .Q(datapath_1_RegisterFile_regfile_mem_30__21_) );
DFFPOSX1 DFFPOSX1_983 ( .CLK(clk_bF_buf34), .D(_1407_), .Q(datapath_1_RegisterFile_regfile_mem_30__22_) );
DFFPOSX1 DFFPOSX1_984 ( .CLK(clk_bF_buf67), .D(_1408_), .Q(datapath_1_RegisterFile_regfile_mem_30__23_) );
DFFPOSX1 DFFPOSX1_985 ( .CLK(clk_bF_buf31), .D(_1856_), .Q(datapath_1_RegisterFile_regfile_mem_30__24_) );
DFFPOSX1 DFFPOSX1_986 ( .CLK(clk_bF_buf78), .D(_1409_), .Q(datapath_1_RegisterFile_regfile_mem_30__25_) );
DFFPOSX1 DFFPOSX1_987 ( .CLK(clk_bF_buf34), .D(_1410_), .Q(datapath_1_RegisterFile_regfile_mem_30__26_) );
DFFPOSX1 DFFPOSX1_988 ( .CLK(clk_bF_buf86), .D(_1411_), .Q(datapath_1_RegisterFile_regfile_mem_30__27_) );
DFFPOSX1 DFFPOSX1_989 ( .CLK(clk_bF_buf40), .D(_1412_), .Q(datapath_1_RegisterFile_regfile_mem_30__28_) );
DFFPOSX1 DFFPOSX1_990 ( .CLK(clk_bF_buf78), .D(_1413_), .Q(datapath_1_RegisterFile_regfile_mem_30__29_) );
DFFPOSX1 DFFPOSX1_991 ( .CLK(clk_bF_buf76), .D(_1414_), .Q(datapath_1_RegisterFile_regfile_mem_30__30_) );
DFFPOSX1 DFFPOSX1_992 ( .CLK(clk_bF_buf48), .D(_1415_), .Q(datapath_1_RegisterFile_regfile_mem_30__31_) );
DFFPOSX1 DFFPOSX1_993 ( .CLK(clk_bF_buf77), .D(_1419_), .Q(datapath_1_RegisterFile_regfile_mem_31__0_) );
DFFPOSX1 DFFPOSX1_994 ( .CLK(clk_bF_buf21), .D(_1857_), .Q(datapath_1_RegisterFile_regfile_mem_31__1_) );
DFFPOSX1 DFFPOSX1_995 ( .CLK(clk_bF_buf2), .D(_1438_), .Q(datapath_1_RegisterFile_regfile_mem_31__2_) );
DFFPOSX1 DFFPOSX1_996 ( .CLK(clk_bF_buf89), .D(_1440_), .Q(datapath_1_RegisterFile_regfile_mem_31__3_) );
DFFPOSX1 DFFPOSX1_997 ( .CLK(clk_bF_buf58), .D(_1441_), .Q(datapath_1_RegisterFile_regfile_mem_31__4_) );
DFFPOSX1 DFFPOSX1_998 ( .CLK(clk_bF_buf13), .D(_1442_), .Q(datapath_1_RegisterFile_regfile_mem_31__5_) );
DFFPOSX1 DFFPOSX1_999 ( .CLK(clk_bF_buf67), .D(_1443_), .Q(datapath_1_RegisterFile_regfile_mem_31__6_) );
DFFPOSX1 DFFPOSX1_1000 ( .CLK(clk_bF_buf98), .D(_1444_), .Q(datapath_1_RegisterFile_regfile_mem_31__7_) );
DFFPOSX1 DFFPOSX1_1001 ( .CLK(clk_bF_buf113), .D(_1445_), .Q(datapath_1_RegisterFile_regfile_mem_31__8_) );
DFFPOSX1 DFFPOSX1_1002 ( .CLK(clk_bF_buf77), .D(_1446_), .Q(datapath_1_RegisterFile_regfile_mem_31__9_) );
DFFPOSX1 DFFPOSX1_1003 ( .CLK(clk_bF_buf13), .D(_1420_), .Q(datapath_1_RegisterFile_regfile_mem_31__10_) );
DFFPOSX1 DFFPOSX1_1004 ( .CLK(clk_bF_buf98), .D(_1858_), .Q(datapath_1_RegisterFile_regfile_mem_31__11_) );
DFFPOSX1 DFFPOSX1_1005 ( .CLK(clk_bF_buf51), .D(_1421_), .Q(datapath_1_RegisterFile_regfile_mem_31__12_) );
DFFPOSX1 DFFPOSX1_1006 ( .CLK(clk_bF_buf34), .D(_1422_), .Q(datapath_1_RegisterFile_regfile_mem_31__13_) );
DFFPOSX1 DFFPOSX1_1007 ( .CLK(clk_bF_buf86), .D(_1423_), .Q(datapath_1_RegisterFile_regfile_mem_31__14_) );
DFFPOSX1 DFFPOSX1_1008 ( .CLK(clk_bF_buf3), .D(_1424_), .Q(datapath_1_RegisterFile_regfile_mem_31__15_) );
DFFPOSX1 DFFPOSX1_1009 ( .CLK(clk_bF_buf31), .D(_1425_), .Q(datapath_1_RegisterFile_regfile_mem_31__16_) );
DFFPOSX1 DFFPOSX1_1010 ( .CLK(clk_bF_buf77), .D(_1426_), .Q(datapath_1_RegisterFile_regfile_mem_31__17_) );
DFFPOSX1 DFFPOSX1_1011 ( .CLK(clk_bF_buf86), .D(_1427_), .Q(datapath_1_RegisterFile_regfile_mem_31__18_) );
DFFPOSX1 DFFPOSX1_1012 ( .CLK(clk_bF_buf51), .D(_1428_), .Q(datapath_1_RegisterFile_regfile_mem_31__19_) );
DFFPOSX1 DFFPOSX1_1013 ( .CLK(clk_bF_buf49), .D(_1429_), .Q(datapath_1_RegisterFile_regfile_mem_31__20_) );
DFFPOSX1 DFFPOSX1_1014 ( .CLK(clk_bF_buf1), .D(_1859_), .Q(datapath_1_RegisterFile_regfile_mem_31__21_) );
DFFPOSX1 DFFPOSX1_1015 ( .CLK(clk_bF_buf66), .D(_1430_), .Q(datapath_1_RegisterFile_regfile_mem_31__22_) );
DFFPOSX1 DFFPOSX1_1016 ( .CLK(clk_bF_buf58), .D(_1431_), .Q(datapath_1_RegisterFile_regfile_mem_31__23_) );
DFFPOSX1 DFFPOSX1_1017 ( .CLK(clk_bF_buf3), .D(_1432_), .Q(datapath_1_RegisterFile_regfile_mem_31__24_) );
DFFPOSX1 DFFPOSX1_1018 ( .CLK(clk_bF_buf58), .D(_1433_), .Q(datapath_1_RegisterFile_regfile_mem_31__25_) );
DFFPOSX1 DFFPOSX1_1019 ( .CLK(clk_bF_buf66), .D(_1434_), .Q(datapath_1_RegisterFile_regfile_mem_31__26_) );
DFFPOSX1 DFFPOSX1_1020 ( .CLK(clk_bF_buf86), .D(_1435_), .Q(datapath_1_RegisterFile_regfile_mem_31__27_) );
DFFPOSX1 DFFPOSX1_1021 ( .CLK(clk_bF_buf40), .D(_1436_), .Q(datapath_1_RegisterFile_regfile_mem_31__28_) );
DFFPOSX1 DFFPOSX1_1022 ( .CLK(clk_bF_buf78), .D(_1437_), .Q(datapath_1_RegisterFile_regfile_mem_31__29_) );
DFFPOSX1 DFFPOSX1_1023 ( .CLK(clk_bF_buf60), .D(_1439_), .Q(datapath_1_RegisterFile_regfile_mem_31__30_) );
DFFPOSX1 DFFPOSX1_1024 ( .CLK(clk_bF_buf86), .D(_1860_), .Q(datapath_1_RegisterFile_regfile_mem_31__31_) );
INVX1 INVX1_109 ( .A(PCSource_1_bF_buf5_), .Y(_6383_) );
NAND3X1 NAND3X1_1163 ( .A(ALUOp_0_bF_buf5_), .B(datapath_1_ALUOut_0_), .C(_6383__bF_buf0), .Y(_6384_) );
INVX1 INVX1_110 ( .A(ALUOp_0_bF_buf4_), .Y(_6385_) );
NAND3X1 NAND3X1_1164 ( .A(PCSource_1_bF_buf4_), .B(gnd), .C(_6385__bF_buf4), .Y(_6386_) );
NOR2X1 NOR2X1_142 ( .A(PCSource_1_bF_buf3_), .B(ALUOp_0_bF_buf3_), .Y(_6387_) );
AND2X2 AND2X2_1 ( .A(PCSource_1_bF_buf2_), .B(ALUOp_0_bF_buf2_), .Y(_6388_) );
AOI22X1 AOI22X1_54 ( .A(_6387__bF_buf0), .B(datapath_1_ALU_aluResult_0_), .C(gnd), .D(_6388__bF_buf3), .Y(_6389_) );
NAND3X1 NAND3X1_1165 ( .A(_6384_), .B(_6386_), .C(_6389_), .Y(datapath_1_PC_prima_0_) );
NAND3X1 NAND3X1_1166 ( .A(ALUOp_0_bF_buf1_), .B(datapath_1_ALUOut_1_), .C(_6383__bF_buf3), .Y(_6390_) );
NAND3X1 NAND3X1_1167 ( .A(PCSource_1_bF_buf1_), .B(gnd), .C(_6385__bF_buf4), .Y(_6391_) );
AOI22X1 AOI22X1_55 ( .A(_6387__bF_buf0), .B(datapath_1_ALU_aluResult_1_), .C(gnd), .D(_6388__bF_buf3), .Y(_6392_) );
NAND3X1 NAND3X1_1168 ( .A(_6390_), .B(_6391_), .C(_6392_), .Y(datapath_1_PC_prima_1_) );
NAND3X1 NAND3X1_1169 ( .A(ALUOp_0_bF_buf0_), .B(datapath_1_ALUOut_2_), .C(_6383__bF_buf0), .Y(_6393_) );
NAND3X1 NAND3X1_1170 ( .A(PCSource_1_bF_buf0_), .B(aluControl_1_inst_0_), .C(_6385__bF_buf4), .Y(_6394_) );
AOI22X1 AOI22X1_56 ( .A(_6387__bF_buf0), .B(datapath_1_ALU_aluResult_2_), .C(gnd), .D(_6388__bF_buf3), .Y(_6395_) );
NAND3X1 NAND3X1_1171 ( .A(_6393_), .B(_6394_), .C(_6395_), .Y(datapath_1_PC_prima_2_) );
NAND3X1 NAND3X1_1172 ( .A(ALUOp_0_bF_buf5_), .B(datapath_1_ALUOut_3_), .C(_6383__bF_buf4), .Y(_6396_) );
NAND3X1 NAND3X1_1173 ( .A(PCSource_1_bF_buf5_), .B(aluControl_1_inst_1_), .C(_6385__bF_buf0), .Y(_6397_) );
AOI22X1 AOI22X1_57 ( .A(_6387__bF_buf0), .B(datapath_1_ALU_aluResult_3_), .C(gnd), .D(_6388__bF_buf1), .Y(_6398_) );
NAND3X1 NAND3X1_1174 ( .A(_6396_), .B(_6397_), .C(_6398_), .Y(datapath_1_PC_prima_3_) );
NAND3X1 NAND3X1_1175 ( .A(ALUOp_0_bF_buf4_), .B(datapath_1_ALUOut_4_), .C(_6383__bF_buf3), .Y(_6399_) );
NAND3X1 NAND3X1_1176 ( .A(PCSource_1_bF_buf4_), .B(aluControl_1_inst_2_), .C(_6385__bF_buf0), .Y(_6400_) );
AOI22X1 AOI22X1_58 ( .A(_6387__bF_buf0), .B(datapath_1_ALU_aluResult_4_), .C(gnd), .D(_6388__bF_buf1), .Y(_6401_) );
NAND3X1 NAND3X1_1177 ( .A(_6399_), .B(_6400_), .C(_6401_), .Y(datapath_1_PC_prima_4_) );
NAND3X1 NAND3X1_1178 ( .A(ALUOp_0_bF_buf3_), .B(datapath_1_ALUOut_5_), .C(_6383__bF_buf3), .Y(_6402_) );
NAND3X1 NAND3X1_1179 ( .A(PCSource_1_bF_buf3_), .B(aluControl_1_inst_3_), .C(_6385__bF_buf0), .Y(_6403_) );
AOI22X1 AOI22X1_59 ( .A(_6387__bF_buf3), .B(datapath_1_ALU_aluResult_5_), .C(gnd), .D(_6388__bF_buf3), .Y(_6404_) );
NAND3X1 NAND3X1_1180 ( .A(_6402_), .B(_6403_), .C(_6404_), .Y(datapath_1_PC_prima_5_) );
NAND3X1 NAND3X1_1181 ( .A(ALUOp_0_bF_buf2_), .B(datapath_1_ALUOut_6_), .C(_6383__bF_buf0), .Y(_6405_) );
NAND3X1 NAND3X1_1182 ( .A(PCSource_1_bF_buf2_), .B(aluControl_1_inst_4_), .C(_6385__bF_buf4), .Y(_6406_) );
AOI22X1 AOI22X1_60 ( .A(_6387__bF_buf3), .B(datapath_1_ALU_aluResult_6_), .C(gnd), .D(_6388__bF_buf3), .Y(_6407_) );
NAND3X1 NAND3X1_1183 ( .A(_6405_), .B(_6406_), .C(_6407_), .Y(datapath_1_PC_prima_6_) );
NAND3X1 NAND3X1_1184 ( .A(ALUOp_0_bF_buf1_), .B(datapath_1_ALUOut_7_), .C(_6383__bF_buf3), .Y(_6408_) );
NAND3X1 NAND3X1_1185 ( .A(PCSource_1_bF_buf1_), .B(aluControl_1_inst_5_), .C(_6385__bF_buf0), .Y(_6409_) );
AOI22X1 AOI22X1_61 ( .A(_6387__bF_buf0), .B(datapath_1_ALU_aluResult_7_), .C(gnd), .D(_6388__bF_buf1), .Y(_6410_) );
NAND3X1 NAND3X1_1186 ( .A(_6408_), .B(_6409_), .C(_6410_), .Y(datapath_1_PC_prima_7_) );
NAND3X1 NAND3X1_1187 ( .A(ALUOp_0_bF_buf0_), .B(datapath_1_ALUOut_8_), .C(_6383__bF_buf2), .Y(_6411_) );
NAND3X1 NAND3X1_1188 ( .A(PCSource_1_bF_buf0_), .B(datapath_1_Instr_6_), .C(_6385__bF_buf2), .Y(_6412_) );
AOI22X1 AOI22X1_62 ( .A(_6387__bF_buf2), .B(datapath_1_ALU_aluResult_8_), .C(gnd), .D(_6388__bF_buf4), .Y(_6413_) );
NAND3X1 NAND3X1_1189 ( .A(_6411_), .B(_6412_), .C(_6413_), .Y(datapath_1_PC_prima_8_) );
NAND3X1 NAND3X1_1190 ( .A(ALUOp_0_bF_buf5_), .B(datapath_1_ALUOut_9_), .C(_6383__bF_buf1), .Y(_6414_) );
NAND3X1 NAND3X1_1191 ( .A(PCSource_1_bF_buf5_), .B(datapath_1_Instr_7_), .C(_6385__bF_buf3), .Y(_6415_) );
AOI22X1 AOI22X1_63 ( .A(_6387__bF_buf1), .B(datapath_1_ALU_aluResult_9_), .C(gnd), .D(_6388__bF_buf2), .Y(_6416_) );
NAND3X1 NAND3X1_1192 ( .A(_6414_), .B(_6415_), .C(_6416_), .Y(datapath_1_PC_prima_9_) );
NAND3X1 NAND3X1_1193 ( .A(ALUOp_0_bF_buf4_), .B(datapath_1_ALUOut_10_), .C(_6383__bF_buf1), .Y(_6417_) );
NAND3X1 NAND3X1_1194 ( .A(PCSource_1_bF_buf4_), .B(datapath_1_Instr_8_), .C(_6385__bF_buf3), .Y(_6418_) );
AOI22X1 AOI22X1_64 ( .A(_6387__bF_buf1), .B(datapath_1_ALU_aluResult_10_), .C(gnd), .D(_6388__bF_buf0), .Y(_6419_) );
NAND3X1 NAND3X1_1195 ( .A(_6417_), .B(_6418_), .C(_6419_), .Y(datapath_1_PC_prima_10_) );
NAND3X1 NAND3X1_1196 ( .A(ALUOp_0_bF_buf3_), .B(datapath_1_ALUOut_11_), .C(_6383__bF_buf4), .Y(_6420_) );
NAND3X1 NAND3X1_1197 ( .A(PCSource_1_bF_buf3_), .B(datapath_1_Instr_9_), .C(_6385__bF_buf1), .Y(_6421_) );
AOI22X1 AOI22X1_65 ( .A(_6387__bF_buf4), .B(datapath_1_ALU_aluResult_11_), .C(gnd), .D(_6388__bF_buf2), .Y(_6422_) );
NAND3X1 NAND3X1_1198 ( .A(_6420_), .B(_6421_), .C(_6422_), .Y(datapath_1_PC_prima_11_) );
NAND3X1 NAND3X1_1199 ( .A(ALUOp_0_bF_buf2_), .B(datapath_1_ALUOut_12_), .C(_6383__bF_buf4), .Y(_6423_) );
NAND3X1 NAND3X1_1200 ( .A(PCSource_1_bF_buf2_), .B(datapath_1_Instr_10_), .C(_6385__bF_buf3), .Y(_6424_) );
AOI22X1 AOI22X1_66 ( .A(_6387__bF_buf4), .B(datapath_1_ALU_aluResult_12_), .C(gnd), .D(_6388__bF_buf2), .Y(_6425_) );
NAND3X1 NAND3X1_1201 ( .A(_6423_), .B(_6424_), .C(_6425_), .Y(datapath_1_PC_prima_12_) );
NAND3X1 NAND3X1_1202 ( .A(ALUOp_0_bF_buf1_), .B(datapath_1_ALUOut_13_), .C(_6383__bF_buf1), .Y(_6426_) );
NAND3X1 NAND3X1_1203 ( .A(PCSource_1_bF_buf1_), .B(datapath_1_Instr_11_), .C(_6385__bF_buf1), .Y(_6427_) );
AOI22X1 AOI22X1_67 ( .A(_6387__bF_buf1), .B(datapath_1_ALU_aluResult_13_), .C(gnd), .D(_6388__bF_buf0), .Y(_6428_) );
NAND3X1 NAND3X1_1204 ( .A(_6426_), .B(_6427_), .C(_6428_), .Y(datapath_1_PC_prima_13_) );
NAND3X1 NAND3X1_1205 ( .A(ALUOp_0_bF_buf0_), .B(datapath_1_ALUOut_14_), .C(_6383__bF_buf2), .Y(_6429_) );
NAND3X1 NAND3X1_1206 ( .A(PCSource_1_bF_buf0_), .B(datapath_1_Instr_12_), .C(_6385__bF_buf2), .Y(_6430_) );
AOI22X1 AOI22X1_68 ( .A(_6387__bF_buf2), .B(datapath_1_ALU_aluResult_14_), .C(gnd), .D(_6388__bF_buf4), .Y(_6431_) );
NAND3X1 NAND3X1_1207 ( .A(_6429_), .B(_6430_), .C(_6431_), .Y(datapath_1_PC_prima_14_) );
NAND3X1 NAND3X1_1208 ( .A(ALUOp_0_bF_buf5_), .B(datapath_1_ALUOut_15_), .C(_6383__bF_buf2), .Y(_6432_) );
NAND3X1 NAND3X1_1209 ( .A(PCSource_1_bF_buf5_), .B(datapath_1_Instr_13_), .C(_6385__bF_buf2), .Y(_6433_) );
AOI22X1 AOI22X1_69 ( .A(_6387__bF_buf3), .B(datapath_1_ALU_aluResult_15_), .C(gnd), .D(_6388__bF_buf4), .Y(_6434_) );
NAND3X1 NAND3X1_1210 ( .A(_6432_), .B(_6433_), .C(_6434_), .Y(datapath_1_PC_prima_15_) );
NAND3X1 NAND3X1_1211 ( .A(ALUOp_0_bF_buf4_), .B(datapath_1_ALUOut_16_), .C(_6383__bF_buf4), .Y(_6435_) );
NAND3X1 NAND3X1_1212 ( .A(PCSource_1_bF_buf4_), .B(datapath_1_Instr_14_), .C(_6385__bF_buf0), .Y(_6436_) );
AOI22X1 AOI22X1_70 ( .A(_6387__bF_buf4), .B(datapath_1_ALU_aluResult_16_), .C(gnd), .D(_6388__bF_buf1), .Y(_6437_) );
NAND3X1 NAND3X1_1213 ( .A(_6435_), .B(_6436_), .C(_6437_), .Y(datapath_1_PC_prima_16_) );
NAND3X1 NAND3X1_1214 ( .A(ALUOp_0_bF_buf3_), .B(datapath_1_ALUOut_17_), .C(_6383__bF_buf4), .Y(_6438_) );
NAND3X1 NAND3X1_1215 ( .A(PCSource_1_bF_buf3_), .B(datapath_1_Instr_15_bF_buf4_), .C(_6385__bF_buf1), .Y(_6439_) );
AOI22X1 AOI22X1_71 ( .A(_6387__bF_buf4), .B(datapath_1_ALU_aluResult_17_), .C(gnd), .D(_6388__bF_buf1), .Y(_6440_) );
NAND3X1 NAND3X1_1216 ( .A(_6438_), .B(_6439_), .C(_6440_), .Y(datapath_1_PC_prima_17_) );
NAND3X1 NAND3X1_1217 ( .A(ALUOp_0_bF_buf2_), .B(datapath_1_ALUOut_18_), .C(_6383__bF_buf0), .Y(_6441_) );
NAND3X1 NAND3X1_1218 ( .A(PCSource_1_bF_buf2_), .B(datapath_1_Instr_16_bF_buf50_), .C(_6385__bF_buf3), .Y(_6442_) );
AOI22X1 AOI22X1_72 ( .A(_6387__bF_buf3), .B(datapath_1_ALU_aluResult_18_), .C(gnd), .D(_6388__bF_buf4), .Y(_6443_) );
NAND3X1 NAND3X1_1219 ( .A(_6441_), .B(_6442_), .C(_6443_), .Y(datapath_1_PC_prima_18_) );
NAND3X1 NAND3X1_1220 ( .A(ALUOp_0_bF_buf1_), .B(datapath_1_ALUOut_19_), .C(_6383__bF_buf3), .Y(_6444_) );
NAND3X1 NAND3X1_1221 ( .A(PCSource_1_bF_buf1_), .B(datapath_1_Instr_17_bF_buf10_), .C(_6385__bF_buf1), .Y(_6445_) );
AOI22X1 AOI22X1_73 ( .A(_6387__bF_buf1), .B(datapath_1_ALU_aluResult_19_), .C(gnd), .D(_6388__bF_buf2), .Y(_6446_) );
NAND3X1 NAND3X1_1222 ( .A(_6444_), .B(_6445_), .C(_6446_), .Y(datapath_1_PC_prima_19_) );
NAND3X1 NAND3X1_1223 ( .A(ALUOp_0_bF_buf0_), .B(datapath_1_ALUOut_20_), .C(_6383__bF_buf0), .Y(_6447_) );
NAND3X1 NAND3X1_1224 ( .A(PCSource_1_bF_buf0_), .B(datapath_1_Instr_18_bF_buf3_), .C(_6385__bF_buf2), .Y(_6448_) );
AOI22X1 AOI22X1_74 ( .A(_6387__bF_buf3), .B(datapath_1_ALU_aluResult_20_), .C(gnd), .D(_6388__bF_buf4), .Y(_6449_) );
NAND3X1 NAND3X1_1225 ( .A(_6447_), .B(_6448_), .C(_6449_), .Y(datapath_1_PC_prima_20_) );
NAND3X1 NAND3X1_1226 ( .A(ALUOp_0_bF_buf5_), .B(datapath_1_ALUOut_21_), .C(_6383__bF_buf0), .Y(_6450_) );
NAND3X1 NAND3X1_1227 ( .A(PCSource_1_bF_buf5_), .B(datapath_1_Instr_19_bF_buf6_), .C(_6385__bF_buf4), .Y(_6451_) );
AOI22X1 AOI22X1_75 ( .A(_6387__bF_buf3), .B(datapath_1_ALU_aluResult_21_), .C(gnd), .D(_6388__bF_buf3), .Y(_6452_) );
NAND3X1 NAND3X1_1228 ( .A(_6450_), .B(_6451_), .C(_6452_), .Y(datapath_1_PC_prima_21_) );
NAND3X1 NAND3X1_1229 ( .A(ALUOp_0_bF_buf4_), .B(datapath_1_ALUOut_22_), .C(_6383__bF_buf3), .Y(_6453_) );
NAND3X1 NAND3X1_1230 ( .A(PCSource_1_bF_buf4_), .B(datapath_1_Instr_20_bF_buf5_), .C(_6385__bF_buf0), .Y(_6454_) );
AOI22X1 AOI22X1_76 ( .A(_6387__bF_buf4), .B(datapath_1_ALU_aluResult_22_), .C(gnd), .D(_6388__bF_buf1), .Y(_6455_) );
NAND3X1 NAND3X1_1231 ( .A(_6453_), .B(_6454_), .C(_6455_), .Y(datapath_1_PC_prima_22_) );
NAND3X1 NAND3X1_1232 ( .A(ALUOp_0_bF_buf3_), .B(datapath_1_ALUOut_23_), .C(_6383__bF_buf4), .Y(_6456_) );
NAND3X1 NAND3X1_1233 ( .A(PCSource_1_bF_buf3_), .B(datapath_1_Instr_21_bF_buf55_), .C(_6385__bF_buf1), .Y(_6457_) );
AOI22X1 AOI22X1_77 ( .A(_6387__bF_buf4), .B(datapath_1_ALU_aluResult_23_), .C(gnd), .D(_6388__bF_buf2), .Y(_6458_) );
NAND3X1 NAND3X1_1234 ( .A(_6456_), .B(_6457_), .C(_6458_), .Y(datapath_1_PC_prima_23_) );
NAND3X1 NAND3X1_1235 ( .A(ALUOp_0_bF_buf2_), .B(datapath_1_ALUOut_24_), .C(_6383__bF_buf2), .Y(_6459_) );
NAND3X1 NAND3X1_1236 ( .A(PCSource_1_bF_buf2_), .B(datapath_1_Instr_22_bF_buf50_), .C(_6385__bF_buf2), .Y(_6460_) );
AOI22X1 AOI22X1_78 ( .A(_6387__bF_buf2), .B(datapath_1_ALU_aluResult_24_), .C(gnd), .D(_6388__bF_buf4), .Y(_6461_) );
NAND3X1 NAND3X1_1237 ( .A(_6459_), .B(_6460_), .C(_6461_), .Y(datapath_1_PC_prima_24_) );
NAND3X1 NAND3X1_1238 ( .A(ALUOp_0_bF_buf1_), .B(datapath_1_ALUOut_25_), .C(_6383__bF_buf3), .Y(_6462_) );
NAND3X1 NAND3X1_1239 ( .A(PCSource_1_bF_buf1_), .B(datapath_1_Instr_23_bF_buf15_bF_buf3_), .C(_6385__bF_buf4), .Y(_6463_) );
AOI22X1 AOI22X1_79 ( .A(_6387__bF_buf3), .B(datapath_1_ALU_aluResult_25_), .C(gnd), .D(_6388__bF_buf3), .Y(_6464_) );
NAND3X1 NAND3X1_1240 ( .A(_6462_), .B(_6463_), .C(_6464_), .Y(datapath_1_PC_prima_25_) );
NAND3X1 NAND3X1_1241 ( .A(ALUOp_0_bF_buf0_), .B(datapath_1_ALUOut_26_), .C(_6383__bF_buf2), .Y(_6465_) );
NAND3X1 NAND3X1_1242 ( .A(PCSource_1_bF_buf0_), .B(datapath_1_Instr_24_bF_buf6_), .C(_6385__bF_buf4), .Y(_6466_) );
AOI22X1 AOI22X1_80 ( .A(_6387__bF_buf2), .B(datapath_1_ALU_aluResult_26_), .C(gnd), .D(_6388__bF_buf0), .Y(_6467_) );
NAND3X1 NAND3X1_1243 ( .A(_6465_), .B(_6466_), .C(_6467_), .Y(datapath_1_PC_prima_26_) );
NAND3X1 NAND3X1_1244 ( .A(ALUOp_0_bF_buf5_), .B(datapath_1_ALUOut_27_), .C(_6383__bF_buf2), .Y(_6468_) );
NAND3X1 NAND3X1_1245 ( .A(PCSource_1_bF_buf5_), .B(datapath_1_Instr_25_bF_buf5_), .C(_6385__bF_buf2), .Y(_6469_) );
AOI22X1 AOI22X1_81 ( .A(_6387__bF_buf2), .B(datapath_1_ALU_aluResult_27_), .C(gnd), .D(_6388__bF_buf4), .Y(_6470_) );
NAND3X1 NAND3X1_1246 ( .A(_6468_), .B(_6469_), .C(_6470_), .Y(datapath_1_PC_prima_27_) );
NAND3X1 NAND3X1_1247 ( .A(ALUOp_0_bF_buf4_), .B(datapath_1_ALUOut_28_), .C(_6383__bF_buf1), .Y(_6471_) );
NAND3X1 NAND3X1_1248 ( .A(PCSource_1_bF_buf4_), .B(datapath_1_PC_28_), .C(_6385__bF_buf3), .Y(_6472_) );
AOI22X1 AOI22X1_82 ( .A(_6387__bF_buf2), .B(datapath_1_ALU_aluResult_28_), .C(gnd), .D(_6388__bF_buf0), .Y(_6473_) );
NAND3X1 NAND3X1_1249 ( .A(_6471_), .B(_6472_), .C(_6473_), .Y(datapath_1_PC_prima_28_) );
NAND3X1 NAND3X1_1250 ( .A(ALUOp_0_bF_buf3_), .B(datapath_1_ALUOut_29_), .C(_6383__bF_buf4), .Y(_6474_) );
NAND3X1 NAND3X1_1251 ( .A(PCSource_1_bF_buf3_), .B(datapath_1_PC_29_), .C(_6385__bF_buf1), .Y(_6475_) );
AOI22X1 AOI22X1_83 ( .A(_6387__bF_buf4), .B(datapath_1_ALU_aluResult_29_), .C(gnd), .D(_6388__bF_buf2), .Y(_6476_) );
NAND3X1 NAND3X1_1252 ( .A(_6474_), .B(_6475_), .C(_6476_), .Y(datapath_1_PC_prima_29_) );
NAND3X1 NAND3X1_1253 ( .A(ALUOp_0_bF_buf2_), .B(datapath_1_ALUOut_30_), .C(_6383__bF_buf1), .Y(_6477_) );
NAND3X1 NAND3X1_1254 ( .A(PCSource_1_bF_buf2_), .B(datapath_1_PC_30_), .C(_6385__bF_buf3), .Y(_6478_) );
AOI22X1 AOI22X1_84 ( .A(_6387__bF_buf1), .B(datapath_1_ALU_aluResult_30_), .C(gnd), .D(_6388__bF_buf0), .Y(_6479_) );
NAND3X1 NAND3X1_1255 ( .A(_6477_), .B(_6478_), .C(_6479_), .Y(datapath_1_PC_prima_30_) );
NAND3X1 NAND3X1_1256 ( .A(ALUOp_0_bF_buf1_), .B(datapath_1_ALUOut_31_), .C(_6383__bF_buf1), .Y(_6480_) );
NAND3X1 NAND3X1_1257 ( .A(PCSource_1_bF_buf1_), .B(datapath_1_PC_31_), .C(_6385__bF_buf3), .Y(_6481_) );
AOI22X1 AOI22X1_85 ( .A(_6387__bF_buf1), .B(datapath_1_ALU_aluResult_31_), .C(gnd), .D(_6388__bF_buf0), .Y(_6482_) );
NAND3X1 NAND3X1_1258 ( .A(_6480_), .B(_6481_), .C(_6482_), .Y(datapath_1_PC_prima_31_) );
INVX1 INVX1_111 ( .A(datapath_1_PC_0_), .Y(_6545_) );
NAND2X1 NAND2X1_424 ( .A(datapath_1_A_0_), .B(ALUSrcA_bF_buf4), .Y(_6546_) );
OAI21X1 OAI21X1_1317 ( .A(ALUSrcA_bF_buf4), .B(_6545_), .C(_6546_), .Y(datapath_1_ALU_aluInA_0_) );
INVX1 INVX1_112 ( .A(datapath_1_PC_1_), .Y(_6483_) );
NAND2X1 NAND2X1_425 ( .A(ALUSrcA_bF_buf2), .B(datapath_1_A_1_), .Y(_6484_) );
OAI21X1 OAI21X1_1318 ( .A(ALUSrcA_bF_buf2), .B(_6483_), .C(_6484_), .Y(datapath_1_ALU_aluInA_1_) );
INVX1 INVX1_113 ( .A(datapath_1_PC_2_), .Y(_6485_) );
NAND2X1 NAND2X1_426 ( .A(ALUSrcA_bF_buf2), .B(datapath_1_A_2_), .Y(_6486_) );
OAI21X1 OAI21X1_1319 ( .A(ALUSrcA_bF_buf2), .B(_6485_), .C(_6486_), .Y(datapath_1_ALU_aluInA_2_) );
INVX1 INVX1_114 ( .A(datapath_1_PC_3_), .Y(_6487_) );
NAND2X1 NAND2X1_427 ( .A(ALUSrcA_bF_buf1), .B(datapath_1_A_3_), .Y(_6488_) );
OAI21X1 OAI21X1_1320 ( .A(ALUSrcA_bF_buf0), .B(_6487_), .C(_6488_), .Y(datapath_1_ALU_aluInA_3_) );
INVX1 INVX1_115 ( .A(datapath_1_PC_4_), .Y(_6489_) );
NAND2X1 NAND2X1_428 ( .A(ALUSrcA_bF_buf4), .B(datapath_1_A_4_), .Y(_6490_) );
OAI21X1 OAI21X1_1321 ( .A(ALUSrcA_bF_buf4), .B(_6489_), .C(_6490_), .Y(datapath_1_ALU_aluInA_4_) );
INVX1 INVX1_116 ( .A(datapath_1_PC_5_), .Y(_6491_) );
NAND2X1 NAND2X1_429 ( .A(ALUSrcA_bF_buf4), .B(datapath_1_A_5_), .Y(_6492_) );
OAI21X1 OAI21X1_1322 ( .A(ALUSrcA_bF_buf4), .B(_6491_), .C(_6492_), .Y(datapath_1_ALU_aluInA_5_) );
INVX1 INVX1_117 ( .A(datapath_1_PC_6_), .Y(_6493_) );
NAND2X1 NAND2X1_430 ( .A(ALUSrcA_bF_buf5), .B(datapath_1_A_6_), .Y(_6494_) );
OAI21X1 OAI21X1_1323 ( .A(ALUSrcA_bF_buf2), .B(_6493_), .C(_6494_), .Y(datapath_1_ALU_aluInA_6_) );
INVX1 INVX1_118 ( .A(datapath_1_PC_7_), .Y(_6495_) );
NAND2X1 NAND2X1_431 ( .A(ALUSrcA_bF_buf1), .B(datapath_1_A_7_), .Y(_6496_) );
OAI21X1 OAI21X1_1324 ( .A(ALUSrcA_bF_buf1), .B(_6495_), .C(_6496_), .Y(datapath_1_ALU_aluInA_7_) );
INVX1 INVX1_119 ( .A(datapath_1_PC_8_), .Y(_6497_) );
NAND2X1 NAND2X1_432 ( .A(ALUSrcA_bF_buf3), .B(datapath_1_A_8_), .Y(_6498_) );
OAI21X1 OAI21X1_1325 ( .A(ALUSrcA_bF_buf3), .B(_6497_), .C(_6498_), .Y(datapath_1_ALU_aluInA_8_) );
INVX1 INVX1_120 ( .A(datapath_1_PC_9_), .Y(_6499_) );
NAND2X1 NAND2X1_433 ( .A(ALUSrcA_bF_buf7), .B(datapath_1_A_9_), .Y(_6500_) );
OAI21X1 OAI21X1_1326 ( .A(ALUSrcA_bF_buf7), .B(_6499_), .C(_6500_), .Y(datapath_1_ALU_aluInA_9_) );
INVX1 INVX1_121 ( .A(datapath_1_PC_10_), .Y(_6501_) );
NAND2X1 NAND2X1_434 ( .A(ALUSrcA_bF_buf7), .B(datapath_1_A_10_), .Y(_6502_) );
OAI21X1 OAI21X1_1327 ( .A(ALUSrcA_bF_buf7), .B(_6501_), .C(_6502_), .Y(datapath_1_ALU_aluInA_10_) );
INVX1 INVX1_122 ( .A(datapath_1_PC_11_), .Y(_6503_) );
NAND2X1 NAND2X1_435 ( .A(ALUSrcA_bF_buf1), .B(datapath_1_A_11_), .Y(_6504_) );
OAI21X1 OAI21X1_1328 ( .A(ALUSrcA_bF_buf6), .B(_6503_), .C(_6504_), .Y(datapath_1_ALU_aluInA_11_) );
INVX1 INVX1_123 ( .A(datapath_1_PC_12_), .Y(_6505_) );
NAND2X1 NAND2X1_436 ( .A(ALUSrcA_bF_buf0), .B(datapath_1_A_12_), .Y(_6506_) );
OAI21X1 OAI21X1_1329 ( .A(ALUSrcA_bF_buf3), .B(_6505_), .C(_6506_), .Y(datapath_1_ALU_aluInA_12_) );
INVX1 INVX1_124 ( .A(datapath_1_PC_13_), .Y(_6507_) );
NAND2X1 NAND2X1_437 ( .A(ALUSrcA_bF_buf5), .B(datapath_1_A_13_), .Y(_6508_) );
OAI21X1 OAI21X1_1330 ( .A(ALUSrcA_bF_buf3), .B(_6507_), .C(_6508_), .Y(datapath_1_ALU_aluInA_13_) );
INVX1 INVX1_125 ( .A(datapath_1_PC_14_), .Y(_6509_) );
NAND2X1 NAND2X1_438 ( .A(ALUSrcA_bF_buf3), .B(datapath_1_A_14_), .Y(_6510_) );
OAI21X1 OAI21X1_1331 ( .A(ALUSrcA_bF_buf7), .B(_6509_), .C(_6510_), .Y(datapath_1_ALU_aluInA_14_) );
INVX1 INVX1_126 ( .A(datapath_1_PC_15_), .Y(_6511_) );
NAND2X1 NAND2X1_439 ( .A(ALUSrcA_bF_buf0), .B(datapath_1_A_15_), .Y(_6512_) );
OAI21X1 OAI21X1_1332 ( .A(ALUSrcA_bF_buf3), .B(_6511_), .C(_6512_), .Y(datapath_1_ALU_aluInA_15_) );
INVX1 INVX1_127 ( .A(datapath_1_PC_16_), .Y(_6513_) );
NAND2X1 NAND2X1_440 ( .A(ALUSrcA_bF_buf1), .B(datapath_1_A_16_), .Y(_6514_) );
OAI21X1 OAI21X1_1333 ( .A(ALUSrcA_bF_buf0), .B(_6513_), .C(_6514_), .Y(datapath_1_ALU_aluInA_16_) );
INVX1 INVX1_128 ( .A(datapath_1_PC_17_), .Y(_6515_) );
NAND2X1 NAND2X1_441 ( .A(ALUSrcA_bF_buf2), .B(datapath_1_A_17_), .Y(_6516_) );
OAI21X1 OAI21X1_1334 ( .A(ALUSrcA_bF_buf0), .B(_6515_), .C(_6516_), .Y(datapath_1_ALU_aluInA_17_) );
INVX1 INVX1_129 ( .A(datapath_1_PC_18_), .Y(_6517_) );
NAND2X1 NAND2X1_442 ( .A(ALUSrcA_bF_buf4), .B(datapath_1_A_18_), .Y(_6518_) );
OAI21X1 OAI21X1_1335 ( .A(ALUSrcA_bF_buf5), .B(_6517_), .C(_6518_), .Y(datapath_1_ALU_aluInA_18_) );
INVX1 INVX1_130 ( .A(datapath_1_PC_19_), .Y(_6519_) );
NAND2X1 NAND2X1_443 ( .A(ALUSrcA_bF_buf1), .B(datapath_1_A_19_), .Y(_6520_) );
OAI21X1 OAI21X1_1336 ( .A(ALUSrcA_bF_buf0), .B(_6519_), .C(_6520_), .Y(datapath_1_ALU_aluInA_19_) );
INVX1 INVX1_131 ( .A(datapath_1_PC_20_), .Y(_6521_) );
NAND2X1 NAND2X1_444 ( .A(ALUSrcA_bF_buf0), .B(datapath_1_A_20_), .Y(_6522_) );
OAI21X1 OAI21X1_1337 ( .A(ALUSrcA_bF_buf0), .B(_6521_), .C(_6522_), .Y(datapath_1_ALU_aluInA_20_) );
INVX1 INVX1_132 ( .A(datapath_1_PC_21_), .Y(_6523_) );
NAND2X1 NAND2X1_445 ( .A(ALUSrcA_bF_buf5), .B(datapath_1_A_21_), .Y(_6524_) );
OAI21X1 OAI21X1_1338 ( .A(ALUSrcA_bF_buf5), .B(_6523_), .C(_6524_), .Y(datapath_1_ALU_aluInA_21_) );
INVX1 INVX1_133 ( .A(datapath_1_PC_22_), .Y(_6525_) );
NAND2X1 NAND2X1_446 ( .A(ALUSrcA_bF_buf5), .B(datapath_1_A_22_), .Y(_6526_) );
OAI21X1 OAI21X1_1339 ( .A(ALUSrcA_bF_buf3), .B(_6525_), .C(_6526_), .Y(datapath_1_ALU_aluInA_22_) );
INVX1 INVX1_134 ( .A(datapath_1_PC_23_), .Y(_6527_) );
NAND2X1 NAND2X1_447 ( .A(ALUSrcA_bF_buf2), .B(datapath_1_A_23_), .Y(_6528_) );
OAI21X1 OAI21X1_1340 ( .A(ALUSrcA_bF_buf6), .B(_6527_), .C(_6528_), .Y(datapath_1_ALU_aluInA_23_) );
INVX1 INVX1_135 ( .A(datapath_1_PC_24_), .Y(_6529_) );
NAND2X1 NAND2X1_448 ( .A(ALUSrcA_bF_buf6), .B(datapath_1_A_24_), .Y(_6530_) );
OAI21X1 OAI21X1_1341 ( .A(ALUSrcA_bF_buf6), .B(_6529_), .C(_6530_), .Y(datapath_1_ALU_aluInA_24_) );
INVX1 INVX1_136 ( .A(datapath_1_PC_25_), .Y(_6531_) );
NAND2X1 NAND2X1_449 ( .A(ALUSrcA_bF_buf1), .B(datapath_1_A_25_), .Y(_6532_) );
OAI21X1 OAI21X1_1342 ( .A(ALUSrcA_bF_buf1), .B(_6531_), .C(_6532_), .Y(datapath_1_ALU_aluInA_25_) );
INVX1 INVX1_137 ( .A(datapath_1_PC_26_), .Y(_6533_) );
NAND2X1 NAND2X1_450 ( .A(ALUSrcA_bF_buf5), .B(datapath_1_A_26_), .Y(_6534_) );
OAI21X1 OAI21X1_1343 ( .A(ALUSrcA_bF_buf7), .B(_6533_), .C(_6534_), .Y(datapath_1_ALU_aluInA_26_) );
INVX1 INVX1_138 ( .A(datapath_1_PC_27_), .Y(_6535_) );
NAND2X1 NAND2X1_451 ( .A(ALUSrcA_bF_buf2), .B(datapath_1_A_27_), .Y(_6536_) );
OAI21X1 OAI21X1_1344 ( .A(ALUSrcA_bF_buf3), .B(_6535_), .C(_6536_), .Y(datapath_1_ALU_aluInA_27_) );
INVX1 INVX1_139 ( .A(datapath_1_PC_28_), .Y(_6537_) );
NAND2X1 NAND2X1_452 ( .A(ALUSrcA_bF_buf6), .B(datapath_1_A_28_), .Y(_6538_) );
OAI21X1 OAI21X1_1345 ( .A(ALUSrcA_bF_buf6), .B(_6537_), .C(_6538_), .Y(datapath_1_ALU_aluInA_28_) );
INVX1 INVX1_140 ( .A(datapath_1_PC_29_), .Y(_6539_) );
NAND2X1 NAND2X1_453 ( .A(ALUSrcA_bF_buf6), .B(datapath_1_A_29_), .Y(_6540_) );
OAI21X1 OAI21X1_1346 ( .A(ALUSrcA_bF_buf6), .B(_6539_), .C(_6540_), .Y(datapath_1_ALU_aluInA_29_) );
INVX1 INVX1_141 ( .A(datapath_1_PC_30_), .Y(_6541_) );
NAND2X1 NAND2X1_454 ( .A(ALUSrcA_bF_buf5), .B(datapath_1_A_30_), .Y(_6542_) );
OAI21X1 OAI21X1_1347 ( .A(ALUSrcA_bF_buf7), .B(_6541_), .C(_6542_), .Y(datapath_1_ALU_aluInA_30_) );
INVX1 INVX1_142 ( .A(datapath_1_PC_31_), .Y(_6543_) );
NAND2X1 NAND2X1_455 ( .A(ALUSrcA_bF_buf4), .B(datapath_1_A_31_), .Y(_6544_) );
OAI21X1 OAI21X1_1348 ( .A(ALUSrcA_bF_buf7), .B(_6543_), .C(_6544_), .Y(datapath_1_ALU_aluInA_31_) );
INVX1 INVX1_143 ( .A(ALUSrcB_1_bF_buf4_), .Y(_6547_) );
NAND3X1 NAND3X1_1259 ( .A(ALUSrcB_0_bF_buf4_), .B(gnd), .C(_6547__bF_buf4), .Y(_6548_) );
INVX1 INVX1_144 ( .A(ALUSrcB_0_bF_buf3_), .Y(_6549_) );
NAND3X1 NAND3X1_1260 ( .A(ALUSrcB_1_bF_buf3_), .B(aluControl_1_inst_0_), .C(_6549__bF_buf1), .Y(_6550_) );
NOR2X1 NOR2X1_143 ( .A(ALUSrcB_1_bF_buf2_), .B(ALUSrcB_0_bF_buf2_), .Y(_6551_) );
AND2X2 AND2X2_2 ( .A(ALUSrcB_1_bF_buf1_), .B(ALUSrcB_0_bF_buf1_), .Y(_6552_) );
AOI22X1 AOI22X1_86 ( .A(_6551__bF_buf3), .B(_2__0_), .C(gnd), .D(_6552__bF_buf0), .Y(_6553_) );
NAND3X1 NAND3X1_1261 ( .A(_6548_), .B(_6550_), .C(_6553_), .Y(datapath_1_ALU_aluInB_0_) );
NAND3X1 NAND3X1_1262 ( .A(ALUSrcB_0_bF_buf0_), .B(gnd), .C(_6547__bF_buf4), .Y(_6554_) );
NAND3X1 NAND3X1_1263 ( .A(ALUSrcB_1_bF_buf0_), .B(aluControl_1_inst_1_), .C(_6549__bF_buf1), .Y(_6555_) );
AOI22X1 AOI22X1_87 ( .A(_6551__bF_buf3), .B(_2__1_), .C(gnd), .D(_6552__bF_buf0), .Y(_6556_) );
NAND3X1 NAND3X1_1264 ( .A(_6554_), .B(_6555_), .C(_6556_), .Y(datapath_1_ALU_aluInB_1_) );
NAND3X1 NAND3X1_1265 ( .A(ALUSrcB_0_bF_buf4_), .B(vdd), .C(_6547__bF_buf4), .Y(_6557_) );
NAND3X1 NAND3X1_1266 ( .A(ALUSrcB_1_bF_buf4_), .B(aluControl_1_inst_2_), .C(_6549__bF_buf4), .Y(_6558_) );
AOI22X1 AOI22X1_88 ( .A(_6551__bF_buf3), .B(_2__2_), .C(aluControl_1_inst_0_), .D(_6552__bF_buf0), .Y(_6559_) );
NAND3X1 NAND3X1_1267 ( .A(_6557_), .B(_6558_), .C(_6559_), .Y(datapath_1_ALU_aluInB_2_) );
NAND3X1 NAND3X1_1268 ( .A(ALUSrcB_0_bF_buf3_), .B(gnd), .C(_6547__bF_buf0), .Y(_6560_) );
NAND3X1 NAND3X1_1269 ( .A(ALUSrcB_1_bF_buf3_), .B(aluControl_1_inst_3_), .C(_6549__bF_buf4), .Y(_6561_) );
AOI22X1 AOI22X1_89 ( .A(_6551__bF_buf3), .B(_2__3_), .C(aluControl_1_inst_1_), .D(_6552__bF_buf0), .Y(_6562_) );
NAND3X1 NAND3X1_1270 ( .A(_6560_), .B(_6561_), .C(_6562_), .Y(datapath_1_ALU_aluInB_3_) );
NAND3X1 NAND3X1_1271 ( .A(ALUSrcB_0_bF_buf2_), .B(gnd), .C(_6547__bF_buf0), .Y(_6563_) );
NAND3X1 NAND3X1_1272 ( .A(ALUSrcB_1_bF_buf2_), .B(aluControl_1_inst_4_), .C(_6549__bF_buf4), .Y(_6564_) );
AOI22X1 AOI22X1_90 ( .A(_6551__bF_buf2), .B(_2__4_), .C(aluControl_1_inst_2_), .D(_6552__bF_buf1), .Y(_6565_) );
NAND3X1 NAND3X1_1273 ( .A(_6563_), .B(_6564_), .C(_6565_), .Y(datapath_1_ALU_aluInB_4_) );
NAND3X1 NAND3X1_1274 ( .A(ALUSrcB_0_bF_buf1_), .B(gnd), .C(_6547__bF_buf4), .Y(_6566_) );
NAND3X1 NAND3X1_1275 ( .A(ALUSrcB_1_bF_buf1_), .B(aluControl_1_inst_5_), .C(_6549__bF_buf1), .Y(_6567_) );
AOI22X1 AOI22X1_91 ( .A(_6551__bF_buf2), .B(_2__5_), .C(aluControl_1_inst_3_), .D(_6552__bF_buf1), .Y(_6568_) );
NAND3X1 NAND3X1_1276 ( .A(_6566_), .B(_6567_), .C(_6568_), .Y(datapath_1_ALU_aluInB_5_) );
NAND3X1 NAND3X1_1277 ( .A(ALUSrcB_0_bF_buf0_), .B(gnd), .C(_6547__bF_buf0), .Y(_6569_) );
NAND3X1 NAND3X1_1278 ( .A(ALUSrcB_1_bF_buf0_), .B(datapath_1_Instr_6_), .C(_6549__bF_buf4), .Y(_6570_) );
AOI22X1 AOI22X1_92 ( .A(_6551__bF_buf2), .B(_2__6_), .C(aluControl_1_inst_4_), .D(_6552__bF_buf1), .Y(_6571_) );
NAND3X1 NAND3X1_1279 ( .A(_6569_), .B(_6570_), .C(_6571_), .Y(datapath_1_ALU_aluInB_6_) );
NAND3X1 NAND3X1_1280 ( .A(ALUSrcB_0_bF_buf4_), .B(gnd), .C(_6547__bF_buf4), .Y(_6572_) );
NAND3X1 NAND3X1_1281 ( .A(ALUSrcB_1_bF_buf4_), .B(datapath_1_Instr_7_), .C(_6549__bF_buf1), .Y(_6573_) );
AOI22X1 AOI22X1_93 ( .A(_6551__bF_buf4), .B(_2__7_), .C(aluControl_1_inst_5_), .D(_6552__bF_buf4), .Y(_6574_) );
NAND3X1 NAND3X1_1282 ( .A(_6572_), .B(_6573_), .C(_6574_), .Y(datapath_1_ALU_aluInB_7_) );
NAND3X1 NAND3X1_1283 ( .A(ALUSrcB_0_bF_buf3_), .B(gnd), .C(_6547__bF_buf2), .Y(_6575_) );
NAND3X1 NAND3X1_1284 ( .A(ALUSrcB_1_bF_buf3_), .B(datapath_1_Instr_8_), .C(_6549__bF_buf3), .Y(_6576_) );
AOI22X1 AOI22X1_94 ( .A(_6551__bF_buf0), .B(_2__8_), .C(datapath_1_Instr_6_), .D(_6552__bF_buf2), .Y(_6577_) );
NAND3X1 NAND3X1_1285 ( .A(_6575_), .B(_6576_), .C(_6577_), .Y(datapath_1_ALU_aluInB_8_) );
NAND3X1 NAND3X1_1286 ( .A(ALUSrcB_0_bF_buf2_), .B(gnd), .C(_6547__bF_buf0), .Y(_6578_) );
NAND3X1 NAND3X1_1287 ( .A(ALUSrcB_1_bF_buf2_), .B(datapath_1_Instr_9_), .C(_6549__bF_buf4), .Y(_6579_) );
AOI22X1 AOI22X1_95 ( .A(_6551__bF_buf3), .B(_2__9_), .C(datapath_1_Instr_7_), .D(_6552__bF_buf3), .Y(_6580_) );
NAND3X1 NAND3X1_1288 ( .A(_6578_), .B(_6579_), .C(_6580_), .Y(datapath_1_ALU_aluInB_9_) );
NAND3X1 NAND3X1_1289 ( .A(ALUSrcB_0_bF_buf1_), .B(gnd), .C(_6547__bF_buf2), .Y(_6581_) );
NAND3X1 NAND3X1_1290 ( .A(ALUSrcB_1_bF_buf1_), .B(datapath_1_Instr_10_), .C(_6549__bF_buf3), .Y(_6582_) );
AOI22X1 AOI22X1_96 ( .A(_6551__bF_buf0), .B(_2__10_), .C(datapath_1_Instr_8_), .D(_6552__bF_buf2), .Y(_6583_) );
NAND3X1 NAND3X1_1291 ( .A(_6581_), .B(_6582_), .C(_6583_), .Y(datapath_1_ALU_aluInB_10_) );
NAND3X1 NAND3X1_1292 ( .A(ALUSrcB_0_bF_buf0_), .B(gnd), .C(_6547__bF_buf3), .Y(_6584_) );
NAND3X1 NAND3X1_1293 ( .A(ALUSrcB_1_bF_buf0_), .B(datapath_1_Instr_11_), .C(_6549__bF_buf3), .Y(_6585_) );
AOI22X1 AOI22X1_97 ( .A(_6551__bF_buf1), .B(_2__11_), .C(datapath_1_Instr_9_), .D(_6552__bF_buf3), .Y(_6586_) );
NAND3X1 NAND3X1_1294 ( .A(_6584_), .B(_6585_), .C(_6586_), .Y(datapath_1_ALU_aluInB_11_) );
NAND3X1 NAND3X1_1295 ( .A(ALUSrcB_0_bF_buf4_), .B(gnd), .C(_6547__bF_buf2), .Y(_6587_) );
NAND3X1 NAND3X1_1296 ( .A(ALUSrcB_1_bF_buf4_), .B(datapath_1_Instr_12_), .C(_6549__bF_buf3), .Y(_6588_) );
AOI22X1 AOI22X1_98 ( .A(_6551__bF_buf1), .B(_2__12_), .C(datapath_1_Instr_10_), .D(_6552__bF_buf3), .Y(_6589_) );
NAND3X1 NAND3X1_1297 ( .A(_6587_), .B(_6588_), .C(_6589_), .Y(datapath_1_ALU_aluInB_12_) );
NAND3X1 NAND3X1_1298 ( .A(ALUSrcB_0_bF_buf3_), .B(gnd), .C(_6547__bF_buf2), .Y(_6590_) );
NAND3X1 NAND3X1_1299 ( .A(ALUSrcB_1_bF_buf3_), .B(datapath_1_Instr_13_), .C(_6549__bF_buf3), .Y(_6591_) );
AOI22X1 AOI22X1_99 ( .A(_6551__bF_buf0), .B(_2__13_), .C(datapath_1_Instr_11_), .D(_6552__bF_buf2), .Y(_6592_) );
NAND3X1 NAND3X1_1300 ( .A(_6590_), .B(_6591_), .C(_6592_), .Y(datapath_1_ALU_aluInB_13_) );
NAND3X1 NAND3X1_1301 ( .A(ALUSrcB_0_bF_buf2_), .B(gnd), .C(_6547__bF_buf0), .Y(_6593_) );
NAND3X1 NAND3X1_1302 ( .A(ALUSrcB_1_bF_buf2_), .B(datapath_1_Instr_14_), .C(_6549__bF_buf3), .Y(_6594_) );
AOI22X1 AOI22X1_100 ( .A(_6551__bF_buf2), .B(_2__14_), .C(datapath_1_Instr_12_), .D(_6552__bF_buf1), .Y(_6595_) );
NAND3X1 NAND3X1_1303 ( .A(_6593_), .B(_6594_), .C(_6595_), .Y(datapath_1_ALU_aluInB_14_) );
NAND3X1 NAND3X1_1304 ( .A(ALUSrcB_0_bF_buf1_), .B(gnd), .C(_6547__bF_buf0), .Y(_6596_) );
NAND3X1 NAND3X1_1305 ( .A(ALUSrcB_1_bF_buf1_), .B(datapath_1_Instr_15_bF_buf3_), .C(_6549__bF_buf4), .Y(_6597_) );
AOI22X1 AOI22X1_101 ( .A(_6551__bF_buf3), .B(_2__15_), .C(datapath_1_Instr_13_), .D(_6552__bF_buf0), .Y(_6598_) );
NAND3X1 NAND3X1_1306 ( .A(_6596_), .B(_6597_), .C(_6598_), .Y(datapath_1_ALU_aluInB_15_) );
NAND3X1 NAND3X1_1307 ( .A(ALUSrcB_0_bF_buf0_), .B(gnd), .C(_6547__bF_buf1), .Y(_6599_) );
NAND3X1 NAND3X1_1308 ( .A(ALUSrcB_1_bF_buf0_), .B(datapath_1_Instr_15_bF_buf2_), .C(_6549__bF_buf4), .Y(_6600_) );
AOI22X1 AOI22X1_102 ( .A(_6551__bF_buf2), .B(_2__16_), .C(datapath_1_Instr_14_), .D(_6552__bF_buf1), .Y(_6601_) );
NAND3X1 NAND3X1_1309 ( .A(_6599_), .B(_6600_), .C(_6601_), .Y(datapath_1_ALU_aluInB_16_) );
NAND3X1 NAND3X1_1310 ( .A(ALUSrcB_0_bF_buf4_), .B(gnd), .C(_6547__bF_buf4), .Y(_6602_) );
NAND3X1 NAND3X1_1311 ( .A(ALUSrcB_1_bF_buf4_), .B(datapath_1_Instr_15_bF_buf1_), .C(_6549__bF_buf1), .Y(_6603_) );
AOI22X1 AOI22X1_103 ( .A(_6551__bF_buf3), .B(_2__17_), .C(datapath_1_Instr_15_bF_buf0_), .D(_6552__bF_buf0), .Y(_6604_) );
NAND3X1 NAND3X1_1312 ( .A(_6602_), .B(_6603_), .C(_6604_), .Y(datapath_1_ALU_aluInB_17_) );
NAND3X1 NAND3X1_1313 ( .A(ALUSrcB_0_bF_buf3_), .B(gnd), .C(_6547__bF_buf3), .Y(_6605_) );
NAND3X1 NAND3X1_1314 ( .A(ALUSrcB_1_bF_buf3_), .B(datapath_1_Instr_15_bF_buf4_), .C(_6549__bF_buf0), .Y(_6606_) );
AOI22X1 AOI22X1_104 ( .A(_6551__bF_buf1), .B(_2__18_), .C(datapath_1_Instr_15_bF_buf3_), .D(_6552__bF_buf3), .Y(_6607_) );
NAND3X1 NAND3X1_1315 ( .A(_6605_), .B(_6606_), .C(_6607_), .Y(datapath_1_ALU_aluInB_18_) );
NAND3X1 NAND3X1_1316 ( .A(ALUSrcB_0_bF_buf2_), .B(gnd), .C(_6547__bF_buf1), .Y(_6608_) );
NAND3X1 NAND3X1_1317 ( .A(ALUSrcB_1_bF_buf2_), .B(datapath_1_Instr_15_bF_buf2_), .C(_6549__bF_buf2), .Y(_6609_) );
AOI22X1 AOI22X1_105 ( .A(_6551__bF_buf4), .B(_2__19_), .C(datapath_1_Instr_15_bF_buf1_), .D(_6552__bF_buf4), .Y(_6610_) );
NAND3X1 NAND3X1_1318 ( .A(_6608_), .B(_6609_), .C(_6610_), .Y(datapath_1_ALU_aluInB_19_) );
NAND3X1 NAND3X1_1319 ( .A(ALUSrcB_0_bF_buf1_), .B(gnd), .C(_6547__bF_buf4), .Y(_6611_) );
NAND3X1 NAND3X1_1320 ( .A(ALUSrcB_1_bF_buf1_), .B(datapath_1_Instr_15_bF_buf0_), .C(_6549__bF_buf1), .Y(_6612_) );
AOI22X1 AOI22X1_106 ( .A(_6551__bF_buf4), .B(_2__20_), .C(datapath_1_Instr_15_bF_buf4_), .D(_6552__bF_buf4), .Y(_6613_) );
NAND3X1 NAND3X1_1321 ( .A(_6611_), .B(_6612_), .C(_6613_), .Y(datapath_1_ALU_aluInB_20_) );
NAND3X1 NAND3X1_1322 ( .A(ALUSrcB_0_bF_buf0_), .B(gnd), .C(_6547__bF_buf1), .Y(_6614_) );
NAND3X1 NAND3X1_1323 ( .A(ALUSrcB_1_bF_buf0_), .B(datapath_1_Instr_15_bF_buf3_), .C(_6549__bF_buf2), .Y(_6615_) );
AOI22X1 AOI22X1_107 ( .A(_6551__bF_buf4), .B(_2__21_), .C(datapath_1_Instr_15_bF_buf2_), .D(_6552__bF_buf4), .Y(_6616_) );
NAND3X1 NAND3X1_1324 ( .A(_6614_), .B(_6615_), .C(_6616_), .Y(datapath_1_ALU_aluInB_21_) );
NAND3X1 NAND3X1_1325 ( .A(ALUSrcB_0_bF_buf4_), .B(gnd), .C(_6547__bF_buf3), .Y(_6617_) );
NAND3X1 NAND3X1_1326 ( .A(ALUSrcB_1_bF_buf4_), .B(datapath_1_Instr_15_bF_buf1_), .C(_6549__bF_buf0), .Y(_6618_) );
AOI22X1 AOI22X1_108 ( .A(_6551__bF_buf0), .B(_2__22_), .C(datapath_1_Instr_15_bF_buf0_), .D(_6552__bF_buf2), .Y(_6619_) );
NAND3X1 NAND3X1_1327 ( .A(_6617_), .B(_6618_), .C(_6619_), .Y(datapath_1_ALU_aluInB_22_) );
NAND3X1 NAND3X1_1328 ( .A(ALUSrcB_0_bF_buf3_), .B(gnd), .C(_6547__bF_buf2), .Y(_6620_) );
NAND3X1 NAND3X1_1329 ( .A(ALUSrcB_1_bF_buf3_), .B(datapath_1_Instr_15_bF_buf4_), .C(_6549__bF_buf0), .Y(_6621_) );
AOI22X1 AOI22X1_109 ( .A(_6551__bF_buf1), .B(_2__23_), .C(datapath_1_Instr_15_bF_buf3_), .D(_6552__bF_buf3), .Y(_6622_) );
NAND3X1 NAND3X1_1330 ( .A(_6620_), .B(_6621_), .C(_6622_), .Y(datapath_1_ALU_aluInB_23_) );
NAND3X1 NAND3X1_1331 ( .A(ALUSrcB_0_bF_buf2_), .B(gnd), .C(_6547__bF_buf1), .Y(_6623_) );
NAND3X1 NAND3X1_1332 ( .A(ALUSrcB_1_bF_buf2_), .B(datapath_1_Instr_15_bF_buf2_), .C(_6549__bF_buf2), .Y(_6624_) );
AOI22X1 AOI22X1_110 ( .A(_6551__bF_buf4), .B(_2__24_), .C(datapath_1_Instr_15_bF_buf1_), .D(_6552__bF_buf4), .Y(_6625_) );
NAND3X1 NAND3X1_1333 ( .A(_6623_), .B(_6624_), .C(_6625_), .Y(datapath_1_ALU_aluInB_24_) );
NAND3X1 NAND3X1_1334 ( .A(ALUSrcB_0_bF_buf1_), .B(gnd), .C(_6547__bF_buf3), .Y(_6626_) );
NAND3X1 NAND3X1_1335 ( .A(ALUSrcB_1_bF_buf1_), .B(datapath_1_Instr_15_bF_buf0_), .C(_6549__bF_buf3), .Y(_6627_) );
AOI22X1 AOI22X1_111 ( .A(_6551__bF_buf1), .B(_2__25_), .C(datapath_1_Instr_15_bF_buf4_), .D(_6552__bF_buf3), .Y(_6628_) );
NAND3X1 NAND3X1_1336 ( .A(_6626_), .B(_6627_), .C(_6628_), .Y(datapath_1_ALU_aluInB_25_) );
NAND3X1 NAND3X1_1337 ( .A(ALUSrcB_0_bF_buf0_), .B(gnd), .C(_6547__bF_buf3), .Y(_6629_) );
NAND3X1 NAND3X1_1338 ( .A(ALUSrcB_1_bF_buf0_), .B(datapath_1_Instr_15_bF_buf3_), .C(_6549__bF_buf0), .Y(_6630_) );
AOI22X1 AOI22X1_112 ( .A(_6551__bF_buf0), .B(_2__26_), .C(datapath_1_Instr_15_bF_buf2_), .D(_6552__bF_buf2), .Y(_6631_) );
NAND3X1 NAND3X1_1339 ( .A(_6629_), .B(_6630_), .C(_6631_), .Y(datapath_1_ALU_aluInB_26_) );
NAND3X1 NAND3X1_1340 ( .A(ALUSrcB_0_bF_buf4_), .B(gnd), .C(_6547__bF_buf2), .Y(_6632_) );
NAND3X1 NAND3X1_1341 ( .A(ALUSrcB_1_bF_buf4_), .B(datapath_1_Instr_15_bF_buf1_), .C(_6549__bF_buf0), .Y(_6633_) );
AOI22X1 AOI22X1_113 ( .A(_6551__bF_buf1), .B(_2__27_), .C(datapath_1_Instr_15_bF_buf0_), .D(_6552__bF_buf3), .Y(_6634_) );
NAND3X1 NAND3X1_1342 ( .A(_6632_), .B(_6633_), .C(_6634_), .Y(datapath_1_ALU_aluInB_27_) );
NAND3X1 NAND3X1_1343 ( .A(ALUSrcB_0_bF_buf3_), .B(gnd), .C(_6547__bF_buf3), .Y(_6635_) );
NAND3X1 NAND3X1_1344 ( .A(ALUSrcB_1_bF_buf3_), .B(datapath_1_Instr_15_bF_buf4_), .C(_6549__bF_buf2), .Y(_6636_) );
AOI22X1 AOI22X1_114 ( .A(_6551__bF_buf4), .B(_2__28_), .C(datapath_1_Instr_15_bF_buf3_), .D(_6552__bF_buf4), .Y(_6637_) );
NAND3X1 NAND3X1_1345 ( .A(_6635_), .B(_6636_), .C(_6637_), .Y(datapath_1_ALU_aluInB_28_) );
NAND3X1 NAND3X1_1346 ( .A(ALUSrcB_0_bF_buf2_), .B(gnd), .C(_6547__bF_buf1), .Y(_6638_) );
NAND3X1 NAND3X1_1347 ( .A(ALUSrcB_1_bF_buf2_), .B(datapath_1_Instr_15_bF_buf2_), .C(_6549__bF_buf2), .Y(_6639_) );
AOI22X1 AOI22X1_115 ( .A(_6551__bF_buf4), .B(_2__29_), .C(datapath_1_Instr_15_bF_buf1_), .D(_6552__bF_buf4), .Y(_6640_) );
NAND3X1 NAND3X1_1348 ( .A(_6638_), .B(_6639_), .C(_6640_), .Y(datapath_1_ALU_aluInB_29_) );
NAND3X1 NAND3X1_1349 ( .A(ALUSrcB_0_bF_buf1_), .B(gnd), .C(_6547__bF_buf3), .Y(_6641_) );
NAND3X1 NAND3X1_1350 ( .A(ALUSrcB_1_bF_buf1_), .B(datapath_1_Instr_15_bF_buf0_), .C(_6549__bF_buf0), .Y(_6642_) );
AOI22X1 AOI22X1_116 ( .A(_6551__bF_buf0), .B(_2__30_), .C(datapath_1_Instr_15_bF_buf4_), .D(_6552__bF_buf2), .Y(_6643_) );
NAND3X1 NAND3X1_1351 ( .A(_6641_), .B(_6642_), .C(_6643_), .Y(datapath_1_ALU_aluInB_30_) );
NAND3X1 NAND3X1_1352 ( .A(ALUSrcB_0_bF_buf0_), .B(gnd), .C(_6547__bF_buf1), .Y(_6644_) );
NAND3X1 NAND3X1_1353 ( .A(ALUSrcB_1_bF_buf0_), .B(datapath_1_Instr_15_bF_buf3_), .C(_6549__bF_buf2), .Y(_6645_) );
AOI22X1 AOI22X1_117 ( .A(_6551__bF_buf2), .B(_2__31_), .C(datapath_1_Instr_15_bF_buf2_), .D(_6552__bF_buf1), .Y(_6646_) );
NAND3X1 NAND3X1_1354 ( .A(_6644_), .B(_6645_), .C(_6646_), .Y(datapath_1_ALU_aluInB_31_) );
INVX1 INVX1_145 ( .A(datapath_1_Instr_16_bF_buf49_), .Y(_6647_) );
NAND2X1 NAND2X1_456 ( .A(datapath_1_Instr_11_), .B(RegDst), .Y(_6648_) );
OAI21X1 OAI21X1_1349 ( .A(RegDst), .B(_6647_), .C(_6648_), .Y(datapath_1_A3_0_) );
INVX1 INVX1_146 ( .A(datapath_1_Instr_17_bF_buf9_), .Y(_6649_) );
NAND2X1 NAND2X1_457 ( .A(RegDst), .B(datapath_1_Instr_12_), .Y(_6650_) );
OAI21X1 OAI21X1_1350 ( .A(RegDst), .B(_6649_), .C(_6650_), .Y(datapath_1_A3_1_) );
INVX1 INVX1_147 ( .A(datapath_1_Instr_18_bF_buf2_), .Y(_6651_) );
NAND2X1 NAND2X1_458 ( .A(RegDst), .B(datapath_1_Instr_13_), .Y(_6652_) );
OAI21X1 OAI21X1_1351 ( .A(RegDst), .B(_6651_), .C(_6652_), .Y(datapath_1_A3_2_) );
INVX1 INVX1_148 ( .A(datapath_1_Instr_19_bF_buf5_), .Y(_6653_) );
NAND2X1 NAND2X1_459 ( .A(RegDst), .B(datapath_1_Instr_14_), .Y(_6654_) );
OAI21X1 OAI21X1_1352 ( .A(RegDst), .B(_6653_), .C(_6654_), .Y(datapath_1_A3_3_) );
INVX1 INVX1_149 ( .A(datapath_1_Instr_20_bF_buf4_), .Y(_6655_) );
NAND2X1 NAND2X1_460 ( .A(RegDst), .B(datapath_1_Instr_15_bF_buf1_), .Y(_6656_) );
OAI21X1 OAI21X1_1353 ( .A(RegDst), .B(_6655_), .C(_6656_), .Y(datapath_1_A3_4_) );
INVX1 INVX1_150 ( .A(datapath_1_PC_0_), .Y(_6719_) );
NAND2X1 NAND2X1_461 ( .A(datapath_1_ALUOut_0_), .B(IorD_bF_buf1), .Y(_6720_) );
OAI21X1 OAI21X1_1354 ( .A(IorD_bF_buf1), .B(_6719_), .C(_6720_), .Y(_0__0_) );
INVX1 INVX1_151 ( .A(datapath_1_PC_1_), .Y(_6657_) );
NAND2X1 NAND2X1_462 ( .A(IorD_bF_buf1), .B(datapath_1_ALUOut_1_), .Y(_6658_) );
OAI21X1 OAI21X1_1355 ( .A(IorD_bF_buf1), .B(_6657_), .C(_6658_), .Y(_0__1_) );
INVX1 INVX1_152 ( .A(datapath_1_PC_2_), .Y(_6659_) );
NAND2X1 NAND2X1_463 ( .A(IorD_bF_buf5), .B(datapath_1_ALUOut_2_), .Y(_6660_) );
OAI21X1 OAI21X1_1356 ( .A(IorD_bF_buf5), .B(_6659_), .C(_6660_), .Y(_0__2_) );
INVX1 INVX1_153 ( .A(datapath_1_PC_3_), .Y(_6661_) );
NAND2X1 NAND2X1_464 ( .A(IorD_bF_buf3), .B(datapath_1_ALUOut_3_), .Y(_6662_) );
OAI21X1 OAI21X1_1357 ( .A(IorD_bF_buf3), .B(_6661_), .C(_6662_), .Y(_0__3_) );
INVX1 INVX1_154 ( .A(datapath_1_PC_4_), .Y(_6663_) );
NAND2X1 NAND2X1_465 ( .A(IorD_bF_buf3), .B(datapath_1_ALUOut_4_), .Y(_6664_) );
OAI21X1 OAI21X1_1358 ( .A(IorD_bF_buf3), .B(_6663_), .C(_6664_), .Y(_0__4_) );
INVX1 INVX1_155 ( .A(datapath_1_PC_5_), .Y(_6665_) );
NAND2X1 NAND2X1_466 ( .A(IorD_bF_buf5), .B(datapath_1_ALUOut_5_), .Y(_6666_) );
OAI21X1 OAI21X1_1359 ( .A(IorD_bF_buf5), .B(_6665_), .C(_6666_), .Y(_0__5_) );
INVX1 INVX1_156 ( .A(datapath_1_PC_6_), .Y(_6667_) );
NAND2X1 NAND2X1_467 ( .A(IorD_bF_buf5), .B(datapath_1_ALUOut_6_), .Y(_6668_) );
OAI21X1 OAI21X1_1360 ( .A(IorD_bF_buf5), .B(_6667_), .C(_6668_), .Y(_0__6_) );
INVX1 INVX1_157 ( .A(datapath_1_PC_7_), .Y(_6669_) );
NAND2X1 NAND2X1_468 ( .A(IorD_bF_buf3), .B(datapath_1_ALUOut_7_), .Y(_6670_) );
OAI21X1 OAI21X1_1361 ( .A(IorD_bF_buf3), .B(_6669_), .C(_6670_), .Y(_0__7_) );
INVX1 INVX1_158 ( .A(datapath_1_PC_8_), .Y(_6671_) );
NAND2X1 NAND2X1_469 ( .A(IorD_bF_buf0), .B(datapath_1_ALUOut_8_), .Y(_6672_) );
OAI21X1 OAI21X1_1362 ( .A(IorD_bF_buf4), .B(_6671_), .C(_6672_), .Y(_0__8_) );
INVX1 INVX1_159 ( .A(datapath_1_PC_9_), .Y(_6673_) );
NAND2X1 NAND2X1_470 ( .A(IorD_bF_buf4), .B(datapath_1_ALUOut_9_), .Y(_6674_) );
OAI21X1 OAI21X1_1363 ( .A(IorD_bF_buf4), .B(_6673_), .C(_6674_), .Y(_0__9_) );
INVX1 INVX1_160 ( .A(datapath_1_PC_10_), .Y(_6675_) );
NAND2X1 NAND2X1_471 ( .A(IorD_bF_buf4), .B(datapath_1_ALUOut_10_), .Y(_6676_) );
OAI21X1 OAI21X1_1364 ( .A(IorD_bF_buf4), .B(_6675_), .C(_6676_), .Y(_0__10_) );
INVX1 INVX1_161 ( .A(datapath_1_PC_11_), .Y(_6677_) );
NAND2X1 NAND2X1_472 ( .A(IorD_bF_buf7), .B(datapath_1_ALUOut_11_), .Y(_6678_) );
OAI21X1 OAI21X1_1365 ( .A(IorD_bF_buf7), .B(_6677_), .C(_6678_), .Y(_0__11_) );
INVX1 INVX1_162 ( .A(datapath_1_PC_12_), .Y(_6679_) );
NAND2X1 NAND2X1_473 ( .A(IorD_bF_buf7), .B(datapath_1_ALUOut_12_), .Y(_6680_) );
OAI21X1 OAI21X1_1366 ( .A(IorD_bF_buf7), .B(_6679_), .C(_6680_), .Y(_0__12_) );
INVX1 INVX1_163 ( .A(datapath_1_PC_13_), .Y(_6681_) );
NAND2X1 NAND2X1_474 ( .A(IorD_bF_buf2), .B(datapath_1_ALUOut_13_), .Y(_6682_) );
OAI21X1 OAI21X1_1367 ( .A(IorD_bF_buf2), .B(_6681_), .C(_6682_), .Y(_0__13_) );
INVX1 INVX1_164 ( .A(datapath_1_PC_14_), .Y(_6683_) );
NAND2X1 NAND2X1_475 ( .A(IorD_bF_buf6), .B(datapath_1_ALUOut_14_), .Y(_6684_) );
OAI21X1 OAI21X1_1368 ( .A(IorD_bF_buf6), .B(_6683_), .C(_6684_), .Y(_0__14_) );
INVX1 INVX1_165 ( .A(datapath_1_PC_15_), .Y(_6685_) );
NAND2X1 NAND2X1_476 ( .A(IorD_bF_buf6), .B(datapath_1_ALUOut_15_), .Y(_6686_) );
OAI21X1 OAI21X1_1369 ( .A(IorD_bF_buf6), .B(_6685_), .C(_6686_), .Y(_0__15_) );
INVX1 INVX1_166 ( .A(datapath_1_PC_16_), .Y(_6687_) );
NAND2X1 NAND2X1_477 ( .A(IorD_bF_buf7), .B(datapath_1_ALUOut_16_), .Y(_6688_) );
OAI21X1 OAI21X1_1370 ( .A(IorD_bF_buf7), .B(_6687_), .C(_6688_), .Y(_0__16_) );
INVX1 INVX1_167 ( .A(datapath_1_PC_17_), .Y(_6689_) );
NAND2X1 NAND2X1_478 ( .A(IorD_bF_buf3), .B(datapath_1_ALUOut_17_), .Y(_6690_) );
OAI21X1 OAI21X1_1371 ( .A(IorD_bF_buf3), .B(_6689_), .C(_6690_), .Y(_0__17_) );
INVX1 INVX1_168 ( .A(datapath_1_PC_18_), .Y(_6691_) );
NAND2X1 NAND2X1_479 ( .A(IorD_bF_buf0), .B(datapath_1_ALUOut_18_), .Y(_6692_) );
OAI21X1 OAI21X1_1372 ( .A(IorD_bF_buf0), .B(_6691_), .C(_6692_), .Y(_0__18_) );
INVX1 INVX1_169 ( .A(datapath_1_PC_19_), .Y(_6693_) );
NAND2X1 NAND2X1_480 ( .A(IorD_bF_buf2), .B(datapath_1_ALUOut_19_), .Y(_6694_) );
OAI21X1 OAI21X1_1373 ( .A(IorD_bF_buf7), .B(_6693_), .C(_6694_), .Y(_0__19_) );
INVX1 INVX1_170 ( .A(datapath_1_PC_20_), .Y(_6695_) );
NAND2X1 NAND2X1_481 ( .A(IorD_bF_buf5), .B(datapath_1_ALUOut_20_), .Y(_6696_) );
OAI21X1 OAI21X1_1374 ( .A(IorD_bF_buf5), .B(_6695_), .C(_6696_), .Y(_0__20_) );
INVX1 INVX1_171 ( .A(datapath_1_PC_21_), .Y(_6697_) );
NAND2X1 NAND2X1_482 ( .A(IorD_bF_buf1), .B(datapath_1_ALUOut_21_), .Y(_6698_) );
OAI21X1 OAI21X1_1375 ( .A(IorD_bF_buf1), .B(_6697_), .C(_6698_), .Y(_0__21_) );
INVX1 INVX1_172 ( .A(datapath_1_PC_22_), .Y(_6699_) );
NAND2X1 NAND2X1_483 ( .A(IorD_bF_buf2), .B(datapath_1_ALUOut_22_), .Y(_6700_) );
OAI21X1 OAI21X1_1376 ( .A(IorD_bF_buf2), .B(_6699_), .C(_6700_), .Y(_0__22_) );
INVX1 INVX1_173 ( .A(datapath_1_PC_23_), .Y(_6701_) );
NAND2X1 NAND2X1_484 ( .A(IorD_bF_buf2), .B(datapath_1_ALUOut_23_), .Y(_6702_) );
OAI21X1 OAI21X1_1377 ( .A(IorD_bF_buf2), .B(_6701_), .C(_6702_), .Y(_0__23_) );
INVX1 INVX1_174 ( .A(datapath_1_PC_24_), .Y(_6703_) );
NAND2X1 NAND2X1_485 ( .A(IorD_bF_buf0), .B(datapath_1_ALUOut_24_), .Y(_6704_) );
OAI21X1 OAI21X1_1378 ( .A(IorD_bF_buf0), .B(_6703_), .C(_6704_), .Y(_0__24_) );
INVX1 INVX1_175 ( .A(datapath_1_PC_25_), .Y(_6705_) );
NAND2X1 NAND2X1_486 ( .A(IorD_bF_buf1), .B(datapath_1_ALUOut_25_), .Y(_6706_) );
OAI21X1 OAI21X1_1379 ( .A(IorD_bF_buf1), .B(_6705_), .C(_6706_), .Y(_0__25_) );
INVX1 INVX1_176 ( .A(datapath_1_PC_26_), .Y(_6707_) );
NAND2X1 NAND2X1_487 ( .A(IorD_bF_buf6), .B(datapath_1_ALUOut_26_), .Y(_6708_) );
OAI21X1 OAI21X1_1380 ( .A(IorD_bF_buf6), .B(_6707_), .C(_6708_), .Y(_0__26_) );
INVX1 INVX1_177 ( .A(datapath_1_PC_27_), .Y(_6709_) );
NAND2X1 NAND2X1_488 ( .A(IorD_bF_buf6), .B(datapath_1_ALUOut_27_), .Y(_6710_) );
OAI21X1 OAI21X1_1381 ( .A(IorD_bF_buf0), .B(_6709_), .C(_6710_), .Y(_0__27_) );
INVX1 INVX1_178 ( .A(datapath_1_PC_28_), .Y(_6711_) );
NAND2X1 NAND2X1_489 ( .A(IorD_bF_buf4), .B(datapath_1_ALUOut_28_), .Y(_6712_) );
OAI21X1 OAI21X1_1382 ( .A(IorD_bF_buf4), .B(_6711_), .C(_6712_), .Y(_0__28_) );
INVX1 INVX1_179 ( .A(datapath_1_PC_29_), .Y(_6713_) );
NAND2X1 NAND2X1_490 ( .A(IorD_bF_buf7), .B(datapath_1_ALUOut_29_), .Y(_6714_) );
OAI21X1 OAI21X1_1383 ( .A(IorD_bF_buf7), .B(_6713_), .C(_6714_), .Y(_0__29_) );
INVX1 INVX1_180 ( .A(datapath_1_PC_30_), .Y(_6715_) );
NAND2X1 NAND2X1_491 ( .A(IorD_bF_buf2), .B(datapath_1_ALUOut_30_), .Y(_6716_) );
OAI21X1 OAI21X1_1384 ( .A(IorD_bF_buf4), .B(_6715_), .C(_6716_), .Y(_0__30_) );
INVX1 INVX1_181 ( .A(datapath_1_PC_31_), .Y(_6717_) );
NAND2X1 NAND2X1_492 ( .A(IorD_bF_buf0), .B(datapath_1_ALUOut_31_), .Y(_6718_) );
OAI21X1 OAI21X1_1385 ( .A(IorD_bF_buf0), .B(_6717_), .C(_6718_), .Y(_0__31_) );
INVX1 INVX1_182 ( .A(datapath_1_ALUOut_0_), .Y(_6783_) );
NAND2X1 NAND2X1_493 ( .A(datapath_1_Data_0_), .B(MemtoReg_bF_buf7), .Y(_6784_) );
OAI21X1 OAI21X1_1386 ( .A(MemtoReg_bF_buf2), .B(_6783_), .C(_6784_), .Y(datapath_1_RegisterFile_dataWrite_0_) );
INVX1 INVX1_183 ( .A(datapath_1_ALUOut_1_), .Y(_6721_) );
NAND2X1 NAND2X1_494 ( .A(MemtoReg_bF_buf7), .B(datapath_1_Data_1_), .Y(_6722_) );
OAI21X1 OAI21X1_1387 ( .A(MemtoReg_bF_buf2), .B(_6721_), .C(_6722_), .Y(datapath_1_RegisterFile_dataWrite_1_) );
INVX1 INVX1_184 ( .A(datapath_1_ALUOut_2_), .Y(_6723_) );
NAND2X1 NAND2X1_495 ( .A(MemtoReg_bF_buf0), .B(datapath_1_Data_2_), .Y(_6724_) );
OAI21X1 OAI21X1_1388 ( .A(MemtoReg_bF_buf2), .B(_6723_), .C(_6724_), .Y(datapath_1_RegisterFile_dataWrite_2_) );
INVX1 INVX1_185 ( .A(datapath_1_ALUOut_3_), .Y(_6725_) );
NAND2X1 NAND2X1_496 ( .A(MemtoReg_bF_buf0), .B(datapath_1_Data_3_), .Y(_6726_) );
OAI21X1 OAI21X1_1389 ( .A(MemtoReg_bF_buf6), .B(_6725_), .C(_6726_), .Y(datapath_1_RegisterFile_dataWrite_3_) );
INVX1 INVX1_186 ( .A(datapath_1_ALUOut_4_), .Y(_6727_) );
NAND2X1 NAND2X1_497 ( .A(MemtoReg_bF_buf0), .B(datapath_1_Data_4_), .Y(_6728_) );
OAI21X1 OAI21X1_1390 ( .A(MemtoReg_bF_buf6), .B(_6727_), .C(_6728_), .Y(datapath_1_RegisterFile_dataWrite_4_) );
INVX1 INVX1_187 ( .A(datapath_1_ALUOut_5_), .Y(_6729_) );
NAND2X1 NAND2X1_498 ( .A(MemtoReg_bF_buf7), .B(datapath_1_Data_5_), .Y(_6730_) );
OAI21X1 OAI21X1_1391 ( .A(MemtoReg_bF_buf7), .B(_6729_), .C(_6730_), .Y(datapath_1_RegisterFile_dataWrite_5_) );
INVX1 INVX1_188 ( .A(datapath_1_ALUOut_6_), .Y(_6731_) );
NAND2X1 NAND2X1_499 ( .A(MemtoReg_bF_buf7), .B(datapath_1_Data_6_), .Y(_6732_) );
OAI21X1 OAI21X1_1392 ( .A(MemtoReg_bF_buf2), .B(_6731_), .C(_6732_), .Y(datapath_1_RegisterFile_dataWrite_6_) );
INVX1 INVX1_189 ( .A(datapath_1_ALUOut_7_), .Y(_6733_) );
NAND2X1 NAND2X1_500 ( .A(MemtoReg_bF_buf1), .B(datapath_1_Data_7_), .Y(_6734_) );
OAI21X1 OAI21X1_1393 ( .A(MemtoReg_bF_buf2), .B(_6733_), .C(_6734_), .Y(datapath_1_RegisterFile_dataWrite_7_) );
INVX1 INVX1_190 ( .A(datapath_1_ALUOut_8_), .Y(_6735_) );
NAND2X1 NAND2X1_501 ( .A(MemtoReg_bF_buf4), .B(datapath_1_Data_8_), .Y(_6736_) );
OAI21X1 OAI21X1_1394 ( .A(MemtoReg_bF_buf5), .B(_6735_), .C(_6736_), .Y(datapath_1_RegisterFile_dataWrite_8_) );
INVX1 INVX1_191 ( .A(datapath_1_ALUOut_9_), .Y(_6737_) );
NAND2X1 NAND2X1_502 ( .A(MemtoReg_bF_buf4), .B(datapath_1_Data_9_), .Y(_6738_) );
OAI21X1 OAI21X1_1395 ( .A(MemtoReg_bF_buf5), .B(_6737_), .C(_6738_), .Y(datapath_1_RegisterFile_dataWrite_9_) );
INVX1 INVX1_192 ( .A(datapath_1_ALUOut_10_), .Y(_6739_) );
NAND2X1 NAND2X1_503 ( .A(MemtoReg_bF_buf5), .B(datapath_1_Data_10_), .Y(_6740_) );
OAI21X1 OAI21X1_1396 ( .A(MemtoReg_bF_buf5), .B(_6739_), .C(_6740_), .Y(datapath_1_RegisterFile_dataWrite_10_) );
INVX1 INVX1_193 ( .A(datapath_1_ALUOut_11_), .Y(_6741_) );
NAND2X1 NAND2X1_504 ( .A(MemtoReg_bF_buf3), .B(datapath_1_Data_11_), .Y(_6742_) );
OAI21X1 OAI21X1_1397 ( .A(MemtoReg_bF_buf6), .B(_6741_), .C(_6742_), .Y(datapath_1_RegisterFile_dataWrite_11_) );
INVX1 INVX1_194 ( .A(datapath_1_ALUOut_12_), .Y(_6743_) );
NAND2X1 NAND2X1_505 ( .A(MemtoReg_bF_buf1), .B(datapath_1_Data_12_), .Y(_6744_) );
OAI21X1 OAI21X1_1398 ( .A(MemtoReg_bF_buf6), .B(_6743_), .C(_6744_), .Y(datapath_1_RegisterFile_dataWrite_12_) );
INVX1 INVX1_195 ( .A(datapath_1_ALUOut_13_), .Y(_6745_) );
NAND2X1 NAND2X1_506 ( .A(MemtoReg_bF_buf5), .B(datapath_1_Data_13_), .Y(_6746_) );
OAI21X1 OAI21X1_1399 ( .A(MemtoReg_bF_buf5), .B(_6745_), .C(_6746_), .Y(datapath_1_RegisterFile_dataWrite_13_) );
INVX1 INVX1_196 ( .A(datapath_1_ALUOut_14_), .Y(_6747_) );
NAND2X1 NAND2X1_507 ( .A(MemtoReg_bF_buf7), .B(datapath_1_Data_14_), .Y(_6748_) );
OAI21X1 OAI21X1_1400 ( .A(MemtoReg_bF_buf7), .B(_6747_), .C(_6748_), .Y(datapath_1_RegisterFile_dataWrite_14_) );
INVX1 INVX1_197 ( .A(datapath_1_ALUOut_15_), .Y(_6749_) );
NAND2X1 NAND2X1_508 ( .A(MemtoReg_bF_buf0), .B(datapath_1_Data_15_), .Y(_6750_) );
OAI21X1 OAI21X1_1401 ( .A(MemtoReg_bF_buf0), .B(_6749_), .C(_6750_), .Y(datapath_1_RegisterFile_dataWrite_15_) );
INVX1 INVX1_198 ( .A(datapath_1_ALUOut_16_), .Y(_6751_) );
NAND2X1 NAND2X1_509 ( .A(MemtoReg_bF_buf1), .B(datapath_1_Data_16_), .Y(_6752_) );
OAI21X1 OAI21X1_1402 ( .A(MemtoReg_bF_buf6), .B(_6751_), .C(_6752_), .Y(datapath_1_RegisterFile_dataWrite_16_) );
INVX1 INVX1_199 ( .A(datapath_1_ALUOut_17_), .Y(_6753_) );
NAND2X1 NAND2X1_510 ( .A(MemtoReg_bF_buf3), .B(datapath_1_Data_17_), .Y(_6754_) );
OAI21X1 OAI21X1_1403 ( .A(MemtoReg_bF_buf6), .B(_6753_), .C(_6754_), .Y(datapath_1_RegisterFile_dataWrite_17_) );
INVX1 INVX1_200 ( .A(datapath_1_ALUOut_18_), .Y(_6755_) );
NAND2X1 NAND2X1_511 ( .A(MemtoReg_bF_buf1), .B(datapath_1_Data_18_), .Y(_6756_) );
OAI21X1 OAI21X1_1404 ( .A(MemtoReg_bF_buf1), .B(_6755_), .C(_6756_), .Y(datapath_1_RegisterFile_dataWrite_18_) );
INVX1 INVX1_201 ( .A(datapath_1_ALUOut_19_), .Y(_6757_) );
NAND2X1 NAND2X1_512 ( .A(MemtoReg_bF_buf3), .B(datapath_1_Data_19_), .Y(_6758_) );
OAI21X1 OAI21X1_1405 ( .A(MemtoReg_bF_buf6), .B(_6757_), .C(_6758_), .Y(datapath_1_RegisterFile_dataWrite_19_) );
INVX1 INVX1_202 ( .A(datapath_1_ALUOut_20_), .Y(_6759_) );
NAND2X1 NAND2X1_513 ( .A(MemtoReg_bF_buf3), .B(datapath_1_Data_20_), .Y(_6760_) );
OAI21X1 OAI21X1_1406 ( .A(MemtoReg_bF_buf3), .B(_6759_), .C(_6760_), .Y(datapath_1_RegisterFile_dataWrite_20_) );
INVX1 INVX1_203 ( .A(datapath_1_ALUOut_21_), .Y(_6761_) );
NAND2X1 NAND2X1_514 ( .A(MemtoReg_bF_buf7), .B(datapath_1_Data_21_), .Y(_6762_) );
OAI21X1 OAI21X1_1407 ( .A(MemtoReg_bF_buf2), .B(_6761_), .C(_6762_), .Y(datapath_1_RegisterFile_dataWrite_21_) );
INVX1 INVX1_204 ( .A(datapath_1_ALUOut_22_), .Y(_6763_) );
NAND2X1 NAND2X1_515 ( .A(MemtoReg_bF_buf1), .B(datapath_1_Data_22_), .Y(_6764_) );
OAI21X1 OAI21X1_1408 ( .A(MemtoReg_bF_buf0), .B(_6763_), .C(_6764_), .Y(datapath_1_RegisterFile_dataWrite_22_) );
INVX1 INVX1_205 ( .A(datapath_1_ALUOut_23_), .Y(_6765_) );
NAND2X1 NAND2X1_516 ( .A(MemtoReg_bF_buf1), .B(datapath_1_Data_23_), .Y(_6766_) );
OAI21X1 OAI21X1_1409 ( .A(MemtoReg_bF_buf0), .B(_6765_), .C(_6766_), .Y(datapath_1_RegisterFile_dataWrite_23_) );
INVX1 INVX1_206 ( .A(datapath_1_ALUOut_24_), .Y(_6767_) );
NAND2X1 NAND2X1_517 ( .A(MemtoReg_bF_buf1), .B(datapath_1_Data_24_), .Y(_6768_) );
OAI21X1 OAI21X1_1410 ( .A(MemtoReg_bF_buf3), .B(_6767_), .C(_6768_), .Y(datapath_1_RegisterFile_dataWrite_24_) );
INVX1 INVX1_207 ( .A(datapath_1_ALUOut_25_), .Y(_6769_) );
NAND2X1 NAND2X1_518 ( .A(MemtoReg_bF_buf3), .B(datapath_1_Data_25_), .Y(_6770_) );
OAI21X1 OAI21X1_1411 ( .A(MemtoReg_bF_buf3), .B(_6769_), .C(_6770_), .Y(datapath_1_RegisterFile_dataWrite_25_) );
INVX1 INVX1_208 ( .A(datapath_1_ALUOut_26_), .Y(_6771_) );
NAND2X1 NAND2X1_519 ( .A(MemtoReg_bF_buf4), .B(datapath_1_Data_26_), .Y(_6772_) );
OAI21X1 OAI21X1_1412 ( .A(MemtoReg_bF_buf5), .B(_6771_), .C(_6772_), .Y(datapath_1_RegisterFile_dataWrite_26_) );
INVX1 INVX1_209 ( .A(datapath_1_ALUOut_27_), .Y(_6773_) );
NAND2X1 NAND2X1_520 ( .A(MemtoReg_bF_buf4), .B(datapath_1_Data_27_), .Y(_6774_) );
OAI21X1 OAI21X1_1413 ( .A(MemtoReg_bF_buf4), .B(_6773_), .C(_6774_), .Y(datapath_1_RegisterFile_dataWrite_27_) );
INVX1 INVX1_210 ( .A(datapath_1_ALUOut_28_), .Y(_6775_) );
NAND2X1 NAND2X1_521 ( .A(MemtoReg_bF_buf7), .B(datapath_1_Data_28_), .Y(_6776_) );
OAI21X1 OAI21X1_1414 ( .A(MemtoReg_bF_buf2), .B(_6775_), .C(_6776_), .Y(datapath_1_RegisterFile_dataWrite_28_) );
INVX1 INVX1_211 ( .A(datapath_1_ALUOut_29_), .Y(_6777_) );
NAND2X1 NAND2X1_522 ( .A(MemtoReg_bF_buf0), .B(datapath_1_Data_29_), .Y(_6778_) );
OAI21X1 OAI21X1_1415 ( .A(MemtoReg_bF_buf6), .B(_6777_), .C(_6778_), .Y(datapath_1_RegisterFile_dataWrite_29_) );
INVX1 INVX1_212 ( .A(datapath_1_ALUOut_30_), .Y(_6779_) );
NAND2X1 NAND2X1_523 ( .A(MemtoReg_bF_buf4), .B(datapath_1_Data_30_), .Y(_6780_) );
OAI21X1 OAI21X1_1416 ( .A(MemtoReg_bF_buf2), .B(_6779_), .C(_6780_), .Y(datapath_1_RegisterFile_dataWrite_30_) );
INVX1 INVX1_213 ( .A(datapath_1_ALUOut_31_), .Y(_6781_) );
NAND2X1 NAND2X1_524 ( .A(MemtoReg_bF_buf4), .B(datapath_1_Data_31_), .Y(_6782_) );
OAI21X1 OAI21X1_1417 ( .A(MemtoReg_bF_buf4), .B(_6781_), .C(_6782_), .Y(datapath_1_RegisterFile_dataWrite_31_) );
NAND2X1 NAND2X1_525 ( .A(datapath_1_ALU_aluResult_0_), .B(vdd), .Y(_6850_) );
INVX1 INVX1_214 ( .A(vdd), .Y(_6786_) );
NAND2X1 NAND2X1_526 ( .A(datapath_1_ALUOut_0_), .B(_6786__bF_buf0), .Y(_6787_) );
AOI21X1 AOI21X1_313 ( .A(_6787_), .B(_6850_), .C(rst_bF_buf10), .Y(_6785__0_) );
NAND2X1 NAND2X1_527 ( .A(vdd), .B(datapath_1_ALU_aluResult_1_), .Y(_6788_) );
NAND2X1 NAND2X1_528 ( .A(datapath_1_ALUOut_1_), .B(_6786__bF_buf0), .Y(_6789_) );
AOI21X1 AOI21X1_314 ( .A(_6789_), .B(_6788_), .C(rst_bF_buf0), .Y(_6785__1_) );
NAND2X1 NAND2X1_529 ( .A(vdd), .B(datapath_1_ALU_aluResult_2_), .Y(_6790_) );
NAND2X1 NAND2X1_530 ( .A(datapath_1_ALUOut_2_), .B(_6786__bF_buf0), .Y(_6791_) );
AOI21X1 AOI21X1_315 ( .A(_6791_), .B(_6790_), .C(rst_bF_buf0), .Y(_6785__2_) );
NAND2X1 NAND2X1_531 ( .A(vdd), .B(datapath_1_ALU_aluResult_3_), .Y(_6792_) );
NAND2X1 NAND2X1_532 ( .A(datapath_1_ALUOut_3_), .B(_6786__bF_buf2), .Y(_6793_) );
AOI21X1 AOI21X1_316 ( .A(_6793_), .B(_6792_), .C(rst_bF_buf13), .Y(_6785__3_) );
NAND2X1 NAND2X1_533 ( .A(vdd), .B(datapath_1_ALU_aluResult_4_), .Y(_6794_) );
NAND2X1 NAND2X1_534 ( .A(datapath_1_ALUOut_4_), .B(_6786__bF_buf2), .Y(_6795_) );
AOI21X1 AOI21X1_317 ( .A(_6795_), .B(_6794_), .C(rst_bF_buf9), .Y(_6785__4_) );
NAND2X1 NAND2X1_535 ( .A(vdd), .B(datapath_1_ALU_aluResult_5_), .Y(_6796_) );
NAND2X1 NAND2X1_536 ( .A(datapath_1_ALUOut_5_), .B(_6786__bF_buf0), .Y(_6797_) );
AOI21X1 AOI21X1_318 ( .A(_6797_), .B(_6796_), .C(rst_bF_buf10), .Y(_6785__5_) );
NAND2X1 NAND2X1_537 ( .A(vdd), .B(datapath_1_ALU_aluResult_6_), .Y(_6798_) );
NAND2X1 NAND2X1_538 ( .A(datapath_1_ALUOut_6_), .B(_6786__bF_buf0), .Y(_6799_) );
AOI21X1 AOI21X1_319 ( .A(_6799_), .B(_6798_), .C(rst_bF_buf0), .Y(_6785__6_) );
NAND2X1 NAND2X1_539 ( .A(vdd), .B(datapath_1_ALU_aluResult_7_), .Y(_6800_) );
NAND2X1 NAND2X1_540 ( .A(datapath_1_ALUOut_7_), .B(_6786__bF_buf2), .Y(_6801_) );
AOI21X1 AOI21X1_320 ( .A(_6801_), .B(_6800_), .C(rst_bF_buf13), .Y(_6785__7_) );
NAND2X1 NAND2X1_541 ( .A(vdd), .B(datapath_1_ALU_aluResult_8_), .Y(_6802_) );
NAND2X1 NAND2X1_542 ( .A(datapath_1_ALUOut_8_), .B(_6786__bF_buf3), .Y(_6803_) );
AOI21X1 AOI21X1_321 ( .A(_6803_), .B(_6802_), .C(rst_bF_buf11), .Y(_6785__8_) );
NAND2X1 NAND2X1_543 ( .A(vdd), .B(datapath_1_ALU_aluResult_9_), .Y(_6804_) );
NAND2X1 NAND2X1_544 ( .A(datapath_1_ALUOut_9_), .B(_6786__bF_buf4), .Y(_6805_) );
AOI21X1 AOI21X1_322 ( .A(_6805_), .B(_6804_), .C(rst_bF_buf5), .Y(_6785__9_) );
NAND2X1 NAND2X1_545 ( .A(vdd), .B(datapath_1_ALU_aluResult_10_), .Y(_6806_) );
NAND2X1 NAND2X1_546 ( .A(datapath_1_ALUOut_10_), .B(_6786__bF_buf3), .Y(_6807_) );
AOI21X1 AOI21X1_323 ( .A(_6807_), .B(_6806_), .C(rst_bF_buf11), .Y(_6785__10_) );
NAND2X1 NAND2X1_547 ( .A(vdd), .B(datapath_1_ALU_aluResult_11_), .Y(_6808_) );
NAND2X1 NAND2X1_548 ( .A(datapath_1_ALUOut_11_), .B(_6786__bF_buf4), .Y(_6809_) );
AOI21X1 AOI21X1_324 ( .A(_6809_), .B(_6808_), .C(rst_bF_buf5), .Y(_6785__11_) );
NAND2X1 NAND2X1_549 ( .A(vdd), .B(datapath_1_ALU_aluResult_12_), .Y(_6810_) );
NAND2X1 NAND2X1_550 ( .A(datapath_1_ALUOut_12_), .B(_6786__bF_buf4), .Y(_6811_) );
AOI21X1 AOI21X1_325 ( .A(_6811_), .B(_6810_), .C(rst_bF_buf7), .Y(_6785__12_) );
NAND2X1 NAND2X1_551 ( .A(vdd), .B(datapath_1_ALU_aluResult_13_), .Y(_6812_) );
NAND2X1 NAND2X1_552 ( .A(datapath_1_ALUOut_13_), .B(_6786__bF_buf3), .Y(_6813_) );
AOI21X1 AOI21X1_326 ( .A(_6813_), .B(_6812_), .C(rst_bF_buf11), .Y(_6785__13_) );
NAND2X1 NAND2X1_553 ( .A(vdd), .B(datapath_1_ALU_aluResult_14_), .Y(_6814_) );
NAND2X1 NAND2X1_554 ( .A(datapath_1_ALUOut_14_), .B(_6786__bF_buf3), .Y(_6815_) );
AOI21X1 AOI21X1_327 ( .A(_6815_), .B(_6814_), .C(rst_bF_buf11), .Y(_6785__14_) );
NAND2X1 NAND2X1_555 ( .A(vdd), .B(datapath_1_ALU_aluResult_15_), .Y(_6816_) );
NAND2X1 NAND2X1_556 ( .A(datapath_1_ALUOut_15_), .B(_6786__bF_buf1), .Y(_6817_) );
AOI21X1 AOI21X1_328 ( .A(_6817_), .B(_6816_), .C(rst_bF_buf11), .Y(_6785__15_) );
NAND2X1 NAND2X1_557 ( .A(vdd), .B(datapath_1_ALU_aluResult_16_), .Y(_6818_) );
NAND2X1 NAND2X1_558 ( .A(datapath_1_ALUOut_16_), .B(_6786__bF_buf2), .Y(_6819_) );
AOI21X1 AOI21X1_329 ( .A(_6819_), .B(_6818_), .C(rst_bF_buf7), .Y(_6785__16_) );
NAND2X1 NAND2X1_559 ( .A(vdd), .B(datapath_1_ALU_aluResult_17_), .Y(_6820_) );
NAND2X1 NAND2X1_560 ( .A(datapath_1_ALUOut_17_), .B(_6786__bF_buf2), .Y(_6821_) );
AOI21X1 AOI21X1_330 ( .A(_6821_), .B(_6820_), .C(rst_bF_buf7), .Y(_6785__17_) );
NAND2X1 NAND2X1_561 ( .A(vdd), .B(datapath_1_ALU_aluResult_18_), .Y(_6822_) );
NAND2X1 NAND2X1_562 ( .A(datapath_1_ALUOut_18_), .B(_6786__bF_buf1), .Y(_6823_) );
AOI21X1 AOI21X1_331 ( .A(_6823_), .B(_6822_), .C(rst_bF_buf11), .Y(_6785__18_) );
NAND2X1 NAND2X1_563 ( .A(vdd), .B(datapath_1_ALU_aluResult_19_), .Y(_6824_) );
NAND2X1 NAND2X1_564 ( .A(datapath_1_ALUOut_19_), .B(_6786__bF_buf4), .Y(_6825_) );
AOI21X1 AOI21X1_332 ( .A(_6825_), .B(_6824_), .C(rst_bF_buf5), .Y(_6785__19_) );
NAND2X1 NAND2X1_565 ( .A(vdd), .B(datapath_1_ALU_aluResult_20_), .Y(_6826_) );
NAND2X1 NAND2X1_566 ( .A(datapath_1_ALUOut_20_), .B(_6786__bF_buf1), .Y(_6827_) );
AOI21X1 AOI21X1_333 ( .A(_6827_), .B(_6826_), .C(rst_bF_buf10), .Y(_6785__20_) );
NAND2X1 NAND2X1_567 ( .A(vdd), .B(datapath_1_ALU_aluResult_21_), .Y(_6828_) );
NAND2X1 NAND2X1_568 ( .A(datapath_1_ALUOut_21_), .B(_6786__bF_buf0), .Y(_6829_) );
AOI21X1 AOI21X1_334 ( .A(_6829_), .B(_6828_), .C(rst_bF_buf10), .Y(_6785__21_) );
NAND2X1 NAND2X1_569 ( .A(vdd), .B(datapath_1_ALU_aluResult_22_), .Y(_6830_) );
NAND2X1 NAND2X1_570 ( .A(datapath_1_ALUOut_22_), .B(_6786__bF_buf2), .Y(_6831_) );
AOI21X1 AOI21X1_335 ( .A(_6831_), .B(_6830_), .C(rst_bF_buf9), .Y(_6785__22_) );
NAND2X1 NAND2X1_571 ( .A(vdd), .B(datapath_1_ALU_aluResult_23_), .Y(_6832_) );
NAND2X1 NAND2X1_572 ( .A(datapath_1_ALUOut_23_), .B(_6786__bF_buf4), .Y(_6833_) );
AOI21X1 AOI21X1_336 ( .A(_6833_), .B(_6832_), .C(rst_bF_buf5), .Y(_6785__23_) );
NAND2X1 NAND2X1_573 ( .A(vdd), .B(datapath_1_ALU_aluResult_24_), .Y(_6834_) );
NAND2X1 NAND2X1_574 ( .A(datapath_1_ALUOut_24_), .B(_6786__bF_buf3), .Y(_6835_) );
AOI21X1 AOI21X1_337 ( .A(_6835_), .B(_6834_), .C(rst_bF_buf11), .Y(_6785__24_) );
NAND2X1 NAND2X1_575 ( .A(vdd), .B(datapath_1_ALU_aluResult_25_), .Y(_6836_) );
NAND2X1 NAND2X1_576 ( .A(datapath_1_ALUOut_25_), .B(_6786__bF_buf1), .Y(_6837_) );
AOI21X1 AOI21X1_338 ( .A(_6837_), .B(_6836_), .C(rst_bF_buf10), .Y(_6785__25_) );
NAND2X1 NAND2X1_577 ( .A(vdd), .B(datapath_1_ALU_aluResult_26_), .Y(_6838_) );
NAND2X1 NAND2X1_578 ( .A(datapath_1_ALUOut_26_), .B(_6786__bF_buf1), .Y(_6839_) );
AOI21X1 AOI21X1_339 ( .A(_6839_), .B(_6838_), .C(rst_bF_buf11), .Y(_6785__26_) );
NAND2X1 NAND2X1_579 ( .A(vdd), .B(datapath_1_ALU_aluResult_27_), .Y(_6840_) );
NAND2X1 NAND2X1_580 ( .A(datapath_1_ALUOut_27_), .B(_6786__bF_buf3), .Y(_6841_) );
AOI21X1 AOI21X1_340 ( .A(_6841_), .B(_6840_), .C(rst_bF_buf11), .Y(_6785__27_) );
NAND2X1 NAND2X1_581 ( .A(vdd), .B(datapath_1_ALU_aluResult_28_), .Y(_6842_) );
NAND2X1 NAND2X1_582 ( .A(datapath_1_ALUOut_28_), .B(_6786__bF_buf1), .Y(_6843_) );
AOI21X1 AOI21X1_341 ( .A(_6843_), .B(_6842_), .C(rst_bF_buf11), .Y(_6785__28_) );
NAND2X1 NAND2X1_583 ( .A(vdd), .B(datapath_1_ALU_aluResult_29_), .Y(_6844_) );
NAND2X1 NAND2X1_584 ( .A(datapath_1_ALUOut_29_), .B(_6786__bF_buf4), .Y(_6845_) );
AOI21X1 AOI21X1_342 ( .A(_6845_), .B(_6844_), .C(rst_bF_buf5), .Y(_6785__29_) );
NAND2X1 NAND2X1_585 ( .A(vdd), .B(datapath_1_ALU_aluResult_30_), .Y(_6846_) );
NAND2X1 NAND2X1_586 ( .A(datapath_1_ALUOut_30_), .B(_6786__bF_buf4), .Y(_6847_) );
AOI21X1 AOI21X1_343 ( .A(_6847_), .B(_6846_), .C(rst_bF_buf5), .Y(_6785__30_) );
NAND2X1 NAND2X1_587 ( .A(vdd), .B(datapath_1_ALU_aluResult_31_), .Y(_6848_) );
NAND2X1 NAND2X1_588 ( .A(datapath_1_ALUOut_31_), .B(_6786__bF_buf3), .Y(_6849_) );
AOI21X1 AOI21X1_344 ( .A(_6849_), .B(_6848_), .C(rst_bF_buf11), .Y(_6785__31_) );
DFFPOSX1 DFFPOSX1_1025 ( .CLK(clk_bF_buf71), .D(_6785__0_), .Q(datapath_1_ALUOut_0_) );
DFFPOSX1 DFFPOSX1_1026 ( .CLK(clk_bF_buf71), .D(_6785__1_), .Q(datapath_1_ALUOut_1_) );
DFFPOSX1 DFFPOSX1_1027 ( .CLK(clk_bF_buf71), .D(_6785__2_), .Q(datapath_1_ALUOut_2_) );
DFFPOSX1 DFFPOSX1_1028 ( .CLK(clk_bF_buf97), .D(_6785__3_), .Q(datapath_1_ALUOut_3_) );
DFFPOSX1 DFFPOSX1_1029 ( .CLK(clk_bF_buf43), .D(_6785__4_), .Q(datapath_1_ALUOut_4_) );
DFFPOSX1 DFFPOSX1_1030 ( .CLK(clk_bF_buf24), .D(_6785__5_), .Q(datapath_1_ALUOut_5_) );
DFFPOSX1 DFFPOSX1_1031 ( .CLK(clk_bF_buf71), .D(_6785__6_), .Q(datapath_1_ALUOut_6_) );
DFFPOSX1 DFFPOSX1_1032 ( .CLK(clk_bF_buf97), .D(_6785__7_), .Q(datapath_1_ALUOut_7_) );
DFFPOSX1 DFFPOSX1_1033 ( .CLK(clk_bF_buf0), .D(_6785__8_), .Q(datapath_1_ALUOut_8_) );
DFFPOSX1 DFFPOSX1_1034 ( .CLK(clk_bF_buf108), .D(_6785__9_), .Q(datapath_1_ALUOut_9_) );
DFFPOSX1 DFFPOSX1_1035 ( .CLK(clk_bF_buf50), .D(_6785__10_), .Q(datapath_1_ALUOut_10_) );
DFFPOSX1 DFFPOSX1_1036 ( .CLK(clk_bF_buf108), .D(_6785__11_), .Q(datapath_1_ALUOut_11_) );
DFFPOSX1 DFFPOSX1_1037 ( .CLK(clk_bF_buf91), .D(_6785__12_), .Q(datapath_1_ALUOut_12_) );
DFFPOSX1 DFFPOSX1_1038 ( .CLK(clk_bF_buf50), .D(_6785__13_), .Q(datapath_1_ALUOut_13_) );
DFFPOSX1 DFFPOSX1_1039 ( .CLK(clk_bF_buf50), .D(_6785__14_), .Q(datapath_1_ALUOut_14_) );
DFFPOSX1 DFFPOSX1_1040 ( .CLK(clk_bF_buf0), .D(_6785__15_), .Q(datapath_1_ALUOut_15_) );
DFFPOSX1 DFFPOSX1_1041 ( .CLK(clk_bF_buf91), .D(_6785__16_), .Q(datapath_1_ALUOut_16_) );
DFFPOSX1 DFFPOSX1_1042 ( .CLK(clk_bF_buf97), .D(_6785__17_), .Q(datapath_1_ALUOut_17_) );
DFFPOSX1 DFFPOSX1_1043 ( .CLK(clk_bF_buf0), .D(_6785__18_), .Q(datapath_1_ALUOut_18_) );
DFFPOSX1 DFFPOSX1_1044 ( .CLK(clk_bF_buf108), .D(_6785__19_), .Q(datapath_1_ALUOut_19_) );
DFFPOSX1 DFFPOSX1_1045 ( .CLK(clk_bF_buf0), .D(_6785__20_), .Q(datapath_1_ALUOut_20_) );
DFFPOSX1 DFFPOSX1_1046 ( .CLK(clk_bF_buf71), .D(_6785__21_), .Q(datapath_1_ALUOut_21_) );
DFFPOSX1 DFFPOSX1_1047 ( .CLK(clk_bF_buf43), .D(_6785__22_), .Q(datapath_1_ALUOut_22_) );
DFFPOSX1 DFFPOSX1_1048 ( .CLK(clk_bF_buf108), .D(_6785__23_), .Q(datapath_1_ALUOut_23_) );
DFFPOSX1 DFFPOSX1_1049 ( .CLK(clk_bF_buf50), .D(_6785__24_), .Q(datapath_1_ALUOut_24_) );
DFFPOSX1 DFFPOSX1_1050 ( .CLK(clk_bF_buf24), .D(_6785__25_), .Q(datapath_1_ALUOut_25_) );
DFFPOSX1 DFFPOSX1_1051 ( .CLK(clk_bF_buf0), .D(_6785__26_), .Q(datapath_1_ALUOut_26_) );
DFFPOSX1 DFFPOSX1_1052 ( .CLK(clk_bF_buf0), .D(_6785__27_), .Q(datapath_1_ALUOut_27_) );
DFFPOSX1 DFFPOSX1_1053 ( .CLK(clk_bF_buf50), .D(_6785__28_), .Q(datapath_1_ALUOut_28_) );
DFFPOSX1 DFFPOSX1_1054 ( .CLK(clk_bF_buf108), .D(_6785__29_), .Q(datapath_1_ALUOut_29_) );
DFFPOSX1 DFFPOSX1_1055 ( .CLK(clk_bF_buf108), .D(_6785__30_), .Q(datapath_1_ALUOut_30_) );
DFFPOSX1 DFFPOSX1_1056 ( .CLK(clk_bF_buf50), .D(_6785__31_), .Q(datapath_1_ALUOut_31_) );
NAND2X1 NAND2X1_589 ( .A(datapath_1_RD1_0_), .B(vdd), .Y(_6916_) );
INVX1 INVX1_215 ( .A(vdd), .Y(_6852_) );
NAND2X1 NAND2X1_590 ( .A(datapath_1_A_0_), .B(_6852__bF_buf1), .Y(_6853_) );
AOI21X1 AOI21X1_345 ( .A(_6853_), .B(_6916_), .C(rst_bF_buf9), .Y(_6851__0_) );
NAND2X1 NAND2X1_591 ( .A(vdd), .B(datapath_1_RD1_1_), .Y(_6854_) );
NAND2X1 NAND2X1_592 ( .A(datapath_1_A_1_), .B(_6852__bF_buf3), .Y(_6855_) );
AOI21X1 AOI21X1_346 ( .A(_6855_), .B(_6854_), .C(rst_bF_buf3), .Y(_6851__1_) );
NAND2X1 NAND2X1_593 ( .A(vdd), .B(datapath_1_RD1_2_), .Y(_6856_) );
NAND2X1 NAND2X1_594 ( .A(datapath_1_A_2_), .B(_6852__bF_buf2), .Y(_6857_) );
AOI21X1 AOI21X1_347 ( .A(_6857_), .B(_6856_), .C(rst_bF_buf3), .Y(_6851__2_) );
NAND2X1 NAND2X1_595 ( .A(vdd), .B(datapath_1_RD1_3_), .Y(_6858_) );
NAND2X1 NAND2X1_596 ( .A(datapath_1_A_3_), .B(_6852__bF_buf3), .Y(_6859_) );
AOI21X1 AOI21X1_348 ( .A(_6859_), .B(_6858_), .C(rst_bF_buf8), .Y(_6851__3_) );
NAND2X1 NAND2X1_597 ( .A(vdd), .B(datapath_1_RD1_4_), .Y(_6860_) );
NAND2X1 NAND2X1_598 ( .A(datapath_1_A_4_), .B(_6852__bF_buf1), .Y(_6861_) );
AOI21X1 AOI21X1_349 ( .A(_6861_), .B(_6860_), .C(rst_bF_buf9), .Y(_6851__4_) );
NAND2X1 NAND2X1_599 ( .A(vdd), .B(datapath_1_RD1_5_), .Y(_6862_) );
NAND2X1 NAND2X1_600 ( .A(datapath_1_A_5_), .B(_6852__bF_buf1), .Y(_6863_) );
AOI21X1 AOI21X1_350 ( .A(_6863_), .B(_6862_), .C(rst_bF_buf9), .Y(_6851__5_) );
NAND2X1 NAND2X1_601 ( .A(vdd), .B(datapath_1_RD1_6_), .Y(_6864_) );
NAND2X1 NAND2X1_602 ( .A(datapath_1_A_6_), .B(_6852__bF_buf4), .Y(_6865_) );
AOI21X1 AOI21X1_351 ( .A(_6865_), .B(_6864_), .C(rst_bF_buf13), .Y(_6851__6_) );
NAND2X1 NAND2X1_603 ( .A(vdd), .B(datapath_1_RD1_7_), .Y(_6866_) );
NAND2X1 NAND2X1_604 ( .A(datapath_1_A_7_), .B(_6852__bF_buf3), .Y(_6867_) );
AOI21X1 AOI21X1_352 ( .A(_6867_), .B(_6866_), .C(rst_bF_buf1), .Y(_6851__7_) );
NAND2X1 NAND2X1_605 ( .A(vdd), .B(datapath_1_RD1_8_), .Y(_6868_) );
NAND2X1 NAND2X1_606 ( .A(datapath_1_A_8_), .B(_6852__bF_buf4), .Y(_6869_) );
AOI21X1 AOI21X1_353 ( .A(_6869_), .B(_6868_), .C(rst_bF_buf7), .Y(_6851__8_) );
NAND2X1 NAND2X1_607 ( .A(vdd), .B(datapath_1_RD1_9_), .Y(_6870_) );
NAND2X1 NAND2X1_608 ( .A(datapath_1_A_9_), .B(_6852__bF_buf4), .Y(_6871_) );
AOI21X1 AOI21X1_354 ( .A(_6871_), .B(_6870_), .C(rst_bF_buf13), .Y(_6851__9_) );
NAND2X1 NAND2X1_609 ( .A(vdd), .B(datapath_1_RD1_10_), .Y(_6872_) );
NAND2X1 NAND2X1_610 ( .A(datapath_1_A_10_), .B(_6852__bF_buf0), .Y(_6873_) );
AOI21X1 AOI21X1_355 ( .A(_6873_), .B(_6872_), .C(rst_bF_buf13), .Y(_6851__10_) );
NAND2X1 NAND2X1_611 ( .A(vdd), .B(datapath_1_RD1_11_), .Y(_6874_) );
NAND2X1 NAND2X1_612 ( .A(datapath_1_A_11_), .B(_6852__bF_buf3), .Y(_6875_) );
AOI21X1 AOI21X1_356 ( .A(_6875_), .B(_6874_), .C(rst_bF_buf8), .Y(_6851__11_) );
NAND2X1 NAND2X1_613 ( .A(vdd), .B(datapath_1_RD1_12_), .Y(_6876_) );
NAND2X1 NAND2X1_614 ( .A(datapath_1_A_12_), .B(_6852__bF_buf4), .Y(_6877_) );
AOI21X1 AOI21X1_357 ( .A(_6877_), .B(_6876_), .C(rst_bF_buf3), .Y(_6851__12_) );
NAND2X1 NAND2X1_615 ( .A(vdd), .B(datapath_1_RD1_13_), .Y(_6878_) );
NAND2X1 NAND2X1_616 ( .A(datapath_1_A_13_), .B(_6852__bF_buf0), .Y(_6879_) );
AOI21X1 AOI21X1_358 ( .A(_6879_), .B(_6878_), .C(rst_bF_buf13), .Y(_6851__13_) );
NAND2X1 NAND2X1_617 ( .A(vdd), .B(datapath_1_RD1_14_), .Y(_6880_) );
NAND2X1 NAND2X1_618 ( .A(datapath_1_A_14_), .B(_6852__bF_buf0), .Y(_6881_) );
AOI21X1 AOI21X1_359 ( .A(_6881_), .B(_6880_), .C(rst_bF_buf13), .Y(_6851__14_) );
NAND2X1 NAND2X1_619 ( .A(vdd), .B(datapath_1_RD1_15_), .Y(_6882_) );
NAND2X1 NAND2X1_620 ( .A(datapath_1_A_15_), .B(_6852__bF_buf2), .Y(_6883_) );
AOI21X1 AOI21X1_360 ( .A(_6883_), .B(_6882_), .C(rst_bF_buf8), .Y(_6851__15_) );
NAND2X1 NAND2X1_621 ( .A(vdd), .B(datapath_1_RD1_16_), .Y(_6884_) );
NAND2X1 NAND2X1_622 ( .A(datapath_1_A_16_), .B(_6852__bF_buf2), .Y(_6885_) );
AOI21X1 AOI21X1_361 ( .A(_6885_), .B(_6884_), .C(rst_bF_buf8), .Y(_6851__16_) );
NAND2X1 NAND2X1_623 ( .A(vdd), .B(datapath_1_RD1_17_), .Y(_6886_) );
NAND2X1 NAND2X1_624 ( .A(datapath_1_A_17_), .B(_6852__bF_buf0), .Y(_6887_) );
AOI21X1 AOI21X1_362 ( .A(_6887_), .B(_6886_), .C(rst_bF_buf3), .Y(_6851__17_) );
NAND2X1 NAND2X1_625 ( .A(vdd), .B(datapath_1_RD1_18_), .Y(_6888_) );
NAND2X1 NAND2X1_626 ( .A(datapath_1_A_18_), .B(_6852__bF_buf1), .Y(_6889_) );
AOI21X1 AOI21X1_363 ( .A(_6889_), .B(_6888_), .C(rst_bF_buf9), .Y(_6851__18_) );
NAND2X1 NAND2X1_627 ( .A(vdd), .B(datapath_1_RD1_19_), .Y(_6890_) );
NAND2X1 NAND2X1_628 ( .A(datapath_1_A_19_), .B(_6852__bF_buf2), .Y(_6891_) );
AOI21X1 AOI21X1_364 ( .A(_6891_), .B(_6890_), .C(rst_bF_buf8), .Y(_6851__19_) );
NAND2X1 NAND2X1_629 ( .A(vdd), .B(datapath_1_RD1_20_), .Y(_6892_) );
NAND2X1 NAND2X1_630 ( .A(datapath_1_A_20_), .B(_6852__bF_buf4), .Y(_6893_) );
AOI21X1 AOI21X1_365 ( .A(_6893_), .B(_6892_), .C(rst_bF_buf3), .Y(_6851__20_) );
NAND2X1 NAND2X1_631 ( .A(vdd), .B(datapath_1_RD1_21_), .Y(_6894_) );
NAND2X1 NAND2X1_632 ( .A(datapath_1_A_21_), .B(_6852__bF_buf0), .Y(_6895_) );
AOI21X1 AOI21X1_366 ( .A(_6895_), .B(_6894_), .C(rst_bF_buf13), .Y(_6851__21_) );
NAND2X1 NAND2X1_633 ( .A(vdd), .B(datapath_1_RD1_22_), .Y(_6896_) );
NAND2X1 NAND2X1_634 ( .A(datapath_1_A_22_), .B(_6852__bF_buf0), .Y(_6897_) );
AOI21X1 AOI21X1_367 ( .A(_6897_), .B(_6896_), .C(rst_bF_buf9), .Y(_6851__22_) );
NAND2X1 NAND2X1_635 ( .A(vdd), .B(datapath_1_RD1_23_), .Y(_6898_) );
NAND2X1 NAND2X1_636 ( .A(datapath_1_A_23_), .B(_6852__bF_buf3), .Y(_6899_) );
AOI21X1 AOI21X1_368 ( .A(_6899_), .B(_6898_), .C(rst_bF_buf3), .Y(_6851__23_) );
NAND2X1 NAND2X1_637 ( .A(vdd), .B(datapath_1_RD1_24_), .Y(_6900_) );
NAND2X1 NAND2X1_638 ( .A(datapath_1_A_24_), .B(_6852__bF_buf3), .Y(_6901_) );
AOI21X1 AOI21X1_369 ( .A(_6901_), .B(_6900_), .C(rst_bF_buf8), .Y(_6851__24_) );
NAND2X1 NAND2X1_639 ( .A(vdd), .B(datapath_1_RD1_25_), .Y(_6902_) );
NAND2X1 NAND2X1_640 ( .A(datapath_1_A_25_), .B(_6852__bF_buf2), .Y(_6903_) );
AOI21X1 AOI21X1_370 ( .A(_6903_), .B(_6902_), .C(rst_bF_buf8), .Y(_6851__25_) );
NAND2X1 NAND2X1_641 ( .A(vdd), .B(datapath_1_RD1_26_), .Y(_6904_) );
NAND2X1 NAND2X1_642 ( .A(datapath_1_A_26_), .B(_6852__bF_buf1), .Y(_6905_) );
AOI21X1 AOI21X1_371 ( .A(_6905_), .B(_6904_), .C(rst_bF_buf9), .Y(_6851__26_) );
NAND2X1 NAND2X1_643 ( .A(vdd), .B(datapath_1_RD1_27_), .Y(_6906_) );
NAND2X1 NAND2X1_644 ( .A(datapath_1_A_27_), .B(_6852__bF_buf4), .Y(_6907_) );
AOI21X1 AOI21X1_372 ( .A(_6907_), .B(_6906_), .C(rst_bF_buf3), .Y(_6851__27_) );
NAND2X1 NAND2X1_645 ( .A(vdd), .B(datapath_1_RD1_28_), .Y(_6908_) );
NAND2X1 NAND2X1_646 ( .A(datapath_1_A_28_), .B(_6852__bF_buf2), .Y(_6909_) );
AOI21X1 AOI21X1_373 ( .A(_6909_), .B(_6908_), .C(rst_bF_buf1), .Y(_6851__28_) );
NAND2X1 NAND2X1_647 ( .A(vdd), .B(datapath_1_RD1_29_), .Y(_6910_) );
NAND2X1 NAND2X1_648 ( .A(datapath_1_A_29_), .B(_6852__bF_buf3), .Y(_6911_) );
AOI21X1 AOI21X1_374 ( .A(_6911_), .B(_6910_), .C(rst_bF_buf8), .Y(_6851__29_) );
NAND2X1 NAND2X1_649 ( .A(vdd), .B(datapath_1_RD1_30_), .Y(_6912_) );
NAND2X1 NAND2X1_650 ( .A(datapath_1_A_30_), .B(_6852__bF_buf4), .Y(_6913_) );
AOI21X1 AOI21X1_375 ( .A(_6913_), .B(_6912_), .C(rst_bF_buf13), .Y(_6851__30_) );
NAND2X1 NAND2X1_651 ( .A(vdd), .B(datapath_1_RD1_31_), .Y(_6914_) );
NAND2X1 NAND2X1_652 ( .A(datapath_1_A_31_), .B(_6852__bF_buf1), .Y(_6915_) );
AOI21X1 AOI21X1_376 ( .A(_6915_), .B(_6914_), .C(rst_bF_buf9), .Y(_6851__31_) );
DFFPOSX1 DFFPOSX1_1057 ( .CLK(clk_bF_buf43), .D(_6851__0_), .Q(datapath_1_A_0_) );
DFFPOSX1 DFFPOSX1_1058 ( .CLK(clk_bF_buf104), .D(_6851__1_), .Q(datapath_1_A_1_) );
DFFPOSX1 DFFPOSX1_1059 ( .CLK(clk_bF_buf104), .D(_6851__2_), .Q(datapath_1_A_2_) );
DFFPOSX1 DFFPOSX1_1060 ( .CLK(clk_bF_buf10), .D(_6851__3_), .Q(datapath_1_A_3_) );
DFFPOSX1 DFFPOSX1_1061 ( .CLK(clk_bF_buf43), .D(_6851__4_), .Q(datapath_1_A_4_) );
DFFPOSX1 DFFPOSX1_1062 ( .CLK(clk_bF_buf88), .D(_6851__5_), .Q(datapath_1_A_5_) );
DFFPOSX1 DFFPOSX1_1063 ( .CLK(clk_bF_buf52), .D(_6851__6_), .Q(datapath_1_A_6_) );
DFFPOSX1 DFFPOSX1_1064 ( .CLK(clk_bF_buf10), .D(_6851__7_), .Q(datapath_1_A_7_) );
DFFPOSX1 DFFPOSX1_1065 ( .CLK(clk_bF_buf91), .D(_6851__8_), .Q(datapath_1_A_8_) );
DFFPOSX1 DFFPOSX1_1066 ( .CLK(clk_bF_buf97), .D(_6851__9_), .Q(datapath_1_A_9_) );
DFFPOSX1 DFFPOSX1_1067 ( .CLK(clk_bF_buf52), .D(_6851__10_), .Q(datapath_1_A_10_) );
DFFPOSX1 DFFPOSX1_1068 ( .CLK(clk_bF_buf10), .D(_6851__11_), .Q(datapath_1_A_11_) );
DFFPOSX1 DFFPOSX1_1069 ( .CLK(clk_bF_buf104), .D(_6851__12_), .Q(datapath_1_A_12_) );
DFFPOSX1 DFFPOSX1_1070 ( .CLK(clk_bF_buf43), .D(_6851__13_), .Q(datapath_1_A_13_) );
DFFPOSX1 DFFPOSX1_1071 ( .CLK(clk_bF_buf57), .D(_6851__14_), .Q(datapath_1_A_14_) );
DFFPOSX1 DFFPOSX1_1072 ( .CLK(clk_bF_buf10), .D(_6851__15_), .Q(datapath_1_A_15_) );
DFFPOSX1 DFFPOSX1_1073 ( .CLK(clk_bF_buf10), .D(_6851__16_), .Q(datapath_1_A_16_) );
DFFPOSX1 DFFPOSX1_1074 ( .CLK(clk_bF_buf52), .D(_6851__17_), .Q(datapath_1_A_17_) );
DFFPOSX1 DFFPOSX1_1075 ( .CLK(clk_bF_buf43), .D(_6851__18_), .Q(datapath_1_A_18_) );
DFFPOSX1 DFFPOSX1_1076 ( .CLK(clk_bF_buf10), .D(_6851__19_), .Q(datapath_1_A_19_) );
DFFPOSX1 DFFPOSX1_1077 ( .CLK(clk_bF_buf104), .D(_6851__20_), .Q(datapath_1_A_20_) );
DFFPOSX1 DFFPOSX1_1078 ( .CLK(clk_bF_buf57), .D(_6851__21_), .Q(datapath_1_A_21_) );
DFFPOSX1 DFFPOSX1_1079 ( .CLK(clk_bF_buf52), .D(_6851__22_), .Q(datapath_1_A_22_) );
DFFPOSX1 DFFPOSX1_1080 ( .CLK(clk_bF_buf104), .D(_6851__23_), .Q(datapath_1_A_23_) );
DFFPOSX1 DFFPOSX1_1081 ( .CLK(clk_bF_buf65), .D(_6851__24_), .Q(datapath_1_A_24_) );
DFFPOSX1 DFFPOSX1_1082 ( .CLK(clk_bF_buf10), .D(_6851__25_), .Q(datapath_1_A_25_) );
DFFPOSX1 DFFPOSX1_1083 ( .CLK(clk_bF_buf43), .D(_6851__26_), .Q(datapath_1_A_26_) );
DFFPOSX1 DFFPOSX1_1084 ( .CLK(clk_bF_buf52), .D(_6851__27_), .Q(datapath_1_A_27_) );
DFFPOSX1 DFFPOSX1_1085 ( .CLK(clk_bF_buf10), .D(_6851__28_), .Q(datapath_1_A_28_) );
DFFPOSX1 DFFPOSX1_1086 ( .CLK(clk_bF_buf10), .D(_6851__29_), .Q(datapath_1_A_29_) );
DFFPOSX1 DFFPOSX1_1087 ( .CLK(clk_bF_buf97), .D(_6851__30_), .Q(datapath_1_A_30_) );
DFFPOSX1 DFFPOSX1_1088 ( .CLK(clk_bF_buf43), .D(_6851__31_), .Q(datapath_1_A_31_) );
NAND2X1 NAND2X1_653 ( .A(datapath_1_RD2_0_), .B(vdd), .Y(_6982_) );
INVX1 INVX1_216 ( .A(vdd), .Y(_6918_) );
NAND2X1 NAND2X1_654 ( .A(_2__0_), .B(_6918__bF_buf0), .Y(_6919_) );
AOI21X1 AOI21X1_377 ( .A(_6919_), .B(_6982_), .C(rst_bF_buf13), .Y(_6917__0_) );
NAND2X1 NAND2X1_655 ( .A(vdd), .B(datapath_1_RD2_1_), .Y(_6920_) );
NAND2X1 NAND2X1_656 ( .A(_2__1_), .B(_6918__bF_buf3), .Y(_6921_) );
AOI21X1 AOI21X1_378 ( .A(_6921_), .B(_6920_), .C(rst_bF_buf8), .Y(_6917__1_) );
NAND2X1 NAND2X1_657 ( .A(vdd), .B(datapath_1_RD2_2_), .Y(_6922_) );
NAND2X1 NAND2X1_658 ( .A(_2__2_), .B(_6918__bF_buf4), .Y(_6923_) );
AOI21X1 AOI21X1_379 ( .A(_6923_), .B(_6922_), .C(rst_bF_buf1), .Y(_6917__2_) );
NAND2X1 NAND2X1_659 ( .A(vdd), .B(datapath_1_RD2_3_), .Y(_6924_) );
NAND2X1 NAND2X1_660 ( .A(_2__3_), .B(_6918__bF_buf4), .Y(_6925_) );
AOI21X1 AOI21X1_380 ( .A(_6925_), .B(_6924_), .C(rst_bF_buf1), .Y(_6917__3_) );
NAND2X1 NAND2X1_661 ( .A(vdd), .B(datapath_1_RD2_4_), .Y(_6926_) );
NAND2X1 NAND2X1_662 ( .A(_2__4_), .B(_6918__bF_buf2), .Y(_6927_) );
AOI21X1 AOI21X1_381 ( .A(_6927_), .B(_6926_), .C(rst_bF_buf8), .Y(_6917__4_) );
NAND2X1 NAND2X1_663 ( .A(vdd), .B(datapath_1_RD2_5_), .Y(_6928_) );
NAND2X1 NAND2X1_664 ( .A(_2__5_), .B(_6918__bF_buf1), .Y(_6929_) );
AOI21X1 AOI21X1_382 ( .A(_6929_), .B(_6928_), .C(rst_bF_buf9), .Y(_6917__5_) );
NAND2X1 NAND2X1_665 ( .A(vdd), .B(datapath_1_RD2_6_), .Y(_6930_) );
NAND2X1 NAND2X1_666 ( .A(_2__6_), .B(_6918__bF_buf2), .Y(_6931_) );
AOI21X1 AOI21X1_383 ( .A(_6931_), .B(_6930_), .C(rst_bF_buf3), .Y(_6917__6_) );
NAND2X1 NAND2X1_667 ( .A(vdd), .B(datapath_1_RD2_7_), .Y(_6932_) );
NAND2X1 NAND2X1_668 ( .A(_2__7_), .B(_6918__bF_buf3), .Y(_6933_) );
AOI21X1 AOI21X1_384 ( .A(_6933_), .B(_6932_), .C(rst_bF_buf1), .Y(_6917__7_) );
NAND2X1 NAND2X1_669 ( .A(vdd), .B(datapath_1_RD2_8_), .Y(_6934_) );
NAND2X1 NAND2X1_670 ( .A(_2__8_), .B(_6918__bF_buf0), .Y(_6935_) );
AOI21X1 AOI21X1_385 ( .A(_6935_), .B(_6934_), .C(rst_bF_buf3), .Y(_6917__8_) );
NAND2X1 NAND2X1_671 ( .A(vdd), .B(datapath_1_RD2_9_), .Y(_6936_) );
NAND2X1 NAND2X1_672 ( .A(_2__9_), .B(_6918__bF_buf2), .Y(_6937_) );
AOI21X1 AOI21X1_386 ( .A(_6937_), .B(_6936_), .C(rst_bF_buf3), .Y(_6917__9_) );
NAND2X1 NAND2X1_673 ( .A(vdd), .B(datapath_1_RD2_10_), .Y(_6938_) );
NAND2X1 NAND2X1_674 ( .A(_2__10_), .B(_6918__bF_buf0), .Y(_6939_) );
AOI21X1 AOI21X1_387 ( .A(_6939_), .B(_6938_), .C(rst_bF_buf3), .Y(_6917__10_) );
NAND2X1 NAND2X1_675 ( .A(vdd), .B(datapath_1_RD2_11_), .Y(_6940_) );
NAND2X1 NAND2X1_676 ( .A(_2__11_), .B(_6918__bF_buf3), .Y(_6941_) );
AOI21X1 AOI21X1_388 ( .A(_6941_), .B(_6940_), .C(rst_bF_buf1), .Y(_6917__11_) );
NAND2X1 NAND2X1_677 ( .A(vdd), .B(datapath_1_RD2_12_), .Y(_6942_) );
NAND2X1 NAND2X1_678 ( .A(_2__12_), .B(_6918__bF_buf3), .Y(_6943_) );
AOI21X1 AOI21X1_389 ( .A(_6943_), .B(_6942_), .C(rst_bF_buf1), .Y(_6917__12_) );
NAND2X1 NAND2X1_679 ( .A(vdd), .B(datapath_1_RD2_13_), .Y(_6944_) );
NAND2X1 NAND2X1_680 ( .A(_2__13_), .B(_6918__bF_buf1), .Y(_6945_) );
AOI21X1 AOI21X1_390 ( .A(_6945_), .B(_6944_), .C(rst_bF_buf9), .Y(_6917__13_) );
NAND2X1 NAND2X1_681 ( .A(vdd), .B(datapath_1_RD2_14_), .Y(_6946_) );
NAND2X1 NAND2X1_682 ( .A(_2__14_), .B(_6918__bF_buf2), .Y(_6947_) );
AOI21X1 AOI21X1_391 ( .A(_6947_), .B(_6946_), .C(rst_bF_buf3), .Y(_6917__14_) );
NAND2X1 NAND2X1_683 ( .A(vdd), .B(datapath_1_RD2_15_), .Y(_6948_) );
NAND2X1 NAND2X1_684 ( .A(_2__15_), .B(_6918__bF_buf4), .Y(_6949_) );
AOI21X1 AOI21X1_392 ( .A(_6949_), .B(_6948_), .C(rst_bF_buf1), .Y(_6917__15_) );
NAND2X1 NAND2X1_685 ( .A(vdd), .B(datapath_1_RD2_16_), .Y(_6950_) );
NAND2X1 NAND2X1_686 ( .A(_2__16_), .B(_6918__bF_buf2), .Y(_6951_) );
AOI21X1 AOI21X1_393 ( .A(_6951_), .B(_6950_), .C(rst_bF_buf8), .Y(_6917__16_) );
NAND2X1 NAND2X1_687 ( .A(vdd), .B(datapath_1_RD2_17_), .Y(_6952_) );
NAND2X1 NAND2X1_688 ( .A(_2__17_), .B(_6918__bF_buf1), .Y(_6953_) );
AOI21X1 AOI21X1_394 ( .A(_6953_), .B(_6952_), .C(rst_bF_buf13), .Y(_6917__17_) );
NAND2X1 NAND2X1_689 ( .A(vdd), .B(datapath_1_RD2_18_), .Y(_6954_) );
NAND2X1 NAND2X1_690 ( .A(_2__18_), .B(_6918__bF_buf0), .Y(_6955_) );
AOI21X1 AOI21X1_395 ( .A(_6955_), .B(_6954_), .C(rst_bF_buf13), .Y(_6917__18_) );
NAND2X1 NAND2X1_691 ( .A(vdd), .B(datapath_1_RD2_19_), .Y(_6956_) );
NAND2X1 NAND2X1_692 ( .A(_2__19_), .B(_6918__bF_buf4), .Y(_6957_) );
AOI21X1 AOI21X1_396 ( .A(_6957_), .B(_6956_), .C(rst_bF_buf1), .Y(_6917__19_) );
NAND2X1 NAND2X1_693 ( .A(vdd), .B(datapath_1_RD2_20_), .Y(_6958_) );
NAND2X1 NAND2X1_694 ( .A(_2__20_), .B(_6918__bF_buf4), .Y(_6959_) );
AOI21X1 AOI21X1_397 ( .A(_6959_), .B(_6958_), .C(rst_bF_buf1), .Y(_6917__20_) );
NAND2X1 NAND2X1_695 ( .A(vdd), .B(datapath_1_RD2_21_), .Y(_6960_) );
NAND2X1 NAND2X1_696 ( .A(_2__21_), .B(_6918__bF_buf3), .Y(_6961_) );
AOI21X1 AOI21X1_398 ( .A(_6961_), .B(_6960_), .C(rst_bF_buf1), .Y(_6917__21_) );
NAND2X1 NAND2X1_697 ( .A(vdd), .B(datapath_1_RD2_22_), .Y(_6962_) );
NAND2X1 NAND2X1_698 ( .A(_2__22_), .B(_6918__bF_buf1), .Y(_6963_) );
AOI21X1 AOI21X1_399 ( .A(_6963_), .B(_6962_), .C(rst_bF_buf13), .Y(_6917__22_) );
NAND2X1 NAND2X1_699 ( .A(vdd), .B(datapath_1_RD2_23_), .Y(_6964_) );
NAND2X1 NAND2X1_700 ( .A(_2__23_), .B(_6918__bF_buf2), .Y(_6965_) );
AOI21X1 AOI21X1_400 ( .A(_6965_), .B(_6964_), .C(rst_bF_buf8), .Y(_6917__23_) );
NAND2X1 NAND2X1_701 ( .A(vdd), .B(datapath_1_RD2_24_), .Y(_6966_) );
NAND2X1 NAND2X1_702 ( .A(_2__24_), .B(_6918__bF_buf4), .Y(_6967_) );
AOI21X1 AOI21X1_401 ( .A(_6967_), .B(_6966_), .C(rst_bF_buf1), .Y(_6917__24_) );
NAND2X1 NAND2X1_703 ( .A(vdd), .B(datapath_1_RD2_25_), .Y(_6968_) );
NAND2X1 NAND2X1_704 ( .A(_2__25_), .B(_6918__bF_buf3), .Y(_6969_) );
AOI21X1 AOI21X1_402 ( .A(_6969_), .B(_6968_), .C(rst_bF_buf8), .Y(_6917__25_) );
NAND2X1 NAND2X1_705 ( .A(vdd), .B(datapath_1_RD2_26_), .Y(_6970_) );
NAND2X1 NAND2X1_706 ( .A(_2__26_), .B(_6918__bF_buf1), .Y(_6971_) );
AOI21X1 AOI21X1_403 ( .A(_6971_), .B(_6970_), .C(rst_bF_buf9), .Y(_6917__26_) );
NAND2X1 NAND2X1_707 ( .A(vdd), .B(datapath_1_RD2_27_), .Y(_6972_) );
NAND2X1 NAND2X1_708 ( .A(_2__27_), .B(_6918__bF_buf0), .Y(_6973_) );
AOI21X1 AOI21X1_404 ( .A(_6973_), .B(_6972_), .C(rst_bF_buf3), .Y(_6917__27_) );
NAND2X1 NAND2X1_709 ( .A(vdd), .B(datapath_1_RD2_28_), .Y(_6974_) );
NAND2X1 NAND2X1_710 ( .A(_2__28_), .B(_6918__bF_buf3), .Y(_6975_) );
AOI21X1 AOI21X1_405 ( .A(_6975_), .B(_6974_), .C(rst_bF_buf1), .Y(_6917__28_) );
NAND2X1 NAND2X1_711 ( .A(vdd), .B(datapath_1_RD2_29_), .Y(_6976_) );
NAND2X1 NAND2X1_712 ( .A(_2__29_), .B(_6918__bF_buf4), .Y(_6977_) );
AOI21X1 AOI21X1_406 ( .A(_6977_), .B(_6976_), .C(rst_bF_buf1), .Y(_6917__29_) );
NAND2X1 NAND2X1_713 ( .A(vdd), .B(datapath_1_RD2_30_), .Y(_6978_) );
NAND2X1 NAND2X1_714 ( .A(_2__30_), .B(_6918__bF_buf0), .Y(_6979_) );
AOI21X1 AOI21X1_407 ( .A(_6979_), .B(_6978_), .C(rst_bF_buf3), .Y(_6917__30_) );
NAND2X1 NAND2X1_715 ( .A(vdd), .B(datapath_1_RD2_31_), .Y(_6980_) );
NAND2X1 NAND2X1_716 ( .A(_2__31_), .B(_6918__bF_buf1), .Y(_6981_) );
AOI21X1 AOI21X1_408 ( .A(_6981_), .B(_6980_), .C(rst_bF_buf13), .Y(_6917__31_) );
DFFPOSX1 DFFPOSX1_1089 ( .CLK(clk_bF_buf97), .D(_6917__0_), .Q(_2__0_) );
DFFPOSX1 DFFPOSX1_1090 ( .CLK(clk_bF_buf65), .D(_6917__1_), .Q(_2__1_) );
DFFPOSX1 DFFPOSX1_1091 ( .CLK(clk_bF_buf83), .D(_6917__2_), .Q(_2__2_) );
DFFPOSX1 DFFPOSX1_1092 ( .CLK(clk_bF_buf95), .D(_6917__3_), .Q(_2__3_) );
DFFPOSX1 DFFPOSX1_1093 ( .CLK(clk_bF_buf104), .D(_6917__4_), .Q(_2__4_) );
DFFPOSX1 DFFPOSX1_1094 ( .CLK(clk_bF_buf43), .D(_6917__5_), .Q(_2__5_) );
DFFPOSX1 DFFPOSX1_1095 ( .CLK(clk_bF_buf57), .D(_6917__6_), .Q(_2__6_) );
DFFPOSX1 DFFPOSX1_1096 ( .CLK(clk_bF_buf83), .D(_6917__7_), .Q(_2__7_) );
DFFPOSX1 DFFPOSX1_1097 ( .CLK(clk_bF_buf104), .D(_6917__8_), .Q(_2__8_) );
DFFPOSX1 DFFPOSX1_1098 ( .CLK(clk_bF_buf52), .D(_6917__9_), .Q(_2__9_) );
DFFPOSX1 DFFPOSX1_1099 ( .CLK(clk_bF_buf52), .D(_6917__10_), .Q(_2__10_) );
DFFPOSX1 DFFPOSX1_1100 ( .CLK(clk_bF_buf83), .D(_6917__11_), .Q(_2__11_) );
DFFPOSX1 DFFPOSX1_1101 ( .CLK(clk_bF_buf83), .D(_6917__12_), .Q(_2__12_) );
DFFPOSX1 DFFPOSX1_1102 ( .CLK(clk_bF_buf97), .D(_6917__13_), .Q(_2__13_) );
DFFPOSX1 DFFPOSX1_1103 ( .CLK(clk_bF_buf104), .D(_6917__14_), .Q(_2__14_) );
DFFPOSX1 DFFPOSX1_1104 ( .CLK(clk_bF_buf95), .D(_6917__15_), .Q(_2__15_) );
DFFPOSX1 DFFPOSX1_1105 ( .CLK(clk_bF_buf104), .D(_6917__16_), .Q(_2__16_) );
DFFPOSX1 DFFPOSX1_1106 ( .CLK(clk_bF_buf52), .D(_6917__17_), .Q(_2__17_) );
DFFPOSX1 DFFPOSX1_1107 ( .CLK(clk_bF_buf97), .D(_6917__18_), .Q(_2__18_) );
DFFPOSX1 DFFPOSX1_1108 ( .CLK(clk_bF_buf83), .D(_6917__19_), .Q(_2__19_) );
DFFPOSX1 DFFPOSX1_1109 ( .CLK(clk_bF_buf95), .D(_6917__20_), .Q(_2__20_) );
DFFPOSX1 DFFPOSX1_1110 ( .CLK(clk_bF_buf83), .D(_6917__21_), .Q(_2__21_) );
DFFPOSX1 DFFPOSX1_1111 ( .CLK(clk_bF_buf52), .D(_6917__22_), .Q(_2__22_) );
DFFPOSX1 DFFPOSX1_1112 ( .CLK(clk_bF_buf104), .D(_6917__23_), .Q(_2__23_) );
DFFPOSX1 DFFPOSX1_1113 ( .CLK(clk_bF_buf83), .D(_6917__24_), .Q(_2__24_) );
DFFPOSX1 DFFPOSX1_1114 ( .CLK(clk_bF_buf10), .D(_6917__25_), .Q(_2__25_) );
DFFPOSX1 DFFPOSX1_1115 ( .CLK(clk_bF_buf88), .D(_6917__26_), .Q(_2__26_) );
DFFPOSX1 DFFPOSX1_1116 ( .CLK(clk_bF_buf52), .D(_6917__27_), .Q(_2__27_) );
DFFPOSX1 DFFPOSX1_1117 ( .CLK(clk_bF_buf83), .D(_6917__28_), .Q(_2__28_) );
DFFPOSX1 DFFPOSX1_1118 ( .CLK(clk_bF_buf83), .D(_6917__29_), .Q(_2__29_) );
DFFPOSX1 DFFPOSX1_1119 ( .CLK(clk_bF_buf104), .D(_6917__30_), .Q(_2__30_) );
DFFPOSX1 DFFPOSX1_1120 ( .CLK(clk_bF_buf52), .D(_6917__31_), .Q(_2__31_) );
NAND2X1 NAND2X1_717 ( .A(MemData[0]), .B(vdd), .Y(_7048_) );
INVX1 INVX1_217 ( .A(vdd), .Y(_6984_) );
NAND2X1 NAND2X1_718 ( .A(datapath_1_Data_0_), .B(_6984__bF_buf3), .Y(_6985_) );
AOI21X1 AOI21X1_409 ( .A(_6985_), .B(_7048_), .C(rst_bF_buf6), .Y(_6983__0_) );
NAND2X1 NAND2X1_719 ( .A(vdd), .B(MemData[1]), .Y(_6986_) );
NAND2X1 NAND2X1_720 ( .A(datapath_1_Data_1_), .B(_6984__bF_buf0), .Y(_6987_) );
AOI21X1 AOI21X1_410 ( .A(_6987_), .B(_6986_), .C(rst_bF_buf12), .Y(_6983__1_) );
NAND2X1 NAND2X1_721 ( .A(vdd), .B(MemData[2]), .Y(_6988_) );
NAND2X1 NAND2X1_722 ( .A(datapath_1_Data_2_), .B(_6984__bF_buf3), .Y(_6989_) );
AOI21X1 AOI21X1_411 ( .A(_6989_), .B(_6988_), .C(rst_bF_buf6), .Y(_6983__2_) );
NAND2X1 NAND2X1_723 ( .A(vdd), .B(MemData[3]), .Y(_6990_) );
NAND2X1 NAND2X1_724 ( .A(datapath_1_Data_3_), .B(_6984__bF_buf2), .Y(_6991_) );
AOI21X1 AOI21X1_412 ( .A(_6991_), .B(_6990_), .C(rst_bF_buf0), .Y(_6983__3_) );
NAND2X1 NAND2X1_725 ( .A(vdd), .B(MemData[4]), .Y(_6992_) );
NAND2X1 NAND2X1_726 ( .A(datapath_1_Data_4_), .B(_6984__bF_buf2), .Y(_6993_) );
AOI21X1 AOI21X1_413 ( .A(_6993_), .B(_6992_), .C(rst_bF_buf10), .Y(_6983__4_) );
NAND2X1 NAND2X1_727 ( .A(vdd), .B(MemData[5]), .Y(_6994_) );
NAND2X1 NAND2X1_728 ( .A(datapath_1_Data_5_), .B(_6984__bF_buf4), .Y(_6995_) );
AOI21X1 AOI21X1_414 ( .A(_6995_), .B(_6994_), .C(rst_bF_buf12), .Y(_6983__5_) );
NAND2X1 NAND2X1_729 ( .A(vdd), .B(MemData[6]), .Y(_6996_) );
NAND2X1 NAND2X1_730 ( .A(datapath_1_Data_6_), .B(_6984__bF_buf0), .Y(_6997_) );
AOI21X1 AOI21X1_415 ( .A(_6997_), .B(_6996_), .C(rst_bF_buf6), .Y(_6983__6_) );
NAND2X1 NAND2X1_731 ( .A(vdd), .B(MemData[7]), .Y(_6998_) );
NAND2X1 NAND2X1_732 ( .A(datapath_1_Data_7_), .B(_6984__bF_buf2), .Y(_6999_) );
AOI21X1 AOI21X1_416 ( .A(_6999_), .B(_6998_), .C(rst_bF_buf12), .Y(_6983__7_) );
NAND2X1 NAND2X1_733 ( .A(vdd), .B(MemData[8]), .Y(_7000_) );
NAND2X1 NAND2X1_734 ( .A(datapath_1_Data_8_), .B(_6984__bF_buf0), .Y(_7001_) );
AOI21X1 AOI21X1_417 ( .A(_7001_), .B(_7000_), .C(rst_bF_buf12), .Y(_6983__8_) );
NAND2X1 NAND2X1_735 ( .A(vdd), .B(MemData[9]), .Y(_7002_) );
NAND2X1 NAND2X1_736 ( .A(datapath_1_Data_9_), .B(_6984__bF_buf4), .Y(_7003_) );
AOI21X1 AOI21X1_418 ( .A(_7003_), .B(_7002_), .C(rst_bF_buf12), .Y(_6983__9_) );
NAND2X1 NAND2X1_737 ( .A(vdd), .B(MemData[10]), .Y(_7004_) );
NAND2X1 NAND2X1_738 ( .A(datapath_1_Data_10_), .B(_6984__bF_buf4), .Y(_7005_) );
AOI21X1 AOI21X1_419 ( .A(_7005_), .B(_7004_), .C(rst_bF_buf12), .Y(_6983__10_) );
NAND2X1 NAND2X1_739 ( .A(vdd), .B(MemData[11]), .Y(_7006_) );
NAND2X1 NAND2X1_740 ( .A(datapath_1_Data_11_), .B(_6984__bF_buf1), .Y(_7007_) );
AOI21X1 AOI21X1_420 ( .A(_7007_), .B(_7006_), .C(rst_bF_buf2), .Y(_6983__11_) );
NAND2X1 NAND2X1_741 ( .A(vdd), .B(MemData[12]), .Y(_7008_) );
NAND2X1 NAND2X1_742 ( .A(datapath_1_Data_12_), .B(_6984__bF_buf1), .Y(_7009_) );
AOI21X1 AOI21X1_421 ( .A(_7009_), .B(_7008_), .C(rst_bF_buf6), .Y(_6983__12_) );
NAND2X1 NAND2X1_743 ( .A(vdd), .B(MemData[13]), .Y(_7010_) );
NAND2X1 NAND2X1_744 ( .A(datapath_1_Data_13_), .B(_6984__bF_buf4), .Y(_7011_) );
AOI21X1 AOI21X1_422 ( .A(_7011_), .B(_7010_), .C(rst_bF_buf12), .Y(_6983__13_) );
NAND2X1 NAND2X1_745 ( .A(vdd), .B(MemData[14]), .Y(_7012_) );
NAND2X1 NAND2X1_746 ( .A(datapath_1_Data_14_), .B(_6984__bF_buf0), .Y(_7013_) );
AOI21X1 AOI21X1_423 ( .A(_7013_), .B(_7012_), .C(rst_bF_buf12), .Y(_6983__14_) );
NAND2X1 NAND2X1_747 ( .A(vdd), .B(MemData[15]), .Y(_7014_) );
NAND2X1 NAND2X1_748 ( .A(datapath_1_Data_15_), .B(_6984__bF_buf2), .Y(_7015_) );
AOI21X1 AOI21X1_424 ( .A(_7015_), .B(_7014_), .C(rst_bF_buf0), .Y(_6983__15_) );
NAND2X1 NAND2X1_749 ( .A(vdd), .B(MemData[16]), .Y(_7016_) );
NAND2X1 NAND2X1_750 ( .A(datapath_1_Data_16_), .B(_6984__bF_buf1), .Y(_7017_) );
AOI21X1 AOI21X1_425 ( .A(_7017_), .B(_7016_), .C(rst_bF_buf6), .Y(_6983__16_) );
NAND2X1 NAND2X1_751 ( .A(vdd), .B(MemData[17]), .Y(_7018_) );
NAND2X1 NAND2X1_752 ( .A(datapath_1_Data_17_), .B(_6984__bF_buf1), .Y(_7019_) );
AOI21X1 AOI21X1_426 ( .A(_7019_), .B(_7018_), .C(rst_bF_buf6), .Y(_6983__17_) );
NAND2X1 NAND2X1_753 ( .A(vdd), .B(MemData[18]), .Y(_7020_) );
NAND2X1 NAND2X1_754 ( .A(datapath_1_Data_18_), .B(_6984__bF_buf1), .Y(_7021_) );
AOI21X1 AOI21X1_427 ( .A(_7021_), .B(_7020_), .C(rst_bF_buf6), .Y(_6983__18_) );
NAND2X1 NAND2X1_755 ( .A(vdd), .B(MemData[19]), .Y(_7022_) );
NAND2X1 NAND2X1_756 ( .A(datapath_1_Data_19_), .B(_6984__bF_buf2), .Y(_7023_) );
AOI21X1 AOI21X1_428 ( .A(_7023_), .B(_7022_), .C(rst_bF_buf0), .Y(_6983__19_) );
NAND2X1 NAND2X1_757 ( .A(vdd), .B(MemData[20]), .Y(_7024_) );
NAND2X1 NAND2X1_758 ( .A(datapath_1_Data_20_), .B(_6984__bF_buf1), .Y(_7025_) );
AOI21X1 AOI21X1_429 ( .A(_7025_), .B(_7024_), .C(rst_bF_buf6), .Y(_6983__20_) );
NAND2X1 NAND2X1_759 ( .A(vdd), .B(MemData[21]), .Y(_7026_) );
NAND2X1 NAND2X1_760 ( .A(datapath_1_Data_21_), .B(_6984__bF_buf3), .Y(_7027_) );
AOI21X1 AOI21X1_430 ( .A(_7027_), .B(_7026_), .C(rst_bF_buf6), .Y(_6983__21_) );
NAND2X1 NAND2X1_761 ( .A(vdd), .B(MemData[22]), .Y(_7028_) );
NAND2X1 NAND2X1_762 ( .A(datapath_1_Data_22_), .B(_6984__bF_buf3), .Y(_7029_) );
AOI21X1 AOI21X1_431 ( .A(_7029_), .B(_7028_), .C(rst_bF_buf6), .Y(_6983__22_) );
NAND2X1 NAND2X1_763 ( .A(vdd), .B(MemData[23]), .Y(_7030_) );
NAND2X1 NAND2X1_764 ( .A(datapath_1_Data_23_), .B(_6984__bF_buf3), .Y(_7031_) );
AOI21X1 AOI21X1_432 ( .A(_7031_), .B(_7030_), .C(rst_bF_buf6), .Y(_6983__23_) );
NAND2X1 NAND2X1_765 ( .A(vdd), .B(MemData[24]), .Y(_7032_) );
NAND2X1 NAND2X1_766 ( .A(datapath_1_Data_24_), .B(_6984__bF_buf3), .Y(_7033_) );
AOI21X1 AOI21X1_433 ( .A(_7033_), .B(_7032_), .C(rst_bF_buf6), .Y(_6983__24_) );
NAND2X1 NAND2X1_767 ( .A(vdd), .B(MemData[25]), .Y(_7034_) );
NAND2X1 NAND2X1_768 ( .A(datapath_1_Data_25_), .B(_6984__bF_buf2), .Y(_7035_) );
AOI21X1 AOI21X1_434 ( .A(_7035_), .B(_7034_), .C(rst_bF_buf2), .Y(_6983__25_) );
NAND2X1 NAND2X1_769 ( .A(vdd), .B(MemData[26]), .Y(_7036_) );
NAND2X1 NAND2X1_770 ( .A(datapath_1_Data_26_), .B(_6984__bF_buf4), .Y(_7037_) );
AOI21X1 AOI21X1_435 ( .A(_7037_), .B(_7036_), .C(rst_bF_buf12), .Y(_6983__26_) );
NAND2X1 NAND2X1_771 ( .A(vdd), .B(MemData[27]), .Y(_7038_) );
NAND2X1 NAND2X1_772 ( .A(datapath_1_Data_27_), .B(_6984__bF_buf4), .Y(_7039_) );
AOI21X1 AOI21X1_436 ( .A(_7039_), .B(_7038_), .C(rst_bF_buf4), .Y(_6983__27_) );
NAND2X1 NAND2X1_773 ( .A(vdd), .B(MemData[28]), .Y(_7040_) );
NAND2X1 NAND2X1_774 ( .A(datapath_1_Data_28_), .B(_6984__bF_buf0), .Y(_7041_) );
AOI21X1 AOI21X1_437 ( .A(_7041_), .B(_7040_), .C(rst_bF_buf6), .Y(_6983__28_) );
NAND2X1 NAND2X1_775 ( .A(vdd), .B(MemData[29]), .Y(_7042_) );
NAND2X1 NAND2X1_776 ( .A(datapath_1_Data_29_), .B(_6984__bF_buf3), .Y(_7043_) );
AOI21X1 AOI21X1_438 ( .A(_7043_), .B(_7042_), .C(rst_bF_buf6), .Y(_6983__29_) );
NAND2X1 NAND2X1_777 ( .A(vdd), .B(MemData[30]), .Y(_7044_) );
NAND2X1 NAND2X1_778 ( .A(datapath_1_Data_30_), .B(_6984__bF_buf0), .Y(_7045_) );
AOI21X1 AOI21X1_439 ( .A(_7045_), .B(_7044_), .C(rst_bF_buf12), .Y(_6983__30_) );
NAND2X1 NAND2X1_779 ( .A(vdd), .B(MemData[31]), .Y(_7046_) );
NAND2X1 NAND2X1_780 ( .A(datapath_1_Data_31_), .B(_6984__bF_buf4), .Y(_7047_) );
AOI21X1 AOI21X1_440 ( .A(_7047_), .B(_7046_), .C(rst_bF_buf4), .Y(_6983__31_) );
DFFPOSX1 DFFPOSX1_1121 ( .CLK(clk_bF_buf27), .D(_6983__0_), .Q(datapath_1_Data_0_) );
DFFPOSX1 DFFPOSX1_1122 ( .CLK(clk_bF_buf8), .D(_6983__1_), .Q(datapath_1_Data_1_) );
DFFPOSX1 DFFPOSX1_1123 ( .CLK(clk_bF_buf8), .D(_6983__2_), .Q(datapath_1_Data_2_) );
DFFPOSX1 DFFPOSX1_1124 ( .CLK(clk_bF_buf8), .D(_6983__3_), .Q(datapath_1_Data_3_) );
DFFPOSX1 DFFPOSX1_1125 ( .CLK(clk_bF_buf8), .D(_6983__4_), .Q(datapath_1_Data_4_) );
DFFPOSX1 DFFPOSX1_1126 ( .CLK(clk_bF_buf18), .D(_6983__5_), .Q(datapath_1_Data_5_) );
DFFPOSX1 DFFPOSX1_1127 ( .CLK(clk_bF_buf8), .D(_6983__6_), .Q(datapath_1_Data_6_) );
DFFPOSX1 DFFPOSX1_1128 ( .CLK(clk_bF_buf8), .D(_6983__7_), .Q(datapath_1_Data_7_) );
DFFPOSX1 DFFPOSX1_1129 ( .CLK(clk_bF_buf27), .D(_6983__8_), .Q(datapath_1_Data_8_) );
DFFPOSX1 DFFPOSX1_1130 ( .CLK(clk_bF_buf18), .D(_6983__9_), .Q(datapath_1_Data_9_) );
DFFPOSX1 DFFPOSX1_1131 ( .CLK(clk_bF_buf18), .D(_6983__10_), .Q(datapath_1_Data_10_) );
DFFPOSX1 DFFPOSX1_1132 ( .CLK(clk_bF_buf4), .D(_6983__11_), .Q(datapath_1_Data_11_) );
DFFPOSX1 DFFPOSX1_1133 ( .CLK(clk_bF_buf8), .D(_6983__12_), .Q(datapath_1_Data_12_) );
DFFPOSX1 DFFPOSX1_1134 ( .CLK(clk_bF_buf18), .D(_6983__13_), .Q(datapath_1_Data_13_) );
DFFPOSX1 DFFPOSX1_1135 ( .CLK(clk_bF_buf8), .D(_6983__14_), .Q(datapath_1_Data_14_) );
DFFPOSX1 DFFPOSX1_1136 ( .CLK(clk_bF_buf24), .D(_6983__15_), .Q(datapath_1_Data_15_) );
DFFPOSX1 DFFPOSX1_1137 ( .CLK(clk_bF_buf9), .D(_6983__16_), .Q(datapath_1_Data_16_) );
DFFPOSX1 DFFPOSX1_1138 ( .CLK(clk_bF_buf9), .D(_6983__17_), .Q(datapath_1_Data_17_) );
DFFPOSX1 DFFPOSX1_1139 ( .CLK(clk_bF_buf27), .D(_6983__18_), .Q(datapath_1_Data_18_) );
DFFPOSX1 DFFPOSX1_1140 ( .CLK(clk_bF_buf8), .D(_6983__19_), .Q(datapath_1_Data_19_) );
DFFPOSX1 DFFPOSX1_1141 ( .CLK(clk_bF_buf4), .D(_6983__20_), .Q(datapath_1_Data_20_) );
DFFPOSX1 DFFPOSX1_1142 ( .CLK(clk_bF_buf27), .D(_6983__21_), .Q(datapath_1_Data_21_) );
DFFPOSX1 DFFPOSX1_1143 ( .CLK(clk_bF_buf9), .D(_6983__22_), .Q(datapath_1_Data_22_) );
DFFPOSX1 DFFPOSX1_1144 ( .CLK(clk_bF_buf9), .D(_6983__23_), .Q(datapath_1_Data_23_) );
DFFPOSX1 DFFPOSX1_1145 ( .CLK(clk_bF_buf9), .D(_6983__24_), .Q(datapath_1_Data_24_) );
DFFPOSX1 DFFPOSX1_1146 ( .CLK(clk_bF_buf8), .D(_6983__25_), .Q(datapath_1_Data_25_) );
DFFPOSX1 DFFPOSX1_1147 ( .CLK(clk_bF_buf18), .D(_6983__26_), .Q(datapath_1_Data_26_) );
DFFPOSX1 DFFPOSX1_1148 ( .CLK(clk_bF_buf18), .D(_6983__27_), .Q(datapath_1_Data_27_) );
DFFPOSX1 DFFPOSX1_1149 ( .CLK(clk_bF_buf27), .D(_6983__28_), .Q(datapath_1_Data_28_) );
DFFPOSX1 DFFPOSX1_1150 ( .CLK(clk_bF_buf27), .D(_6983__29_), .Q(datapath_1_Data_29_) );
DFFPOSX1 DFFPOSX1_1151 ( .CLK(clk_bF_buf27), .D(_6983__30_), .Q(datapath_1_Data_30_) );
DFFPOSX1 DFFPOSX1_1152 ( .CLK(clk_bF_buf68), .D(_6983__31_), .Q(datapath_1_Data_31_) );
NAND2X1 NAND2X1_781 ( .A(MemData[0]), .B(IRWrite_bF_buf4), .Y(_7114_) );
INVX1 INVX1_218 ( .A(IRWrite_bF_buf0), .Y(_7050_) );
NAND2X1 NAND2X1_782 ( .A(aluControl_1_inst_0_), .B(_7050__bF_buf0), .Y(_7051_) );
AOI21X1 AOI21X1_441 ( .A(_7051_), .B(_7114_), .C(rst_bF_buf12), .Y(_7049__0_) );
NAND2X1 NAND2X1_783 ( .A(IRWrite_bF_buf3), .B(MemData[1]), .Y(_7052_) );
NAND2X1 NAND2X1_784 ( .A(aluControl_1_inst_1_), .B(_7050__bF_buf2), .Y(_7053_) );
AOI21X1 AOI21X1_442 ( .A(_7053_), .B(_7052_), .C(rst_bF_buf0), .Y(_7049__1_) );
NAND2X1 NAND2X1_785 ( .A(IRWrite_bF_buf4), .B(MemData[2]), .Y(_7054_) );
NAND2X1 NAND2X1_786 ( .A(aluControl_1_inst_2_), .B(_7050__bF_buf0), .Y(_7055_) );
AOI21X1 AOI21X1_443 ( .A(_7055_), .B(_7054_), .C(rst_bF_buf12), .Y(_7049__2_) );
NAND2X1 NAND2X1_787 ( .A(IRWrite_bF_buf4), .B(MemData[3]), .Y(_7056_) );
NAND2X1 NAND2X1_788 ( .A(aluControl_1_inst_3_), .B(_7050__bF_buf0), .Y(_7057_) );
AOI21X1 AOI21X1_444 ( .A(_7057_), .B(_7056_), .C(rst_bF_buf12), .Y(_7049__3_) );
NAND2X1 NAND2X1_789 ( .A(IRWrite_bF_buf0), .B(MemData[4]), .Y(_7058_) );
NAND2X1 NAND2X1_790 ( .A(aluControl_1_inst_4_), .B(_7050__bF_buf2), .Y(_7059_) );
AOI21X1 AOI21X1_445 ( .A(_7059_), .B(_7058_), .C(rst_bF_buf10), .Y(_7049__4_) );
NAND2X1 NAND2X1_791 ( .A(IRWrite_bF_buf3), .B(MemData[5]), .Y(_7060_) );
NAND2X1 NAND2X1_792 ( .A(aluControl_1_inst_5_), .B(_7050__bF_buf2), .Y(_7061_) );
AOI21X1 AOI21X1_446 ( .A(_7061_), .B(_7060_), .C(rst_bF_buf0), .Y(_7049__5_) );
NAND2X1 NAND2X1_793 ( .A(IRWrite_bF_buf4), .B(MemData[6]), .Y(_7062_) );
NAND2X1 NAND2X1_794 ( .A(datapath_1_Instr_6_), .B(_7050__bF_buf0), .Y(_7063_) );
AOI21X1 AOI21X1_447 ( .A(_7063_), .B(_7062_), .C(rst_bF_buf12), .Y(_7049__6_) );
NAND2X1 NAND2X1_795 ( .A(IRWrite_bF_buf0), .B(MemData[7]), .Y(_7064_) );
NAND2X1 NAND2X1_796 ( .A(datapath_1_Instr_7_), .B(_7050__bF_buf4), .Y(_7065_) );
AOI21X1 AOI21X1_448 ( .A(_7065_), .B(_7064_), .C(rst_bF_buf10), .Y(_7049__7_) );
NAND2X1 NAND2X1_797 ( .A(IRWrite_bF_buf4), .B(MemData[8]), .Y(_7066_) );
NAND2X1 NAND2X1_798 ( .A(datapath_1_Instr_8_), .B(_7050__bF_buf0), .Y(_7067_) );
AOI21X1 AOI21X1_449 ( .A(_7067_), .B(_7066_), .C(rst_bF_buf12), .Y(_7049__8_) );
NAND2X1 NAND2X1_799 ( .A(IRWrite_bF_buf4), .B(MemData[9]), .Y(_7068_) );
NAND2X1 NAND2X1_800 ( .A(datapath_1_Instr_9_), .B(_7050__bF_buf0), .Y(_7069_) );
AOI21X1 AOI21X1_450 ( .A(_7069_), .B(_7068_), .C(rst_bF_buf4), .Y(_7049__9_) );
NAND2X1 NAND2X1_801 ( .A(IRWrite_bF_buf1), .B(MemData[10]), .Y(_7070_) );
NAND2X1 NAND2X1_802 ( .A(datapath_1_Instr_10_), .B(_7050__bF_buf2), .Y(_7071_) );
AOI21X1 AOI21X1_451 ( .A(_7071_), .B(_7070_), .C(rst_bF_buf4), .Y(_7049__10_) );
NAND2X1 NAND2X1_803 ( .A(IRWrite_bF_buf3), .B(MemData[11]), .Y(_7072_) );
NAND2X1 NAND2X1_804 ( .A(datapath_1_Instr_11_), .B(_7050__bF_buf3), .Y(_7073_) );
AOI21X1 AOI21X1_452 ( .A(_7073_), .B(_7072_), .C(rst_bF_buf2), .Y(_7049__11_) );
NAND2X1 NAND2X1_805 ( .A(IRWrite_bF_buf3), .B(MemData[12]), .Y(_7074_) );
NAND2X1 NAND2X1_806 ( .A(datapath_1_Instr_12_), .B(_7050__bF_buf2), .Y(_7075_) );
AOI21X1 AOI21X1_453 ( .A(_7075_), .B(_7074_), .C(rst_bF_buf0), .Y(_7049__12_) );
NAND2X1 NAND2X1_807 ( .A(IRWrite_bF_buf0), .B(MemData[13]), .Y(_7076_) );
NAND2X1 NAND2X1_808 ( .A(datapath_1_Instr_13_), .B(_7050__bF_buf2), .Y(_7077_) );
AOI21X1 AOI21X1_454 ( .A(_7077_), .B(_7076_), .C(rst_bF_buf10), .Y(_7049__13_) );
NAND2X1 NAND2X1_809 ( .A(IRWrite_bF_buf0), .B(MemData[14]), .Y(_7078_) );
NAND2X1 NAND2X1_810 ( .A(datapath_1_Instr_14_), .B(_7050__bF_buf4), .Y(_7079_) );
AOI21X1 AOI21X1_455 ( .A(_7079_), .B(_7078_), .C(rst_bF_buf10), .Y(_7049__14_) );
NAND2X1 NAND2X1_811 ( .A(IRWrite_bF_buf0), .B(MemData[15]), .Y(_7080_) );
NAND2X1 NAND2X1_812 ( .A(datapath_1_Instr_15_bF_buf0_), .B(_7050__bF_buf4), .Y(_7081_) );
AOI21X1 AOI21X1_456 ( .A(_7081_), .B(_7080_), .C(rst_bF_buf13), .Y(_7049__15_) );
NAND2X1 NAND2X1_813 ( .A(IRWrite_bF_buf2), .B(MemData[16]), .Y(_7082_) );
NAND2X1 NAND2X1_814 ( .A(datapath_1_Instr_16_bF_buf48_), .B(_7050__bF_buf3), .Y(_7083_) );
AOI21X1 AOI21X1_457 ( .A(_7083_), .B(_7082_), .C(rst_bF_buf2), .Y(_7049__16_) );
NAND2X1 NAND2X1_815 ( .A(IRWrite_bF_buf2), .B(MemData[17]), .Y(_7084_) );
NAND2X1 NAND2X1_816 ( .A(datapath_1_Instr_17_bF_buf8_), .B(_7050__bF_buf3), .Y(_7085_) );
AOI21X1 AOI21X1_458 ( .A(_7085_), .B(_7084_), .C(rst_bF_buf2), .Y(_7049__17_) );
NAND2X1 NAND2X1_817 ( .A(IRWrite_bF_buf2), .B(MemData[18]), .Y(_7086_) );
NAND2X1 NAND2X1_818 ( .A(datapath_1_Instr_18_bF_buf1_), .B(_7050__bF_buf3), .Y(_7087_) );
AOI21X1 AOI21X1_459 ( .A(_7087_), .B(_7086_), .C(rst_bF_buf2), .Y(_7049__18_) );
NAND2X1 NAND2X1_819 ( .A(IRWrite_bF_buf3), .B(MemData[19]), .Y(_7088_) );
NAND2X1 NAND2X1_820 ( .A(datapath_1_Instr_19_bF_buf4_), .B(_7050__bF_buf3), .Y(_7089_) );
AOI21X1 AOI21X1_460 ( .A(_7089_), .B(_7088_), .C(rst_bF_buf2), .Y(_7049__19_) );
NAND2X1 NAND2X1_821 ( .A(IRWrite_bF_buf2), .B(MemData[20]), .Y(_7090_) );
NAND2X1 NAND2X1_822 ( .A(datapath_1_Instr_20_bF_buf3_), .B(_7050__bF_buf4), .Y(_7091_) );
AOI21X1 AOI21X1_461 ( .A(_7091_), .B(_7090_), .C(rst_bF_buf2), .Y(_7049__20_) );
NAND2X1 NAND2X1_823 ( .A(IRWrite_bF_buf3), .B(MemData[21]), .Y(_7092_) );
NAND2X1 NAND2X1_824 ( .A(datapath_1_Instr_21_bF_buf54_), .B(_7050__bF_buf4), .Y(_7093_) );
AOI21X1 AOI21X1_462 ( .A(_7093_), .B(_7092_), .C(rst_bF_buf2), .Y(_7049__21_) );
NAND2X1 NAND2X1_825 ( .A(IRWrite_bF_buf2), .B(MemData[22]), .Y(_7094_) );
NAND2X1 NAND2X1_826 ( .A(datapath_1_Instr_22_bF_buf49_), .B(_7050__bF_buf3), .Y(_7095_) );
AOI21X1 AOI21X1_463 ( .A(_7095_), .B(_7094_), .C(rst_bF_buf2), .Y(_7049__22_) );
NAND2X1 NAND2X1_827 ( .A(IRWrite_bF_buf2), .B(MemData[23]), .Y(_7096_) );
NAND2X1 NAND2X1_828 ( .A(datapath_1_Instr_23_bF_buf14_bF_buf3_), .B(_7050__bF_buf3), .Y(_7097_) );
AOI21X1 AOI21X1_464 ( .A(_7097_), .B(_7096_), .C(rst_bF_buf2), .Y(_7049__23_) );
NAND2X1 NAND2X1_829 ( .A(IRWrite_bF_buf2), .B(MemData[24]), .Y(_7098_) );
NAND2X1 NAND2X1_830 ( .A(datapath_1_Instr_24_bF_buf5_), .B(_7050__bF_buf4), .Y(_7099_) );
AOI21X1 AOI21X1_465 ( .A(_7099_), .B(_7098_), .C(rst_bF_buf2), .Y(_7049__24_) );
NAND2X1 NAND2X1_831 ( .A(IRWrite_bF_buf3), .B(MemData[25]), .Y(_7100_) );
NAND2X1 NAND2X1_832 ( .A(datapath_1_Instr_25_bF_buf4_), .B(_7050__bF_buf4), .Y(_7101_) );
AOI21X1 AOI21X1_466 ( .A(_7101_), .B(_7100_), .C(rst_bF_buf2), .Y(_7049__25_) );
NAND2X1 NAND2X1_833 ( .A(IRWrite_bF_buf1), .B(MemData[26]), .Y(_7102_) );
NAND2X1 NAND2X1_834 ( .A(control_1_op_0_), .B(_7050__bF_buf1), .Y(_7103_) );
AOI21X1 AOI21X1_467 ( .A(_7103_), .B(_7102_), .C(rst_bF_buf4), .Y(_7049__26_) );
NAND2X1 NAND2X1_835 ( .A(IRWrite_bF_buf1), .B(MemData[27]), .Y(_7104_) );
NAND2X1 NAND2X1_836 ( .A(control_1_op_1_), .B(_7050__bF_buf1), .Y(_7105_) );
AOI21X1 AOI21X1_468 ( .A(_7105_), .B(_7104_), .C(rst_bF_buf4), .Y(_7049__27_) );
NAND2X1 NAND2X1_837 ( .A(IRWrite_bF_buf1), .B(MemData[28]), .Y(_7106_) );
NAND2X1 NAND2X1_838 ( .A(control_1_op_2_), .B(_7050__bF_buf1), .Y(_7107_) );
AOI21X1 AOI21X1_469 ( .A(_7107_), .B(_7106_), .C(rst_bF_buf4), .Y(_7049__28_) );
NAND2X1 NAND2X1_839 ( .A(IRWrite_bF_buf4), .B(MemData[29]), .Y(_7108_) );
NAND2X1 NAND2X1_840 ( .A(control_1_op_3_), .B(_7050__bF_buf1), .Y(_7109_) );
AOI21X1 AOI21X1_470 ( .A(_7109_), .B(_7108_), .C(rst_bF_buf4), .Y(_7049__29_) );
NAND2X1 NAND2X1_841 ( .A(IRWrite_bF_buf1), .B(MemData[30]), .Y(_7110_) );
NAND2X1 NAND2X1_842 ( .A(control_1_op_4_), .B(_7050__bF_buf1), .Y(_7111_) );
AOI21X1 AOI21X1_471 ( .A(_7111_), .B(_7110_), .C(rst_bF_buf4), .Y(_7049__30_) );
NAND2X1 NAND2X1_843 ( .A(IRWrite_bF_buf1), .B(MemData[31]), .Y(_7112_) );
NAND2X1 NAND2X1_844 ( .A(control_1_op_5_), .B(_7050__bF_buf1), .Y(_7113_) );
AOI21X1 AOI21X1_472 ( .A(_7113_), .B(_7112_), .C(rst_bF_buf4), .Y(_7049__31_) );
DFFPOSX1 DFFPOSX1_1153 ( .CLK(clk_bF_buf27), .D(_7049__0_), .Q(aluControl_1_inst_0_) );
DFFPOSX1 DFFPOSX1_1154 ( .CLK(clk_bF_buf18), .D(_7049__1_), .Q(aluControl_1_inst_1_) );
DFFPOSX1 DFFPOSX1_1155 ( .CLK(clk_bF_buf27), .D(_7049__2_), .Q(aluControl_1_inst_2_) );
DFFPOSX1 DFFPOSX1_1156 ( .CLK(clk_bF_buf27), .D(_7049__3_), .Q(aluControl_1_inst_3_) );
DFFPOSX1 DFFPOSX1_1157 ( .CLK(clk_bF_buf24), .D(_7049__4_), .Q(aluControl_1_inst_4_) );
DFFPOSX1 DFFPOSX1_1158 ( .CLK(clk_bF_buf18), .D(_7049__5_), .Q(aluControl_1_inst_5_) );
DFFPOSX1 DFFPOSX1_1159 ( .CLK(clk_bF_buf18), .D(_7049__6_), .Q(datapath_1_Instr_6_) );
DFFPOSX1 DFFPOSX1_1160 ( .CLK(clk_bF_buf24), .D(_7049__7_), .Q(datapath_1_Instr_7_) );
DFFPOSX1 DFFPOSX1_1161 ( .CLK(clk_bF_buf68), .D(_7049__8_), .Q(datapath_1_Instr_8_) );
DFFPOSX1 DFFPOSX1_1162 ( .CLK(clk_bF_buf68), .D(_7049__9_), .Q(datapath_1_Instr_9_) );
DFFPOSX1 DFFPOSX1_1163 ( .CLK(clk_bF_buf24), .D(_7049__10_), .Q(datapath_1_Instr_10_) );
DFFPOSX1 DFFPOSX1_1164 ( .CLK(clk_bF_buf4), .D(_7049__11_), .Q(datapath_1_Instr_11_) );
DFFPOSX1 DFFPOSX1_1165 ( .CLK(clk_bF_buf18), .D(_7049__12_), .Q(datapath_1_Instr_12_) );
DFFPOSX1 DFFPOSX1_1166 ( .CLK(clk_bF_buf24), .D(_7049__13_), .Q(datapath_1_Instr_13_) );
DFFPOSX1 DFFPOSX1_1167 ( .CLK(clk_bF_buf24), .D(_7049__14_), .Q(datapath_1_Instr_14_) );
DFFPOSX1 DFFPOSX1_1168 ( .CLK(clk_bF_buf97), .D(_7049__15_), .Q(datapath_1_Instr_15_) );
DFFPOSX1 DFFPOSX1_1169 ( .CLK(clk_bF_buf4), .D(_7049__16_), .Q(datapath_1_Instr_16_) );
DFFPOSX1 DFFPOSX1_1170 ( .CLK(clk_bF_buf4), .D(_7049__17_), .Q(datapath_1_Instr_17_) );
DFFPOSX1 DFFPOSX1_1171 ( .CLK(clk_bF_buf80), .D(_7049__18_), .Q(datapath_1_Instr_18_) );
DFFPOSX1 DFFPOSX1_1172 ( .CLK(clk_bF_buf4), .D(_7049__19_), .Q(datapath_1_Instr_19_) );
DFFPOSX1 DFFPOSX1_1173 ( .CLK(clk_bF_buf47), .D(_7049__20_), .Q(datapath_1_Instr_20_) );
DFFPOSX1 DFFPOSX1_1174 ( .CLK(clk_bF_buf4), .D(_7049__21_), .Q(datapath_1_Instr_21_) );
DFFPOSX1 DFFPOSX1_1175 ( .CLK(clk_bF_buf4), .D(_7049__22_), .Q(datapath_1_Instr_22_) );
DFFPOSX1 DFFPOSX1_1176 ( .CLK(clk_bF_buf80), .D(_7049__23_), .Q(datapath_1_Instr_23_) );
DFFPOSX1 DFFPOSX1_1177 ( .CLK(clk_bF_buf47), .D(_7049__24_), .Q(datapath_1_Instr_24_) );
DFFPOSX1 DFFPOSX1_1178 ( .CLK(clk_bF_buf47), .D(_7049__25_), .Q(datapath_1_Instr_25_) );
DFFPOSX1 DFFPOSX1_1179 ( .CLK(clk_bF_buf68), .D(_7049__26_), .Q(control_1_op_0_) );
DFFPOSX1 DFFPOSX1_1180 ( .CLK(clk_bF_buf68), .D(_7049__27_), .Q(control_1_op_1_) );
DFFPOSX1 DFFPOSX1_1181 ( .CLK(clk_bF_buf68), .D(_7049__28_), .Q(control_1_op_2_) );
DFFPOSX1 DFFPOSX1_1182 ( .CLK(clk_bF_buf68), .D(_7049__29_), .Q(control_1_op_3_) );
DFFPOSX1 DFFPOSX1_1183 ( .CLK(clk_bF_buf68), .D(_7049__30_), .Q(control_1_op_4_) );
DFFPOSX1 DFFPOSX1_1184 ( .CLK(clk_bF_buf68), .D(_7049__31_), .Q(control_1_op_5_) );
NAND2X1 NAND2X1_845 ( .A(datapath_1_PC_prima_0_), .B(datapath_1_PCEn_bF_buf1), .Y(_7180_) );
INVX1 INVX1_219 ( .A(datapath_1_PCEn_bF_buf0), .Y(_7116_) );
NAND2X1 NAND2X1_846 ( .A(datapath_1_PC_0_), .B(_7116__bF_buf0), .Y(_7117_) );
AOI21X1 AOI21X1_473 ( .A(_7117_), .B(_7180_), .C(rst_bF_buf0), .Y(_7115__0_) );
NAND2X1 NAND2X1_847 ( .A(datapath_1_PCEn_bF_buf1), .B(datapath_1_PC_prima_1_), .Y(_7118_) );
NAND2X1 NAND2X1_848 ( .A(datapath_1_PC_1_), .B(_7116__bF_buf0), .Y(_7119_) );
AOI21X1 AOI21X1_474 ( .A(_7119_), .B(_7118_), .C(rst_bF_buf0), .Y(_7115__1_) );
NAND2X1 NAND2X1_849 ( .A(datapath_1_PCEn_bF_buf1), .B(datapath_1_PC_prima_2_), .Y(_7120_) );
NAND2X1 NAND2X1_850 ( .A(datapath_1_PC_2_), .B(_7116__bF_buf0), .Y(_7121_) );
AOI21X1 AOI21X1_475 ( .A(_7121_), .B(_7120_), .C(rst_bF_buf0), .Y(_7115__2_) );
NAND2X1 NAND2X1_851 ( .A(datapath_1_PCEn_bF_buf0), .B(datapath_1_PC_prima_3_), .Y(_7122_) );
NAND2X1 NAND2X1_852 ( .A(datapath_1_PC_3_), .B(_7116__bF_buf4), .Y(_7123_) );
AOI21X1 AOI21X1_476 ( .A(_7123_), .B(_7122_), .C(rst_bF_buf7), .Y(_7115__3_) );
NAND2X1 NAND2X1_853 ( .A(datapath_1_PCEn_bF_buf0), .B(datapath_1_PC_prima_4_), .Y(_7124_) );
NAND2X1 NAND2X1_854 ( .A(datapath_1_PC_4_), .B(_7116__bF_buf0), .Y(_7125_) );
AOI21X1 AOI21X1_477 ( .A(_7125_), .B(_7124_), .C(rst_bF_buf9), .Y(_7115__4_) );
NAND2X1 NAND2X1_855 ( .A(datapath_1_PCEn_bF_buf4), .B(datapath_1_PC_prima_5_), .Y(_7126_) );
NAND2X1 NAND2X1_856 ( .A(datapath_1_PC_5_), .B(_7116__bF_buf3), .Y(_7127_) );
AOI21X1 AOI21X1_478 ( .A(_7127_), .B(_7126_), .C(rst_bF_buf10), .Y(_7115__5_) );
NAND2X1 NAND2X1_857 ( .A(datapath_1_PCEn_bF_buf4), .B(datapath_1_PC_prima_6_), .Y(_7128_) );
NAND2X1 NAND2X1_858 ( .A(datapath_1_PC_6_), .B(_7116__bF_buf3), .Y(_7129_) );
AOI21X1 AOI21X1_479 ( .A(_7129_), .B(_7128_), .C(rst_bF_buf10), .Y(_7115__6_) );
NAND2X1 NAND2X1_859 ( .A(datapath_1_PCEn_bF_buf1), .B(datapath_1_PC_prima_7_), .Y(_7130_) );
NAND2X1 NAND2X1_860 ( .A(datapath_1_PC_7_), .B(_7116__bF_buf0), .Y(_7131_) );
AOI21X1 AOI21X1_480 ( .A(_7131_), .B(_7130_), .C(rst_bF_buf9), .Y(_7115__7_) );
NAND2X1 NAND2X1_861 ( .A(datapath_1_PCEn_bF_buf4), .B(datapath_1_PC_prima_8_), .Y(_7132_) );
NAND2X1 NAND2X1_862 ( .A(datapath_1_PC_8_), .B(_7116__bF_buf1), .Y(_7133_) );
AOI21X1 AOI21X1_481 ( .A(_7133_), .B(_7132_), .C(rst_bF_buf11), .Y(_7115__8_) );
NAND2X1 NAND2X1_863 ( .A(datapath_1_PCEn_bF_buf3), .B(datapath_1_PC_prima_9_), .Y(_7134_) );
NAND2X1 NAND2X1_864 ( .A(datapath_1_PC_9_), .B(_7116__bF_buf2), .Y(_7135_) );
AOI21X1 AOI21X1_482 ( .A(_7135_), .B(_7134_), .C(rst_bF_buf5), .Y(_7115__9_) );
NAND2X1 NAND2X1_865 ( .A(datapath_1_PCEn_bF_buf3), .B(datapath_1_PC_prima_10_), .Y(_7136_) );
NAND2X1 NAND2X1_866 ( .A(datapath_1_PC_10_), .B(_7116__bF_buf2), .Y(_7137_) );
AOI21X1 AOI21X1_483 ( .A(_7137_), .B(_7136_), .C(rst_bF_buf5), .Y(_7115__10_) );
NAND2X1 NAND2X1_867 ( .A(datapath_1_PCEn_bF_buf2), .B(datapath_1_PC_prima_11_), .Y(_7138_) );
NAND2X1 NAND2X1_868 ( .A(datapath_1_PC_11_), .B(_7116__bF_buf4), .Y(_7139_) );
AOI21X1 AOI21X1_484 ( .A(_7139_), .B(_7138_), .C(rst_bF_buf7), .Y(_7115__11_) );
NAND2X1 NAND2X1_869 ( .A(datapath_1_PCEn_bF_buf2), .B(datapath_1_PC_prima_12_), .Y(_7140_) );
NAND2X1 NAND2X1_870 ( .A(datapath_1_PC_12_), .B(_7116__bF_buf2), .Y(_7141_) );
AOI21X1 AOI21X1_485 ( .A(_7141_), .B(_7140_), .C(rst_bF_buf7), .Y(_7115__12_) );
NAND2X1 NAND2X1_871 ( .A(datapath_1_PCEn_bF_buf2), .B(datapath_1_PC_prima_13_), .Y(_7142_) );
NAND2X1 NAND2X1_872 ( .A(datapath_1_PC_13_), .B(_7116__bF_buf4), .Y(_7143_) );
AOI21X1 AOI21X1_486 ( .A(_7143_), .B(_7142_), .C(rst_bF_buf7), .Y(_7115__13_) );
NAND2X1 NAND2X1_873 ( .A(datapath_1_PCEn_bF_buf4), .B(datapath_1_PC_prima_14_), .Y(_7144_) );
NAND2X1 NAND2X1_874 ( .A(datapath_1_PC_14_), .B(_7116__bF_buf1), .Y(_7145_) );
AOI21X1 AOI21X1_487 ( .A(_7145_), .B(_7144_), .C(rst_bF_buf5), .Y(_7115__14_) );
NAND2X1 NAND2X1_875 ( .A(datapath_1_PCEn_bF_buf4), .B(datapath_1_PC_prima_15_), .Y(_7146_) );
NAND2X1 NAND2X1_876 ( .A(datapath_1_PC_15_), .B(_7116__bF_buf3), .Y(_7147_) );
AOI21X1 AOI21X1_488 ( .A(_7147_), .B(_7146_), .C(rst_bF_buf10), .Y(_7115__15_) );
NAND2X1 NAND2X1_877 ( .A(datapath_1_PCEn_bF_buf0), .B(datapath_1_PC_prima_16_), .Y(_7148_) );
NAND2X1 NAND2X1_878 ( .A(datapath_1_PC_16_), .B(_7116__bF_buf4), .Y(_7149_) );
AOI21X1 AOI21X1_489 ( .A(_7149_), .B(_7148_), .C(rst_bF_buf7), .Y(_7115__16_) );
NAND2X1 NAND2X1_879 ( .A(datapath_1_PCEn_bF_buf0), .B(datapath_1_PC_prima_17_), .Y(_7150_) );
NAND2X1 NAND2X1_880 ( .A(datapath_1_PC_17_), .B(_7116__bF_buf4), .Y(_7151_) );
AOI21X1 AOI21X1_490 ( .A(_7151_), .B(_7150_), .C(rst_bF_buf7), .Y(_7115__17_) );
NAND2X1 NAND2X1_881 ( .A(datapath_1_PCEn_bF_buf3), .B(datapath_1_PC_prima_18_), .Y(_7152_) );
NAND2X1 NAND2X1_882 ( .A(datapath_1_PC_18_), .B(_7116__bF_buf1), .Y(_7153_) );
AOI21X1 AOI21X1_491 ( .A(_7153_), .B(_7152_), .C(rst_bF_buf5), .Y(_7115__18_) );
NAND2X1 NAND2X1_883 ( .A(datapath_1_PCEn_bF_buf0), .B(datapath_1_PC_prima_19_), .Y(_7154_) );
NAND2X1 NAND2X1_884 ( .A(datapath_1_PC_19_), .B(_7116__bF_buf4), .Y(_7155_) );
AOI21X1 AOI21X1_492 ( .A(_7155_), .B(_7154_), .C(rst_bF_buf7), .Y(_7115__19_) );
NAND2X1 NAND2X1_885 ( .A(datapath_1_PCEn_bF_buf4), .B(datapath_1_PC_prima_20_), .Y(_7156_) );
NAND2X1 NAND2X1_886 ( .A(datapath_1_PC_20_), .B(_7116__bF_buf3), .Y(_7157_) );
AOI21X1 AOI21X1_493 ( .A(_7157_), .B(_7156_), .C(rst_bF_buf10), .Y(_7115__20_) );
NAND2X1 NAND2X1_887 ( .A(datapath_1_PCEn_bF_buf1), .B(datapath_1_PC_prima_21_), .Y(_7158_) );
NAND2X1 NAND2X1_888 ( .A(datapath_1_PC_21_), .B(_7116__bF_buf3), .Y(_7159_) );
AOI21X1 AOI21X1_494 ( .A(_7159_), .B(_7158_), .C(rst_bF_buf0), .Y(_7115__21_) );
NAND2X1 NAND2X1_889 ( .A(datapath_1_PCEn_bF_buf2), .B(datapath_1_PC_prima_22_), .Y(_7160_) );
NAND2X1 NAND2X1_890 ( .A(datapath_1_PC_22_), .B(_7116__bF_buf2), .Y(_7161_) );
AOI21X1 AOI21X1_495 ( .A(_7161_), .B(_7160_), .C(rst_bF_buf7), .Y(_7115__22_) );
NAND2X1 NAND2X1_891 ( .A(datapath_1_PCEn_bF_buf2), .B(datapath_1_PC_prima_23_), .Y(_7162_) );
NAND2X1 NAND2X1_892 ( .A(datapath_1_PC_23_), .B(_7116__bF_buf2), .Y(_7163_) );
AOI21X1 AOI21X1_496 ( .A(_7163_), .B(_7162_), .C(rst_bF_buf7), .Y(_7115__23_) );
NAND2X1 NAND2X1_893 ( .A(datapath_1_PCEn_bF_buf3), .B(datapath_1_PC_prima_24_), .Y(_7164_) );
NAND2X1 NAND2X1_894 ( .A(datapath_1_PC_24_), .B(_7116__bF_buf1), .Y(_7165_) );
AOI21X1 AOI21X1_497 ( .A(_7165_), .B(_7164_), .C(rst_bF_buf5), .Y(_7115__24_) );
NAND2X1 NAND2X1_895 ( .A(datapath_1_PCEn_bF_buf1), .B(datapath_1_PC_prima_25_), .Y(_7166_) );
NAND2X1 NAND2X1_896 ( .A(datapath_1_PC_25_), .B(_7116__bF_buf0), .Y(_7167_) );
AOI21X1 AOI21X1_498 ( .A(_7167_), .B(_7166_), .C(rst_bF_buf0), .Y(_7115__25_) );
NAND2X1 NAND2X1_897 ( .A(datapath_1_PCEn_bF_buf3), .B(datapath_1_PC_prima_26_), .Y(_7168_) );
NAND2X1 NAND2X1_898 ( .A(datapath_1_PC_26_), .B(_7116__bF_buf1), .Y(_7169_) );
AOI21X1 AOI21X1_499 ( .A(_7169_), .B(_7168_), .C(rst_bF_buf11), .Y(_7115__26_) );
NAND2X1 NAND2X1_899 ( .A(datapath_1_PCEn_bF_buf4), .B(datapath_1_PC_prima_27_), .Y(_7170_) );
NAND2X1 NAND2X1_900 ( .A(datapath_1_PC_27_), .B(_7116__bF_buf3), .Y(_7171_) );
AOI21X1 AOI21X1_500 ( .A(_7171_), .B(_7170_), .C(rst_bF_buf11), .Y(_7115__27_) );
NAND2X1 NAND2X1_901 ( .A(datapath_1_PCEn_bF_buf3), .B(datapath_1_PC_prima_28_), .Y(_7172_) );
NAND2X1 NAND2X1_902 ( .A(datapath_1_PC_28_), .B(_7116__bF_buf1), .Y(_7173_) );
AOI21X1 AOI21X1_501 ( .A(_7173_), .B(_7172_), .C(rst_bF_buf5), .Y(_7115__28_) );
NAND2X1 NAND2X1_903 ( .A(datapath_1_PCEn_bF_buf2), .B(datapath_1_PC_prima_29_), .Y(_7174_) );
NAND2X1 NAND2X1_904 ( .A(datapath_1_PC_29_), .B(_7116__bF_buf4), .Y(_7175_) );
AOI21X1 AOI21X1_502 ( .A(_7175_), .B(_7174_), .C(rst_bF_buf7), .Y(_7115__29_) );
NAND2X1 NAND2X1_905 ( .A(datapath_1_PCEn_bF_buf2), .B(datapath_1_PC_prima_30_), .Y(_7176_) );
NAND2X1 NAND2X1_906 ( .A(datapath_1_PC_30_), .B(_7116__bF_buf2), .Y(_7177_) );
AOI21X1 AOI21X1_503 ( .A(_7177_), .B(_7176_), .C(rst_bF_buf5), .Y(_7115__30_) );
NAND2X1 NAND2X1_907 ( .A(datapath_1_PCEn_bF_buf3), .B(datapath_1_PC_prima_31_), .Y(_7178_) );
NAND2X1 NAND2X1_908 ( .A(datapath_1_PC_31_), .B(_7116__bF_buf3), .Y(_7179_) );
AOI21X1 AOI21X1_504 ( .A(_7179_), .B(_7178_), .C(rst_bF_buf5), .Y(_7115__31_) );
DFFPOSX1 DFFPOSX1_1185 ( .CLK(clk_bF_buf71), .D(_7115__0_), .Q(datapath_1_PC_0_) );
DFFPOSX1 DFFPOSX1_1186 ( .CLK(clk_bF_buf71), .D(_7115__1_), .Q(datapath_1_PC_1_) );
DFFPOSX1 DFFPOSX1_1187 ( .CLK(clk_bF_buf71), .D(_7115__2_), .Q(datapath_1_PC_2_) );
DFFPOSX1 DFFPOSX1_1188 ( .CLK(clk_bF_buf97), .D(_7115__3_), .Q(datapath_1_PC_3_) );
DFFPOSX1 DFFPOSX1_1189 ( .CLK(clk_bF_buf43), .D(_7115__4_), .Q(datapath_1_PC_4_) );
DFFPOSX1 DFFPOSX1_1190 ( .CLK(clk_bF_buf71), .D(_7115__5_), .Q(datapath_1_PC_5_) );
DFFPOSX1 DFFPOSX1_1191 ( .CLK(clk_bF_buf24), .D(_7115__6_), .Q(datapath_1_PC_6_) );
DFFPOSX1 DFFPOSX1_1192 ( .CLK(clk_bF_buf43), .D(_7115__7_), .Q(datapath_1_PC_7_) );
DFFPOSX1 DFFPOSX1_1193 ( .CLK(clk_bF_buf50), .D(_7115__8_), .Q(datapath_1_PC_8_) );
DFFPOSX1 DFFPOSX1_1194 ( .CLK(clk_bF_buf108), .D(_7115__9_), .Q(datapath_1_PC_9_) );
DFFPOSX1 DFFPOSX1_1195 ( .CLK(clk_bF_buf108), .D(_7115__10_), .Q(datapath_1_PC_10_) );
DFFPOSX1 DFFPOSX1_1196 ( .CLK(clk_bF_buf91), .D(_7115__11_), .Q(datapath_1_PC_11_) );
DFFPOSX1 DFFPOSX1_1197 ( .CLK(clk_bF_buf91), .D(_7115__12_), .Q(datapath_1_PC_12_) );
DFFPOSX1 DFFPOSX1_1198 ( .CLK(clk_bF_buf91), .D(_7115__13_), .Q(datapath_1_PC_13_) );
DFFPOSX1 DFFPOSX1_1199 ( .CLK(clk_bF_buf50), .D(_7115__14_), .Q(datapath_1_PC_14_) );
DFFPOSX1 DFFPOSX1_1200 ( .CLK(clk_bF_buf0), .D(_7115__15_), .Q(datapath_1_PC_15_) );
DFFPOSX1 DFFPOSX1_1201 ( .CLK(clk_bF_buf91), .D(_7115__16_), .Q(datapath_1_PC_16_) );
DFFPOSX1 DFFPOSX1_1202 ( .CLK(clk_bF_buf97), .D(_7115__17_), .Q(datapath_1_PC_17_) );
DFFPOSX1 DFFPOSX1_1203 ( .CLK(clk_bF_buf108), .D(_7115__18_), .Q(datapath_1_PC_18_) );
DFFPOSX1 DFFPOSX1_1204 ( .CLK(clk_bF_buf91), .D(_7115__19_), .Q(datapath_1_PC_19_) );
DFFPOSX1 DFFPOSX1_1205 ( .CLK(clk_bF_buf24), .D(_7115__20_), .Q(datapath_1_PC_20_) );
DFFPOSX1 DFFPOSX1_1206 ( .CLK(clk_bF_buf71), .D(_7115__21_), .Q(datapath_1_PC_21_) );
DFFPOSX1 DFFPOSX1_1207 ( .CLK(clk_bF_buf91), .D(_7115__22_), .Q(datapath_1_PC_22_) );
DFFPOSX1 DFFPOSX1_1208 ( .CLK(clk_bF_buf91), .D(_7115__23_), .Q(datapath_1_PC_23_) );
DFFPOSX1 DFFPOSX1_1209 ( .CLK(clk_bF_buf50), .D(_7115__24_), .Q(datapath_1_PC_24_) );
DFFPOSX1 DFFPOSX1_1210 ( .CLK(clk_bF_buf71), .D(_7115__25_), .Q(datapath_1_PC_25_) );
DFFPOSX1 DFFPOSX1_1211 ( .CLK(clk_bF_buf50), .D(_7115__26_), .Q(datapath_1_PC_26_) );
DFFPOSX1 DFFPOSX1_1212 ( .CLK(clk_bF_buf0), .D(_7115__27_), .Q(datapath_1_PC_27_) );
DFFPOSX1 DFFPOSX1_1213 ( .CLK(clk_bF_buf108), .D(_7115__28_), .Q(datapath_1_PC_28_) );
DFFPOSX1 DFFPOSX1_1214 ( .CLK(clk_bF_buf91), .D(_7115__29_), .Q(datapath_1_PC_29_) );
DFFPOSX1 DFFPOSX1_1215 ( .CLK(clk_bF_buf108), .D(_7115__30_), .Q(datapath_1_PC_30_) );
DFFPOSX1 DFFPOSX1_1216 ( .CLK(clk_bF_buf50), .D(_7115__31_), .Q(datapath_1_PC_31_) );
BUFX2 BUFX2_1297 ( .A(_0__0_), .Y(MemAddr[0]) );
BUFX2 BUFX2_1298 ( .A(_0__1_), .Y(MemAddr[1]) );
BUFX2 BUFX2_1299 ( .A(_0__2_), .Y(MemAddr[2]) );
BUFX2 BUFX2_1300 ( .A(_0__3_), .Y(MemAddr[3]) );
BUFX2 BUFX2_1301 ( .A(_0__4_), .Y(MemAddr[4]) );
BUFX2 BUFX2_1302 ( .A(_0__5_), .Y(MemAddr[5]) );
BUFX2 BUFX2_1303 ( .A(_0__6_), .Y(MemAddr[6]) );
BUFX2 BUFX2_1304 ( .A(_0__7_), .Y(MemAddr[7]) );
BUFX2 BUFX2_1305 ( .A(_0__8_), .Y(MemAddr[8]) );
BUFX2 BUFX2_1306 ( .A(_0__9_), .Y(MemAddr[9]) );
BUFX2 BUFX2_1307 ( .A(_0__10_), .Y(MemAddr[10]) );
BUFX2 BUFX2_1308 ( .A(_0__11_), .Y(MemAddr[11]) );
BUFX2 BUFX2_1309 ( .A(_0__12_), .Y(MemAddr[12]) );
BUFX2 BUFX2_1310 ( .A(_0__13_), .Y(MemAddr[13]) );
BUFX2 BUFX2_1311 ( .A(_0__14_), .Y(MemAddr[14]) );
BUFX2 BUFX2_1312 ( .A(_0__15_), .Y(MemAddr[15]) );
BUFX2 BUFX2_1313 ( .A(_0__16_), .Y(MemAddr[16]) );
BUFX2 BUFX2_1314 ( .A(_0__17_), .Y(MemAddr[17]) );
BUFX2 BUFX2_1315 ( .A(_0__18_), .Y(MemAddr[18]) );
BUFX2 BUFX2_1316 ( .A(_0__19_), .Y(MemAddr[19]) );
BUFX2 BUFX2_1317 ( .A(_0__20_), .Y(MemAddr[20]) );
BUFX2 BUFX2_1318 ( .A(_0__21_), .Y(MemAddr[21]) );
BUFX2 BUFX2_1319 ( .A(_0__22_), .Y(MemAddr[22]) );
BUFX2 BUFX2_1320 ( .A(_0__23_), .Y(MemAddr[23]) );
BUFX2 BUFX2_1321 ( .A(_0__24_), .Y(MemAddr[24]) );
BUFX2 BUFX2_1322 ( .A(_0__25_), .Y(MemAddr[25]) );
BUFX2 BUFX2_1323 ( .A(_0__26_), .Y(MemAddr[26]) );
BUFX2 BUFX2_1324 ( .A(_0__27_), .Y(MemAddr[27]) );
BUFX2 BUFX2_1325 ( .A(_0__28_), .Y(MemAddr[28]) );
BUFX2 BUFX2_1326 ( .A(_0__29_), .Y(MemAddr[29]) );
BUFX2 BUFX2_1327 ( .A(_0__30_), .Y(MemAddr[30]) );
BUFX2 BUFX2_1328 ( .A(_0__31_), .Y(MemAddr[31]) );
BUFX2 BUFX2_1329 ( .A(vdd), .Y(MemRead) );
BUFX2 BUFX2_1330 ( .A(_1_), .Y(MemWrite) );
BUFX2 BUFX2_1331 ( .A(_2__0_), .Y(MemWriteData[0]) );
BUFX2 BUFX2_1332 ( .A(_2__1_), .Y(MemWriteData[1]) );
BUFX2 BUFX2_1333 ( .A(_2__2_), .Y(MemWriteData[2]) );
BUFX2 BUFX2_1334 ( .A(_2__3_), .Y(MemWriteData[3]) );
BUFX2 BUFX2_1335 ( .A(_2__4_), .Y(MemWriteData[4]) );
BUFX2 BUFX2_1336 ( .A(_2__5_), .Y(MemWriteData[5]) );
BUFX2 BUFX2_1337 ( .A(_2__6_), .Y(MemWriteData[6]) );
BUFX2 BUFX2_1338 ( .A(_2__7_), .Y(MemWriteData[7]) );
BUFX2 BUFX2_1339 ( .A(_2__8_), .Y(MemWriteData[8]) );
BUFX2 BUFX2_1340 ( .A(_2__9_), .Y(MemWriteData[9]) );
BUFX2 BUFX2_1341 ( .A(_2__10_), .Y(MemWriteData[10]) );
BUFX2 BUFX2_1342 ( .A(_2__11_), .Y(MemWriteData[11]) );
BUFX2 BUFX2_1343 ( .A(_2__12_), .Y(MemWriteData[12]) );
BUFX2 BUFX2_1344 ( .A(_2__13_), .Y(MemWriteData[13]) );
BUFX2 BUFX2_1345 ( .A(_2__14_), .Y(MemWriteData[14]) );
BUFX2 BUFX2_1346 ( .A(_2__15_), .Y(MemWriteData[15]) );
BUFX2 BUFX2_1347 ( .A(_2__16_), .Y(MemWriteData[16]) );
BUFX2 BUFX2_1348 ( .A(_2__17_), .Y(MemWriteData[17]) );
BUFX2 BUFX2_1349 ( .A(_2__18_), .Y(MemWriteData[18]) );
BUFX2 BUFX2_1350 ( .A(_2__19_), .Y(MemWriteData[19]) );
BUFX2 BUFX2_1351 ( .A(_2__20_), .Y(MemWriteData[20]) );
BUFX2 BUFX2_1352 ( .A(_2__21_), .Y(MemWriteData[21]) );
BUFX2 BUFX2_1353 ( .A(_2__22_), .Y(MemWriteData[22]) );
BUFX2 BUFX2_1354 ( .A(_2__23_), .Y(MemWriteData[23]) );
BUFX2 BUFX2_1355 ( .A(_2__24_), .Y(MemWriteData[24]) );
BUFX2 BUFX2_1356 ( .A(_2__25_), .Y(MemWriteData[25]) );
BUFX2 BUFX2_1357 ( .A(_2__26_), .Y(MemWriteData[26]) );
BUFX2 BUFX2_1358 ( .A(_2__27_), .Y(MemWriteData[27]) );
BUFX2 BUFX2_1359 ( .A(_2__28_), .Y(MemWriteData[28]) );
BUFX2 BUFX2_1360 ( .A(_2__29_), .Y(MemWriteData[29]) );
BUFX2 BUFX2_1361 ( .A(_2__30_), .Y(MemWriteData[30]) );
BUFX2 BUFX2_1362 ( .A(_2__31_), .Y(MemWriteData[31]) );
NAND2X1 NAND2X1_909 ( .A(ALUOp_0_bF_buf0_), .B(ALUOp_1_), .Y(_3_) );
NOR2X1 NOR2X1_144 ( .A(aluControl_1_inst_4_), .B(ALUOp_0_bF_buf5_), .Y(_4_) );
NAND2X1 NAND2X1_910 ( .A(aluControl_1_inst_5_), .B(ALUOp_1_), .Y(_5_) );
INVX1 INVX1_220 ( .A(_5_), .Y(_6_) );
INVX1 INVX1_221 ( .A(aluControl_1_inst_2_), .Y(_7_) );
NOR2X1 NOR2X1_145 ( .A(aluControl_1_inst_3_), .B(_7_), .Y(_8_) );
NAND3X1 NAND3X1_1355 ( .A(_4_), .B(_6_), .C(_8_), .Y(_9_) );
XNOR2X1 XNOR2X1_1 ( .A(aluControl_1_inst_0_), .B(aluControl_1_inst_1_), .Y(_10_) );
OAI21X1 OAI21X1_1418 ( .A(_10_), .B(_9_), .C(_3_), .Y(aluControl_0_) );
NOR3X1 NOR3X1_1 ( .A(aluControl_1_inst_4_), .B(ALUOp_0_bF_buf4_), .C(_5_), .Y(_11_) );
AOI21X1 AOI21X1_505 ( .A(_11_), .B(_8_), .C(ALUOp_0_bF_buf3_), .Y(aluControl_1_) );
NAND2X1 NAND2X1_911 ( .A(_4_), .B(_6_), .Y(_12_) );
INVX1 INVX1_222 ( .A(aluControl_1_inst_1_), .Y(_13_) );
NOR2X1 NOR2X1_146 ( .A(aluControl_1_inst_0_), .B(_13_), .Y(_14_) );
AND2X2 AND2X2_3 ( .A(aluControl_1_inst_0_), .B(aluControl_1_inst_1_), .Y(_15_) );
OAI21X1 OAI21X1_1419 ( .A(_15_), .B(_14_), .C(_8_), .Y(_16_) );
NOR2X1 NOR2X1_147 ( .A(aluControl_1_inst_3_), .B(aluControl_1_inst_2_), .Y(_17_) );
NAND3X1 NAND3X1_1356 ( .A(_14_), .B(_17_), .C(_11_), .Y(_18_) );
OAI21X1 OAI21X1_1420 ( .A(_12_), .B(_16_), .C(_18_), .Y(aluControl_2_) );
INVX1 INVX1_223 ( .A(ALUOp_0_bF_buf2_), .Y(_19_) );
OAI21X1 OAI21X1_1421 ( .A(_12_), .B(_16_), .C(_19_), .Y(aluControl_3_) );
INVX1 INVX1_224 ( .A(control_1_state_3_), .Y(_23_) );
NAND2X1 NAND2X1_912 ( .A(control_1_state_2_), .B(_23_), .Y(_24_) );
NAND2X1 NAND2X1_913 ( .A(control_1_state_1_), .B(control_1_state_0_), .Y(_25_) );
NOR2X1 NOR2X1_148 ( .A(_25_), .B(_24_), .Y(RegDst) );
NOR2X1 NOR2X1_149 ( .A(control_1_state_1_), .B(control_1_state_0_), .Y(_26_) );
INVX1 INVX1_225 ( .A(_26_), .Y(_27_) );
NOR2X1 NOR2X1_150 ( .A(_24_), .B(_27_), .Y(MemtoReg) );
INVX1 INVX1_226 ( .A(control_1_state_1_), .Y(_28_) );
NAND2X1 NAND2X1_914 ( .A(control_1_state_0_), .B(_28_), .Y(_29_) );
NOR2X1 NOR2X1_151 ( .A(_24_), .B(_29_), .Y(_1_) );
INVX1 INVX1_227 ( .A(control_1_state_2_), .Y(_30_) );
NAND2X1 NAND2X1_915 ( .A(_23_), .B(_30_), .Y(_31_) );
OAI22X1 OAI22X1_109 ( .A(control_1_state_1_), .B(_24_), .C(_25_), .D(_31_), .Y(IorD) );
INVX1 INVX1_228 ( .A(control_1_state_0_), .Y(_32_) );
NAND2X1 NAND2X1_916 ( .A(control_1_state_1_), .B(_32_), .Y(_33_) );
NOR2X1 NOR2X1_152 ( .A(control_1_state_1_), .B(_32_), .Y(_34_) );
NOR2X1 NOR2X1_153 ( .A(control_1_state_2_), .B(_23_), .Y(_35_) );
NAND2X1 NAND2X1_917 ( .A(_34_), .B(_35_), .Y(_36_) );
OAI21X1 OAI21X1_1422 ( .A(control_1_state_2_), .B(_33_), .C(_36_), .Y(_37_) );
NOR2X1 NOR2X1_154 ( .A(IorD_bF_buf6), .B(_37_), .Y(_38_) );
NOR2X1 NOR2X1_155 ( .A(_28_), .B(_24_), .Y(_39_) );
INVX1 INVX1_229 ( .A(_35_), .Y(_40_) );
NAND3X1 NAND3X1_1357 ( .A(control_1_state_3_), .B(control_1_state_2_), .C(_26_), .Y(_41_) );
OAI21X1 OAI21X1_1423 ( .A(_27_), .B(_40_), .C(_41_), .Y(PCWriteCond) );
NOR2X1 NOR2X1_156 ( .A(_39_), .B(PCWriteCond), .Y(_42_) );
NAND2X1 NAND2X1_918 ( .A(_38_), .B(_42_), .Y(ALUSrcA) );
NOR2X1 NOR2X1_157 ( .A(RegDst), .B(MemtoReg_bF_buf5), .Y(_43_) );
OAI21X1 OAI21X1_1424 ( .A(_33_), .B(_40_), .C(_43_), .Y(RegWrite) );
NOR2X1 NOR2X1_158 ( .A(_31_), .B(_27_), .Y(IRWrite) );
NOR2X1 NOR2X1_159 ( .A(_25_), .B(_40_), .Y(PCSource_1_) );
OR2X2 OR2X2_3 ( .A(PCSource_1_bF_buf0_), .B(IRWrite_bF_buf0), .Y(PCWrite) );
NOR2X1 NOR2X1_160 ( .A(_29_), .B(_31_), .Y(_44_) );
NOR2X1 NOR2X1_161 ( .A(control_1_op_4_), .B(control_1_op_5_), .Y(_45_) );
INVX1 INVX1_230 ( .A(_45_), .Y(_46_) );
INVX1 INVX1_231 ( .A(control_1_op_0_), .Y(_47_) );
NOR2X1 NOR2X1_162 ( .A(control_1_op_2_), .B(control_1_op_3_), .Y(_48_) );
NAND3X1 NAND3X1_1358 ( .A(_47_), .B(control_1_op_1_), .C(_48_), .Y(_49_) );
INVX1 INVX1_232 ( .A(control_1_op_2_), .Y(_50_) );
NOR2X1 NOR2X1_163 ( .A(control_1_op_0_), .B(control_1_op_1_), .Y(_51_) );
NAND3X1 NAND3X1_1359 ( .A(_50_), .B(control_1_op_3_), .C(_51_), .Y(_52_) );
AOI21X1 AOI21X1_506 ( .A(_49_), .B(_52_), .C(_46_), .Y(_53_) );
AOI21X1 AOI21X1_507 ( .A(_53_), .B(_44_), .C(IRWrite_bF_buf1), .Y(_54_) );
NOR2X1 NOR2X1_164 ( .A(_33_), .B(_31_), .Y(_55_) );
AND2X2 AND2X2_4 ( .A(control_1_op_0_), .B(control_1_op_1_), .Y(_56_) );
INVX1 INVX1_233 ( .A(_56_), .Y(_57_) );
INVX1 INVX1_234 ( .A(control_1_op_4_), .Y(_58_) );
NAND2X1 NAND2X1_919 ( .A(control_1_op_5_), .B(_58_), .Y(_59_) );
NAND3X1 NAND3X1_1360 ( .A(_50_), .B(control_1_op_3_), .C(_56_), .Y(_60_) );
NAND3X1 NAND3X1_1361 ( .A(_58_), .B(control_1_op_5_), .C(_48_), .Y(_61_) );
OAI22X1 OAI22X1_110 ( .A(_57_), .B(_61_), .C(_59_), .D(_60_), .Y(_62_) );
AOI22X1 AOI22X1_118 ( .A(_32_), .B(_39_), .C(_55_), .D(_62_), .Y(_63_) );
AOI21X1 AOI21X1_508 ( .A(_54_), .B(_63_), .C(rst_bF_buf4), .Y(_20__0_) );
NAND3X1 NAND3X1_1362 ( .A(_47_), .B(_45_), .C(_48_), .Y(_64_) );
INVX1 INVX1_235 ( .A(_64_), .Y(_65_) );
OAI21X1 OAI21X1_1425 ( .A(_65_), .B(_62_), .C(_44_), .Y(_66_) );
OAI21X1 OAI21X1_1426 ( .A(_24_), .B(_33_), .C(_36_), .Y(_67_) );
NOR2X1 NOR2X1_165 ( .A(_57_), .B(_61_), .Y(_68_) );
AOI21X1 AOI21X1_509 ( .A(_55_), .B(_68_), .C(_67_), .Y(_69_) );
AOI21X1 AOI21X1_510 ( .A(_66_), .B(_69_), .C(rst_bF_buf4), .Y(_20__1_) );
NOR2X1 NOR2X1_166 ( .A(_59_), .B(_60_), .Y(_70_) );
OAI22X1 OAI22X1_111 ( .A(_24_), .B(_33_), .C(_25_), .D(_31_), .Y(_71_) );
AOI21X1 AOI21X1_511 ( .A(_70_), .B(_55_), .C(_71_), .Y(_72_) );
NOR3X1 NOR3X1_2 ( .A(control_1_op_1_), .B(_29_), .C(_31_), .Y(_73_) );
NOR2X1 NOR2X1_167 ( .A(control_1_op_3_), .B(_50_), .Y(_74_) );
NAND2X1 NAND2X1_920 ( .A(_45_), .B(_74_), .Y(_75_) );
OAI21X1 OAI21X1_1427 ( .A(_47_), .B(_75_), .C(_64_), .Y(_76_) );
NAND2X1 NAND2X1_921 ( .A(_73_), .B(_76_), .Y(_77_) );
AOI21X1 AOI21X1_512 ( .A(_77_), .B(_72_), .C(rst_bF_buf4), .Y(_20__2_) );
NAND2X1 NAND2X1_922 ( .A(_44_), .B(_53_), .Y(_78_) );
INVX1 INVX1_236 ( .A(_75_), .Y(_79_) );
AOI22X1 AOI22X1_119 ( .A(_34_), .B(_35_), .C(_73_), .D(_79_), .Y(_21_) );
AOI21X1 AOI21X1_513 ( .A(_21_), .B(_78_), .C(rst_bF_buf4), .Y(_20__3_) );
NOR2X1 NOR2X1_168 ( .A(_44_), .B(PCSource_1_bF_buf5_), .Y(_22_) );
OAI21X1 OAI21X1_1428 ( .A(_27_), .B(_31_), .C(_22_), .Y(ALUSrcB_0_) );
NAND2X1 NAND2X1_923 ( .A(_22_), .B(_38_), .Y(ALUSrcB_1_) );
OAI21X1 OAI21X1_1429 ( .A(_28_), .B(_24_), .C(_41_), .Y(ALUOp_1_) );
OAI21X1 OAI21X1_1430 ( .A(_27_), .B(_40_), .C(_41_), .Y(ALUOp_0_) );
DFFPOSX1 DFFPOSX1_1217 ( .CLK(clk_bF_buf68), .D(_20__0_), .Q(control_1_state_0_) );
DFFPOSX1 DFFPOSX1_1218 ( .CLK(clk_bF_buf0), .D(_20__1_), .Q(control_1_state_1_) );
DFFPOSX1 DFFPOSX1_1219 ( .CLK(clk_bF_buf68), .D(_20__2_), .Q(control_1_state_2_) );
DFFPOSX1 DFFPOSX1_1220 ( .CLK(clk_bF_buf0), .D(_20__3_), .Q(control_1_state_3_) );
OR2X2 OR2X2_4 ( .A(datapath_1_ALU_aluInA_23_), .B(datapath_1_ALU_aluInB_23_), .Y(_80_) );
NAND2X1 NAND2X1_924 ( .A(datapath_1_ALU_aluInA_23_), .B(datapath_1_ALU_aluInB_23_), .Y(_81_) );
NAND2X1 NAND2X1_925 ( .A(_81_), .B(_80_), .Y(_82_) );
INVX1 INVX1_237 ( .A(_82_), .Y(_83_) );
INVX1 INVX1_238 ( .A(datapath_1_ALU_aluInA_22_), .Y(_84_) );
INVX1 INVX1_239 ( .A(datapath_1_ALU_aluInB_22_), .Y(_85_) );
NAND2X1 NAND2X1_926 ( .A(_84_), .B(_85_), .Y(_86_) );
NAND2X1 NAND2X1_927 ( .A(datapath_1_ALU_aluInA_22_), .B(datapath_1_ALU_aluInB_22_), .Y(_87_) );
NAND2X1 NAND2X1_928 ( .A(_87_), .B(_86_), .Y(_88_) );
INVX1 INVX1_240 ( .A(_88_), .Y(_89_) );
NOR2X1 NOR2X1_169 ( .A(_83_), .B(_89_), .Y(_90_) );
INVX1 INVX1_241 ( .A(datapath_1_ALU_aluInA_20_), .Y(_91_) );
INVX1 INVX1_242 ( .A(datapath_1_ALU_aluInB_20_), .Y(_92_) );
NAND2X1 NAND2X1_929 ( .A(_91_), .B(_92_), .Y(_93_) );
NAND2X1 NAND2X1_930 ( .A(datapath_1_ALU_aluInA_20_), .B(datapath_1_ALU_aluInB_20_), .Y(_94_) );
NAND2X1 NAND2X1_931 ( .A(_94_), .B(_93_), .Y(_95_) );
INVX1 INVX1_243 ( .A(_95_), .Y(_96_) );
INVX1 INVX1_244 ( .A(datapath_1_ALU_aluInA_21_), .Y(_97_) );
INVX1 INVX1_245 ( .A(datapath_1_ALU_aluInB_21_), .Y(_98_) );
NAND2X1 NAND2X1_932 ( .A(_97_), .B(_98_), .Y(_99_) );
NAND2X1 NAND2X1_933 ( .A(datapath_1_ALU_aluInA_21_), .B(datapath_1_ALU_aluInB_21_), .Y(_100_) );
NAND2X1 NAND2X1_934 ( .A(_100_), .B(_99_), .Y(_101_) );
INVX1 INVX1_246 ( .A(_101_), .Y(_102_) );
NOR2X1 NOR2X1_170 ( .A(_96_), .B(_102_), .Y(_103_) );
NAND2X1 NAND2X1_935 ( .A(_90_), .B(_103_), .Y(_104_) );
INVX1 INVX1_247 ( .A(datapath_1_ALU_aluInA_17_), .Y(_105_) );
INVX1 INVX1_248 ( .A(datapath_1_ALU_aluInB_17_), .Y(_106_) );
NAND2X1 NAND2X1_936 ( .A(_105_), .B(_106_), .Y(_107_) );
INVX1 INVX1_249 ( .A(_107_), .Y(_108_) );
NAND2X1 NAND2X1_937 ( .A(datapath_1_ALU_aluInA_17_), .B(datapath_1_ALU_aluInB_17_), .Y(_109_) );
INVX1 INVX1_250 ( .A(_109_), .Y(_110_) );
INVX1 INVX1_251 ( .A(datapath_1_ALU_aluInA_16_), .Y(_111_) );
INVX1 INVX1_252 ( .A(datapath_1_ALU_aluInB_16_), .Y(_112_) );
NAND2X1 NAND2X1_938 ( .A(_111_), .B(_112_), .Y(_113_) );
NAND2X1 NAND2X1_939 ( .A(datapath_1_ALU_aluInA_16_), .B(datapath_1_ALU_aluInB_16_), .Y(_114_) );
NAND2X1 NAND2X1_940 ( .A(_114_), .B(_113_), .Y(_115_) );
OAI21X1 OAI21X1_1431 ( .A(_110_), .B(_108_), .C(_115_), .Y(_116_) );
NOR2X1 NOR2X1_171 ( .A(datapath_1_ALU_aluInA_19_), .B(datapath_1_ALU_aluInB_19_), .Y(_117_) );
AND2X2 AND2X2_5 ( .A(datapath_1_ALU_aluInA_19_), .B(datapath_1_ALU_aluInB_19_), .Y(_118_) );
NOR2X1 NOR2X1_172 ( .A(_117_), .B(_118_), .Y(_119_) );
INVX1 INVX1_253 ( .A(_119_), .Y(_120_) );
NOR2X1 NOR2X1_173 ( .A(datapath_1_ALU_aluInA_18_), .B(datapath_1_ALU_aluInB_18_), .Y(_121_) );
INVX1 INVX1_254 ( .A(datapath_1_ALU_aluInA_18_), .Y(_122_) );
INVX1 INVX1_255 ( .A(datapath_1_ALU_aluInB_18_), .Y(_123_) );
NOR2X1 NOR2X1_174 ( .A(_122_), .B(_123_), .Y(_124_) );
OAI21X1 OAI21X1_1432 ( .A(_121_), .B(_124_), .C(_120_), .Y(_125_) );
OR2X2 OR2X2_5 ( .A(_125_), .B(_116_), .Y(_126_) );
NOR2X1 NOR2X1_175 ( .A(_104_), .B(_126_), .Y(_127_) );
NOR2X1 NOR2X1_176 ( .A(datapath_1_ALU_aluInA_27_), .B(datapath_1_ALU_aluInB_27_), .Y(_128_) );
NAND2X1 NAND2X1_941 ( .A(datapath_1_ALU_aluInA_27_), .B(datapath_1_ALU_aluInB_27_), .Y(_129_) );
INVX1 INVX1_256 ( .A(_129_), .Y(_130_) );
NOR2X1 NOR2X1_177 ( .A(_128_), .B(_130_), .Y(_131_) );
NOR2X1 NOR2X1_178 ( .A(datapath_1_ALU_aluInA_26_), .B(datapath_1_ALU_aluInB_26_), .Y(_132_) );
INVX1 INVX1_257 ( .A(datapath_1_ALU_aluInA_26_), .Y(_133_) );
INVX1 INVX1_258 ( .A(datapath_1_ALU_aluInB_26_), .Y(_134_) );
NOR2X1 NOR2X1_179 ( .A(_133_), .B(_134_), .Y(_135_) );
NOR2X1 NOR2X1_180 ( .A(_132_), .B(_135_), .Y(_136_) );
NOR2X1 NOR2X1_181 ( .A(_131_), .B(_136_), .Y(_137_) );
NOR2X1 NOR2X1_182 ( .A(datapath_1_ALU_aluInA_24_), .B(datapath_1_ALU_aluInB_24_), .Y(_138_) );
NAND2X1 NAND2X1_942 ( .A(datapath_1_ALU_aluInA_24_), .B(datapath_1_ALU_aluInB_24_), .Y(_139_) );
INVX1 INVX1_259 ( .A(_139_), .Y(_140_) );
INVX1 INVX1_260 ( .A(datapath_1_ALU_aluInB_25_), .Y(_141_) );
NOR2X1 NOR2X1_183 ( .A(datapath_1_ALU_aluInA_25_), .B(_141_), .Y(_142_) );
INVX1 INVX1_261 ( .A(datapath_1_ALU_aluInA_25_), .Y(_143_) );
NOR2X1 NOR2X1_184 ( .A(datapath_1_ALU_aluInB_25_), .B(_143_), .Y(_144_) );
NOR2X1 NOR2X1_185 ( .A(_142_), .B(_144_), .Y(_145_) );
OAI21X1 OAI21X1_1433 ( .A(_138_), .B(_140_), .C(_145_), .Y(_146_) );
INVX1 INVX1_262 ( .A(_146_), .Y(_147_) );
NAND2X1 NAND2X1_943 ( .A(_137_), .B(_147_), .Y(_148_) );
NOR2X1 NOR2X1_186 ( .A(datapath_1_ALU_aluInA_30_), .B(datapath_1_ALU_aluInB_30_), .Y(_149_) );
INVX1 INVX1_263 ( .A(datapath_1_ALU_aluInA_30_), .Y(_150_) );
INVX1 INVX1_264 ( .A(datapath_1_ALU_aluInB_30_), .Y(_151_) );
NOR2X1 NOR2X1_187 ( .A(_150_), .B(_151_), .Y(_152_) );
NOR2X1 NOR2X1_188 ( .A(_149_), .B(_152_), .Y(_153_) );
INVX1 INVX1_265 ( .A(_153_), .Y(_154_) );
NOR2X1 NOR2X1_189 ( .A(datapath_1_ALU_aluInA_31_), .B(datapath_1_ALU_aluInB_31_), .Y(_155_) );
NAND2X1 NAND2X1_944 ( .A(datapath_1_ALU_aluInA_31_), .B(datapath_1_ALU_aluInB_31_), .Y(_156_) );
INVX1 INVX1_266 ( .A(_156_), .Y(_157_) );
NOR2X1 NOR2X1_190 ( .A(_155_), .B(_157_), .Y(_158_) );
INVX1 INVX1_267 ( .A(_158_), .Y(_159_) );
NOR2X1 NOR2X1_191 ( .A(datapath_1_ALU_aluInA_29_), .B(datapath_1_ALU_aluInB_29_), .Y(_160_) );
NAND2X1 NAND2X1_945 ( .A(datapath_1_ALU_aluInA_29_), .B(datapath_1_ALU_aluInB_29_), .Y(_161_) );
INVX1 INVX1_268 ( .A(_161_), .Y(_162_) );
NOR2X1 NOR2X1_192 ( .A(_160_), .B(_162_), .Y(_163_) );
INVX1 INVX1_269 ( .A(_163_), .Y(_164_) );
NOR2X1 NOR2X1_193 ( .A(datapath_1_ALU_aluInA_28_), .B(datapath_1_ALU_aluInB_28_), .Y(_165_) );
INVX1 INVX1_270 ( .A(datapath_1_ALU_aluInA_28_), .Y(_166_) );
INVX1 INVX1_271 ( .A(datapath_1_ALU_aluInB_28_), .Y(_167_) );
NOR2X1 NOR2X1_194 ( .A(_166_), .B(_167_), .Y(_168_) );
OAI21X1 OAI21X1_1434 ( .A(_165_), .B(_168_), .C(_164_), .Y(_169_) );
INVX1 INVX1_272 ( .A(_169_), .Y(_170_) );
NAND3X1 NAND3X1_1363 ( .A(_154_), .B(_159_), .C(_170_), .Y(_171_) );
NOR2X1 NOR2X1_195 ( .A(_148_), .B(_171_), .Y(_172_) );
NOR2X1 NOR2X1_196 ( .A(datapath_1_ALU_aluInA_15_), .B(datapath_1_ALU_aluInB_15_), .Y(_173_) );
AND2X2 AND2X2_6 ( .A(datapath_1_ALU_aluInA_15_), .B(datapath_1_ALU_aluInB_15_), .Y(_174_) );
NOR2X1 NOR2X1_197 ( .A(_173_), .B(_174_), .Y(_175_) );
NOR2X1 NOR2X1_198 ( .A(datapath_1_ALU_aluInA_14_), .B(datapath_1_ALU_aluInB_14_), .Y(_176_) );
AND2X2 AND2X2_7 ( .A(datapath_1_ALU_aluInA_14_), .B(datapath_1_ALU_aluInB_14_), .Y(_177_) );
NOR2X1 NOR2X1_199 ( .A(_176_), .B(_177_), .Y(_178_) );
NOR2X1 NOR2X1_200 ( .A(_175_), .B(_178_), .Y(_179_) );
NOR2X1 NOR2X1_201 ( .A(datapath_1_ALU_aluInA_12_), .B(datapath_1_ALU_aluInB_12_), .Y(_180_) );
AND2X2 AND2X2_8 ( .A(datapath_1_ALU_aluInA_12_), .B(datapath_1_ALU_aluInB_12_), .Y(_181_) );
NOR2X1 NOR2X1_202 ( .A(_180_), .B(_181_), .Y(_182_) );
NOR2X1 NOR2X1_203 ( .A(datapath_1_ALU_aluInA_13_), .B(datapath_1_ALU_aluInB_13_), .Y(_183_) );
AND2X2 AND2X2_9 ( .A(datapath_1_ALU_aluInA_13_), .B(datapath_1_ALU_aluInB_13_), .Y(_184_) );
NOR2X1 NOR2X1_204 ( .A(_183_), .B(_184_), .Y(_185_) );
NOR2X1 NOR2X1_205 ( .A(_182_), .B(_185_), .Y(_186_) );
INVX1 INVX1_273 ( .A(datapath_1_ALU_aluInA_9_), .Y(_187_) );
INVX1 INVX1_274 ( .A(datapath_1_ALU_aluInB_9_), .Y(_188_) );
NAND2X1 NAND2X1_946 ( .A(_187_), .B(_188_), .Y(_189_) );
NAND2X1 NAND2X1_947 ( .A(datapath_1_ALU_aluInA_9_), .B(datapath_1_ALU_aluInB_9_), .Y(_190_) );
NAND2X1 NAND2X1_948 ( .A(_190_), .B(_189_), .Y(_191_) );
NOR2X1 NOR2X1_206 ( .A(datapath_1_ALU_aluInA_8_), .B(datapath_1_ALU_aluInB_8_), .Y(_192_) );
NAND2X1 NAND2X1_949 ( .A(datapath_1_ALU_aluInA_8_), .B(datapath_1_ALU_aluInB_8_), .Y(_193_) );
INVX1 INVX1_275 ( .A(_193_), .Y(_194_) );
OAI21X1 OAI21X1_1435 ( .A(_192_), .B(_194_), .C(_191_), .Y(_195_) );
XNOR2X1 XNOR2X1_2 ( .A(datapath_1_ALU_aluInA_10_), .B(datapath_1_ALU_aluInB_10_), .Y(_196_) );
NOR2X1 NOR2X1_207 ( .A(datapath_1_ALU_aluInA_11_), .B(datapath_1_ALU_aluInB_11_), .Y(_197_) );
AND2X2 AND2X2_10 ( .A(datapath_1_ALU_aluInA_11_), .B(datapath_1_ALU_aluInB_11_), .Y(_198_) );
OAI21X1 OAI21X1_1436 ( .A(_197_), .B(_198_), .C(_196_), .Y(_199_) );
NOR2X1 NOR2X1_208 ( .A(_199_), .B(_195_), .Y(_200_) );
NAND3X1 NAND3X1_1364 ( .A(_179_), .B(_186_), .C(_200_), .Y(_201_) );
XOR2X1 XOR2X1_1 ( .A(datapath_1_ALU_aluInA_2_), .B(datapath_1_ALU_aluInB_2_), .Y(_202_) );
OR2X2 OR2X2_6 ( .A(datapath_1_ALU_aluInA_3_), .B(datapath_1_ALU_aluInB_3_), .Y(_203_) );
NAND2X1 NAND2X1_950 ( .A(datapath_1_ALU_aluInA_3_), .B(datapath_1_ALU_aluInB_3_), .Y(_204_) );
AOI21X1 AOI21X1_514 ( .A(_203_), .B(_204_), .C(_202_), .Y(_205_) );
XNOR2X1 XNOR2X1_3 ( .A(datapath_1_ALU_aluInA_7_), .B(datapath_1_ALU_aluInB_7_), .Y(_206_) );
NOR2X1 NOR2X1_209 ( .A(datapath_1_ALU_aluInA_6_), .B(datapath_1_ALU_aluInB_6_), .Y(_207_) );
AND2X2 AND2X2_11 ( .A(datapath_1_ALU_aluInA_6_), .B(datapath_1_ALU_aluInB_6_), .Y(_208_) );
OAI21X1 OAI21X1_1437 ( .A(_207_), .B(_208_), .C(_206_), .Y(_209_) );
OR2X2 OR2X2_7 ( .A(datapath_1_ALU_aluInA_4_), .B(datapath_1_ALU_aluInB_4_), .Y(_210_) );
NAND2X1 NAND2X1_951 ( .A(datapath_1_ALU_aluInA_4_), .B(datapath_1_ALU_aluInB_4_), .Y(_211_) );
NAND2X1 NAND2X1_952 ( .A(_211_), .B(_210_), .Y(_212_) );
NOR2X1 NOR2X1_210 ( .A(datapath_1_ALU_aluInA_5_), .B(datapath_1_ALU_aluInB_5_), .Y(_213_) );
AND2X2 AND2X2_12 ( .A(datapath_1_ALU_aluInA_5_), .B(datapath_1_ALU_aluInB_5_), .Y(_214_) );
OAI21X1 OAI21X1_1438 ( .A(_213_), .B(_214_), .C(_212_), .Y(_215_) );
NOR2X1 NOR2X1_211 ( .A(_215_), .B(_209_), .Y(_216_) );
NOR2X1 NOR2X1_212 ( .A(datapath_1_ALU_aluInA_0_), .B(datapath_1_ALU_aluInB_0_), .Y(_217_) );
NAND2X1 NAND2X1_953 ( .A(datapath_1_ALU_aluInA_0_), .B(datapath_1_ALU_aluInB_0_), .Y(_218_) );
INVX1 INVX1_276 ( .A(_218_), .Y(_219_) );
NOR2X1 NOR2X1_213 ( .A(_217_), .B(_219_), .Y(_220_) );
NOR2X1 NOR2X1_214 ( .A(datapath_1_ALU_aluInA_1_), .B(datapath_1_ALU_aluInB_1_), .Y(_221_) );
AND2X2 AND2X2_13 ( .A(datapath_1_ALU_aluInA_1_), .B(datapath_1_ALU_aluInB_1_), .Y(_222_) );
NOR2X1 NOR2X1_215 ( .A(_221_), .B(_222_), .Y(_223_) );
NOR2X1 NOR2X1_216 ( .A(_223_), .B(_220_), .Y(_224_) );
NAND3X1 NAND3X1_1365 ( .A(_205_), .B(_224_), .C(_216_), .Y(_225_) );
NOR2X1 NOR2X1_217 ( .A(_225_), .B(_201_), .Y(_226_) );
NAND3X1 NAND3X1_1366 ( .A(_127_), .B(_226_), .C(_172_), .Y(_227_) );
INVX1 INVX1_277 ( .A(aluControl_0_), .Y(_228_) );
NOR2X1 NOR2X1_218 ( .A(aluControl_1_), .B(_228_), .Y(_229_) );
INVX1 INVX1_278 ( .A(_229_), .Y(_230_) );
INVX1 INVX1_279 ( .A(aluControl_3_), .Y(_231_) );
NOR2X1 NOR2X1_219 ( .A(aluControl_2_), .B(_231_), .Y(_232_) );
NOR2X1 NOR2X1_220 ( .A(aluControl_0_), .B(aluControl_1_), .Y(_233_) );
OAI21X1 OAI21X1_1439 ( .A(_233_), .B(_227_), .C(_232_), .Y(_234_) );
AOI21X1 AOI21X1_515 ( .A(_227_), .B(_230_), .C(_234_), .Y(datapath_1_ALU_aluZero) );
NOR2X1 NOR2X1_221 ( .A(aluControl_3_), .B(aluControl_2_), .Y(_235_) );
INVX1 INVX1_280 ( .A(_235_), .Y(_236_) );
NOR2X1 NOR2X1_222 ( .A(_236_), .B(_230_), .Y(_237_) );
INVX1 INVX1_281 ( .A(_237__bF_buf3), .Y(_238_) );
AND2X2 AND2X2_14 ( .A(aluControl_3_), .B(aluControl_2_), .Y(_239_) );
NAND2X1 NAND2X1_954 ( .A(_239_), .B(_229_), .Y(_240_) );
INVX1 INVX1_282 ( .A(_240__bF_buf4), .Y(_241_) );
NAND2X1 NAND2X1_955 ( .A(aluControl_1_), .B(_228_), .Y(_242_) );
NOR2X1 NOR2X1_223 ( .A(aluControl_3_), .B(_242_), .Y(_243_) );
OAI21X1 OAI21X1_1440 ( .A(_243_), .B(_241_), .C(_220_), .Y(_244_) );
NAND2X1 NAND2X1_956 ( .A(_233_), .B(_235_), .Y(_245_) );
INVX1 INVX1_283 ( .A(_245__bF_buf0), .Y(_246_) );
NAND2X1 NAND2X1_957 ( .A(_233_), .B(_239_), .Y(_247_) );
INVX1 INVX1_284 ( .A(_247_), .Y(_248_) );
AOI22X1 AOI22X1_120 ( .A(_246_), .B(_219_), .C(_217_), .D(_248__bF_buf2), .Y(_249_) );
AND2X2 AND2X2_15 ( .A(_244_), .B(_249_), .Y(_250_) );
OAI21X1 OAI21X1_1441 ( .A(_217_), .B(_238_), .C(_250_), .Y(datapath_1_ALU_aluResult_0_) );
INVX1 INVX1_285 ( .A(datapath_1_ALU_aluInA_0_), .Y(_251_) );
NAND2X1 NAND2X1_958 ( .A(datapath_1_ALU_aluInB_0_), .B(_251_), .Y(_252_) );
OAI21X1 OAI21X1_1442 ( .A(_221_), .B(_222_), .C(_252_), .Y(_253_) );
INVX1 INVX1_286 ( .A(_253_), .Y(_254_) );
INVX1 INVX1_287 ( .A(_223_), .Y(_255_) );
NAND2X1 NAND2X1_959 ( .A(aluControl_2_), .B(_243_), .Y(_256_) );
INVX1 INVX1_288 ( .A(_256__bF_buf2), .Y(_257_) );
OAI21X1 OAI21X1_1443 ( .A(_255_), .B(_252_), .C(_257_), .Y(_258_) );
NOR2X1 NOR2X1_224 ( .A(_218_), .B(_255_), .Y(_259_) );
NOR2X1 NOR2X1_225 ( .A(_242_), .B(_236_), .Y(_260_) );
OAI21X1 OAI21X1_1444 ( .A(_219_), .B(_223_), .C(_260_), .Y(_261_) );
NAND2X1 NAND2X1_960 ( .A(datapath_1_ALU_aluInA_1_), .B(datapath_1_ALU_aluInB_1_), .Y(_262_) );
OAI22X1 OAI22X1_112 ( .A(_262_), .B(_245__bF_buf1), .C(_240__bF_buf0), .D(_255_), .Y(_263_) );
NAND2X1 NAND2X1_961 ( .A(_221_), .B(_248__bF_buf2), .Y(_264_) );
OAI21X1 OAI21X1_1445 ( .A(_221_), .B(_238_), .C(_264_), .Y(_265_) );
NOR2X1 NOR2X1_226 ( .A(_263_), .B(_265_), .Y(_266_) );
OAI21X1 OAI21X1_1446 ( .A(_259_), .B(_261_), .C(_266_), .Y(_267_) );
INVX1 INVX1_289 ( .A(_267_), .Y(_268_) );
OAI21X1 OAI21X1_1447 ( .A(_254_), .B(_258_), .C(_268_), .Y(datapath_1_ALU_aluResult_1_) );
XNOR2X1 XNOR2X1_4 ( .A(datapath_1_ALU_aluInA_2_), .B(datapath_1_ALU_aluInB_2_), .Y(_269_) );
INVX1 INVX1_290 ( .A(datapath_1_ALU_aluInB_1_), .Y(_270_) );
NAND2X1 NAND2X1_962 ( .A(datapath_1_ALU_aluInA_1_), .B(_270_), .Y(_271_) );
NAND2X1 NAND2X1_963 ( .A(_271_), .B(_253_), .Y(_272_) );
NAND2X1 NAND2X1_964 ( .A(_269_), .B(_272_), .Y(_273_) );
INVX1 INVX1_291 ( .A(_273_), .Y(_274_) );
OAI21X1 OAI21X1_1448 ( .A(_269_), .B(_272_), .C(_257_), .Y(_275_) );
OAI21X1 OAI21X1_1449 ( .A(_218_), .B(_221_), .C(_262_), .Y(_276_) );
INVX1 INVX1_292 ( .A(_260_), .Y(_277_) );
OAI21X1 OAI21X1_1450 ( .A(_222_), .B(_259_), .C(_202_), .Y(_278_) );
INVX1 INVX1_293 ( .A(_278_), .Y(_279_) );
NOR2X1 NOR2X1_227 ( .A(_277__bF_buf0), .B(_279_), .Y(_280_) );
OAI21X1 OAI21X1_1451 ( .A(_202_), .B(_276_), .C(_280_), .Y(_281_) );
INVX1 INVX1_294 ( .A(datapath_1_ALU_aluInA_2_), .Y(_282_) );
INVX1 INVX1_295 ( .A(datapath_1_ALU_aluInB_2_), .Y(_283_) );
NOR2X1 NOR2X1_228 ( .A(_282_), .B(_283_), .Y(_284_) );
INVX1 INVX1_296 ( .A(_284_), .Y(_285_) );
OAI22X1 OAI22X1_113 ( .A(_245__bF_buf1), .B(_285_), .C(_269_), .D(_240__bF_buf0), .Y(_286_) );
NAND2X1 NAND2X1_965 ( .A(_282_), .B(_283_), .Y(_287_) );
OAI21X1 OAI21X1_1452 ( .A(datapath_1_ALU_aluInA_2_), .B(datapath_1_ALU_aluInB_2_), .C(_237__bF_buf2), .Y(_288_) );
OAI21X1 OAI21X1_1453 ( .A(_247_), .B(_287_), .C(_288_), .Y(_289_) );
NOR2X1 NOR2X1_229 ( .A(_286_), .B(_289_), .Y(_290_) );
AND2X2 AND2X2_16 ( .A(_281_), .B(_290_), .Y(_291_) );
OAI21X1 OAI21X1_1454 ( .A(_274_), .B(_275_), .C(_291_), .Y(datapath_1_ALU_aluResult_2_) );
NAND2X1 NAND2X1_966 ( .A(_204_), .B(_203_), .Y(_292_) );
OAI21X1 OAI21X1_1455 ( .A(_282_), .B(datapath_1_ALU_aluInB_2_), .C(_273_), .Y(_293_) );
NAND2X1 NAND2X1_967 ( .A(_292_), .B(_269_), .Y(_294_) );
AOI21X1 AOI21X1_516 ( .A(_253_), .B(_271_), .C(_294_), .Y(_295_) );
NAND2X1 NAND2X1_968 ( .A(datapath_1_ALU_aluInA_2_), .B(_283_), .Y(_296_) );
NOR2X1 NOR2X1_230 ( .A(datapath_1_ALU_aluInA_3_), .B(datapath_1_ALU_aluInB_3_), .Y(_297_) );
AND2X2 AND2X2_17 ( .A(datapath_1_ALU_aluInA_3_), .B(datapath_1_ALU_aluInB_3_), .Y(_298_) );
NOR2X1 NOR2X1_231 ( .A(_297_), .B(_298_), .Y(_299_) );
OAI21X1 OAI21X1_1456 ( .A(_296_), .B(_299_), .C(_257_), .Y(_300_) );
NOR2X1 NOR2X1_232 ( .A(_295_), .B(_300_), .Y(_301_) );
OAI21X1 OAI21X1_1457 ( .A(_292_), .B(_293_), .C(_301_), .Y(_302_) );
NAND3X1 NAND3X1_1367 ( .A(_292_), .B(_285_), .C(_278_), .Y(_303_) );
OAI21X1 OAI21X1_1458 ( .A(_284_), .B(_279_), .C(_299_), .Y(_304_) );
NAND3X1 NAND3X1_1368 ( .A(_260_), .B(_303_), .C(_304_), .Y(_305_) );
OAI22X1 OAI22X1_114 ( .A(_204_), .B(_245__bF_buf1), .C(_297_), .D(_238_), .Y(_306_) );
OAI22X1 OAI22X1_115 ( .A(_203_), .B(_247_), .C(_292_), .D(_240__bF_buf0), .Y(_307_) );
NOR2X1 NOR2X1_233 ( .A(_307_), .B(_306_), .Y(_308_) );
NAND3X1 NAND3X1_1369 ( .A(_302_), .B(_308_), .C(_305_), .Y(datapath_1_ALU_aluResult_3_) );
NOR2X1 NOR2X1_234 ( .A(datapath_1_ALU_aluInA_4_), .B(datapath_1_ALU_aluInB_4_), .Y(_309_) );
AND2X2 AND2X2_18 ( .A(datapath_1_ALU_aluInA_4_), .B(datapath_1_ALU_aluInB_4_), .Y(_310_) );
NOR2X1 NOR2X1_235 ( .A(_309_), .B(_310_), .Y(_311_) );
NAND3X1 NAND3X1_1370 ( .A(_299_), .B(_202_), .C(_276_), .Y(_312_) );
AOI21X1 AOI21X1_517 ( .A(_284_), .B(_203_), .C(_298_), .Y(_313_) );
NAND2X1 NAND2X1_969 ( .A(_313_), .B(_312_), .Y(_314_) );
NAND2X1 NAND2X1_970 ( .A(_311_), .B(_314_), .Y(_315_) );
NAND2X1 NAND2X1_971 ( .A(_260_), .B(_315_), .Y(_316_) );
OAI21X1 OAI21X1_1459 ( .A(_212_), .B(_240__bF_buf1), .C(_316_), .Y(_317_) );
OAI21X1 OAI21X1_1460 ( .A(_311_), .B(_314_), .C(_317_), .Y(_318_) );
INVX1 INVX1_297 ( .A(datapath_1_ALU_aluInB_3_), .Y(_319_) );
NAND2X1 NAND2X1_972 ( .A(datapath_1_ALU_aluInA_3_), .B(_319_), .Y(_320_) );
OAI21X1 OAI21X1_1461 ( .A(_296_), .B(_299_), .C(_320_), .Y(_321_) );
AOI21X1 AOI21X1_518 ( .A(_205_), .B(_272_), .C(_321_), .Y(_322_) );
NAND2X1 NAND2X1_973 ( .A(_311_), .B(_322_), .Y(_323_) );
OAI21X1 OAI21X1_1462 ( .A(_321_), .B(_295_), .C(_212_), .Y(_324_) );
NAND3X1 NAND3X1_1371 ( .A(_257_), .B(_324_), .C(_323_), .Y(_325_) );
OAI21X1 OAI21X1_1463 ( .A(datapath_1_ALU_aluInA_4_), .B(datapath_1_ALU_aluInB_4_), .C(_237__bF_buf2), .Y(_326_) );
OAI21X1 OAI21X1_1464 ( .A(_210_), .B(_247_), .C(_326_), .Y(_327_) );
AOI21X1 AOI21X1_519 ( .A(_310_), .B(_246_), .C(_327_), .Y(_328_) );
NAND3X1 NAND3X1_1372 ( .A(_325_), .B(_328_), .C(_318_), .Y(datapath_1_ALU_aluResult_4_) );
OR2X2 OR2X2_8 ( .A(datapath_1_ALU_aluInA_5_), .B(datapath_1_ALU_aluInB_5_), .Y(_329_) );
NAND2X1 NAND2X1_974 ( .A(datapath_1_ALU_aluInA_5_), .B(datapath_1_ALU_aluInB_5_), .Y(_330_) );
NAND2X1 NAND2X1_975 ( .A(_330_), .B(_329_), .Y(_331_) );
INVX1 INVX1_298 ( .A(datapath_1_ALU_aluInB_4_), .Y(_332_) );
NAND2X1 NAND2X1_976 ( .A(datapath_1_ALU_aluInA_4_), .B(_332_), .Y(_333_) );
OAI21X1 OAI21X1_1465 ( .A(_311_), .B(_322_), .C(_333_), .Y(_334_) );
XNOR2X1 XNOR2X1_5 ( .A(_334_), .B(_331_), .Y(_335_) );
NOR2X1 NOR2X1_236 ( .A(_213_), .B(_214_), .Y(_336_) );
NAND2X1 NAND2X1_977 ( .A(_211_), .B(_315_), .Y(_337_) );
NOR2X1 NOR2X1_237 ( .A(_331_), .B(_315_), .Y(_338_) );
OAI21X1 OAI21X1_1466 ( .A(_211_), .B(_331_), .C(_260_), .Y(_339_) );
NOR2X1 NOR2X1_238 ( .A(_339_), .B(_338_), .Y(_340_) );
OAI21X1 OAI21X1_1467 ( .A(_336_), .B(_337_), .C(_340_), .Y(_341_) );
MUX2X1 MUX2X1_126 ( .A(_237__bF_buf2), .B(_248__bF_buf2), .S(_329_), .Y(_342_) );
OAI21X1 OAI21X1_1468 ( .A(_330_), .B(_245__bF_buf2), .C(_342_), .Y(_343_) );
AOI21X1 AOI21X1_520 ( .A(_336_), .B(_241_), .C(_343_), .Y(_344_) );
AND2X2 AND2X2_19 ( .A(_341_), .B(_344_), .Y(_345_) );
OAI21X1 OAI21X1_1469 ( .A(_256__bF_buf3), .B(_335_), .C(_345_), .Y(datapath_1_ALU_aluResult_5_) );
INVX1 INVX1_299 ( .A(datapath_1_ALU_aluInA_6_), .Y(_346_) );
INVX1 INVX1_300 ( .A(datapath_1_ALU_aluInB_6_), .Y(_347_) );
NAND2X1 NAND2X1_978 ( .A(_346_), .B(_347_), .Y(_348_) );
NAND2X1 NAND2X1_979 ( .A(datapath_1_ALU_aluInA_6_), .B(datapath_1_ALU_aluInB_6_), .Y(_349_) );
NAND2X1 NAND2X1_980 ( .A(_349_), .B(_348_), .Y(_350_) );
INVX1 INVX1_301 ( .A(datapath_1_ALU_aluInB_5_), .Y(_351_) );
NAND2X1 NAND2X1_981 ( .A(datapath_1_ALU_aluInA_5_), .B(_351_), .Y(_352_) );
OAI21X1 OAI21X1_1470 ( .A(_333_), .B(_336_), .C(_352_), .Y(_353_) );
INVX1 INVX1_302 ( .A(_353_), .Y(_354_) );
OAI21X1 OAI21X1_1471 ( .A(_215_), .B(_322_), .C(_354_), .Y(_355_) );
AOI21X1 AOI21X1_521 ( .A(_355_), .B(_350_), .C(_256__bF_buf0), .Y(_356_) );
OAI21X1 OAI21X1_1472 ( .A(_350_), .B(_355_), .C(_356_), .Y(_357_) );
OAI21X1 OAI21X1_1473 ( .A(_211_), .B(_213_), .C(_330_), .Y(_358_) );
NOR2X1 NOR2X1_239 ( .A(_358_), .B(_338_), .Y(_359_) );
OAI21X1 OAI21X1_1474 ( .A(_207_), .B(_208_), .C(_359_), .Y(_360_) );
NOR2X1 NOR2X1_240 ( .A(_207_), .B(_208_), .Y(_361_) );
OAI21X1 OAI21X1_1475 ( .A(_358_), .B(_338_), .C(_361_), .Y(_362_) );
NAND3X1 NAND3X1_1373 ( .A(_260_), .B(_362_), .C(_360_), .Y(_363_) );
OAI21X1 OAI21X1_1476 ( .A(datapath_1_ALU_aluInA_6_), .B(datapath_1_ALU_aluInB_6_), .C(_237__bF_buf1), .Y(_364_) );
OAI21X1 OAI21X1_1477 ( .A(_348_), .B(_247_), .C(_364_), .Y(_365_) );
OAI22X1 OAI22X1_116 ( .A(_349_), .B(_245__bF_buf2), .C(_350_), .D(_240__bF_buf1), .Y(_366_) );
NOR2X1 NOR2X1_241 ( .A(_366_), .B(_365_), .Y(_367_) );
NAND3X1 NAND3X1_1374 ( .A(_357_), .B(_367_), .C(_363_), .Y(datapath_1_ALU_aluResult_6_) );
OAI21X1 OAI21X1_1478 ( .A(_207_), .B(_208_), .C(_355_), .Y(_368_) );
OAI21X1 OAI21X1_1479 ( .A(_346_), .B(datapath_1_ALU_aluInB_6_), .C(_368_), .Y(_369_) );
AOI21X1 AOI21X1_522 ( .A(_369_), .B(_206_), .C(_256__bF_buf0), .Y(_370_) );
OAI21X1 OAI21X1_1480 ( .A(_206_), .B(_369_), .C(_370_), .Y(_371_) );
NOR2X1 NOR2X1_242 ( .A(datapath_1_ALU_aluInA_7_), .B(datapath_1_ALU_aluInB_7_), .Y(_372_) );
AND2X2 AND2X2_20 ( .A(datapath_1_ALU_aluInA_7_), .B(datapath_1_ALU_aluInB_7_), .Y(_373_) );
NOR2X1 NOR2X1_243 ( .A(_372_), .B(_373_), .Y(_374_) );
OAI21X1 OAI21X1_1481 ( .A(_346_), .B(_347_), .C(_362_), .Y(_375_) );
AOI21X1 AOI21X1_523 ( .A(_375_), .B(_374_), .C(_277__bF_buf0), .Y(_376_) );
OAI21X1 OAI21X1_1482 ( .A(_374_), .B(_375_), .C(_376_), .Y(_377_) );
NAND2X1 NAND2X1_982 ( .A(_373_), .B(_246_), .Y(_378_) );
OAI21X1 OAI21X1_1483 ( .A(_206_), .B(_240__bF_buf1), .C(_378_), .Y(_379_) );
NAND2X1 NAND2X1_983 ( .A(_372_), .B(_248__bF_buf2), .Y(_380_) );
OAI21X1 OAI21X1_1484 ( .A(_372_), .B(_238_), .C(_380_), .Y(_381_) );
NOR2X1 NOR2X1_244 ( .A(_379_), .B(_381_), .Y(_382_) );
NAND3X1 NAND3X1_1375 ( .A(_371_), .B(_382_), .C(_377_), .Y(datapath_1_ALU_aluResult_7_) );
NAND2X1 NAND2X1_984 ( .A(_311_), .B(_336_), .Y(_383_) );
NAND2X1 NAND2X1_985 ( .A(_374_), .B(_361_), .Y(_384_) );
NOR2X1 NOR2X1_245 ( .A(_383_), .B(_384_), .Y(_385_) );
INVX1 INVX1_303 ( .A(_358_), .Y(_386_) );
AOI21X1 AOI21X1_524 ( .A(_374_), .B(_208_), .C(_373_), .Y(_387_) );
OAI21X1 OAI21X1_1485 ( .A(_386_), .B(_384_), .C(_387_), .Y(_388_) );
AOI21X1 AOI21X1_525 ( .A(_385_), .B(_314_), .C(_388_), .Y(_389_) );
OAI21X1 OAI21X1_1486 ( .A(_192_), .B(_194_), .C(_389_), .Y(_390_) );
INVX1 INVX1_304 ( .A(_192_), .Y(_391_) );
NAND2X1 NAND2X1_986 ( .A(_193_), .B(_391_), .Y(_392_) );
NOR2X1 NOR2X1_246 ( .A(_392_), .B(_389_), .Y(_393_) );
OAI22X1 OAI22X1_117 ( .A(_392_), .B(_240__bF_buf2), .C(_277__bF_buf2), .D(_393_), .Y(_394_) );
NAND2X1 NAND2X1_987 ( .A(_390_), .B(_394_), .Y(_395_) );
NOR2X1 NOR2X1_247 ( .A(_374_), .B(_361_), .Y(_396_) );
NAND3X1 NAND3X1_1376 ( .A(_212_), .B(_331_), .C(_396_), .Y(_397_) );
NAND2X1 NAND2X1_988 ( .A(datapath_1_ALU_aluInA_6_), .B(_347_), .Y(_398_) );
INVX1 INVX1_305 ( .A(datapath_1_ALU_aluInB_7_), .Y(_399_) );
NAND2X1 NAND2X1_989 ( .A(datapath_1_ALU_aluInA_7_), .B(_399_), .Y(_400_) );
OAI21X1 OAI21X1_1487 ( .A(_398_), .B(_374_), .C(_400_), .Y(_401_) );
AOI21X1 AOI21X1_526 ( .A(_353_), .B(_396_), .C(_401_), .Y(_402_) );
OAI21X1 OAI21X1_1488 ( .A(_397_), .B(_322_), .C(_402_), .Y(_403_) );
OAI21X1 OAI21X1_1489 ( .A(_192_), .B(_194_), .C(_403_), .Y(_404_) );
INVX1 INVX1_306 ( .A(_404_), .Y(_405_) );
NOR2X1 NOR2X1_248 ( .A(_256__bF_buf1), .B(_405_), .Y(_406_) );
OAI21X1 OAI21X1_1490 ( .A(_392_), .B(_403_), .C(_406_), .Y(_407_) );
OAI21X1 OAI21X1_1491 ( .A(datapath_1_ALU_aluInA_8_), .B(datapath_1_ALU_aluInB_8_), .C(_237__bF_buf3), .Y(_408_) );
OAI21X1 OAI21X1_1492 ( .A(_391_), .B(_247_), .C(_408_), .Y(_409_) );
AOI21X1 AOI21X1_527 ( .A(_194_), .B(_246_), .C(_409_), .Y(_410_) );
NAND3X1 NAND3X1_1377 ( .A(_395_), .B(_410_), .C(_407_), .Y(datapath_1_ALU_aluResult_8_) );
NOR2X1 NOR2X1_249 ( .A(datapath_1_ALU_aluInA_9_), .B(datapath_1_ALU_aluInB_9_), .Y(_411_) );
AND2X2 AND2X2_21 ( .A(datapath_1_ALU_aluInA_9_), .B(datapath_1_ALU_aluInB_9_), .Y(_412_) );
OAI21X1 OAI21X1_1493 ( .A(_411_), .B(_412_), .C(_193_), .Y(_413_) );
NOR2X1 NOR2X1_250 ( .A(_411_), .B(_412_), .Y(_414_) );
OAI21X1 OAI21X1_1494 ( .A(_194_), .B(_393_), .C(_414_), .Y(_415_) );
OAI21X1 OAI21X1_1495 ( .A(_393_), .B(_413_), .C(_415_), .Y(_416_) );
INVX1 INVX1_307 ( .A(datapath_1_ALU_aluInB_8_), .Y(_417_) );
NAND2X1 NAND2X1_990 ( .A(datapath_1_ALU_aluInA_8_), .B(_417_), .Y(_418_) );
NAND2X1 NAND2X1_991 ( .A(_418_), .B(_404_), .Y(_419_) );
NOR2X1 NOR2X1_251 ( .A(_414_), .B(_404_), .Y(_420_) );
OAI21X1 OAI21X1_1496 ( .A(_414_), .B(_418_), .C(_257_), .Y(_421_) );
NOR2X1 NOR2X1_252 ( .A(_421_), .B(_420_), .Y(_422_) );
OAI21X1 OAI21X1_1497 ( .A(_191_), .B(_419_), .C(_422_), .Y(_423_) );
OAI22X1 OAI22X1_118 ( .A(_190_), .B(_245__bF_buf3), .C(_191_), .D(_240__bF_buf4), .Y(_424_) );
OAI21X1 OAI21X1_1498 ( .A(datapath_1_ALU_aluInA_9_), .B(datapath_1_ALU_aluInB_9_), .C(_237__bF_buf3), .Y(_425_) );
OAI21X1 OAI21X1_1499 ( .A(_189_), .B(_247_), .C(_425_), .Y(_426_) );
NOR2X1 NOR2X1_253 ( .A(_424_), .B(_426_), .Y(_427_) );
AND2X2 AND2X2_22 ( .A(_423_), .B(_427_), .Y(_428_) );
OAI21X1 OAI21X1_1500 ( .A(_277__bF_buf3), .B(_416_), .C(_428_), .Y(datapath_1_ALU_aluResult_9_) );
INVX1 INVX1_308 ( .A(datapath_1_ALU_aluInA_10_), .Y(_429_) );
NAND2X1 NAND2X1_992 ( .A(datapath_1_ALU_aluInB_10_), .B(_429_), .Y(_430_) );
INVX1 INVX1_309 ( .A(datapath_1_ALU_aluInB_10_), .Y(_431_) );
NAND2X1 NAND2X1_993 ( .A(datapath_1_ALU_aluInA_10_), .B(_431_), .Y(_432_) );
NAND2X1 NAND2X1_994 ( .A(_430_), .B(_432_), .Y(_433_) );
NAND3X1 NAND3X1_1378 ( .A(_391_), .B(_193_), .C(_414_), .Y(_434_) );
OAI21X1 OAI21X1_1501 ( .A(_193_), .B(_411_), .C(_190_), .Y(_435_) );
INVX1 INVX1_310 ( .A(_435_), .Y(_436_) );
OAI21X1 OAI21X1_1502 ( .A(_434_), .B(_389_), .C(_436_), .Y(_437_) );
AOI21X1 AOI21X1_528 ( .A(_437_), .B(_433_), .C(_277__bF_buf3), .Y(_438_) );
OAI21X1 OAI21X1_1503 ( .A(_433_), .B(_437_), .C(_438_), .Y(_439_) );
NAND2X1 NAND2X1_995 ( .A(datapath_1_ALU_aluInA_9_), .B(_188_), .Y(_440_) );
OAI21X1 OAI21X1_1504 ( .A(_418_), .B(_414_), .C(_440_), .Y(_441_) );
NOR2X1 NOR2X1_254 ( .A(_441_), .B(_420_), .Y(_442_) );
NAND2X1 NAND2X1_996 ( .A(_433_), .B(_442_), .Y(_443_) );
OAI21X1 OAI21X1_1505 ( .A(_441_), .B(_420_), .C(_196_), .Y(_444_) );
NAND3X1 NAND3X1_1379 ( .A(_257_), .B(_444_), .C(_443_), .Y(_445_) );
NAND2X1 NAND2X1_997 ( .A(datapath_1_ALU_aluInA_10_), .B(datapath_1_ALU_aluInB_10_), .Y(_446_) );
OAI22X1 OAI22X1_119 ( .A(_245__bF_buf3), .B(_446_), .C(_196_), .D(_240__bF_buf2), .Y(_447_) );
NAND2X1 NAND2X1_998 ( .A(_429_), .B(_431_), .Y(_448_) );
OAI21X1 OAI21X1_1506 ( .A(datapath_1_ALU_aluInA_10_), .B(datapath_1_ALU_aluInB_10_), .C(_237__bF_buf3), .Y(_449_) );
OAI21X1 OAI21X1_1507 ( .A(_247_), .B(_448_), .C(_449_), .Y(_450_) );
NOR2X1 NOR2X1_255 ( .A(_447_), .B(_450_), .Y(_451_) );
NAND3X1 NAND3X1_1380 ( .A(_439_), .B(_451_), .C(_445_), .Y(datapath_1_ALU_aluResult_10_) );
NOR2X1 NOR2X1_256 ( .A(_197_), .B(_198_), .Y(_452_) );
NAND2X1 NAND2X1_999 ( .A(_433_), .B(_437_), .Y(_453_) );
OAI21X1 OAI21X1_1508 ( .A(_429_), .B(_431_), .C(_453_), .Y(_454_) );
AOI21X1 AOI21X1_529 ( .A(_454_), .B(_452_), .C(_277__bF_buf2), .Y(_455_) );
OAI21X1 OAI21X1_1509 ( .A(_452_), .B(_454_), .C(_455_), .Y(_456_) );
INVX1 INVX1_311 ( .A(_452_), .Y(_457_) );
OAI21X1 OAI21X1_1510 ( .A(_429_), .B(datapath_1_ALU_aluInB_10_), .C(_444_), .Y(_458_) );
AOI21X1 AOI21X1_530 ( .A(_458_), .B(_457_), .C(_256__bF_buf1), .Y(_459_) );
OAI21X1 OAI21X1_1511 ( .A(_457_), .B(_458_), .C(_459_), .Y(_460_) );
INVX1 INVX1_312 ( .A(_198_), .Y(_461_) );
OAI22X1 OAI22X1_120 ( .A(_461_), .B(_245__bF_buf3), .C(_240__bF_buf2), .D(_457_), .Y(_462_) );
NAND2X1 NAND2X1_1000 ( .A(_197_), .B(_248__bF_buf1), .Y(_463_) );
OAI21X1 OAI21X1_1512 ( .A(_197_), .B(_238_), .C(_463_), .Y(_464_) );
NOR2X1 NOR2X1_257 ( .A(_462_), .B(_464_), .Y(_465_) );
NAND3X1 NAND3X1_1381 ( .A(_456_), .B(_465_), .C(_460_), .Y(datapath_1_ALU_aluResult_11_) );
INVX1 INVX1_313 ( .A(_181_), .Y(_466_) );
OAI22X1 OAI22X1_121 ( .A(_466_), .B(_245__bF_buf3), .C(_180_), .D(_238_), .Y(_467_) );
NOR2X1 NOR2X1_258 ( .A(_452_), .B(_433_), .Y(_468_) );
INVX1 INVX1_314 ( .A(datapath_1_ALU_aluInB_11_), .Y(_469_) );
NAND2X1 NAND2X1_1001 ( .A(datapath_1_ALU_aluInA_11_), .B(_469_), .Y(_470_) );
OAI21X1 OAI21X1_1513 ( .A(_432_), .B(_452_), .C(_470_), .Y(_471_) );
AOI21X1 AOI21X1_531 ( .A(_468_), .B(_441_), .C(_471_), .Y(_472_) );
INVX1 INVX1_315 ( .A(_472_), .Y(_473_) );
AOI21X1 AOI21X1_532 ( .A(_403_), .B(_200_), .C(_473_), .Y(_474_) );
NAND2X1 NAND2X1_1002 ( .A(_182_), .B(_474_), .Y(_475_) );
NOR2X1 NOR2X1_259 ( .A(_182_), .B(_474_), .Y(_476_) );
INVX1 INVX1_316 ( .A(_476_), .Y(_477_) );
NAND3X1 NAND3X1_1382 ( .A(_257_), .B(_475_), .C(_477_), .Y(_478_) );
NAND2X1 NAND2X1_1003 ( .A(_452_), .B(_433_), .Y(_479_) );
OAI21X1 OAI21X1_1514 ( .A(_446_), .B(_197_), .C(_461_), .Y(_480_) );
INVX1 INVX1_317 ( .A(_480_), .Y(_481_) );
OAI21X1 OAI21X1_1515 ( .A(_436_), .B(_479_), .C(_481_), .Y(_482_) );
INVX1 INVX1_318 ( .A(_482_), .Y(_483_) );
NOR2X1 NOR2X1_260 ( .A(_479_), .B(_434_), .Y(_484_) );
INVX1 INVX1_319 ( .A(_484_), .Y(_485_) );
OAI21X1 OAI21X1_1516 ( .A(_485_), .B(_389_), .C(_483_), .Y(_486_) );
AOI21X1 AOI21X1_533 ( .A(_486_), .B(_182_), .C(_277__bF_buf2), .Y(_487_) );
OAI21X1 OAI21X1_1517 ( .A(_182_), .B(_486_), .C(_487_), .Y(_488_) );
AOI22X1 AOI22X1_121 ( .A(_180_), .B(_248__bF_buf0), .C(_182_), .D(_241_), .Y(_489_) );
NAND3X1 NAND3X1_1383 ( .A(_488_), .B(_489_), .C(_478_), .Y(_490_) );
OR2X2 OR2X2_9 ( .A(_490_), .B(_467_), .Y(datapath_1_ALU_aluResult_12_) );
INVX1 INVX1_320 ( .A(_185_), .Y(_491_) );
INVX1 INVX1_321 ( .A(datapath_1_ALU_aluInB_12_), .Y(_492_) );
NAND2X1 NAND2X1_1004 ( .A(datapath_1_ALU_aluInA_12_), .B(_492_), .Y(_493_) );
OAI21X1 OAI21X1_1518 ( .A(_182_), .B(_474_), .C(_493_), .Y(_494_) );
XNOR2X1 XNOR2X1_6 ( .A(_494_), .B(_491_), .Y(_495_) );
AOI22X1 AOI22X1_122 ( .A(_184_), .B(_246_), .C(_185_), .D(_241_), .Y(_496_) );
OAI21X1 OAI21X1_1519 ( .A(_183_), .B(_238_), .C(_496_), .Y(_497_) );
NAND2X1 NAND2X1_1005 ( .A(_182_), .B(_486_), .Y(_498_) );
NAND2X1 NAND2X1_1006 ( .A(_466_), .B(_498_), .Y(_499_) );
NOR2X1 NOR2X1_261 ( .A(_491_), .B(_498_), .Y(_500_) );
OAI21X1 OAI21X1_1520 ( .A(_466_), .B(_491_), .C(_260_), .Y(_501_) );
NOR2X1 NOR2X1_262 ( .A(_501_), .B(_500_), .Y(_502_) );
OAI21X1 OAI21X1_1521 ( .A(_185_), .B(_499_), .C(_502_), .Y(_503_) );
NAND2X1 NAND2X1_1007 ( .A(_183_), .B(_248__bF_buf0), .Y(_504_) );
NAND2X1 NAND2X1_1008 ( .A(_504_), .B(_503_), .Y(_505_) );
NOR2X1 NOR2X1_263 ( .A(_497_), .B(_505_), .Y(_506_) );
OAI21X1 OAI21X1_1522 ( .A(_256__bF_buf1), .B(_495_), .C(_506_), .Y(datapath_1_ALU_aluResult_13_) );
INVX1 INVX1_322 ( .A(_178_), .Y(_507_) );
INVX1 INVX1_323 ( .A(datapath_1_ALU_aluInB_13_), .Y(_508_) );
NAND2X1 NAND2X1_1009 ( .A(datapath_1_ALU_aluInA_13_), .B(_508_), .Y(_509_) );
OAI21X1 OAI21X1_1523 ( .A(_493_), .B(_185_), .C(_509_), .Y(_510_) );
INVX1 INVX1_324 ( .A(_510_), .Y(_511_) );
OAI21X1 OAI21X1_1524 ( .A(_185_), .B(_477_), .C(_511_), .Y(_512_) );
AND2X2 AND2X2_23 ( .A(_512_), .B(_507_), .Y(_513_) );
NOR2X1 NOR2X1_264 ( .A(_256__bF_buf1), .B(_513_), .Y(_514_) );
OAI21X1 OAI21X1_1525 ( .A(_507_), .B(_512_), .C(_514_), .Y(_515_) );
AOI21X1 AOI21X1_534 ( .A(_185_), .B(_181_), .C(_184_), .Y(_516_) );
INVX1 INVX1_325 ( .A(_516_), .Y(_517_) );
NOR2X1 NOR2X1_265 ( .A(_517_), .B(_500_), .Y(_518_) );
AOI21X1 AOI21X1_535 ( .A(_518_), .B(_507_), .C(_277__bF_buf2), .Y(_519_) );
OAI21X1 OAI21X1_1526 ( .A(_507_), .B(_518_), .C(_519_), .Y(_520_) );
INVX1 INVX1_326 ( .A(_177_), .Y(_521_) );
OAI22X1 OAI22X1_122 ( .A(_521_), .B(_245__bF_buf3), .C(_240__bF_buf2), .D(_507_), .Y(_522_) );
NAND2X1 NAND2X1_1010 ( .A(_176_), .B(_248__bF_buf0), .Y(_523_) );
OAI21X1 OAI21X1_1527 ( .A(_176_), .B(_238_), .C(_523_), .Y(_524_) );
NOR2X1 NOR2X1_266 ( .A(_522_), .B(_524_), .Y(_525_) );
NAND3X1 NAND3X1_1384 ( .A(_520_), .B(_525_), .C(_515_), .Y(datapath_1_ALU_aluResult_14_) );
OAI21X1 OAI21X1_1528 ( .A(_176_), .B(_177_), .C(_512_), .Y(_526_) );
INVX1 INVX1_327 ( .A(datapath_1_ALU_aluInB_14_), .Y(_527_) );
NAND2X1 NAND2X1_1011 ( .A(datapath_1_ALU_aluInA_14_), .B(_527_), .Y(_528_) );
NAND3X1 NAND3X1_1385 ( .A(_175_), .B(_528_), .C(_526_), .Y(_529_) );
INVX1 INVX1_328 ( .A(_175_), .Y(_530_) );
INVX1 INVX1_329 ( .A(_528_), .Y(_531_) );
OAI21X1 OAI21X1_1529 ( .A(_531_), .B(_513_), .C(_530_), .Y(_532_) );
NAND3X1 NAND3X1_1386 ( .A(_257_), .B(_529_), .C(_532_), .Y(_533_) );
OAI21X1 OAI21X1_1530 ( .A(_176_), .B(_518_), .C(_521_), .Y(_534_) );
AOI21X1 AOI21X1_536 ( .A(_534_), .B(_175_), .C(_277__bF_buf2), .Y(_535_) );
OAI21X1 OAI21X1_1531 ( .A(_175_), .B(_534_), .C(_535_), .Y(_536_) );
NAND2X1 NAND2X1_1012 ( .A(_174_), .B(_246_), .Y(_537_) );
OAI21X1 OAI21X1_1532 ( .A(_530_), .B(_240__bF_buf2), .C(_537_), .Y(_538_) );
NAND2X1 NAND2X1_1013 ( .A(_173_), .B(_248__bF_buf0), .Y(_539_) );
OAI21X1 OAI21X1_1533 ( .A(_173_), .B(_238_), .C(_539_), .Y(_540_) );
NOR2X1 NOR2X1_267 ( .A(_538_), .B(_540_), .Y(_541_) );
NAND3X1 NAND3X1_1387 ( .A(_536_), .B(_541_), .C(_533_), .Y(datapath_1_ALU_aluResult_15_) );
INVX1 INVX1_330 ( .A(_115_), .Y(_542_) );
NAND2X1 NAND2X1_1014 ( .A(_179_), .B(_186_), .Y(_543_) );
OR2X2 OR2X2_10 ( .A(_195_), .B(_199_), .Y(_544_) );
NOR2X1 NOR2X1_268 ( .A(_543_), .B(_544_), .Y(_545_) );
INVX1 INVX1_331 ( .A(datapath_1_ALU_aluInB_15_), .Y(_546_) );
NAND2X1 NAND2X1_1015 ( .A(datapath_1_ALU_aluInA_15_), .B(_546_), .Y(_547_) );
OAI21X1 OAI21X1_1534 ( .A(_528_), .B(_175_), .C(_547_), .Y(_548_) );
AOI21X1 AOI21X1_537 ( .A(_510_), .B(_179_), .C(_548_), .Y(_549_) );
OAI21X1 OAI21X1_1535 ( .A(_543_), .B(_472_), .C(_549_), .Y(_550_) );
AOI21X1 AOI21X1_538 ( .A(_403_), .B(_545_), .C(_550_), .Y(_551_) );
NAND2X1 NAND2X1_1016 ( .A(_542_), .B(_551_), .Y(_552_) );
NOR2X1 NOR2X1_269 ( .A(_542_), .B(_551_), .Y(_553_) );
NOR2X1 NOR2X1_270 ( .A(_256__bF_buf2), .B(_553_), .Y(_554_) );
NAND2X1 NAND2X1_1017 ( .A(_552_), .B(_554_), .Y(_555_) );
NAND2X1 NAND2X1_1018 ( .A(_182_), .B(_185_), .Y(_556_) );
NAND2X1 NAND2X1_1019 ( .A(_175_), .B(_178_), .Y(_557_) );
NOR2X1 NOR2X1_271 ( .A(_556_), .B(_557_), .Y(_558_) );
NAND2X1 NAND2X1_1020 ( .A(_558_), .B(_484_), .Y(_559_) );
AOI21X1 AOI21X1_539 ( .A(_175_), .B(_177_), .C(_174_), .Y(_560_) );
OAI21X1 OAI21X1_1536 ( .A(_557_), .B(_516_), .C(_560_), .Y(_561_) );
AOI21X1 AOI21X1_540 ( .A(_558_), .B(_482_), .C(_561_), .Y(_562_) );
OAI21X1 OAI21X1_1537 ( .A(_559_), .B(_389_), .C(_562_), .Y(_563_) );
INVX1 INVX1_332 ( .A(_563_), .Y(_564_) );
NOR2X1 NOR2X1_272 ( .A(_115_), .B(_564_), .Y(_565_) );
NOR2X1 NOR2X1_273 ( .A(_277__bF_buf0), .B(_565_), .Y(_566_) );
OAI21X1 OAI21X1_1538 ( .A(_542_), .B(_563_), .C(_566_), .Y(_567_) );
OAI22X1 OAI22X1_123 ( .A(_114_), .B(_245__bF_buf2), .C(_115_), .D(_240__bF_buf1), .Y(_568_) );
OAI21X1 OAI21X1_1539 ( .A(datapath_1_ALU_aluInA_16_), .B(datapath_1_ALU_aluInB_16_), .C(_237__bF_buf2), .Y(_569_) );
OAI21X1 OAI21X1_1540 ( .A(_113_), .B(_247_), .C(_569_), .Y(_570_) );
NOR2X1 NOR2X1_274 ( .A(_568_), .B(_570_), .Y(_571_) );
NAND3X1 NAND3X1_1388 ( .A(_555_), .B(_571_), .C(_567_), .Y(datapath_1_ALU_aluResult_16_) );
NAND2X1 NAND2X1_1021 ( .A(_109_), .B(_107_), .Y(_572_) );
OAI21X1 OAI21X1_1541 ( .A(_111_), .B(_112_), .C(_572_), .Y(_573_) );
INVX1 INVX1_333 ( .A(_572_), .Y(_574_) );
INVX1 INVX1_334 ( .A(_114_), .Y(_575_) );
OAI21X1 OAI21X1_1542 ( .A(_575_), .B(_565_), .C(_574_), .Y(_576_) );
OAI21X1 OAI21X1_1543 ( .A(_565_), .B(_573_), .C(_576_), .Y(_577_) );
OAI21X1 OAI21X1_1544 ( .A(_111_), .B(datapath_1_ALU_aluInB_16_), .C(_574_), .Y(_578_) );
NAND2X1 NAND2X1_1022 ( .A(datapath_1_ALU_aluInA_16_), .B(_112_), .Y(_579_) );
OAI21X1 OAI21X1_1545 ( .A(_574_), .B(_579_), .C(_257_), .Y(_580_) );
AOI21X1 AOI21X1_541 ( .A(_553_), .B(_572_), .C(_580_), .Y(_581_) );
OAI21X1 OAI21X1_1546 ( .A(_553_), .B(_578_), .C(_581_), .Y(_582_) );
AOI22X1 AOI22X1_123 ( .A(_110_), .B(_246_), .C(_574_), .D(_241_), .Y(_583_) );
OAI21X1 OAI21X1_1547 ( .A(_108_), .B(_238_), .C(_583_), .Y(_584_) );
AOI21X1 AOI21X1_542 ( .A(_108_), .B(_248__bF_buf3), .C(_584_), .Y(_585_) );
AND2X2 AND2X2_24 ( .A(_582_), .B(_585_), .Y(_586_) );
OAI21X1 OAI21X1_1548 ( .A(_277__bF_buf1), .B(_577_), .C(_586_), .Y(datapath_1_ALU_aluResult_17_) );
NOR2X1 NOR2X1_275 ( .A(_121_), .B(_124_), .Y(_587_) );
INVX1 INVX1_335 ( .A(_587_), .Y(_588_) );
AOI21X1 AOI21X1_543 ( .A(_107_), .B(_109_), .C(_579_), .Y(_589_) );
NOR2X1 NOR2X1_276 ( .A(datapath_1_ALU_aluInB_17_), .B(_105_), .Y(_590_) );
NOR2X1 NOR2X1_277 ( .A(_590_), .B(_589_), .Y(_591_) );
OAI21X1 OAI21X1_1549 ( .A(_116_), .B(_551_), .C(_591_), .Y(_592_) );
AOI21X1 AOI21X1_544 ( .A(_592_), .B(_588_), .C(_256__bF_buf0), .Y(_593_) );
OAI21X1 OAI21X1_1550 ( .A(_588_), .B(_592_), .C(_593_), .Y(_594_) );
NOR2X1 NOR2X1_278 ( .A(_572_), .B(_115_), .Y(_595_) );
INVX1 INVX1_336 ( .A(_595_), .Y(_596_) );
NOR2X1 NOR2X1_279 ( .A(_596_), .B(_564_), .Y(_597_) );
AOI21X1 AOI21X1_545 ( .A(_575_), .B(_107_), .C(_110_), .Y(_598_) );
INVX1 INVX1_337 ( .A(_598_), .Y(_599_) );
NOR2X1 NOR2X1_280 ( .A(_599_), .B(_597_), .Y(_600_) );
AOI21X1 AOI21X1_546 ( .A(_600_), .B(_588_), .C(_277__bF_buf1), .Y(_601_) );
OAI21X1 OAI21X1_1551 ( .A(_588_), .B(_600_), .C(_601_), .Y(_602_) );
NAND2X1 NAND2X1_1023 ( .A(_124_), .B(_246_), .Y(_603_) );
OAI21X1 OAI21X1_1552 ( .A(_240__bF_buf3), .B(_588_), .C(_603_), .Y(_604_) );
NAND2X1 NAND2X1_1024 ( .A(_121_), .B(_248__bF_buf3), .Y(_605_) );
OAI21X1 OAI21X1_1553 ( .A(_121_), .B(_238_), .C(_605_), .Y(_606_) );
NOR2X1 NOR2X1_281 ( .A(_604_), .B(_606_), .Y(_607_) );
NAND3X1 NAND3X1_1389 ( .A(_594_), .B(_607_), .C(_602_), .Y(datapath_1_ALU_aluResult_18_) );
OAI21X1 OAI21X1_1554 ( .A(_121_), .B(_124_), .C(_592_), .Y(_608_) );
OAI21X1 OAI21X1_1555 ( .A(_122_), .B(datapath_1_ALU_aluInB_18_), .C(_608_), .Y(_609_) );
AOI21X1 AOI21X1_547 ( .A(_609_), .B(_120_), .C(_256__bF_buf0), .Y(_610_) );
OAI21X1 OAI21X1_1556 ( .A(_120_), .B(_609_), .C(_610_), .Y(_611_) );
OAI21X1 OAI21X1_1557 ( .A(_599_), .B(_597_), .C(_587_), .Y(_612_) );
OAI21X1 OAI21X1_1558 ( .A(_122_), .B(_123_), .C(_612_), .Y(_613_) );
AOI21X1 AOI21X1_548 ( .A(_613_), .B(_119_), .C(_277__bF_buf1), .Y(_614_) );
OAI21X1 OAI21X1_1559 ( .A(_119_), .B(_613_), .C(_614_), .Y(_615_) );
NAND2X1 NAND2X1_1025 ( .A(_118_), .B(_246_), .Y(_616_) );
OAI21X1 OAI21X1_1560 ( .A(_120_), .B(_240__bF_buf1), .C(_616_), .Y(_617_) );
NAND2X1 NAND2X1_1026 ( .A(_117_), .B(_248__bF_buf2), .Y(_618_) );
OAI21X1 OAI21X1_1561 ( .A(_117_), .B(_238_), .C(_618_), .Y(_619_) );
NOR2X1 NOR2X1_282 ( .A(_617_), .B(_619_), .Y(_620_) );
NAND3X1 NAND3X1_1390 ( .A(_611_), .B(_620_), .C(_615_), .Y(datapath_1_ALU_aluResult_19_) );
NOR2X1 NOR2X1_283 ( .A(_119_), .B(_587_), .Y(_621_) );
OAI21X1 OAI21X1_1562 ( .A(_589_), .B(_590_), .C(_621_), .Y(_622_) );
INVX1 INVX1_338 ( .A(datapath_1_ALU_aluInB_19_), .Y(_623_) );
NAND2X1 NAND2X1_1027 ( .A(datapath_1_ALU_aluInA_19_), .B(_623_), .Y(_624_) );
NAND3X1 NAND3X1_1391 ( .A(datapath_1_ALU_aluInA_18_), .B(_123_), .C(_120_), .Y(_625_) );
NAND3X1 NAND3X1_1392 ( .A(_624_), .B(_625_), .C(_622_), .Y(_626_) );
INVX1 INVX1_339 ( .A(_626_), .Y(_627_) );
OAI21X1 OAI21X1_1563 ( .A(_126_), .B(_551_), .C(_627_), .Y(_628_) );
AND2X2 AND2X2_25 ( .A(_628_), .B(_95_), .Y(_629_) );
NOR2X1 NOR2X1_284 ( .A(_256__bF_buf3), .B(_629_), .Y(_630_) );
OAI21X1 OAI21X1_1564 ( .A(_95_), .B(_628_), .C(_630_), .Y(_631_) );
NAND2X1 NAND2X1_1028 ( .A(_119_), .B(_587_), .Y(_632_) );
AOI21X1 AOI21X1_549 ( .A(_119_), .B(_124_), .C(_118_), .Y(_633_) );
OAI21X1 OAI21X1_1565 ( .A(_598_), .B(_632_), .C(_633_), .Y(_634_) );
NOR2X1 NOR2X1_285 ( .A(_632_), .B(_596_), .Y(_635_) );
AOI21X1 AOI21X1_550 ( .A(_563_), .B(_635_), .C(_634_), .Y(_636_) );
AOI21X1 AOI21X1_551 ( .A(_636_), .B(_95_), .C(_277__bF_buf0), .Y(_637_) );
OAI21X1 OAI21X1_1566 ( .A(_95_), .B(_636_), .C(_637_), .Y(_638_) );
OAI22X1 OAI22X1_124 ( .A(_94_), .B(_245__bF_buf2), .C(_95_), .D(_240__bF_buf0), .Y(_639_) );
OAI21X1 OAI21X1_1567 ( .A(datapath_1_ALU_aluInA_20_), .B(datapath_1_ALU_aluInB_20_), .C(_237__bF_buf0), .Y(_640_) );
OAI21X1 OAI21X1_1568 ( .A(_93_), .B(_247_), .C(_640_), .Y(_641_) );
NOR2X1 NOR2X1_286 ( .A(_639_), .B(_641_), .Y(_642_) );
NAND3X1 NAND3X1_1393 ( .A(_638_), .B(_642_), .C(_631_), .Y(datapath_1_ALU_aluResult_20_) );
OAI21X1 OAI21X1_1569 ( .A(_95_), .B(_636_), .C(_94_), .Y(_643_) );
AOI21X1 AOI21X1_552 ( .A(_643_), .B(_102_), .C(_277__bF_buf0), .Y(_644_) );
OAI21X1 OAI21X1_1570 ( .A(_102_), .B(_643_), .C(_644_), .Y(_645_) );
OAI21X1 OAI21X1_1571 ( .A(_91_), .B(datapath_1_ALU_aluInB_20_), .C(_102_), .Y(_646_) );
NAND3X1 NAND3X1_1394 ( .A(datapath_1_ALU_aluInA_20_), .B(_92_), .C(_101_), .Y(_647_) );
NAND2X1 NAND2X1_1029 ( .A(_647_), .B(_257_), .Y(_648_) );
AOI21X1 AOI21X1_553 ( .A(_628_), .B(_103_), .C(_648_), .Y(_649_) );
OAI21X1 OAI21X1_1572 ( .A(_646_), .B(_629_), .C(_649_), .Y(_650_) );
OAI21X1 OAI21X1_1573 ( .A(datapath_1_ALU_aluInA_21_), .B(datapath_1_ALU_aluInB_21_), .C(_237__bF_buf0), .Y(_651_) );
OAI21X1 OAI21X1_1574 ( .A(_99_), .B(_247_), .C(_651_), .Y(_652_) );
OAI22X1 OAI22X1_125 ( .A(_100_), .B(_245__bF_buf1), .C(_101_), .D(_240__bF_buf0), .Y(_653_) );
NOR2X1 NOR2X1_287 ( .A(_653_), .B(_652_), .Y(_654_) );
NAND3X1 NAND3X1_1395 ( .A(_650_), .B(_654_), .C(_645_), .Y(datapath_1_ALU_aluResult_21_) );
NAND2X1 NAND2X1_1030 ( .A(_103_), .B(_628_), .Y(_655_) );
OAI21X1 OAI21X1_1575 ( .A(_97_), .B(datapath_1_ALU_aluInB_21_), .C(_647_), .Y(_656_) );
INVX1 INVX1_340 ( .A(_656_), .Y(_657_) );
NAND2X1 NAND2X1_1031 ( .A(_657_), .B(_655_), .Y(_658_) );
AOI21X1 AOI21X1_554 ( .A(_655_), .B(_657_), .C(_89_), .Y(_659_) );
NOR2X1 NOR2X1_288 ( .A(_256__bF_buf3), .B(_659_), .Y(_660_) );
OAI21X1 OAI21X1_1576 ( .A(_88_), .B(_658_), .C(_660_), .Y(_661_) );
NAND2X1 NAND2X1_1032 ( .A(_96_), .B(_102_), .Y(_662_) );
INVX1 INVX1_341 ( .A(_100_), .Y(_663_) );
NOR2X1 NOR2X1_289 ( .A(_94_), .B(_101_), .Y(_664_) );
NOR2X1 NOR2X1_290 ( .A(_663_), .B(_664_), .Y(_665_) );
OAI21X1 OAI21X1_1577 ( .A(_662_), .B(_636_), .C(_665_), .Y(_666_) );
AND2X2 AND2X2_26 ( .A(_666_), .B(_89_), .Y(_667_) );
OAI21X1 OAI21X1_1578 ( .A(_89_), .B(_666_), .C(_260_), .Y(_668_) );
OR2X2 OR2X2_11 ( .A(_668_), .B(_667_), .Y(_669_) );
OAI22X1 OAI22X1_126 ( .A(_87_), .B(_245__bF_buf1), .C(_88_), .D(_240__bF_buf4), .Y(_670_) );
OAI21X1 OAI21X1_1579 ( .A(datapath_1_ALU_aluInA_22_), .B(datapath_1_ALU_aluInB_22_), .C(_237__bF_buf0), .Y(_671_) );
OAI21X1 OAI21X1_1580 ( .A(_86_), .B(_247_), .C(_671_), .Y(_672_) );
NOR2X1 NOR2X1_291 ( .A(_670_), .B(_672_), .Y(_673_) );
NAND3X1 NAND3X1_1396 ( .A(_669_), .B(_673_), .C(_661_), .Y(datapath_1_ALU_aluResult_22_) );
NOR2X1 NOR2X1_292 ( .A(datapath_1_ALU_aluInB_22_), .B(_84_), .Y(_674_) );
NOR2X1 NOR2X1_293 ( .A(_674_), .B(_659_), .Y(_675_) );
NAND2X1 NAND2X1_1033 ( .A(_83_), .B(_675_), .Y(_676_) );
OAI21X1 OAI21X1_1581 ( .A(_674_), .B(_659_), .C(_82_), .Y(_677_) );
NAND3X1 NAND3X1_1397 ( .A(_257_), .B(_677_), .C(_676_), .Y(_678_) );
INVX1 INVX1_342 ( .A(_87_), .Y(_679_) );
NOR2X1 NOR2X1_294 ( .A(_679_), .B(_667_), .Y(_680_) );
NAND2X1 NAND2X1_1034 ( .A(_82_), .B(_680_), .Y(_681_) );
OAI21X1 OAI21X1_1582 ( .A(_679_), .B(_667_), .C(_83_), .Y(_682_) );
NAND3X1 NAND3X1_1398 ( .A(_260_), .B(_682_), .C(_681_), .Y(_683_) );
OAI22X1 OAI22X1_127 ( .A(_81_), .B(_245__bF_buf3), .C(_82_), .D(_240__bF_buf4), .Y(_684_) );
OAI21X1 OAI21X1_1583 ( .A(datapath_1_ALU_aluInA_23_), .B(datapath_1_ALU_aluInB_23_), .C(_237__bF_buf0), .Y(_685_) );
OAI21X1 OAI21X1_1584 ( .A(_80_), .B(_247_), .C(_685_), .Y(_686_) );
NOR2X1 NOR2X1_295 ( .A(_684_), .B(_686_), .Y(_687_) );
NAND3X1 NAND3X1_1399 ( .A(_687_), .B(_678_), .C(_683_), .Y(datapath_1_ALU_aluResult_23_) );
NOR2X1 NOR2X1_296 ( .A(_138_), .B(_140_), .Y(_688_) );
INVX1 INVX1_343 ( .A(_688_), .Y(_689_) );
OR2X2 OR2X2_12 ( .A(_126_), .B(_104_), .Y(_690_) );
INVX1 INVX1_344 ( .A(_104_), .Y(_691_) );
NAND2X1 NAND2X1_1035 ( .A(_90_), .B(_656_), .Y(_692_) );
NAND2X1 NAND2X1_1036 ( .A(_674_), .B(_82_), .Y(_693_) );
INVX1 INVX1_345 ( .A(datapath_1_ALU_aluInB_23_), .Y(_694_) );
NAND2X1 NAND2X1_1037 ( .A(datapath_1_ALU_aluInA_23_), .B(_694_), .Y(_695_) );
NAND3X1 NAND3X1_1400 ( .A(_693_), .B(_695_), .C(_692_), .Y(_696_) );
AOI21X1 AOI21X1_555 ( .A(_626_), .B(_691_), .C(_696_), .Y(_697_) );
OAI21X1 OAI21X1_1585 ( .A(_690_), .B(_551_), .C(_697_), .Y(_698_) );
OAI21X1 OAI21X1_1586 ( .A(_138_), .B(_140_), .C(_698_), .Y(_699_) );
INVX1 INVX1_346 ( .A(_699_), .Y(_700_) );
NOR2X1 NOR2X1_297 ( .A(_256__bF_buf2), .B(_700_), .Y(_701_) );
OAI21X1 OAI21X1_1587 ( .A(_689_), .B(_698_), .C(_701_), .Y(_702_) );
NOR2X1 NOR2X1_298 ( .A(_82_), .B(_88_), .Y(_703_) );
INVX1 INVX1_347 ( .A(_703_), .Y(_704_) );
NOR2X1 NOR2X1_299 ( .A(_662_), .B(_704_), .Y(_705_) );
NAND2X1 NAND2X1_1038 ( .A(_634_), .B(_705_), .Y(_706_) );
OAI21X1 OAI21X1_1588 ( .A(_94_), .B(_101_), .C(_100_), .Y(_707_) );
OAI21X1 OAI21X1_1589 ( .A(_87_), .B(_82_), .C(_81_), .Y(_708_) );
AOI21X1 AOI21X1_556 ( .A(_707_), .B(_703_), .C(_708_), .Y(_709_) );
NAND2X1 NAND2X1_1039 ( .A(_709_), .B(_706_), .Y(_710_) );
AND2X2 AND2X2_27 ( .A(_635_), .B(_705_), .Y(_711_) );
AOI21X1 AOI21X1_557 ( .A(_563_), .B(_711_), .C(_710_), .Y(_712_) );
AOI21X1 AOI21X1_558 ( .A(_712_), .B(_689_), .C(_277__bF_buf1), .Y(_713_) );
OAI21X1 OAI21X1_1590 ( .A(_689_), .B(_712_), .C(_713_), .Y(_714_) );
OAI22X1 OAI22X1_128 ( .A(_139_), .B(_245__bF_buf2), .C(_240__bF_buf3), .D(_689_), .Y(_715_) );
NAND2X1 NAND2X1_1040 ( .A(_138_), .B(_248__bF_buf3), .Y(_716_) );
OAI21X1 OAI21X1_1591 ( .A(_138_), .B(_238_), .C(_716_), .Y(_717_) );
NOR2X1 NOR2X1_300 ( .A(_715_), .B(_717_), .Y(_718_) );
NAND3X1 NAND3X1_1401 ( .A(_714_), .B(_718_), .C(_702_), .Y(datapath_1_ALU_aluResult_24_) );
INVX1 INVX1_348 ( .A(_145_), .Y(_719_) );
OAI21X1 OAI21X1_1592 ( .A(_138_), .B(_712_), .C(_139_), .Y(_720_) );
AOI21X1 AOI21X1_559 ( .A(_720_), .B(_719_), .C(_277__bF_buf1), .Y(_721_) );
OAI21X1 OAI21X1_1593 ( .A(_719_), .B(_720_), .C(_721_), .Y(_722_) );
INVX1 INVX1_349 ( .A(datapath_1_ALU_aluInB_24_), .Y(_723_) );
NAND2X1 NAND2X1_1041 ( .A(datapath_1_ALU_aluInA_24_), .B(_723_), .Y(_724_) );
OAI21X1 OAI21X1_1594 ( .A(_142_), .B(_144_), .C(_724_), .Y(_725_) );
OAI21X1 OAI21X1_1595 ( .A(_719_), .B(_724_), .C(_257_), .Y(_726_) );
AOI21X1 AOI21X1_560 ( .A(_698_), .B(_147_), .C(_726_), .Y(_727_) );
OAI21X1 OAI21X1_1596 ( .A(_725_), .B(_700_), .C(_727_), .Y(_728_) );
NOR2X1 NOR2X1_301 ( .A(_143_), .B(_141_), .Y(_729_) );
NAND2X1 NAND2X1_1042 ( .A(_729_), .B(_246_), .Y(_730_) );
OAI21X1 OAI21X1_1597 ( .A(_145_), .B(_240__bF_buf3), .C(_730_), .Y(_731_) );
NAND2X1 NAND2X1_1043 ( .A(_143_), .B(_141_), .Y(_732_) );
OAI21X1 OAI21X1_1598 ( .A(datapath_1_ALU_aluInA_25_), .B(datapath_1_ALU_aluInB_25_), .C(_237__bF_buf1), .Y(_733_) );
OAI21X1 OAI21X1_1599 ( .A(_247_), .B(_732_), .C(_733_), .Y(_734_) );
NOR2X1 NOR2X1_302 ( .A(_731_), .B(_734_), .Y(_735_) );
NAND3X1 NAND3X1_1402 ( .A(_728_), .B(_735_), .C(_722_), .Y(datapath_1_ALU_aluResult_25_) );
OAI21X1 OAI21X1_1600 ( .A(_142_), .B(_144_), .C(_688_), .Y(_736_) );
AOI21X1 AOI21X1_561 ( .A(_719_), .B(_140_), .C(_729_), .Y(_737_) );
OAI21X1 OAI21X1_1601 ( .A(_736_), .B(_712_), .C(_737_), .Y(_738_) );
AND2X2 AND2X2_28 ( .A(_738_), .B(_136_), .Y(_739_) );
OAI21X1 OAI21X1_1602 ( .A(_136_), .B(_738_), .C(_260_), .Y(_740_) );
INVX1 INVX1_350 ( .A(_136_), .Y(_741_) );
INVX1 INVX1_351 ( .A(_144_), .Y(_742_) );
OAI21X1 OAI21X1_1603 ( .A(_142_), .B(_724_), .C(_742_), .Y(_743_) );
INVX1 INVX1_352 ( .A(_743_), .Y(_744_) );
OAI21X1 OAI21X1_1604 ( .A(_719_), .B(_699_), .C(_744_), .Y(_745_) );
NAND2X1 NAND2X1_1044 ( .A(_147_), .B(_698_), .Y(_746_) );
AOI21X1 AOI21X1_562 ( .A(_746_), .B(_744_), .C(_136_), .Y(_747_) );
NOR2X1 NOR2X1_303 ( .A(_256__bF_buf2), .B(_747_), .Y(_748_) );
OAI21X1 OAI21X1_1605 ( .A(_741_), .B(_745_), .C(_748_), .Y(_749_) );
INVX1 INVX1_353 ( .A(_135_), .Y(_750_) );
OAI22X1 OAI22X1_129 ( .A(_750_), .B(_245__bF_buf2), .C(_240__bF_buf3), .D(_741_), .Y(_751_) );
NAND2X1 NAND2X1_1045 ( .A(_132_), .B(_248__bF_buf3), .Y(_752_) );
OAI21X1 OAI21X1_1606 ( .A(_132_), .B(_238_), .C(_752_), .Y(_753_) );
NOR2X1 NOR2X1_304 ( .A(_751_), .B(_753_), .Y(_754_) );
AND2X2 AND2X2_29 ( .A(_749_), .B(_754_), .Y(_755_) );
OAI21X1 OAI21X1_1607 ( .A(_739_), .B(_740_), .C(_755_), .Y(datapath_1_ALU_aluResult_26_) );
NOR2X1 NOR2X1_305 ( .A(datapath_1_ALU_aluInB_26_), .B(_133_), .Y(_756_) );
NOR2X1 NOR2X1_306 ( .A(_756_), .B(_747_), .Y(_757_) );
AOI21X1 AOI21X1_563 ( .A(_757_), .B(_131_), .C(_256__bF_buf2), .Y(_758_) );
OAI21X1 OAI21X1_1608 ( .A(_131_), .B(_757_), .C(_758_), .Y(_759_) );
NOR2X1 NOR2X1_307 ( .A(_135_), .B(_739_), .Y(_760_) );
OAI21X1 OAI21X1_1609 ( .A(_128_), .B(_130_), .C(_760_), .Y(_761_) );
OAI21X1 OAI21X1_1610 ( .A(_135_), .B(_739_), .C(_131_), .Y(_762_) );
NAND3X1 NAND3X1_1403 ( .A(_260_), .B(_762_), .C(_761_), .Y(_763_) );
NAND2X1 NAND2X1_1046 ( .A(_131_), .B(_241_), .Y(_764_) );
OAI21X1 OAI21X1_1611 ( .A(_129_), .B(_245__bF_buf0), .C(_764_), .Y(_765_) );
NAND2X1 NAND2X1_1047 ( .A(_128_), .B(_248__bF_buf3), .Y(_766_) );
OAI21X1 OAI21X1_1612 ( .A(_128_), .B(_238_), .C(_766_), .Y(_767_) );
NOR2X1 NOR2X1_308 ( .A(_765_), .B(_767_), .Y(_768_) );
NAND3X1 NAND3X1_1404 ( .A(_763_), .B(_768_), .C(_759_), .Y(datapath_1_ALU_aluResult_27_) );
NOR2X1 NOR2X1_309 ( .A(_165_), .B(_168_), .Y(_769_) );
INVX1 INVX1_354 ( .A(_148_), .Y(_770_) );
NAND2X1 NAND2X1_1048 ( .A(_743_), .B(_137_), .Y(_771_) );
OAI21X1 OAI21X1_1613 ( .A(_128_), .B(_130_), .C(_756_), .Y(_772_) );
INVX1 INVX1_355 ( .A(datapath_1_ALU_aluInB_27_), .Y(_773_) );
NAND2X1 NAND2X1_1049 ( .A(datapath_1_ALU_aluInA_27_), .B(_773_), .Y(_774_) );
NAND3X1 NAND3X1_1405 ( .A(_772_), .B(_774_), .C(_771_), .Y(_775_) );
AOI21X1 AOI21X1_564 ( .A(_698_), .B(_770_), .C(_775_), .Y(_776_) );
AND2X2 AND2X2_30 ( .A(_776_), .B(_769_), .Y(_777_) );
OAI21X1 OAI21X1_1614 ( .A(_769_), .B(_776_), .C(_257_), .Y(_778_) );
NAND2X1 NAND2X1_1050 ( .A(_131_), .B(_136_), .Y(_779_) );
NOR2X1 NOR2X1_310 ( .A(_736_), .B(_779_), .Y(_780_) );
INVX1 INVX1_356 ( .A(_780_), .Y(_781_) );
NOR2X1 NOR2X1_311 ( .A(_779_), .B(_737_), .Y(_782_) );
OAI21X1 OAI21X1_1615 ( .A(_128_), .B(_750_), .C(_129_), .Y(_783_) );
NOR2X1 NOR2X1_312 ( .A(_783_), .B(_782_), .Y(_784_) );
OAI21X1 OAI21X1_1616 ( .A(_781_), .B(_712_), .C(_784_), .Y(_785_) );
INVX1 INVX1_357 ( .A(_769_), .Y(_786_) );
NOR2X1 NOR2X1_313 ( .A(_212_), .B(_331_), .Y(_787_) );
NOR2X1 NOR2X1_314 ( .A(_206_), .B(_350_), .Y(_788_) );
NAND2X1 NAND2X1_1051 ( .A(_787_), .B(_788_), .Y(_789_) );
AOI21X1 AOI21X1_565 ( .A(_312_), .B(_313_), .C(_789_), .Y(_790_) );
AND2X2 AND2X2_31 ( .A(_484_), .B(_558_), .Y(_791_) );
OAI21X1 OAI21X1_1617 ( .A(_388_), .B(_790_), .C(_791_), .Y(_792_) );
NAND2X1 NAND2X1_1052 ( .A(_705_), .B(_635_), .Y(_793_) );
AOI21X1 AOI21X1_566 ( .A(_792_), .B(_562_), .C(_793_), .Y(_794_) );
OAI21X1 OAI21X1_1618 ( .A(_710_), .B(_794_), .C(_780_), .Y(_795_) );
AOI21X1 AOI21X1_567 ( .A(_795_), .B(_784_), .C(_786_), .Y(_796_) );
NOR2X1 NOR2X1_315 ( .A(_277__bF_buf3), .B(_796_), .Y(_797_) );
OAI21X1 OAI21X1_1619 ( .A(_769_), .B(_785_), .C(_797_), .Y(_798_) );
INVX1 INVX1_358 ( .A(_165_), .Y(_799_) );
AOI22X1 AOI22X1_124 ( .A(_168_), .B(_246_), .C(_799_), .D(_237__bF_buf1), .Y(_800_) );
OAI21X1 OAI21X1_1620 ( .A(_786_), .B(_240__bF_buf3), .C(_800_), .Y(_801_) );
AOI21X1 AOI21X1_568 ( .A(_165_), .B(_248__bF_buf1), .C(_801_), .Y(_802_) );
AND2X2 AND2X2_32 ( .A(_798_), .B(_802_), .Y(_803_) );
OAI21X1 OAI21X1_1621 ( .A(_777_), .B(_778_), .C(_803_), .Y(datapath_1_ALU_aluResult_28_) );
INVX1 INVX1_359 ( .A(_168_), .Y(_804_) );
OAI21X1 OAI21X1_1622 ( .A(_160_), .B(_162_), .C(_804_), .Y(_805_) );
OAI21X1 OAI21X1_1623 ( .A(_168_), .B(_796_), .C(_163_), .Y(_806_) );
OAI21X1 OAI21X1_1624 ( .A(_796_), .B(_805_), .C(_806_), .Y(_807_) );
NAND2X1 NAND2X1_1053 ( .A(datapath_1_ALU_aluInA_28_), .B(_167_), .Y(_808_) );
OAI21X1 OAI21X1_1625 ( .A(_769_), .B(_776_), .C(_808_), .Y(_809_) );
OAI21X1 OAI21X1_1626 ( .A(_321_), .B(_295_), .C(_216_), .Y(_810_) );
AOI21X1 AOI21X1_569 ( .A(_810_), .B(_402_), .C(_201_), .Y(_811_) );
OAI21X1 OAI21X1_1627 ( .A(_550_), .B(_811_), .C(_127_), .Y(_812_) );
AOI21X1 AOI21X1_570 ( .A(_812_), .B(_697_), .C(_148_), .Y(_813_) );
OAI21X1 OAI21X1_1628 ( .A(_775_), .B(_813_), .C(_170_), .Y(_814_) );
NOR2X1 NOR2X1_316 ( .A(_808_), .B(_163_), .Y(_815_) );
NOR2X1 NOR2X1_317 ( .A(_256__bF_buf3), .B(_815_), .Y(_816_) );
AND2X2 AND2X2_33 ( .A(_814_), .B(_816_), .Y(_817_) );
OAI21X1 OAI21X1_1629 ( .A(_164_), .B(_809_), .C(_817_), .Y(_818_) );
MUX2X1 MUX2X1_127 ( .A(_248__bF_buf1), .B(_237__bF_buf1), .S(_160_), .Y(_819_) );
OAI21X1 OAI21X1_1630 ( .A(_161_), .B(_245__bF_buf0), .C(_819_), .Y(_820_) );
AOI21X1 AOI21X1_571 ( .A(_163_), .B(_241_), .C(_820_), .Y(_821_) );
AND2X2 AND2X2_34 ( .A(_818_), .B(_821_), .Y(_822_) );
OAI21X1 OAI21X1_1631 ( .A(_277__bF_buf3), .B(_807_), .C(_822_), .Y(datapath_1_ALU_aluResult_29_) );
INVX1 INVX1_360 ( .A(datapath_1_ALU_aluInB_29_), .Y(_823_) );
AOI21X1 AOI21X1_572 ( .A(datapath_1_ALU_aluInA_29_), .B(_823_), .C(_815_), .Y(_824_) );
OAI21X1 OAI21X1_1632 ( .A(_169_), .B(_776_), .C(_824_), .Y(_825_) );
INVX1 INVX1_361 ( .A(_149_), .Y(_826_) );
INVX1 INVX1_362 ( .A(_152_), .Y(_827_) );
AOI22X1 AOI22X1_125 ( .A(_826_), .B(_827_), .C(_824_), .D(_814_), .Y(_828_) );
NOR2X1 NOR2X1_318 ( .A(_256__bF_buf3), .B(_828_), .Y(_829_) );
OAI21X1 OAI21X1_1633 ( .A(_154_), .B(_825_), .C(_829_), .Y(_830_) );
NOR2X1 NOR2X1_319 ( .A(_164_), .B(_786_), .Y(_831_) );
OAI21X1 OAI21X1_1634 ( .A(_160_), .B(_804_), .C(_161_), .Y(_832_) );
AOI21X1 AOI21X1_573 ( .A(_785_), .B(_831_), .C(_832_), .Y(_833_) );
AOI21X1 AOI21X1_574 ( .A(_833_), .B(_154_), .C(_277__bF_buf3), .Y(_834_) );
OAI21X1 OAI21X1_1635 ( .A(_154_), .B(_833_), .C(_834_), .Y(_835_) );
OAI22X1 OAI22X1_130 ( .A(_827_), .B(_245__bF_buf0), .C(_240__bF_buf4), .D(_154_), .Y(_836_) );
OAI21X1 OAI21X1_1636 ( .A(datapath_1_ALU_aluInA_30_), .B(datapath_1_ALU_aluInB_30_), .C(_237__bF_buf3), .Y(_837_) );
OAI21X1 OAI21X1_1637 ( .A(_826_), .B(_247_), .C(_837_), .Y(_838_) );
NOR2X1 NOR2X1_320 ( .A(_836_), .B(_838_), .Y(_839_) );
NAND3X1 NAND3X1_1406 ( .A(_835_), .B(_839_), .C(_830_), .Y(datapath_1_ALU_aluResult_30_) );
NAND2X1 NAND2X1_1054 ( .A(_154_), .B(_825_), .Y(_840_) );
NOR2X1 NOR2X1_321 ( .A(datapath_1_ALU_aluInB_30_), .B(_150_), .Y(_841_) );
INVX1 INVX1_363 ( .A(_841_), .Y(_842_) );
NAND3X1 NAND3X1_1407 ( .A(_158_), .B(_842_), .C(_840_), .Y(_843_) );
OAI21X1 OAI21X1_1638 ( .A(_841_), .B(_828_), .C(_159_), .Y(_844_) );
NAND3X1 NAND3X1_1408 ( .A(_257_), .B(_843_), .C(_844_), .Y(_845_) );
INVX1 INVX1_364 ( .A(_831_), .Y(_846_) );
AOI21X1 AOI21X1_575 ( .A(_795_), .B(_784_), .C(_846_), .Y(_847_) );
OAI21X1 OAI21X1_1639 ( .A(_832_), .B(_847_), .C(_153_), .Y(_848_) );
NAND3X1 NAND3X1_1409 ( .A(_827_), .B(_159_), .C(_848_), .Y(_849_) );
OAI21X1 OAI21X1_1640 ( .A(_154_), .B(_833_), .C(_827_), .Y(_850_) );
NAND2X1 NAND2X1_1055 ( .A(_158_), .B(_850_), .Y(_851_) );
NAND3X1 NAND3X1_1410 ( .A(_260_), .B(_849_), .C(_851_), .Y(_852_) );
OAI22X1 OAI22X1_131 ( .A(_156_), .B(_245__bF_buf0), .C(_240__bF_buf4), .D(_159_), .Y(_853_) );
NAND2X1 NAND2X1_1056 ( .A(_155_), .B(_248__bF_buf1), .Y(_854_) );
OAI21X1 OAI21X1_1641 ( .A(_155_), .B(_238_), .C(_854_), .Y(_855_) );
NOR2X1 NOR2X1_322 ( .A(_853_), .B(_855_), .Y(_856_) );
NAND3X1 NAND3X1_1411 ( .A(_856_), .B(_852_), .C(_845_), .Y(datapath_1_ALU_aluResult_31_) );
INVX1 INVX1_365 ( .A(PCWrite), .Y(_857_) );
NAND2X1 NAND2X1_1057 ( .A(datapath_1_ALU_aluZero), .B(PCWriteCond), .Y(_858_) );
NAND2X1 NAND2X1_1058 ( .A(_857_), .B(_858_), .Y(datapath_1_PCEn) );
NOR2X1 NOR2X1_323 ( .A(datapath_1_Instr_25_bF_buf3_), .B(datapath_1_Instr_21_bF_buf53_), .Y(_1883_) );
INVX1 INVX1_366 ( .A(datapath_1_Instr_22_bF_buf48_), .Y(_1884_) );
INVX1 INVX1_367 ( .A(datapath_1_Instr_23_bF_buf13_bF_buf3_), .Y(_1885_) );
NAND2X1 NAND2X1_1059 ( .A(_1884__bF_buf2), .B(_1885__bF_buf7), .Y(_1886_) );
NOR2X1 NOR2X1_324 ( .A(datapath_1_Instr_24_bF_buf4_), .B(_1886_), .Y(_1887_) );
INVX1 INVX1_368 ( .A(datapath_1_Instr_24_bF_buf3_), .Y(_1888_) );
NAND2X1 NAND2X1_1060 ( .A(datapath_1_Instr_21_bF_buf52_), .B(datapath_1_RegisterFile_regfile_mem_27__0_), .Y(_1889_) );
INVX1 INVX1_369 ( .A(datapath_1_Instr_21_bF_buf51_), .Y(_1890_) );
NAND2X1 NAND2X1_1061 ( .A(datapath_1_RegisterFile_regfile_mem_26__0_), .B(_1890__bF_buf1), .Y(_1891_) );
NAND3X1 NAND3X1_1412 ( .A(datapath_1_Instr_22_bF_buf47_), .B(_1889_), .C(_1891_), .Y(_1892_) );
NAND2X1 NAND2X1_1062 ( .A(datapath_1_Instr_21_bF_buf50_), .B(datapath_1_RegisterFile_regfile_mem_25__0_), .Y(_1893_) );
AOI21X1 AOI21X1_576 ( .A(_1890__bF_buf1), .B(datapath_1_RegisterFile_regfile_mem_24__0_), .C(datapath_1_Instr_22_bF_buf46_), .Y(_1894_) );
NAND2X1 NAND2X1_1063 ( .A(_1893_), .B(_1894_), .Y(_1895_) );
NAND3X1 NAND3X1_1413 ( .A(_1885__bF_buf4), .B(_1892_), .C(_1895_), .Y(_1896_) );
NAND2X1 NAND2X1_1064 ( .A(datapath_1_Instr_21_bF_buf49_), .B(datapath_1_RegisterFile_regfile_mem_31__0_), .Y(_1897_) );
AOI21X1 AOI21X1_577 ( .A(_1890__bF_buf7), .B(datapath_1_RegisterFile_regfile_mem_30__0_), .C(_1884__bF_buf9), .Y(_1898_) );
NAND2X1 NAND2X1_1065 ( .A(_1897_), .B(_1898_), .Y(_1899_) );
INVX1 INVX1_370 ( .A(datapath_1_RegisterFile_regfile_mem_28__0_), .Y(_1900_) );
AOI21X1 AOI21X1_578 ( .A(datapath_1_Instr_21_bF_buf48_), .B(datapath_1_RegisterFile_regfile_mem_29__0_), .C(datapath_1_Instr_22_bF_buf45_), .Y(_1901_) );
OAI21X1 OAI21X1_1642 ( .A(datapath_1_Instr_21_bF_buf47_), .B(_1900_), .C(_1901_), .Y(_1902_) );
NAND3X1 NAND3X1_1414 ( .A(datapath_1_Instr_23_bF_buf12_bF_buf3_), .B(_1902_), .C(_1899_), .Y(_1903_) );
AOI21X1 AOI21X1_579 ( .A(_1896_), .B(_1903_), .C(_1888__bF_buf1), .Y(_1904_) );
MUX2X1 MUX2X1_128 ( .A(datapath_1_RegisterFile_regfile_mem_18__0_), .B(datapath_1_RegisterFile_regfile_mem_16__0_), .S(datapath_1_Instr_22_bF_buf44_), .Y(_1905_) );
NAND2X1 NAND2X1_1066 ( .A(_1890__bF_buf9), .B(_1905_), .Y(_1906_) );
MUX2X1 MUX2X1_129 ( .A(datapath_1_RegisterFile_regfile_mem_19__0_), .B(datapath_1_RegisterFile_regfile_mem_17__0_), .S(datapath_1_Instr_22_bF_buf43_), .Y(_1907_) );
NAND2X1 NAND2X1_1067 ( .A(datapath_1_Instr_21_bF_buf46_), .B(_1907_), .Y(_1908_) );
NAND3X1 NAND3X1_1415 ( .A(_1885__bF_buf9), .B(_1906_), .C(_1908_), .Y(_1909_) );
MUX2X1 MUX2X1_130 ( .A(datapath_1_RegisterFile_regfile_mem_22__0_), .B(datapath_1_RegisterFile_regfile_mem_20__0_), .S(datapath_1_Instr_22_bF_buf42_), .Y(_1910_) );
NAND2X1 NAND2X1_1068 ( .A(_1890__bF_buf37), .B(_1910_), .Y(_1911_) );
MUX2X1 MUX2X1_131 ( .A(datapath_1_RegisterFile_regfile_mem_23__0_), .B(datapath_1_RegisterFile_regfile_mem_21__0_), .S(datapath_1_Instr_22_bF_buf41_), .Y(_1912_) );
NAND2X1 NAND2X1_1069 ( .A(datapath_1_Instr_21_bF_buf45_), .B(_1912_), .Y(_1913_) );
NAND3X1 NAND3X1_1416 ( .A(datapath_1_Instr_23_bF_buf11_bF_buf3_), .B(_1911_), .C(_1913_), .Y(_1914_) );
AOI21X1 AOI21X1_580 ( .A(_1909_), .B(_1914_), .C(datapath_1_Instr_24_bF_buf2_), .Y(_1915_) );
OAI21X1 OAI21X1_1643 ( .A(_1915_), .B(_1904_), .C(datapath_1_Instr_25_bF_buf2_), .Y(_1916_) );
INVX1 INVX1_371 ( .A(datapath_1_Instr_25_bF_buf1_), .Y(_1917_) );
INVX1 INVX1_372 ( .A(datapath_1_RegisterFile_regfile_mem_9__0_), .Y(_1918_) );
AOI21X1 AOI21X1_581 ( .A(datapath_1_Instr_23_bF_buf10_bF_buf3_), .B(datapath_1_RegisterFile_regfile_mem_13__0_), .C(_1890__bF_buf20), .Y(_1919_) );
OAI21X1 OAI21X1_1644 ( .A(datapath_1_Instr_23_bF_buf9_bF_buf3_), .B(_1918_), .C(_1919_), .Y(_1920_) );
INVX1 INVX1_373 ( .A(datapath_1_RegisterFile_regfile_mem_8__0_), .Y(_1921_) );
AOI21X1 AOI21X1_582 ( .A(datapath_1_Instr_23_bF_buf8_bF_buf3_), .B(datapath_1_RegisterFile_regfile_mem_12__0_), .C(datapath_1_Instr_21_bF_buf44_), .Y(_1922_) );
OAI21X1 OAI21X1_1645 ( .A(datapath_1_Instr_23_bF_buf7_bF_buf3_), .B(_1921_), .C(_1922_), .Y(_1923_) );
NAND3X1 NAND3X1_1417 ( .A(_1884__bF_buf4), .B(_1923_), .C(_1920_), .Y(_1924_) );
INVX1 INVX1_374 ( .A(datapath_1_RegisterFile_regfile_mem_11__0_), .Y(_1925_) );
AOI21X1 AOI21X1_583 ( .A(datapath_1_Instr_23_bF_buf6_bF_buf3_), .B(datapath_1_RegisterFile_regfile_mem_15__0_), .C(_1890__bF_buf20), .Y(_1926_) );
OAI21X1 OAI21X1_1646 ( .A(datapath_1_Instr_23_bF_buf5_bF_buf3_), .B(_1925_), .C(_1926_), .Y(_1927_) );
INVX1 INVX1_375 ( .A(datapath_1_RegisterFile_regfile_mem_10__0_), .Y(_1928_) );
AOI21X1 AOI21X1_584 ( .A(datapath_1_Instr_23_bF_buf4_bF_buf3_), .B(datapath_1_RegisterFile_regfile_mem_14__0_), .C(datapath_1_Instr_21_bF_buf43_), .Y(_1929_) );
OAI21X1 OAI21X1_1647 ( .A(datapath_1_Instr_23_bF_buf3_bF_buf3_), .B(_1928_), .C(_1929_), .Y(_1930_) );
NAND3X1 NAND3X1_1418 ( .A(datapath_1_Instr_22_bF_buf40_), .B(_1930_), .C(_1927_), .Y(_1931_) );
AOI21X1 AOI21X1_585 ( .A(_1924_), .B(_1931_), .C(_1888__bF_buf5), .Y(_1932_) );
MUX2X1 MUX2X1_132 ( .A(datapath_1_RegisterFile_regfile_mem_1__0_), .B(datapath_1_RegisterFile_regfile_mem_0__0_), .S(datapath_1_Instr_21_bF_buf42_), .Y(_1933_) );
NOR2X1 NOR2X1_325 ( .A(datapath_1_RegisterFile_regfile_mem_3__0_), .B(_1890__bF_buf30), .Y(_1934_) );
OAI21X1 OAI21X1_1648 ( .A(datapath_1_Instr_21_bF_buf41_), .B(datapath_1_RegisterFile_regfile_mem_2__0_), .C(datapath_1_Instr_22_bF_buf39_), .Y(_1935_) );
OAI22X1 OAI22X1_132 ( .A(_1935_), .B(_1934_), .C(datapath_1_Instr_22_bF_buf38_), .D(_1933_), .Y(_1936_) );
NAND2X1 NAND2X1_1070 ( .A(_1885__bF_buf4), .B(_1936_), .Y(_1937_) );
MUX2X1 MUX2X1_133 ( .A(datapath_1_RegisterFile_regfile_mem_5__0_), .B(datapath_1_RegisterFile_regfile_mem_4__0_), .S(datapath_1_Instr_21_bF_buf40_), .Y(_1938_) );
NOR2X1 NOR2X1_326 ( .A(datapath_1_RegisterFile_regfile_mem_7__0_), .B(_1890__bF_buf30), .Y(_1939_) );
OAI21X1 OAI21X1_1649 ( .A(datapath_1_Instr_21_bF_buf39_), .B(datapath_1_RegisterFile_regfile_mem_6__0_), .C(datapath_1_Instr_22_bF_buf37_), .Y(_1940_) );
OAI22X1 OAI22X1_133 ( .A(_1940_), .B(_1939_), .C(datapath_1_Instr_22_bF_buf36_), .D(_1938_), .Y(_1941_) );
NAND2X1 NAND2X1_1071 ( .A(datapath_1_Instr_23_bF_buf2_bF_buf3_), .B(_1941_), .Y(_1942_) );
AOI21X1 AOI21X1_586 ( .A(_1937_), .B(_1942_), .C(datapath_1_Instr_24_bF_buf1_), .Y(_1943_) );
OAI21X1 OAI21X1_1650 ( .A(_1932_), .B(_1943_), .C(_1917__bF_buf0), .Y(_1944_) );
AOI22X1 AOI22X1_126 ( .A(_1883__bF_buf2), .B(_1887__bF_buf4), .C(_1916_), .D(_1944_), .Y(datapath_1_RD1_0_) );
MUX2X1 MUX2X1_134 ( .A(datapath_1_RegisterFile_regfile_mem_9__1_), .B(datapath_1_RegisterFile_regfile_mem_8__1_), .S(datapath_1_Instr_21_bF_buf38_), .Y(_1945_) );
NOR2X1 NOR2X1_327 ( .A(datapath_1_RegisterFile_regfile_mem_11__1_), .B(_1890__bF_buf12), .Y(_1946_) );
OAI21X1 OAI21X1_1651 ( .A(datapath_1_Instr_21_bF_buf37_), .B(datapath_1_RegisterFile_regfile_mem_10__1_), .C(datapath_1_Instr_22_bF_buf35_), .Y(_1947_) );
OAI22X1 OAI22X1_134 ( .A(_1947_), .B(_1946_), .C(datapath_1_Instr_22_bF_buf34_), .D(_1945_), .Y(_1948_) );
INVX1 INVX1_376 ( .A(datapath_1_RegisterFile_regfile_mem_15__1_), .Y(_1949_) );
AOI21X1 AOI21X1_587 ( .A(_1890__bF_buf12), .B(datapath_1_RegisterFile_regfile_mem_14__1_), .C(_1884__bF_buf8), .Y(_1950_) );
OAI21X1 OAI21X1_1652 ( .A(_1890__bF_buf12), .B(_1949_), .C(_1950_), .Y(_1951_) );
NAND2X1 NAND2X1_1072 ( .A(datapath_1_RegisterFile_regfile_mem_12__1_), .B(_1890__bF_buf12), .Y(_1952_) );
AOI21X1 AOI21X1_588 ( .A(datapath_1_Instr_21_bF_buf36_), .B(datapath_1_RegisterFile_regfile_mem_13__1_), .C(datapath_1_Instr_22_bF_buf33_), .Y(_1953_) );
AOI21X1 AOI21X1_589 ( .A(_1952_), .B(_1953_), .C(_1885__bF_buf0), .Y(_1954_) );
AOI22X1 AOI22X1_127 ( .A(_1951_), .B(_1954_), .C(_1885__bF_buf0), .D(_1948_), .Y(_1955_) );
NOR2X1 NOR2X1_328 ( .A(datapath_1_Instr_21_bF_buf35_), .B(datapath_1_RegisterFile_regfile_mem_0__1_), .Y(_1956_) );
OAI21X1 OAI21X1_1653 ( .A(datapath_1_RegisterFile_regfile_mem_1__1_), .B(_1890__bF_buf41), .C(_1884__bF_buf8), .Y(_1957_) );
NOR2X1 NOR2X1_329 ( .A(datapath_1_RegisterFile_regfile_mem_3__1_), .B(_1890__bF_buf38), .Y(_1958_) );
OAI21X1 OAI21X1_1654 ( .A(datapath_1_Instr_21_bF_buf34_), .B(datapath_1_RegisterFile_regfile_mem_2__1_), .C(datapath_1_Instr_22_bF_buf32_), .Y(_1959_) );
OAI22X1 OAI22X1_135 ( .A(_1958_), .B(_1959_), .C(_1956_), .D(_1957_), .Y(_1960_) );
NOR2X1 NOR2X1_330 ( .A(datapath_1_Instr_23_bF_buf1_), .B(_1960_), .Y(_1961_) );
MUX2X1 MUX2X1_135 ( .A(datapath_1_RegisterFile_regfile_mem_5__1_), .B(datapath_1_RegisterFile_regfile_mem_4__1_), .S(datapath_1_Instr_21_bF_buf33_), .Y(_1962_) );
NOR2X1 NOR2X1_331 ( .A(datapath_1_RegisterFile_regfile_mem_7__1_), .B(_1890__bF_buf38), .Y(_1963_) );
OAI21X1 OAI21X1_1655 ( .A(datapath_1_Instr_21_bF_buf32_), .B(datapath_1_RegisterFile_regfile_mem_6__1_), .C(datapath_1_Instr_22_bF_buf31_), .Y(_1964_) );
OAI22X1 OAI22X1_136 ( .A(_1964_), .B(_1963_), .C(datapath_1_Instr_22_bF_buf30_), .D(_1962_), .Y(_1965_) );
OAI21X1 OAI21X1_1656 ( .A(_1885__bF_buf4), .B(_1965_), .C(_1888__bF_buf6), .Y(_1966_) );
OAI22X1 OAI22X1_137 ( .A(_1888__bF_buf6), .B(_1955_), .C(_1961_), .D(_1966_), .Y(_1967_) );
NAND2X1 NAND2X1_1073 ( .A(_1917__bF_buf3), .B(_1967_), .Y(_1968_) );
INVX1 INVX1_377 ( .A(datapath_1_RegisterFile_regfile_mem_27__1_), .Y(_1969_) );
AOI21X1 AOI21X1_590 ( .A(datapath_1_Instr_23_bF_buf0_), .B(datapath_1_RegisterFile_regfile_mem_31__1_), .C(_1890__bF_buf11), .Y(_1970_) );
OAI21X1 OAI21X1_1657 ( .A(datapath_1_Instr_23_bF_buf15_bF_buf2_), .B(_1969_), .C(_1970_), .Y(_1971_) );
INVX1 INVX1_378 ( .A(datapath_1_RegisterFile_regfile_mem_26__1_), .Y(_1972_) );
AOI21X1 AOI21X1_591 ( .A(datapath_1_Instr_23_bF_buf14_bF_buf2_), .B(datapath_1_RegisterFile_regfile_mem_30__1_), .C(datapath_1_Instr_21_bF_buf31_), .Y(_1973_) );
OAI21X1 OAI21X1_1658 ( .A(datapath_1_Instr_23_bF_buf13_bF_buf2_), .B(_1972_), .C(_1973_), .Y(_1974_) );
NAND3X1 NAND3X1_1419 ( .A(datapath_1_Instr_22_bF_buf29_), .B(_1974_), .C(_1971_), .Y(_1975_) );
INVX1 INVX1_379 ( .A(datapath_1_RegisterFile_regfile_mem_25__1_), .Y(_1976_) );
AOI21X1 AOI21X1_592 ( .A(datapath_1_Instr_23_bF_buf12_bF_buf2_), .B(datapath_1_RegisterFile_regfile_mem_29__1_), .C(_1890__bF_buf11), .Y(_1977_) );
OAI21X1 OAI21X1_1659 ( .A(datapath_1_Instr_23_bF_buf11_bF_buf2_), .B(_1976_), .C(_1977_), .Y(_1978_) );
INVX1 INVX1_380 ( .A(datapath_1_RegisterFile_regfile_mem_24__1_), .Y(_1979_) );
AOI21X1 AOI21X1_593 ( .A(datapath_1_Instr_23_bF_buf10_bF_buf2_), .B(datapath_1_RegisterFile_regfile_mem_28__1_), .C(datapath_1_Instr_21_bF_buf30_), .Y(_1980_) );
OAI21X1 OAI21X1_1660 ( .A(datapath_1_Instr_23_bF_buf9_bF_buf2_), .B(_1979_), .C(_1980_), .Y(_1981_) );
NAND3X1 NAND3X1_1420 ( .A(_1884__bF_buf2), .B(_1981_), .C(_1978_), .Y(_1982_) );
AOI21X1 AOI21X1_594 ( .A(_1975_), .B(_1982_), .C(_1888__bF_buf0), .Y(_1983_) );
MUX2X1 MUX2X1_136 ( .A(datapath_1_RegisterFile_regfile_mem_18__1_), .B(datapath_1_RegisterFile_regfile_mem_16__1_), .S(datapath_1_Instr_22_bF_buf28_), .Y(_1984_) );
NAND2X1 NAND2X1_1074 ( .A(_1890__bF_buf43), .B(_1984_), .Y(_1985_) );
MUX2X1 MUX2X1_137 ( .A(datapath_1_RegisterFile_regfile_mem_19__1_), .B(datapath_1_RegisterFile_regfile_mem_17__1_), .S(datapath_1_Instr_22_bF_buf27_), .Y(_1986_) );
NAND2X1 NAND2X1_1075 ( .A(datapath_1_Instr_21_bF_buf29_), .B(_1986_), .Y(_1987_) );
NAND3X1 NAND3X1_1421 ( .A(_1885__bF_buf3), .B(_1985_), .C(_1987_), .Y(_1988_) );
MUX2X1 MUX2X1_138 ( .A(datapath_1_RegisterFile_regfile_mem_22__1_), .B(datapath_1_RegisterFile_regfile_mem_20__1_), .S(datapath_1_Instr_22_bF_buf26_), .Y(_1989_) );
NAND2X1 NAND2X1_1076 ( .A(_1890__bF_buf11), .B(_1989_), .Y(_1990_) );
MUX2X1 MUX2X1_139 ( .A(datapath_1_RegisterFile_regfile_mem_23__1_), .B(datapath_1_RegisterFile_regfile_mem_21__1_), .S(datapath_1_Instr_22_bF_buf25_), .Y(_1991_) );
NAND2X1 NAND2X1_1077 ( .A(datapath_1_Instr_21_bF_buf28_), .B(_1991_), .Y(_1992_) );
NAND3X1 NAND3X1_1422 ( .A(datapath_1_Instr_23_bF_buf8_bF_buf2_), .B(_1990_), .C(_1992_), .Y(_1993_) );
AOI21X1 AOI21X1_595 ( .A(_1988_), .B(_1993_), .C(datapath_1_Instr_24_bF_buf0_), .Y(_1994_) );
OAI21X1 OAI21X1_1661 ( .A(_1983_), .B(_1994_), .C(datapath_1_Instr_25_bF_buf0_), .Y(_1995_) );
AOI22X1 AOI22X1_128 ( .A(_1883__bF_buf0), .B(_1887__bF_buf2), .C(_1995_), .D(_1968_), .Y(datapath_1_RD1_1_) );
MUX2X1 MUX2X1_140 ( .A(datapath_1_RegisterFile_regfile_mem_2__2_), .B(datapath_1_RegisterFile_regfile_mem_0__2_), .S(datapath_1_Instr_22_bF_buf24_), .Y(_1996_) );
NAND2X1 NAND2X1_1078 ( .A(_1890__bF_buf12), .B(_1996_), .Y(_1997_) );
MUX2X1 MUX2X1_141 ( .A(datapath_1_RegisterFile_regfile_mem_3__2_), .B(datapath_1_RegisterFile_regfile_mem_1__2_), .S(datapath_1_Instr_22_bF_buf23_), .Y(_1998_) );
NAND2X1 NAND2X1_1079 ( .A(datapath_1_Instr_21_bF_buf27_), .B(_1998_), .Y(_1999_) );
NAND3X1 NAND3X1_1423 ( .A(_1885__bF_buf0), .B(_1997_), .C(_1999_), .Y(_2000_) );
MUX2X1 MUX2X1_142 ( .A(datapath_1_RegisterFile_regfile_mem_6__2_), .B(datapath_1_RegisterFile_regfile_mem_4__2_), .S(datapath_1_Instr_22_bF_buf22_), .Y(_2001_) );
NAND2X1 NAND2X1_1080 ( .A(_1890__bF_buf8), .B(_2001_), .Y(_2002_) );
MUX2X1 MUX2X1_143 ( .A(datapath_1_RegisterFile_regfile_mem_7__2_), .B(datapath_1_RegisterFile_regfile_mem_5__2_), .S(datapath_1_Instr_22_bF_buf21_), .Y(_2003_) );
NAND2X1 NAND2X1_1081 ( .A(datapath_1_Instr_21_bF_buf26_), .B(_2003_), .Y(_2004_) );
NAND3X1 NAND3X1_1424 ( .A(datapath_1_Instr_23_bF_buf7_bF_buf2_), .B(_2002_), .C(_2004_), .Y(_2005_) );
AOI21X1 AOI21X1_596 ( .A(_2000_), .B(_2005_), .C(datapath_1_Instr_24_bF_buf6_), .Y(_2006_) );
INVX1 INVX1_381 ( .A(datapath_1_RegisterFile_regfile_mem_9__2_), .Y(_2007_) );
AOI21X1 AOI21X1_597 ( .A(datapath_1_Instr_23_bF_buf6_bF_buf2_), .B(datapath_1_RegisterFile_regfile_mem_13__2_), .C(_1890__bF_buf41), .Y(_2008_) );
OAI21X1 OAI21X1_1662 ( .A(datapath_1_Instr_23_bF_buf5_bF_buf2_), .B(_2007_), .C(_2008_), .Y(_2009_) );
INVX1 INVX1_382 ( .A(datapath_1_RegisterFile_regfile_mem_8__2_), .Y(_2010_) );
AOI21X1 AOI21X1_598 ( .A(datapath_1_Instr_23_bF_buf4_bF_buf2_), .B(datapath_1_RegisterFile_regfile_mem_12__2_), .C(datapath_1_Instr_21_bF_buf25_), .Y(_2011_) );
OAI21X1 OAI21X1_1663 ( .A(datapath_1_Instr_23_bF_buf3_bF_buf2_), .B(_2010_), .C(_2011_), .Y(_2012_) );
NAND3X1 NAND3X1_1425 ( .A(_1884__bF_buf4), .B(_2012_), .C(_2009_), .Y(_2013_) );
INVX1 INVX1_383 ( .A(datapath_1_RegisterFile_regfile_mem_11__2_), .Y(_2014_) );
AOI21X1 AOI21X1_599 ( .A(datapath_1_Instr_23_bF_buf2_bF_buf2_), .B(datapath_1_RegisterFile_regfile_mem_15__2_), .C(_1890__bF_buf41), .Y(_2015_) );
OAI21X1 OAI21X1_1664 ( .A(datapath_1_Instr_23_bF_buf1_), .B(_2014_), .C(_2015_), .Y(_2016_) );
INVX1 INVX1_384 ( .A(datapath_1_RegisterFile_regfile_mem_10__2_), .Y(_2017_) );
AOI21X1 AOI21X1_600 ( .A(datapath_1_Instr_23_bF_buf0_), .B(datapath_1_RegisterFile_regfile_mem_14__2_), .C(datapath_1_Instr_21_bF_buf24_), .Y(_2018_) );
OAI21X1 OAI21X1_1665 ( .A(datapath_1_Instr_23_bF_buf15_bF_buf1_), .B(_2017_), .C(_2018_), .Y(_2019_) );
NAND3X1 NAND3X1_1426 ( .A(datapath_1_Instr_22_bF_buf20_), .B(_2019_), .C(_2016_), .Y(_2020_) );
AOI21X1 AOI21X1_601 ( .A(_2013_), .B(_2020_), .C(_1888__bF_buf6), .Y(_2021_) );
OAI21X1 OAI21X1_1666 ( .A(_2021_), .B(_2006_), .C(_1917__bF_buf2), .Y(_2022_) );
NOR2X1 NOR2X1_332 ( .A(datapath_1_Instr_21_bF_buf23_), .B(datapath_1_RegisterFile_regfile_mem_24__2_), .Y(_2023_) );
OAI21X1 OAI21X1_1667 ( .A(datapath_1_RegisterFile_regfile_mem_25__2_), .B(_1890__bF_buf35), .C(_1884__bF_buf6), .Y(_2024_) );
NOR2X1 NOR2X1_333 ( .A(datapath_1_RegisterFile_regfile_mem_27__2_), .B(_1890__bF_buf35), .Y(_2025_) );
OAI21X1 OAI21X1_1668 ( .A(datapath_1_Instr_21_bF_buf22_), .B(datapath_1_RegisterFile_regfile_mem_26__2_), .C(datapath_1_Instr_22_bF_buf19_), .Y(_2026_) );
OAI22X1 OAI22X1_138 ( .A(_2025_), .B(_2026_), .C(_2023_), .D(_2024_), .Y(_2027_) );
NOR2X1 NOR2X1_334 ( .A(datapath_1_Instr_23_bF_buf14_bF_buf1_), .B(_2027_), .Y(_2028_) );
MUX2X1 MUX2X1_144 ( .A(datapath_1_RegisterFile_regfile_mem_29__2_), .B(datapath_1_RegisterFile_regfile_mem_28__2_), .S(datapath_1_Instr_21_bF_buf21_), .Y(_2029_) );
NOR2X1 NOR2X1_335 ( .A(datapath_1_RegisterFile_regfile_mem_31__2_), .B(_1890__bF_buf32), .Y(_2030_) );
OAI21X1 OAI21X1_1669 ( .A(datapath_1_Instr_21_bF_buf20_), .B(datapath_1_RegisterFile_regfile_mem_30__2_), .C(datapath_1_Instr_22_bF_buf18_), .Y(_2031_) );
OAI22X1 OAI22X1_139 ( .A(_2031_), .B(_2030_), .C(datapath_1_Instr_22_bF_buf17_), .D(_2029_), .Y(_2032_) );
OAI21X1 OAI21X1_1670 ( .A(_1885__bF_buf10), .B(_2032_), .C(datapath_1_Instr_24_bF_buf5_), .Y(_2033_) );
INVX1 INVX1_385 ( .A(datapath_1_RegisterFile_regfile_mem_19__2_), .Y(_2034_) );
AOI21X1 AOI21X1_602 ( .A(datapath_1_Instr_23_bF_buf13_bF_buf1_), .B(datapath_1_RegisterFile_regfile_mem_23__2_), .C(_1890__bF_buf32), .Y(_2035_) );
OAI21X1 OAI21X1_1671 ( .A(datapath_1_Instr_23_bF_buf12_bF_buf1_), .B(_2034_), .C(_2035_), .Y(_2036_) );
NAND2X1 NAND2X1_1082 ( .A(datapath_1_RegisterFile_regfile_mem_18__2_), .B(_1885__bF_buf3), .Y(_2037_) );
AOI21X1 AOI21X1_603 ( .A(datapath_1_Instr_23_bF_buf11_bF_buf1_), .B(datapath_1_RegisterFile_regfile_mem_22__2_), .C(datapath_1_Instr_21_bF_buf19_), .Y(_2038_) );
AOI21X1 AOI21X1_604 ( .A(_2037_), .B(_2038_), .C(_1884__bF_buf6), .Y(_2039_) );
INVX1 INVX1_386 ( .A(datapath_1_RegisterFile_regfile_mem_17__2_), .Y(_2040_) );
AOI21X1 AOI21X1_605 ( .A(datapath_1_Instr_23_bF_buf10_bF_buf1_), .B(datapath_1_RegisterFile_regfile_mem_21__2_), .C(_1890__bF_buf32), .Y(_2041_) );
OAI21X1 OAI21X1_1672 ( .A(datapath_1_Instr_23_bF_buf9_bF_buf1_), .B(_2040_), .C(_2041_), .Y(_2042_) );
NAND2X1 NAND2X1_1083 ( .A(datapath_1_RegisterFile_regfile_mem_16__2_), .B(_1885__bF_buf3), .Y(_2043_) );
AOI21X1 AOI21X1_606 ( .A(datapath_1_Instr_23_bF_buf8_bF_buf1_), .B(datapath_1_RegisterFile_regfile_mem_20__2_), .C(datapath_1_Instr_21_bF_buf18_), .Y(_2044_) );
AOI21X1 AOI21X1_607 ( .A(_2043_), .B(_2044_), .C(datapath_1_Instr_22_bF_buf16_), .Y(_2045_) );
AOI22X1 AOI22X1_129 ( .A(_2039_), .B(_2036_), .C(_2042_), .D(_2045_), .Y(_2046_) );
OAI22X1 OAI22X1_140 ( .A(datapath_1_Instr_24_bF_buf4_), .B(_2046_), .C(_2028_), .D(_2033_), .Y(_2047_) );
NAND2X1 NAND2X1_1084 ( .A(datapath_1_Instr_25_bF_buf5_), .B(_2047_), .Y(_2048_) );
AOI22X1 AOI22X1_130 ( .A(_1883__bF_buf1), .B(_1887__bF_buf2), .C(_2022_), .D(_2048_), .Y(datapath_1_RD1_2_) );
NAND2X1 NAND2X1_1085 ( .A(datapath_1_Instr_21_bF_buf17_), .B(datapath_1_RegisterFile_regfile_mem_27__3_), .Y(_2049_) );
NAND2X1 NAND2X1_1086 ( .A(datapath_1_RegisterFile_regfile_mem_26__3_), .B(_1890__bF_buf17), .Y(_2050_) );
NAND3X1 NAND3X1_1427 ( .A(datapath_1_Instr_22_bF_buf15_), .B(_2049_), .C(_2050_), .Y(_2051_) );
NAND2X1 NAND2X1_1087 ( .A(datapath_1_Instr_21_bF_buf16_), .B(datapath_1_RegisterFile_regfile_mem_25__3_), .Y(_2052_) );
AOI21X1 AOI21X1_608 ( .A(_1890__bF_buf17), .B(datapath_1_RegisterFile_regfile_mem_24__3_), .C(datapath_1_Instr_22_bF_buf14_), .Y(_2053_) );
NAND2X1 NAND2X1_1088 ( .A(_2052_), .B(_2053_), .Y(_2054_) );
NAND3X1 NAND3X1_1428 ( .A(_1885__bF_buf10), .B(_2051_), .C(_2054_), .Y(_2055_) );
NAND2X1 NAND2X1_1089 ( .A(datapath_1_Instr_21_bF_buf15_), .B(datapath_1_RegisterFile_regfile_mem_31__3_), .Y(_2056_) );
AOI21X1 AOI21X1_609 ( .A(_1890__bF_buf19), .B(datapath_1_RegisterFile_regfile_mem_30__3_), .C(_1884__bF_buf6), .Y(_2057_) );
NAND2X1 NAND2X1_1090 ( .A(_2056_), .B(_2057_), .Y(_2058_) );
INVX1 INVX1_387 ( .A(datapath_1_RegisterFile_regfile_mem_28__3_), .Y(_2059_) );
AOI21X1 AOI21X1_610 ( .A(datapath_1_Instr_21_bF_buf14_), .B(datapath_1_RegisterFile_regfile_mem_29__3_), .C(datapath_1_Instr_22_bF_buf13_), .Y(_2060_) );
OAI21X1 OAI21X1_1673 ( .A(datapath_1_Instr_21_bF_buf13_), .B(_2059_), .C(_2060_), .Y(_2061_) );
NAND3X1 NAND3X1_1429 ( .A(datapath_1_Instr_23_bF_buf7_bF_buf1_), .B(_2061_), .C(_2058_), .Y(_2062_) );
AOI21X1 AOI21X1_611 ( .A(_2055_), .B(_2062_), .C(_1888__bF_buf3), .Y(_2063_) );
MUX2X1 MUX2X1_145 ( .A(datapath_1_RegisterFile_regfile_mem_17__3_), .B(datapath_1_RegisterFile_regfile_mem_16__3_), .S(datapath_1_Instr_21_bF_buf12_), .Y(_2064_) );
NOR2X1 NOR2X1_336 ( .A(datapath_1_RegisterFile_regfile_mem_19__3_), .B(_1890__bF_buf19), .Y(_2065_) );
OAI21X1 OAI21X1_1674 ( .A(datapath_1_Instr_21_bF_buf11_), .B(datapath_1_RegisterFile_regfile_mem_18__3_), .C(datapath_1_Instr_22_bF_buf12_), .Y(_2066_) );
OAI22X1 OAI22X1_141 ( .A(_2066_), .B(_2065_), .C(datapath_1_Instr_22_bF_buf11_), .D(_2064_), .Y(_2067_) );
NAND2X1 NAND2X1_1091 ( .A(_1885__bF_buf10), .B(_2067_), .Y(_2068_) );
MUX2X1 MUX2X1_146 ( .A(datapath_1_RegisterFile_regfile_mem_21__3_), .B(datapath_1_RegisterFile_regfile_mem_20__3_), .S(datapath_1_Instr_21_bF_buf10_), .Y(_2069_) );
NOR2X1 NOR2X1_337 ( .A(datapath_1_RegisterFile_regfile_mem_23__3_), .B(_1890__bF_buf19), .Y(_2070_) );
OAI21X1 OAI21X1_1675 ( .A(datapath_1_Instr_21_bF_buf9_), .B(datapath_1_RegisterFile_regfile_mem_22__3_), .C(datapath_1_Instr_22_bF_buf10_), .Y(_2071_) );
OAI22X1 OAI22X1_142 ( .A(_2071_), .B(_2070_), .C(datapath_1_Instr_22_bF_buf9_), .D(_2069_), .Y(_2072_) );
NAND2X1 NAND2X1_1092 ( .A(datapath_1_Instr_23_bF_buf6_bF_buf1_), .B(_2072_), .Y(_2073_) );
AOI21X1 AOI21X1_612 ( .A(_2068_), .B(_2073_), .C(datapath_1_Instr_24_bF_buf3_), .Y(_2074_) );
OAI21X1 OAI21X1_1676 ( .A(_2063_), .B(_2074_), .C(datapath_1_Instr_25_bF_buf4_), .Y(_2075_) );
NAND2X1 NAND2X1_1093 ( .A(datapath_1_Instr_22_bF_buf8_), .B(datapath_1_RegisterFile_regfile_mem_11__3_), .Y(_2076_) );
NAND2X1 NAND2X1_1094 ( .A(datapath_1_RegisterFile_regfile_mem_9__3_), .B(_1884__bF_buf8), .Y(_2077_) );
NAND3X1 NAND3X1_1430 ( .A(datapath_1_Instr_21_bF_buf8_), .B(_2076_), .C(_2077_), .Y(_2078_) );
NAND2X1 NAND2X1_1095 ( .A(datapath_1_Instr_22_bF_buf7_), .B(datapath_1_RegisterFile_regfile_mem_10__3_), .Y(_2079_) );
AOI21X1 AOI21X1_613 ( .A(_1884__bF_buf8), .B(datapath_1_RegisterFile_regfile_mem_8__3_), .C(datapath_1_Instr_21_bF_buf7_), .Y(_2080_) );
NAND2X1 NAND2X1_1096 ( .A(_2079_), .B(_2080_), .Y(_2081_) );
NAND3X1 NAND3X1_1431 ( .A(_1885__bF_buf0), .B(_2078_), .C(_2081_), .Y(_2082_) );
NAND2X1 NAND2X1_1097 ( .A(datapath_1_Instr_22_bF_buf6_), .B(datapath_1_RegisterFile_regfile_mem_15__3_), .Y(_2083_) );
NAND2X1 NAND2X1_1098 ( .A(datapath_1_RegisterFile_regfile_mem_13__3_), .B(_1884__bF_buf8), .Y(_2084_) );
NAND3X1 NAND3X1_1432 ( .A(datapath_1_Instr_21_bF_buf6_), .B(_2083_), .C(_2084_), .Y(_2085_) );
NAND2X1 NAND2X1_1099 ( .A(datapath_1_Instr_22_bF_buf5_), .B(datapath_1_RegisterFile_regfile_mem_14__3_), .Y(_2086_) );
AOI21X1 AOI21X1_614 ( .A(_1884__bF_buf8), .B(datapath_1_RegisterFile_regfile_mem_12__3_), .C(datapath_1_Instr_21_bF_buf5_), .Y(_2087_) );
NAND2X1 NAND2X1_1100 ( .A(_2086_), .B(_2087_), .Y(_2088_) );
NAND3X1 NAND3X1_1433 ( .A(datapath_1_Instr_23_bF_buf5_bF_buf1_), .B(_2085_), .C(_2088_), .Y(_2089_) );
AOI21X1 AOI21X1_615 ( .A(_2082_), .B(_2089_), .C(_1888__bF_buf7), .Y(_2090_) );
INVX1 INVX1_388 ( .A(datapath_1_RegisterFile_regfile_mem_1__3_), .Y(_2091_) );
AOI21X1 AOI21X1_616 ( .A(datapath_1_Instr_23_bF_buf4_bF_buf1_), .B(datapath_1_RegisterFile_regfile_mem_5__3_), .C(_1890__bF_buf8), .Y(_2092_) );
OAI21X1 OAI21X1_1677 ( .A(datapath_1_Instr_23_bF_buf3_bF_buf1_), .B(_2091_), .C(_2092_), .Y(_2093_) );
INVX1 INVX1_389 ( .A(datapath_1_RegisterFile_regfile_mem_0__3_), .Y(_2094_) );
AOI21X1 AOI21X1_617 ( .A(datapath_1_Instr_23_bF_buf2_bF_buf1_), .B(datapath_1_RegisterFile_regfile_mem_4__3_), .C(datapath_1_Instr_21_bF_buf4_), .Y(_2095_) );
OAI21X1 OAI21X1_1678 ( .A(datapath_1_Instr_23_bF_buf1_), .B(_2094_), .C(_2095_), .Y(_2096_) );
NAND3X1 NAND3X1_1434 ( .A(_1884__bF_buf8), .B(_2096_), .C(_2093_), .Y(_2097_) );
INVX1 INVX1_390 ( .A(datapath_1_RegisterFile_regfile_mem_3__3_), .Y(_2098_) );
AOI21X1 AOI21X1_618 ( .A(datapath_1_Instr_23_bF_buf0_), .B(datapath_1_RegisterFile_regfile_mem_7__3_), .C(_1890__bF_buf8), .Y(_2099_) );
OAI21X1 OAI21X1_1679 ( .A(datapath_1_Instr_23_bF_buf15_bF_buf0_), .B(_2098_), .C(_2099_), .Y(_2100_) );
INVX1 INVX1_391 ( .A(datapath_1_RegisterFile_regfile_mem_2__3_), .Y(_2101_) );
AOI21X1 AOI21X1_619 ( .A(datapath_1_Instr_23_bF_buf14_bF_buf0_), .B(datapath_1_RegisterFile_regfile_mem_6__3_), .C(datapath_1_Instr_21_bF_buf3_), .Y(_2102_) );
OAI21X1 OAI21X1_1680 ( .A(datapath_1_Instr_23_bF_buf13_bF_buf0_), .B(_2101_), .C(_2102_), .Y(_2103_) );
NAND3X1 NAND3X1_1435 ( .A(datapath_1_Instr_22_bF_buf4_), .B(_2103_), .C(_2100_), .Y(_2104_) );
AOI21X1 AOI21X1_620 ( .A(_2097_), .B(_2104_), .C(datapath_1_Instr_24_bF_buf2_), .Y(_2105_) );
OAI21X1 OAI21X1_1681 ( .A(_2105_), .B(_2090_), .C(_1917__bF_buf2), .Y(_2106_) );
AOI22X1 AOI22X1_131 ( .A(_1883__bF_buf1), .B(_1887__bF_buf0), .C(_2106_), .D(_2075_), .Y(datapath_1_RD1_3_) );
MUX2X1 MUX2X1_147 ( .A(datapath_1_RegisterFile_regfile_mem_9__4_), .B(datapath_1_RegisterFile_regfile_mem_8__4_), .S(datapath_1_Instr_21_bF_buf2_), .Y(_2107_) );
NOR2X1 NOR2X1_338 ( .A(datapath_1_RegisterFile_regfile_mem_11__4_), .B(_1890__bF_buf28), .Y(_2108_) );
OAI21X1 OAI21X1_1682 ( .A(datapath_1_Instr_21_bF_buf1_), .B(datapath_1_RegisterFile_regfile_mem_10__4_), .C(datapath_1_Instr_22_bF_buf3_), .Y(_2109_) );
OAI22X1 OAI22X1_143 ( .A(_2109_), .B(_2108_), .C(datapath_1_Instr_22_bF_buf2_), .D(_2107_), .Y(_2110_) );
INVX1 INVX1_392 ( .A(datapath_1_RegisterFile_regfile_mem_15__4_), .Y(_2111_) );
AOI21X1 AOI21X1_621 ( .A(_1890__bF_buf28), .B(datapath_1_RegisterFile_regfile_mem_14__4_), .C(_1884__bF_buf4), .Y(_2112_) );
OAI21X1 OAI21X1_1683 ( .A(_1890__bF_buf28), .B(_2111_), .C(_2112_), .Y(_2113_) );
NAND2X1 NAND2X1_1101 ( .A(datapath_1_RegisterFile_regfile_mem_12__4_), .B(_1890__bF_buf28), .Y(_2114_) );
AOI21X1 AOI21X1_622 ( .A(datapath_1_Instr_21_bF_buf0_), .B(datapath_1_RegisterFile_regfile_mem_13__4_), .C(datapath_1_Instr_22_bF_buf1_), .Y(_2115_) );
AOI21X1 AOI21X1_623 ( .A(_2114_), .B(_2115_), .C(_1885__bF_buf4), .Y(_2116_) );
AOI22X1 AOI22X1_132 ( .A(_2113_), .B(_2116_), .C(_1885__bF_buf4), .D(_2110_), .Y(_2117_) );
NOR2X1 NOR2X1_339 ( .A(datapath_1_Instr_21_bF_buf55_), .B(datapath_1_RegisterFile_regfile_mem_0__4_), .Y(_2118_) );
OAI21X1 OAI21X1_1684 ( .A(datapath_1_RegisterFile_regfile_mem_1__4_), .B(_1890__bF_buf27), .C(_1884__bF_buf4), .Y(_2119_) );
NOR2X1 NOR2X1_340 ( .A(datapath_1_RegisterFile_regfile_mem_3__4_), .B(_1890__bF_buf27), .Y(_2120_) );
OAI21X1 OAI21X1_1685 ( .A(datapath_1_Instr_21_bF_buf54_), .B(datapath_1_RegisterFile_regfile_mem_2__4_), .C(datapath_1_Instr_22_bF_buf0_), .Y(_2121_) );
OAI22X1 OAI22X1_144 ( .A(_2120_), .B(_2121_), .C(_2118_), .D(_2119_), .Y(_2122_) );
NOR2X1 NOR2X1_341 ( .A(datapath_1_Instr_23_bF_buf12_bF_buf0_), .B(_2122_), .Y(_2123_) );
MUX2X1 MUX2X1_148 ( .A(datapath_1_RegisterFile_regfile_mem_5__4_), .B(datapath_1_RegisterFile_regfile_mem_4__4_), .S(datapath_1_Instr_21_bF_buf53_), .Y(_2124_) );
NOR2X1 NOR2X1_342 ( .A(datapath_1_RegisterFile_regfile_mem_7__4_), .B(_1890__bF_buf27), .Y(_2125_) );
OAI21X1 OAI21X1_1686 ( .A(datapath_1_Instr_21_bF_buf52_), .B(datapath_1_RegisterFile_regfile_mem_6__4_), .C(datapath_1_Instr_22_bF_buf50_), .Y(_2126_) );
OAI22X1 OAI22X1_145 ( .A(_2126_), .B(_2125_), .C(datapath_1_Instr_22_bF_buf49_), .D(_2124_), .Y(_2127_) );
OAI21X1 OAI21X1_1687 ( .A(_1885__bF_buf4), .B(_2127_), .C(_1888__bF_buf6), .Y(_2128_) );
OAI22X1 OAI22X1_146 ( .A(_1888__bF_buf6), .B(_2117_), .C(_2123_), .D(_2128_), .Y(_2129_) );
NAND2X1 NAND2X1_1102 ( .A(_1917__bF_buf3), .B(_2129_), .Y(_2130_) );
INVX1 INVX1_393 ( .A(datapath_1_RegisterFile_regfile_mem_27__4_), .Y(_2131_) );
AOI21X1 AOI21X1_624 ( .A(datapath_1_Instr_23_bF_buf11_bF_buf0_), .B(datapath_1_RegisterFile_regfile_mem_31__4_), .C(_1890__bF_buf25), .Y(_2132_) );
OAI21X1 OAI21X1_1688 ( .A(datapath_1_Instr_23_bF_buf10_bF_buf0_), .B(_2131_), .C(_2132_), .Y(_2133_) );
INVX1 INVX1_394 ( .A(datapath_1_RegisterFile_regfile_mem_26__4_), .Y(_2134_) );
AOI21X1 AOI21X1_625 ( .A(datapath_1_Instr_23_bF_buf9_bF_buf0_), .B(datapath_1_RegisterFile_regfile_mem_30__4_), .C(datapath_1_Instr_21_bF_buf51_), .Y(_2135_) );
OAI21X1 OAI21X1_1689 ( .A(datapath_1_Instr_23_bF_buf8_bF_buf0_), .B(_2134_), .C(_2135_), .Y(_2136_) );
NAND3X1 NAND3X1_1436 ( .A(datapath_1_Instr_22_bF_buf48_), .B(_2136_), .C(_2133_), .Y(_2137_) );
INVX1 INVX1_395 ( .A(datapath_1_RegisterFile_regfile_mem_25__4_), .Y(_2138_) );
AOI21X1 AOI21X1_626 ( .A(datapath_1_Instr_23_bF_buf7_bF_buf0_), .B(datapath_1_RegisterFile_regfile_mem_29__4_), .C(_1890__bF_buf25), .Y(_2139_) );
OAI21X1 OAI21X1_1690 ( .A(datapath_1_Instr_23_bF_buf6_bF_buf0_), .B(_2138_), .C(_2139_), .Y(_2140_) );
INVX1 INVX1_396 ( .A(datapath_1_RegisterFile_regfile_mem_24__4_), .Y(_2141_) );
AOI21X1 AOI21X1_627 ( .A(datapath_1_Instr_23_bF_buf5_bF_buf0_), .B(datapath_1_RegisterFile_regfile_mem_28__4_), .C(datapath_1_Instr_21_bF_buf50_), .Y(_2142_) );
OAI21X1 OAI21X1_1691 ( .A(datapath_1_Instr_23_bF_buf4_bF_buf0_), .B(_2141_), .C(_2142_), .Y(_2143_) );
NAND3X1 NAND3X1_1437 ( .A(_1884__bF_buf2), .B(_2143_), .C(_2140_), .Y(_2144_) );
AOI21X1 AOI21X1_628 ( .A(_2137_), .B(_2144_), .C(_1888__bF_buf0), .Y(_2145_) );
MUX2X1 MUX2X1_149 ( .A(datapath_1_RegisterFile_regfile_mem_18__4_), .B(datapath_1_RegisterFile_regfile_mem_16__4_), .S(datapath_1_Instr_22_bF_buf47_), .Y(_2146_) );
NAND2X1 NAND2X1_1103 ( .A(_1890__bF_buf40), .B(_2146_), .Y(_2147_) );
MUX2X1 MUX2X1_150 ( .A(datapath_1_RegisterFile_regfile_mem_19__4_), .B(datapath_1_RegisterFile_regfile_mem_17__4_), .S(datapath_1_Instr_22_bF_buf46_), .Y(_2148_) );
NAND2X1 NAND2X1_1104 ( .A(datapath_1_Instr_21_bF_buf49_), .B(_2148_), .Y(_2149_) );
NAND3X1 NAND3X1_1438 ( .A(_1885__bF_buf11), .B(_2147_), .C(_2149_), .Y(_2150_) );
MUX2X1 MUX2X1_151 ( .A(datapath_1_RegisterFile_regfile_mem_22__4_), .B(datapath_1_RegisterFile_regfile_mem_20__4_), .S(datapath_1_Instr_22_bF_buf45_), .Y(_2151_) );
NAND2X1 NAND2X1_1105 ( .A(_1890__bF_buf40), .B(_2151_), .Y(_2152_) );
MUX2X1 MUX2X1_152 ( .A(datapath_1_RegisterFile_regfile_mem_23__4_), .B(datapath_1_RegisterFile_regfile_mem_21__4_), .S(datapath_1_Instr_22_bF_buf44_), .Y(_2153_) );
NAND2X1 NAND2X1_1106 ( .A(datapath_1_Instr_21_bF_buf48_), .B(_2153_), .Y(_2154_) );
NAND3X1 NAND3X1_1439 ( .A(datapath_1_Instr_23_bF_buf3_bF_buf0_), .B(_2152_), .C(_2154_), .Y(_2155_) );
AOI21X1 AOI21X1_629 ( .A(_2150_), .B(_2155_), .C(datapath_1_Instr_24_bF_buf1_), .Y(_2156_) );
OAI21X1 OAI21X1_1692 ( .A(_2145_), .B(_2156_), .C(datapath_1_Instr_25_bF_buf3_), .Y(_2157_) );
AOI22X1 AOI22X1_133 ( .A(_1883__bF_buf2), .B(_1887__bF_buf4), .C(_2157_), .D(_2130_), .Y(datapath_1_RD1_4_) );
MUX2X1 MUX2X1_153 ( .A(datapath_1_RegisterFile_regfile_mem_9__5_), .B(datapath_1_RegisterFile_regfile_mem_8__5_), .S(datapath_1_Instr_21_bF_buf47_), .Y(_2158_) );
NOR2X1 NOR2X1_343 ( .A(datapath_1_RegisterFile_regfile_mem_11__5_), .B(_1890__bF_buf15), .Y(_2159_) );
OAI21X1 OAI21X1_1693 ( .A(datapath_1_Instr_21_bF_buf46_), .B(datapath_1_RegisterFile_regfile_mem_10__5_), .C(datapath_1_Instr_22_bF_buf43_), .Y(_2160_) );
OAI22X1 OAI22X1_147 ( .A(_2160_), .B(_2159_), .C(datapath_1_Instr_22_bF_buf42_), .D(_2158_), .Y(_2161_) );
INVX1 INVX1_397 ( .A(datapath_1_RegisterFile_regfile_mem_15__5_), .Y(_2162_) );
AOI21X1 AOI21X1_630 ( .A(_1890__bF_buf15), .B(datapath_1_RegisterFile_regfile_mem_14__5_), .C(_1884__bF_buf5), .Y(_2163_) );
OAI21X1 OAI21X1_1694 ( .A(_1890__bF_buf15), .B(_2162_), .C(_2163_), .Y(_2164_) );
NAND2X1 NAND2X1_1107 ( .A(datapath_1_RegisterFile_regfile_mem_12__5_), .B(_1890__bF_buf15), .Y(_2165_) );
AOI21X1 AOI21X1_631 ( .A(datapath_1_Instr_21_bF_buf45_), .B(datapath_1_RegisterFile_regfile_mem_13__5_), .C(datapath_1_Instr_22_bF_buf41_), .Y(_2166_) );
AOI21X1 AOI21X1_632 ( .A(_2165_), .B(_2166_), .C(_1885__bF_buf1), .Y(_2167_) );
AOI22X1 AOI22X1_134 ( .A(_2164_), .B(_2167_), .C(_1885__bF_buf1), .D(_2161_), .Y(_2168_) );
NOR2X1 NOR2X1_344 ( .A(datapath_1_Instr_21_bF_buf44_), .B(datapath_1_RegisterFile_regfile_mem_0__5_), .Y(_2169_) );
OAI21X1 OAI21X1_1695 ( .A(datapath_1_RegisterFile_regfile_mem_1__5_), .B(_1890__bF_buf30), .C(_1884__bF_buf3), .Y(_2170_) );
NOR2X1 NOR2X1_345 ( .A(datapath_1_RegisterFile_regfile_mem_3__5_), .B(_1890__bF_buf33), .Y(_2171_) );
OAI21X1 OAI21X1_1696 ( .A(datapath_1_Instr_21_bF_buf43_), .B(datapath_1_RegisterFile_regfile_mem_2__5_), .C(datapath_1_Instr_22_bF_buf40_), .Y(_2172_) );
OAI22X1 OAI22X1_148 ( .A(_2171_), .B(_2172_), .C(_2169_), .D(_2170_), .Y(_2173_) );
NOR2X1 NOR2X1_346 ( .A(datapath_1_Instr_23_bF_buf2_bF_buf0_), .B(_2173_), .Y(_2174_) );
MUX2X1 MUX2X1_154 ( .A(datapath_1_RegisterFile_regfile_mem_5__5_), .B(datapath_1_RegisterFile_regfile_mem_4__5_), .S(datapath_1_Instr_21_bF_buf42_), .Y(_2175_) );
NOR2X1 NOR2X1_347 ( .A(datapath_1_RegisterFile_regfile_mem_7__5_), .B(_1890__bF_buf13), .Y(_2176_) );
OAI21X1 OAI21X1_1697 ( .A(datapath_1_Instr_21_bF_buf41_), .B(datapath_1_RegisterFile_regfile_mem_6__5_), .C(datapath_1_Instr_22_bF_buf39_), .Y(_2177_) );
OAI22X1 OAI22X1_149 ( .A(_2177_), .B(_2176_), .C(datapath_1_Instr_22_bF_buf38_), .D(_2175_), .Y(_2178_) );
OAI21X1 OAI21X1_1698 ( .A(_1885__bF_buf1), .B(_2178_), .C(_1888__bF_buf2), .Y(_2179_) );
OAI22X1 OAI22X1_150 ( .A(_1888__bF_buf2), .B(_2168_), .C(_2174_), .D(_2179_), .Y(_2180_) );
NAND2X1 NAND2X1_1108 ( .A(_1917__bF_buf4), .B(_2180_), .Y(_2181_) );
INVX1 INVX1_398 ( .A(datapath_1_RegisterFile_regfile_mem_19__5_), .Y(_2182_) );
AOI21X1 AOI21X1_633 ( .A(datapath_1_Instr_23_bF_buf1_), .B(datapath_1_RegisterFile_regfile_mem_23__5_), .C(_1890__bF_buf24), .Y(_2183_) );
OAI21X1 OAI21X1_1699 ( .A(datapath_1_Instr_23_bF_buf0_), .B(_2182_), .C(_2183_), .Y(_2184_) );
NAND2X1 NAND2X1_1109 ( .A(datapath_1_RegisterFile_regfile_mem_18__5_), .B(_1885__bF_buf9), .Y(_2185_) );
AOI21X1 AOI21X1_634 ( .A(datapath_1_Instr_23_bF_buf15_bF_buf3_), .B(datapath_1_RegisterFile_regfile_mem_22__5_), .C(datapath_1_Instr_21_bF_buf40_), .Y(_2186_) );
AOI21X1 AOI21X1_635 ( .A(_2185_), .B(_2186_), .C(_1884__bF_buf3), .Y(_2187_) );
INVX1 INVX1_399 ( .A(datapath_1_RegisterFile_regfile_mem_17__5_), .Y(_2188_) );
AOI21X1 AOI21X1_636 ( .A(datapath_1_Instr_23_bF_buf14_bF_buf3_), .B(datapath_1_RegisterFile_regfile_mem_21__5_), .C(_1890__bF_buf24), .Y(_2189_) );
OAI21X1 OAI21X1_1700 ( .A(datapath_1_Instr_23_bF_buf13_bF_buf3_), .B(_2188_), .C(_2189_), .Y(_2190_) );
NAND2X1 NAND2X1_1110 ( .A(datapath_1_RegisterFile_regfile_mem_16__5_), .B(_1885__bF_buf6), .Y(_2191_) );
AOI21X1 AOI21X1_637 ( .A(datapath_1_Instr_23_bF_buf12_bF_buf3_), .B(datapath_1_RegisterFile_regfile_mem_20__5_), .C(datapath_1_Instr_21_bF_buf39_), .Y(_2192_) );
AOI21X1 AOI21X1_638 ( .A(_2191_), .B(_2192_), .C(datapath_1_Instr_22_bF_buf37_), .Y(_2193_) );
AOI22X1 AOI22X1_135 ( .A(_2187_), .B(_2184_), .C(_2190_), .D(_2193_), .Y(_2194_) );
NOR2X1 NOR2X1_348 ( .A(datapath_1_Instr_21_bF_buf38_), .B(datapath_1_RegisterFile_regfile_mem_24__5_), .Y(_2195_) );
OAI21X1 OAI21X1_1701 ( .A(datapath_1_RegisterFile_regfile_mem_25__5_), .B(_1890__bF_buf22), .C(_1884__bF_buf3), .Y(_2196_) );
NOR2X1 NOR2X1_349 ( .A(datapath_1_RegisterFile_regfile_mem_27__5_), .B(_1890__bF_buf22), .Y(_2197_) );
OAI21X1 OAI21X1_1702 ( .A(datapath_1_Instr_21_bF_buf37_), .B(datapath_1_RegisterFile_regfile_mem_26__5_), .C(datapath_1_Instr_22_bF_buf36_), .Y(_2198_) );
OAI22X1 OAI22X1_151 ( .A(_2197_), .B(_2198_), .C(_2195_), .D(_2196_), .Y(_2199_) );
NOR2X1 NOR2X1_350 ( .A(datapath_1_Instr_23_bF_buf11_bF_buf3_), .B(_2199_), .Y(_2200_) );
MUX2X1 MUX2X1_155 ( .A(datapath_1_RegisterFile_regfile_mem_29__5_), .B(datapath_1_RegisterFile_regfile_mem_28__5_), .S(datapath_1_Instr_21_bF_buf36_), .Y(_2201_) );
NOR2X1 NOR2X1_351 ( .A(datapath_1_RegisterFile_regfile_mem_31__5_), .B(_1890__bF_buf4), .Y(_2202_) );
OAI21X1 OAI21X1_1703 ( .A(datapath_1_Instr_21_bF_buf35_), .B(datapath_1_RegisterFile_regfile_mem_30__5_), .C(datapath_1_Instr_22_bF_buf35_), .Y(_2203_) );
OAI22X1 OAI22X1_152 ( .A(_2203_), .B(_2202_), .C(datapath_1_Instr_22_bF_buf34_), .D(_2201_), .Y(_2204_) );
OAI21X1 OAI21X1_1704 ( .A(_1885__bF_buf6), .B(_2204_), .C(datapath_1_Instr_24_bF_buf0_), .Y(_2205_) );
OAI22X1 OAI22X1_153 ( .A(datapath_1_Instr_24_bF_buf6_), .B(_2194_), .C(_2200_), .D(_2205_), .Y(_2206_) );
NAND2X1 NAND2X1_1111 ( .A(datapath_1_Instr_25_bF_buf2_), .B(_2206_), .Y(_2207_) );
AOI22X1 AOI22X1_136 ( .A(_1883__bF_buf4), .B(_1887__bF_buf3), .C(_2207_), .D(_2181_), .Y(datapath_1_RD1_5_) );
NAND2X1 NAND2X1_1112 ( .A(datapath_1_Instr_21_bF_buf34_), .B(datapath_1_RegisterFile_regfile_mem_27__6_), .Y(_2208_) );
NAND2X1 NAND2X1_1113 ( .A(datapath_1_RegisterFile_regfile_mem_26__6_), .B(_1890__bF_buf10), .Y(_2209_) );
NAND3X1 NAND3X1_1440 ( .A(datapath_1_Instr_22_bF_buf33_), .B(_2208_), .C(_2209_), .Y(_2210_) );
NAND2X1 NAND2X1_1114 ( .A(datapath_1_Instr_21_bF_buf33_), .B(datapath_1_RegisterFile_regfile_mem_25__6_), .Y(_2211_) );
AOI21X1 AOI21X1_639 ( .A(_1890__bF_buf7), .B(datapath_1_RegisterFile_regfile_mem_24__6_), .C(datapath_1_Instr_22_bF_buf32_), .Y(_2212_) );
NAND2X1 NAND2X1_1115 ( .A(_2211_), .B(_2212_), .Y(_2213_) );
NAND3X1 NAND3X1_1441 ( .A(_1885__bF_buf11), .B(_2210_), .C(_2213_), .Y(_2214_) );
NAND2X1 NAND2X1_1116 ( .A(datapath_1_Instr_21_bF_buf32_), .B(datapath_1_RegisterFile_regfile_mem_31__6_), .Y(_2215_) );
AOI21X1 AOI21X1_640 ( .A(_1890__bF_buf10), .B(datapath_1_RegisterFile_regfile_mem_30__6_), .C(_1884__bF_buf2), .Y(_2216_) );
NAND2X1 NAND2X1_1117 ( .A(_2215_), .B(_2216_), .Y(_2217_) );
INVX1 INVX1_400 ( .A(datapath_1_RegisterFile_regfile_mem_28__6_), .Y(_2218_) );
AOI21X1 AOI21X1_641 ( .A(datapath_1_Instr_21_bF_buf31_), .B(datapath_1_RegisterFile_regfile_mem_29__6_), .C(datapath_1_Instr_22_bF_buf31_), .Y(_2219_) );
OAI21X1 OAI21X1_1705 ( .A(datapath_1_Instr_21_bF_buf30_), .B(_2218_), .C(_2219_), .Y(_2220_) );
NAND3X1 NAND3X1_1442 ( .A(datapath_1_Instr_23_bF_buf10_bF_buf3_), .B(_2220_), .C(_2217_), .Y(_2221_) );
AOI21X1 AOI21X1_642 ( .A(_2214_), .B(_2221_), .C(_1888__bF_buf0), .Y(_2222_) );
MUX2X1 MUX2X1_156 ( .A(datapath_1_RegisterFile_regfile_mem_17__6_), .B(datapath_1_RegisterFile_regfile_mem_16__6_), .S(datapath_1_Instr_21_bF_buf29_), .Y(_2223_) );
NOR2X1 NOR2X1_352 ( .A(datapath_1_RegisterFile_regfile_mem_19__6_), .B(_1890__bF_buf25), .Y(_2224_) );
OAI21X1 OAI21X1_1706 ( .A(datapath_1_Instr_21_bF_buf28_), .B(datapath_1_RegisterFile_regfile_mem_18__6_), .C(datapath_1_Instr_22_bF_buf30_), .Y(_2225_) );
OAI22X1 OAI22X1_154 ( .A(_2225_), .B(_2224_), .C(datapath_1_Instr_22_bF_buf29_), .D(_2223_), .Y(_2226_) );
NAND2X1 NAND2X1_1118 ( .A(_1885__bF_buf7), .B(_2226_), .Y(_2227_) );
MUX2X1 MUX2X1_157 ( .A(datapath_1_RegisterFile_regfile_mem_21__6_), .B(datapath_1_RegisterFile_regfile_mem_20__6_), .S(datapath_1_Instr_21_bF_buf27_), .Y(_2228_) );
NOR2X1 NOR2X1_353 ( .A(datapath_1_RegisterFile_regfile_mem_23__6_), .B(_1890__bF_buf25), .Y(_2229_) );
OAI21X1 OAI21X1_1707 ( .A(datapath_1_Instr_21_bF_buf26_), .B(datapath_1_RegisterFile_regfile_mem_22__6_), .C(datapath_1_Instr_22_bF_buf28_), .Y(_2230_) );
OAI22X1 OAI22X1_155 ( .A(_2230_), .B(_2229_), .C(datapath_1_Instr_22_bF_buf27_), .D(_2228_), .Y(_2231_) );
NAND2X1 NAND2X1_1119 ( .A(datapath_1_Instr_23_bF_buf9_bF_buf3_), .B(_2231_), .Y(_2232_) );
AOI21X1 AOI21X1_643 ( .A(_2227_), .B(_2232_), .C(datapath_1_Instr_24_bF_buf5_), .Y(_2233_) );
OAI21X1 OAI21X1_1708 ( .A(_2222_), .B(_2233_), .C(datapath_1_Instr_25_bF_buf1_), .Y(_2234_) );
NAND2X1 NAND2X1_1120 ( .A(datapath_1_Instr_22_bF_buf26_), .B(datapath_1_RegisterFile_regfile_mem_11__6_), .Y(_2235_) );
NAND2X1 NAND2X1_1121 ( .A(datapath_1_RegisterFile_regfile_mem_9__6_), .B(_1884__bF_buf1), .Y(_2236_) );
NAND3X1 NAND3X1_1443 ( .A(datapath_1_Instr_21_bF_buf25_), .B(_2235_), .C(_2236_), .Y(_2237_) );
NAND2X1 NAND2X1_1122 ( .A(datapath_1_Instr_22_bF_buf25_), .B(datapath_1_RegisterFile_regfile_mem_10__6_), .Y(_2238_) );
AOI21X1 AOI21X1_644 ( .A(_1884__bF_buf1), .B(datapath_1_RegisterFile_regfile_mem_8__6_), .C(datapath_1_Instr_21_bF_buf24_), .Y(_2239_) );
NAND2X1 NAND2X1_1123 ( .A(_2238_), .B(_2239_), .Y(_2240_) );
NAND3X1 NAND3X1_1444 ( .A(_1885__bF_buf0), .B(_2237_), .C(_2240_), .Y(_2241_) );
NAND2X1 NAND2X1_1124 ( .A(datapath_1_Instr_22_bF_buf24_), .B(datapath_1_RegisterFile_regfile_mem_15__6_), .Y(_2242_) );
NAND2X1 NAND2X1_1125 ( .A(datapath_1_RegisterFile_regfile_mem_13__6_), .B(_1884__bF_buf8), .Y(_2243_) );
NAND3X1 NAND3X1_1445 ( .A(datapath_1_Instr_21_bF_buf23_), .B(_2242_), .C(_2243_), .Y(_2244_) );
NAND2X1 NAND2X1_1126 ( .A(datapath_1_Instr_22_bF_buf23_), .B(datapath_1_RegisterFile_regfile_mem_14__6_), .Y(_2245_) );
AOI21X1 AOI21X1_645 ( .A(_1884__bF_buf8), .B(datapath_1_RegisterFile_regfile_mem_12__6_), .C(datapath_1_Instr_21_bF_buf22_), .Y(_2246_) );
NAND2X1 NAND2X1_1127 ( .A(_2245_), .B(_2246_), .Y(_2247_) );
NAND3X1 NAND3X1_1446 ( .A(datapath_1_Instr_23_bF_buf8_bF_buf3_), .B(_2244_), .C(_2247_), .Y(_2248_) );
AOI21X1 AOI21X1_646 ( .A(_2241_), .B(_2248_), .C(_1888__bF_buf7), .Y(_2249_) );
INVX1 INVX1_401 ( .A(datapath_1_RegisterFile_regfile_mem_1__6_), .Y(_2250_) );
AOI21X1 AOI21X1_647 ( .A(datapath_1_Instr_23_bF_buf7_bF_buf3_), .B(datapath_1_RegisterFile_regfile_mem_5__6_), .C(_1890__bF_buf41), .Y(_2251_) );
OAI21X1 OAI21X1_1709 ( .A(datapath_1_Instr_23_bF_buf6_bF_buf3_), .B(_2250_), .C(_2251_), .Y(_2252_) );
INVX1 INVX1_402 ( .A(datapath_1_RegisterFile_regfile_mem_0__6_), .Y(_2253_) );
AOI21X1 AOI21X1_648 ( .A(datapath_1_Instr_23_bF_buf5_bF_buf3_), .B(datapath_1_RegisterFile_regfile_mem_4__6_), .C(datapath_1_Instr_21_bF_buf21_), .Y(_2254_) );
OAI21X1 OAI21X1_1710 ( .A(datapath_1_Instr_23_bF_buf4_bF_buf3_), .B(_2253_), .C(_2254_), .Y(_2255_) );
NAND3X1 NAND3X1_1447 ( .A(_1884__bF_buf4), .B(_2255_), .C(_2252_), .Y(_2256_) );
INVX1 INVX1_403 ( .A(datapath_1_RegisterFile_regfile_mem_3__6_), .Y(_2257_) );
AOI21X1 AOI21X1_649 ( .A(datapath_1_Instr_23_bF_buf3_bF_buf3_), .B(datapath_1_RegisterFile_regfile_mem_7__6_), .C(_1890__bF_buf41), .Y(_2258_) );
OAI21X1 OAI21X1_1711 ( .A(datapath_1_Instr_23_bF_buf2_bF_buf3_), .B(_2257_), .C(_2258_), .Y(_2259_) );
INVX1 INVX1_404 ( .A(datapath_1_RegisterFile_regfile_mem_2__6_), .Y(_2260_) );
AOI21X1 AOI21X1_650 ( .A(datapath_1_Instr_23_bF_buf1_), .B(datapath_1_RegisterFile_regfile_mem_6__6_), .C(datapath_1_Instr_21_bF_buf20_), .Y(_2261_) );
OAI21X1 OAI21X1_1712 ( .A(datapath_1_Instr_23_bF_buf0_), .B(_2260_), .C(_2261_), .Y(_2262_) );
NAND3X1 NAND3X1_1448 ( .A(datapath_1_Instr_22_bF_buf22_), .B(_2262_), .C(_2259_), .Y(_2263_) );
AOI21X1 AOI21X1_651 ( .A(_2256_), .B(_2263_), .C(datapath_1_Instr_24_bF_buf4_), .Y(_2264_) );
OAI21X1 OAI21X1_1713 ( .A(_2264_), .B(_2249_), .C(_1917__bF_buf3), .Y(_2265_) );
AOI22X1 AOI22X1_137 ( .A(_1883__bF_buf0), .B(_1887__bF_buf2), .C(_2265_), .D(_2234_), .Y(datapath_1_RD1_6_) );
NAND2X1 NAND2X1_1128 ( .A(datapath_1_Instr_21_bF_buf19_), .B(datapath_1_RegisterFile_regfile_mem_27__7_), .Y(_2266_) );
NAND2X1 NAND2X1_1129 ( .A(datapath_1_RegisterFile_regfile_mem_26__7_), .B(_1890__bF_buf17), .Y(_2267_) );
NAND3X1 NAND3X1_1449 ( .A(datapath_1_Instr_22_bF_buf21_), .B(_2266_), .C(_2267_), .Y(_2268_) );
NAND2X1 NAND2X1_1130 ( .A(datapath_1_Instr_21_bF_buf18_), .B(datapath_1_RegisterFile_regfile_mem_25__7_), .Y(_2269_) );
AOI21X1 AOI21X1_652 ( .A(_1890__bF_buf17), .B(datapath_1_RegisterFile_regfile_mem_24__7_), .C(datapath_1_Instr_22_bF_buf20_), .Y(_2270_) );
NAND2X1 NAND2X1_1131 ( .A(_2269_), .B(_2270_), .Y(_2271_) );
NAND3X1 NAND3X1_1450 ( .A(_1885__bF_buf10), .B(_2268_), .C(_2271_), .Y(_2272_) );
NAND2X1 NAND2X1_1132 ( .A(datapath_1_Instr_21_bF_buf17_), .B(datapath_1_RegisterFile_regfile_mem_31__7_), .Y(_2273_) );
AOI21X1 AOI21X1_653 ( .A(_1890__bF_buf17), .B(datapath_1_RegisterFile_regfile_mem_30__7_), .C(_1884__bF_buf6), .Y(_2274_) );
NAND2X1 NAND2X1_1133 ( .A(_2273_), .B(_2274_), .Y(_2275_) );
INVX1 INVX1_405 ( .A(datapath_1_RegisterFile_regfile_mem_28__7_), .Y(_2276_) );
AOI21X1 AOI21X1_654 ( .A(datapath_1_Instr_21_bF_buf16_), .B(datapath_1_RegisterFile_regfile_mem_29__7_), .C(datapath_1_Instr_22_bF_buf19_), .Y(_2277_) );
OAI21X1 OAI21X1_1714 ( .A(datapath_1_Instr_21_bF_buf15_), .B(_2276_), .C(_2277_), .Y(_2278_) );
NAND3X1 NAND3X1_1451 ( .A(datapath_1_Instr_23_bF_buf15_bF_buf2_), .B(_2278_), .C(_2275_), .Y(_2279_) );
AOI21X1 AOI21X1_655 ( .A(_2272_), .B(_2279_), .C(_1888__bF_buf3), .Y(_2280_) );
MUX2X1 MUX2X1_158 ( .A(datapath_1_RegisterFile_regfile_mem_18__7_), .B(datapath_1_RegisterFile_regfile_mem_16__7_), .S(datapath_1_Instr_22_bF_buf18_), .Y(_2281_) );
NAND2X1 NAND2X1_1134 ( .A(_1890__bF_buf31), .B(_2281_), .Y(_2282_) );
MUX2X1 MUX2X1_159 ( .A(datapath_1_RegisterFile_regfile_mem_19__7_), .B(datapath_1_RegisterFile_regfile_mem_17__7_), .S(datapath_1_Instr_22_bF_buf17_), .Y(_2283_) );
NAND2X1 NAND2X1_1135 ( .A(datapath_1_Instr_21_bF_buf14_), .B(_2283_), .Y(_2284_) );
NAND3X1 NAND3X1_1452 ( .A(_1885__bF_buf7), .B(_2282_), .C(_2284_), .Y(_2285_) );
MUX2X1 MUX2X1_160 ( .A(datapath_1_RegisterFile_regfile_mem_22__7_), .B(datapath_1_RegisterFile_regfile_mem_20__7_), .S(datapath_1_Instr_22_bF_buf16_), .Y(_2286_) );
NAND2X1 NAND2X1_1136 ( .A(_1890__bF_buf31), .B(_2286_), .Y(_2287_) );
MUX2X1 MUX2X1_161 ( .A(datapath_1_RegisterFile_regfile_mem_23__7_), .B(datapath_1_RegisterFile_regfile_mem_21__7_), .S(datapath_1_Instr_22_bF_buf15_), .Y(_2288_) );
NAND2X1 NAND2X1_1137 ( .A(datapath_1_Instr_21_bF_buf13_), .B(_2288_), .Y(_2289_) );
NAND3X1 NAND3X1_1453 ( .A(datapath_1_Instr_23_bF_buf14_bF_buf2_), .B(_2287_), .C(_2289_), .Y(_2290_) );
AOI21X1 AOI21X1_656 ( .A(_2285_), .B(_2290_), .C(datapath_1_Instr_24_bF_buf3_), .Y(_2291_) );
OAI21X1 OAI21X1_1715 ( .A(_2291_), .B(_2280_), .C(datapath_1_Instr_25_bF_buf0_), .Y(_2292_) );
MUX2X1 MUX2X1_162 ( .A(datapath_1_RegisterFile_regfile_mem_9__7_), .B(datapath_1_RegisterFile_regfile_mem_8__7_), .S(datapath_1_Instr_21_bF_buf12_), .Y(_2293_) );
NOR2X1 NOR2X1_354 ( .A(datapath_1_RegisterFile_regfile_mem_11__7_), .B(_1890__bF_buf42), .Y(_2294_) );
OAI21X1 OAI21X1_1716 ( .A(datapath_1_Instr_21_bF_buf11_), .B(datapath_1_RegisterFile_regfile_mem_10__7_), .C(datapath_1_Instr_22_bF_buf14_), .Y(_2295_) );
OAI22X1 OAI22X1_156 ( .A(_2295_), .B(_2294_), .C(datapath_1_Instr_22_bF_buf13_), .D(_2293_), .Y(_2296_) );
INVX1 INVX1_406 ( .A(datapath_1_RegisterFile_regfile_mem_15__7_), .Y(_2297_) );
AOI21X1 AOI21X1_657 ( .A(_1890__bF_buf23), .B(datapath_1_RegisterFile_regfile_mem_14__7_), .C(_1884__bF_buf7), .Y(_2298_) );
OAI21X1 OAI21X1_1717 ( .A(_1890__bF_buf42), .B(_2297_), .C(_2298_), .Y(_2299_) );
NAND2X1 NAND2X1_1138 ( .A(datapath_1_RegisterFile_regfile_mem_12__7_), .B(_1890__bF_buf42), .Y(_2300_) );
AOI21X1 AOI21X1_658 ( .A(datapath_1_Instr_21_bF_buf10_), .B(datapath_1_RegisterFile_regfile_mem_13__7_), .C(datapath_1_Instr_22_bF_buf12_), .Y(_2301_) );
AOI21X1 AOI21X1_659 ( .A(_2300_), .B(_2301_), .C(_1885__bF_buf8), .Y(_2302_) );
AOI22X1 AOI22X1_138 ( .A(_2299_), .B(_2302_), .C(_1885__bF_buf8), .D(_2296_), .Y(_2303_) );
NOR2X1 NOR2X1_355 ( .A(datapath_1_Instr_21_bF_buf9_), .B(datapath_1_RegisterFile_regfile_mem_0__7_), .Y(_2304_) );
OAI21X1 OAI21X1_1718 ( .A(datapath_1_RegisterFile_regfile_mem_1__7_), .B(_1890__bF_buf0), .C(_1884__bF_buf7), .Y(_2305_) );
NOR2X1 NOR2X1_356 ( .A(datapath_1_RegisterFile_regfile_mem_3__7_), .B(_1890__bF_buf0), .Y(_2306_) );
OAI21X1 OAI21X1_1719 ( .A(datapath_1_Instr_21_bF_buf8_), .B(datapath_1_RegisterFile_regfile_mem_2__7_), .C(datapath_1_Instr_22_bF_buf11_), .Y(_2307_) );
OAI22X1 OAI22X1_157 ( .A(_2306_), .B(_2307_), .C(_2304_), .D(_2305_), .Y(_2308_) );
NOR2X1 NOR2X1_357 ( .A(datapath_1_Instr_23_bF_buf13_bF_buf2_), .B(_2308_), .Y(_2309_) );
MUX2X1 MUX2X1_163 ( .A(datapath_1_RegisterFile_regfile_mem_5__7_), .B(datapath_1_RegisterFile_regfile_mem_4__7_), .S(datapath_1_Instr_21_bF_buf7_), .Y(_2310_) );
NOR2X1 NOR2X1_358 ( .A(datapath_1_RegisterFile_regfile_mem_7__7_), .B(_1890__bF_buf42), .Y(_2311_) );
OAI21X1 OAI21X1_1720 ( .A(datapath_1_Instr_21_bF_buf6_), .B(datapath_1_RegisterFile_regfile_mem_6__7_), .C(datapath_1_Instr_22_bF_buf10_), .Y(_2312_) );
OAI22X1 OAI22X1_158 ( .A(_2312_), .B(_2311_), .C(datapath_1_Instr_22_bF_buf9_), .D(_2310_), .Y(_2313_) );
OAI21X1 OAI21X1_1721 ( .A(_1885__bF_buf8), .B(_2313_), .C(_1888__bF_buf4), .Y(_2314_) );
OAI22X1 OAI22X1_159 ( .A(_1888__bF_buf4), .B(_2303_), .C(_2309_), .D(_2314_), .Y(_2315_) );
NAND2X1 NAND2X1_1139 ( .A(_1917__bF_buf1), .B(_2315_), .Y(_2316_) );
AOI22X1 AOI22X1_139 ( .A(_1883__bF_buf3), .B(_1887__bF_buf1), .C(_2292_), .D(_2316_), .Y(datapath_1_RD1_7_) );
MUX2X1 MUX2X1_164 ( .A(datapath_1_RegisterFile_regfile_mem_9__8_), .B(datapath_1_RegisterFile_regfile_mem_8__8_), .S(datapath_1_Instr_21_bF_buf5_), .Y(_2317_) );
NOR2X1 NOR2X1_359 ( .A(datapath_1_RegisterFile_regfile_mem_11__8_), .B(_1890__bF_buf21), .Y(_2318_) );
OAI21X1 OAI21X1_1722 ( .A(datapath_1_Instr_21_bF_buf4_), .B(datapath_1_RegisterFile_regfile_mem_10__8_), .C(datapath_1_Instr_22_bF_buf8_), .Y(_2319_) );
OAI22X1 OAI22X1_160 ( .A(_2319_), .B(_2318_), .C(datapath_1_Instr_22_bF_buf7_), .D(_2317_), .Y(_2320_) );
INVX1 INVX1_407 ( .A(datapath_1_RegisterFile_regfile_mem_15__8_), .Y(_2321_) );
AOI21X1 AOI21X1_660 ( .A(_1890__bF_buf21), .B(datapath_1_RegisterFile_regfile_mem_14__8_), .C(_1884__bF_buf1), .Y(_2322_) );
OAI21X1 OAI21X1_1723 ( .A(_1890__bF_buf21), .B(_2321_), .C(_2322_), .Y(_2323_) );
NAND2X1 NAND2X1_1140 ( .A(datapath_1_RegisterFile_regfile_mem_12__8_), .B(_1890__bF_buf21), .Y(_2324_) );
AOI21X1 AOI21X1_661 ( .A(datapath_1_Instr_21_bF_buf3_), .B(datapath_1_RegisterFile_regfile_mem_13__8_), .C(datapath_1_Instr_22_bF_buf6_), .Y(_2325_) );
AOI21X1 AOI21X1_662 ( .A(_2324_), .B(_2325_), .C(_1885__bF_buf0), .Y(_2326_) );
AOI22X1 AOI22X1_140 ( .A(_2323_), .B(_2326_), .C(_1885__bF_buf0), .D(_2320_), .Y(_2327_) );
NOR2X1 NOR2X1_360 ( .A(datapath_1_Instr_21_bF_buf2_), .B(datapath_1_RegisterFile_regfile_mem_0__8_), .Y(_2328_) );
OAI21X1 OAI21X1_1724 ( .A(datapath_1_RegisterFile_regfile_mem_1__8_), .B(_1890__bF_buf38), .C(_1884__bF_buf4), .Y(_2329_) );
NOR2X1 NOR2X1_361 ( .A(datapath_1_RegisterFile_regfile_mem_3__8_), .B(_1890__bF_buf38), .Y(_2330_) );
OAI21X1 OAI21X1_1725 ( .A(datapath_1_Instr_21_bF_buf1_), .B(datapath_1_RegisterFile_regfile_mem_2__8_), .C(datapath_1_Instr_22_bF_buf5_), .Y(_2331_) );
OAI22X1 OAI22X1_161 ( .A(_2330_), .B(_2331_), .C(_2328_), .D(_2329_), .Y(_2332_) );
NOR2X1 NOR2X1_362 ( .A(datapath_1_Instr_23_bF_buf12_bF_buf2_), .B(_2332_), .Y(_2333_) );
MUX2X1 MUX2X1_165 ( .A(datapath_1_RegisterFile_regfile_mem_5__8_), .B(datapath_1_RegisterFile_regfile_mem_4__8_), .S(datapath_1_Instr_21_bF_buf0_), .Y(_2334_) );
NOR2X1 NOR2X1_363 ( .A(datapath_1_RegisterFile_regfile_mem_7__8_), .B(_1890__bF_buf27), .Y(_2335_) );
OAI21X1 OAI21X1_1726 ( .A(datapath_1_Instr_21_bF_buf55_), .B(datapath_1_RegisterFile_regfile_mem_6__8_), .C(datapath_1_Instr_22_bF_buf4_), .Y(_2336_) );
OAI22X1 OAI22X1_162 ( .A(_2336_), .B(_2335_), .C(datapath_1_Instr_22_bF_buf3_), .D(_2334_), .Y(_2337_) );
OAI21X1 OAI21X1_1727 ( .A(_1885__bF_buf4), .B(_2337_), .C(_1888__bF_buf6), .Y(_2338_) );
OAI22X1 OAI22X1_163 ( .A(_1888__bF_buf6), .B(_2327_), .C(_2333_), .D(_2338_), .Y(_2339_) );
NAND2X1 NAND2X1_1141 ( .A(_1917__bF_buf3), .B(_2339_), .Y(_2340_) );
INVX1 INVX1_408 ( .A(datapath_1_RegisterFile_regfile_mem_19__8_), .Y(_2341_) );
AOI21X1 AOI21X1_663 ( .A(datapath_1_Instr_23_bF_buf11_bF_buf2_), .B(datapath_1_RegisterFile_regfile_mem_23__8_), .C(_1890__bF_buf25), .Y(_2342_) );
OAI21X1 OAI21X1_1728 ( .A(datapath_1_Instr_23_bF_buf10_bF_buf2_), .B(_2341_), .C(_2342_), .Y(_2343_) );
NAND2X1 NAND2X1_1142 ( .A(datapath_1_RegisterFile_regfile_mem_18__8_), .B(_1885__bF_buf11), .Y(_2344_) );
AOI21X1 AOI21X1_664 ( .A(datapath_1_Instr_23_bF_buf9_bF_buf2_), .B(datapath_1_RegisterFile_regfile_mem_22__8_), .C(datapath_1_Instr_21_bF_buf54_), .Y(_2345_) );
AOI21X1 AOI21X1_665 ( .A(_2344_), .B(_2345_), .C(_1884__bF_buf2), .Y(_2346_) );
INVX1 INVX1_409 ( .A(datapath_1_RegisterFile_regfile_mem_17__8_), .Y(_2347_) );
AOI21X1 AOI21X1_666 ( .A(datapath_1_Instr_23_bF_buf8_bF_buf2_), .B(datapath_1_RegisterFile_regfile_mem_21__8_), .C(_1890__bF_buf36), .Y(_2348_) );
OAI21X1 OAI21X1_1729 ( .A(datapath_1_Instr_23_bF_buf7_bF_buf2_), .B(_2347_), .C(_2348_), .Y(_2349_) );
NAND2X1 NAND2X1_1143 ( .A(datapath_1_RegisterFile_regfile_mem_16__8_), .B(_1885__bF_buf11), .Y(_2350_) );
AOI21X1 AOI21X1_667 ( .A(datapath_1_Instr_23_bF_buf6_bF_buf2_), .B(datapath_1_RegisterFile_regfile_mem_20__8_), .C(datapath_1_Instr_21_bF_buf53_), .Y(_2351_) );
AOI21X1 AOI21X1_668 ( .A(_2350_), .B(_2351_), .C(datapath_1_Instr_22_bF_buf2_), .Y(_2352_) );
AOI22X1 AOI22X1_141 ( .A(_2346_), .B(_2343_), .C(_2349_), .D(_2352_), .Y(_2353_) );
NOR2X1 NOR2X1_364 ( .A(datapath_1_Instr_21_bF_buf52_), .B(datapath_1_RegisterFile_regfile_mem_24__8_), .Y(_2354_) );
OAI21X1 OAI21X1_1730 ( .A(datapath_1_RegisterFile_regfile_mem_25__8_), .B(_1890__bF_buf25), .C(_1884__bF_buf2), .Y(_2355_) );
NOR2X1 NOR2X1_365 ( .A(datapath_1_RegisterFile_regfile_mem_27__8_), .B(_1890__bF_buf25), .Y(_2356_) );
OAI21X1 OAI21X1_1731 ( .A(datapath_1_Instr_21_bF_buf51_), .B(datapath_1_RegisterFile_regfile_mem_26__8_), .C(datapath_1_Instr_22_bF_buf1_), .Y(_2357_) );
OAI22X1 OAI22X1_164 ( .A(_2356_), .B(_2357_), .C(_2354_), .D(_2355_), .Y(_2358_) );
NOR2X1 NOR2X1_366 ( .A(datapath_1_Instr_23_bF_buf5_bF_buf2_), .B(_2358_), .Y(_2359_) );
MUX2X1 MUX2X1_166 ( .A(datapath_1_RegisterFile_regfile_mem_29__8_), .B(datapath_1_RegisterFile_regfile_mem_28__8_), .S(datapath_1_Instr_21_bF_buf50_), .Y(_2360_) );
NOR2X1 NOR2X1_367 ( .A(datapath_1_RegisterFile_regfile_mem_31__8_), .B(_1890__bF_buf36), .Y(_2361_) );
OAI21X1 OAI21X1_1732 ( .A(datapath_1_Instr_21_bF_buf49_), .B(datapath_1_RegisterFile_regfile_mem_30__8_), .C(datapath_1_Instr_22_bF_buf0_), .Y(_2362_) );
OAI22X1 OAI22X1_165 ( .A(_2362_), .B(_2361_), .C(datapath_1_Instr_22_bF_buf50_), .D(_2360_), .Y(_2363_) );
OAI21X1 OAI21X1_1733 ( .A(_1885__bF_buf11), .B(_2363_), .C(datapath_1_Instr_24_bF_buf2_), .Y(_2364_) );
OAI22X1 OAI22X1_166 ( .A(datapath_1_Instr_24_bF_buf1_), .B(_2353_), .C(_2359_), .D(_2364_), .Y(_2365_) );
NAND2X1 NAND2X1_1144 ( .A(datapath_1_Instr_25_bF_buf5_), .B(_2365_), .Y(_2366_) );
AOI22X1 AOI22X1_142 ( .A(_1883__bF_buf0), .B(_1887__bF_buf2), .C(_2366_), .D(_2340_), .Y(datapath_1_RD1_8_) );
INVX1 INVX1_410 ( .A(datapath_1_RegisterFile_regfile_mem_1__9_), .Y(_2367_) );
AOI21X1 AOI21X1_669 ( .A(datapath_1_Instr_23_bF_buf4_bF_buf2_), .B(datapath_1_RegisterFile_regfile_mem_5__9_), .C(_1890__bF_buf5), .Y(_2368_) );
OAI21X1 OAI21X1_1734 ( .A(datapath_1_Instr_23_bF_buf3_bF_buf2_), .B(_2367_), .C(_2368_), .Y(_2369_) );
INVX1 INVX1_411 ( .A(datapath_1_RegisterFile_regfile_mem_0__9_), .Y(_2370_) );
AOI21X1 AOI21X1_670 ( .A(datapath_1_Instr_23_bF_buf2_bF_buf2_), .B(datapath_1_RegisterFile_regfile_mem_4__9_), .C(datapath_1_Instr_21_bF_buf48_), .Y(_2371_) );
OAI21X1 OAI21X1_1735 ( .A(datapath_1_Instr_23_bF_buf1_), .B(_2370_), .C(_2371_), .Y(_2372_) );
NAND3X1 NAND3X1_1454 ( .A(_1884__bF_buf3), .B(_2372_), .C(_2369_), .Y(_2373_) );
INVX1 INVX1_412 ( .A(datapath_1_RegisterFile_regfile_mem_3__9_), .Y(_2374_) );
AOI21X1 AOI21X1_671 ( .A(datapath_1_Instr_23_bF_buf0_), .B(datapath_1_RegisterFile_regfile_mem_7__9_), .C(_1890__bF_buf5), .Y(_2375_) );
OAI21X1 OAI21X1_1736 ( .A(datapath_1_Instr_23_bF_buf15_bF_buf1_), .B(_2374_), .C(_2375_), .Y(_2376_) );
INVX1 INVX1_413 ( .A(datapath_1_RegisterFile_regfile_mem_2__9_), .Y(_2377_) );
AOI21X1 AOI21X1_672 ( .A(datapath_1_Instr_23_bF_buf14_bF_buf1_), .B(datapath_1_RegisterFile_regfile_mem_6__9_), .C(datapath_1_Instr_21_bF_buf47_), .Y(_2378_) );
OAI21X1 OAI21X1_1737 ( .A(datapath_1_Instr_23_bF_buf13_bF_buf1_), .B(_2377_), .C(_2378_), .Y(_2379_) );
NAND3X1 NAND3X1_1455 ( .A(datapath_1_Instr_22_bF_buf49_), .B(_2379_), .C(_2376_), .Y(_2380_) );
AOI21X1 AOI21X1_673 ( .A(_2373_), .B(_2380_), .C(datapath_1_Instr_24_bF_buf0_), .Y(_2381_) );
NAND2X1 NAND2X1_1145 ( .A(datapath_1_Instr_22_bF_buf48_), .B(datapath_1_RegisterFile_regfile_mem_11__9_), .Y(_2382_) );
NAND2X1 NAND2X1_1146 ( .A(datapath_1_RegisterFile_regfile_mem_9__9_), .B(_1884__bF_buf5), .Y(_2383_) );
NAND3X1 NAND3X1_1456 ( .A(datapath_1_Instr_21_bF_buf46_), .B(_2382_), .C(_2383_), .Y(_2384_) );
NAND2X1 NAND2X1_1147 ( .A(datapath_1_Instr_22_bF_buf47_), .B(datapath_1_RegisterFile_regfile_mem_10__9_), .Y(_2385_) );
AOI21X1 AOI21X1_674 ( .A(_1884__bF_buf5), .B(datapath_1_RegisterFile_regfile_mem_8__9_), .C(datapath_1_Instr_21_bF_buf45_), .Y(_2386_) );
NAND2X1 NAND2X1_1148 ( .A(_2385_), .B(_2386_), .Y(_2387_) );
NAND3X1 NAND3X1_1457 ( .A(_1885__bF_buf1), .B(_2384_), .C(_2387_), .Y(_2388_) );
NAND2X1 NAND2X1_1149 ( .A(datapath_1_Instr_22_bF_buf46_), .B(datapath_1_RegisterFile_regfile_mem_15__9_), .Y(_2389_) );
NAND2X1 NAND2X1_1150 ( .A(datapath_1_RegisterFile_regfile_mem_13__9_), .B(_1884__bF_buf5), .Y(_2390_) );
NAND3X1 NAND3X1_1458 ( .A(datapath_1_Instr_21_bF_buf44_), .B(_2389_), .C(_2390_), .Y(_2391_) );
NAND2X1 NAND2X1_1151 ( .A(datapath_1_Instr_22_bF_buf45_), .B(datapath_1_RegisterFile_regfile_mem_14__9_), .Y(_2392_) );
AOI21X1 AOI21X1_675 ( .A(_1884__bF_buf5), .B(datapath_1_RegisterFile_regfile_mem_12__9_), .C(datapath_1_Instr_21_bF_buf43_), .Y(_2393_) );
NAND2X1 NAND2X1_1152 ( .A(_2392_), .B(_2393_), .Y(_2394_) );
NAND3X1 NAND3X1_1459 ( .A(datapath_1_Instr_23_bF_buf12_bF_buf1_), .B(_2391_), .C(_2394_), .Y(_2395_) );
AOI21X1 AOI21X1_676 ( .A(_2388_), .B(_2395_), .C(_1888__bF_buf5), .Y(_2396_) );
OAI21X1 OAI21X1_1738 ( .A(_2381_), .B(_2396_), .C(_1917__bF_buf4), .Y(_2397_) );
MUX2X1 MUX2X1_167 ( .A(datapath_1_RegisterFile_regfile_mem_17__9_), .B(datapath_1_RegisterFile_regfile_mem_16__9_), .S(datapath_1_Instr_21_bF_buf42_), .Y(_2398_) );
NOR2X1 NOR2X1_368 ( .A(datapath_1_RegisterFile_regfile_mem_19__9_), .B(_1890__bF_buf39), .Y(_2399_) );
OAI21X1 OAI21X1_1739 ( .A(datapath_1_Instr_21_bF_buf41_), .B(datapath_1_RegisterFile_regfile_mem_18__9_), .C(datapath_1_Instr_22_bF_buf44_), .Y(_2400_) );
OAI22X1 OAI22X1_167 ( .A(_2400_), .B(_2399_), .C(datapath_1_Instr_22_bF_buf43_), .D(_2398_), .Y(_2401_) );
NAND2X1 NAND2X1_1153 ( .A(_1885__bF_buf6), .B(_2401_), .Y(_2402_) );
MUX2X1 MUX2X1_168 ( .A(datapath_1_RegisterFile_regfile_mem_21__9_), .B(datapath_1_RegisterFile_regfile_mem_20__9_), .S(datapath_1_Instr_21_bF_buf40_), .Y(_2403_) );
NOR2X1 NOR2X1_369 ( .A(datapath_1_RegisterFile_regfile_mem_23__9_), .B(_1890__bF_buf39), .Y(_2404_) );
OAI21X1 OAI21X1_1740 ( .A(datapath_1_Instr_21_bF_buf39_), .B(datapath_1_RegisterFile_regfile_mem_22__9_), .C(datapath_1_Instr_22_bF_buf42_), .Y(_2405_) );
OAI22X1 OAI22X1_168 ( .A(_2405_), .B(_2404_), .C(datapath_1_Instr_22_bF_buf41_), .D(_2403_), .Y(_2406_) );
NAND2X1 NAND2X1_1154 ( .A(datapath_1_Instr_23_bF_buf11_bF_buf1_), .B(_2406_), .Y(_2407_) );
AOI21X1 AOI21X1_677 ( .A(_2402_), .B(_2407_), .C(datapath_1_Instr_24_bF_buf6_), .Y(_2408_) );
INVX1 INVX1_414 ( .A(datapath_1_RegisterFile_regfile_mem_27__9_), .Y(_2409_) );
AOI21X1 AOI21X1_678 ( .A(datapath_1_Instr_23_bF_buf10_bF_buf1_), .B(datapath_1_RegisterFile_regfile_mem_31__9_), .C(_1890__bF_buf4), .Y(_2410_) );
OAI21X1 OAI21X1_1741 ( .A(datapath_1_Instr_23_bF_buf9_bF_buf1_), .B(_2409_), .C(_2410_), .Y(_2411_) );
INVX1 INVX1_415 ( .A(datapath_1_RegisterFile_regfile_mem_26__9_), .Y(_2412_) );
AOI21X1 AOI21X1_679 ( .A(datapath_1_Instr_23_bF_buf8_bF_buf1_), .B(datapath_1_RegisterFile_regfile_mem_30__9_), .C(datapath_1_Instr_21_bF_buf38_), .Y(_2413_) );
OAI21X1 OAI21X1_1742 ( .A(datapath_1_Instr_23_bF_buf7_bF_buf1_), .B(_2412_), .C(_2413_), .Y(_2414_) );
NAND3X1 NAND3X1_1460 ( .A(datapath_1_Instr_22_bF_buf40_), .B(_2414_), .C(_2411_), .Y(_2415_) );
INVX1 INVX1_416 ( .A(datapath_1_RegisterFile_regfile_mem_25__9_), .Y(_2416_) );
AOI21X1 AOI21X1_680 ( .A(datapath_1_Instr_23_bF_buf6_bF_buf1_), .B(datapath_1_RegisterFile_regfile_mem_29__9_), .C(_1890__bF_buf1), .Y(_2417_) );
OAI21X1 OAI21X1_1743 ( .A(datapath_1_Instr_23_bF_buf5_bF_buf1_), .B(_2416_), .C(_2417_), .Y(_2418_) );
INVX1 INVX1_417 ( .A(datapath_1_RegisterFile_regfile_mem_24__9_), .Y(_2419_) );
AOI21X1 AOI21X1_681 ( .A(datapath_1_Instr_23_bF_buf4_bF_buf1_), .B(datapath_1_RegisterFile_regfile_mem_28__9_), .C(datapath_1_Instr_21_bF_buf37_), .Y(_2420_) );
OAI21X1 OAI21X1_1744 ( .A(datapath_1_Instr_23_bF_buf3_bF_buf1_), .B(_2419_), .C(_2420_), .Y(_2421_) );
NAND3X1 NAND3X1_1461 ( .A(_1884__bF_buf9), .B(_2421_), .C(_2418_), .Y(_2422_) );
AOI21X1 AOI21X1_682 ( .A(_2415_), .B(_2422_), .C(_1888__bF_buf1), .Y(_2423_) );
OAI21X1 OAI21X1_1745 ( .A(_2423_), .B(_2408_), .C(datapath_1_Instr_25_bF_buf4_), .Y(_2424_) );
AOI22X1 AOI22X1_143 ( .A(_1883__bF_buf4), .B(_1887__bF_buf3), .C(_2397_), .D(_2424_), .Y(datapath_1_RD1_9_) );
NAND2X1 NAND2X1_1155 ( .A(datapath_1_Instr_21_bF_buf36_), .B(datapath_1_RegisterFile_regfile_mem_27__10_), .Y(_2425_) );
NAND2X1 NAND2X1_1156 ( .A(datapath_1_RegisterFile_regfile_mem_26__10_), .B(_1890__bF_buf4), .Y(_2426_) );
NAND3X1 NAND3X1_1462 ( .A(datapath_1_Instr_22_bF_buf39_), .B(_2425_), .C(_2426_), .Y(_2427_) );
NAND2X1 NAND2X1_1157 ( .A(datapath_1_Instr_21_bF_buf35_), .B(datapath_1_RegisterFile_regfile_mem_25__10_), .Y(_2428_) );
AOI21X1 AOI21X1_683 ( .A(_1890__bF_buf4), .B(datapath_1_RegisterFile_regfile_mem_24__10_), .C(datapath_1_Instr_22_bF_buf38_), .Y(_2429_) );
NAND2X1 NAND2X1_1158 ( .A(_2428_), .B(_2429_), .Y(_2430_) );
NAND3X1 NAND3X1_1463 ( .A(_1885__bF_buf6), .B(_2427_), .C(_2430_), .Y(_2431_) );
NAND2X1 NAND2X1_1159 ( .A(datapath_1_Instr_21_bF_buf34_), .B(datapath_1_RegisterFile_regfile_mem_31__10_), .Y(_2432_) );
AOI21X1 AOI21X1_684 ( .A(_1890__bF_buf4), .B(datapath_1_RegisterFile_regfile_mem_30__10_), .C(_1884__bF_buf3), .Y(_2433_) );
NAND2X1 NAND2X1_1160 ( .A(_2432_), .B(_2433_), .Y(_2434_) );
INVX1 INVX1_418 ( .A(datapath_1_RegisterFile_regfile_mem_28__10_), .Y(_2435_) );
AOI21X1 AOI21X1_685 ( .A(datapath_1_Instr_21_bF_buf33_), .B(datapath_1_RegisterFile_regfile_mem_29__10_), .C(datapath_1_Instr_22_bF_buf37_), .Y(_2436_) );
OAI21X1 OAI21X1_1746 ( .A(datapath_1_Instr_21_bF_buf32_), .B(_2435_), .C(_2436_), .Y(_2437_) );
NAND3X1 NAND3X1_1464 ( .A(datapath_1_Instr_23_bF_buf2_bF_buf1_), .B(_2437_), .C(_2434_), .Y(_2438_) );
AOI21X1 AOI21X1_686 ( .A(_2431_), .B(_2438_), .C(_1888__bF_buf1), .Y(_2439_) );
MUX2X1 MUX2X1_169 ( .A(datapath_1_RegisterFile_regfile_mem_18__10_), .B(datapath_1_RegisterFile_regfile_mem_16__10_), .S(datapath_1_Instr_22_bF_buf36_), .Y(_2440_) );
NAND2X1 NAND2X1_1161 ( .A(_1890__bF_buf24), .B(_2440_), .Y(_2441_) );
MUX2X1 MUX2X1_170 ( .A(datapath_1_RegisterFile_regfile_mem_19__10_), .B(datapath_1_RegisterFile_regfile_mem_17__10_), .S(datapath_1_Instr_22_bF_buf35_), .Y(_2442_) );
NAND2X1 NAND2X1_1162 ( .A(datapath_1_Instr_21_bF_buf31_), .B(_2442_), .Y(_2443_) );
NAND3X1 NAND3X1_1465 ( .A(_1885__bF_buf6), .B(_2441_), .C(_2443_), .Y(_2444_) );
MUX2X1 MUX2X1_171 ( .A(datapath_1_RegisterFile_regfile_mem_22__10_), .B(datapath_1_RegisterFile_regfile_mem_20__10_), .S(datapath_1_Instr_22_bF_buf34_), .Y(_2445_) );
NAND2X1 NAND2X1_1163 ( .A(_1890__bF_buf4), .B(_2445_), .Y(_2446_) );
MUX2X1 MUX2X1_172 ( .A(datapath_1_RegisterFile_regfile_mem_23__10_), .B(datapath_1_RegisterFile_regfile_mem_21__10_), .S(datapath_1_Instr_22_bF_buf33_), .Y(_2447_) );
NAND2X1 NAND2X1_1164 ( .A(datapath_1_Instr_21_bF_buf30_), .B(_2447_), .Y(_2448_) );
NAND3X1 NAND3X1_1466 ( .A(datapath_1_Instr_23_bF_buf1_), .B(_2446_), .C(_2448_), .Y(_2449_) );
AOI21X1 AOI21X1_687 ( .A(_2444_), .B(_2449_), .C(datapath_1_Instr_24_bF_buf5_), .Y(_2450_) );
OAI21X1 OAI21X1_1747 ( .A(_2450_), .B(_2439_), .C(datapath_1_Instr_25_bF_buf3_), .Y(_2451_) );
MUX2X1 MUX2X1_173 ( .A(datapath_1_RegisterFile_regfile_mem_9__10_), .B(datapath_1_RegisterFile_regfile_mem_8__10_), .S(datapath_1_Instr_21_bF_buf29_), .Y(_2452_) );
NOR2X1 NOR2X1_370 ( .A(datapath_1_RegisterFile_regfile_mem_11__10_), .B(_1890__bF_buf26), .Y(_2453_) );
OAI21X1 OAI21X1_1748 ( .A(datapath_1_Instr_21_bF_buf28_), .B(datapath_1_RegisterFile_regfile_mem_10__10_), .C(datapath_1_Instr_22_bF_buf32_), .Y(_2454_) );
OAI22X1 OAI22X1_169 ( .A(_2454_), .B(_2453_), .C(datapath_1_Instr_22_bF_buf31_), .D(_2452_), .Y(_2455_) );
INVX1 INVX1_419 ( .A(datapath_1_RegisterFile_regfile_mem_15__10_), .Y(_2456_) );
AOI21X1 AOI21X1_688 ( .A(_1890__bF_buf26), .B(datapath_1_RegisterFile_regfile_mem_14__10_), .C(_1884__bF_buf1), .Y(_2457_) );
OAI21X1 OAI21X1_1749 ( .A(_1890__bF_buf26), .B(_2456_), .C(_2457_), .Y(_2458_) );
NAND2X1 NAND2X1_1165 ( .A(datapath_1_RegisterFile_regfile_mem_12__10_), .B(_1890__bF_buf26), .Y(_2459_) );
AOI21X1 AOI21X1_689 ( .A(datapath_1_Instr_21_bF_buf27_), .B(datapath_1_RegisterFile_regfile_mem_13__10_), .C(datapath_1_Instr_22_bF_buf30_), .Y(_2460_) );
AOI21X1 AOI21X1_690 ( .A(_2459_), .B(_2460_), .C(_1885__bF_buf0), .Y(_2461_) );
AOI22X1 AOI22X1_144 ( .A(_2458_), .B(_2461_), .C(_1885__bF_buf0), .D(_2455_), .Y(_2462_) );
NOR2X1 NOR2X1_371 ( .A(datapath_1_Instr_21_bF_buf26_), .B(datapath_1_RegisterFile_regfile_mem_0__10_), .Y(_2463_) );
OAI21X1 OAI21X1_1750 ( .A(datapath_1_RegisterFile_regfile_mem_1__10_), .B(_1890__bF_buf44), .C(_1884__bF_buf4), .Y(_2464_) );
NOR2X1 NOR2X1_372 ( .A(datapath_1_RegisterFile_regfile_mem_3__10_), .B(_1890__bF_buf44), .Y(_2465_) );
OAI21X1 OAI21X1_1751 ( .A(datapath_1_Instr_21_bF_buf25_), .B(datapath_1_RegisterFile_regfile_mem_2__10_), .C(datapath_1_Instr_22_bF_buf29_), .Y(_2466_) );
OAI22X1 OAI22X1_170 ( .A(_2465_), .B(_2466_), .C(_2463_), .D(_2464_), .Y(_2467_) );
NOR2X1 NOR2X1_373 ( .A(datapath_1_Instr_23_bF_buf0_), .B(_2467_), .Y(_2468_) );
MUX2X1 MUX2X1_174 ( .A(datapath_1_RegisterFile_regfile_mem_5__10_), .B(datapath_1_RegisterFile_regfile_mem_4__10_), .S(datapath_1_Instr_21_bF_buf24_), .Y(_2469_) );
NOR2X1 NOR2X1_374 ( .A(datapath_1_RegisterFile_regfile_mem_7__10_), .B(_1890__bF_buf44), .Y(_2470_) );
OAI21X1 OAI21X1_1752 ( .A(datapath_1_Instr_21_bF_buf23_), .B(datapath_1_RegisterFile_regfile_mem_6__10_), .C(datapath_1_Instr_22_bF_buf28_), .Y(_2471_) );
OAI22X1 OAI22X1_171 ( .A(_2471_), .B(_2470_), .C(datapath_1_Instr_22_bF_buf27_), .D(_2469_), .Y(_2472_) );
OAI21X1 OAI21X1_1753 ( .A(_1885__bF_buf10), .B(_2472_), .C(_1888__bF_buf0), .Y(_2473_) );
OAI22X1 OAI22X1_172 ( .A(_1888__bF_buf6), .B(_2462_), .C(_2468_), .D(_2473_), .Y(_2474_) );
NAND2X1 NAND2X1_1166 ( .A(_1917__bF_buf3), .B(_2474_), .Y(_2475_) );
AOI22X1 AOI22X1_145 ( .A(_1883__bF_buf0), .B(_1887__bF_buf2), .C(_2451_), .D(_2475_), .Y(datapath_1_RD1_10_) );
NAND2X1 NAND2X1_1167 ( .A(datapath_1_Instr_22_bF_buf26_), .B(datapath_1_RegisterFile_regfile_mem_11__11_), .Y(_2476_) );
NAND2X1 NAND2X1_1168 ( .A(datapath_1_RegisterFile_regfile_mem_9__11_), .B(_1884__bF_buf7), .Y(_2477_) );
NAND3X1 NAND3X1_1467 ( .A(datapath_1_Instr_21_bF_buf22_), .B(_2476_), .C(_2477_), .Y(_2478_) );
NAND2X1 NAND2X1_1169 ( .A(datapath_1_Instr_22_bF_buf25_), .B(datapath_1_RegisterFile_regfile_mem_10__11_), .Y(_2479_) );
AOI21X1 AOI21X1_691 ( .A(_1884__bF_buf7), .B(datapath_1_RegisterFile_regfile_mem_8__11_), .C(datapath_1_Instr_21_bF_buf21_), .Y(_2480_) );
NAND2X1 NAND2X1_1170 ( .A(_2479_), .B(_2480_), .Y(_2481_) );
NAND3X1 NAND3X1_1468 ( .A(_1885__bF_buf8), .B(_2478_), .C(_2481_), .Y(_2482_) );
NAND2X1 NAND2X1_1171 ( .A(datapath_1_Instr_22_bF_buf24_), .B(datapath_1_RegisterFile_regfile_mem_15__11_), .Y(_2483_) );
NAND2X1 NAND2X1_1172 ( .A(datapath_1_RegisterFile_regfile_mem_13__11_), .B(_1884__bF_buf7), .Y(_2484_) );
NAND3X1 NAND3X1_1469 ( .A(datapath_1_Instr_21_bF_buf20_), .B(_2483_), .C(_2484_), .Y(_2485_) );
NAND2X1 NAND2X1_1173 ( .A(datapath_1_Instr_22_bF_buf23_), .B(datapath_1_RegisterFile_regfile_mem_14__11_), .Y(_2486_) );
AOI21X1 AOI21X1_692 ( .A(_1884__bF_buf7), .B(datapath_1_RegisterFile_regfile_mem_12__11_), .C(datapath_1_Instr_21_bF_buf19_), .Y(_2487_) );
NAND2X1 NAND2X1_1174 ( .A(_2486_), .B(_2487_), .Y(_2488_) );
NAND3X1 NAND3X1_1470 ( .A(datapath_1_Instr_23_bF_buf15_bF_buf0_), .B(_2485_), .C(_2488_), .Y(_2489_) );
AOI21X1 AOI21X1_693 ( .A(_2482_), .B(_2489_), .C(_1888__bF_buf4), .Y(_2490_) );
INVX1 INVX1_420 ( .A(datapath_1_RegisterFile_regfile_mem_1__11_), .Y(_2491_) );
AOI21X1 AOI21X1_694 ( .A(datapath_1_Instr_23_bF_buf14_bF_buf0_), .B(datapath_1_RegisterFile_regfile_mem_5__11_), .C(_1890__bF_buf8), .Y(_2492_) );
OAI21X1 OAI21X1_1754 ( .A(datapath_1_Instr_23_bF_buf13_bF_buf0_), .B(_2491_), .C(_2492_), .Y(_2493_) );
INVX1 INVX1_421 ( .A(datapath_1_RegisterFile_regfile_mem_0__11_), .Y(_2494_) );
AOI21X1 AOI21X1_695 ( .A(datapath_1_Instr_23_bF_buf12_bF_buf0_), .B(datapath_1_RegisterFile_regfile_mem_4__11_), .C(datapath_1_Instr_21_bF_buf18_), .Y(_2495_) );
OAI21X1 OAI21X1_1755 ( .A(datapath_1_Instr_23_bF_buf11_bF_buf0_), .B(_2494_), .C(_2495_), .Y(_2496_) );
NAND3X1 NAND3X1_1471 ( .A(_1884__bF_buf6), .B(_2496_), .C(_2493_), .Y(_2497_) );
INVX1 INVX1_422 ( .A(datapath_1_RegisterFile_regfile_mem_3__11_), .Y(_2498_) );
AOI21X1 AOI21X1_696 ( .A(datapath_1_Instr_23_bF_buf10_bF_buf0_), .B(datapath_1_RegisterFile_regfile_mem_7__11_), .C(_1890__bF_buf6), .Y(_2499_) );
OAI21X1 OAI21X1_1756 ( .A(datapath_1_Instr_23_bF_buf9_bF_buf0_), .B(_2498_), .C(_2499_), .Y(_2500_) );
INVX1 INVX1_423 ( .A(datapath_1_RegisterFile_regfile_mem_2__11_), .Y(_2501_) );
AOI21X1 AOI21X1_697 ( .A(datapath_1_Instr_23_bF_buf8_bF_buf0_), .B(datapath_1_RegisterFile_regfile_mem_6__11_), .C(datapath_1_Instr_21_bF_buf17_), .Y(_2502_) );
OAI21X1 OAI21X1_1757 ( .A(datapath_1_Instr_23_bF_buf7_bF_buf0_), .B(_2501_), .C(_2502_), .Y(_2503_) );
NAND3X1 NAND3X1_1472 ( .A(datapath_1_Instr_22_bF_buf22_), .B(_2503_), .C(_2500_), .Y(_2504_) );
AOI21X1 AOI21X1_698 ( .A(_2497_), .B(_2504_), .C(datapath_1_Instr_24_bF_buf4_), .Y(_2505_) );
OAI21X1 OAI21X1_1758 ( .A(_2505_), .B(_2490_), .C(_1917__bF_buf1), .Y(_2506_) );
INVX1 INVX1_424 ( .A(datapath_1_RegisterFile_regfile_mem_19__11_), .Y(_2507_) );
AOI21X1 AOI21X1_699 ( .A(datapath_1_Instr_23_bF_buf6_bF_buf0_), .B(datapath_1_RegisterFile_regfile_mem_23__11_), .C(_1890__bF_buf2), .Y(_2508_) );
OAI21X1 OAI21X1_1759 ( .A(datapath_1_Instr_23_bF_buf5_bF_buf0_), .B(_2507_), .C(_2508_), .Y(_2509_) );
NAND2X1 NAND2X1_1175 ( .A(datapath_1_RegisterFile_regfile_mem_18__11_), .B(_1885__bF_buf3), .Y(_2510_) );
AOI21X1 AOI21X1_700 ( .A(datapath_1_Instr_23_bF_buf4_bF_buf0_), .B(datapath_1_RegisterFile_regfile_mem_22__11_), .C(datapath_1_Instr_21_bF_buf16_), .Y(_2511_) );
AOI21X1 AOI21X1_701 ( .A(_2510_), .B(_2511_), .C(_1884__bF_buf6), .Y(_2512_) );
INVX1 INVX1_425 ( .A(datapath_1_RegisterFile_regfile_mem_17__11_), .Y(_2513_) );
AOI21X1 AOI21X1_702 ( .A(datapath_1_Instr_23_bF_buf3_bF_buf0_), .B(datapath_1_RegisterFile_regfile_mem_21__11_), .C(_1890__bF_buf2), .Y(_2514_) );
OAI21X1 OAI21X1_1760 ( .A(datapath_1_Instr_23_bF_buf2_bF_buf0_), .B(_2513_), .C(_2514_), .Y(_2515_) );
NAND2X1 NAND2X1_1176 ( .A(datapath_1_RegisterFile_regfile_mem_16__11_), .B(_1885__bF_buf7), .Y(_2516_) );
AOI21X1 AOI21X1_703 ( .A(datapath_1_Instr_23_bF_buf1_), .B(datapath_1_RegisterFile_regfile_mem_20__11_), .C(datapath_1_Instr_21_bF_buf15_), .Y(_2517_) );
AOI21X1 AOI21X1_704 ( .A(_2516_), .B(_2517_), .C(datapath_1_Instr_22_bF_buf21_), .Y(_2518_) );
AOI22X1 AOI22X1_146 ( .A(_2512_), .B(_2509_), .C(_2515_), .D(_2518_), .Y(_2519_) );
NOR2X1 NOR2X1_375 ( .A(datapath_1_Instr_21_bF_buf14_), .B(datapath_1_RegisterFile_regfile_mem_24__11_), .Y(_2520_) );
OAI21X1 OAI21X1_1761 ( .A(datapath_1_RegisterFile_regfile_mem_25__11_), .B(_1890__bF_buf19), .C(_1884__bF_buf6), .Y(_2521_) );
NOR2X1 NOR2X1_376 ( .A(datapath_1_RegisterFile_regfile_mem_27__11_), .B(_1890__bF_buf19), .Y(_2522_) );
OAI21X1 OAI21X1_1762 ( .A(datapath_1_Instr_21_bF_buf13_), .B(datapath_1_RegisterFile_regfile_mem_26__11_), .C(datapath_1_Instr_22_bF_buf20_), .Y(_2523_) );
OAI22X1 OAI22X1_173 ( .A(_2522_), .B(_2523_), .C(_2520_), .D(_2521_), .Y(_2524_) );
NOR2X1 NOR2X1_377 ( .A(datapath_1_Instr_23_bF_buf0_), .B(_2524_), .Y(_2525_) );
MUX2X1 MUX2X1_175 ( .A(datapath_1_RegisterFile_regfile_mem_29__11_), .B(datapath_1_RegisterFile_regfile_mem_28__11_), .S(datapath_1_Instr_21_bF_buf12_), .Y(_2526_) );
NOR2X1 NOR2X1_378 ( .A(datapath_1_RegisterFile_regfile_mem_31__11_), .B(_1890__bF_buf17), .Y(_2527_) );
OAI21X1 OAI21X1_1763 ( .A(datapath_1_Instr_21_bF_buf11_), .B(datapath_1_RegisterFile_regfile_mem_30__11_), .C(datapath_1_Instr_22_bF_buf19_), .Y(_2528_) );
OAI22X1 OAI22X1_174 ( .A(_2528_), .B(_2527_), .C(datapath_1_Instr_22_bF_buf18_), .D(_2526_), .Y(_2529_) );
OAI21X1 OAI21X1_1764 ( .A(_1885__bF_buf7), .B(_2529_), .C(datapath_1_Instr_24_bF_buf3_), .Y(_2530_) );
OAI22X1 OAI22X1_175 ( .A(datapath_1_Instr_24_bF_buf2_), .B(_2519_), .C(_2525_), .D(_2530_), .Y(_2531_) );
NAND2X1 NAND2X1_1177 ( .A(datapath_1_Instr_25_bF_buf2_), .B(_2531_), .Y(_2532_) );
AOI22X1 AOI22X1_147 ( .A(_1883__bF_buf3), .B(_1887__bF_buf1), .C(_2506_), .D(_2532_), .Y(datapath_1_RD1_11_) );
NAND2X1 NAND2X1_1178 ( .A(datapath_1_Instr_21_bF_buf10_), .B(datapath_1_RegisterFile_regfile_mem_27__12_), .Y(_2533_) );
NAND2X1 NAND2X1_1179 ( .A(datapath_1_RegisterFile_regfile_mem_26__12_), .B(_1890__bF_buf6), .Y(_2534_) );
NAND3X1 NAND3X1_1473 ( .A(datapath_1_Instr_22_bF_buf17_), .B(_2533_), .C(_2534_), .Y(_2535_) );
NAND2X1 NAND2X1_1180 ( .A(datapath_1_Instr_21_bF_buf9_), .B(datapath_1_RegisterFile_regfile_mem_25__12_), .Y(_2536_) );
AOI21X1 AOI21X1_705 ( .A(_1890__bF_buf6), .B(datapath_1_RegisterFile_regfile_mem_24__12_), .C(datapath_1_Instr_22_bF_buf16_), .Y(_2537_) );
NAND2X1 NAND2X1_1181 ( .A(_2536_), .B(_2537_), .Y(_2538_) );
NAND3X1 NAND3X1_1474 ( .A(_1885__bF_buf10), .B(_2535_), .C(_2538_), .Y(_2539_) );
NAND2X1 NAND2X1_1182 ( .A(datapath_1_Instr_21_bF_buf8_), .B(datapath_1_RegisterFile_regfile_mem_31__12_), .Y(_2540_) );
AOI21X1 AOI21X1_706 ( .A(_1890__bF_buf44), .B(datapath_1_RegisterFile_regfile_mem_30__12_), .C(_1884__bF_buf4), .Y(_2541_) );
NAND2X1 NAND2X1_1183 ( .A(_2540_), .B(_2541_), .Y(_2542_) );
INVX1 INVX1_426 ( .A(datapath_1_RegisterFile_regfile_mem_28__12_), .Y(_2543_) );
AOI21X1 AOI21X1_707 ( .A(datapath_1_Instr_21_bF_buf7_), .B(datapath_1_RegisterFile_regfile_mem_29__12_), .C(datapath_1_Instr_22_bF_buf15_), .Y(_2544_) );
OAI21X1 OAI21X1_1765 ( .A(datapath_1_Instr_21_bF_buf6_), .B(_2543_), .C(_2544_), .Y(_2545_) );
NAND3X1 NAND3X1_1475 ( .A(datapath_1_Instr_23_bF_buf15_bF_buf3_), .B(_2545_), .C(_2542_), .Y(_2546_) );
AOI21X1 AOI21X1_708 ( .A(_2539_), .B(_2546_), .C(_1888__bF_buf0), .Y(_2547_) );
MUX2X1 MUX2X1_176 ( .A(datapath_1_RegisterFile_regfile_mem_18__12_), .B(datapath_1_RegisterFile_regfile_mem_16__12_), .S(datapath_1_Instr_22_bF_buf14_), .Y(_2548_) );
NAND2X1 NAND2X1_1184 ( .A(_1890__bF_buf6), .B(_2548_), .Y(_2549_) );
MUX2X1 MUX2X1_177 ( .A(datapath_1_RegisterFile_regfile_mem_19__12_), .B(datapath_1_RegisterFile_regfile_mem_17__12_), .S(datapath_1_Instr_22_bF_buf13_), .Y(_2550_) );
NAND2X1 NAND2X1_1185 ( .A(datapath_1_Instr_21_bF_buf5_), .B(_2550_), .Y(_2551_) );
NAND3X1 NAND3X1_1476 ( .A(_1885__bF_buf10), .B(_2549_), .C(_2551_), .Y(_2552_) );
MUX2X1 MUX2X1_178 ( .A(datapath_1_RegisterFile_regfile_mem_22__12_), .B(datapath_1_RegisterFile_regfile_mem_20__12_), .S(datapath_1_Instr_22_bF_buf12_), .Y(_2553_) );
NAND2X1 NAND2X1_1186 ( .A(_1890__bF_buf32), .B(_2553_), .Y(_2554_) );
MUX2X1 MUX2X1_179 ( .A(datapath_1_RegisterFile_regfile_mem_23__12_), .B(datapath_1_RegisterFile_regfile_mem_21__12_), .S(datapath_1_Instr_22_bF_buf11_), .Y(_2555_) );
NAND2X1 NAND2X1_1187 ( .A(datapath_1_Instr_21_bF_buf4_), .B(_2555_), .Y(_2556_) );
NAND3X1 NAND3X1_1477 ( .A(datapath_1_Instr_23_bF_buf14_bF_buf3_), .B(_2554_), .C(_2556_), .Y(_2557_) );
AOI21X1 AOI21X1_709 ( .A(_2552_), .B(_2557_), .C(datapath_1_Instr_24_bF_buf1_), .Y(_2558_) );
OAI21X1 OAI21X1_1766 ( .A(_2558_), .B(_2547_), .C(datapath_1_Instr_25_bF_buf1_), .Y(_2559_) );
MUX2X1 MUX2X1_180 ( .A(datapath_1_RegisterFile_regfile_mem_9__12_), .B(datapath_1_RegisterFile_regfile_mem_8__12_), .S(datapath_1_Instr_21_bF_buf3_), .Y(_2560_) );
NOR2X1 NOR2X1_379 ( .A(datapath_1_RegisterFile_regfile_mem_11__12_), .B(_1890__bF_buf41), .Y(_2561_) );
OAI21X1 OAI21X1_1767 ( .A(datapath_1_Instr_21_bF_buf2_), .B(datapath_1_RegisterFile_regfile_mem_10__12_), .C(datapath_1_Instr_22_bF_buf10_), .Y(_2562_) );
OAI22X1 OAI22X1_176 ( .A(_2562_), .B(_2561_), .C(datapath_1_Instr_22_bF_buf9_), .D(_2560_), .Y(_2563_) );
INVX1 INVX1_427 ( .A(datapath_1_RegisterFile_regfile_mem_15__12_), .Y(_2564_) );
AOI21X1 AOI21X1_710 ( .A(_1890__bF_buf21), .B(datapath_1_RegisterFile_regfile_mem_14__12_), .C(_1884__bF_buf1), .Y(_2565_) );
OAI21X1 OAI21X1_1768 ( .A(_1890__bF_buf21), .B(_2564_), .C(_2565_), .Y(_2566_) );
NAND2X1 NAND2X1_1188 ( .A(datapath_1_RegisterFile_regfile_mem_12__12_), .B(_1890__bF_buf21), .Y(_2567_) );
AOI21X1 AOI21X1_711 ( .A(datapath_1_Instr_21_bF_buf1_), .B(datapath_1_RegisterFile_regfile_mem_13__12_), .C(datapath_1_Instr_22_bF_buf8_), .Y(_2568_) );
AOI21X1 AOI21X1_712 ( .A(_2567_), .B(_2568_), .C(_1885__bF_buf0), .Y(_2569_) );
AOI22X1 AOI22X1_148 ( .A(_2566_), .B(_2569_), .C(_1885__bF_buf0), .D(_2563_), .Y(_2570_) );
NOR2X1 NOR2X1_380 ( .A(datapath_1_Instr_21_bF_buf0_), .B(datapath_1_RegisterFile_regfile_mem_0__12_), .Y(_2571_) );
OAI21X1 OAI21X1_1769 ( .A(datapath_1_RegisterFile_regfile_mem_1__12_), .B(_1890__bF_buf12), .C(_1884__bF_buf8), .Y(_2572_) );
NOR2X1 NOR2X1_381 ( .A(datapath_1_RegisterFile_regfile_mem_3__12_), .B(_1890__bF_buf12), .Y(_2573_) );
OAI21X1 OAI21X1_1770 ( .A(datapath_1_Instr_21_bF_buf55_), .B(datapath_1_RegisterFile_regfile_mem_2__12_), .C(datapath_1_Instr_22_bF_buf7_), .Y(_2574_) );
OAI22X1 OAI22X1_177 ( .A(_2573_), .B(_2574_), .C(_2571_), .D(_2572_), .Y(_2575_) );
NOR2X1 NOR2X1_382 ( .A(datapath_1_Instr_23_bF_buf13_bF_buf3_), .B(_2575_), .Y(_2576_) );
MUX2X1 MUX2X1_181 ( .A(datapath_1_RegisterFile_regfile_mem_5__12_), .B(datapath_1_RegisterFile_regfile_mem_4__12_), .S(datapath_1_Instr_21_bF_buf54_), .Y(_2577_) );
NOR2X1 NOR2X1_383 ( .A(datapath_1_RegisterFile_regfile_mem_7__12_), .B(_1890__bF_buf41), .Y(_2578_) );
OAI21X1 OAI21X1_1771 ( .A(datapath_1_Instr_21_bF_buf53_), .B(datapath_1_RegisterFile_regfile_mem_6__12_), .C(datapath_1_Instr_22_bF_buf6_), .Y(_2579_) );
OAI22X1 OAI22X1_178 ( .A(_2579_), .B(_2578_), .C(datapath_1_Instr_22_bF_buf5_), .D(_2577_), .Y(_2580_) );
OAI21X1 OAI21X1_1772 ( .A(_1885__bF_buf0), .B(_2580_), .C(_1888__bF_buf7), .Y(_2581_) );
OAI22X1 OAI22X1_179 ( .A(_1888__bF_buf7), .B(_2570_), .C(_2576_), .D(_2581_), .Y(_2582_) );
NAND2X1 NAND2X1_1189 ( .A(_1917__bF_buf3), .B(_2582_), .Y(_2583_) );
AOI22X1 AOI22X1_149 ( .A(_1883__bF_buf1), .B(_1887__bF_buf0), .C(_2559_), .D(_2583_), .Y(datapath_1_RD1_12_) );
NAND2X1 NAND2X1_1190 ( .A(datapath_1_Instr_21_bF_buf52_), .B(datapath_1_RegisterFile_regfile_mem_27__13_), .Y(_2584_) );
NAND2X1 NAND2X1_1191 ( .A(datapath_1_RegisterFile_regfile_mem_26__13_), .B(_1890__bF_buf37), .Y(_2585_) );
NAND3X1 NAND3X1_1478 ( .A(datapath_1_Instr_22_bF_buf4_), .B(_2584_), .C(_2585_), .Y(_2586_) );
NAND2X1 NAND2X1_1192 ( .A(datapath_1_Instr_21_bF_buf51_), .B(datapath_1_RegisterFile_regfile_mem_25__13_), .Y(_2587_) );
AOI21X1 AOI21X1_713 ( .A(_1890__bF_buf37), .B(datapath_1_RegisterFile_regfile_mem_24__13_), .C(datapath_1_Instr_22_bF_buf3_), .Y(_2588_) );
NAND2X1 NAND2X1_1193 ( .A(_2587_), .B(_2588_), .Y(_2589_) );
NAND3X1 NAND3X1_1479 ( .A(_1885__bF_buf9), .B(_2586_), .C(_2589_), .Y(_2590_) );
NAND2X1 NAND2X1_1194 ( .A(datapath_1_Instr_21_bF_buf50_), .B(datapath_1_RegisterFile_regfile_mem_31__13_), .Y(_2591_) );
AOI21X1 AOI21X1_714 ( .A(_1890__bF_buf9), .B(datapath_1_RegisterFile_regfile_mem_30__13_), .C(_1884__bF_buf9), .Y(_2592_) );
NAND2X1 NAND2X1_1195 ( .A(_2591_), .B(_2592_), .Y(_2593_) );
INVX1 INVX1_428 ( .A(datapath_1_RegisterFile_regfile_mem_28__13_), .Y(_2594_) );
AOI21X1 AOI21X1_715 ( .A(datapath_1_Instr_21_bF_buf49_), .B(datapath_1_RegisterFile_regfile_mem_29__13_), .C(datapath_1_Instr_22_bF_buf2_), .Y(_2595_) );
OAI21X1 OAI21X1_1773 ( .A(datapath_1_Instr_21_bF_buf48_), .B(_2594_), .C(_2595_), .Y(_2596_) );
NAND3X1 NAND3X1_1480 ( .A(datapath_1_Instr_23_bF_buf12_bF_buf3_), .B(_2596_), .C(_2593_), .Y(_2597_) );
AOI21X1 AOI21X1_716 ( .A(_2590_), .B(_2597_), .C(_1888__bF_buf1), .Y(_2598_) );
MUX2X1 MUX2X1_182 ( .A(datapath_1_RegisterFile_regfile_mem_18__13_), .B(datapath_1_RegisterFile_regfile_mem_16__13_), .S(datapath_1_Instr_22_bF_buf1_), .Y(_2599_) );
NAND2X1 NAND2X1_1196 ( .A(_1890__bF_buf24), .B(_2599_), .Y(_2600_) );
MUX2X1 MUX2X1_183 ( .A(datapath_1_RegisterFile_regfile_mem_19__13_), .B(datapath_1_RegisterFile_regfile_mem_17__13_), .S(datapath_1_Instr_22_bF_buf0_), .Y(_2601_) );
NAND2X1 NAND2X1_1197 ( .A(datapath_1_Instr_21_bF_buf47_), .B(_2601_), .Y(_2602_) );
NAND3X1 NAND3X1_1481 ( .A(_1885__bF_buf9), .B(_2600_), .C(_2602_), .Y(_2603_) );
MUX2X1 MUX2X1_184 ( .A(datapath_1_RegisterFile_regfile_mem_22__13_), .B(datapath_1_RegisterFile_regfile_mem_20__13_), .S(datapath_1_Instr_22_bF_buf50_), .Y(_2604_) );
NAND2X1 NAND2X1_1198 ( .A(_1890__bF_buf24), .B(_2604_), .Y(_2605_) );
MUX2X1 MUX2X1_185 ( .A(datapath_1_RegisterFile_regfile_mem_23__13_), .B(datapath_1_RegisterFile_regfile_mem_21__13_), .S(datapath_1_Instr_22_bF_buf49_), .Y(_2606_) );
NAND2X1 NAND2X1_1199 ( .A(datapath_1_Instr_21_bF_buf46_), .B(_2606_), .Y(_2607_) );
NAND3X1 NAND3X1_1482 ( .A(datapath_1_Instr_23_bF_buf11_bF_buf3_), .B(_2605_), .C(_2607_), .Y(_2608_) );
AOI21X1 AOI21X1_717 ( .A(_2603_), .B(_2608_), .C(datapath_1_Instr_24_bF_buf0_), .Y(_2609_) );
OAI21X1 OAI21X1_1774 ( .A(_2609_), .B(_2598_), .C(datapath_1_Instr_25_bF_buf0_), .Y(_2610_) );
MUX2X1 MUX2X1_186 ( .A(datapath_1_RegisterFile_regfile_mem_9__13_), .B(datapath_1_RegisterFile_regfile_mem_8__13_), .S(datapath_1_Instr_21_bF_buf45_), .Y(_2611_) );
NOR2X1 NOR2X1_384 ( .A(datapath_1_RegisterFile_regfile_mem_11__13_), .B(_1890__bF_buf15), .Y(_2612_) );
OAI21X1 OAI21X1_1775 ( .A(datapath_1_Instr_21_bF_buf44_), .B(datapath_1_RegisterFile_regfile_mem_10__13_), .C(datapath_1_Instr_22_bF_buf48_), .Y(_2613_) );
OAI22X1 OAI22X1_180 ( .A(_2613_), .B(_2612_), .C(datapath_1_Instr_22_bF_buf47_), .D(_2611_), .Y(_2614_) );
INVX1 INVX1_429 ( .A(datapath_1_RegisterFile_regfile_mem_15__13_), .Y(_2615_) );
AOI21X1 AOI21X1_718 ( .A(_1890__bF_buf15), .B(datapath_1_RegisterFile_regfile_mem_14__13_), .C(_1884__bF_buf5), .Y(_2616_) );
OAI21X1 OAI21X1_1776 ( .A(_1890__bF_buf15), .B(_2615_), .C(_2616_), .Y(_2617_) );
NAND2X1 NAND2X1_1200 ( .A(datapath_1_RegisterFile_regfile_mem_12__13_), .B(_1890__bF_buf46), .Y(_2618_) );
AOI21X1 AOI21X1_719 ( .A(datapath_1_Instr_21_bF_buf43_), .B(datapath_1_RegisterFile_regfile_mem_13__13_), .C(datapath_1_Instr_22_bF_buf46_), .Y(_2619_) );
AOI21X1 AOI21X1_720 ( .A(_2618_), .B(_2619_), .C(_1885__bF_buf1), .Y(_2620_) );
AOI22X1 AOI22X1_150 ( .A(_2617_), .B(_2620_), .C(_1885__bF_buf1), .D(_2614_), .Y(_2621_) );
NOR2X1 NOR2X1_385 ( .A(datapath_1_Instr_21_bF_buf42_), .B(datapath_1_RegisterFile_regfile_mem_0__13_), .Y(_2622_) );
OAI21X1 OAI21X1_1777 ( .A(datapath_1_RegisterFile_regfile_mem_1__13_), .B(_1890__bF_buf33), .C(_1884__bF_buf3), .Y(_2623_) );
NOR2X1 NOR2X1_386 ( .A(datapath_1_RegisterFile_regfile_mem_3__13_), .B(_1890__bF_buf33), .Y(_2624_) );
OAI21X1 OAI21X1_1778 ( .A(datapath_1_Instr_21_bF_buf41_), .B(datapath_1_RegisterFile_regfile_mem_2__13_), .C(datapath_1_Instr_22_bF_buf45_), .Y(_2625_) );
OAI22X1 OAI22X1_181 ( .A(_2624_), .B(_2625_), .C(_2622_), .D(_2623_), .Y(_2626_) );
NOR2X1 NOR2X1_387 ( .A(datapath_1_Instr_23_bF_buf10_bF_buf3_), .B(_2626_), .Y(_2627_) );
MUX2X1 MUX2X1_187 ( .A(datapath_1_RegisterFile_regfile_mem_5__13_), .B(datapath_1_RegisterFile_regfile_mem_4__13_), .S(datapath_1_Instr_21_bF_buf40_), .Y(_2628_) );
NOR2X1 NOR2X1_388 ( .A(datapath_1_RegisterFile_regfile_mem_7__13_), .B(_1890__bF_buf33), .Y(_2629_) );
OAI21X1 OAI21X1_1779 ( .A(datapath_1_Instr_21_bF_buf39_), .B(datapath_1_RegisterFile_regfile_mem_6__13_), .C(datapath_1_Instr_22_bF_buf44_), .Y(_2630_) );
OAI22X1 OAI22X1_182 ( .A(_2630_), .B(_2629_), .C(datapath_1_Instr_22_bF_buf43_), .D(_2628_), .Y(_2631_) );
OAI21X1 OAI21X1_1780 ( .A(_1885__bF_buf1), .B(_2631_), .C(_1888__bF_buf2), .Y(_2632_) );
OAI22X1 OAI22X1_183 ( .A(_1888__bF_buf2), .B(_2621_), .C(_2627_), .D(_2632_), .Y(_2633_) );
NAND2X1 NAND2X1_1201 ( .A(_1917__bF_buf4), .B(_2633_), .Y(_2634_) );
AOI22X1 AOI22X1_151 ( .A(_1883__bF_buf4), .B(_1887__bF_buf3), .C(_2610_), .D(_2634_), .Y(datapath_1_RD1_13_) );
NAND2X1 NAND2X1_1202 ( .A(datapath_1_Instr_21_bF_buf38_), .B(datapath_1_RegisterFile_regfile_mem_27__14_), .Y(_2635_) );
NAND2X1 NAND2X1_1203 ( .A(datapath_1_RegisterFile_regfile_mem_26__14_), .B(_1890__bF_buf22), .Y(_2636_) );
NAND3X1 NAND3X1_1483 ( .A(datapath_1_Instr_22_bF_buf42_), .B(_2635_), .C(_2636_), .Y(_2637_) );
NAND2X1 NAND2X1_1204 ( .A(datapath_1_Instr_21_bF_buf37_), .B(datapath_1_RegisterFile_regfile_mem_25__14_), .Y(_2638_) );
AOI21X1 AOI21X1_721 ( .A(_1890__bF_buf22), .B(datapath_1_RegisterFile_regfile_mem_24__14_), .C(datapath_1_Instr_22_bF_buf41_), .Y(_2639_) );
NAND2X1 NAND2X1_1205 ( .A(_2638_), .B(_2639_), .Y(_2640_) );
NAND3X1 NAND3X1_1484 ( .A(_1885__bF_buf6), .B(_2637_), .C(_2640_), .Y(_2641_) );
NAND2X1 NAND2X1_1206 ( .A(datapath_1_Instr_21_bF_buf36_), .B(datapath_1_RegisterFile_regfile_mem_31__14_), .Y(_2642_) );
AOI21X1 AOI21X1_722 ( .A(_1890__bF_buf34), .B(datapath_1_RegisterFile_regfile_mem_30__14_), .C(_1884__bF_buf3), .Y(_2643_) );
NAND2X1 NAND2X1_1207 ( .A(_2642_), .B(_2643_), .Y(_2644_) );
INVX1 INVX1_430 ( .A(datapath_1_RegisterFile_regfile_mem_28__14_), .Y(_2645_) );
AOI21X1 AOI21X1_723 ( .A(datapath_1_Instr_21_bF_buf35_), .B(datapath_1_RegisterFile_regfile_mem_29__14_), .C(datapath_1_Instr_22_bF_buf40_), .Y(_2646_) );
OAI21X1 OAI21X1_1781 ( .A(datapath_1_Instr_21_bF_buf34_), .B(_2645_), .C(_2646_), .Y(_2647_) );
NAND3X1 NAND3X1_1485 ( .A(datapath_1_Instr_23_bF_buf9_bF_buf3_), .B(_2647_), .C(_2644_), .Y(_2648_) );
AOI21X1 AOI21X1_724 ( .A(_2641_), .B(_2648_), .C(_1888__bF_buf1), .Y(_2649_) );
MUX2X1 MUX2X1_188 ( .A(datapath_1_RegisterFile_regfile_mem_18__14_), .B(datapath_1_RegisterFile_regfile_mem_16__14_), .S(datapath_1_Instr_22_bF_buf39_), .Y(_2650_) );
NAND2X1 NAND2X1_1208 ( .A(_1890__bF_buf22), .B(_2650_), .Y(_2651_) );
MUX2X1 MUX2X1_189 ( .A(datapath_1_RegisterFile_regfile_mem_19__14_), .B(datapath_1_RegisterFile_regfile_mem_17__14_), .S(datapath_1_Instr_22_bF_buf38_), .Y(_2652_) );
NAND2X1 NAND2X1_1209 ( .A(datapath_1_Instr_21_bF_buf33_), .B(_2652_), .Y(_2653_) );
NAND3X1 NAND3X1_1486 ( .A(_1885__bF_buf6), .B(_2651_), .C(_2653_), .Y(_2654_) );
MUX2X1 MUX2X1_190 ( .A(datapath_1_RegisterFile_regfile_mem_22__14_), .B(datapath_1_RegisterFile_regfile_mem_20__14_), .S(datapath_1_Instr_22_bF_buf37_), .Y(_2655_) );
NAND2X1 NAND2X1_1210 ( .A(_1890__bF_buf39), .B(_2655_), .Y(_2656_) );
MUX2X1 MUX2X1_191 ( .A(datapath_1_RegisterFile_regfile_mem_23__14_), .B(datapath_1_RegisterFile_regfile_mem_21__14_), .S(datapath_1_Instr_22_bF_buf36_), .Y(_2657_) );
NAND2X1 NAND2X1_1211 ( .A(datapath_1_Instr_21_bF_buf32_), .B(_2657_), .Y(_2658_) );
NAND3X1 NAND3X1_1487 ( .A(datapath_1_Instr_23_bF_buf8_bF_buf3_), .B(_2656_), .C(_2658_), .Y(_2659_) );
AOI21X1 AOI21X1_725 ( .A(_2654_), .B(_2659_), .C(datapath_1_Instr_24_bF_buf6_), .Y(_2660_) );
OAI21X1 OAI21X1_1782 ( .A(_2660_), .B(_2649_), .C(datapath_1_Instr_25_bF_buf5_), .Y(_2661_) );
MUX2X1 MUX2X1_192 ( .A(datapath_1_RegisterFile_regfile_mem_9__14_), .B(datapath_1_RegisterFile_regfile_mem_8__14_), .S(datapath_1_Instr_21_bF_buf31_), .Y(_2662_) );
NOR2X1 NOR2X1_389 ( .A(datapath_1_RegisterFile_regfile_mem_11__14_), .B(_1890__bF_buf45), .Y(_2663_) );
OAI21X1 OAI21X1_1783 ( .A(datapath_1_Instr_21_bF_buf30_), .B(datapath_1_RegisterFile_regfile_mem_10__14_), .C(datapath_1_Instr_22_bF_buf35_), .Y(_2664_) );
OAI22X1 OAI22X1_184 ( .A(_2664_), .B(_2663_), .C(datapath_1_Instr_22_bF_buf34_), .D(_2662_), .Y(_2665_) );
INVX1 INVX1_431 ( .A(datapath_1_RegisterFile_regfile_mem_15__14_), .Y(_2666_) );
AOI21X1 AOI21X1_726 ( .A(_1890__bF_buf45), .B(datapath_1_RegisterFile_regfile_mem_14__14_), .C(_1884__bF_buf1), .Y(_2667_) );
OAI21X1 OAI21X1_1784 ( .A(_1890__bF_buf45), .B(_2666_), .C(_2667_), .Y(_2668_) );
NAND2X1 NAND2X1_1212 ( .A(datapath_1_RegisterFile_regfile_mem_12__14_), .B(_1890__bF_buf45), .Y(_2669_) );
AOI21X1 AOI21X1_727 ( .A(datapath_1_Instr_21_bF_buf29_), .B(datapath_1_RegisterFile_regfile_mem_13__14_), .C(datapath_1_Instr_22_bF_buf33_), .Y(_2670_) );
AOI21X1 AOI21X1_728 ( .A(_2669_), .B(_2670_), .C(_1885__bF_buf5), .Y(_2671_) );
AOI22X1 AOI22X1_152 ( .A(_2668_), .B(_2671_), .C(_1885__bF_buf5), .D(_2665_), .Y(_2672_) );
NOR2X1 NOR2X1_390 ( .A(datapath_1_Instr_21_bF_buf28_), .B(datapath_1_RegisterFile_regfile_mem_0__14_), .Y(_2673_) );
OAI21X1 OAI21X1_1785 ( .A(datapath_1_RegisterFile_regfile_mem_1__14_), .B(_1890__bF_buf45), .C(_1884__bF_buf1), .Y(_2674_) );
NOR2X1 NOR2X1_391 ( .A(datapath_1_RegisterFile_regfile_mem_3__14_), .B(_1890__bF_buf14), .Y(_2675_) );
OAI21X1 OAI21X1_1786 ( .A(datapath_1_Instr_21_bF_buf27_), .B(datapath_1_RegisterFile_regfile_mem_2__14_), .C(datapath_1_Instr_22_bF_buf32_), .Y(_2676_) );
OAI22X1 OAI22X1_185 ( .A(_2675_), .B(_2676_), .C(_2673_), .D(_2674_), .Y(_2677_) );
NOR2X1 NOR2X1_392 ( .A(datapath_1_Instr_23_bF_buf7_bF_buf3_), .B(_2677_), .Y(_2678_) );
MUX2X1 MUX2X1_193 ( .A(datapath_1_RegisterFile_regfile_mem_5__14_), .B(datapath_1_RegisterFile_regfile_mem_4__14_), .S(datapath_1_Instr_21_bF_buf26_), .Y(_2679_) );
NOR2X1 NOR2X1_393 ( .A(datapath_1_RegisterFile_regfile_mem_7__14_), .B(_1890__bF_buf45), .Y(_2680_) );
OAI21X1 OAI21X1_1787 ( .A(datapath_1_Instr_21_bF_buf25_), .B(datapath_1_RegisterFile_regfile_mem_6__14_), .C(datapath_1_Instr_22_bF_buf31_), .Y(_2681_) );
OAI22X1 OAI22X1_186 ( .A(_2681_), .B(_2680_), .C(datapath_1_Instr_22_bF_buf30_), .D(_2679_), .Y(_2682_) );
OAI21X1 OAI21X1_1788 ( .A(_1885__bF_buf5), .B(_2682_), .C(_1888__bF_buf5), .Y(_2683_) );
OAI22X1 OAI22X1_187 ( .A(_1888__bF_buf5), .B(_2672_), .C(_2678_), .D(_2683_), .Y(_2684_) );
NAND2X1 NAND2X1_1213 ( .A(_1917__bF_buf0), .B(_2684_), .Y(_2685_) );
AOI22X1 AOI22X1_153 ( .A(_1883__bF_buf4), .B(_1887__bF_buf3), .C(_2661_), .D(_2685_), .Y(datapath_1_RD1_14_) );
NAND2X1 NAND2X1_1214 ( .A(datapath_1_Instr_21_bF_buf24_), .B(datapath_1_RegisterFile_regfile_mem_27__15_), .Y(_2686_) );
NAND2X1 NAND2X1_1215 ( .A(datapath_1_RegisterFile_regfile_mem_26__15_), .B(_1890__bF_buf6), .Y(_2687_) );
NAND3X1 NAND3X1_1488 ( .A(datapath_1_Instr_22_bF_buf29_), .B(_2686_), .C(_2687_), .Y(_2688_) );
NAND2X1 NAND2X1_1216 ( .A(datapath_1_Instr_21_bF_buf23_), .B(datapath_1_RegisterFile_regfile_mem_25__15_), .Y(_2689_) );
AOI21X1 AOI21X1_729 ( .A(_1890__bF_buf6), .B(datapath_1_RegisterFile_regfile_mem_24__15_), .C(datapath_1_Instr_22_bF_buf28_), .Y(_2690_) );
NAND2X1 NAND2X1_1217 ( .A(_2689_), .B(_2690_), .Y(_2691_) );
NAND3X1 NAND3X1_1489 ( .A(_1885__bF_buf10), .B(_2688_), .C(_2691_), .Y(_2692_) );
NAND2X1 NAND2X1_1218 ( .A(datapath_1_Instr_21_bF_buf22_), .B(datapath_1_RegisterFile_regfile_mem_31__15_), .Y(_2693_) );
AOI21X1 AOI21X1_730 ( .A(_1890__bF_buf2), .B(datapath_1_RegisterFile_regfile_mem_30__15_), .C(_1884__bF_buf6), .Y(_2694_) );
NAND2X1 NAND2X1_1219 ( .A(_2693_), .B(_2694_), .Y(_2695_) );
INVX1 INVX1_432 ( .A(datapath_1_RegisterFile_regfile_mem_28__15_), .Y(_2696_) );
AOI21X1 AOI21X1_731 ( .A(datapath_1_Instr_21_bF_buf21_), .B(datapath_1_RegisterFile_regfile_mem_29__15_), .C(datapath_1_Instr_22_bF_buf27_), .Y(_2697_) );
OAI21X1 OAI21X1_1789 ( .A(datapath_1_Instr_21_bF_buf20_), .B(_2696_), .C(_2697_), .Y(_2698_) );
NAND3X1 NAND3X1_1490 ( .A(datapath_1_Instr_23_bF_buf6_bF_buf3_), .B(_2698_), .C(_2695_), .Y(_2699_) );
AOI21X1 AOI21X1_732 ( .A(_2692_), .B(_2699_), .C(_1888__bF_buf3), .Y(_2700_) );
MUX2X1 MUX2X1_194 ( .A(datapath_1_RegisterFile_regfile_mem_18__15_), .B(datapath_1_RegisterFile_regfile_mem_16__15_), .S(datapath_1_Instr_22_bF_buf26_), .Y(_2701_) );
NAND2X1 NAND2X1_1220 ( .A(_1890__bF_buf43), .B(_2701_), .Y(_2702_) );
MUX2X1 MUX2X1_195 ( .A(datapath_1_RegisterFile_regfile_mem_19__15_), .B(datapath_1_RegisterFile_regfile_mem_17__15_), .S(datapath_1_Instr_22_bF_buf25_), .Y(_2703_) );
NAND2X1 NAND2X1_1221 ( .A(datapath_1_Instr_21_bF_buf19_), .B(_2703_), .Y(_2704_) );
NAND3X1 NAND3X1_1491 ( .A(_1885__bF_buf3), .B(_2702_), .C(_2704_), .Y(_2705_) );
MUX2X1 MUX2X1_196 ( .A(datapath_1_RegisterFile_regfile_mem_22__15_), .B(datapath_1_RegisterFile_regfile_mem_20__15_), .S(datapath_1_Instr_22_bF_buf24_), .Y(_2706_) );
NAND2X1 NAND2X1_1222 ( .A(_1890__bF_buf19), .B(_2706_), .Y(_2707_) );
MUX2X1 MUX2X1_197 ( .A(datapath_1_RegisterFile_regfile_mem_23__15_), .B(datapath_1_RegisterFile_regfile_mem_21__15_), .S(datapath_1_Instr_22_bF_buf23_), .Y(_2708_) );
NAND2X1 NAND2X1_1223 ( .A(datapath_1_Instr_21_bF_buf18_), .B(_2708_), .Y(_2709_) );
NAND3X1 NAND3X1_1492 ( .A(datapath_1_Instr_23_bF_buf5_bF_buf3_), .B(_2707_), .C(_2709_), .Y(_2710_) );
AOI21X1 AOI21X1_733 ( .A(_2705_), .B(_2710_), .C(datapath_1_Instr_24_bF_buf5_), .Y(_2711_) );
OAI21X1 OAI21X1_1790 ( .A(_2711_), .B(_2700_), .C(datapath_1_Instr_25_bF_buf4_), .Y(_2712_) );
MUX2X1 MUX2X1_198 ( .A(datapath_1_RegisterFile_regfile_mem_9__15_), .B(datapath_1_RegisterFile_regfile_mem_8__15_), .S(datapath_1_Instr_21_bF_buf17_), .Y(_2713_) );
NOR2X1 NOR2X1_394 ( .A(datapath_1_RegisterFile_regfile_mem_11__15_), .B(_1890__bF_buf42), .Y(_2714_) );
OAI21X1 OAI21X1_1791 ( .A(datapath_1_Instr_21_bF_buf16_), .B(datapath_1_RegisterFile_regfile_mem_10__15_), .C(datapath_1_Instr_22_bF_buf22_), .Y(_2715_) );
OAI22X1 OAI22X1_188 ( .A(_2715_), .B(_2714_), .C(datapath_1_Instr_22_bF_buf21_), .D(_2713_), .Y(_2716_) );
INVX1 INVX1_433 ( .A(datapath_1_RegisterFile_regfile_mem_15__15_), .Y(_2717_) );
AOI21X1 AOI21X1_734 ( .A(_1890__bF_buf23), .B(datapath_1_RegisterFile_regfile_mem_14__15_), .C(_1884__bF_buf7), .Y(_2718_) );
OAI21X1 OAI21X1_1792 ( .A(_1890__bF_buf23), .B(_2717_), .C(_2718_), .Y(_2719_) );
NAND2X1 NAND2X1_1224 ( .A(datapath_1_RegisterFile_regfile_mem_12__15_), .B(_1890__bF_buf42), .Y(_2720_) );
AOI21X1 AOI21X1_735 ( .A(datapath_1_Instr_21_bF_buf15_), .B(datapath_1_RegisterFile_regfile_mem_13__15_), .C(datapath_1_Instr_22_bF_buf20_), .Y(_2721_) );
AOI21X1 AOI21X1_736 ( .A(_2720_), .B(_2721_), .C(_1885__bF_buf8), .Y(_2722_) );
AOI22X1 AOI22X1_154 ( .A(_2719_), .B(_2722_), .C(_1885__bF_buf8), .D(_2716_), .Y(_2723_) );
NOR2X1 NOR2X1_395 ( .A(datapath_1_Instr_21_bF_buf14_), .B(datapath_1_RegisterFile_regfile_mem_0__15_), .Y(_2724_) );
OAI21X1 OAI21X1_1793 ( .A(datapath_1_RegisterFile_regfile_mem_1__15_), .B(_1890__bF_buf0), .C(_1884__bF_buf7), .Y(_2725_) );
NOR2X1 NOR2X1_396 ( .A(datapath_1_RegisterFile_regfile_mem_3__15_), .B(_1890__bF_buf0), .Y(_2726_) );
OAI21X1 OAI21X1_1794 ( .A(datapath_1_Instr_21_bF_buf13_), .B(datapath_1_RegisterFile_regfile_mem_2__15_), .C(datapath_1_Instr_22_bF_buf19_), .Y(_2727_) );
OAI22X1 OAI22X1_189 ( .A(_2726_), .B(_2727_), .C(_2724_), .D(_2725_), .Y(_2728_) );
NOR2X1 NOR2X1_397 ( .A(datapath_1_Instr_23_bF_buf4_bF_buf3_), .B(_2728_), .Y(_2729_) );
MUX2X1 MUX2X1_199 ( .A(datapath_1_RegisterFile_regfile_mem_5__15_), .B(datapath_1_RegisterFile_regfile_mem_4__15_), .S(datapath_1_Instr_21_bF_buf12_), .Y(_2730_) );
NOR2X1 NOR2X1_398 ( .A(datapath_1_RegisterFile_regfile_mem_7__15_), .B(_1890__bF_buf29), .Y(_2731_) );
OAI21X1 OAI21X1_1795 ( .A(datapath_1_Instr_21_bF_buf11_), .B(datapath_1_RegisterFile_regfile_mem_6__15_), .C(datapath_1_Instr_22_bF_buf18_), .Y(_2732_) );
OAI22X1 OAI22X1_190 ( .A(_2732_), .B(_2731_), .C(datapath_1_Instr_22_bF_buf17_), .D(_2730_), .Y(_2733_) );
OAI21X1 OAI21X1_1796 ( .A(_1885__bF_buf8), .B(_2733_), .C(_1888__bF_buf4), .Y(_2734_) );
OAI22X1 OAI22X1_191 ( .A(_1888__bF_buf4), .B(_2723_), .C(_2729_), .D(_2734_), .Y(_2735_) );
NAND2X1 NAND2X1_1225 ( .A(_1917__bF_buf1), .B(_2735_), .Y(_2736_) );
AOI22X1 AOI22X1_155 ( .A(_1883__bF_buf3), .B(_1887__bF_buf1), .C(_2712_), .D(_2736_), .Y(datapath_1_RD1_15_) );
MUX2X1 MUX2X1_200 ( .A(datapath_1_RegisterFile_regfile_mem_9__16_), .B(datapath_1_RegisterFile_regfile_mem_8__16_), .S(datapath_1_Instr_21_bF_buf10_), .Y(_2737_) );
NOR2X1 NOR2X1_399 ( .A(datapath_1_RegisterFile_regfile_mem_11__16_), .B(_1890__bF_buf23), .Y(_2738_) );
OAI21X1 OAI21X1_1797 ( .A(datapath_1_Instr_21_bF_buf9_), .B(datapath_1_RegisterFile_regfile_mem_10__16_), .C(datapath_1_Instr_22_bF_buf16_), .Y(_2739_) );
OAI22X1 OAI22X1_192 ( .A(_2739_), .B(_2738_), .C(datapath_1_Instr_22_bF_buf15_), .D(_2737_), .Y(_2740_) );
INVX1 INVX1_434 ( .A(datapath_1_RegisterFile_regfile_mem_15__16_), .Y(_2741_) );
AOI21X1 AOI21X1_737 ( .A(_1890__bF_buf23), .B(datapath_1_RegisterFile_regfile_mem_14__16_), .C(_1884__bF_buf7), .Y(_2742_) );
OAI21X1 OAI21X1_1798 ( .A(_1890__bF_buf0), .B(_2741_), .C(_2742_), .Y(_2743_) );
NAND2X1 NAND2X1_1226 ( .A(datapath_1_RegisterFile_regfile_mem_12__16_), .B(_1890__bF_buf47), .Y(_2744_) );
AOI21X1 AOI21X1_738 ( .A(datapath_1_Instr_21_bF_buf8_), .B(datapath_1_RegisterFile_regfile_mem_13__16_), .C(datapath_1_Instr_22_bF_buf14_), .Y(_2745_) );
AOI21X1 AOI21X1_739 ( .A(_2744_), .B(_2745_), .C(_1885__bF_buf8), .Y(_2746_) );
AOI22X1 AOI22X1_156 ( .A(_2743_), .B(_2746_), .C(_1885__bF_buf8), .D(_2740_), .Y(_2747_) );
NOR2X1 NOR2X1_400 ( .A(datapath_1_Instr_21_bF_buf7_), .B(datapath_1_RegisterFile_regfile_mem_0__16_), .Y(_2748_) );
OAI21X1 OAI21X1_1799 ( .A(datapath_1_RegisterFile_regfile_mem_1__16_), .B(_1890__bF_buf18), .C(_1884__bF_buf8), .Y(_2749_) );
NOR2X1 NOR2X1_401 ( .A(datapath_1_RegisterFile_regfile_mem_3__16_), .B(_1890__bF_buf18), .Y(_2750_) );
OAI21X1 OAI21X1_1800 ( .A(datapath_1_Instr_21_bF_buf6_), .B(datapath_1_RegisterFile_regfile_mem_2__16_), .C(datapath_1_Instr_22_bF_buf13_), .Y(_2751_) );
OAI22X1 OAI22X1_193 ( .A(_2750_), .B(_2751_), .C(_2748_), .D(_2749_), .Y(_2752_) );
NOR2X1 NOR2X1_402 ( .A(datapath_1_Instr_23_bF_buf3_bF_buf3_), .B(_2752_), .Y(_2753_) );
MUX2X1 MUX2X1_201 ( .A(datapath_1_RegisterFile_regfile_mem_5__16_), .B(datapath_1_RegisterFile_regfile_mem_4__16_), .S(datapath_1_Instr_21_bF_buf5_), .Y(_2754_) );
NOR2X1 NOR2X1_403 ( .A(datapath_1_RegisterFile_regfile_mem_7__16_), .B(_1890__bF_buf16), .Y(_2755_) );
OAI21X1 OAI21X1_1801 ( .A(datapath_1_Instr_21_bF_buf4_), .B(datapath_1_RegisterFile_regfile_mem_6__16_), .C(datapath_1_Instr_22_bF_buf12_), .Y(_2756_) );
OAI22X1 OAI22X1_194 ( .A(_2756_), .B(_2755_), .C(datapath_1_Instr_22_bF_buf11_), .D(_2754_), .Y(_2757_) );
OAI21X1 OAI21X1_1802 ( .A(_1885__bF_buf2), .B(_2757_), .C(_1888__bF_buf7), .Y(_2758_) );
OAI22X1 OAI22X1_195 ( .A(_1888__bF_buf7), .B(_2747_), .C(_2753_), .D(_2758_), .Y(_2759_) );
NAND2X1 NAND2X1_1227 ( .A(_1917__bF_buf2), .B(_2759_), .Y(_2760_) );
INVX1 INVX1_435 ( .A(datapath_1_RegisterFile_regfile_mem_19__16_), .Y(_2761_) );
AOI21X1 AOI21X1_740 ( .A(datapath_1_Instr_23_bF_buf2_bF_buf3_), .B(datapath_1_RegisterFile_regfile_mem_23__16_), .C(_1890__bF_buf11), .Y(_2762_) );
OAI21X1 OAI21X1_1803 ( .A(datapath_1_Instr_23_bF_buf1_), .B(_2761_), .C(_2762_), .Y(_2763_) );
NAND2X1 NAND2X1_1228 ( .A(datapath_1_RegisterFile_regfile_mem_18__16_), .B(_1885__bF_buf3), .Y(_2764_) );
AOI21X1 AOI21X1_741 ( .A(datapath_1_Instr_23_bF_buf0_), .B(datapath_1_RegisterFile_regfile_mem_22__16_), .C(datapath_1_Instr_21_bF_buf3_), .Y(_2765_) );
AOI21X1 AOI21X1_742 ( .A(_2764_), .B(_2765_), .C(_1884__bF_buf2), .Y(_2766_) );
INVX1 INVX1_436 ( .A(datapath_1_RegisterFile_regfile_mem_17__16_), .Y(_2767_) );
AOI21X1 AOI21X1_743 ( .A(datapath_1_Instr_23_bF_buf15_bF_buf2_), .B(datapath_1_RegisterFile_regfile_mem_21__16_), .C(_1890__bF_buf43), .Y(_2768_) );
OAI21X1 OAI21X1_1804 ( .A(datapath_1_Instr_23_bF_buf14_bF_buf2_), .B(_2767_), .C(_2768_), .Y(_2769_) );
NAND2X1 NAND2X1_1229 ( .A(datapath_1_RegisterFile_regfile_mem_16__16_), .B(_1885__bF_buf3), .Y(_2770_) );
AOI21X1 AOI21X1_744 ( .A(datapath_1_Instr_23_bF_buf13_bF_buf2_), .B(datapath_1_RegisterFile_regfile_mem_20__16_), .C(datapath_1_Instr_21_bF_buf2_), .Y(_2771_) );
AOI21X1 AOI21X1_745 ( .A(_2770_), .B(_2771_), .C(datapath_1_Instr_22_bF_buf10_), .Y(_2772_) );
AOI22X1 AOI22X1_157 ( .A(_2766_), .B(_2763_), .C(_2769_), .D(_2772_), .Y(_2773_) );
NOR2X1 NOR2X1_404 ( .A(datapath_1_Instr_21_bF_buf1_), .B(datapath_1_RegisterFile_regfile_mem_24__16_), .Y(_2774_) );
OAI21X1 OAI21X1_1805 ( .A(datapath_1_RegisterFile_regfile_mem_25__16_), .B(_1890__bF_buf35), .C(_1884__bF_buf6), .Y(_2775_) );
NOR2X1 NOR2X1_405 ( .A(datapath_1_RegisterFile_regfile_mem_27__16_), .B(_1890__bF_buf35), .Y(_2776_) );
OAI21X1 OAI21X1_1806 ( .A(datapath_1_Instr_21_bF_buf0_), .B(datapath_1_RegisterFile_regfile_mem_26__16_), .C(datapath_1_Instr_22_bF_buf9_), .Y(_2777_) );
OAI22X1 OAI22X1_196 ( .A(_2776_), .B(_2777_), .C(_2774_), .D(_2775_), .Y(_2778_) );
NOR2X1 NOR2X1_406 ( .A(datapath_1_Instr_23_bF_buf12_bF_buf2_), .B(_2778_), .Y(_2779_) );
MUX2X1 MUX2X1_202 ( .A(datapath_1_RegisterFile_regfile_mem_29__16_), .B(datapath_1_RegisterFile_regfile_mem_28__16_), .S(datapath_1_Instr_21_bF_buf55_), .Y(_2780_) );
NOR2X1 NOR2X1_407 ( .A(datapath_1_RegisterFile_regfile_mem_31__16_), .B(_1890__bF_buf35), .Y(_2781_) );
OAI21X1 OAI21X1_1807 ( .A(datapath_1_Instr_21_bF_buf54_), .B(datapath_1_RegisterFile_regfile_mem_30__16_), .C(datapath_1_Instr_22_bF_buf8_), .Y(_2782_) );
OAI22X1 OAI22X1_197 ( .A(_2782_), .B(_2781_), .C(datapath_1_Instr_22_bF_buf7_), .D(_2780_), .Y(_2783_) );
OAI21X1 OAI21X1_1808 ( .A(_1885__bF_buf7), .B(_2783_), .C(datapath_1_Instr_24_bF_buf4_), .Y(_2784_) );
OAI22X1 OAI22X1_198 ( .A(datapath_1_Instr_24_bF_buf3_), .B(_2773_), .C(_2779_), .D(_2784_), .Y(_2785_) );
NAND2X1 NAND2X1_1230 ( .A(datapath_1_Instr_25_bF_buf3_), .B(_2785_), .Y(_2786_) );
AOI22X1 AOI22X1_158 ( .A(_1883__bF_buf3), .B(_1887__bF_buf0), .C(_2786_), .D(_2760_), .Y(datapath_1_RD1_16_) );
MUX2X1 MUX2X1_203 ( .A(datapath_1_RegisterFile_regfile_mem_9__17_), .B(datapath_1_RegisterFile_regfile_mem_8__17_), .S(datapath_1_Instr_21_bF_buf53_), .Y(_2787_) );
NOR2X1 NOR2X1_408 ( .A(datapath_1_RegisterFile_regfile_mem_11__17_), .B(_1890__bF_buf20), .Y(_2788_) );
OAI21X1 OAI21X1_1809 ( .A(datapath_1_Instr_21_bF_buf52_), .B(datapath_1_RegisterFile_regfile_mem_10__17_), .C(datapath_1_Instr_22_bF_buf6_), .Y(_2789_) );
OAI22X1 OAI22X1_199 ( .A(_2789_), .B(_2788_), .C(datapath_1_Instr_22_bF_buf5_), .D(_2787_), .Y(_2790_) );
INVX1 INVX1_437 ( .A(datapath_1_RegisterFile_regfile_mem_15__17_), .Y(_2791_) );
AOI21X1 AOI21X1_746 ( .A(_1890__bF_buf5), .B(datapath_1_RegisterFile_regfile_mem_14__17_), .C(_1884__bF_buf5), .Y(_2792_) );
OAI21X1 OAI21X1_1810 ( .A(_1890__bF_buf5), .B(_2791_), .C(_2792_), .Y(_2793_) );
NAND2X1 NAND2X1_1231 ( .A(datapath_1_RegisterFile_regfile_mem_12__17_), .B(_1890__bF_buf20), .Y(_2794_) );
AOI21X1 AOI21X1_747 ( .A(datapath_1_Instr_21_bF_buf51_), .B(datapath_1_RegisterFile_regfile_mem_13__17_), .C(datapath_1_Instr_22_bF_buf4_), .Y(_2795_) );
AOI21X1 AOI21X1_748 ( .A(_2794_), .B(_2795_), .C(_1885__bF_buf5), .Y(_2796_) );
AOI22X1 AOI22X1_159 ( .A(_2793_), .B(_2796_), .C(_1885__bF_buf5), .D(_2790_), .Y(_2797_) );
NOR2X1 NOR2X1_409 ( .A(datapath_1_Instr_21_bF_buf50_), .B(datapath_1_RegisterFile_regfile_mem_0__17_), .Y(_2798_) );
OAI21X1 OAI21X1_1811 ( .A(datapath_1_RegisterFile_regfile_mem_1__17_), .B(_1890__bF_buf1), .C(_1884__bF_buf4), .Y(_2799_) );
NOR2X1 NOR2X1_410 ( .A(datapath_1_RegisterFile_regfile_mem_3__17_), .B(_1890__bF_buf1), .Y(_2800_) );
OAI21X1 OAI21X1_1812 ( .A(datapath_1_Instr_21_bF_buf49_), .B(datapath_1_RegisterFile_regfile_mem_2__17_), .C(datapath_1_Instr_22_bF_buf3_), .Y(_2801_) );
OAI22X1 OAI22X1_200 ( .A(_2800_), .B(_2801_), .C(_2798_), .D(_2799_), .Y(_2802_) );
NOR2X1 NOR2X1_411 ( .A(datapath_1_Instr_23_bF_buf11_bF_buf2_), .B(_2802_), .Y(_2803_) );
MUX2X1 MUX2X1_204 ( .A(datapath_1_RegisterFile_regfile_mem_5__17_), .B(datapath_1_RegisterFile_regfile_mem_4__17_), .S(datapath_1_Instr_21_bF_buf48_), .Y(_2804_) );
NOR2X1 NOR2X1_412 ( .A(datapath_1_RegisterFile_regfile_mem_7__17_), .B(_1890__bF_buf27), .Y(_2805_) );
OAI21X1 OAI21X1_1813 ( .A(datapath_1_Instr_21_bF_buf47_), .B(datapath_1_RegisterFile_regfile_mem_6__17_), .C(datapath_1_Instr_22_bF_buf2_), .Y(_2806_) );
OAI22X1 OAI22X1_201 ( .A(_2806_), .B(_2805_), .C(datapath_1_Instr_22_bF_buf1_), .D(_2804_), .Y(_2807_) );
OAI21X1 OAI21X1_1814 ( .A(_1885__bF_buf4), .B(_2807_), .C(_1888__bF_buf2), .Y(_2808_) );
OAI22X1 OAI22X1_202 ( .A(_1888__bF_buf2), .B(_2797_), .C(_2803_), .D(_2808_), .Y(_2809_) );
NAND2X1 NAND2X1_1232 ( .A(_1917__bF_buf0), .B(_2809_), .Y(_2810_) );
INVX1 INVX1_438 ( .A(datapath_1_RegisterFile_regfile_mem_19__17_), .Y(_2811_) );
AOI21X1 AOI21X1_749 ( .A(datapath_1_Instr_23_bF_buf10_bF_buf2_), .B(datapath_1_RegisterFile_regfile_mem_23__17_), .C(_1890__bF_buf36), .Y(_2812_) );
OAI21X1 OAI21X1_1815 ( .A(datapath_1_Instr_23_bF_buf9_bF_buf2_), .B(_2811_), .C(_2812_), .Y(_2813_) );
NAND2X1 NAND2X1_1233 ( .A(datapath_1_RegisterFile_regfile_mem_18__17_), .B(_1885__bF_buf11), .Y(_2814_) );
AOI21X1 AOI21X1_750 ( .A(datapath_1_Instr_23_bF_buf8_bF_buf2_), .B(datapath_1_RegisterFile_regfile_mem_22__17_), .C(datapath_1_Instr_21_bF_buf46_), .Y(_2815_) );
AOI21X1 AOI21X1_751 ( .A(_2814_), .B(_2815_), .C(_1884__bF_buf9), .Y(_2816_) );
INVX1 INVX1_439 ( .A(datapath_1_RegisterFile_regfile_mem_17__17_), .Y(_2817_) );
AOI21X1 AOI21X1_752 ( .A(datapath_1_Instr_23_bF_buf7_bF_buf2_), .B(datapath_1_RegisterFile_regfile_mem_21__17_), .C(_1890__bF_buf36), .Y(_2818_) );
OAI21X1 OAI21X1_1816 ( .A(datapath_1_Instr_23_bF_buf6_bF_buf2_), .B(_2817_), .C(_2818_), .Y(_2819_) );
NAND2X1 NAND2X1_1234 ( .A(datapath_1_RegisterFile_regfile_mem_16__17_), .B(_1885__bF_buf11), .Y(_2820_) );
AOI21X1 AOI21X1_753 ( .A(datapath_1_Instr_23_bF_buf5_bF_buf2_), .B(datapath_1_RegisterFile_regfile_mem_20__17_), .C(datapath_1_Instr_21_bF_buf45_), .Y(_2821_) );
AOI21X1 AOI21X1_754 ( .A(_2820_), .B(_2821_), .C(datapath_1_Instr_22_bF_buf0_), .Y(_2822_) );
AOI22X1 AOI22X1_160 ( .A(_2816_), .B(_2813_), .C(_2819_), .D(_2822_), .Y(_2823_) );
NOR2X1 NOR2X1_413 ( .A(datapath_1_Instr_21_bF_buf44_), .B(datapath_1_RegisterFile_regfile_mem_24__17_), .Y(_2824_) );
OAI21X1 OAI21X1_1817 ( .A(datapath_1_RegisterFile_regfile_mem_25__17_), .B(_1890__bF_buf40), .C(_1884__bF_buf9), .Y(_2825_) );
NOR2X1 NOR2X1_414 ( .A(datapath_1_RegisterFile_regfile_mem_27__17_), .B(_1890__bF_buf40), .Y(_2826_) );
OAI21X1 OAI21X1_1818 ( .A(datapath_1_Instr_21_bF_buf43_), .B(datapath_1_RegisterFile_regfile_mem_26__17_), .C(datapath_1_Instr_22_bF_buf50_), .Y(_2827_) );
OAI22X1 OAI22X1_203 ( .A(_2826_), .B(_2827_), .C(_2824_), .D(_2825_), .Y(_2828_) );
NOR2X1 NOR2X1_415 ( .A(datapath_1_Instr_23_bF_buf4_bF_buf2_), .B(_2828_), .Y(_2829_) );
MUX2X1 MUX2X1_205 ( .A(datapath_1_RegisterFile_regfile_mem_29__17_), .B(datapath_1_RegisterFile_regfile_mem_28__17_), .S(datapath_1_Instr_21_bF_buf42_), .Y(_2830_) );
NOR2X1 NOR2X1_416 ( .A(datapath_1_RegisterFile_regfile_mem_31__17_), .B(_1890__bF_buf7), .Y(_2831_) );
OAI21X1 OAI21X1_1819 ( .A(datapath_1_Instr_21_bF_buf41_), .B(datapath_1_RegisterFile_regfile_mem_30__17_), .C(datapath_1_Instr_22_bF_buf49_), .Y(_2832_) );
OAI22X1 OAI22X1_204 ( .A(_2832_), .B(_2831_), .C(datapath_1_Instr_22_bF_buf48_), .D(_2830_), .Y(_2833_) );
OAI21X1 OAI21X1_1820 ( .A(_1885__bF_buf11), .B(_2833_), .C(datapath_1_Instr_24_bF_buf2_), .Y(_2834_) );
OAI22X1 OAI22X1_205 ( .A(datapath_1_Instr_24_bF_buf1_), .B(_2823_), .C(_2829_), .D(_2834_), .Y(_2835_) );
NAND2X1 NAND2X1_1235 ( .A(datapath_1_Instr_25_bF_buf2_), .B(_2835_), .Y(_2836_) );
AOI22X1 AOI22X1_161 ( .A(_1883__bF_buf2), .B(_1887__bF_buf4), .C(_2836_), .D(_2810_), .Y(datapath_1_RD1_17_) );
NAND2X1 NAND2X1_1236 ( .A(datapath_1_Instr_21_bF_buf40_), .B(datapath_1_RegisterFile_regfile_mem_27__18_), .Y(_2837_) );
NAND2X1 NAND2X1_1237 ( .A(datapath_1_RegisterFile_regfile_mem_26__18_), .B(_1890__bF_buf22), .Y(_2838_) );
NAND3X1 NAND3X1_1493 ( .A(datapath_1_Instr_22_bF_buf47_), .B(_2837_), .C(_2838_), .Y(_2839_) );
NAND2X1 NAND2X1_1238 ( .A(datapath_1_Instr_21_bF_buf39_), .B(datapath_1_RegisterFile_regfile_mem_25__18_), .Y(_2840_) );
AOI21X1 AOI21X1_755 ( .A(_1890__bF_buf22), .B(datapath_1_RegisterFile_regfile_mem_24__18_), .C(datapath_1_Instr_22_bF_buf46_), .Y(_2841_) );
NAND2X1 NAND2X1_1239 ( .A(_2840_), .B(_2841_), .Y(_2842_) );
NAND3X1 NAND3X1_1494 ( .A(_1885__bF_buf6), .B(_2839_), .C(_2842_), .Y(_2843_) );
NAND2X1 NAND2X1_1240 ( .A(datapath_1_Instr_21_bF_buf38_), .B(datapath_1_RegisterFile_regfile_mem_31__18_), .Y(_2844_) );
AOI21X1 AOI21X1_756 ( .A(_1890__bF_buf34), .B(datapath_1_RegisterFile_regfile_mem_30__18_), .C(_1884__bF_buf3), .Y(_2845_) );
NAND2X1 NAND2X1_1241 ( .A(_2844_), .B(_2845_), .Y(_2846_) );
INVX1 INVX1_440 ( .A(datapath_1_RegisterFile_regfile_mem_28__18_), .Y(_2847_) );
AOI21X1 AOI21X1_757 ( .A(datapath_1_Instr_21_bF_buf37_), .B(datapath_1_RegisterFile_regfile_mem_29__18_), .C(datapath_1_Instr_22_bF_buf45_), .Y(_2848_) );
OAI21X1 OAI21X1_1821 ( .A(datapath_1_Instr_21_bF_buf36_), .B(_2847_), .C(_2848_), .Y(_2849_) );
NAND3X1 NAND3X1_1495 ( .A(datapath_1_Instr_23_bF_buf3_bF_buf2_), .B(_2849_), .C(_2846_), .Y(_2850_) );
AOI21X1 AOI21X1_758 ( .A(_2843_), .B(_2850_), .C(_1888__bF_buf1), .Y(_2851_) );
MUX2X1 MUX2X1_206 ( .A(datapath_1_RegisterFile_regfile_mem_18__18_), .B(datapath_1_RegisterFile_regfile_mem_16__18_), .S(datapath_1_Instr_22_bF_buf44_), .Y(_2852_) );
NAND2X1 NAND2X1_1242 ( .A(_1890__bF_buf24), .B(_2852_), .Y(_2853_) );
MUX2X1 MUX2X1_207 ( .A(datapath_1_RegisterFile_regfile_mem_19__18_), .B(datapath_1_RegisterFile_regfile_mem_17__18_), .S(datapath_1_Instr_22_bF_buf43_), .Y(_2854_) );
NAND2X1 NAND2X1_1243 ( .A(datapath_1_Instr_21_bF_buf35_), .B(_2854_), .Y(_2855_) );
NAND3X1 NAND3X1_1496 ( .A(_1885__bF_buf9), .B(_2853_), .C(_2855_), .Y(_2856_) );
MUX2X1 MUX2X1_208 ( .A(datapath_1_RegisterFile_regfile_mem_22__18_), .B(datapath_1_RegisterFile_regfile_mem_20__18_), .S(datapath_1_Instr_22_bF_buf42_), .Y(_2857_) );
NAND2X1 NAND2X1_1244 ( .A(_1890__bF_buf24), .B(_2857_), .Y(_2858_) );
MUX2X1 MUX2X1_209 ( .A(datapath_1_RegisterFile_regfile_mem_23__18_), .B(datapath_1_RegisterFile_regfile_mem_21__18_), .S(datapath_1_Instr_22_bF_buf41_), .Y(_2859_) );
NAND2X1 NAND2X1_1245 ( .A(datapath_1_Instr_21_bF_buf34_), .B(_2859_), .Y(_2860_) );
NAND3X1 NAND3X1_1497 ( .A(datapath_1_Instr_23_bF_buf2_bF_buf2_), .B(_2858_), .C(_2860_), .Y(_2861_) );
AOI21X1 AOI21X1_759 ( .A(_2856_), .B(_2861_), .C(datapath_1_Instr_24_bF_buf0_), .Y(_2862_) );
OAI21X1 OAI21X1_1822 ( .A(_2862_), .B(_2851_), .C(datapath_1_Instr_25_bF_buf1_), .Y(_2863_) );
INVX1 INVX1_441 ( .A(datapath_1_RegisterFile_regfile_mem_9__18_), .Y(_2864_) );
AOI21X1 AOI21X1_760 ( .A(datapath_1_Instr_23_bF_buf1_), .B(datapath_1_RegisterFile_regfile_mem_13__18_), .C(_1890__bF_buf46), .Y(_2865_) );
OAI21X1 OAI21X1_1823 ( .A(datapath_1_Instr_23_bF_buf0_), .B(_2864_), .C(_2865_), .Y(_2866_) );
INVX1 INVX1_442 ( .A(datapath_1_RegisterFile_regfile_mem_8__18_), .Y(_2867_) );
AOI21X1 AOI21X1_761 ( .A(datapath_1_Instr_23_bF_buf15_bF_buf1_), .B(datapath_1_RegisterFile_regfile_mem_12__18_), .C(datapath_1_Instr_21_bF_buf33_), .Y(_2868_) );
OAI21X1 OAI21X1_1824 ( .A(datapath_1_Instr_23_bF_buf14_bF_buf1_), .B(_2867_), .C(_2868_), .Y(_2869_) );
NAND3X1 NAND3X1_1498 ( .A(_1884__bF_buf5), .B(_2869_), .C(_2866_), .Y(_2870_) );
INVX1 INVX1_443 ( .A(datapath_1_RegisterFile_regfile_mem_11__18_), .Y(_2871_) );
AOI21X1 AOI21X1_762 ( .A(datapath_1_Instr_23_bF_buf13_bF_buf1_), .B(datapath_1_RegisterFile_regfile_mem_15__18_), .C(_1890__bF_buf13), .Y(_2872_) );
OAI21X1 OAI21X1_1825 ( .A(datapath_1_Instr_23_bF_buf12_bF_buf1_), .B(_2871_), .C(_2872_), .Y(_2873_) );
INVX1 INVX1_444 ( .A(datapath_1_RegisterFile_regfile_mem_10__18_), .Y(_2874_) );
AOI21X1 AOI21X1_763 ( .A(datapath_1_Instr_23_bF_buf11_bF_buf1_), .B(datapath_1_RegisterFile_regfile_mem_14__18_), .C(datapath_1_Instr_21_bF_buf32_), .Y(_2875_) );
OAI21X1 OAI21X1_1826 ( .A(datapath_1_Instr_23_bF_buf10_bF_buf1_), .B(_2874_), .C(_2875_), .Y(_2876_) );
NAND3X1 NAND3X1_1499 ( .A(datapath_1_Instr_22_bF_buf40_), .B(_2876_), .C(_2873_), .Y(_2877_) );
AOI21X1 AOI21X1_764 ( .A(_2870_), .B(_2877_), .C(_1888__bF_buf2), .Y(_2878_) );
MUX2X1 MUX2X1_210 ( .A(datapath_1_RegisterFile_regfile_mem_1__18_), .B(datapath_1_RegisterFile_regfile_mem_0__18_), .S(datapath_1_Instr_21_bF_buf31_), .Y(_2879_) );
NOR2X1 NOR2X1_417 ( .A(datapath_1_RegisterFile_regfile_mem_3__18_), .B(_1890__bF_buf33), .Y(_2880_) );
OAI21X1 OAI21X1_1827 ( .A(datapath_1_Instr_21_bF_buf30_), .B(datapath_1_RegisterFile_regfile_mem_2__18_), .C(datapath_1_Instr_22_bF_buf39_), .Y(_2881_) );
OAI22X1 OAI22X1_206 ( .A(_2881_), .B(_2880_), .C(datapath_1_Instr_22_bF_buf38_), .D(_2879_), .Y(_2882_) );
NAND2X1 NAND2X1_1246 ( .A(_1885__bF_buf1), .B(_2882_), .Y(_2883_) );
MUX2X1 MUX2X1_211 ( .A(datapath_1_RegisterFile_regfile_mem_5__18_), .B(datapath_1_RegisterFile_regfile_mem_4__18_), .S(datapath_1_Instr_21_bF_buf29_), .Y(_2884_) );
NOR2X1 NOR2X1_418 ( .A(datapath_1_RegisterFile_regfile_mem_7__18_), .B(_1890__bF_buf13), .Y(_2885_) );
OAI21X1 OAI21X1_1828 ( .A(datapath_1_Instr_21_bF_buf28_), .B(datapath_1_RegisterFile_regfile_mem_6__18_), .C(datapath_1_Instr_22_bF_buf37_), .Y(_2886_) );
OAI22X1 OAI22X1_207 ( .A(_2886_), .B(_2885_), .C(datapath_1_Instr_22_bF_buf36_), .D(_2884_), .Y(_2887_) );
NAND2X1 NAND2X1_1247 ( .A(datapath_1_Instr_23_bF_buf9_bF_buf1_), .B(_2887_), .Y(_2888_) );
AOI21X1 AOI21X1_765 ( .A(_2883_), .B(_2888_), .C(datapath_1_Instr_24_bF_buf6_), .Y(_2889_) );
OAI21X1 OAI21X1_1829 ( .A(_2878_), .B(_2889_), .C(_1917__bF_buf4), .Y(_2890_) );
AOI22X1 AOI22X1_162 ( .A(_1883__bF_buf4), .B(_1887__bF_buf3), .C(_2863_), .D(_2890_), .Y(datapath_1_RD1_18_) );
NAND2X1 NAND2X1_1248 ( .A(datapath_1_Instr_21_bF_buf27_), .B(datapath_1_RegisterFile_regfile_mem_27__19_), .Y(_2891_) );
NAND2X1 NAND2X1_1249 ( .A(datapath_1_RegisterFile_regfile_mem_26__19_), .B(_1890__bF_buf32), .Y(_2892_) );
NAND3X1 NAND3X1_1500 ( .A(datapath_1_Instr_22_bF_buf35_), .B(_2891_), .C(_2892_), .Y(_2893_) );
NAND2X1 NAND2X1_1250 ( .A(datapath_1_Instr_21_bF_buf26_), .B(datapath_1_RegisterFile_regfile_mem_25__19_), .Y(_2894_) );
AOI21X1 AOI21X1_766 ( .A(_1890__bF_buf44), .B(datapath_1_RegisterFile_regfile_mem_24__19_), .C(datapath_1_Instr_22_bF_buf34_), .Y(_2895_) );
NAND2X1 NAND2X1_1251 ( .A(_2894_), .B(_2895_), .Y(_2896_) );
NAND3X1 NAND3X1_1501 ( .A(_1885__bF_buf7), .B(_2893_), .C(_2896_), .Y(_2897_) );
NAND2X1 NAND2X1_1252 ( .A(datapath_1_Instr_21_bF_buf25_), .B(datapath_1_RegisterFile_regfile_mem_31__19_), .Y(_2898_) );
AOI21X1 AOI21X1_767 ( .A(_1890__bF_buf32), .B(datapath_1_RegisterFile_regfile_mem_30__19_), .C(_1884__bF_buf2), .Y(_2899_) );
NAND2X1 NAND2X1_1253 ( .A(_2898_), .B(_2899_), .Y(_2900_) );
INVX1 INVX1_445 ( .A(datapath_1_RegisterFile_regfile_mem_28__19_), .Y(_2901_) );
AOI21X1 AOI21X1_768 ( .A(datapath_1_Instr_21_bF_buf24_), .B(datapath_1_RegisterFile_regfile_mem_29__19_), .C(datapath_1_Instr_22_bF_buf33_), .Y(_2902_) );
OAI21X1 OAI21X1_1830 ( .A(datapath_1_Instr_21_bF_buf23_), .B(_2901_), .C(_2902_), .Y(_2903_) );
NAND3X1 NAND3X1_1502 ( .A(datapath_1_Instr_23_bF_buf8_bF_buf1_), .B(_2903_), .C(_2900_), .Y(_2904_) );
AOI21X1 AOI21X1_769 ( .A(_2897_), .B(_2904_), .C(_1888__bF_buf0), .Y(_2905_) );
MUX2X1 MUX2X1_212 ( .A(datapath_1_RegisterFile_regfile_mem_18__19_), .B(datapath_1_RegisterFile_regfile_mem_16__19_), .S(datapath_1_Instr_22_bF_buf32_), .Y(_2906_) );
NAND2X1 NAND2X1_1254 ( .A(_1890__bF_buf31), .B(_2906_), .Y(_2907_) );
MUX2X1 MUX2X1_213 ( .A(datapath_1_RegisterFile_regfile_mem_19__19_), .B(datapath_1_RegisterFile_regfile_mem_17__19_), .S(datapath_1_Instr_22_bF_buf31_), .Y(_2908_) );
NAND2X1 NAND2X1_1255 ( .A(datapath_1_Instr_21_bF_buf22_), .B(_2908_), .Y(_2909_) );
NAND3X1 NAND3X1_1503 ( .A(_1885__bF_buf7), .B(_2907_), .C(_2909_), .Y(_2910_) );
MUX2X1 MUX2X1_214 ( .A(datapath_1_RegisterFile_regfile_mem_22__19_), .B(datapath_1_RegisterFile_regfile_mem_20__19_), .S(datapath_1_Instr_22_bF_buf30_), .Y(_2911_) );
NAND2X1 NAND2X1_1256 ( .A(_1890__bF_buf35), .B(_2911_), .Y(_2912_) );
MUX2X1 MUX2X1_215 ( .A(datapath_1_RegisterFile_regfile_mem_23__19_), .B(datapath_1_RegisterFile_regfile_mem_21__19_), .S(datapath_1_Instr_22_bF_buf29_), .Y(_2913_) );
NAND2X1 NAND2X1_1257 ( .A(datapath_1_Instr_21_bF_buf21_), .B(_2913_), .Y(_2914_) );
NAND3X1 NAND3X1_1504 ( .A(datapath_1_Instr_23_bF_buf7_bF_buf1_), .B(_2912_), .C(_2914_), .Y(_2915_) );
AOI21X1 AOI21X1_770 ( .A(_2910_), .B(_2915_), .C(datapath_1_Instr_24_bF_buf5_), .Y(_2916_) );
OAI21X1 OAI21X1_1831 ( .A(_2916_), .B(_2905_), .C(datapath_1_Instr_25_bF_buf0_), .Y(_2917_) );
MUX2X1 MUX2X1_216 ( .A(datapath_1_RegisterFile_regfile_mem_9__19_), .B(datapath_1_RegisterFile_regfile_mem_8__19_), .S(datapath_1_Instr_21_bF_buf20_), .Y(_2918_) );
NOR2X1 NOR2X1_419 ( .A(datapath_1_RegisterFile_regfile_mem_11__19_), .B(_1890__bF_buf16), .Y(_2919_) );
OAI21X1 OAI21X1_1832 ( .A(datapath_1_Instr_21_bF_buf19_), .B(datapath_1_RegisterFile_regfile_mem_10__19_), .C(datapath_1_Instr_22_bF_buf28_), .Y(_2920_) );
OAI22X1 OAI22X1_208 ( .A(_2920_), .B(_2919_), .C(datapath_1_Instr_22_bF_buf27_), .D(_2918_), .Y(_2921_) );
INVX1 INVX1_446 ( .A(datapath_1_RegisterFile_regfile_mem_15__19_), .Y(_2922_) );
AOI21X1 AOI21X1_771 ( .A(_1890__bF_buf16), .B(datapath_1_RegisterFile_regfile_mem_14__19_), .C(_1884__bF_buf0), .Y(_2923_) );
OAI21X1 OAI21X1_1833 ( .A(_1890__bF_buf16), .B(_2922_), .C(_2923_), .Y(_2924_) );
NAND2X1 NAND2X1_1258 ( .A(datapath_1_RegisterFile_regfile_mem_12__19_), .B(_1890__bF_buf16), .Y(_2925_) );
AOI21X1 AOI21X1_772 ( .A(datapath_1_Instr_21_bF_buf18_), .B(datapath_1_RegisterFile_regfile_mem_13__19_), .C(datapath_1_Instr_22_bF_buf26_), .Y(_2926_) );
AOI21X1 AOI21X1_773 ( .A(_2925_), .B(_2926_), .C(_1885__bF_buf2), .Y(_2927_) );
AOI22X1 AOI22X1_163 ( .A(_2924_), .B(_2927_), .C(_1885__bF_buf2), .D(_2921_), .Y(_2928_) );
NOR2X1 NOR2X1_420 ( .A(datapath_1_Instr_21_bF_buf17_), .B(datapath_1_RegisterFile_regfile_mem_0__19_), .Y(_2929_) );
OAI21X1 OAI21X1_1834 ( .A(datapath_1_RegisterFile_regfile_mem_1__19_), .B(_1890__bF_buf3), .C(_1884__bF_buf0), .Y(_2930_) );
NOR2X1 NOR2X1_421 ( .A(datapath_1_RegisterFile_regfile_mem_3__19_), .B(_1890__bF_buf3), .Y(_2931_) );
OAI21X1 OAI21X1_1835 ( .A(datapath_1_Instr_21_bF_buf16_), .B(datapath_1_RegisterFile_regfile_mem_2__19_), .C(datapath_1_Instr_22_bF_buf25_), .Y(_2932_) );
OAI22X1 OAI22X1_209 ( .A(_2931_), .B(_2932_), .C(_2929_), .D(_2930_), .Y(_2933_) );
NOR2X1 NOR2X1_422 ( .A(datapath_1_Instr_23_bF_buf6_bF_buf1_), .B(_2933_), .Y(_2934_) );
MUX2X1 MUX2X1_217 ( .A(datapath_1_RegisterFile_regfile_mem_5__19_), .B(datapath_1_RegisterFile_regfile_mem_4__19_), .S(datapath_1_Instr_21_bF_buf15_), .Y(_2935_) );
NOR2X1 NOR2X1_423 ( .A(datapath_1_RegisterFile_regfile_mem_7__19_), .B(_1890__bF_buf17), .Y(_2936_) );
OAI21X1 OAI21X1_1836 ( .A(datapath_1_Instr_21_bF_buf14_), .B(datapath_1_RegisterFile_regfile_mem_6__19_), .C(datapath_1_Instr_22_bF_buf24_), .Y(_2937_) );
OAI22X1 OAI22X1_210 ( .A(_2937_), .B(_2936_), .C(datapath_1_Instr_22_bF_buf23_), .D(_2935_), .Y(_2938_) );
OAI21X1 OAI21X1_1837 ( .A(_1885__bF_buf10), .B(_2938_), .C(_1888__bF_buf3), .Y(_2939_) );
OAI22X1 OAI22X1_211 ( .A(_1888__bF_buf3), .B(_2928_), .C(_2934_), .D(_2939_), .Y(_2940_) );
NAND2X1 NAND2X1_1259 ( .A(_1917__bF_buf1), .B(_2940_), .Y(_2941_) );
AOI22X1 AOI22X1_164 ( .A(_1883__bF_buf3), .B(_1887__bF_buf1), .C(_2917_), .D(_2941_), .Y(datapath_1_RD1_19_) );
NAND2X1 NAND2X1_1260 ( .A(datapath_1_Instr_21_bF_buf13_), .B(datapath_1_RegisterFile_regfile_mem_27__20_), .Y(_2942_) );
NAND2X1 NAND2X1_1261 ( .A(datapath_1_RegisterFile_regfile_mem_26__20_), .B(_1890__bF_buf29), .Y(_2943_) );
NAND3X1 NAND3X1_1505 ( .A(datapath_1_Instr_22_bF_buf22_), .B(_2942_), .C(_2943_), .Y(_2944_) );
NAND2X1 NAND2X1_1262 ( .A(datapath_1_Instr_21_bF_buf12_), .B(datapath_1_RegisterFile_regfile_mem_25__20_), .Y(_2945_) );
AOI21X1 AOI21X1_774 ( .A(_1890__bF_buf29), .B(datapath_1_RegisterFile_regfile_mem_24__20_), .C(datapath_1_Instr_22_bF_buf21_), .Y(_2946_) );
NAND2X1 NAND2X1_1263 ( .A(_2945_), .B(_2946_), .Y(_2947_) );
NAND3X1 NAND3X1_1506 ( .A(_1885__bF_buf10), .B(_2944_), .C(_2947_), .Y(_2948_) );
NAND2X1 NAND2X1_1264 ( .A(datapath_1_Instr_21_bF_buf11_), .B(datapath_1_RegisterFile_regfile_mem_31__20_), .Y(_2949_) );
AOI21X1 AOI21X1_775 ( .A(_1890__bF_buf29), .B(datapath_1_RegisterFile_regfile_mem_30__20_), .C(_1884__bF_buf7), .Y(_2950_) );
NAND2X1 NAND2X1_1265 ( .A(_2949_), .B(_2950_), .Y(_2951_) );
INVX1 INVX1_447 ( .A(datapath_1_RegisterFile_regfile_mem_28__20_), .Y(_2952_) );
AOI21X1 AOI21X1_776 ( .A(datapath_1_Instr_21_bF_buf10_), .B(datapath_1_RegisterFile_regfile_mem_29__20_), .C(datapath_1_Instr_22_bF_buf20_), .Y(_2953_) );
OAI21X1 OAI21X1_1838 ( .A(datapath_1_Instr_21_bF_buf9_), .B(_2952_), .C(_2953_), .Y(_2954_) );
NAND3X1 NAND3X1_1507 ( .A(datapath_1_Instr_23_bF_buf5_bF_buf1_), .B(_2954_), .C(_2951_), .Y(_2955_) );
AOI21X1 AOI21X1_777 ( .A(_2948_), .B(_2955_), .C(_1888__bF_buf4), .Y(_2956_) );
MUX2X1 MUX2X1_218 ( .A(datapath_1_RegisterFile_regfile_mem_18__20_), .B(datapath_1_RegisterFile_regfile_mem_16__20_), .S(datapath_1_Instr_22_bF_buf19_), .Y(_2957_) );
NAND2X1 NAND2X1_1266 ( .A(_1890__bF_buf31), .B(_2957_), .Y(_2958_) );
MUX2X1 MUX2X1_219 ( .A(datapath_1_RegisterFile_regfile_mem_19__20_), .B(datapath_1_RegisterFile_regfile_mem_17__20_), .S(datapath_1_Instr_22_bF_buf18_), .Y(_2959_) );
NAND2X1 NAND2X1_1267 ( .A(datapath_1_Instr_21_bF_buf8_), .B(_2959_), .Y(_2960_) );
NAND3X1 NAND3X1_1508 ( .A(_1885__bF_buf7), .B(_2958_), .C(_2960_), .Y(_2961_) );
MUX2X1 MUX2X1_220 ( .A(datapath_1_RegisterFile_regfile_mem_22__20_), .B(datapath_1_RegisterFile_regfile_mem_20__20_), .S(datapath_1_Instr_22_bF_buf17_), .Y(_2962_) );
NAND2X1 NAND2X1_1268 ( .A(_1890__bF_buf31), .B(_2962_), .Y(_2963_) );
MUX2X1 MUX2X1_221 ( .A(datapath_1_RegisterFile_regfile_mem_23__20_), .B(datapath_1_RegisterFile_regfile_mem_21__20_), .S(datapath_1_Instr_22_bF_buf16_), .Y(_2964_) );
NAND2X1 NAND2X1_1269 ( .A(datapath_1_Instr_21_bF_buf7_), .B(_2964_), .Y(_2965_) );
NAND3X1 NAND3X1_1509 ( .A(datapath_1_Instr_23_bF_buf4_bF_buf1_), .B(_2963_), .C(_2965_), .Y(_2966_) );
AOI21X1 AOI21X1_778 ( .A(_2961_), .B(_2966_), .C(datapath_1_Instr_24_bF_buf4_), .Y(_2967_) );
OAI21X1 OAI21X1_1839 ( .A(_2967_), .B(_2956_), .C(datapath_1_Instr_25_bF_buf5_), .Y(_2968_) );
MUX2X1 MUX2X1_222 ( .A(datapath_1_RegisterFile_regfile_mem_9__20_), .B(datapath_1_RegisterFile_regfile_mem_8__20_), .S(datapath_1_Instr_21_bF_buf6_), .Y(_2969_) );
NOR2X1 NOR2X1_424 ( .A(datapath_1_RegisterFile_regfile_mem_11__20_), .B(_1890__bF_buf3), .Y(_2970_) );
OAI21X1 OAI21X1_1840 ( .A(datapath_1_Instr_21_bF_buf5_), .B(datapath_1_RegisterFile_regfile_mem_10__20_), .C(datapath_1_Instr_22_bF_buf15_), .Y(_2971_) );
OAI22X1 OAI22X1_212 ( .A(_2971_), .B(_2970_), .C(datapath_1_Instr_22_bF_buf14_), .D(_2969_), .Y(_2972_) );
INVX1 INVX1_448 ( .A(datapath_1_RegisterFile_regfile_mem_15__20_), .Y(_2973_) );
AOI21X1 AOI21X1_779 ( .A(_1890__bF_buf3), .B(datapath_1_RegisterFile_regfile_mem_14__20_), .C(_1884__bF_buf0), .Y(_2974_) );
OAI21X1 OAI21X1_1841 ( .A(_1890__bF_buf3), .B(_2973_), .C(_2974_), .Y(_2975_) );
NAND2X1 NAND2X1_1270 ( .A(datapath_1_RegisterFile_regfile_mem_12__20_), .B(_1890__bF_buf3), .Y(_2976_) );
AOI21X1 AOI21X1_780 ( .A(datapath_1_Instr_21_bF_buf4_), .B(datapath_1_RegisterFile_regfile_mem_13__20_), .C(datapath_1_Instr_22_bF_buf13_), .Y(_2977_) );
AOI21X1 AOI21X1_781 ( .A(_2976_), .B(_2977_), .C(_1885__bF_buf2), .Y(_2978_) );
AOI22X1 AOI22X1_165 ( .A(_2975_), .B(_2978_), .C(_1885__bF_buf2), .D(_2972_), .Y(_2979_) );
NOR2X1 NOR2X1_425 ( .A(datapath_1_Instr_21_bF_buf3_), .B(datapath_1_RegisterFile_regfile_mem_0__20_), .Y(_2980_) );
OAI21X1 OAI21X1_1842 ( .A(datapath_1_RegisterFile_regfile_mem_1__20_), .B(_1890__bF_buf18), .C(_1884__bF_buf0), .Y(_2981_) );
NOR2X1 NOR2X1_426 ( .A(datapath_1_RegisterFile_regfile_mem_3__20_), .B(_1890__bF_buf18), .Y(_2982_) );
OAI21X1 OAI21X1_1843 ( .A(datapath_1_Instr_21_bF_buf2_), .B(datapath_1_RegisterFile_regfile_mem_2__20_), .C(datapath_1_Instr_22_bF_buf12_), .Y(_2983_) );
OAI22X1 OAI22X1_213 ( .A(_2982_), .B(_2983_), .C(_2980_), .D(_2981_), .Y(_2984_) );
NOR2X1 NOR2X1_427 ( .A(datapath_1_Instr_23_bF_buf3_bF_buf1_), .B(_2984_), .Y(_2985_) );
MUX2X1 MUX2X1_223 ( .A(datapath_1_RegisterFile_regfile_mem_5__20_), .B(datapath_1_RegisterFile_regfile_mem_4__20_), .S(datapath_1_Instr_21_bF_buf1_), .Y(_2986_) );
NOR2X1 NOR2X1_428 ( .A(datapath_1_RegisterFile_regfile_mem_7__20_), .B(_1890__bF_buf16), .Y(_2987_) );
OAI21X1 OAI21X1_1844 ( .A(datapath_1_Instr_21_bF_buf0_), .B(datapath_1_RegisterFile_regfile_mem_6__20_), .C(datapath_1_Instr_22_bF_buf11_), .Y(_2988_) );
OAI22X1 OAI22X1_214 ( .A(_2988_), .B(_2987_), .C(datapath_1_Instr_22_bF_buf10_), .D(_2986_), .Y(_2989_) );
OAI21X1 OAI21X1_1845 ( .A(_1885__bF_buf2), .B(_2989_), .C(_1888__bF_buf7), .Y(_2990_) );
OAI22X1 OAI22X1_215 ( .A(_1888__bF_buf7), .B(_2979_), .C(_2985_), .D(_2990_), .Y(_2991_) );
NAND2X1 NAND2X1_1271 ( .A(_1917__bF_buf2), .B(_2991_), .Y(_2992_) );
AOI22X1 AOI22X1_166 ( .A(_1883__bF_buf1), .B(_1887__bF_buf0), .C(_2968_), .D(_2992_), .Y(datapath_1_RD1_20_) );
MUX2X1 MUX2X1_224 ( .A(datapath_1_RegisterFile_regfile_mem_9__21_), .B(datapath_1_RegisterFile_regfile_mem_8__21_), .S(datapath_1_Instr_21_bF_buf55_), .Y(_2993_) );
NOR2X1 NOR2X1_429 ( .A(datapath_1_RegisterFile_regfile_mem_11__21_), .B(_1890__bF_buf28), .Y(_2994_) );
OAI21X1 OAI21X1_1846 ( .A(datapath_1_Instr_21_bF_buf54_), .B(datapath_1_RegisterFile_regfile_mem_10__21_), .C(datapath_1_Instr_22_bF_buf9_), .Y(_2995_) );
OAI22X1 OAI22X1_216 ( .A(_2995_), .B(_2994_), .C(datapath_1_Instr_22_bF_buf8_), .D(_2993_), .Y(_2996_) );
INVX1 INVX1_449 ( .A(datapath_1_RegisterFile_regfile_mem_15__21_), .Y(_2997_) );
AOI21X1 AOI21X1_782 ( .A(_1890__bF_buf26), .B(datapath_1_RegisterFile_regfile_mem_14__21_), .C(_1884__bF_buf1), .Y(_2998_) );
OAI21X1 OAI21X1_1847 ( .A(_1890__bF_buf26), .B(_2997_), .C(_2998_), .Y(_2999_) );
NAND2X1 NAND2X1_1272 ( .A(datapath_1_RegisterFile_regfile_mem_12__21_), .B(_1890__bF_buf26), .Y(_3000_) );
AOI21X1 AOI21X1_783 ( .A(datapath_1_Instr_21_bF_buf53_), .B(datapath_1_RegisterFile_regfile_mem_13__21_), .C(datapath_1_Instr_22_bF_buf7_), .Y(_3001_) );
AOI21X1 AOI21X1_784 ( .A(_3000_), .B(_3001_), .C(_1885__bF_buf5), .Y(_3002_) );
AOI22X1 AOI22X1_167 ( .A(_2999_), .B(_3002_), .C(_1885__bF_buf5), .D(_2996_), .Y(_3003_) );
NOR2X1 NOR2X1_430 ( .A(datapath_1_Instr_21_bF_buf52_), .B(datapath_1_RegisterFile_regfile_mem_0__21_), .Y(_3004_) );
OAI21X1 OAI21X1_1848 ( .A(datapath_1_RegisterFile_regfile_mem_1__21_), .B(_1890__bF_buf38), .C(_1884__bF_buf4), .Y(_3005_) );
NOR2X1 NOR2X1_431 ( .A(datapath_1_RegisterFile_regfile_mem_3__21_), .B(_1890__bF_buf38), .Y(_3006_) );
OAI21X1 OAI21X1_1849 ( .A(datapath_1_Instr_21_bF_buf51_), .B(datapath_1_RegisterFile_regfile_mem_2__21_), .C(datapath_1_Instr_22_bF_buf6_), .Y(_3007_) );
OAI22X1 OAI22X1_217 ( .A(_3006_), .B(_3007_), .C(_3004_), .D(_3005_), .Y(_3008_) );
NOR2X1 NOR2X1_432 ( .A(datapath_1_Instr_23_bF_buf2_bF_buf1_), .B(_3008_), .Y(_3009_) );
MUX2X1 MUX2X1_225 ( .A(datapath_1_RegisterFile_regfile_mem_5__21_), .B(datapath_1_RegisterFile_regfile_mem_4__21_), .S(datapath_1_Instr_21_bF_buf50_), .Y(_3010_) );
NOR2X1 NOR2X1_433 ( .A(datapath_1_RegisterFile_regfile_mem_7__21_), .B(_1890__bF_buf38), .Y(_3011_) );
OAI21X1 OAI21X1_1850 ( .A(datapath_1_Instr_21_bF_buf49_), .B(datapath_1_RegisterFile_regfile_mem_6__21_), .C(datapath_1_Instr_22_bF_buf5_), .Y(_3012_) );
OAI22X1 OAI22X1_218 ( .A(_3012_), .B(_3011_), .C(datapath_1_Instr_22_bF_buf4_), .D(_3010_), .Y(_3013_) );
OAI21X1 OAI21X1_1851 ( .A(_1885__bF_buf4), .B(_3013_), .C(_1888__bF_buf6), .Y(_3014_) );
OAI22X1 OAI22X1_219 ( .A(_1888__bF_buf6), .B(_3003_), .C(_3009_), .D(_3014_), .Y(_3015_) );
NAND2X1 NAND2X1_1273 ( .A(_1917__bF_buf3), .B(_3015_), .Y(_3016_) );
INVX1 INVX1_450 ( .A(datapath_1_RegisterFile_regfile_mem_19__21_), .Y(_3017_) );
AOI21X1 AOI21X1_785 ( .A(datapath_1_Instr_23_bF_buf1_), .B(datapath_1_RegisterFile_regfile_mem_23__21_), .C(_1890__bF_buf36), .Y(_3018_) );
OAI21X1 OAI21X1_1852 ( .A(datapath_1_Instr_23_bF_buf0_), .B(_3017_), .C(_3018_), .Y(_3019_) );
NAND2X1 NAND2X1_1274 ( .A(datapath_1_RegisterFile_regfile_mem_18__21_), .B(_1885__bF_buf11), .Y(_3020_) );
AOI21X1 AOI21X1_786 ( .A(datapath_1_Instr_23_bF_buf15_bF_buf0_), .B(datapath_1_RegisterFile_regfile_mem_22__21_), .C(datapath_1_Instr_21_bF_buf48_), .Y(_3021_) );
AOI21X1 AOI21X1_787 ( .A(_3020_), .B(_3021_), .C(_1884__bF_buf9), .Y(_3022_) );
INVX1 INVX1_451 ( .A(datapath_1_RegisterFile_regfile_mem_17__21_), .Y(_3023_) );
AOI21X1 AOI21X1_788 ( .A(datapath_1_Instr_23_bF_buf14_bF_buf0_), .B(datapath_1_RegisterFile_regfile_mem_21__21_), .C(_1890__bF_buf36), .Y(_3024_) );
OAI21X1 OAI21X1_1853 ( .A(datapath_1_Instr_23_bF_buf13_bF_buf0_), .B(_3023_), .C(_3024_), .Y(_3025_) );
NAND2X1 NAND2X1_1275 ( .A(datapath_1_RegisterFile_regfile_mem_16__21_), .B(_1885__bF_buf11), .Y(_3026_) );
AOI21X1 AOI21X1_789 ( .A(datapath_1_Instr_23_bF_buf12_bF_buf0_), .B(datapath_1_RegisterFile_regfile_mem_20__21_), .C(datapath_1_Instr_21_bF_buf47_), .Y(_3027_) );
AOI21X1 AOI21X1_790 ( .A(_3026_), .B(_3027_), .C(datapath_1_Instr_22_bF_buf3_), .Y(_3028_) );
AOI22X1 AOI22X1_168 ( .A(_3022_), .B(_3019_), .C(_3025_), .D(_3028_), .Y(_3029_) );
NOR2X1 NOR2X1_434 ( .A(datapath_1_Instr_21_bF_buf46_), .B(datapath_1_RegisterFile_regfile_mem_24__21_), .Y(_3030_) );
OAI21X1 OAI21X1_1854 ( .A(datapath_1_RegisterFile_regfile_mem_25__21_), .B(_1890__bF_buf7), .C(_1884__bF_buf9), .Y(_3031_) );
NOR2X1 NOR2X1_435 ( .A(datapath_1_RegisterFile_regfile_mem_27__21_), .B(_1890__bF_buf36), .Y(_3032_) );
OAI21X1 OAI21X1_1855 ( .A(datapath_1_Instr_21_bF_buf45_), .B(datapath_1_RegisterFile_regfile_mem_26__21_), .C(datapath_1_Instr_22_bF_buf2_), .Y(_3033_) );
OAI22X1 OAI22X1_220 ( .A(_3032_), .B(_3033_), .C(_3030_), .D(_3031_), .Y(_3034_) );
NOR2X1 NOR2X1_436 ( .A(datapath_1_Instr_23_bF_buf11_bF_buf0_), .B(_3034_), .Y(_3035_) );
MUX2X1 MUX2X1_226 ( .A(datapath_1_RegisterFile_regfile_mem_29__21_), .B(datapath_1_RegisterFile_regfile_mem_28__21_), .S(datapath_1_Instr_21_bF_buf44_), .Y(_3036_) );
NOR2X1 NOR2X1_437 ( .A(datapath_1_RegisterFile_regfile_mem_31__21_), .B(_1890__bF_buf7), .Y(_3037_) );
OAI21X1 OAI21X1_1856 ( .A(datapath_1_Instr_21_bF_buf43_), .B(datapath_1_RegisterFile_regfile_mem_30__21_), .C(datapath_1_Instr_22_bF_buf1_), .Y(_3038_) );
OAI22X1 OAI22X1_221 ( .A(_3038_), .B(_3037_), .C(datapath_1_Instr_22_bF_buf0_), .D(_3036_), .Y(_3039_) );
OAI21X1 OAI21X1_1857 ( .A(_1885__bF_buf11), .B(_3039_), .C(datapath_1_Instr_24_bF_buf3_), .Y(_3040_) );
OAI22X1 OAI22X1_222 ( .A(datapath_1_Instr_24_bF_buf2_), .B(_3029_), .C(_3035_), .D(_3040_), .Y(_3041_) );
NAND2X1 NAND2X1_1276 ( .A(datapath_1_Instr_25_bF_buf4_), .B(_3041_), .Y(_3042_) );
AOI22X1 AOI22X1_169 ( .A(_1883__bF_buf0), .B(_1887__bF_buf4), .C(_3042_), .D(_3016_), .Y(datapath_1_RD1_21_) );
MUX2X1 MUX2X1_227 ( .A(datapath_1_RegisterFile_regfile_mem_9__22_), .B(datapath_1_RegisterFile_regfile_mem_8__22_), .S(datapath_1_Instr_21_bF_buf42_), .Y(_3043_) );
NOR2X1 NOR2X1_438 ( .A(datapath_1_RegisterFile_regfile_mem_11__22_), .B(_1890__bF_buf13), .Y(_3044_) );
OAI21X1 OAI21X1_1858 ( .A(datapath_1_Instr_21_bF_buf41_), .B(datapath_1_RegisterFile_regfile_mem_10__22_), .C(datapath_1_Instr_22_bF_buf50_), .Y(_3045_) );
OAI22X1 OAI22X1_223 ( .A(_3045_), .B(_3044_), .C(datapath_1_Instr_22_bF_buf49_), .D(_3043_), .Y(_3046_) );
INVX1 INVX1_452 ( .A(datapath_1_RegisterFile_regfile_mem_15__22_), .Y(_3047_) );
AOI21X1 AOI21X1_791 ( .A(_1890__bF_buf13), .B(datapath_1_RegisterFile_regfile_mem_14__22_), .C(_1884__bF_buf5), .Y(_3048_) );
OAI21X1 OAI21X1_1859 ( .A(_1890__bF_buf13), .B(_3047_), .C(_3048_), .Y(_3049_) );
NAND2X1 NAND2X1_1277 ( .A(datapath_1_RegisterFile_regfile_mem_12__22_), .B(_1890__bF_buf13), .Y(_3050_) );
AOI21X1 AOI21X1_792 ( .A(datapath_1_Instr_21_bF_buf40_), .B(datapath_1_RegisterFile_regfile_mem_13__22_), .C(datapath_1_Instr_22_bF_buf48_), .Y(_3051_) );
AOI21X1 AOI21X1_793 ( .A(_3050_), .B(_3051_), .C(_1885__bF_buf1), .Y(_3052_) );
AOI22X1 AOI22X1_170 ( .A(_3049_), .B(_3052_), .C(_1885__bF_buf1), .D(_3046_), .Y(_3053_) );
NOR2X1 NOR2X1_439 ( .A(datapath_1_Instr_21_bF_buf39_), .B(datapath_1_RegisterFile_regfile_mem_0__22_), .Y(_3054_) );
OAI21X1 OAI21X1_1860 ( .A(datapath_1_RegisterFile_regfile_mem_1__22_), .B(_1890__bF_buf30), .C(_1884__bF_buf3), .Y(_3055_) );
NOR2X1 NOR2X1_440 ( .A(datapath_1_RegisterFile_regfile_mem_3__22_), .B(_1890__bF_buf30), .Y(_3056_) );
OAI21X1 OAI21X1_1861 ( .A(datapath_1_Instr_21_bF_buf38_), .B(datapath_1_RegisterFile_regfile_mem_2__22_), .C(datapath_1_Instr_22_bF_buf47_), .Y(_3057_) );
OAI22X1 OAI22X1_224 ( .A(_3056_), .B(_3057_), .C(_3054_), .D(_3055_), .Y(_3058_) );
NOR2X1 NOR2X1_441 ( .A(datapath_1_Instr_23_bF_buf10_bF_buf0_), .B(_3058_), .Y(_3059_) );
MUX2X1 MUX2X1_228 ( .A(datapath_1_RegisterFile_regfile_mem_5__22_), .B(datapath_1_RegisterFile_regfile_mem_4__22_), .S(datapath_1_Instr_21_bF_buf37_), .Y(_3060_) );
NOR2X1 NOR2X1_442 ( .A(datapath_1_RegisterFile_regfile_mem_7__22_), .B(_1890__bF_buf33), .Y(_3061_) );
OAI21X1 OAI21X1_1862 ( .A(datapath_1_Instr_21_bF_buf36_), .B(datapath_1_RegisterFile_regfile_mem_6__22_), .C(datapath_1_Instr_22_bF_buf46_), .Y(_3062_) );
OAI22X1 OAI22X1_225 ( .A(_3062_), .B(_3061_), .C(datapath_1_Instr_22_bF_buf45_), .D(_3060_), .Y(_3063_) );
OAI21X1 OAI21X1_1863 ( .A(_1885__bF_buf1), .B(_3063_), .C(_1888__bF_buf2), .Y(_3064_) );
OAI22X1 OAI22X1_226 ( .A(_1888__bF_buf2), .B(_3053_), .C(_3059_), .D(_3064_), .Y(_3065_) );
NAND2X1 NAND2X1_1278 ( .A(_1917__bF_buf0), .B(_3065_), .Y(_3066_) );
INVX1 INVX1_453 ( .A(datapath_1_RegisterFile_regfile_mem_19__22_), .Y(_3067_) );
AOI21X1 AOI21X1_794 ( .A(datapath_1_Instr_23_bF_buf9_bF_buf0_), .B(datapath_1_RegisterFile_regfile_mem_23__22_), .C(_1890__bF_buf9), .Y(_3068_) );
OAI21X1 OAI21X1_1864 ( .A(datapath_1_Instr_23_bF_buf8_bF_buf0_), .B(_3067_), .C(_3068_), .Y(_3069_) );
NAND2X1 NAND2X1_1279 ( .A(datapath_1_RegisterFile_regfile_mem_18__22_), .B(_1885__bF_buf9), .Y(_3070_) );
AOI21X1 AOI21X1_795 ( .A(datapath_1_Instr_23_bF_buf7_bF_buf0_), .B(datapath_1_RegisterFile_regfile_mem_22__22_), .C(datapath_1_Instr_21_bF_buf35_), .Y(_3071_) );
AOI21X1 AOI21X1_796 ( .A(_3070_), .B(_3071_), .C(_1884__bF_buf9), .Y(_3072_) );
INVX1 INVX1_454 ( .A(datapath_1_RegisterFile_regfile_mem_17__22_), .Y(_3073_) );
AOI21X1 AOI21X1_797 ( .A(datapath_1_Instr_23_bF_buf6_bF_buf0_), .B(datapath_1_RegisterFile_regfile_mem_21__22_), .C(_1890__bF_buf9), .Y(_3074_) );
OAI21X1 OAI21X1_1865 ( .A(datapath_1_Instr_23_bF_buf5_bF_buf0_), .B(_3073_), .C(_3074_), .Y(_3075_) );
NAND2X1 NAND2X1_1280 ( .A(datapath_1_RegisterFile_regfile_mem_16__22_), .B(_1885__bF_buf9), .Y(_3076_) );
AOI21X1 AOI21X1_798 ( .A(datapath_1_Instr_23_bF_buf4_bF_buf0_), .B(datapath_1_RegisterFile_regfile_mem_20__22_), .C(datapath_1_Instr_21_bF_buf34_), .Y(_3077_) );
AOI21X1 AOI21X1_799 ( .A(_3076_), .B(_3077_), .C(datapath_1_Instr_22_bF_buf44_), .Y(_3078_) );
AOI22X1 AOI22X1_171 ( .A(_3072_), .B(_3069_), .C(_3075_), .D(_3078_), .Y(_3079_) );
NOR2X1 NOR2X1_443 ( .A(datapath_1_Instr_21_bF_buf33_), .B(datapath_1_RegisterFile_regfile_mem_24__22_), .Y(_3080_) );
OAI21X1 OAI21X1_1866 ( .A(datapath_1_RegisterFile_regfile_mem_25__22_), .B(_1890__bF_buf37), .C(_1884__bF_buf3), .Y(_3081_) );
NOR2X1 NOR2X1_444 ( .A(datapath_1_RegisterFile_regfile_mem_27__22_), .B(_1890__bF_buf37), .Y(_3082_) );
OAI21X1 OAI21X1_1867 ( .A(datapath_1_Instr_21_bF_buf32_), .B(datapath_1_RegisterFile_regfile_mem_26__22_), .C(datapath_1_Instr_22_bF_buf43_), .Y(_3083_) );
OAI22X1 OAI22X1_227 ( .A(_3082_), .B(_3083_), .C(_3080_), .D(_3081_), .Y(_3084_) );
NOR2X1 NOR2X1_445 ( .A(datapath_1_Instr_23_bF_buf3_bF_buf0_), .B(_3084_), .Y(_3085_) );
MUX2X1 MUX2X1_229 ( .A(datapath_1_RegisterFile_regfile_mem_29__22_), .B(datapath_1_RegisterFile_regfile_mem_28__22_), .S(datapath_1_Instr_21_bF_buf31_), .Y(_3086_) );
NOR2X1 NOR2X1_446 ( .A(datapath_1_RegisterFile_regfile_mem_31__22_), .B(_1890__bF_buf37), .Y(_3087_) );
OAI21X1 OAI21X1_1868 ( .A(datapath_1_Instr_21_bF_buf30_), .B(datapath_1_RegisterFile_regfile_mem_30__22_), .C(datapath_1_Instr_22_bF_buf42_), .Y(_3088_) );
OAI22X1 OAI22X1_228 ( .A(_3088_), .B(_3087_), .C(datapath_1_Instr_22_bF_buf41_), .D(_3086_), .Y(_3089_) );
OAI21X1 OAI21X1_1869 ( .A(_1885__bF_buf9), .B(_3089_), .C(datapath_1_Instr_24_bF_buf1_), .Y(_3090_) );
OAI22X1 OAI22X1_229 ( .A(datapath_1_Instr_24_bF_buf0_), .B(_3079_), .C(_3085_), .D(_3090_), .Y(_3091_) );
NAND2X1 NAND2X1_1281 ( .A(datapath_1_Instr_25_bF_buf3_), .B(_3091_), .Y(_3092_) );
AOI22X1 AOI22X1_172 ( .A(_1883__bF_buf2), .B(_1887__bF_buf4), .C(_3092_), .D(_3066_), .Y(datapath_1_RD1_22_) );
MUX2X1 MUX2X1_230 ( .A(datapath_1_RegisterFile_regfile_mem_2__23_), .B(datapath_1_RegisterFile_regfile_mem_0__23_), .S(datapath_1_Instr_22_bF_buf40_), .Y(_3093_) );
NAND2X1 NAND2X1_1282 ( .A(_1890__bF_buf46), .B(_3093_), .Y(_3094_) );
MUX2X1 MUX2X1_231 ( .A(datapath_1_RegisterFile_regfile_mem_3__23_), .B(datapath_1_RegisterFile_regfile_mem_1__23_), .S(datapath_1_Instr_22_bF_buf39_), .Y(_3095_) );
NAND2X1 NAND2X1_1283 ( .A(datapath_1_Instr_21_bF_buf29_), .B(_3095_), .Y(_3096_) );
NAND3X1 NAND3X1_1510 ( .A(_1885__bF_buf1), .B(_3094_), .C(_3096_), .Y(_3097_) );
MUX2X1 MUX2X1_232 ( .A(datapath_1_RegisterFile_regfile_mem_6__23_), .B(datapath_1_RegisterFile_regfile_mem_4__23_), .S(datapath_1_Instr_22_bF_buf38_), .Y(_3098_) );
NAND2X1 NAND2X1_1284 ( .A(_1890__bF_buf46), .B(_3098_), .Y(_3099_) );
MUX2X1 MUX2X1_233 ( .A(datapath_1_RegisterFile_regfile_mem_7__23_), .B(datapath_1_RegisterFile_regfile_mem_5__23_), .S(datapath_1_Instr_22_bF_buf37_), .Y(_3100_) );
NAND2X1 NAND2X1_1285 ( .A(datapath_1_Instr_21_bF_buf28_), .B(_3100_), .Y(_3101_) );
NAND3X1 NAND3X1_1511 ( .A(datapath_1_Instr_23_bF_buf2_bF_buf0_), .B(_3099_), .C(_3101_), .Y(_3102_) );
AOI21X1 AOI21X1_800 ( .A(_3097_), .B(_3102_), .C(datapath_1_Instr_24_bF_buf6_), .Y(_3103_) );
INVX1 INVX1_455 ( .A(datapath_1_RegisterFile_regfile_mem_9__23_), .Y(_3104_) );
AOI21X1 AOI21X1_801 ( .A(datapath_1_Instr_23_bF_buf1_), .B(datapath_1_RegisterFile_regfile_mem_13__23_), .C(_1890__bF_buf46), .Y(_3105_) );
OAI21X1 OAI21X1_1870 ( .A(datapath_1_Instr_23_bF_buf0_), .B(_3104_), .C(_3105_), .Y(_3106_) );
INVX1 INVX1_456 ( .A(datapath_1_RegisterFile_regfile_mem_8__23_), .Y(_3107_) );
AOI21X1 AOI21X1_802 ( .A(datapath_1_Instr_23_bF_buf15_bF_buf3_), .B(datapath_1_RegisterFile_regfile_mem_12__23_), .C(datapath_1_Instr_21_bF_buf27_), .Y(_3108_) );
OAI21X1 OAI21X1_1871 ( .A(datapath_1_Instr_23_bF_buf14_bF_buf3_), .B(_3107_), .C(_3108_), .Y(_3109_) );
NAND3X1 NAND3X1_1512 ( .A(_1884__bF_buf5), .B(_3109_), .C(_3106_), .Y(_3110_) );
INVX1 INVX1_457 ( .A(datapath_1_RegisterFile_regfile_mem_11__23_), .Y(_3111_) );
AOI21X1 AOI21X1_803 ( .A(datapath_1_Instr_23_bF_buf13_bF_buf3_), .B(datapath_1_RegisterFile_regfile_mem_15__23_), .C(_1890__bF_buf46), .Y(_3112_) );
OAI21X1 OAI21X1_1872 ( .A(datapath_1_Instr_23_bF_buf12_bF_buf3_), .B(_3111_), .C(_3112_), .Y(_3113_) );
INVX1 INVX1_458 ( .A(datapath_1_RegisterFile_regfile_mem_10__23_), .Y(_3114_) );
AOI21X1 AOI21X1_804 ( .A(datapath_1_Instr_23_bF_buf11_bF_buf3_), .B(datapath_1_RegisterFile_regfile_mem_14__23_), .C(datapath_1_Instr_21_bF_buf26_), .Y(_3115_) );
OAI21X1 OAI21X1_1873 ( .A(datapath_1_Instr_23_bF_buf10_bF_buf3_), .B(_3114_), .C(_3115_), .Y(_3116_) );
NAND3X1 NAND3X1_1513 ( .A(datapath_1_Instr_22_bF_buf36_), .B(_3116_), .C(_3113_), .Y(_3117_) );
AOI21X1 AOI21X1_805 ( .A(_3110_), .B(_3117_), .C(_1888__bF_buf5), .Y(_3118_) );
OAI21X1 OAI21X1_1874 ( .A(_3118_), .B(_3103_), .C(_1917__bF_buf4), .Y(_3119_) );
NOR2X1 NOR2X1_447 ( .A(datapath_1_Instr_21_bF_buf25_), .B(datapath_1_RegisterFile_regfile_mem_24__23_), .Y(_3120_) );
OAI21X1 OAI21X1_1875 ( .A(datapath_1_RegisterFile_regfile_mem_25__23_), .B(_1890__bF_buf10), .C(_1884__bF_buf9), .Y(_3121_) );
NOR2X1 NOR2X1_448 ( .A(datapath_1_RegisterFile_regfile_mem_27__23_), .B(_1890__bF_buf10), .Y(_3122_) );
OAI21X1 OAI21X1_1876 ( .A(datapath_1_Instr_21_bF_buf24_), .B(datapath_1_RegisterFile_regfile_mem_26__23_), .C(datapath_1_Instr_22_bF_buf35_), .Y(_3123_) );
OAI22X1 OAI22X1_230 ( .A(_3122_), .B(_3123_), .C(_3120_), .D(_3121_), .Y(_3124_) );
NOR2X1 NOR2X1_449 ( .A(datapath_1_Instr_23_bF_buf9_bF_buf3_), .B(_3124_), .Y(_3125_) );
MUX2X1 MUX2X1_234 ( .A(datapath_1_RegisterFile_regfile_mem_29__23_), .B(datapath_1_RegisterFile_regfile_mem_28__23_), .S(datapath_1_Instr_21_bF_buf23_), .Y(_3126_) );
NOR2X1 NOR2X1_450 ( .A(datapath_1_RegisterFile_regfile_mem_31__23_), .B(_1890__bF_buf10), .Y(_3127_) );
OAI21X1 OAI21X1_1877 ( .A(datapath_1_Instr_21_bF_buf22_), .B(datapath_1_RegisterFile_regfile_mem_30__23_), .C(datapath_1_Instr_22_bF_buf34_), .Y(_3128_) );
OAI22X1 OAI22X1_231 ( .A(_3128_), .B(_3127_), .C(datapath_1_Instr_22_bF_buf33_), .D(_3126_), .Y(_3129_) );
OAI21X1 OAI21X1_1878 ( .A(_1885__bF_buf10), .B(_3129_), .C(datapath_1_Instr_24_bF_buf5_), .Y(_3130_) );
INVX1 INVX1_459 ( .A(datapath_1_RegisterFile_regfile_mem_19__23_), .Y(_3131_) );
AOI21X1 AOI21X1_806 ( .A(datapath_1_Instr_23_bF_buf8_bF_buf3_), .B(datapath_1_RegisterFile_regfile_mem_23__23_), .C(_1890__bF_buf10), .Y(_3132_) );
OAI21X1 OAI21X1_1879 ( .A(datapath_1_Instr_23_bF_buf7_bF_buf3_), .B(_3131_), .C(_3132_), .Y(_3133_) );
NAND2X1 NAND2X1_1286 ( .A(datapath_1_RegisterFile_regfile_mem_18__23_), .B(_1885__bF_buf7), .Y(_3134_) );
AOI21X1 AOI21X1_807 ( .A(datapath_1_Instr_23_bF_buf6_bF_buf3_), .B(datapath_1_RegisterFile_regfile_mem_22__23_), .C(datapath_1_Instr_21_bF_buf21_), .Y(_3135_) );
AOI21X1 AOI21X1_808 ( .A(_3134_), .B(_3135_), .C(_1884__bF_buf2), .Y(_3136_) );
INVX1 INVX1_460 ( .A(datapath_1_RegisterFile_regfile_mem_17__23_), .Y(_3137_) );
AOI21X1 AOI21X1_809 ( .A(datapath_1_Instr_23_bF_buf5_bF_buf3_), .B(datapath_1_RegisterFile_regfile_mem_21__23_), .C(_1890__bF_buf10), .Y(_3138_) );
OAI21X1 OAI21X1_1880 ( .A(datapath_1_Instr_23_bF_buf4_bF_buf3_), .B(_3137_), .C(_3138_), .Y(_3139_) );
NAND2X1 NAND2X1_1287 ( .A(datapath_1_RegisterFile_regfile_mem_16__23_), .B(_1885__bF_buf11), .Y(_3140_) );
AOI21X1 AOI21X1_810 ( .A(datapath_1_Instr_23_bF_buf3_bF_buf3_), .B(datapath_1_RegisterFile_regfile_mem_20__23_), .C(datapath_1_Instr_21_bF_buf20_), .Y(_3141_) );
AOI21X1 AOI21X1_811 ( .A(_3140_), .B(_3141_), .C(datapath_1_Instr_22_bF_buf32_), .Y(_3142_) );
AOI22X1 AOI22X1_173 ( .A(_3136_), .B(_3133_), .C(_3139_), .D(_3142_), .Y(_3143_) );
OAI22X1 OAI22X1_232 ( .A(datapath_1_Instr_24_bF_buf4_), .B(_3143_), .C(_3125_), .D(_3130_), .Y(_3144_) );
NAND2X1 NAND2X1_1288 ( .A(datapath_1_Instr_25_bF_buf2_), .B(_3144_), .Y(_3145_) );
AOI22X1 AOI22X1_174 ( .A(_1883__bF_buf0), .B(_1887__bF_buf2), .C(_3119_), .D(_3145_), .Y(datapath_1_RD1_23_) );
NAND2X1 NAND2X1_1289 ( .A(datapath_1_Instr_21_bF_buf19_), .B(datapath_1_RegisterFile_regfile_mem_27__24_), .Y(_3146_) );
NAND2X1 NAND2X1_1290 ( .A(datapath_1_RegisterFile_regfile_mem_26__24_), .B(_1890__bF_buf31), .Y(_3147_) );
NAND3X1 NAND3X1_1514 ( .A(datapath_1_Instr_22_bF_buf31_), .B(_3146_), .C(_3147_), .Y(_3148_) );
NAND2X1 NAND2X1_1291 ( .A(datapath_1_Instr_21_bF_buf18_), .B(datapath_1_RegisterFile_regfile_mem_25__24_), .Y(_3149_) );
AOI21X1 AOI21X1_812 ( .A(_1890__bF_buf31), .B(datapath_1_RegisterFile_regfile_mem_24__24_), .C(datapath_1_Instr_22_bF_buf30_), .Y(_3150_) );
NAND2X1 NAND2X1_1292 ( .A(_3149_), .B(_3150_), .Y(_3151_) );
NAND3X1 NAND3X1_1515 ( .A(_1885__bF_buf7), .B(_3148_), .C(_3151_), .Y(_3152_) );
NAND2X1 NAND2X1_1293 ( .A(datapath_1_Instr_21_bF_buf17_), .B(datapath_1_RegisterFile_regfile_mem_31__24_), .Y(_3153_) );
AOI21X1 AOI21X1_813 ( .A(_1890__bF_buf2), .B(datapath_1_RegisterFile_regfile_mem_30__24_), .C(_1884__bF_buf6), .Y(_3154_) );
NAND2X1 NAND2X1_1294 ( .A(_3153_), .B(_3154_), .Y(_3155_) );
INVX1 INVX1_461 ( .A(datapath_1_RegisterFile_regfile_mem_28__24_), .Y(_3156_) );
AOI21X1 AOI21X1_814 ( .A(datapath_1_Instr_21_bF_buf16_), .B(datapath_1_RegisterFile_regfile_mem_29__24_), .C(datapath_1_Instr_22_bF_buf29_), .Y(_3157_) );
OAI21X1 OAI21X1_1881 ( .A(datapath_1_Instr_21_bF_buf15_), .B(_3156_), .C(_3157_), .Y(_3158_) );
NAND3X1 NAND3X1_1516 ( .A(datapath_1_Instr_23_bF_buf2_bF_buf3_), .B(_3158_), .C(_3155_), .Y(_3159_) );
AOI21X1 AOI21X1_815 ( .A(_3152_), .B(_3159_), .C(_1888__bF_buf3), .Y(_3160_) );
MUX2X1 MUX2X1_235 ( .A(datapath_1_RegisterFile_regfile_mem_18__24_), .B(datapath_1_RegisterFile_regfile_mem_16__24_), .S(datapath_1_Instr_22_bF_buf28_), .Y(_3161_) );
NAND2X1 NAND2X1_1295 ( .A(_1890__bF_buf43), .B(_3161_), .Y(_3162_) );
MUX2X1 MUX2X1_236 ( .A(datapath_1_RegisterFile_regfile_mem_19__24_), .B(datapath_1_RegisterFile_regfile_mem_17__24_), .S(datapath_1_Instr_22_bF_buf27_), .Y(_3163_) );
NAND2X1 NAND2X1_1296 ( .A(datapath_1_Instr_21_bF_buf14_), .B(_3163_), .Y(_3164_) );
NAND3X1 NAND3X1_1517 ( .A(_1885__bF_buf3), .B(_3162_), .C(_3164_), .Y(_3165_) );
MUX2X1 MUX2X1_237 ( .A(datapath_1_RegisterFile_regfile_mem_22__24_), .B(datapath_1_RegisterFile_regfile_mem_20__24_), .S(datapath_1_Instr_22_bF_buf26_), .Y(_3166_) );
NAND2X1 NAND2X1_1297 ( .A(_1890__bF_buf2), .B(_3166_), .Y(_3167_) );
MUX2X1 MUX2X1_238 ( .A(datapath_1_RegisterFile_regfile_mem_23__24_), .B(datapath_1_RegisterFile_regfile_mem_21__24_), .S(datapath_1_Instr_22_bF_buf25_), .Y(_3168_) );
NAND2X1 NAND2X1_1298 ( .A(datapath_1_Instr_21_bF_buf13_), .B(_3168_), .Y(_3169_) );
NAND3X1 NAND3X1_1518 ( .A(datapath_1_Instr_23_bF_buf1_), .B(_3167_), .C(_3169_), .Y(_3170_) );
AOI21X1 AOI21X1_816 ( .A(_3165_), .B(_3170_), .C(datapath_1_Instr_24_bF_buf3_), .Y(_3171_) );
OAI21X1 OAI21X1_1882 ( .A(_3171_), .B(_3160_), .C(datapath_1_Instr_25_bF_buf1_), .Y(_3172_) );
MUX2X1 MUX2X1_239 ( .A(datapath_1_RegisterFile_regfile_mem_9__24_), .B(datapath_1_RegisterFile_regfile_mem_8__24_), .S(datapath_1_Instr_21_bF_buf12_), .Y(_3173_) );
NOR2X1 NOR2X1_451 ( .A(datapath_1_RegisterFile_regfile_mem_11__24_), .B(_1890__bF_buf0), .Y(_3174_) );
OAI21X1 OAI21X1_1883 ( .A(datapath_1_Instr_21_bF_buf11_), .B(datapath_1_RegisterFile_regfile_mem_10__24_), .C(datapath_1_Instr_22_bF_buf24_), .Y(_3175_) );
OAI22X1 OAI22X1_233 ( .A(_3175_), .B(_3174_), .C(datapath_1_Instr_22_bF_buf23_), .D(_3173_), .Y(_3176_) );
INVX1 INVX1_462 ( .A(datapath_1_RegisterFile_regfile_mem_15__24_), .Y(_3177_) );
AOI21X1 AOI21X1_817 ( .A(_1890__bF_buf23), .B(datapath_1_RegisterFile_regfile_mem_14__24_), .C(_1884__bF_buf7), .Y(_3178_) );
OAI21X1 OAI21X1_1884 ( .A(_1890__bF_buf23), .B(_3177_), .C(_3178_), .Y(_3179_) );
NAND2X1 NAND2X1_1299 ( .A(datapath_1_RegisterFile_regfile_mem_12__24_), .B(_1890__bF_buf0), .Y(_3180_) );
AOI21X1 AOI21X1_818 ( .A(datapath_1_Instr_21_bF_buf10_), .B(datapath_1_RegisterFile_regfile_mem_13__24_), .C(datapath_1_Instr_22_bF_buf22_), .Y(_3181_) );
AOI21X1 AOI21X1_819 ( .A(_3180_), .B(_3181_), .C(_1885__bF_buf8), .Y(_3182_) );
AOI22X1 AOI22X1_175 ( .A(_3179_), .B(_3182_), .C(_1885__bF_buf8), .D(_3176_), .Y(_3183_) );
NOR2X1 NOR2X1_452 ( .A(datapath_1_Instr_21_bF_buf9_), .B(datapath_1_RegisterFile_regfile_mem_0__24_), .Y(_3184_) );
OAI21X1 OAI21X1_1885 ( .A(datapath_1_RegisterFile_regfile_mem_1__24_), .B(_1890__bF_buf47), .C(_1884__bF_buf7), .Y(_3185_) );
NOR2X1 NOR2X1_453 ( .A(datapath_1_RegisterFile_regfile_mem_3__24_), .B(_1890__bF_buf47), .Y(_3186_) );
OAI21X1 OAI21X1_1886 ( .A(datapath_1_Instr_21_bF_buf8_), .B(datapath_1_RegisterFile_regfile_mem_2__24_), .C(datapath_1_Instr_22_bF_buf21_), .Y(_3187_) );
OAI22X1 OAI22X1_234 ( .A(_3186_), .B(_3187_), .C(_3184_), .D(_3185_), .Y(_3188_) );
NOR2X1 NOR2X1_454 ( .A(datapath_1_Instr_23_bF_buf0_), .B(_3188_), .Y(_3189_) );
MUX2X1 MUX2X1_240 ( .A(datapath_1_RegisterFile_regfile_mem_5__24_), .B(datapath_1_RegisterFile_regfile_mem_4__24_), .S(datapath_1_Instr_21_bF_buf7_), .Y(_3190_) );
NOR2X1 NOR2X1_455 ( .A(datapath_1_RegisterFile_regfile_mem_7__24_), .B(_1890__bF_buf29), .Y(_3191_) );
OAI21X1 OAI21X1_1887 ( .A(datapath_1_Instr_21_bF_buf6_), .B(datapath_1_RegisterFile_regfile_mem_6__24_), .C(datapath_1_Instr_22_bF_buf20_), .Y(_3192_) );
OAI22X1 OAI22X1_235 ( .A(_3192_), .B(_3191_), .C(datapath_1_Instr_22_bF_buf19_), .D(_3190_), .Y(_3193_) );
OAI21X1 OAI21X1_1888 ( .A(_1885__bF_buf8), .B(_3193_), .C(_1888__bF_buf4), .Y(_3194_) );
OAI22X1 OAI22X1_236 ( .A(_1888__bF_buf4), .B(_3183_), .C(_3189_), .D(_3194_), .Y(_3195_) );
NAND2X1 NAND2X1_1300 ( .A(_1917__bF_buf1), .B(_3195_), .Y(_3196_) );
AOI22X1 AOI22X1_176 ( .A(_1883__bF_buf3), .B(_1887__bF_buf1), .C(_3172_), .D(_3196_), .Y(datapath_1_RD1_24_) );
MUX2X1 MUX2X1_241 ( .A(datapath_1_RegisterFile_regfile_mem_9__25_), .B(datapath_1_RegisterFile_regfile_mem_8__25_), .S(datapath_1_Instr_21_bF_buf5_), .Y(_3197_) );
NOR2X1 NOR2X1_456 ( .A(datapath_1_RegisterFile_regfile_mem_11__25_), .B(_1890__bF_buf18), .Y(_3198_) );
OAI21X1 OAI21X1_1889 ( .A(datapath_1_Instr_21_bF_buf4_), .B(datapath_1_RegisterFile_regfile_mem_10__25_), .C(datapath_1_Instr_22_bF_buf18_), .Y(_3199_) );
OAI22X1 OAI22X1_237 ( .A(_3199_), .B(_3198_), .C(datapath_1_Instr_22_bF_buf17_), .D(_3197_), .Y(_3200_) );
INVX1 INVX1_463 ( .A(datapath_1_RegisterFile_regfile_mem_15__25_), .Y(_3201_) );
AOI21X1 AOI21X1_820 ( .A(_1890__bF_buf16), .B(datapath_1_RegisterFile_regfile_mem_14__25_), .C(_1884__bF_buf0), .Y(_3202_) );
OAI21X1 OAI21X1_1890 ( .A(_1890__bF_buf18), .B(_3201_), .C(_3202_), .Y(_3203_) );
NAND2X1 NAND2X1_1301 ( .A(datapath_1_RegisterFile_regfile_mem_12__25_), .B(_1890__bF_buf18), .Y(_3204_) );
AOI21X1 AOI21X1_821 ( .A(datapath_1_Instr_21_bF_buf3_), .B(datapath_1_RegisterFile_regfile_mem_13__25_), .C(datapath_1_Instr_22_bF_buf16_), .Y(_3205_) );
AOI21X1 AOI21X1_822 ( .A(_3204_), .B(_3205_), .C(_1885__bF_buf2), .Y(_3206_) );
AOI22X1 AOI22X1_177 ( .A(_3203_), .B(_3206_), .C(_1885__bF_buf2), .D(_3200_), .Y(_3207_) );
NOR2X1 NOR2X1_457 ( .A(datapath_1_Instr_21_bF_buf2_), .B(datapath_1_RegisterFile_regfile_mem_0__25_), .Y(_3208_) );
OAI21X1 OAI21X1_1891 ( .A(datapath_1_RegisterFile_regfile_mem_1__25_), .B(_1890__bF_buf8), .C(_1884__bF_buf4), .Y(_3209_) );
NOR2X1 NOR2X1_458 ( .A(datapath_1_RegisterFile_regfile_mem_3__25_), .B(_1890__bF_buf44), .Y(_3210_) );
OAI21X1 OAI21X1_1892 ( .A(datapath_1_Instr_21_bF_buf1_), .B(datapath_1_RegisterFile_regfile_mem_2__25_), .C(datapath_1_Instr_22_bF_buf15_), .Y(_3211_) );
OAI22X1 OAI22X1_238 ( .A(_3210_), .B(_3211_), .C(_3208_), .D(_3209_), .Y(_3212_) );
NOR2X1 NOR2X1_459 ( .A(datapath_1_Instr_23_bF_buf15_bF_buf2_), .B(_3212_), .Y(_3213_) );
MUX2X1 MUX2X1_242 ( .A(datapath_1_RegisterFile_regfile_mem_5__25_), .B(datapath_1_RegisterFile_regfile_mem_4__25_), .S(datapath_1_Instr_21_bF_buf0_), .Y(_3214_) );
NOR2X1 NOR2X1_460 ( .A(datapath_1_RegisterFile_regfile_mem_7__25_), .B(_1890__bF_buf44), .Y(_3215_) );
OAI21X1 OAI21X1_1893 ( .A(datapath_1_Instr_21_bF_buf55_), .B(datapath_1_RegisterFile_regfile_mem_6__25_), .C(datapath_1_Instr_22_bF_buf14_), .Y(_3216_) );
OAI22X1 OAI22X1_239 ( .A(_3216_), .B(_3215_), .C(datapath_1_Instr_22_bF_buf13_), .D(_3214_), .Y(_3217_) );
OAI21X1 OAI21X1_1894 ( .A(_1885__bF_buf10), .B(_3217_), .C(_1888__bF_buf3), .Y(_3218_) );
OAI22X1 OAI22X1_240 ( .A(_1888__bF_buf3), .B(_3207_), .C(_3213_), .D(_3218_), .Y(_3219_) );
NAND2X1 NAND2X1_1302 ( .A(_1917__bF_buf2), .B(_3219_), .Y(_3220_) );
INVX1 INVX1_464 ( .A(datapath_1_RegisterFile_regfile_mem_27__25_), .Y(_3221_) );
AOI21X1 AOI21X1_823 ( .A(datapath_1_Instr_23_bF_buf14_bF_buf2_), .B(datapath_1_RegisterFile_regfile_mem_31__25_), .C(_1890__bF_buf11), .Y(_3222_) );
OAI21X1 OAI21X1_1895 ( .A(datapath_1_Instr_23_bF_buf13_bF_buf2_), .B(_3221_), .C(_3222_), .Y(_3223_) );
INVX1 INVX1_465 ( .A(datapath_1_RegisterFile_regfile_mem_26__25_), .Y(_3224_) );
AOI21X1 AOI21X1_824 ( .A(datapath_1_Instr_23_bF_buf12_bF_buf2_), .B(datapath_1_RegisterFile_regfile_mem_30__25_), .C(datapath_1_Instr_21_bF_buf54_), .Y(_3225_) );
OAI21X1 OAI21X1_1896 ( .A(datapath_1_Instr_23_bF_buf11_bF_buf2_), .B(_3224_), .C(_3225_), .Y(_3226_) );
NAND3X1 NAND3X1_1519 ( .A(datapath_1_Instr_22_bF_buf12_), .B(_3226_), .C(_3223_), .Y(_3227_) );
INVX1 INVX1_466 ( .A(datapath_1_RegisterFile_regfile_mem_25__25_), .Y(_3228_) );
AOI21X1 AOI21X1_825 ( .A(datapath_1_Instr_23_bF_buf10_bF_buf2_), .B(datapath_1_RegisterFile_regfile_mem_29__25_), .C(_1890__bF_buf11), .Y(_3229_) );
OAI21X1 OAI21X1_1897 ( .A(datapath_1_Instr_23_bF_buf9_bF_buf2_), .B(_3228_), .C(_3229_), .Y(_3230_) );
INVX1 INVX1_467 ( .A(datapath_1_RegisterFile_regfile_mem_24__25_), .Y(_3231_) );
AOI21X1 AOI21X1_826 ( .A(datapath_1_Instr_23_bF_buf8_bF_buf2_), .B(datapath_1_RegisterFile_regfile_mem_28__25_), .C(datapath_1_Instr_21_bF_buf53_), .Y(_3232_) );
OAI21X1 OAI21X1_1898 ( .A(datapath_1_Instr_23_bF_buf7_bF_buf2_), .B(_3231_), .C(_3232_), .Y(_3233_) );
NAND3X1 NAND3X1_1520 ( .A(_1884__bF_buf2), .B(_3233_), .C(_3230_), .Y(_3234_) );
AOI21X1 AOI21X1_827 ( .A(_3227_), .B(_3234_), .C(_1888__bF_buf0), .Y(_3235_) );
MUX2X1 MUX2X1_243 ( .A(datapath_1_RegisterFile_regfile_mem_18__25_), .B(datapath_1_RegisterFile_regfile_mem_16__25_), .S(datapath_1_Instr_22_bF_buf11_), .Y(_3236_) );
NAND2X1 NAND2X1_1303 ( .A(_1890__bF_buf43), .B(_3236_), .Y(_3237_) );
MUX2X1 MUX2X1_244 ( .A(datapath_1_RegisterFile_regfile_mem_19__25_), .B(datapath_1_RegisterFile_regfile_mem_17__25_), .S(datapath_1_Instr_22_bF_buf10_), .Y(_3238_) );
NAND2X1 NAND2X1_1304 ( .A(datapath_1_Instr_21_bF_buf52_), .B(_3238_), .Y(_3239_) );
NAND3X1 NAND3X1_1521 ( .A(_1885__bF_buf3), .B(_3237_), .C(_3239_), .Y(_3240_) );
MUX2X1 MUX2X1_245 ( .A(datapath_1_RegisterFile_regfile_mem_22__25_), .B(datapath_1_RegisterFile_regfile_mem_20__25_), .S(datapath_1_Instr_22_bF_buf9_), .Y(_3241_) );
NAND2X1 NAND2X1_1305 ( .A(_1890__bF_buf32), .B(_3241_), .Y(_3242_) );
MUX2X1 MUX2X1_246 ( .A(datapath_1_RegisterFile_regfile_mem_23__25_), .B(datapath_1_RegisterFile_regfile_mem_21__25_), .S(datapath_1_Instr_22_bF_buf8_), .Y(_3243_) );
NAND2X1 NAND2X1_1306 ( .A(datapath_1_Instr_21_bF_buf51_), .B(_3243_), .Y(_3244_) );
NAND3X1 NAND3X1_1522 ( .A(datapath_1_Instr_23_bF_buf6_bF_buf2_), .B(_3242_), .C(_3244_), .Y(_3245_) );
AOI21X1 AOI21X1_828 ( .A(_3240_), .B(_3245_), .C(datapath_1_Instr_24_bF_buf2_), .Y(_3246_) );
OAI21X1 OAI21X1_1899 ( .A(_3235_), .B(_3246_), .C(datapath_1_Instr_25_bF_buf0_), .Y(_3247_) );
AOI22X1 AOI22X1_178 ( .A(_1883__bF_buf1), .B(_1887__bF_buf0), .C(_3247_), .D(_3220_), .Y(datapath_1_RD1_25_) );
NAND2X1 NAND2X1_1307 ( .A(datapath_1_Instr_21_bF_buf50_), .B(datapath_1_RegisterFile_regfile_mem_27__26_), .Y(_3248_) );
NAND2X1 NAND2X1_1308 ( .A(datapath_1_RegisterFile_regfile_mem_26__26_), .B(_1890__bF_buf40), .Y(_3249_) );
NAND3X1 NAND3X1_1523 ( .A(datapath_1_Instr_22_bF_buf7_), .B(_3248_), .C(_3249_), .Y(_3250_) );
NAND2X1 NAND2X1_1309 ( .A(datapath_1_Instr_21_bF_buf49_), .B(datapath_1_RegisterFile_regfile_mem_25__26_), .Y(_3251_) );
AOI21X1 AOI21X1_829 ( .A(_1890__bF_buf1), .B(datapath_1_RegisterFile_regfile_mem_24__26_), .C(datapath_1_Instr_22_bF_buf6_), .Y(_3252_) );
NAND2X1 NAND2X1_1310 ( .A(_3251_), .B(_3252_), .Y(_3253_) );
NAND3X1 NAND3X1_1524 ( .A(_1885__bF_buf9), .B(_3250_), .C(_3253_), .Y(_3254_) );
NAND2X1 NAND2X1_1311 ( .A(datapath_1_Instr_21_bF_buf48_), .B(datapath_1_RegisterFile_regfile_mem_31__26_), .Y(_3255_) );
AOI21X1 AOI21X1_830 ( .A(_1890__bF_buf9), .B(datapath_1_RegisterFile_regfile_mem_30__26_), .C(_1884__bF_buf9), .Y(_3256_) );
NAND2X1 NAND2X1_1312 ( .A(_3255_), .B(_3256_), .Y(_3257_) );
INVX1 INVX1_468 ( .A(datapath_1_RegisterFile_regfile_mem_28__26_), .Y(_3258_) );
AOI21X1 AOI21X1_831 ( .A(datapath_1_Instr_21_bF_buf47_), .B(datapath_1_RegisterFile_regfile_mem_29__26_), .C(datapath_1_Instr_22_bF_buf5_), .Y(_3259_) );
OAI21X1 OAI21X1_1900 ( .A(datapath_1_Instr_21_bF_buf46_), .B(_3258_), .C(_3259_), .Y(_3260_) );
NAND3X1 NAND3X1_1525 ( .A(datapath_1_Instr_23_bF_buf5_bF_buf2_), .B(_3260_), .C(_3257_), .Y(_3261_) );
AOI21X1 AOI21X1_832 ( .A(_3254_), .B(_3261_), .C(_1888__bF_buf1), .Y(_3262_) );
MUX2X1 MUX2X1_247 ( .A(datapath_1_RegisterFile_regfile_mem_18__26_), .B(datapath_1_RegisterFile_regfile_mem_16__26_), .S(datapath_1_Instr_22_bF_buf4_), .Y(_3263_) );
NAND2X1 NAND2X1_1313 ( .A(_1890__bF_buf9), .B(_3263_), .Y(_3264_) );
MUX2X1 MUX2X1_248 ( .A(datapath_1_RegisterFile_regfile_mem_19__26_), .B(datapath_1_RegisterFile_regfile_mem_17__26_), .S(datapath_1_Instr_22_bF_buf3_), .Y(_3265_) );
NAND2X1 NAND2X1_1314 ( .A(datapath_1_Instr_21_bF_buf45_), .B(_3265_), .Y(_3266_) );
NAND3X1 NAND3X1_1526 ( .A(_1885__bF_buf9), .B(_3264_), .C(_3266_), .Y(_3267_) );
MUX2X1 MUX2X1_249 ( .A(datapath_1_RegisterFile_regfile_mem_22__26_), .B(datapath_1_RegisterFile_regfile_mem_20__26_), .S(datapath_1_Instr_22_bF_buf2_), .Y(_3268_) );
NAND2X1 NAND2X1_1315 ( .A(_1890__bF_buf37), .B(_3268_), .Y(_3269_) );
MUX2X1 MUX2X1_250 ( .A(datapath_1_RegisterFile_regfile_mem_23__26_), .B(datapath_1_RegisterFile_regfile_mem_21__26_), .S(datapath_1_Instr_22_bF_buf1_), .Y(_3270_) );
NAND2X1 NAND2X1_1316 ( .A(datapath_1_Instr_21_bF_buf44_), .B(_3270_), .Y(_3271_) );
NAND3X1 NAND3X1_1527 ( .A(datapath_1_Instr_23_bF_buf4_bF_buf2_), .B(_3269_), .C(_3271_), .Y(_3272_) );
AOI21X1 AOI21X1_833 ( .A(_3267_), .B(_3272_), .C(datapath_1_Instr_24_bF_buf1_), .Y(_3273_) );
OAI21X1 OAI21X1_1901 ( .A(_3273_), .B(_3262_), .C(datapath_1_Instr_25_bF_buf5_), .Y(_3274_) );
INVX1 INVX1_469 ( .A(datapath_1_RegisterFile_regfile_mem_9__26_), .Y(_3275_) );
AOI21X1 AOI21X1_834 ( .A(datapath_1_Instr_23_bF_buf3_bF_buf2_), .B(datapath_1_RegisterFile_regfile_mem_13__26_), .C(_1890__bF_buf5), .Y(_3276_) );
OAI21X1 OAI21X1_1902 ( .A(datapath_1_Instr_23_bF_buf2_bF_buf2_), .B(_3275_), .C(_3276_), .Y(_3277_) );
INVX1 INVX1_470 ( .A(datapath_1_RegisterFile_regfile_mem_8__26_), .Y(_3278_) );
AOI21X1 AOI21X1_835 ( .A(datapath_1_Instr_23_bF_buf1_), .B(datapath_1_RegisterFile_regfile_mem_12__26_), .C(datapath_1_Instr_21_bF_buf43_), .Y(_3279_) );
OAI21X1 OAI21X1_1903 ( .A(datapath_1_Instr_23_bF_buf0_), .B(_3278_), .C(_3279_), .Y(_3280_) );
NAND3X1 NAND3X1_1528 ( .A(_1884__bF_buf5), .B(_3280_), .C(_3277_), .Y(_3281_) );
INVX1 INVX1_471 ( .A(datapath_1_RegisterFile_regfile_mem_11__26_), .Y(_3282_) );
AOI21X1 AOI21X1_836 ( .A(datapath_1_Instr_23_bF_buf15_bF_buf1_), .B(datapath_1_RegisterFile_regfile_mem_15__26_), .C(_1890__bF_buf5), .Y(_3283_) );
OAI21X1 OAI21X1_1904 ( .A(datapath_1_Instr_23_bF_buf14_bF_buf1_), .B(_3282_), .C(_3283_), .Y(_3284_) );
INVX1 INVX1_472 ( .A(datapath_1_RegisterFile_regfile_mem_10__26_), .Y(_3285_) );
AOI21X1 AOI21X1_837 ( .A(datapath_1_Instr_23_bF_buf13_bF_buf1_), .B(datapath_1_RegisterFile_regfile_mem_14__26_), .C(datapath_1_Instr_21_bF_buf42_), .Y(_3286_) );
OAI21X1 OAI21X1_1905 ( .A(datapath_1_Instr_23_bF_buf12_bF_buf1_), .B(_3285_), .C(_3286_), .Y(_3287_) );
NAND3X1 NAND3X1_1529 ( .A(datapath_1_Instr_22_bF_buf0_), .B(_3287_), .C(_3284_), .Y(_3288_) );
AOI21X1 AOI21X1_838 ( .A(_3281_), .B(_3288_), .C(_1888__bF_buf5), .Y(_3289_) );
MUX2X1 MUX2X1_251 ( .A(datapath_1_RegisterFile_regfile_mem_1__26_), .B(datapath_1_RegisterFile_regfile_mem_0__26_), .S(datapath_1_Instr_21_bF_buf41_), .Y(_3290_) );
NOR2X1 NOR2X1_461 ( .A(datapath_1_RegisterFile_regfile_mem_3__26_), .B(_1890__bF_buf30), .Y(_3291_) );
OAI21X1 OAI21X1_1906 ( .A(datapath_1_Instr_21_bF_buf40_), .B(datapath_1_RegisterFile_regfile_mem_2__26_), .C(datapath_1_Instr_22_bF_buf50_), .Y(_3292_) );
OAI22X1 OAI22X1_241 ( .A(_3292_), .B(_3291_), .C(datapath_1_Instr_22_bF_buf49_), .D(_3290_), .Y(_3293_) );
NAND2X1 NAND2X1_1317 ( .A(_1885__bF_buf4), .B(_3293_), .Y(_3294_) );
MUX2X1 MUX2X1_252 ( .A(datapath_1_RegisterFile_regfile_mem_5__26_), .B(datapath_1_RegisterFile_regfile_mem_4__26_), .S(datapath_1_Instr_21_bF_buf39_), .Y(_3295_) );
NOR2X1 NOR2X1_462 ( .A(datapath_1_RegisterFile_regfile_mem_7__26_), .B(_1890__bF_buf30), .Y(_3296_) );
OAI21X1 OAI21X1_1907 ( .A(datapath_1_Instr_21_bF_buf38_), .B(datapath_1_RegisterFile_regfile_mem_6__26_), .C(datapath_1_Instr_22_bF_buf48_), .Y(_3297_) );
OAI22X1 OAI22X1_242 ( .A(_3297_), .B(_3296_), .C(datapath_1_Instr_22_bF_buf47_), .D(_3295_), .Y(_3298_) );
NAND2X1 NAND2X1_1318 ( .A(datapath_1_Instr_23_bF_buf11_bF_buf1_), .B(_3298_), .Y(_3299_) );
AOI21X1 AOI21X1_839 ( .A(_3294_), .B(_3299_), .C(datapath_1_Instr_24_bF_buf0_), .Y(_3300_) );
OAI21X1 OAI21X1_1908 ( .A(_3289_), .B(_3300_), .C(_1917__bF_buf4), .Y(_3301_) );
AOI22X1 AOI22X1_179 ( .A(_1883__bF_buf2), .B(_1887__bF_buf4), .C(_3274_), .D(_3301_), .Y(datapath_1_RD1_26_) );
NAND2X1 NAND2X1_1319 ( .A(datapath_1_Instr_21_bF_buf37_), .B(datapath_1_RegisterFile_regfile_mem_27__27_), .Y(_3302_) );
NAND2X1 NAND2X1_1320 ( .A(datapath_1_RegisterFile_regfile_mem_26__27_), .B(_1890__bF_buf34), .Y(_3303_) );
NAND3X1 NAND3X1_1530 ( .A(datapath_1_Instr_22_bF_buf46_), .B(_3302_), .C(_3303_), .Y(_3304_) );
NAND2X1 NAND2X1_1321 ( .A(datapath_1_Instr_21_bF_buf36_), .B(datapath_1_RegisterFile_regfile_mem_25__27_), .Y(_3305_) );
AOI21X1 AOI21X1_840 ( .A(_1890__bF_buf34), .B(datapath_1_RegisterFile_regfile_mem_24__27_), .C(datapath_1_Instr_22_bF_buf45_), .Y(_3306_) );
NAND2X1 NAND2X1_1322 ( .A(_3305_), .B(_3306_), .Y(_3307_) );
NAND3X1 NAND3X1_1531 ( .A(_1885__bF_buf6), .B(_3304_), .C(_3307_), .Y(_3308_) );
NAND2X1 NAND2X1_1323 ( .A(datapath_1_Instr_21_bF_buf35_), .B(datapath_1_RegisterFile_regfile_mem_31__27_), .Y(_3309_) );
AOI21X1 AOI21X1_841 ( .A(_1890__bF_buf34), .B(datapath_1_RegisterFile_regfile_mem_30__27_), .C(_1884__bF_buf3), .Y(_3310_) );
NAND2X1 NAND2X1_1324 ( .A(_3309_), .B(_3310_), .Y(_3311_) );
INVX1 INVX1_473 ( .A(datapath_1_RegisterFile_regfile_mem_28__27_), .Y(_3312_) );
AOI21X1 AOI21X1_842 ( .A(datapath_1_Instr_21_bF_buf34_), .B(datapath_1_RegisterFile_regfile_mem_29__27_), .C(datapath_1_Instr_22_bF_buf44_), .Y(_3313_) );
OAI21X1 OAI21X1_1909 ( .A(datapath_1_Instr_21_bF_buf33_), .B(_3312_), .C(_3313_), .Y(_3314_) );
NAND3X1 NAND3X1_1532 ( .A(datapath_1_Instr_23_bF_buf10_bF_buf1_), .B(_3314_), .C(_3311_), .Y(_3315_) );
AOI21X1 AOI21X1_843 ( .A(_3308_), .B(_3315_), .C(_1888__bF_buf1), .Y(_3316_) );
MUX2X1 MUX2X1_253 ( .A(datapath_1_RegisterFile_regfile_mem_18__27_), .B(datapath_1_RegisterFile_regfile_mem_16__27_), .S(datapath_1_Instr_22_bF_buf43_), .Y(_3317_) );
NAND2X1 NAND2X1_1325 ( .A(_1890__bF_buf39), .B(_3317_), .Y(_3318_) );
MUX2X1 MUX2X1_254 ( .A(datapath_1_RegisterFile_regfile_mem_19__27_), .B(datapath_1_RegisterFile_regfile_mem_17__27_), .S(datapath_1_Instr_22_bF_buf42_), .Y(_3319_) );
NAND2X1 NAND2X1_1326 ( .A(datapath_1_Instr_21_bF_buf32_), .B(_3319_), .Y(_3320_) );
NAND3X1 NAND3X1_1533 ( .A(_1885__bF_buf6), .B(_3318_), .C(_3320_), .Y(_3321_) );
MUX2X1 MUX2X1_255 ( .A(datapath_1_RegisterFile_regfile_mem_22__27_), .B(datapath_1_RegisterFile_regfile_mem_20__27_), .S(datapath_1_Instr_22_bF_buf41_), .Y(_3322_) );
NAND2X1 NAND2X1_1327 ( .A(_1890__bF_buf39), .B(_3322_), .Y(_3323_) );
MUX2X1 MUX2X1_256 ( .A(datapath_1_RegisterFile_regfile_mem_23__27_), .B(datapath_1_RegisterFile_regfile_mem_21__27_), .S(datapath_1_Instr_22_bF_buf40_), .Y(_3324_) );
NAND2X1 NAND2X1_1328 ( .A(datapath_1_Instr_21_bF_buf31_), .B(_3324_), .Y(_3325_) );
NAND3X1 NAND3X1_1534 ( .A(datapath_1_Instr_23_bF_buf9_bF_buf1_), .B(_3323_), .C(_3325_), .Y(_3326_) );
AOI21X1 AOI21X1_844 ( .A(_3321_), .B(_3326_), .C(datapath_1_Instr_24_bF_buf6_), .Y(_3327_) );
OAI21X1 OAI21X1_1910 ( .A(_3327_), .B(_3316_), .C(datapath_1_Instr_25_bF_buf4_), .Y(_3328_) );
MUX2X1 MUX2X1_257 ( .A(datapath_1_RegisterFile_regfile_mem_9__27_), .B(datapath_1_RegisterFile_regfile_mem_8__27_), .S(datapath_1_Instr_21_bF_buf30_), .Y(_3329_) );
NOR2X1 NOR2X1_463 ( .A(datapath_1_RegisterFile_regfile_mem_11__27_), .B(_1890__bF_buf14), .Y(_3330_) );
OAI21X1 OAI21X1_1911 ( .A(datapath_1_Instr_21_bF_buf29_), .B(datapath_1_RegisterFile_regfile_mem_10__27_), .C(datapath_1_Instr_22_bF_buf39_), .Y(_3331_) );
OAI22X1 OAI22X1_243 ( .A(_3331_), .B(_3330_), .C(datapath_1_Instr_22_bF_buf38_), .D(_3329_), .Y(_3332_) );
INVX1 INVX1_474 ( .A(datapath_1_RegisterFile_regfile_mem_15__27_), .Y(_3333_) );
AOI21X1 AOI21X1_845 ( .A(_1890__bF_buf14), .B(datapath_1_RegisterFile_regfile_mem_14__27_), .C(_1884__bF_buf1), .Y(_3334_) );
OAI21X1 OAI21X1_1912 ( .A(_1890__bF_buf14), .B(_3333_), .C(_3334_), .Y(_3335_) );
NAND2X1 NAND2X1_1329 ( .A(datapath_1_RegisterFile_regfile_mem_12__27_), .B(_1890__bF_buf45), .Y(_3336_) );
AOI21X1 AOI21X1_846 ( .A(datapath_1_Instr_21_bF_buf28_), .B(datapath_1_RegisterFile_regfile_mem_13__27_), .C(datapath_1_Instr_22_bF_buf37_), .Y(_3337_) );
AOI21X1 AOI21X1_847 ( .A(_3336_), .B(_3337_), .C(_1885__bF_buf5), .Y(_3338_) );
AOI22X1 AOI22X1_180 ( .A(_3335_), .B(_3338_), .C(_1885__bF_buf5), .D(_3332_), .Y(_3339_) );
NOR2X1 NOR2X1_464 ( .A(datapath_1_Instr_21_bF_buf27_), .B(datapath_1_RegisterFile_regfile_mem_0__27_), .Y(_3340_) );
OAI21X1 OAI21X1_1913 ( .A(datapath_1_RegisterFile_regfile_mem_1__27_), .B(_1890__bF_buf14), .C(_1884__bF_buf1), .Y(_3341_) );
NOR2X1 NOR2X1_465 ( .A(datapath_1_RegisterFile_regfile_mem_3__27_), .B(_1890__bF_buf14), .Y(_3342_) );
OAI21X1 OAI21X1_1914 ( .A(datapath_1_Instr_21_bF_buf26_), .B(datapath_1_RegisterFile_regfile_mem_2__27_), .C(datapath_1_Instr_22_bF_buf36_), .Y(_3343_) );
OAI22X1 OAI22X1_244 ( .A(_3342_), .B(_3343_), .C(_3340_), .D(_3341_), .Y(_3344_) );
NOR2X1 NOR2X1_466 ( .A(datapath_1_Instr_23_bF_buf8_bF_buf1_), .B(_3344_), .Y(_3345_) );
MUX2X1 MUX2X1_258 ( .A(datapath_1_RegisterFile_regfile_mem_5__27_), .B(datapath_1_RegisterFile_regfile_mem_4__27_), .S(datapath_1_Instr_21_bF_buf25_), .Y(_3346_) );
NOR2X1 NOR2X1_467 ( .A(datapath_1_RegisterFile_regfile_mem_7__27_), .B(_1890__bF_buf14), .Y(_3347_) );
OAI21X1 OAI21X1_1915 ( .A(datapath_1_Instr_21_bF_buf24_), .B(datapath_1_RegisterFile_regfile_mem_6__27_), .C(datapath_1_Instr_22_bF_buf35_), .Y(_3348_) );
OAI22X1 OAI22X1_245 ( .A(_3348_), .B(_3347_), .C(datapath_1_Instr_22_bF_buf34_), .D(_3346_), .Y(_3349_) );
OAI21X1 OAI21X1_1916 ( .A(_1885__bF_buf5), .B(_3349_), .C(_1888__bF_buf5), .Y(_3350_) );
OAI22X1 OAI22X1_246 ( .A(_1888__bF_buf5), .B(_3339_), .C(_3345_), .D(_3350_), .Y(_3351_) );
NAND2X1 NAND2X1_1330 ( .A(_1917__bF_buf0), .B(_3351_), .Y(_3352_) );
AOI22X1 AOI22X1_181 ( .A(_1883__bF_buf4), .B(_1887__bF_buf3), .C(_3328_), .D(_3352_), .Y(datapath_1_RD1_27_) );
NAND2X1 NAND2X1_1331 ( .A(datapath_1_Instr_21_bF_buf23_), .B(datapath_1_RegisterFile_regfile_mem_27__28_), .Y(_3353_) );
NAND2X1 NAND2X1_1332 ( .A(datapath_1_RegisterFile_regfile_mem_26__28_), .B(_1890__bF_buf29), .Y(_3354_) );
NAND3X1 NAND3X1_1535 ( .A(datapath_1_Instr_22_bF_buf33_), .B(_3353_), .C(_3354_), .Y(_3355_) );
NAND2X1 NAND2X1_1333 ( .A(datapath_1_Instr_21_bF_buf22_), .B(datapath_1_RegisterFile_regfile_mem_25__28_), .Y(_3356_) );
AOI21X1 AOI21X1_848 ( .A(_1890__bF_buf29), .B(datapath_1_RegisterFile_regfile_mem_24__28_), .C(datapath_1_Instr_22_bF_buf32_), .Y(_3357_) );
NAND2X1 NAND2X1_1334 ( .A(_3356_), .B(_3357_), .Y(_3358_) );
NAND3X1 NAND3X1_1536 ( .A(_1885__bF_buf10), .B(_3355_), .C(_3358_), .Y(_3359_) );
NAND2X1 NAND2X1_1335 ( .A(datapath_1_Instr_21_bF_buf21_), .B(datapath_1_RegisterFile_regfile_mem_31__28_), .Y(_3360_) );
AOI21X1 AOI21X1_849 ( .A(_1890__bF_buf19), .B(datapath_1_RegisterFile_regfile_mem_30__28_), .C(_1884__bF_buf6), .Y(_3361_) );
NAND2X1 NAND2X1_1336 ( .A(_3360_), .B(_3361_), .Y(_3362_) );
INVX1 INVX1_475 ( .A(datapath_1_RegisterFile_regfile_mem_28__28_), .Y(_3363_) );
AOI21X1 AOI21X1_850 ( .A(datapath_1_Instr_21_bF_buf20_), .B(datapath_1_RegisterFile_regfile_mem_29__28_), .C(datapath_1_Instr_22_bF_buf31_), .Y(_3364_) );
OAI21X1 OAI21X1_1917 ( .A(datapath_1_Instr_21_bF_buf19_), .B(_3363_), .C(_3364_), .Y(_3365_) );
NAND3X1 NAND3X1_1537 ( .A(datapath_1_Instr_23_bF_buf7_bF_buf1_), .B(_3365_), .C(_3362_), .Y(_3366_) );
AOI21X1 AOI21X1_851 ( .A(_3359_), .B(_3366_), .C(_1888__bF_buf3), .Y(_3367_) );
MUX2X1 MUX2X1_259 ( .A(datapath_1_RegisterFile_regfile_mem_18__28_), .B(datapath_1_RegisterFile_regfile_mem_16__28_), .S(datapath_1_Instr_22_bF_buf30_), .Y(_3368_) );
NAND2X1 NAND2X1_1337 ( .A(_1890__bF_buf2), .B(_3368_), .Y(_3369_) );
MUX2X1 MUX2X1_260 ( .A(datapath_1_RegisterFile_regfile_mem_19__28_), .B(datapath_1_RegisterFile_regfile_mem_17__28_), .S(datapath_1_Instr_22_bF_buf29_), .Y(_3370_) );
NAND2X1 NAND2X1_1338 ( .A(datapath_1_Instr_21_bF_buf18_), .B(_3370_), .Y(_3371_) );
NAND3X1 NAND3X1_1538 ( .A(_1885__bF_buf7), .B(_3369_), .C(_3371_), .Y(_3372_) );
MUX2X1 MUX2X1_261 ( .A(datapath_1_RegisterFile_regfile_mem_22__28_), .B(datapath_1_RegisterFile_regfile_mem_20__28_), .S(datapath_1_Instr_22_bF_buf28_), .Y(_3373_) );
NAND2X1 NAND2X1_1339 ( .A(_1890__bF_buf2), .B(_3373_), .Y(_3374_) );
MUX2X1 MUX2X1_262 ( .A(datapath_1_RegisterFile_regfile_mem_23__28_), .B(datapath_1_RegisterFile_regfile_mem_21__28_), .S(datapath_1_Instr_22_bF_buf27_), .Y(_3375_) );
NAND2X1 NAND2X1_1340 ( .A(datapath_1_Instr_21_bF_buf17_), .B(_3375_), .Y(_3376_) );
NAND3X1 NAND3X1_1539 ( .A(datapath_1_Instr_23_bF_buf6_bF_buf1_), .B(_3374_), .C(_3376_), .Y(_3377_) );
AOI21X1 AOI21X1_852 ( .A(_3372_), .B(_3377_), .C(datapath_1_Instr_24_bF_buf5_), .Y(_3378_) );
OAI21X1 OAI21X1_1918 ( .A(_3378_), .B(_3367_), .C(datapath_1_Instr_25_bF_buf3_), .Y(_3379_) );
MUX2X1 MUX2X1_263 ( .A(datapath_1_RegisterFile_regfile_mem_9__28_), .B(datapath_1_RegisterFile_regfile_mem_8__28_), .S(datapath_1_Instr_21_bF_buf16_), .Y(_3380_) );
NOR2X1 NOR2X1_468 ( .A(datapath_1_RegisterFile_regfile_mem_11__28_), .B(_1890__bF_buf47), .Y(_3381_) );
OAI21X1 OAI21X1_1919 ( .A(datapath_1_Instr_21_bF_buf15_), .B(datapath_1_RegisterFile_regfile_mem_10__28_), .C(datapath_1_Instr_22_bF_buf26_), .Y(_3382_) );
OAI22X1 OAI22X1_247 ( .A(_3382_), .B(_3381_), .C(datapath_1_Instr_22_bF_buf25_), .D(_3380_), .Y(_3383_) );
INVX1 INVX1_476 ( .A(datapath_1_RegisterFile_regfile_mem_15__28_), .Y(_3384_) );
AOI21X1 AOI21X1_853 ( .A(_1890__bF_buf47), .B(datapath_1_RegisterFile_regfile_mem_14__28_), .C(_1884__bF_buf0), .Y(_3385_) );
OAI21X1 OAI21X1_1920 ( .A(_1890__bF_buf47), .B(_3384_), .C(_3385_), .Y(_3386_) );
NAND2X1 NAND2X1_1341 ( .A(datapath_1_RegisterFile_regfile_mem_12__28_), .B(_1890__bF_buf47), .Y(_3387_) );
AOI21X1 AOI21X1_854 ( .A(datapath_1_Instr_21_bF_buf14_), .B(datapath_1_RegisterFile_regfile_mem_13__28_), .C(datapath_1_Instr_22_bF_buf24_), .Y(_3388_) );
AOI21X1 AOI21X1_855 ( .A(_3387_), .B(_3388_), .C(_1885__bF_buf2), .Y(_3389_) );
AOI22X1 AOI22X1_182 ( .A(_3386_), .B(_3389_), .C(_1885__bF_buf2), .D(_3383_), .Y(_3390_) );
NOR2X1 NOR2X1_469 ( .A(datapath_1_Instr_21_bF_buf13_), .B(datapath_1_RegisterFile_regfile_mem_0__28_), .Y(_3391_) );
OAI21X1 OAI21X1_1921 ( .A(datapath_1_RegisterFile_regfile_mem_1__28_), .B(_1890__bF_buf47), .C(_1884__bF_buf0), .Y(_3392_) );
NOR2X1 NOR2X1_470 ( .A(datapath_1_RegisterFile_regfile_mem_3__28_), .B(_1890__bF_buf3), .Y(_3393_) );
OAI21X1 OAI21X1_1922 ( .A(datapath_1_Instr_21_bF_buf12_), .B(datapath_1_RegisterFile_regfile_mem_2__28_), .C(datapath_1_Instr_22_bF_buf23_), .Y(_3394_) );
OAI22X1 OAI22X1_248 ( .A(_3393_), .B(_3394_), .C(_3391_), .D(_3392_), .Y(_3395_) );
NOR2X1 NOR2X1_471 ( .A(datapath_1_Instr_23_bF_buf5_bF_buf1_), .B(_3395_), .Y(_3396_) );
MUX2X1 MUX2X1_264 ( .A(datapath_1_RegisterFile_regfile_mem_5__28_), .B(datapath_1_RegisterFile_regfile_mem_4__28_), .S(datapath_1_Instr_21_bF_buf11_), .Y(_3397_) );
NOR2X1 NOR2X1_472 ( .A(datapath_1_RegisterFile_regfile_mem_7__28_), .B(_1890__bF_buf42), .Y(_3398_) );
OAI21X1 OAI21X1_1923 ( .A(datapath_1_Instr_21_bF_buf10_), .B(datapath_1_RegisterFile_regfile_mem_6__28_), .C(datapath_1_Instr_22_bF_buf22_), .Y(_3399_) );
OAI22X1 OAI22X1_249 ( .A(_3399_), .B(_3398_), .C(datapath_1_Instr_22_bF_buf21_), .D(_3397_), .Y(_3400_) );
OAI21X1 OAI21X1_1924 ( .A(_1885__bF_buf2), .B(_3400_), .C(_1888__bF_buf7), .Y(_3401_) );
OAI22X1 OAI22X1_250 ( .A(_1888__bF_buf4), .B(_3390_), .C(_3396_), .D(_3401_), .Y(_3402_) );
NAND2X1 NAND2X1_1342 ( .A(_1917__bF_buf1), .B(_3402_), .Y(_3403_) );
AOI22X1 AOI22X1_183 ( .A(_1883__bF_buf3), .B(_1887__bF_buf1), .C(_3379_), .D(_3403_), .Y(datapath_1_RD1_28_) );
NAND2X1 NAND2X1_1343 ( .A(datapath_1_Instr_22_bF_buf20_), .B(datapath_1_RegisterFile_regfile_mem_11__29_), .Y(_3404_) );
NAND2X1 NAND2X1_1344 ( .A(datapath_1_RegisterFile_regfile_mem_9__29_), .B(_1884__bF_buf0), .Y(_3405_) );
NAND3X1 NAND3X1_1540 ( .A(datapath_1_Instr_21_bF_buf9_), .B(_3404_), .C(_3405_), .Y(_3406_) );
NAND2X1 NAND2X1_1345 ( .A(datapath_1_Instr_22_bF_buf19_), .B(datapath_1_RegisterFile_regfile_mem_10__29_), .Y(_3407_) );
AOI21X1 AOI21X1_856 ( .A(_1884__bF_buf0), .B(datapath_1_RegisterFile_regfile_mem_8__29_), .C(datapath_1_Instr_21_bF_buf8_), .Y(_3408_) );
NAND2X1 NAND2X1_1346 ( .A(_3407_), .B(_3408_), .Y(_3409_) );
NAND3X1 NAND3X1_1541 ( .A(_1885__bF_buf2), .B(_3406_), .C(_3409_), .Y(_3410_) );
NAND2X1 NAND2X1_1347 ( .A(datapath_1_Instr_22_bF_buf18_), .B(datapath_1_RegisterFile_regfile_mem_15__29_), .Y(_3411_) );
NAND2X1 NAND2X1_1348 ( .A(datapath_1_RegisterFile_regfile_mem_13__29_), .B(_1884__bF_buf0), .Y(_3412_) );
NAND3X1 NAND3X1_1542 ( .A(datapath_1_Instr_21_bF_buf7_), .B(_3411_), .C(_3412_), .Y(_3413_) );
NAND2X1 NAND2X1_1349 ( .A(datapath_1_Instr_22_bF_buf17_), .B(datapath_1_RegisterFile_regfile_mem_14__29_), .Y(_3414_) );
AOI21X1 AOI21X1_857 ( .A(_1884__bF_buf0), .B(datapath_1_RegisterFile_regfile_mem_12__29_), .C(datapath_1_Instr_21_bF_buf6_), .Y(_3415_) );
NAND2X1 NAND2X1_1350 ( .A(_3414_), .B(_3415_), .Y(_3416_) );
NAND3X1 NAND3X1_1543 ( .A(datapath_1_Instr_23_bF_buf4_bF_buf1_), .B(_3413_), .C(_3416_), .Y(_3417_) );
AOI21X1 AOI21X1_858 ( .A(_3410_), .B(_3417_), .C(_1888__bF_buf7), .Y(_3418_) );
INVX1 INVX1_477 ( .A(datapath_1_RegisterFile_regfile_mem_1__29_), .Y(_3419_) );
AOI21X1 AOI21X1_859 ( .A(datapath_1_Instr_23_bF_buf3_bF_buf1_), .B(datapath_1_RegisterFile_regfile_mem_5__29_), .C(_1890__bF_buf8), .Y(_3420_) );
OAI21X1 OAI21X1_1925 ( .A(datapath_1_Instr_23_bF_buf2_bF_buf1_), .B(_3419_), .C(_3420_), .Y(_3421_) );
INVX1 INVX1_478 ( .A(datapath_1_RegisterFile_regfile_mem_0__29_), .Y(_3422_) );
AOI21X1 AOI21X1_860 ( .A(datapath_1_Instr_23_bF_buf1_), .B(datapath_1_RegisterFile_regfile_mem_4__29_), .C(datapath_1_Instr_21_bF_buf5_), .Y(_3423_) );
OAI21X1 OAI21X1_1926 ( .A(datapath_1_Instr_23_bF_buf0_), .B(_3422_), .C(_3423_), .Y(_3424_) );
NAND3X1 NAND3X1_1544 ( .A(_1884__bF_buf8), .B(_3424_), .C(_3421_), .Y(_3425_) );
INVX1 INVX1_479 ( .A(datapath_1_RegisterFile_regfile_mem_3__29_), .Y(_3426_) );
AOI21X1 AOI21X1_861 ( .A(datapath_1_Instr_23_bF_buf15_bF_buf0_), .B(datapath_1_RegisterFile_regfile_mem_7__29_), .C(_1890__bF_buf8), .Y(_3427_) );
OAI21X1 OAI21X1_1927 ( .A(datapath_1_Instr_23_bF_buf14_bF_buf0_), .B(_3426_), .C(_3427_), .Y(_3428_) );
INVX1 INVX1_480 ( .A(datapath_1_RegisterFile_regfile_mem_2__29_), .Y(_3429_) );
AOI21X1 AOI21X1_862 ( .A(datapath_1_Instr_23_bF_buf13_bF_buf0_), .B(datapath_1_RegisterFile_regfile_mem_6__29_), .C(datapath_1_Instr_21_bF_buf4_), .Y(_3430_) );
OAI21X1 OAI21X1_1928 ( .A(datapath_1_Instr_23_bF_buf12_bF_buf0_), .B(_3429_), .C(_3430_), .Y(_3431_) );
NAND3X1 NAND3X1_1545 ( .A(datapath_1_Instr_22_bF_buf16_), .B(_3431_), .C(_3428_), .Y(_3432_) );
AOI21X1 AOI21X1_863 ( .A(_3425_), .B(_3432_), .C(datapath_1_Instr_24_bF_buf4_), .Y(_3433_) );
OAI21X1 OAI21X1_1929 ( .A(_3433_), .B(_3418_), .C(_1917__bF_buf2), .Y(_3434_) );
INVX1 INVX1_481 ( .A(datapath_1_RegisterFile_regfile_mem_19__29_), .Y(_3435_) );
AOI21X1 AOI21X1_864 ( .A(datapath_1_Instr_23_bF_buf11_bF_buf0_), .B(datapath_1_RegisterFile_regfile_mem_23__29_), .C(_1890__bF_buf43), .Y(_3436_) );
OAI21X1 OAI21X1_1930 ( .A(datapath_1_Instr_23_bF_buf10_bF_buf0_), .B(_3435_), .C(_3436_), .Y(_3437_) );
NAND2X1 NAND2X1_1351 ( .A(datapath_1_RegisterFile_regfile_mem_18__29_), .B(_1885__bF_buf3), .Y(_3438_) );
AOI21X1 AOI21X1_865 ( .A(datapath_1_Instr_23_bF_buf9_bF_buf0_), .B(datapath_1_RegisterFile_regfile_mem_22__29_), .C(datapath_1_Instr_21_bF_buf3_), .Y(_3439_) );
AOI21X1 AOI21X1_866 ( .A(_3438_), .B(_3439_), .C(_1884__bF_buf2), .Y(_3440_) );
INVX1 INVX1_482 ( .A(datapath_1_RegisterFile_regfile_mem_17__29_), .Y(_3441_) );
AOI21X1 AOI21X1_867 ( .A(datapath_1_Instr_23_bF_buf8_bF_buf0_), .B(datapath_1_RegisterFile_regfile_mem_21__29_), .C(_1890__bF_buf43), .Y(_3442_) );
OAI21X1 OAI21X1_1931 ( .A(datapath_1_Instr_23_bF_buf7_bF_buf0_), .B(_3441_), .C(_3442_), .Y(_3443_) );
NAND2X1 NAND2X1_1352 ( .A(datapath_1_RegisterFile_regfile_mem_16__29_), .B(_1885__bF_buf3), .Y(_3444_) );
AOI21X1 AOI21X1_868 ( .A(datapath_1_Instr_23_bF_buf6_bF_buf0_), .B(datapath_1_RegisterFile_regfile_mem_20__29_), .C(datapath_1_Instr_21_bF_buf2_), .Y(_3445_) );
AOI21X1 AOI21X1_869 ( .A(_3444_), .B(_3445_), .C(datapath_1_Instr_22_bF_buf15_), .Y(_3446_) );
AOI22X1 AOI22X1_184 ( .A(_3440_), .B(_3437_), .C(_3443_), .D(_3446_), .Y(_3447_) );
NOR2X1 NOR2X1_473 ( .A(datapath_1_Instr_21_bF_buf1_), .B(datapath_1_RegisterFile_regfile_mem_24__29_), .Y(_3448_) );
OAI21X1 OAI21X1_1932 ( .A(datapath_1_RegisterFile_regfile_mem_25__29_), .B(_1890__bF_buf35), .C(_1884__bF_buf6), .Y(_3449_) );
NOR2X1 NOR2X1_474 ( .A(datapath_1_RegisterFile_regfile_mem_27__29_), .B(_1890__bF_buf6), .Y(_3450_) );
OAI21X1 OAI21X1_1933 ( .A(datapath_1_Instr_21_bF_buf0_), .B(datapath_1_RegisterFile_regfile_mem_26__29_), .C(datapath_1_Instr_22_bF_buf14_), .Y(_3451_) );
OAI22X1 OAI22X1_251 ( .A(_3450_), .B(_3451_), .C(_3448_), .D(_3449_), .Y(_3452_) );
NOR2X1 NOR2X1_475 ( .A(datapath_1_Instr_23_bF_buf5_bF_buf0_), .B(_3452_), .Y(_3453_) );
MUX2X1 MUX2X1_265 ( .A(datapath_1_RegisterFile_regfile_mem_29__29_), .B(datapath_1_RegisterFile_regfile_mem_28__29_), .S(datapath_1_Instr_21_bF_buf55_), .Y(_3454_) );
NOR2X1 NOR2X1_476 ( .A(datapath_1_RegisterFile_regfile_mem_31__29_), .B(_1890__bF_buf11), .Y(_3455_) );
OAI21X1 OAI21X1_1934 ( .A(datapath_1_Instr_21_bF_buf54_), .B(datapath_1_RegisterFile_regfile_mem_30__29_), .C(datapath_1_Instr_22_bF_buf13_), .Y(_3456_) );
OAI22X1 OAI22X1_252 ( .A(_3456_), .B(_3455_), .C(datapath_1_Instr_22_bF_buf12_), .D(_3454_), .Y(_3457_) );
OAI21X1 OAI21X1_1935 ( .A(_1885__bF_buf3), .B(_3457_), .C(datapath_1_Instr_24_bF_buf3_), .Y(_3458_) );
OAI22X1 OAI22X1_253 ( .A(datapath_1_Instr_24_bF_buf2_), .B(_3447_), .C(_3453_), .D(_3458_), .Y(_3459_) );
NAND2X1 NAND2X1_1353 ( .A(datapath_1_Instr_25_bF_buf2_), .B(_3459_), .Y(_3460_) );
AOI22X1 AOI22X1_185 ( .A(_1883__bF_buf1), .B(_1887__bF_buf0), .C(_3434_), .D(_3460_), .Y(datapath_1_RD1_29_) );
MUX2X1 MUX2X1_266 ( .A(datapath_1_RegisterFile_regfile_mem_9__30_), .B(datapath_1_RegisterFile_regfile_mem_8__30_), .S(datapath_1_Instr_21_bF_buf53_), .Y(_3461_) );
NOR2X1 NOR2X1_477 ( .A(datapath_1_RegisterFile_regfile_mem_11__30_), .B(_1890__bF_buf20), .Y(_3462_) );
OAI21X1 OAI21X1_1936 ( .A(datapath_1_Instr_21_bF_buf52_), .B(datapath_1_RegisterFile_regfile_mem_10__30_), .C(datapath_1_Instr_22_bF_buf11_), .Y(_3463_) );
OAI22X1 OAI22X1_254 ( .A(_3463_), .B(_3462_), .C(datapath_1_Instr_22_bF_buf10_), .D(_3461_), .Y(_3464_) );
INVX1 INVX1_483 ( .A(datapath_1_RegisterFile_regfile_mem_15__30_), .Y(_3465_) );
AOI21X1 AOI21X1_870 ( .A(_1890__bF_buf28), .B(datapath_1_RegisterFile_regfile_mem_14__30_), .C(_1884__bF_buf1), .Y(_3466_) );
OAI21X1 OAI21X1_1937 ( .A(_1890__bF_buf28), .B(_3465_), .C(_3466_), .Y(_3467_) );
NAND2X1 NAND2X1_1354 ( .A(datapath_1_RegisterFile_regfile_mem_12__30_), .B(_1890__bF_buf20), .Y(_3468_) );
AOI21X1 AOI21X1_871 ( .A(datapath_1_Instr_21_bF_buf51_), .B(datapath_1_RegisterFile_regfile_mem_13__30_), .C(datapath_1_Instr_22_bF_buf9_), .Y(_3469_) );
AOI21X1 AOI21X1_872 ( .A(_3468_), .B(_3469_), .C(_1885__bF_buf5), .Y(_3470_) );
AOI22X1 AOI22X1_186 ( .A(_3467_), .B(_3470_), .C(_1885__bF_buf5), .D(_3464_), .Y(_3471_) );
NOR2X1 NOR2X1_478 ( .A(datapath_1_Instr_21_bF_buf50_), .B(datapath_1_RegisterFile_regfile_mem_0__30_), .Y(_3472_) );
OAI21X1 OAI21X1_1938 ( .A(datapath_1_RegisterFile_regfile_mem_1__30_), .B(_1890__bF_buf1), .C(_1884__bF_buf4), .Y(_3473_) );
NOR2X1 NOR2X1_479 ( .A(datapath_1_RegisterFile_regfile_mem_3__30_), .B(_1890__bF_buf27), .Y(_3474_) );
OAI21X1 OAI21X1_1939 ( .A(datapath_1_Instr_21_bF_buf49_), .B(datapath_1_RegisterFile_regfile_mem_2__30_), .C(datapath_1_Instr_22_bF_buf8_), .Y(_3475_) );
OAI22X1 OAI22X1_255 ( .A(_3474_), .B(_3475_), .C(_3472_), .D(_3473_), .Y(_3476_) );
NOR2X1 NOR2X1_480 ( .A(datapath_1_Instr_23_bF_buf4_bF_buf0_), .B(_3476_), .Y(_3477_) );
MUX2X1 MUX2X1_267 ( .A(datapath_1_RegisterFile_regfile_mem_5__30_), .B(datapath_1_RegisterFile_regfile_mem_4__30_), .S(datapath_1_Instr_21_bF_buf48_), .Y(_3478_) );
NOR2X1 NOR2X1_481 ( .A(datapath_1_RegisterFile_regfile_mem_7__30_), .B(_1890__bF_buf27), .Y(_3479_) );
OAI21X1 OAI21X1_1940 ( .A(datapath_1_Instr_21_bF_buf47_), .B(datapath_1_RegisterFile_regfile_mem_6__30_), .C(datapath_1_Instr_22_bF_buf7_), .Y(_3480_) );
OAI22X1 OAI22X1_256 ( .A(_3480_), .B(_3479_), .C(datapath_1_Instr_22_bF_buf6_), .D(_3478_), .Y(_3481_) );
OAI21X1 OAI21X1_1941 ( .A(_1885__bF_buf4), .B(_3481_), .C(_1888__bF_buf0), .Y(_3482_) );
OAI22X1 OAI22X1_257 ( .A(_1888__bF_buf0), .B(_3471_), .C(_3477_), .D(_3482_), .Y(_3483_) );
NAND2X1 NAND2X1_1355 ( .A(_1917__bF_buf0), .B(_3483_), .Y(_3484_) );
INVX1 INVX1_484 ( .A(datapath_1_RegisterFile_regfile_mem_19__30_), .Y(_3485_) );
AOI21X1 AOI21X1_873 ( .A(datapath_1_Instr_23_bF_buf3_bF_buf0_), .B(datapath_1_RegisterFile_regfile_mem_23__30_), .C(_1890__bF_buf40), .Y(_3486_) );
OAI21X1 OAI21X1_1942 ( .A(datapath_1_Instr_23_bF_buf2_bF_buf0_), .B(_3485_), .C(_3486_), .Y(_3487_) );
NAND2X1 NAND2X1_1356 ( .A(datapath_1_RegisterFile_regfile_mem_18__30_), .B(_1885__bF_buf9), .Y(_3488_) );
AOI21X1 AOI21X1_874 ( .A(datapath_1_Instr_23_bF_buf1_), .B(datapath_1_RegisterFile_regfile_mem_22__30_), .C(datapath_1_Instr_21_bF_buf46_), .Y(_3489_) );
AOI21X1 AOI21X1_875 ( .A(_3488_), .B(_3489_), .C(_1884__bF_buf9), .Y(_3490_) );
INVX1 INVX1_485 ( .A(datapath_1_RegisterFile_regfile_mem_17__30_), .Y(_3491_) );
AOI21X1 AOI21X1_876 ( .A(datapath_1_Instr_23_bF_buf0_), .B(datapath_1_RegisterFile_regfile_mem_21__30_), .C(_1890__bF_buf9), .Y(_3492_) );
OAI21X1 OAI21X1_1943 ( .A(datapath_1_Instr_23_bF_buf15_bF_buf3_), .B(_3491_), .C(_3492_), .Y(_3493_) );
NAND2X1 NAND2X1_1357 ( .A(datapath_1_RegisterFile_regfile_mem_16__30_), .B(_1885__bF_buf11), .Y(_3494_) );
AOI21X1 AOI21X1_877 ( .A(datapath_1_Instr_23_bF_buf14_bF_buf3_), .B(datapath_1_RegisterFile_regfile_mem_20__30_), .C(datapath_1_Instr_21_bF_buf45_), .Y(_3495_) );
AOI21X1 AOI21X1_878 ( .A(_3494_), .B(_3495_), .C(datapath_1_Instr_22_bF_buf5_), .Y(_3496_) );
AOI22X1 AOI22X1_187 ( .A(_3490_), .B(_3487_), .C(_3493_), .D(_3496_), .Y(_3497_) );
NOR2X1 NOR2X1_482 ( .A(datapath_1_Instr_21_bF_buf44_), .B(datapath_1_RegisterFile_regfile_mem_24__30_), .Y(_3498_) );
OAI21X1 OAI21X1_1944 ( .A(datapath_1_RegisterFile_regfile_mem_25__30_), .B(_1890__bF_buf7), .C(_1884__bF_buf9), .Y(_3499_) );
NOR2X1 NOR2X1_483 ( .A(datapath_1_RegisterFile_regfile_mem_27__30_), .B(_1890__bF_buf7), .Y(_3500_) );
OAI21X1 OAI21X1_1945 ( .A(datapath_1_Instr_21_bF_buf43_), .B(datapath_1_RegisterFile_regfile_mem_26__30_), .C(datapath_1_Instr_22_bF_buf4_), .Y(_3501_) );
OAI22X1 OAI22X1_258 ( .A(_3500_), .B(_3501_), .C(_3498_), .D(_3499_), .Y(_3502_) );
NOR2X1 NOR2X1_484 ( .A(datapath_1_Instr_23_bF_buf13_bF_buf3_), .B(_3502_), .Y(_3503_) );
MUX2X1 MUX2X1_268 ( .A(datapath_1_RegisterFile_regfile_mem_29__30_), .B(datapath_1_RegisterFile_regfile_mem_28__30_), .S(datapath_1_Instr_21_bF_buf42_), .Y(_3504_) );
NOR2X1 NOR2X1_485 ( .A(datapath_1_RegisterFile_regfile_mem_31__30_), .B(_1890__bF_buf40), .Y(_3505_) );
OAI21X1 OAI21X1_1946 ( .A(datapath_1_Instr_21_bF_buf41_), .B(datapath_1_RegisterFile_regfile_mem_30__30_), .C(datapath_1_Instr_22_bF_buf3_), .Y(_3506_) );
OAI22X1 OAI22X1_259 ( .A(_3506_), .B(_3505_), .C(datapath_1_Instr_22_bF_buf2_), .D(_3504_), .Y(_3507_) );
OAI21X1 OAI21X1_1947 ( .A(_1885__bF_buf9), .B(_3507_), .C(datapath_1_Instr_24_bF_buf1_), .Y(_3508_) );
OAI22X1 OAI22X1_260 ( .A(datapath_1_Instr_24_bF_buf0_), .B(_3497_), .C(_3503_), .D(_3508_), .Y(_3509_) );
NAND2X1 NAND2X1_1358 ( .A(datapath_1_Instr_25_bF_buf1_), .B(_3509_), .Y(_3510_) );
AOI22X1 AOI22X1_188 ( .A(_1883__bF_buf2), .B(_1887__bF_buf4), .C(_3510_), .D(_3484_), .Y(datapath_1_RD1_30_) );
NAND2X1 NAND2X1_1359 ( .A(datapath_1_Instr_21_bF_buf40_), .B(datapath_1_RegisterFile_regfile_mem_27__31_), .Y(_3511_) );
NAND2X1 NAND2X1_1360 ( .A(datapath_1_RegisterFile_regfile_mem_26__31_), .B(_1890__bF_buf34), .Y(_3512_) );
NAND3X1 NAND3X1_1546 ( .A(datapath_1_Instr_22_bF_buf1_), .B(_3511_), .C(_3512_), .Y(_3513_) );
NAND2X1 NAND2X1_1361 ( .A(datapath_1_Instr_21_bF_buf39_), .B(datapath_1_RegisterFile_regfile_mem_25__31_), .Y(_3514_) );
AOI21X1 AOI21X1_879 ( .A(_1890__bF_buf4), .B(datapath_1_RegisterFile_regfile_mem_24__31_), .C(datapath_1_Instr_22_bF_buf0_), .Y(_3515_) );
NAND2X1 NAND2X1_1362 ( .A(_3514_), .B(_3515_), .Y(_3516_) );
NAND3X1 NAND3X1_1547 ( .A(_1885__bF_buf6), .B(_3513_), .C(_3516_), .Y(_3517_) );
NAND2X1 NAND2X1_1363 ( .A(datapath_1_Instr_21_bF_buf38_), .B(datapath_1_RegisterFile_regfile_mem_31__31_), .Y(_3518_) );
AOI21X1 AOI21X1_880 ( .A(_1890__bF_buf34), .B(datapath_1_RegisterFile_regfile_mem_30__31_), .C(_1884__bF_buf3), .Y(_3519_) );
NAND2X1 NAND2X1_1364 ( .A(_3518_), .B(_3519_), .Y(_3520_) );
INVX1 INVX1_486 ( .A(datapath_1_RegisterFile_regfile_mem_28__31_), .Y(_3521_) );
AOI21X1 AOI21X1_881 ( .A(datapath_1_Instr_21_bF_buf37_), .B(datapath_1_RegisterFile_regfile_mem_29__31_), .C(datapath_1_Instr_22_bF_buf50_), .Y(_3522_) );
OAI21X1 OAI21X1_1948 ( .A(datapath_1_Instr_21_bF_buf36_), .B(_3521_), .C(_3522_), .Y(_3523_) );
NAND3X1 NAND3X1_1548 ( .A(datapath_1_Instr_23_bF_buf12_bF_buf3_), .B(_3523_), .C(_3520_), .Y(_3524_) );
AOI21X1 AOI21X1_882 ( .A(_3517_), .B(_3524_), .C(_1888__bF_buf1), .Y(_3525_) );
MUX2X1 MUX2X1_269 ( .A(datapath_1_RegisterFile_regfile_mem_18__31_), .B(datapath_1_RegisterFile_regfile_mem_16__31_), .S(datapath_1_Instr_22_bF_buf49_), .Y(_3526_) );
NAND2X1 NAND2X1_1365 ( .A(_1890__bF_buf39), .B(_3526_), .Y(_3527_) );
MUX2X1 MUX2X1_270 ( .A(datapath_1_RegisterFile_regfile_mem_19__31_), .B(datapath_1_RegisterFile_regfile_mem_17__31_), .S(datapath_1_Instr_22_bF_buf48_), .Y(_3528_) );
NAND2X1 NAND2X1_1366 ( .A(datapath_1_Instr_21_bF_buf35_), .B(_3528_), .Y(_3529_) );
NAND3X1 NAND3X1_1549 ( .A(_1885__bF_buf6), .B(_3527_), .C(_3529_), .Y(_3530_) );
MUX2X1 MUX2X1_271 ( .A(datapath_1_RegisterFile_regfile_mem_22__31_), .B(datapath_1_RegisterFile_regfile_mem_20__31_), .S(datapath_1_Instr_22_bF_buf47_), .Y(_3531_) );
NAND2X1 NAND2X1_1367 ( .A(_1890__bF_buf39), .B(_3531_), .Y(_3532_) );
MUX2X1 MUX2X1_272 ( .A(datapath_1_RegisterFile_regfile_mem_23__31_), .B(datapath_1_RegisterFile_regfile_mem_21__31_), .S(datapath_1_Instr_22_bF_buf46_), .Y(_3533_) );
NAND2X1 NAND2X1_1368 ( .A(datapath_1_Instr_21_bF_buf34_), .B(_3533_), .Y(_3534_) );
NAND3X1 NAND3X1_1550 ( .A(datapath_1_Instr_23_bF_buf11_bF_buf3_), .B(_3532_), .C(_3534_), .Y(_3535_) );
AOI21X1 AOI21X1_883 ( .A(_3530_), .B(_3535_), .C(datapath_1_Instr_24_bF_buf6_), .Y(_3536_) );
OAI21X1 OAI21X1_1949 ( .A(_3536_), .B(_3525_), .C(datapath_1_Instr_25_bF_buf0_), .Y(_3537_) );
INVX1 INVX1_487 ( .A(datapath_1_RegisterFile_regfile_mem_9__31_), .Y(_3538_) );
AOI21X1 AOI21X1_884 ( .A(datapath_1_Instr_23_bF_buf10_bF_buf3_), .B(datapath_1_RegisterFile_regfile_mem_13__31_), .C(_1890__bF_buf5), .Y(_3539_) );
OAI21X1 OAI21X1_1950 ( .A(datapath_1_Instr_23_bF_buf9_bF_buf3_), .B(_3538_), .C(_3539_), .Y(_3540_) );
INVX1 INVX1_488 ( .A(datapath_1_RegisterFile_regfile_mem_8__31_), .Y(_3541_) );
AOI21X1 AOI21X1_885 ( .A(datapath_1_Instr_23_bF_buf8_bF_buf3_), .B(datapath_1_RegisterFile_regfile_mem_12__31_), .C(datapath_1_Instr_21_bF_buf33_), .Y(_3542_) );
OAI21X1 OAI21X1_1951 ( .A(datapath_1_Instr_23_bF_buf7_bF_buf3_), .B(_3541_), .C(_3542_), .Y(_3543_) );
NAND3X1 NAND3X1_1551 ( .A(_1884__bF_buf5), .B(_3543_), .C(_3540_), .Y(_3544_) );
INVX1 INVX1_489 ( .A(datapath_1_RegisterFile_regfile_mem_11__31_), .Y(_3545_) );
AOI21X1 AOI21X1_886 ( .A(datapath_1_Instr_23_bF_buf6_bF_buf3_), .B(datapath_1_RegisterFile_regfile_mem_15__31_), .C(_1890__bF_buf20), .Y(_3546_) );
OAI21X1 OAI21X1_1952 ( .A(datapath_1_Instr_23_bF_buf5_bF_buf3_), .B(_3545_), .C(_3546_), .Y(_3547_) );
INVX1 INVX1_490 ( .A(datapath_1_RegisterFile_regfile_mem_10__31_), .Y(_3548_) );
AOI21X1 AOI21X1_887 ( .A(datapath_1_Instr_23_bF_buf4_bF_buf3_), .B(datapath_1_RegisterFile_regfile_mem_14__31_), .C(datapath_1_Instr_21_bF_buf32_), .Y(_3549_) );
OAI21X1 OAI21X1_1953 ( .A(datapath_1_Instr_23_bF_buf3_bF_buf3_), .B(_3548_), .C(_3549_), .Y(_3550_) );
NAND3X1 NAND3X1_1552 ( .A(datapath_1_Instr_22_bF_buf45_), .B(_3550_), .C(_3547_), .Y(_3551_) );
AOI21X1 AOI21X1_888 ( .A(_3544_), .B(_3551_), .C(_1888__bF_buf5), .Y(_3552_) );
MUX2X1 MUX2X1_273 ( .A(datapath_1_RegisterFile_regfile_mem_1__31_), .B(datapath_1_RegisterFile_regfile_mem_0__31_), .S(datapath_1_Instr_21_bF_buf31_), .Y(_3553_) );
NOR2X1 NOR2X1_486 ( .A(datapath_1_RegisterFile_regfile_mem_3__31_), .B(_1890__bF_buf33), .Y(_3554_) );
OAI21X1 OAI21X1_1954 ( .A(datapath_1_Instr_21_bF_buf30_), .B(datapath_1_RegisterFile_regfile_mem_2__31_), .C(datapath_1_Instr_22_bF_buf44_), .Y(_3555_) );
OAI22X1 OAI22X1_261 ( .A(_3555_), .B(_3554_), .C(datapath_1_Instr_22_bF_buf43_), .D(_3553_), .Y(_3556_) );
NAND2X1 NAND2X1_1369 ( .A(_1885__bF_buf4), .B(_3556_), .Y(_3557_) );
MUX2X1 MUX2X1_274 ( .A(datapath_1_RegisterFile_regfile_mem_5__31_), .B(datapath_1_RegisterFile_regfile_mem_4__31_), .S(datapath_1_Instr_21_bF_buf29_), .Y(_3558_) );
NOR2X1 NOR2X1_487 ( .A(datapath_1_RegisterFile_regfile_mem_7__31_), .B(_1890__bF_buf46), .Y(_3559_) );
OAI21X1 OAI21X1_1955 ( .A(datapath_1_Instr_21_bF_buf28_), .B(datapath_1_RegisterFile_regfile_mem_6__31_), .C(datapath_1_Instr_22_bF_buf42_), .Y(_3560_) );
OAI22X1 OAI22X1_262 ( .A(_3560_), .B(_3559_), .C(datapath_1_Instr_22_bF_buf41_), .D(_3558_), .Y(_3561_) );
NAND2X1 NAND2X1_1370 ( .A(datapath_1_Instr_23_bF_buf2_bF_buf3_), .B(_3561_), .Y(_3562_) );
AOI21X1 AOI21X1_889 ( .A(_3557_), .B(_3562_), .C(datapath_1_Instr_24_bF_buf5_), .Y(_3563_) );
OAI21X1 OAI21X1_1956 ( .A(_3552_), .B(_3563_), .C(_1917__bF_buf4), .Y(_3564_) );
AOI22X1 AOI22X1_189 ( .A(_1883__bF_buf4), .B(_1887__bF_buf3), .C(_3537_), .D(_3564_), .Y(datapath_1_RD1_31_) );
NOR2X1 NOR2X1_488 ( .A(datapath_1_Instr_20_bF_buf2_), .B(datapath_1_Instr_16_bF_buf47_), .Y(_3565_) );
INVX1 INVX1_491 ( .A(datapath_1_Instr_17_bF_buf7_), .Y(_3566_) );
INVX1 INVX1_492 ( .A(datapath_1_Instr_18_bF_buf0_), .Y(_3567_) );
NAND2X1 NAND2X1_1371 ( .A(_3566__bF_buf10), .B(_3567__bF_buf2), .Y(_3568_) );
NOR2X1 NOR2X1_489 ( .A(datapath_1_Instr_19_bF_buf3_), .B(_3568_), .Y(_3569_) );
INVX1 INVX1_493 ( .A(datapath_1_Instr_20_bF_buf1_), .Y(_3570_) );
INVX1 INVX1_494 ( .A(datapath_1_Instr_19_bF_buf2_), .Y(_3571_) );
NAND2X1 NAND2X1_1372 ( .A(datapath_1_RegisterFile_regfile_mem_11__0_), .B(datapath_1_Instr_17_bF_buf6_), .Y(_3572_) );
NAND2X1 NAND2X1_1373 ( .A(datapath_1_RegisterFile_regfile_mem_9__0_), .B(_3566__bF_buf5), .Y(_3573_) );
NAND3X1 NAND3X1_1553 ( .A(datapath_1_Instr_16_bF_buf46_), .B(_3572_), .C(_3573_), .Y(_3574_) );
NAND2X1 NAND2X1_1374 ( .A(datapath_1_RegisterFile_regfile_mem_10__0_), .B(datapath_1_Instr_17_bF_buf5_), .Y(_3575_) );
AOI21X1 AOI21X1_890 ( .A(_3566__bF_buf5), .B(datapath_1_RegisterFile_regfile_mem_8__0_), .C(datapath_1_Instr_16_bF_buf45_), .Y(_3576_) );
NAND2X1 NAND2X1_1375 ( .A(_3575_), .B(_3576_), .Y(_3577_) );
NAND3X1 NAND3X1_1554 ( .A(_3567__bF_buf8), .B(_3574_), .C(_3577_), .Y(_3578_) );
NAND2X1 NAND2X1_1376 ( .A(datapath_1_RegisterFile_regfile_mem_15__0_), .B(datapath_1_Instr_17_bF_buf4_), .Y(_3579_) );
NAND2X1 NAND2X1_1377 ( .A(datapath_1_RegisterFile_regfile_mem_13__0_), .B(_3566__bF_buf8), .Y(_3580_) );
NAND3X1 NAND3X1_1555 ( .A(datapath_1_Instr_16_bF_buf44_), .B(_3579_), .C(_3580_), .Y(_3581_) );
NAND2X1 NAND2X1_1378 ( .A(datapath_1_RegisterFile_regfile_mem_14__0_), .B(datapath_1_Instr_17_bF_buf3_), .Y(_3582_) );
AOI21X1 AOI21X1_891 ( .A(_3566__bF_buf8), .B(datapath_1_RegisterFile_regfile_mem_12__0_), .C(datapath_1_Instr_16_bF_buf43_), .Y(_3583_) );
NAND2X1 NAND2X1_1379 ( .A(_3582_), .B(_3583_), .Y(_3584_) );
NAND3X1 NAND3X1_1556 ( .A(datapath_1_Instr_18_bF_buf44_), .B(_3581_), .C(_3584_), .Y(_3585_) );
AOI21X1 AOI21X1_892 ( .A(_3578_), .B(_3585_), .C(_3571__bF_buf3), .Y(_3586_) );
INVX1 INVX1_495 ( .A(datapath_1_RegisterFile_regfile_mem_1__0_), .Y(_3587_) );
INVX1 INVX1_496 ( .A(datapath_1_Instr_16_bF_buf42_), .Y(_3588_) );
AOI21X1 AOI21X1_893 ( .A(datapath_1_RegisterFile_regfile_mem_5__0_), .B(datapath_1_Instr_18_bF_buf43_), .C(_3588__bF_buf21), .Y(_3589_) );
OAI21X1 OAI21X1_1957 ( .A(_3587_), .B(datapath_1_Instr_18_bF_buf42_), .C(_3589_), .Y(_3590_) );
INVX1 INVX1_497 ( .A(datapath_1_RegisterFile_regfile_mem_0__0_), .Y(_3591_) );
AOI21X1 AOI21X1_894 ( .A(datapath_1_RegisterFile_regfile_mem_4__0_), .B(datapath_1_Instr_18_bF_buf41_), .C(datapath_1_Instr_16_bF_buf41_), .Y(_3592_) );
OAI21X1 OAI21X1_1958 ( .A(_3591_), .B(datapath_1_Instr_18_bF_buf40_), .C(_3592_), .Y(_3593_) );
NAND3X1 NAND3X1_1557 ( .A(_3566__bF_buf4), .B(_3593_), .C(_3590_), .Y(_3594_) );
INVX1 INVX1_498 ( .A(datapath_1_RegisterFile_regfile_mem_3__0_), .Y(_3595_) );
AOI21X1 AOI21X1_895 ( .A(datapath_1_RegisterFile_regfile_mem_7__0_), .B(datapath_1_Instr_18_bF_buf39_), .C(_3588__bF_buf21), .Y(_3596_) );
OAI21X1 OAI21X1_1959 ( .A(_3595_), .B(datapath_1_Instr_18_bF_buf38_), .C(_3596_), .Y(_3597_) );
INVX1 INVX1_499 ( .A(datapath_1_RegisterFile_regfile_mem_2__0_), .Y(_3598_) );
AOI21X1 AOI21X1_896 ( .A(datapath_1_RegisterFile_regfile_mem_6__0_), .B(datapath_1_Instr_18_bF_buf37_), .C(datapath_1_Instr_16_bF_buf40_), .Y(_3599_) );
OAI21X1 OAI21X1_1960 ( .A(_3598_), .B(datapath_1_Instr_18_bF_buf36_), .C(_3599_), .Y(_3600_) );
NAND3X1 NAND3X1_1558 ( .A(datapath_1_Instr_17_bF_buf2_), .B(_3600_), .C(_3597_), .Y(_3601_) );
AOI21X1 AOI21X1_897 ( .A(_3594_), .B(_3601_), .C(datapath_1_Instr_19_bF_buf1_), .Y(_3602_) );
OAI21X1 OAI21X1_1961 ( .A(_3602_), .B(_3586_), .C(_3570__bF_buf4), .Y(_3603_) );
INVX1 INVX1_500 ( .A(datapath_1_RegisterFile_regfile_mem_19__0_), .Y(_3604_) );
AOI21X1 AOI21X1_898 ( .A(datapath_1_RegisterFile_regfile_mem_23__0_), .B(datapath_1_Instr_18_bF_buf35_), .C(_3588__bF_buf29), .Y(_3605_) );
OAI21X1 OAI21X1_1962 ( .A(_3604_), .B(datapath_1_Instr_18_bF_buf34_), .C(_3605_), .Y(_3606_) );
NAND2X1 NAND2X1_1380 ( .A(datapath_1_RegisterFile_regfile_mem_18__0_), .B(_3567__bF_buf3), .Y(_3607_) );
AOI21X1 AOI21X1_899 ( .A(datapath_1_RegisterFile_regfile_mem_22__0_), .B(datapath_1_Instr_18_bF_buf33_), .C(datapath_1_Instr_16_bF_buf39_), .Y(_3608_) );
AOI21X1 AOI21X1_900 ( .A(_3607_), .B(_3608_), .C(_3566__bF_buf4), .Y(_3609_) );
INVX1 INVX1_501 ( .A(datapath_1_RegisterFile_regfile_mem_17__0_), .Y(_3610_) );
AOI21X1 AOI21X1_901 ( .A(datapath_1_RegisterFile_regfile_mem_21__0_), .B(datapath_1_Instr_18_bF_buf32_), .C(_3588__bF_buf29), .Y(_3611_) );
OAI21X1 OAI21X1_1963 ( .A(_3610_), .B(datapath_1_Instr_18_bF_buf31_), .C(_3611_), .Y(_3612_) );
NAND2X1 NAND2X1_1381 ( .A(datapath_1_RegisterFile_regfile_mem_16__0_), .B(_3567__bF_buf3), .Y(_3613_) );
AOI21X1 AOI21X1_902 ( .A(datapath_1_RegisterFile_regfile_mem_20__0_), .B(datapath_1_Instr_18_bF_buf30_), .C(datapath_1_Instr_16_bF_buf38_), .Y(_3614_) );
AOI21X1 AOI21X1_903 ( .A(_3613_), .B(_3614_), .C(datapath_1_Instr_17_bF_buf1_), .Y(_3615_) );
AOI22X1 AOI22X1_190 ( .A(_3609_), .B(_3606_), .C(_3612_), .D(_3615_), .Y(_3616_) );
NOR2X1 NOR2X1_490 ( .A(datapath_1_RegisterFile_regfile_mem_24__0_), .B(datapath_1_Instr_16_bF_buf37_), .Y(_3617_) );
OAI21X1 OAI21X1_1964 ( .A(datapath_1_RegisterFile_regfile_mem_25__0_), .B(_3588__bF_buf37), .C(_3566__bF_buf4), .Y(_3618_) );
NOR2X1 NOR2X1_491 ( .A(datapath_1_RegisterFile_regfile_mem_27__0_), .B(_3588__bF_buf37), .Y(_3619_) );
OAI21X1 OAI21X1_1965 ( .A(datapath_1_RegisterFile_regfile_mem_26__0_), .B(datapath_1_Instr_16_bF_buf36_), .C(datapath_1_Instr_17_bF_buf0_), .Y(_3620_) );
OAI22X1 OAI22X1_263 ( .A(_3619_), .B(_3620_), .C(_3617_), .D(_3618_), .Y(_3621_) );
NOR2X1 NOR2X1_492 ( .A(datapath_1_Instr_18_bF_buf29_), .B(_3621_), .Y(_3622_) );
MUX2X1 MUX2X1_275 ( .A(datapath_1_RegisterFile_regfile_mem_29__0_), .B(datapath_1_RegisterFile_regfile_mem_28__0_), .S(datapath_1_Instr_16_bF_buf35_), .Y(_3623_) );
NOR2X1 NOR2X1_493 ( .A(datapath_1_RegisterFile_regfile_mem_31__0_), .B(_3588__bF_buf37), .Y(_3624_) );
OAI21X1 OAI21X1_1966 ( .A(datapath_1_RegisterFile_regfile_mem_30__0_), .B(datapath_1_Instr_16_bF_buf34_), .C(datapath_1_Instr_17_bF_buf50_), .Y(_3625_) );
OAI22X1 OAI22X1_264 ( .A(_3625_), .B(_3624_), .C(datapath_1_Instr_17_bF_buf49_), .D(_3623_), .Y(_3626_) );
OAI21X1 OAI21X1_1967 ( .A(_3567__bF_buf3), .B(_3626_), .C(datapath_1_Instr_19_bF_buf0_), .Y(_3627_) );
OAI22X1 OAI22X1_265 ( .A(datapath_1_Instr_19_bF_buf6_), .B(_3616_), .C(_3622_), .D(_3627_), .Y(_3628_) );
NAND2X1 NAND2X1_1382 ( .A(datapath_1_Instr_20_bF_buf0_), .B(_3628_), .Y(_3629_) );
AOI22X1 AOI22X1_191 ( .A(_3565__bF_buf2), .B(_3569__bF_buf2), .C(_3603_), .D(_3629_), .Y(datapath_1_RD2_0_) );
INVX1 INVX1_502 ( .A(datapath_1_RegisterFile_regfile_mem_1__1_), .Y(_3630_) );
AOI21X1 AOI21X1_904 ( .A(datapath_1_RegisterFile_regfile_mem_5__1_), .B(datapath_1_Instr_18_bF_buf28_), .C(_3588__bF_buf9), .Y(_3631_) );
OAI21X1 OAI21X1_1968 ( .A(_3630_), .B(datapath_1_Instr_18_bF_buf27_), .C(_3631_), .Y(_3632_) );
INVX1 INVX1_503 ( .A(datapath_1_RegisterFile_regfile_mem_0__1_), .Y(_3633_) );
AOI21X1 AOI21X1_905 ( .A(datapath_1_RegisterFile_regfile_mem_4__1_), .B(datapath_1_Instr_18_bF_buf26_), .C(datapath_1_Instr_16_bF_buf33_), .Y(_3634_) );
OAI21X1 OAI21X1_1969 ( .A(_3633_), .B(datapath_1_Instr_18_bF_buf25_), .C(_3634_), .Y(_3635_) );
NAND3X1 NAND3X1_1559 ( .A(_3566__bF_buf7), .B(_3635_), .C(_3632_), .Y(_3636_) );
INVX1 INVX1_504 ( .A(datapath_1_RegisterFile_regfile_mem_3__1_), .Y(_3637_) );
AOI21X1 AOI21X1_906 ( .A(datapath_1_RegisterFile_regfile_mem_7__1_), .B(datapath_1_Instr_18_bF_buf24_), .C(_3588__bF_buf9), .Y(_3638_) );
OAI21X1 OAI21X1_1970 ( .A(_3637_), .B(datapath_1_Instr_18_bF_buf23_), .C(_3638_), .Y(_3639_) );
INVX1 INVX1_505 ( .A(datapath_1_RegisterFile_regfile_mem_2__1_), .Y(_3640_) );
AOI21X1 AOI21X1_907 ( .A(datapath_1_RegisterFile_regfile_mem_6__1_), .B(datapath_1_Instr_18_bF_buf22_), .C(datapath_1_Instr_16_bF_buf32_), .Y(_3641_) );
OAI21X1 OAI21X1_1971 ( .A(_3640_), .B(datapath_1_Instr_18_bF_buf21_), .C(_3641_), .Y(_3642_) );
NAND3X1 NAND3X1_1560 ( .A(datapath_1_Instr_17_bF_buf48_), .B(_3642_), .C(_3639_), .Y(_3643_) );
AOI21X1 AOI21X1_908 ( .A(_3636_), .B(_3643_), .C(datapath_1_Instr_19_bF_buf5_), .Y(_3644_) );
NAND2X1 NAND2X1_1383 ( .A(datapath_1_RegisterFile_regfile_mem_11__1_), .B(datapath_1_Instr_17_bF_buf47_), .Y(_3645_) );
NAND2X1 NAND2X1_1384 ( .A(datapath_1_RegisterFile_regfile_mem_9__1_), .B(_3566__bF_buf7), .Y(_3646_) );
NAND3X1 NAND3X1_1561 ( .A(datapath_1_Instr_16_bF_buf31_), .B(_3645_), .C(_3646_), .Y(_3647_) );
NAND2X1 NAND2X1_1385 ( .A(datapath_1_RegisterFile_regfile_mem_10__1_), .B(datapath_1_Instr_17_bF_buf46_), .Y(_3648_) );
AOI21X1 AOI21X1_909 ( .A(_3566__bF_buf7), .B(datapath_1_RegisterFile_regfile_mem_8__1_), .C(datapath_1_Instr_16_bF_buf30_), .Y(_3649_) );
NAND2X1 NAND2X1_1386 ( .A(_3648_), .B(_3649_), .Y(_3650_) );
NAND3X1 NAND3X1_1562 ( .A(_3567__bF_buf4), .B(_3647_), .C(_3650_), .Y(_3651_) );
NAND2X1 NAND2X1_1387 ( .A(datapath_1_RegisterFile_regfile_mem_15__1_), .B(datapath_1_Instr_17_bF_buf45_), .Y(_3652_) );
NAND2X1 NAND2X1_1388 ( .A(datapath_1_RegisterFile_regfile_mem_13__1_), .B(_3566__bF_buf0), .Y(_3653_) );
NAND3X1 NAND3X1_1563 ( .A(datapath_1_Instr_16_bF_buf29_), .B(_3652_), .C(_3653_), .Y(_3654_) );
NAND2X1 NAND2X1_1389 ( .A(datapath_1_RegisterFile_regfile_mem_14__1_), .B(datapath_1_Instr_17_bF_buf44_), .Y(_3655_) );
AOI21X1 AOI21X1_910 ( .A(_3566__bF_buf1), .B(datapath_1_RegisterFile_regfile_mem_12__1_), .C(datapath_1_Instr_16_bF_buf28_), .Y(_3656_) );
NAND2X1 NAND2X1_1390 ( .A(_3655_), .B(_3656_), .Y(_3657_) );
NAND3X1 NAND3X1_1564 ( .A(datapath_1_Instr_18_bF_buf20_), .B(_3654_), .C(_3657_), .Y(_3658_) );
AOI21X1 AOI21X1_911 ( .A(_3651_), .B(_3658_), .C(_3571__bF_buf1), .Y(_3659_) );
OAI21X1 OAI21X1_1972 ( .A(_3644_), .B(_3659_), .C(_3570__bF_buf3), .Y(_3660_) );
MUX2X1 MUX2X1_276 ( .A(datapath_1_RegisterFile_regfile_mem_17__1_), .B(datapath_1_RegisterFile_regfile_mem_16__1_), .S(datapath_1_Instr_16_bF_buf27_), .Y(_3661_) );
NOR2X1 NOR2X1_494 ( .A(datapath_1_RegisterFile_regfile_mem_19__1_), .B(_3588__bF_buf15), .Y(_3662_) );
OAI21X1 OAI21X1_1973 ( .A(datapath_1_RegisterFile_regfile_mem_18__1_), .B(datapath_1_Instr_16_bF_buf26_), .C(datapath_1_Instr_17_bF_buf43_), .Y(_3663_) );
OAI22X1 OAI22X1_266 ( .A(_3663_), .B(_3662_), .C(datapath_1_Instr_17_bF_buf42_), .D(_3661_), .Y(_3664_) );
NAND2X1 NAND2X1_1391 ( .A(_3567__bF_buf0), .B(_3664_), .Y(_3665_) );
MUX2X1 MUX2X1_277 ( .A(datapath_1_RegisterFile_regfile_mem_21__1_), .B(datapath_1_RegisterFile_regfile_mem_20__1_), .S(datapath_1_Instr_16_bF_buf25_), .Y(_3666_) );
NOR2X1 NOR2X1_495 ( .A(datapath_1_RegisterFile_regfile_mem_23__1_), .B(_3588__bF_buf39), .Y(_3667_) );
OAI21X1 OAI21X1_1974 ( .A(datapath_1_RegisterFile_regfile_mem_22__1_), .B(datapath_1_Instr_16_bF_buf24_), .C(datapath_1_Instr_17_bF_buf41_), .Y(_3668_) );
OAI22X1 OAI22X1_267 ( .A(_3668_), .B(_3667_), .C(datapath_1_Instr_17_bF_buf40_), .D(_3666_), .Y(_3669_) );
NAND2X1 NAND2X1_1392 ( .A(datapath_1_Instr_18_bF_buf19_), .B(_3669_), .Y(_3670_) );
AOI21X1 AOI21X1_912 ( .A(_3665_), .B(_3670_), .C(datapath_1_Instr_19_bF_buf4_), .Y(_3671_) );
AOI21X1 AOI21X1_913 ( .A(datapath_1_RegisterFile_regfile_mem_31__1_), .B(datapath_1_Instr_18_bF_buf18_), .C(_3588__bF_buf33), .Y(_3672_) );
OAI21X1 OAI21X1_1975 ( .A(_1969_), .B(datapath_1_Instr_18_bF_buf17_), .C(_3672_), .Y(_3673_) );
AOI21X1 AOI21X1_914 ( .A(datapath_1_RegisterFile_regfile_mem_30__1_), .B(datapath_1_Instr_18_bF_buf16_), .C(datapath_1_Instr_16_bF_buf23_), .Y(_3674_) );
OAI21X1 OAI21X1_1976 ( .A(_1972_), .B(datapath_1_Instr_18_bF_buf15_), .C(_3674_), .Y(_3675_) );
NAND3X1 NAND3X1_1565 ( .A(datapath_1_Instr_17_bF_buf39_), .B(_3675_), .C(_3673_), .Y(_3676_) );
AOI21X1 AOI21X1_915 ( .A(datapath_1_RegisterFile_regfile_mem_29__1_), .B(datapath_1_Instr_18_bF_buf14_), .C(_3588__bF_buf33), .Y(_3677_) );
OAI21X1 OAI21X1_1977 ( .A(_1976_), .B(datapath_1_Instr_18_bF_buf13_), .C(_3677_), .Y(_3678_) );
AOI21X1 AOI21X1_916 ( .A(datapath_1_RegisterFile_regfile_mem_28__1_), .B(datapath_1_Instr_18_bF_buf12_), .C(datapath_1_Instr_16_bF_buf22_), .Y(_3679_) );
OAI21X1 OAI21X1_1978 ( .A(_1979_), .B(datapath_1_Instr_18_bF_buf11_), .C(_3679_), .Y(_3680_) );
NAND3X1 NAND3X1_1566 ( .A(_3566__bF_buf10), .B(_3680_), .C(_3678_), .Y(_3681_) );
AOI21X1 AOI21X1_917 ( .A(_3676_), .B(_3681_), .C(_3571__bF_buf7), .Y(_3682_) );
OAI21X1 OAI21X1_1979 ( .A(_3682_), .B(_3671_), .C(datapath_1_Instr_20_bF_buf5_), .Y(_3683_) );
AOI22X1 AOI22X1_192 ( .A(_3565__bF_buf4), .B(_3569__bF_buf4), .C(_3660_), .D(_3683_), .Y(datapath_1_RD2_1_) );
MUX2X1 MUX2X1_278 ( .A(datapath_1_RegisterFile_regfile_mem_9__2_), .B(datapath_1_RegisterFile_regfile_mem_8__2_), .S(datapath_1_Instr_16_bF_buf21_), .Y(_3684_) );
NOR2X1 NOR2X1_496 ( .A(datapath_1_RegisterFile_regfile_mem_11__2_), .B(_3588__bF_buf1), .Y(_3685_) );
OAI21X1 OAI21X1_1980 ( .A(datapath_1_RegisterFile_regfile_mem_10__2_), .B(datapath_1_Instr_16_bF_buf20_), .C(datapath_1_Instr_17_bF_buf38_), .Y(_3686_) );
FILL FILL_0_0_0 ( );
FILL FILL_0_0_1 ( );
FILL FILL_0_0_2 ( );
FILL FILL_0_1_0 ( );
FILL FILL_0_1_1 ( );
FILL FILL_0_1_2 ( );
FILL FILL_0_2_0 ( );
FILL FILL_0_2_1 ( );
FILL FILL_0_2_2 ( );
FILL FILL_0_3_0 ( );
FILL FILL_0_3_1 ( );
FILL FILL_0_3_2 ( );
FILL FILL_0_4_0 ( );
FILL FILL_0_4_1 ( );
FILL FILL_0_4_2 ( );
FILL FILL_0_5_0 ( );
FILL FILL_0_5_1 ( );
FILL FILL_0_5_2 ( );
FILL FILL_0_6_0 ( );
FILL FILL_0_6_1 ( );
FILL FILL_0_6_2 ( );
FILL FILL_0_7_0 ( );
FILL FILL_0_7_1 ( );
FILL FILL_0_7_2 ( );
FILL FILL_0_8_0 ( );
FILL FILL_0_8_1 ( );
FILL FILL_0_8_2 ( );
FILL FILL_1_1 ( );
FILL FILL_1_2 ( );
FILL FILL_1_3 ( );
FILL FILL_1_0_0 ( );
FILL FILL_1_0_1 ( );
FILL FILL_1_0_2 ( );
FILL FILL_1_1_0 ( );
FILL FILL_1_1_1 ( );
FILL FILL_1_1_2 ( );
FILL FILL_1_2_0 ( );
FILL FILL_1_2_1 ( );
FILL FILL_1_2_2 ( );
FILL FILL_1_3_0 ( );
FILL FILL_1_3_1 ( );
FILL FILL_1_3_2 ( );
FILL FILL_1_4_0 ( );
FILL FILL_1_4_1 ( );
FILL FILL_1_4_2 ( );
FILL FILL_1_5_0 ( );
FILL FILL_1_5_1 ( );
FILL FILL_1_5_2 ( );
FILL FILL_1_6_0 ( );
FILL FILL_1_6_1 ( );
FILL FILL_1_6_2 ( );
FILL FILL_1_7_0 ( );
FILL FILL_1_7_1 ( );
FILL FILL_1_7_2 ( );
FILL FILL_1_8_0 ( );
FILL FILL_1_8_1 ( );
FILL FILL_1_8_2 ( );
FILL FILL_2_1 ( );
FILL FILL_2_2 ( );
FILL FILL_2_0_0 ( );
FILL FILL_2_0_1 ( );
FILL FILL_2_0_2 ( );
FILL FILL_2_1_0 ( );
FILL FILL_2_1_1 ( );
FILL FILL_2_1_2 ( );
FILL FILL_2_2_0 ( );
FILL FILL_2_2_1 ( );
FILL FILL_2_2_2 ( );
FILL FILL_2_3_0 ( );
FILL FILL_2_3_1 ( );
FILL FILL_2_3_2 ( );
FILL FILL_2_4_0 ( );
FILL FILL_2_4_1 ( );
FILL FILL_2_4_2 ( );
FILL FILL_2_5_0 ( );
FILL FILL_2_5_1 ( );
FILL FILL_2_5_2 ( );
FILL FILL_2_6_0 ( );
FILL FILL_2_6_1 ( );
FILL FILL_2_6_2 ( );
FILL FILL_2_7_0 ( );
FILL FILL_2_7_1 ( );
FILL FILL_2_7_2 ( );
FILL FILL_2_8_0 ( );
FILL FILL_2_8_1 ( );
FILL FILL_2_8_2 ( );
FILL FILL_3_1 ( );
FILL FILL_3_2 ( );
FILL FILL_3_3 ( );
FILL FILL_3_4 ( );
FILL FILL_3_0_0 ( );
FILL FILL_3_0_1 ( );
FILL FILL_3_0_2 ( );
FILL FILL_3_1_0 ( );
FILL FILL_3_1_1 ( );
FILL FILL_3_1_2 ( );
FILL FILL_3_2_0 ( );
FILL FILL_3_2_1 ( );
FILL FILL_3_2_2 ( );
FILL FILL_3_3_0 ( );
FILL FILL_3_3_1 ( );
FILL FILL_3_3_2 ( );
FILL FILL_3_4_0 ( );
FILL FILL_3_4_1 ( );
FILL FILL_3_4_2 ( );
FILL FILL_3_5_0 ( );
FILL FILL_3_5_1 ( );
FILL FILL_3_5_2 ( );
FILL FILL_3_6_0 ( );
FILL FILL_3_6_1 ( );
FILL FILL_3_6_2 ( );
FILL FILL_3_7_0 ( );
FILL FILL_3_7_1 ( );
FILL FILL_3_7_2 ( );
FILL FILL_3_8_0 ( );
FILL FILL_3_8_1 ( );
FILL FILL_3_8_2 ( );
FILL FILL_4_1 ( );
FILL FILL_4_2 ( );
FILL FILL_4_3 ( );
FILL FILL_4_0_0 ( );
FILL FILL_4_0_1 ( );
FILL FILL_4_0_2 ( );
FILL FILL_4_1_0 ( );
FILL FILL_4_1_1 ( );
FILL FILL_4_1_2 ( );
FILL FILL_4_2_0 ( );
FILL FILL_4_2_1 ( );
FILL FILL_4_2_2 ( );
FILL FILL_4_3_0 ( );
FILL FILL_4_3_1 ( );
FILL FILL_4_3_2 ( );
FILL FILL_4_4_0 ( );
FILL FILL_4_4_1 ( );
FILL FILL_4_4_2 ( );
FILL FILL_4_5_0 ( );
FILL FILL_4_5_1 ( );
FILL FILL_4_5_2 ( );
FILL FILL_4_6_0 ( );
FILL FILL_4_6_1 ( );
FILL FILL_4_6_2 ( );
FILL FILL_4_7_0 ( );
FILL FILL_4_7_1 ( );
FILL FILL_4_7_2 ( );
FILL FILL_4_8_0 ( );
FILL FILL_4_8_1 ( );
FILL FILL_4_8_2 ( );
FILL FILL_5_1 ( );
FILL FILL_5_0_0 ( );
FILL FILL_5_0_1 ( );
FILL FILL_5_0_2 ( );
FILL FILL_5_1_0 ( );
FILL FILL_5_1_1 ( );
FILL FILL_5_1_2 ( );
FILL FILL_5_2_0 ( );
FILL FILL_5_2_1 ( );
FILL FILL_5_2_2 ( );
FILL FILL_5_3_0 ( );
FILL FILL_5_3_1 ( );
FILL FILL_5_3_2 ( );
FILL FILL_5_4_0 ( );
FILL FILL_5_4_1 ( );
FILL FILL_5_4_2 ( );
FILL FILL_5_5_0 ( );
FILL FILL_5_5_1 ( );
FILL FILL_5_5_2 ( );
FILL FILL_5_6_0 ( );
FILL FILL_5_6_1 ( );
FILL FILL_5_6_2 ( );
FILL FILL_5_7_0 ( );
FILL FILL_5_7_1 ( );
FILL FILL_5_7_2 ( );
FILL FILL_5_8_0 ( );
FILL FILL_5_8_1 ( );
FILL FILL_5_8_2 ( );
FILL FILL_6_0_0 ( );
FILL FILL_6_0_1 ( );
FILL FILL_6_0_2 ( );
FILL FILL_6_1_0 ( );
FILL FILL_6_1_1 ( );
FILL FILL_6_1_2 ( );
FILL FILL_6_2_0 ( );
FILL FILL_6_2_1 ( );
FILL FILL_6_2_2 ( );
FILL FILL_6_3_0 ( );
FILL FILL_6_3_1 ( );
FILL FILL_6_3_2 ( );
FILL FILL_6_4_0 ( );
FILL FILL_6_4_1 ( );
FILL FILL_6_4_2 ( );
FILL FILL_6_5_0 ( );
FILL FILL_6_5_1 ( );
FILL FILL_6_5_2 ( );
FILL FILL_6_6_0 ( );
FILL FILL_6_6_1 ( );
FILL FILL_6_6_2 ( );
FILL FILL_6_7_0 ( );
FILL FILL_6_7_1 ( );
FILL FILL_6_7_2 ( );
FILL FILL_6_8_0 ( );
FILL FILL_6_8_1 ( );
FILL FILL_6_8_2 ( );
FILL FILL_7_1 ( );
FILL FILL_7_2 ( );
FILL FILL_7_3 ( );
FILL FILL_7_4 ( );
FILL FILL_7_0_0 ( );
FILL FILL_7_0_1 ( );
FILL FILL_7_0_2 ( );
FILL FILL_7_1_0 ( );
FILL FILL_7_1_1 ( );
FILL FILL_7_1_2 ( );
FILL FILL_7_2_0 ( );
FILL FILL_7_2_1 ( );
FILL FILL_7_2_2 ( );
FILL FILL_7_3_0 ( );
FILL FILL_7_3_1 ( );
FILL FILL_7_3_2 ( );
FILL FILL_7_4_0 ( );
FILL FILL_7_4_1 ( );
FILL FILL_7_4_2 ( );
FILL FILL_7_5_0 ( );
FILL FILL_7_5_1 ( );
FILL FILL_7_5_2 ( );
FILL FILL_7_6_0 ( );
FILL FILL_7_6_1 ( );
FILL FILL_7_6_2 ( );
FILL FILL_7_7_0 ( );
FILL FILL_7_7_1 ( );
FILL FILL_7_7_2 ( );
FILL FILL_7_8_0 ( );
FILL FILL_7_8_1 ( );
FILL FILL_7_8_2 ( );
FILL FILL_8_1 ( );
FILL FILL_8_2 ( );
FILL FILL_8_3 ( );
FILL FILL_8_4 ( );
FILL FILL_8_0_0 ( );
FILL FILL_8_0_1 ( );
FILL FILL_8_0_2 ( );
FILL FILL_8_1_0 ( );
FILL FILL_8_1_1 ( );
FILL FILL_8_1_2 ( );
FILL FILL_8_2_0 ( );
FILL FILL_8_2_1 ( );
FILL FILL_8_2_2 ( );
FILL FILL_8_3_0 ( );
FILL FILL_8_3_1 ( );
FILL FILL_8_3_2 ( );
FILL FILL_8_4_0 ( );
FILL FILL_8_4_1 ( );
FILL FILL_8_4_2 ( );
FILL FILL_8_5_0 ( );
FILL FILL_8_5_1 ( );
FILL FILL_8_5_2 ( );
FILL FILL_8_6_0 ( );
FILL FILL_8_6_1 ( );
FILL FILL_8_6_2 ( );
FILL FILL_8_7_0 ( );
FILL FILL_8_7_1 ( );
FILL FILL_8_7_2 ( );
FILL FILL_8_8_0 ( );
FILL FILL_8_8_1 ( );
FILL FILL_8_8_2 ( );
FILL FILL_9_1 ( );
FILL FILL_9_0_0 ( );
FILL FILL_9_0_1 ( );
FILL FILL_9_0_2 ( );
FILL FILL_9_1_0 ( );
FILL FILL_9_1_1 ( );
FILL FILL_9_1_2 ( );
FILL FILL_9_2_0 ( );
FILL FILL_9_2_1 ( );
FILL FILL_9_2_2 ( );
FILL FILL_9_3_0 ( );
FILL FILL_9_3_1 ( );
FILL FILL_9_3_2 ( );
FILL FILL_9_4_0 ( );
FILL FILL_9_4_1 ( );
FILL FILL_9_4_2 ( );
FILL FILL_9_5_0 ( );
FILL FILL_9_5_1 ( );
FILL FILL_9_5_2 ( );
FILL FILL_9_6_0 ( );
FILL FILL_9_6_1 ( );
FILL FILL_9_6_2 ( );
FILL FILL_9_7_0 ( );
FILL FILL_9_7_1 ( );
FILL FILL_9_7_2 ( );
FILL FILL_9_8_0 ( );
FILL FILL_9_8_1 ( );
FILL FILL_9_8_2 ( );
FILL FILL_10_1 ( );
FILL FILL_10_2 ( );
FILL FILL_10_3 ( );
FILL FILL_10_4 ( );
FILL FILL_10_0_0 ( );
FILL FILL_10_0_1 ( );
FILL FILL_10_0_2 ( );
FILL FILL_10_1_0 ( );
FILL FILL_10_1_1 ( );
FILL FILL_10_1_2 ( );
FILL FILL_10_2_0 ( );
FILL FILL_10_2_1 ( );
FILL FILL_10_2_2 ( );
FILL FILL_10_3_0 ( );
FILL FILL_10_3_1 ( );
FILL FILL_10_3_2 ( );
FILL FILL_10_4_0 ( );
FILL FILL_10_4_1 ( );
FILL FILL_10_4_2 ( );
FILL FILL_10_5_0 ( );
FILL FILL_10_5_1 ( );
FILL FILL_10_5_2 ( );
FILL FILL_10_6_0 ( );
FILL FILL_10_6_1 ( );
FILL FILL_10_6_2 ( );
FILL FILL_10_7_0 ( );
FILL FILL_10_7_1 ( );
FILL FILL_10_7_2 ( );
FILL FILL_10_8_0 ( );
FILL FILL_10_8_1 ( );
FILL FILL_10_8_2 ( );
FILL FILL_11_1 ( );
FILL FILL_11_0_0 ( );
FILL FILL_11_0_1 ( );
FILL FILL_11_0_2 ( );
FILL FILL_11_1_0 ( );
FILL FILL_11_1_1 ( );
FILL FILL_11_1_2 ( );
FILL FILL_11_2_0 ( );
FILL FILL_11_2_1 ( );
FILL FILL_11_2_2 ( );
FILL FILL_11_3_0 ( );
FILL FILL_11_3_1 ( );
FILL FILL_11_3_2 ( );
FILL FILL_11_4_0 ( );
FILL FILL_11_4_1 ( );
FILL FILL_11_4_2 ( );
FILL FILL_11_5_0 ( );
FILL FILL_11_5_1 ( );
FILL FILL_11_5_2 ( );
FILL FILL_11_6_0 ( );
FILL FILL_11_6_1 ( );
FILL FILL_11_6_2 ( );
FILL FILL_11_7_0 ( );
FILL FILL_11_7_1 ( );
FILL FILL_11_7_2 ( );
FILL FILL_11_8_0 ( );
FILL FILL_11_8_1 ( );
FILL FILL_11_8_2 ( );
FILL FILL_12_1 ( );
FILL FILL_12_2 ( );
FILL FILL_12_3 ( );
FILL FILL_12_0_0 ( );
FILL FILL_12_0_1 ( );
FILL FILL_12_0_2 ( );
FILL FILL_12_1_0 ( );
FILL FILL_12_1_1 ( );
FILL FILL_12_1_2 ( );
FILL FILL_12_2_0 ( );
FILL FILL_12_2_1 ( );
FILL FILL_12_2_2 ( );
FILL FILL_12_3_0 ( );
FILL FILL_12_3_1 ( );
FILL FILL_12_3_2 ( );
FILL FILL_12_4_0 ( );
FILL FILL_12_4_1 ( );
FILL FILL_12_4_2 ( );
FILL FILL_12_5_0 ( );
FILL FILL_12_5_1 ( );
FILL FILL_12_5_2 ( );
FILL FILL_12_6_0 ( );
FILL FILL_12_6_1 ( );
FILL FILL_12_6_2 ( );
FILL FILL_12_7_0 ( );
FILL FILL_12_7_1 ( );
FILL FILL_12_7_2 ( );
FILL FILL_12_8_0 ( );
FILL FILL_12_8_1 ( );
FILL FILL_12_8_2 ( );
FILL FILL_13_1 ( );
FILL FILL_13_2 ( );
FILL FILL_13_0_0 ( );
FILL FILL_13_0_1 ( );
FILL FILL_13_0_2 ( );
FILL FILL_13_1_0 ( );
FILL FILL_13_1_1 ( );
FILL FILL_13_1_2 ( );
FILL FILL_13_2_0 ( );
FILL FILL_13_2_1 ( );
FILL FILL_13_2_2 ( );
FILL FILL_13_3_0 ( );
FILL FILL_13_3_1 ( );
FILL FILL_13_3_2 ( );
FILL FILL_13_4_0 ( );
FILL FILL_13_4_1 ( );
FILL FILL_13_4_2 ( );
FILL FILL_13_5_0 ( );
FILL FILL_13_5_1 ( );
FILL FILL_13_5_2 ( );
FILL FILL_13_6_0 ( );
FILL FILL_13_6_1 ( );
FILL FILL_13_6_2 ( );
FILL FILL_13_7_0 ( );
FILL FILL_13_7_1 ( );
FILL FILL_13_7_2 ( );
FILL FILL_13_8_0 ( );
FILL FILL_13_8_1 ( );
FILL FILL_13_8_2 ( );
FILL FILL_14_1 ( );
FILL FILL_14_2 ( );
FILL FILL_14_3 ( );
FILL FILL_14_4 ( );
FILL FILL_14_0_0 ( );
FILL FILL_14_0_1 ( );
FILL FILL_14_0_2 ( );
FILL FILL_14_1_0 ( );
FILL FILL_14_1_1 ( );
FILL FILL_14_1_2 ( );
FILL FILL_14_2_0 ( );
FILL FILL_14_2_1 ( );
FILL FILL_14_2_2 ( );
FILL FILL_14_3_0 ( );
FILL FILL_14_3_1 ( );
FILL FILL_14_3_2 ( );
FILL FILL_14_4_0 ( );
FILL FILL_14_4_1 ( );
FILL FILL_14_4_2 ( );
FILL FILL_14_5_0 ( );
FILL FILL_14_5_1 ( );
FILL FILL_14_5_2 ( );
FILL FILL_14_6_0 ( );
FILL FILL_14_6_1 ( );
FILL FILL_14_6_2 ( );
FILL FILL_14_7_0 ( );
FILL FILL_14_7_1 ( );
FILL FILL_14_7_2 ( );
FILL FILL_14_8_0 ( );
FILL FILL_14_8_1 ( );
FILL FILL_14_8_2 ( );
FILL FILL_15_1 ( );
FILL FILL_15_0_0 ( );
FILL FILL_15_0_1 ( );
FILL FILL_15_0_2 ( );
FILL FILL_15_1_0 ( );
FILL FILL_15_1_1 ( );
FILL FILL_15_1_2 ( );
FILL FILL_15_2_0 ( );
FILL FILL_15_2_1 ( );
FILL FILL_15_2_2 ( );
FILL FILL_15_3_0 ( );
FILL FILL_15_3_1 ( );
FILL FILL_15_3_2 ( );
FILL FILL_15_4_0 ( );
FILL FILL_15_4_1 ( );
FILL FILL_15_4_2 ( );
FILL FILL_15_5_0 ( );
FILL FILL_15_5_1 ( );
FILL FILL_15_5_2 ( );
FILL FILL_15_6_0 ( );
FILL FILL_15_6_1 ( );
FILL FILL_15_6_2 ( );
FILL FILL_15_7_0 ( );
FILL FILL_15_7_1 ( );
FILL FILL_15_7_2 ( );
FILL FILL_15_8_0 ( );
FILL FILL_15_8_1 ( );
FILL FILL_15_8_2 ( );
FILL FILL_16_1 ( );
FILL FILL_16_2 ( );
FILL FILL_16_3 ( );
FILL FILL_16_0_0 ( );
FILL FILL_16_0_1 ( );
FILL FILL_16_0_2 ( );
FILL FILL_16_1_0 ( );
FILL FILL_16_1_1 ( );
FILL FILL_16_1_2 ( );
FILL FILL_16_2_0 ( );
FILL FILL_16_2_1 ( );
FILL FILL_16_2_2 ( );
FILL FILL_16_3_0 ( );
FILL FILL_16_3_1 ( );
FILL FILL_16_3_2 ( );
FILL FILL_16_4_0 ( );
FILL FILL_16_4_1 ( );
FILL FILL_16_4_2 ( );
FILL FILL_16_5_0 ( );
FILL FILL_16_5_1 ( );
FILL FILL_16_5_2 ( );
FILL FILL_16_6_0 ( );
FILL FILL_16_6_1 ( );
FILL FILL_16_6_2 ( );
FILL FILL_16_7_0 ( );
FILL FILL_16_7_1 ( );
FILL FILL_16_7_2 ( );
FILL FILL_16_8_0 ( );
FILL FILL_16_8_1 ( );
FILL FILL_16_8_2 ( );
FILL FILL_17_1 ( );
FILL FILL_17_2 ( );
FILL FILL_17_3 ( );
FILL FILL_17_4 ( );
FILL FILL_17_0_0 ( );
FILL FILL_17_0_1 ( );
FILL FILL_17_0_2 ( );
FILL FILL_17_1_0 ( );
FILL FILL_17_1_1 ( );
FILL FILL_17_1_2 ( );
FILL FILL_17_2_0 ( );
FILL FILL_17_2_1 ( );
FILL FILL_17_2_2 ( );
FILL FILL_17_3_0 ( );
FILL FILL_17_3_1 ( );
FILL FILL_17_3_2 ( );
FILL FILL_17_4_0 ( );
FILL FILL_17_4_1 ( );
FILL FILL_17_4_2 ( );
FILL FILL_17_5_0 ( );
FILL FILL_17_5_1 ( );
FILL FILL_17_5_2 ( );
FILL FILL_17_6_0 ( );
FILL FILL_17_6_1 ( );
FILL FILL_17_6_2 ( );
FILL FILL_17_7_0 ( );
FILL FILL_17_7_1 ( );
FILL FILL_17_7_2 ( );
FILL FILL_17_8_0 ( );
FILL FILL_17_8_1 ( );
FILL FILL_17_8_2 ( );
FILL FILL_18_0_0 ( );
FILL FILL_18_0_1 ( );
FILL FILL_18_0_2 ( );
FILL FILL_18_1_0 ( );
FILL FILL_18_1_1 ( );
FILL FILL_18_1_2 ( );
FILL FILL_18_2_0 ( );
FILL FILL_18_2_1 ( );
FILL FILL_18_2_2 ( );
FILL FILL_18_3_0 ( );
FILL FILL_18_3_1 ( );
FILL FILL_18_3_2 ( );
FILL FILL_18_4_0 ( );
FILL FILL_18_4_1 ( );
FILL FILL_18_4_2 ( );
FILL FILL_18_5_0 ( );
FILL FILL_18_5_1 ( );
FILL FILL_18_5_2 ( );
FILL FILL_18_6_0 ( );
FILL FILL_18_6_1 ( );
FILL FILL_18_6_2 ( );
FILL FILL_18_7_0 ( );
FILL FILL_18_7_1 ( );
FILL FILL_18_7_2 ( );
FILL FILL_18_8_0 ( );
FILL FILL_18_8_1 ( );
FILL FILL_18_8_2 ( );
FILL FILL_19_1 ( );
FILL FILL_19_2 ( );
FILL FILL_19_3 ( );
FILL FILL_19_0_0 ( );
FILL FILL_19_0_1 ( );
FILL FILL_19_0_2 ( );
FILL FILL_19_1_0 ( );
FILL FILL_19_1_1 ( );
FILL FILL_19_1_2 ( );
FILL FILL_19_2_0 ( );
FILL FILL_19_2_1 ( );
FILL FILL_19_2_2 ( );
FILL FILL_19_3_0 ( );
FILL FILL_19_3_1 ( );
FILL FILL_19_3_2 ( );
FILL FILL_19_4_0 ( );
FILL FILL_19_4_1 ( );
FILL FILL_19_4_2 ( );
FILL FILL_19_5_0 ( );
FILL FILL_19_5_1 ( );
FILL FILL_19_5_2 ( );
FILL FILL_19_6_0 ( );
FILL FILL_19_6_1 ( );
FILL FILL_19_6_2 ( );
FILL FILL_19_7_0 ( );
FILL FILL_19_7_1 ( );
FILL FILL_19_7_2 ( );
FILL FILL_19_8_0 ( );
FILL FILL_19_8_1 ( );
FILL FILL_19_8_2 ( );
FILL FILL_20_1 ( );
FILL FILL_20_0_0 ( );
FILL FILL_20_0_1 ( );
FILL FILL_20_0_2 ( );
FILL FILL_20_1_0 ( );
FILL FILL_20_1_1 ( );
FILL FILL_20_1_2 ( );
FILL FILL_20_2_0 ( );
FILL FILL_20_2_1 ( );
FILL FILL_20_2_2 ( );
FILL FILL_20_3_0 ( );
FILL FILL_20_3_1 ( );
FILL FILL_20_3_2 ( );
FILL FILL_20_4_0 ( );
FILL FILL_20_4_1 ( );
FILL FILL_20_4_2 ( );
FILL FILL_20_5_0 ( );
FILL FILL_20_5_1 ( );
FILL FILL_20_5_2 ( );
FILL FILL_20_6_0 ( );
FILL FILL_20_6_1 ( );
FILL FILL_20_6_2 ( );
FILL FILL_20_7_0 ( );
FILL FILL_20_7_1 ( );
FILL FILL_20_7_2 ( );
FILL FILL_20_8_0 ( );
FILL FILL_20_8_1 ( );
FILL FILL_20_8_2 ( );
FILL FILL_21_1 ( );
FILL FILL_21_2 ( );
FILL FILL_21_0_0 ( );
FILL FILL_21_0_1 ( );
FILL FILL_21_0_2 ( );
FILL FILL_21_1_0 ( );
FILL FILL_21_1_1 ( );
FILL FILL_21_1_2 ( );
FILL FILL_21_2_0 ( );
FILL FILL_21_2_1 ( );
FILL FILL_21_2_2 ( );
FILL FILL_21_3_0 ( );
FILL FILL_21_3_1 ( );
FILL FILL_21_3_2 ( );
FILL FILL_21_4_0 ( );
FILL FILL_21_4_1 ( );
FILL FILL_21_4_2 ( );
FILL FILL_21_5_0 ( );
FILL FILL_21_5_1 ( );
FILL FILL_21_5_2 ( );
FILL FILL_21_6_0 ( );
FILL FILL_21_6_1 ( );
FILL FILL_21_6_2 ( );
FILL FILL_21_7_0 ( );
FILL FILL_21_7_1 ( );
FILL FILL_21_7_2 ( );
FILL FILL_21_8_0 ( );
FILL FILL_21_8_1 ( );
FILL FILL_21_8_2 ( );
FILL FILL_22_1 ( );
FILL FILL_22_2 ( );
FILL FILL_22_0_0 ( );
FILL FILL_22_0_1 ( );
FILL FILL_22_0_2 ( );
FILL FILL_22_1_0 ( );
FILL FILL_22_1_1 ( );
FILL FILL_22_1_2 ( );
FILL FILL_22_2_0 ( );
FILL FILL_22_2_1 ( );
FILL FILL_22_2_2 ( );
FILL FILL_22_3_0 ( );
FILL FILL_22_3_1 ( );
FILL FILL_22_3_2 ( );
FILL FILL_22_4_0 ( );
FILL FILL_22_4_1 ( );
FILL FILL_22_4_2 ( );
FILL FILL_22_5_0 ( );
FILL FILL_22_5_1 ( );
FILL FILL_22_5_2 ( );
FILL FILL_22_6_0 ( );
FILL FILL_22_6_1 ( );
FILL FILL_22_6_2 ( );
FILL FILL_22_7_0 ( );
FILL FILL_22_7_1 ( );
FILL FILL_22_7_2 ( );
FILL FILL_22_8_0 ( );
FILL FILL_22_8_1 ( );
FILL FILL_22_8_2 ( );
FILL FILL_23_1 ( );
FILL FILL_23_2 ( );
FILL FILL_23_0_0 ( );
FILL FILL_23_0_1 ( );
FILL FILL_23_0_2 ( );
FILL FILL_23_1_0 ( );
FILL FILL_23_1_1 ( );
FILL FILL_23_1_2 ( );
FILL FILL_23_2_0 ( );
FILL FILL_23_2_1 ( );
FILL FILL_23_2_2 ( );
FILL FILL_23_3_0 ( );
FILL FILL_23_3_1 ( );
FILL FILL_23_3_2 ( );
FILL FILL_23_4_0 ( );
FILL FILL_23_4_1 ( );
FILL FILL_23_4_2 ( );
FILL FILL_23_5_0 ( );
FILL FILL_23_5_1 ( );
FILL FILL_23_5_2 ( );
FILL FILL_23_6_0 ( );
FILL FILL_23_6_1 ( );
FILL FILL_23_6_2 ( );
FILL FILL_23_7_0 ( );
FILL FILL_23_7_1 ( );
FILL FILL_23_7_2 ( );
FILL FILL_23_8_0 ( );
FILL FILL_23_8_1 ( );
FILL FILL_23_8_2 ( );
FILL FILL_24_0_0 ( );
FILL FILL_24_0_1 ( );
FILL FILL_24_0_2 ( );
FILL FILL_24_1_0 ( );
FILL FILL_24_1_1 ( );
FILL FILL_24_1_2 ( );
FILL FILL_24_2_0 ( );
FILL FILL_24_2_1 ( );
FILL FILL_24_2_2 ( );
FILL FILL_24_3_0 ( );
FILL FILL_24_3_1 ( );
FILL FILL_24_3_2 ( );
FILL FILL_24_4_0 ( );
FILL FILL_24_4_1 ( );
FILL FILL_24_4_2 ( );
FILL FILL_24_5_0 ( );
FILL FILL_24_5_1 ( );
FILL FILL_24_5_2 ( );
FILL FILL_24_6_0 ( );
FILL FILL_24_6_1 ( );
FILL FILL_24_6_2 ( );
FILL FILL_24_7_0 ( );
FILL FILL_24_7_1 ( );
FILL FILL_24_7_2 ( );
FILL FILL_24_8_0 ( );
FILL FILL_24_8_1 ( );
FILL FILL_24_8_2 ( );
FILL FILL_25_1 ( );
FILL FILL_25_2 ( );
FILL FILL_25_3 ( );
FILL FILL_25_0_0 ( );
FILL FILL_25_0_1 ( );
FILL FILL_25_0_2 ( );
FILL FILL_25_1_0 ( );
FILL FILL_25_1_1 ( );
FILL FILL_25_1_2 ( );
FILL FILL_25_2_0 ( );
FILL FILL_25_2_1 ( );
FILL FILL_25_2_2 ( );
FILL FILL_25_3_0 ( );
FILL FILL_25_3_1 ( );
FILL FILL_25_3_2 ( );
FILL FILL_25_4_0 ( );
FILL FILL_25_4_1 ( );
FILL FILL_25_4_2 ( );
FILL FILL_25_5_0 ( );
FILL FILL_25_5_1 ( );
FILL FILL_25_5_2 ( );
FILL FILL_25_6_0 ( );
FILL FILL_25_6_1 ( );
FILL FILL_25_6_2 ( );
FILL FILL_25_7_0 ( );
FILL FILL_25_7_1 ( );
FILL FILL_25_7_2 ( );
FILL FILL_25_8_0 ( );
FILL FILL_25_8_1 ( );
FILL FILL_25_8_2 ( );
FILL FILL_26_1 ( );
FILL FILL_26_2 ( );
FILL FILL_26_0_0 ( );
FILL FILL_26_0_1 ( );
FILL FILL_26_0_2 ( );
FILL FILL_26_1_0 ( );
FILL FILL_26_1_1 ( );
FILL FILL_26_1_2 ( );
FILL FILL_26_2_0 ( );
FILL FILL_26_2_1 ( );
FILL FILL_26_2_2 ( );
FILL FILL_26_3_0 ( );
FILL FILL_26_3_1 ( );
FILL FILL_26_3_2 ( );
FILL FILL_26_4_0 ( );
FILL FILL_26_4_1 ( );
FILL FILL_26_4_2 ( );
FILL FILL_26_5_0 ( );
FILL FILL_26_5_1 ( );
FILL FILL_26_5_2 ( );
FILL FILL_26_6_0 ( );
FILL FILL_26_6_1 ( );
FILL FILL_26_6_2 ( );
FILL FILL_26_7_0 ( );
FILL FILL_26_7_1 ( );
FILL FILL_26_7_2 ( );
FILL FILL_26_8_0 ( );
FILL FILL_26_8_1 ( );
FILL FILL_26_8_2 ( );
FILL FILL_27_1 ( );
FILL FILL_27_2 ( );
FILL FILL_27_3 ( );
FILL FILL_27_0_0 ( );
FILL FILL_27_0_1 ( );
FILL FILL_27_0_2 ( );
FILL FILL_27_1_0 ( );
FILL FILL_27_1_1 ( );
FILL FILL_27_1_2 ( );
FILL FILL_27_2_0 ( );
FILL FILL_27_2_1 ( );
FILL FILL_27_2_2 ( );
FILL FILL_27_3_0 ( );
FILL FILL_27_3_1 ( );
FILL FILL_27_3_2 ( );
FILL FILL_27_4_0 ( );
FILL FILL_27_4_1 ( );
FILL FILL_27_4_2 ( );
FILL FILL_27_5_0 ( );
FILL FILL_27_5_1 ( );
FILL FILL_27_5_2 ( );
FILL FILL_27_6_0 ( );
FILL FILL_27_6_1 ( );
FILL FILL_27_6_2 ( );
FILL FILL_27_7_0 ( );
FILL FILL_27_7_1 ( );
FILL FILL_27_7_2 ( );
FILL FILL_27_8_0 ( );
FILL FILL_27_8_1 ( );
FILL FILL_27_8_2 ( );
FILL FILL_28_1 ( );
FILL FILL_28_2 ( );
FILL FILL_28_0_0 ( );
FILL FILL_28_0_1 ( );
FILL FILL_28_0_2 ( );
FILL FILL_28_1_0 ( );
FILL FILL_28_1_1 ( );
FILL FILL_28_1_2 ( );
FILL FILL_28_2_0 ( );
FILL FILL_28_2_1 ( );
FILL FILL_28_2_2 ( );
FILL FILL_28_3_0 ( );
FILL FILL_28_3_1 ( );
FILL FILL_28_3_2 ( );
FILL FILL_28_4_0 ( );
FILL FILL_28_4_1 ( );
FILL FILL_28_4_2 ( );
FILL FILL_28_5_0 ( );
FILL FILL_28_5_1 ( );
FILL FILL_28_5_2 ( );
FILL FILL_28_6_0 ( );
FILL FILL_28_6_1 ( );
FILL FILL_28_6_2 ( );
FILL FILL_28_7_0 ( );
FILL FILL_28_7_1 ( );
FILL FILL_28_7_2 ( );
FILL FILL_28_8_0 ( );
FILL FILL_28_8_1 ( );
FILL FILL_28_8_2 ( );
FILL FILL_29_1 ( );
FILL FILL_29_2 ( );
FILL FILL_29_3 ( );
FILL FILL_29_0_0 ( );
FILL FILL_29_0_1 ( );
FILL FILL_29_0_2 ( );
FILL FILL_29_1_0 ( );
FILL FILL_29_1_1 ( );
FILL FILL_29_1_2 ( );
FILL FILL_29_2_0 ( );
FILL FILL_29_2_1 ( );
FILL FILL_29_2_2 ( );
FILL FILL_29_3_0 ( );
FILL FILL_29_3_1 ( );
FILL FILL_29_3_2 ( );
FILL FILL_29_4_0 ( );
FILL FILL_29_4_1 ( );
FILL FILL_29_4_2 ( );
FILL FILL_29_5_0 ( );
FILL FILL_29_5_1 ( );
FILL FILL_29_5_2 ( );
FILL FILL_29_6_0 ( );
FILL FILL_29_6_1 ( );
FILL FILL_29_6_2 ( );
FILL FILL_29_7_0 ( );
FILL FILL_29_7_1 ( );
FILL FILL_29_7_2 ( );
FILL FILL_29_8_0 ( );
FILL FILL_29_8_1 ( );
FILL FILL_29_8_2 ( );
FILL FILL_30_1 ( );
FILL FILL_30_2 ( );
FILL FILL_30_0_0 ( );
FILL FILL_30_0_1 ( );
FILL FILL_30_0_2 ( );
FILL FILL_30_1_0 ( );
FILL FILL_30_1_1 ( );
FILL FILL_30_1_2 ( );
FILL FILL_30_2_0 ( );
FILL FILL_30_2_1 ( );
FILL FILL_30_2_2 ( );
FILL FILL_30_3_0 ( );
FILL FILL_30_3_1 ( );
FILL FILL_30_3_2 ( );
FILL FILL_30_4_0 ( );
FILL FILL_30_4_1 ( );
FILL FILL_30_4_2 ( );
FILL FILL_30_5_0 ( );
FILL FILL_30_5_1 ( );
FILL FILL_30_5_2 ( );
FILL FILL_30_6_0 ( );
FILL FILL_30_6_1 ( );
FILL FILL_30_6_2 ( );
FILL FILL_30_7_0 ( );
FILL FILL_30_7_1 ( );
FILL FILL_30_7_2 ( );
FILL FILL_30_8_0 ( );
FILL FILL_30_8_1 ( );
FILL FILL_30_8_2 ( );
FILL FILL_31_1 ( );
FILL FILL_31_0_0 ( );
FILL FILL_31_0_1 ( );
FILL FILL_31_0_2 ( );
FILL FILL_31_1_0 ( );
FILL FILL_31_1_1 ( );
FILL FILL_31_1_2 ( );
FILL FILL_31_2_0 ( );
FILL FILL_31_2_1 ( );
FILL FILL_31_2_2 ( );
FILL FILL_31_3_0 ( );
FILL FILL_31_3_1 ( );
FILL FILL_31_3_2 ( );
FILL FILL_31_4_0 ( );
FILL FILL_31_4_1 ( );
FILL FILL_31_4_2 ( );
FILL FILL_31_5_0 ( );
FILL FILL_31_5_1 ( );
FILL FILL_31_5_2 ( );
FILL FILL_31_6_0 ( );
FILL FILL_31_6_1 ( );
FILL FILL_31_6_2 ( );
FILL FILL_31_7_0 ( );
FILL FILL_31_7_1 ( );
FILL FILL_31_7_2 ( );
FILL FILL_31_8_0 ( );
FILL FILL_31_8_1 ( );
FILL FILL_31_8_2 ( );
FILL FILL_32_1 ( );
FILL FILL_32_2 ( );
FILL FILL_32_3 ( );
FILL FILL_32_4 ( );
FILL FILL_32_0_0 ( );
FILL FILL_32_0_1 ( );
FILL FILL_32_0_2 ( );
FILL FILL_32_1_0 ( );
FILL FILL_32_1_1 ( );
FILL FILL_32_1_2 ( );
FILL FILL_32_2_0 ( );
FILL FILL_32_2_1 ( );
FILL FILL_32_2_2 ( );
FILL FILL_32_3_0 ( );
FILL FILL_32_3_1 ( );
FILL FILL_32_3_2 ( );
FILL FILL_32_4_0 ( );
FILL FILL_32_4_1 ( );
FILL FILL_32_4_2 ( );
FILL FILL_32_5_0 ( );
FILL FILL_32_5_1 ( );
FILL FILL_32_5_2 ( );
FILL FILL_32_6_0 ( );
FILL FILL_32_6_1 ( );
FILL FILL_32_6_2 ( );
FILL FILL_32_7_0 ( );
FILL FILL_32_7_1 ( );
FILL FILL_32_7_2 ( );
FILL FILL_32_8_0 ( );
FILL FILL_32_8_1 ( );
FILL FILL_32_8_2 ( );
FILL FILL_33_1 ( );
FILL FILL_33_2 ( );
FILL FILL_33_3 ( );
FILL FILL_33_4 ( );
FILL FILL_33_0_0 ( );
FILL FILL_33_0_1 ( );
FILL FILL_33_0_2 ( );
FILL FILL_33_1_0 ( );
FILL FILL_33_1_1 ( );
FILL FILL_33_1_2 ( );
FILL FILL_33_2_0 ( );
FILL FILL_33_2_1 ( );
FILL FILL_33_2_2 ( );
FILL FILL_33_3_0 ( );
FILL FILL_33_3_1 ( );
FILL FILL_33_3_2 ( );
FILL FILL_33_4_0 ( );
FILL FILL_33_4_1 ( );
FILL FILL_33_4_2 ( );
FILL FILL_33_5_0 ( );
FILL FILL_33_5_1 ( );
FILL FILL_33_5_2 ( );
FILL FILL_33_6_0 ( );
FILL FILL_33_6_1 ( );
FILL FILL_33_6_2 ( );
FILL FILL_33_7_0 ( );
FILL FILL_33_7_1 ( );
FILL FILL_33_7_2 ( );
FILL FILL_33_8_0 ( );
FILL FILL_33_8_1 ( );
FILL FILL_33_8_2 ( );
FILL FILL_34_1 ( );
FILL FILL_34_2 ( );
FILL FILL_34_3 ( );
FILL FILL_34_0_0 ( );
FILL FILL_34_0_1 ( );
FILL FILL_34_0_2 ( );
FILL FILL_34_1_0 ( );
FILL FILL_34_1_1 ( );
FILL FILL_34_1_2 ( );
FILL FILL_34_2_0 ( );
FILL FILL_34_2_1 ( );
FILL FILL_34_2_2 ( );
FILL FILL_34_3_0 ( );
FILL FILL_34_3_1 ( );
FILL FILL_34_3_2 ( );
FILL FILL_34_4_0 ( );
FILL FILL_34_4_1 ( );
FILL FILL_34_4_2 ( );
FILL FILL_34_5_0 ( );
FILL FILL_34_5_1 ( );
FILL FILL_34_5_2 ( );
FILL FILL_34_6_0 ( );
FILL FILL_34_6_1 ( );
FILL FILL_34_6_2 ( );
FILL FILL_34_7_0 ( );
FILL FILL_34_7_1 ( );
FILL FILL_34_7_2 ( );
FILL FILL_34_8_0 ( );
FILL FILL_34_8_1 ( );
FILL FILL_34_8_2 ( );
FILL FILL_35_1 ( );
FILL FILL_35_2 ( );
FILL FILL_35_0_0 ( );
FILL FILL_35_0_1 ( );
FILL FILL_35_0_2 ( );
FILL FILL_35_1_0 ( );
FILL FILL_35_1_1 ( );
FILL FILL_35_1_2 ( );
FILL FILL_35_2_0 ( );
FILL FILL_35_2_1 ( );
FILL FILL_35_2_2 ( );
FILL FILL_35_3_0 ( );
FILL FILL_35_3_1 ( );
FILL FILL_35_3_2 ( );
FILL FILL_35_4_0 ( );
FILL FILL_35_4_1 ( );
FILL FILL_35_4_2 ( );
FILL FILL_35_5_0 ( );
FILL FILL_35_5_1 ( );
FILL FILL_35_5_2 ( );
FILL FILL_35_6_0 ( );
FILL FILL_35_6_1 ( );
FILL FILL_35_6_2 ( );
FILL FILL_35_7_0 ( );
FILL FILL_35_7_1 ( );
FILL FILL_35_7_2 ( );
FILL FILL_35_8_0 ( );
FILL FILL_35_8_1 ( );
FILL FILL_35_8_2 ( );
FILL FILL_36_1 ( );
FILL FILL_36_2 ( );
FILL FILL_36_0_0 ( );
FILL FILL_36_0_1 ( );
FILL FILL_36_0_2 ( );
FILL FILL_36_1_0 ( );
FILL FILL_36_1_1 ( );
FILL FILL_36_1_2 ( );
FILL FILL_36_2_0 ( );
FILL FILL_36_2_1 ( );
FILL FILL_36_2_2 ( );
FILL FILL_36_3_0 ( );
FILL FILL_36_3_1 ( );
FILL FILL_36_3_2 ( );
FILL FILL_36_4_0 ( );
FILL FILL_36_4_1 ( );
FILL FILL_36_4_2 ( );
FILL FILL_36_5_0 ( );
FILL FILL_36_5_1 ( );
FILL FILL_36_5_2 ( );
FILL FILL_36_6_0 ( );
FILL FILL_36_6_1 ( );
FILL FILL_36_6_2 ( );
FILL FILL_36_7_0 ( );
FILL FILL_36_7_1 ( );
FILL FILL_36_7_2 ( );
FILL FILL_36_8_0 ( );
FILL FILL_36_8_1 ( );
FILL FILL_36_8_2 ( );
FILL FILL_37_1 ( );
FILL FILL_37_2 ( );
FILL FILL_37_0_0 ( );
FILL FILL_37_0_1 ( );
FILL FILL_37_0_2 ( );
FILL FILL_37_1_0 ( );
FILL FILL_37_1_1 ( );
FILL FILL_37_1_2 ( );
FILL FILL_37_2_0 ( );
FILL FILL_37_2_1 ( );
FILL FILL_37_2_2 ( );
FILL FILL_37_3_0 ( );
FILL FILL_37_3_1 ( );
FILL FILL_37_3_2 ( );
FILL FILL_37_4_0 ( );
FILL FILL_37_4_1 ( );
FILL FILL_37_4_2 ( );
FILL FILL_37_5_0 ( );
FILL FILL_37_5_1 ( );
FILL FILL_37_5_2 ( );
FILL FILL_37_6_0 ( );
FILL FILL_37_6_1 ( );
FILL FILL_37_6_2 ( );
FILL FILL_37_7_0 ( );
FILL FILL_37_7_1 ( );
FILL FILL_37_7_2 ( );
FILL FILL_37_8_0 ( );
FILL FILL_37_8_1 ( );
FILL FILL_37_8_2 ( );
FILL FILL_38_0_0 ( );
FILL FILL_38_0_1 ( );
FILL FILL_38_0_2 ( );
FILL FILL_38_1_0 ( );
FILL FILL_38_1_1 ( );
FILL FILL_38_1_2 ( );
FILL FILL_38_2_0 ( );
FILL FILL_38_2_1 ( );
FILL FILL_38_2_2 ( );
FILL FILL_38_3_0 ( );
FILL FILL_38_3_1 ( );
FILL FILL_38_3_2 ( );
FILL FILL_38_4_0 ( );
FILL FILL_38_4_1 ( );
FILL FILL_38_4_2 ( );
FILL FILL_38_5_0 ( );
FILL FILL_38_5_1 ( );
FILL FILL_38_5_2 ( );
FILL FILL_38_6_0 ( );
FILL FILL_38_6_1 ( );
FILL FILL_38_6_2 ( );
FILL FILL_38_7_0 ( );
FILL FILL_38_7_1 ( );
FILL FILL_38_7_2 ( );
FILL FILL_38_8_0 ( );
FILL FILL_38_8_1 ( );
FILL FILL_38_8_2 ( );
FILL FILL_39_1 ( );
FILL FILL_39_2 ( );
FILL FILL_39_3 ( );
FILL FILL_39_0_0 ( );
FILL FILL_39_0_1 ( );
FILL FILL_39_0_2 ( );
FILL FILL_39_1_0 ( );
FILL FILL_39_1_1 ( );
FILL FILL_39_1_2 ( );
FILL FILL_39_2_0 ( );
FILL FILL_39_2_1 ( );
FILL FILL_39_2_2 ( );
FILL FILL_39_3_0 ( );
FILL FILL_39_3_1 ( );
FILL FILL_39_3_2 ( );
FILL FILL_39_4_0 ( );
FILL FILL_39_4_1 ( );
FILL FILL_39_4_2 ( );
FILL FILL_39_5_0 ( );
FILL FILL_39_5_1 ( );
FILL FILL_39_5_2 ( );
FILL FILL_39_6_0 ( );
FILL FILL_39_6_1 ( );
FILL FILL_39_6_2 ( );
FILL FILL_39_7_0 ( );
FILL FILL_39_7_1 ( );
FILL FILL_39_7_2 ( );
FILL FILL_39_8_0 ( );
FILL FILL_39_8_1 ( );
FILL FILL_39_8_2 ( );
FILL FILL_40_1 ( );
FILL FILL_40_2 ( );
FILL FILL_40_3 ( );
FILL FILL_40_0_0 ( );
FILL FILL_40_0_1 ( );
FILL FILL_40_0_2 ( );
FILL FILL_40_1_0 ( );
FILL FILL_40_1_1 ( );
FILL FILL_40_1_2 ( );
FILL FILL_40_2_0 ( );
FILL FILL_40_2_1 ( );
FILL FILL_40_2_2 ( );
FILL FILL_40_3_0 ( );
FILL FILL_40_3_1 ( );
FILL FILL_40_3_2 ( );
FILL FILL_40_4_0 ( );
FILL FILL_40_4_1 ( );
FILL FILL_40_4_2 ( );
FILL FILL_40_5_0 ( );
FILL FILL_40_5_1 ( );
FILL FILL_40_5_2 ( );
FILL FILL_40_6_0 ( );
FILL FILL_40_6_1 ( );
FILL FILL_40_6_2 ( );
FILL FILL_40_7_0 ( );
FILL FILL_40_7_1 ( );
FILL FILL_40_7_2 ( );
FILL FILL_40_8_0 ( );
FILL FILL_40_8_1 ( );
FILL FILL_40_8_2 ( );
FILL FILL_41_0_0 ( );
FILL FILL_41_0_1 ( );
FILL FILL_41_0_2 ( );
FILL FILL_41_1_0 ( );
FILL FILL_41_1_1 ( );
FILL FILL_41_1_2 ( );
FILL FILL_41_2_0 ( );
FILL FILL_41_2_1 ( );
FILL FILL_41_2_2 ( );
FILL FILL_41_3_0 ( );
FILL FILL_41_3_1 ( );
FILL FILL_41_3_2 ( );
FILL FILL_41_4_0 ( );
FILL FILL_41_4_1 ( );
FILL FILL_41_4_2 ( );
FILL FILL_41_5_0 ( );
FILL FILL_41_5_1 ( );
FILL FILL_41_5_2 ( );
FILL FILL_41_6_0 ( );
FILL FILL_41_6_1 ( );
FILL FILL_41_6_2 ( );
FILL FILL_41_7_0 ( );
FILL FILL_41_7_1 ( );
FILL FILL_41_7_2 ( );
FILL FILL_41_8_0 ( );
FILL FILL_41_8_1 ( );
FILL FILL_41_8_2 ( );
FILL FILL_42_1 ( );
FILL FILL_42_2 ( );
FILL FILL_42_0_0 ( );
FILL FILL_42_0_1 ( );
FILL FILL_42_0_2 ( );
FILL FILL_42_1_0 ( );
FILL FILL_42_1_1 ( );
FILL FILL_42_1_2 ( );
FILL FILL_42_2_0 ( );
FILL FILL_42_2_1 ( );
FILL FILL_42_2_2 ( );
FILL FILL_42_3_0 ( );
FILL FILL_42_3_1 ( );
FILL FILL_42_3_2 ( );
FILL FILL_42_4_0 ( );
FILL FILL_42_4_1 ( );
FILL FILL_42_4_2 ( );
FILL FILL_42_5_0 ( );
FILL FILL_42_5_1 ( );
FILL FILL_42_5_2 ( );
FILL FILL_42_6_0 ( );
FILL FILL_42_6_1 ( );
FILL FILL_42_6_2 ( );
FILL FILL_42_7_0 ( );
FILL FILL_42_7_1 ( );
FILL FILL_42_7_2 ( );
FILL FILL_42_8_0 ( );
FILL FILL_42_8_1 ( );
FILL FILL_42_8_2 ( );
FILL FILL_43_1 ( );
FILL FILL_43_0_0 ( );
FILL FILL_43_0_1 ( );
FILL FILL_43_0_2 ( );
FILL FILL_43_1_0 ( );
FILL FILL_43_1_1 ( );
FILL FILL_43_1_2 ( );
FILL FILL_43_2_0 ( );
FILL FILL_43_2_1 ( );
FILL FILL_43_2_2 ( );
FILL FILL_43_3_0 ( );
FILL FILL_43_3_1 ( );
FILL FILL_43_3_2 ( );
FILL FILL_43_4_0 ( );
FILL FILL_43_4_1 ( );
FILL FILL_43_4_2 ( );
FILL FILL_43_5_0 ( );
FILL FILL_43_5_1 ( );
FILL FILL_43_5_2 ( );
FILL FILL_43_6_0 ( );
FILL FILL_43_6_1 ( );
FILL FILL_43_6_2 ( );
FILL FILL_43_7_0 ( );
FILL FILL_43_7_1 ( );
FILL FILL_43_7_2 ( );
FILL FILL_43_8_0 ( );
FILL FILL_43_8_1 ( );
FILL FILL_43_8_2 ( );
FILL FILL_44_1 ( );
FILL FILL_44_2 ( );
FILL FILL_44_3 ( );
FILL FILL_44_0_0 ( );
FILL FILL_44_0_1 ( );
FILL FILL_44_0_2 ( );
FILL FILL_44_1_0 ( );
FILL FILL_44_1_1 ( );
FILL FILL_44_1_2 ( );
FILL FILL_44_2_0 ( );
FILL FILL_44_2_1 ( );
FILL FILL_44_2_2 ( );
FILL FILL_44_3_0 ( );
FILL FILL_44_3_1 ( );
FILL FILL_44_3_2 ( );
FILL FILL_44_4_0 ( );
FILL FILL_44_4_1 ( );
FILL FILL_44_4_2 ( );
FILL FILL_44_5_0 ( );
FILL FILL_44_5_1 ( );
FILL FILL_44_5_2 ( );
FILL FILL_44_6_0 ( );
FILL FILL_44_6_1 ( );
FILL FILL_44_6_2 ( );
FILL FILL_44_7_0 ( );
FILL FILL_44_7_1 ( );
FILL FILL_44_7_2 ( );
FILL FILL_44_8_0 ( );
FILL FILL_44_8_1 ( );
FILL FILL_44_8_2 ( );
FILL FILL_45_0_0 ( );
FILL FILL_45_0_1 ( );
FILL FILL_45_0_2 ( );
FILL FILL_45_1_0 ( );
FILL FILL_45_1_1 ( );
FILL FILL_45_1_2 ( );
FILL FILL_45_2_0 ( );
FILL FILL_45_2_1 ( );
FILL FILL_45_2_2 ( );
FILL FILL_45_3_0 ( );
FILL FILL_45_3_1 ( );
FILL FILL_45_3_2 ( );
FILL FILL_45_4_0 ( );
FILL FILL_45_4_1 ( );
FILL FILL_45_4_2 ( );
FILL FILL_45_5_0 ( );
FILL FILL_45_5_1 ( );
FILL FILL_45_5_2 ( );
FILL FILL_45_6_0 ( );
FILL FILL_45_6_1 ( );
FILL FILL_45_6_2 ( );
FILL FILL_45_7_0 ( );
FILL FILL_45_7_1 ( );
FILL FILL_45_7_2 ( );
FILL FILL_45_8_0 ( );
FILL FILL_45_8_1 ( );
FILL FILL_45_8_2 ( );
FILL FILL_46_1 ( );
FILL FILL_46_0_0 ( );
FILL FILL_46_0_1 ( );
FILL FILL_46_0_2 ( );
FILL FILL_46_1_0 ( );
FILL FILL_46_1_1 ( );
FILL FILL_46_1_2 ( );
FILL FILL_46_2_0 ( );
FILL FILL_46_2_1 ( );
FILL FILL_46_2_2 ( );
FILL FILL_46_3_0 ( );
FILL FILL_46_3_1 ( );
FILL FILL_46_3_2 ( );
FILL FILL_46_4_0 ( );
FILL FILL_46_4_1 ( );
FILL FILL_46_4_2 ( );
FILL FILL_46_5_0 ( );
FILL FILL_46_5_1 ( );
FILL FILL_46_5_2 ( );
FILL FILL_46_6_0 ( );
FILL FILL_46_6_1 ( );
FILL FILL_46_6_2 ( );
FILL FILL_46_7_0 ( );
FILL FILL_46_7_1 ( );
FILL FILL_46_7_2 ( );
FILL FILL_46_8_0 ( );
FILL FILL_46_8_1 ( );
FILL FILL_46_8_2 ( );
FILL FILL_47_1 ( );
FILL FILL_47_0_0 ( );
FILL FILL_47_0_1 ( );
FILL FILL_47_0_2 ( );
FILL FILL_47_1_0 ( );
FILL FILL_47_1_1 ( );
FILL FILL_47_1_2 ( );
FILL FILL_47_2_0 ( );
FILL FILL_47_2_1 ( );
FILL FILL_47_2_2 ( );
FILL FILL_47_3_0 ( );
FILL FILL_47_3_1 ( );
FILL FILL_47_3_2 ( );
FILL FILL_47_4_0 ( );
FILL FILL_47_4_1 ( );
FILL FILL_47_4_2 ( );
FILL FILL_47_5_0 ( );
FILL FILL_47_5_1 ( );
FILL FILL_47_5_2 ( );
FILL FILL_47_6_0 ( );
FILL FILL_47_6_1 ( );
FILL FILL_47_6_2 ( );
FILL FILL_47_7_0 ( );
FILL FILL_47_7_1 ( );
FILL FILL_47_7_2 ( );
FILL FILL_47_8_0 ( );
FILL FILL_47_8_1 ( );
FILL FILL_47_8_2 ( );
FILL FILL_48_1 ( );
FILL FILL_48_2 ( );
FILL FILL_48_3 ( );
FILL FILL_48_0_0 ( );
FILL FILL_48_0_1 ( );
FILL FILL_48_0_2 ( );
FILL FILL_48_1_0 ( );
FILL FILL_48_1_1 ( );
FILL FILL_48_1_2 ( );
FILL FILL_48_2_0 ( );
FILL FILL_48_2_1 ( );
FILL FILL_48_2_2 ( );
FILL FILL_48_3_0 ( );
FILL FILL_48_3_1 ( );
FILL FILL_48_3_2 ( );
FILL FILL_48_4_0 ( );
FILL FILL_48_4_1 ( );
FILL FILL_48_4_2 ( );
FILL FILL_48_5_0 ( );
FILL FILL_48_5_1 ( );
FILL FILL_48_5_2 ( );
FILL FILL_48_6_0 ( );
FILL FILL_48_6_1 ( );
FILL FILL_48_6_2 ( );
FILL FILL_48_7_0 ( );
FILL FILL_48_7_1 ( );
FILL FILL_48_7_2 ( );
FILL FILL_48_8_0 ( );
FILL FILL_48_8_1 ( );
FILL FILL_48_8_2 ( );
FILL FILL_49_0_0 ( );
FILL FILL_49_0_1 ( );
FILL FILL_49_0_2 ( );
FILL FILL_49_1_0 ( );
FILL FILL_49_1_1 ( );
FILL FILL_49_1_2 ( );
FILL FILL_49_2_0 ( );
FILL FILL_49_2_1 ( );
FILL FILL_49_2_2 ( );
FILL FILL_49_3_0 ( );
FILL FILL_49_3_1 ( );
FILL FILL_49_3_2 ( );
FILL FILL_49_4_0 ( );
FILL FILL_49_4_1 ( );
FILL FILL_49_4_2 ( );
FILL FILL_49_5_0 ( );
FILL FILL_49_5_1 ( );
FILL FILL_49_5_2 ( );
FILL FILL_49_6_0 ( );
FILL FILL_49_6_1 ( );
FILL FILL_49_6_2 ( );
FILL FILL_49_7_0 ( );
FILL FILL_49_7_1 ( );
FILL FILL_49_7_2 ( );
FILL FILL_49_8_0 ( );
FILL FILL_49_8_1 ( );
FILL FILL_49_8_2 ( );
FILL FILL_50_0_0 ( );
FILL FILL_50_0_1 ( );
FILL FILL_50_0_2 ( );
FILL FILL_50_1_0 ( );
FILL FILL_50_1_1 ( );
FILL FILL_50_1_2 ( );
FILL FILL_50_2_0 ( );
FILL FILL_50_2_1 ( );
FILL FILL_50_2_2 ( );
FILL FILL_50_3_0 ( );
FILL FILL_50_3_1 ( );
FILL FILL_50_3_2 ( );
FILL FILL_50_4_0 ( );
FILL FILL_50_4_1 ( );
FILL FILL_50_4_2 ( );
FILL FILL_50_5_0 ( );
FILL FILL_50_5_1 ( );
FILL FILL_50_5_2 ( );
FILL FILL_50_6_0 ( );
FILL FILL_50_6_1 ( );
FILL FILL_50_6_2 ( );
FILL FILL_50_7_0 ( );
FILL FILL_50_7_1 ( );
FILL FILL_50_7_2 ( );
FILL FILL_50_8_0 ( );
FILL FILL_50_8_1 ( );
FILL FILL_50_8_2 ( );
FILL FILL_51_0_0 ( );
FILL FILL_51_0_1 ( );
FILL FILL_51_0_2 ( );
FILL FILL_51_1_0 ( );
FILL FILL_51_1_1 ( );
FILL FILL_51_1_2 ( );
FILL FILL_51_2_0 ( );
FILL FILL_51_2_1 ( );
FILL FILL_51_2_2 ( );
FILL FILL_51_3_0 ( );
FILL FILL_51_3_1 ( );
FILL FILL_51_3_2 ( );
FILL FILL_51_4_0 ( );
FILL FILL_51_4_1 ( );
FILL FILL_51_4_2 ( );
FILL FILL_51_5_0 ( );
FILL FILL_51_5_1 ( );
FILL FILL_51_5_2 ( );
FILL FILL_51_6_0 ( );
FILL FILL_51_6_1 ( );
FILL FILL_51_6_2 ( );
FILL FILL_51_7_0 ( );
FILL FILL_51_7_1 ( );
FILL FILL_51_7_2 ( );
FILL FILL_51_8_0 ( );
FILL FILL_51_8_1 ( );
FILL FILL_51_8_2 ( );
FILL FILL_52_1 ( );
FILL FILL_52_0_0 ( );
FILL FILL_52_0_1 ( );
FILL FILL_52_0_2 ( );
FILL FILL_52_1_0 ( );
FILL FILL_52_1_1 ( );
FILL FILL_52_1_2 ( );
FILL FILL_52_2_0 ( );
FILL FILL_52_2_1 ( );
FILL FILL_52_2_2 ( );
FILL FILL_52_3_0 ( );
FILL FILL_52_3_1 ( );
FILL FILL_52_3_2 ( );
FILL FILL_52_4_0 ( );
FILL FILL_52_4_1 ( );
FILL FILL_52_4_2 ( );
FILL FILL_52_5_0 ( );
FILL FILL_52_5_1 ( );
FILL FILL_52_5_2 ( );
FILL FILL_52_6_0 ( );
FILL FILL_52_6_1 ( );
FILL FILL_52_6_2 ( );
FILL FILL_52_7_0 ( );
FILL FILL_52_7_1 ( );
FILL FILL_52_7_2 ( );
FILL FILL_52_8_0 ( );
FILL FILL_52_8_1 ( );
FILL FILL_52_8_2 ( );
FILL FILL_53_1 ( );
FILL FILL_53_2 ( );
FILL FILL_53_0_0 ( );
FILL FILL_53_0_1 ( );
FILL FILL_53_0_2 ( );
FILL FILL_53_1_0 ( );
FILL FILL_53_1_1 ( );
FILL FILL_53_1_2 ( );
FILL FILL_53_2_0 ( );
FILL FILL_53_2_1 ( );
FILL FILL_53_2_2 ( );
FILL FILL_53_3_0 ( );
FILL FILL_53_3_1 ( );
FILL FILL_53_3_2 ( );
FILL FILL_53_4_0 ( );
FILL FILL_53_4_1 ( );
FILL FILL_53_4_2 ( );
FILL FILL_53_5_0 ( );
FILL FILL_53_5_1 ( );
FILL FILL_53_5_2 ( );
FILL FILL_53_6_0 ( );
FILL FILL_53_6_1 ( );
FILL FILL_53_6_2 ( );
FILL FILL_53_7_0 ( );
FILL FILL_53_7_1 ( );
FILL FILL_53_7_2 ( );
FILL FILL_53_8_0 ( );
FILL FILL_53_8_1 ( );
FILL FILL_53_8_2 ( );
FILL FILL_54_1 ( );
FILL FILL_54_2 ( );
FILL FILL_54_3 ( );
endmodule
