VERSION 5.3 ;
   NAMESCASESENSITIVE ON ;
   NOWIREEXTENSIONATPIN ON ;
   DIVIDERCHAR "/" ;
   BUSBITCHARS "[]" ;
UNITS
   DATABASE MICRONS 1000 ;
END UNITS

MACRO FIR
   CLASS BLOCK ;
   FOREIGN FIR ;
   ORIGIN -1.2000 3.4500 ;
   SIZE 1571.5500 BY 1479.9000 ;
   PIN clk
      PORT
         LAYER metal1 ;
	    RECT 762.6000 1395.4501 763.8000 1395.6000 ;
	    RECT 793.8000 1395.4501 795.0000 1395.6000 ;
	    RECT 762.6000 1394.5500 795.0000 1395.4501 ;
	    RECT 762.6000 1394.4000 763.8000 1394.5500 ;
	    RECT 793.8000 1394.4000 795.0000 1394.5500 ;
	    RECT 762.6000 1301.4000 763.8000 1302.6000 ;
	    RECT 1108.2001 1100.4000 1109.4000 1101.6000 ;
	    RECT 606.6000 1041.4501 607.8000 1041.6000 ;
	    RECT 630.6000 1041.4501 631.8000 1041.6000 ;
	    RECT 606.6000 1040.5500 631.8000 1041.4501 ;
	    RECT 606.6000 1040.4000 607.8000 1040.5500 ;
	    RECT 630.6000 1040.4000 631.8000 1040.5500 ;
	    RECT 1041.0000 1041.4501 1042.2001 1041.6000 ;
	    RECT 1091.4000 1041.4501 1092.6000 1041.6000 ;
	    RECT 1041.0000 1040.5500 1092.6000 1041.4501 ;
	    RECT 1041.0000 1040.4000 1042.2001 1040.5500 ;
	    RECT 1091.4000 1040.4000 1092.6000 1040.5500 ;
	    RECT 630.6000 756.4500 631.8000 756.6000 ;
	    RECT 649.8000 756.4500 651.0000 756.6000 ;
	    RECT 630.6000 755.5500 651.0000 756.4500 ;
	    RECT 630.6000 755.4000 631.8000 755.5500 ;
	    RECT 649.8000 755.4000 651.0000 755.5500 ;
	    RECT 625.8000 522.4500 627.0000 522.6000 ;
	    RECT 630.6000 522.4500 631.8000 522.6000 ;
	    RECT 625.8000 521.5500 631.8000 522.4500 ;
	    RECT 625.8000 521.4000 627.0000 521.5500 ;
	    RECT 630.6000 521.4000 631.8000 521.5500 ;
	    RECT 1009.8000 380.4000 1011.0000 381.6000 ;
	    RECT 472.2000 281.4000 473.4000 282.6000 ;
	    RECT 801.0000 282.4500 802.2000 282.6000 ;
	    RECT 815.4000 282.4500 816.6000 282.6000 ;
	    RECT 825.0000 282.4500 826.2000 282.6000 ;
	    RECT 801.0000 281.5500 826.2000 282.4500 ;
	    RECT 801.0000 281.4000 802.2000 281.5500 ;
	    RECT 815.4000 281.4000 816.6000 281.5500 ;
	    RECT 825.0000 281.4000 826.2000 281.5500 ;
         LAYER metal2 ;
	    RECT 793.9500 1395.6000 794.8500 1476.4501 ;
	    RECT 762.6000 1394.4000 763.8000 1395.6000 ;
	    RECT 793.8000 1394.4000 795.0000 1395.6000 ;
	    RECT 762.7500 1302.6000 763.6500 1394.4000 ;
	    RECT 762.6000 1301.4000 763.8000 1302.6000 ;
	    RECT 762.7500 1212.6000 763.6500 1301.4000 ;
	    RECT 630.6000 1211.4000 631.8000 1212.6000 ;
	    RECT 762.6000 1211.4000 763.8000 1212.6000 ;
	    RECT 810.6000 1211.4000 811.8000 1212.6000 ;
	    RECT 630.7500 1041.6000 631.6500 1211.4000 ;
	    RECT 810.7500 1044.6000 811.6500 1211.4000 ;
	    RECT 1108.2001 1100.4000 1109.4000 1101.6000 ;
	    RECT 1108.3500 1050.6000 1109.2500 1100.4000 ;
	    RECT 1091.4000 1049.4000 1092.6000 1050.6000 ;
	    RECT 1108.2001 1049.4000 1109.4000 1050.6000 ;
	    RECT 810.6000 1043.4000 811.8000 1044.6000 ;
	    RECT 1041.0000 1043.4000 1042.2001 1044.6000 ;
	    RECT 1041.1500 1041.6000 1042.0500 1043.4000 ;
	    RECT 1091.5500 1041.6000 1092.4501 1049.4000 ;
	    RECT 630.6000 1040.4000 631.8000 1041.6000 ;
	    RECT 1041.0000 1040.4000 1042.2001 1041.6000 ;
	    RECT 1091.4000 1040.4000 1092.6000 1041.6000 ;
	    RECT 630.7500 1032.6000 631.6500 1040.4000 ;
	    RECT 630.6000 1031.4000 631.8000 1032.6000 ;
	    RECT 649.8000 1031.4000 651.0000 1032.6000 ;
	    RECT 649.9500 756.6000 650.8500 1031.4000 ;
	    RECT 630.6000 755.4000 631.8000 756.6000 ;
	    RECT 649.8000 755.4000 651.0000 756.6000 ;
	    RECT 630.7500 684.6000 631.6500 755.4000 ;
	    RECT 625.8000 683.4000 627.0000 684.6000 ;
	    RECT 630.6000 683.4000 631.8000 684.6000 ;
	    RECT 625.9500 522.6000 626.8500 683.4000 ;
	    RECT 625.8000 521.4000 627.0000 522.6000 ;
	    RECT 625.9500 516.6000 626.8500 521.4000 ;
	    RECT 472.2000 515.4000 473.4000 516.6000 ;
	    RECT 625.8000 515.4000 627.0000 516.6000 ;
	    RECT 472.3500 312.6000 473.2500 515.4000 ;
	    RECT 1009.8000 380.4000 1011.0000 381.6000 ;
	    RECT 1009.9500 372.6000 1010.8500 380.4000 ;
	    RECT 815.4000 371.4000 816.6000 372.6000 ;
	    RECT 1009.8000 371.4000 1011.0000 372.6000 ;
	    RECT 472.2000 311.4000 473.4000 312.6000 ;
	    RECT 801.0000 311.4000 802.2000 312.6000 ;
	    RECT 472.3500 282.6000 473.2500 311.4000 ;
	    RECT 801.1500 282.6000 802.0500 311.4000 ;
	    RECT 815.5500 282.6000 816.4500 371.4000 ;
	    RECT 472.2000 281.4000 473.4000 282.6000 ;
	    RECT 801.0000 281.4000 802.2000 282.6000 ;
	    RECT 815.4000 281.4000 816.6000 282.6000 ;
         LAYER metal3 ;
	    RECT 630.3000 1212.7500 632.1000 1212.9000 ;
	    RECT 762.3000 1212.7500 764.1000 1212.9000 ;
	    RECT 810.3000 1212.7500 812.1000 1212.9000 ;
	    RECT 630.3000 1211.2500 812.1000 1212.7500 ;
	    RECT 630.3000 1211.1000 632.1000 1211.2500 ;
	    RECT 762.3000 1211.1000 764.1000 1211.2500 ;
	    RECT 810.3000 1211.1000 812.1000 1211.2500 ;
	    RECT 1091.1000 1050.7500 1092.9000 1050.9000 ;
	    RECT 1107.9000 1050.7500 1109.7001 1050.9000 ;
	    RECT 1091.1000 1049.2500 1109.7001 1050.7500 ;
	    RECT 1091.1000 1049.1000 1092.9000 1049.2500 ;
	    RECT 1107.9000 1049.1000 1109.7001 1049.2500 ;
	    RECT 810.3000 1044.7500 812.1000 1044.9000 ;
	    RECT 1040.7001 1044.7500 1042.5000 1044.9000 ;
	    RECT 810.3000 1043.2500 1042.5000 1044.7500 ;
	    RECT 810.3000 1043.1000 812.1000 1043.2500 ;
	    RECT 1040.7001 1043.1000 1042.5000 1043.2500 ;
	    RECT 630.3000 1032.7500 632.1000 1032.9000 ;
	    RECT 649.5000 1032.7500 651.3000 1032.9000 ;
	    RECT 630.3000 1031.2500 651.3000 1032.7500 ;
	    RECT 630.3000 1031.1000 632.1000 1031.2500 ;
	    RECT 649.5000 1031.1000 651.3000 1031.2500 ;
	    RECT 625.5000 684.7500 627.3000 684.9000 ;
	    RECT 630.3000 684.7500 632.1000 684.9000 ;
	    RECT 625.5000 683.2500 632.1000 684.7500 ;
	    RECT 625.5000 683.1000 627.3000 683.2500 ;
	    RECT 630.3000 683.1000 632.1000 683.2500 ;
	    RECT 471.9000 516.7500 473.7000 516.9000 ;
	    RECT 625.5000 516.7500 627.3000 516.9000 ;
	    RECT 471.9000 515.2500 627.3000 516.7500 ;
	    RECT 471.9000 515.1000 473.7000 515.2500 ;
	    RECT 625.5000 515.1000 627.3000 515.2500 ;
	    RECT 815.1000 372.7500 816.9000 372.9000 ;
	    RECT 1009.5000 372.7500 1011.3000 372.9000 ;
	    RECT 815.1000 371.2500 1011.3000 372.7500 ;
	    RECT 815.1000 371.1000 816.9000 371.2500 ;
	    RECT 1009.5000 371.1000 1011.3000 371.2500 ;
	    RECT 471.9000 312.7500 473.7000 312.9000 ;
	    RECT 800.7000 312.7500 802.5000 312.9000 ;
	    RECT 471.9000 311.2500 802.5000 312.7500 ;
	    RECT 471.9000 311.1000 473.7000 311.2500 ;
	    RECT 800.7000 311.1000 802.5000 311.2500 ;
      END
   END clk
   PIN rst
      PORT
         LAYER metal1 ;
	    RECT 462.6000 704.4000 463.8000 705.6000 ;
	    RECT 462.6000 651.4500 463.8000 651.6000 ;
	    RECT 469.8000 651.4500 471.0000 651.6000 ;
	    RECT 462.6000 650.5500 471.0000 651.4500 ;
	    RECT 462.6000 650.4000 463.8000 650.5500 ;
	    RECT 469.8000 650.4000 471.0000 650.5500 ;
	    RECT 544.2000 497.4000 545.4000 498.6000 ;
	    RECT 597.0000 497.4000 598.2000 498.6000 ;
	    RECT 465.0000 438.4500 466.2000 438.6000 ;
	    RECT 469.8000 438.4500 471.0000 438.6000 ;
	    RECT 465.0000 437.5500 471.0000 438.4500 ;
	    RECT 465.0000 437.4000 466.2000 437.5500 ;
	    RECT 469.8000 437.4000 471.0000 437.5500 ;
	    RECT 503.4000 317.4000 504.6000 318.6000 ;
	    RECT 630.6000 164.4000 631.8000 165.6000 ;
         LAYER metal2 ;
	    RECT 462.6000 704.4000 463.8000 705.6000 ;
	    RECT 462.7500 651.6000 463.6500 704.4000 ;
	    RECT 462.6000 650.4000 463.8000 651.6000 ;
	    RECT 469.8000 650.4000 471.0000 651.6000 ;
	    RECT 469.9500 486.6000 470.8500 650.4000 ;
	    RECT 544.2000 497.4000 545.4000 498.6000 ;
	    RECT 597.0000 497.4000 598.2000 498.6000 ;
	    RECT 544.3500 486.6000 545.2500 497.4000 ;
	    RECT 597.1500 486.6000 598.0500 497.4000 ;
	    RECT 465.0000 485.4000 466.2000 486.6000 ;
	    RECT 469.8000 485.4000 471.0000 486.6000 ;
	    RECT 544.2000 485.4000 545.4000 486.6000 ;
	    RECT 597.0000 485.4000 598.2000 486.6000 ;
	    RECT 465.1500 438.6000 466.0500 485.4000 ;
	    RECT 465.0000 437.4000 466.2000 438.6000 ;
	    RECT 465.1500 360.6000 466.0500 437.4000 ;
	    RECT 465.0000 359.4000 466.2000 360.6000 ;
	    RECT 503.4000 359.4000 504.6000 360.6000 ;
	    RECT 503.5500 318.6000 504.4500 359.4000 ;
	    RECT 503.4000 317.4000 504.6000 318.6000 ;
	    RECT 503.5500 180.6000 504.4500 317.4000 ;
	    RECT 503.4000 179.4000 504.6000 180.6000 ;
	    RECT 592.2000 179.4000 593.4000 180.6000 ;
	    RECT 630.6000 179.4000 631.8000 180.6000 ;
	    RECT 592.3500 -3.4500 593.2500 179.4000 ;
	    RECT 630.7500 165.6000 631.6500 179.4000 ;
	    RECT 630.6000 164.4000 631.8000 165.6000 ;
         LAYER metal3 ;
	    RECT 464.7000 486.7500 466.5000 486.9000 ;
	    RECT 469.5000 486.7500 471.3000 486.9000 ;
	    RECT 543.9000 486.7500 545.7000 486.9000 ;
	    RECT 596.7000 486.7500 598.5000 486.9000 ;
	    RECT 464.7000 485.2500 598.5000 486.7500 ;
	    RECT 464.7000 485.1000 466.5000 485.2500 ;
	    RECT 469.5000 485.1000 471.3000 485.2500 ;
	    RECT 543.9000 485.1000 545.7000 485.2500 ;
	    RECT 596.7000 485.1000 598.5000 485.2500 ;
	    RECT 464.7000 360.7500 466.5000 360.9000 ;
	    RECT 503.1000 360.7500 504.9000 360.9000 ;
	    RECT 464.7000 359.2500 504.9000 360.7500 ;
	    RECT 464.7000 359.1000 466.5000 359.2500 ;
	    RECT 503.1000 359.1000 504.9000 359.2500 ;
	    RECT 503.1000 180.7500 504.9000 180.9000 ;
	    RECT 591.9000 180.7500 593.7000 180.9000 ;
	    RECT 630.3000 180.7500 632.1000 180.9000 ;
	    RECT 503.1000 179.2500 632.1000 180.7500 ;
	    RECT 503.1000 179.1000 504.9000 179.2500 ;
	    RECT 591.9000 179.1000 593.7000 179.2500 ;
	    RECT 630.3000 179.1000 632.1000 179.2500 ;
      END
   END rst
   PIN din[0]
      PORT
         LAYER metal1 ;
	    RECT 1554.6000 1242.4501 1555.8000 1242.6000 ;
	    RECT 1566.6000 1242.4501 1567.8000 1242.6000 ;
	    RECT 1554.6000 1241.5500 1567.8000 1242.4501 ;
	    RECT 1554.6000 1241.4000 1555.8000 1241.5500 ;
	    RECT 1566.6000 1241.4000 1567.8000 1241.5500 ;
         LAYER metal2 ;
	    RECT 1566.6000 1241.4000 1567.8000 1242.6000 ;
         LAYER metal3 ;
	    RECT 1566.3000 1242.7500 1568.1000 1242.9000 ;
	    RECT 1571.2500 1242.7500 1572.7500 1245.7500 ;
	    RECT 1566.3000 1241.2500 1572.7500 1242.7500 ;
	    RECT 1566.3000 1241.1000 1568.1000 1241.2500 ;
      END
   END din[0]
   PIN din[1]
      PORT
         LAYER metal1 ;
	    RECT 1564.2001 915.4500 1565.4000 915.6000 ;
	    RECT 1566.6000 915.4500 1567.8000 915.6000 ;
	    RECT 1564.2001 914.5500 1567.8000 915.4500 ;
	    RECT 1564.2001 914.4000 1565.4000 914.5500 ;
	    RECT 1566.6000 914.4000 1567.8000 914.5500 ;
         LAYER metal2 ;
	    RECT 1566.6000 914.4000 1567.8000 915.6000 ;
	    RECT 1566.7500 912.6000 1567.6500 914.4000 ;
	    RECT 1566.6000 911.4000 1567.8000 912.6000 ;
         LAYER metal3 ;
	    RECT 1566.3000 912.7500 1568.1000 912.9000 ;
	    RECT 1571.2500 912.7500 1572.7500 915.7500 ;
	    RECT 1566.3000 911.2500 1572.7500 912.7500 ;
	    RECT 1566.3000 911.1000 1568.1000 911.2500 ;
      END
   END din[1]
   PIN din[2]
      PORT
         LAYER metal1 ;
	    RECT 1151.4000 1454.4000 1152.6000 1455.6000 ;
         LAYER metal2 ;
	    RECT 1149.1500 1475.5500 1152.4501 1476.4501 ;
	    RECT 1151.5500 1455.6000 1152.4501 1475.5500 ;
	    RECT 1151.4000 1454.4000 1152.6000 1455.6000 ;
      END
   END din[2]
   PIN din[3]
      PORT
         LAYER metal1 ;
	    RECT 1319.4000 1454.4000 1320.6000 1455.6000 ;
         LAYER metal2 ;
	    RECT 1317.1500 1475.5500 1320.4501 1476.4501 ;
	    RECT 1319.5500 1455.6000 1320.4501 1475.5500 ;
	    RECT 1319.4000 1454.4000 1320.6000 1455.6000 ;
      END
   END din[3]
   PIN din[4]
      PORT
         LAYER metal1 ;
	    RECT 1547.4000 1128.4501 1548.6000 1128.6000 ;
	    RECT 1566.6000 1128.4501 1567.8000 1128.6000 ;
	    RECT 1547.4000 1127.5500 1567.8000 1128.4501 ;
	    RECT 1547.4000 1127.4000 1548.6000 1127.5500 ;
	    RECT 1566.6000 1127.4000 1567.8000 1127.5500 ;
         LAYER metal2 ;
	    RECT 1566.6000 1127.4000 1567.8000 1128.6000 ;
         LAYER metal3 ;
	    RECT 1566.3000 1128.7500 1568.1000 1128.9000 ;
	    RECT 1566.3000 1127.2500 1572.7500 1128.7500 ;
	    RECT 1566.3000 1127.1000 1568.1000 1127.2500 ;
	    RECT 1571.2500 1124.2500 1572.7500 1127.2500 ;
      END
   END din[4]
   PIN din[5]
      PORT
         LAYER metal1 ;
	    RECT 525.0000 48.4500 526.2000 48.6000 ;
	    RECT 532.2000 48.4500 533.4000 48.6000 ;
	    RECT 525.0000 47.5500 533.4000 48.4500 ;
	    RECT 525.0000 47.4000 526.2000 47.5500 ;
	    RECT 532.2000 47.4000 533.4000 47.5500 ;
         LAYER metal2 ;
	    RECT 532.2000 47.4000 533.4000 48.6000 ;
	    RECT 532.3500 6.6000 533.2500 47.4000 ;
	    RECT 522.6000 5.4000 523.8000 6.6000 ;
	    RECT 532.2000 5.4000 533.4000 6.6000 ;
	    RECT 522.7500 -3.4500 523.6500 5.4000 ;
         LAYER metal3 ;
	    RECT 522.3000 6.7500 524.1000 6.9000 ;
	    RECT 531.9000 6.7500 533.7000 6.9000 ;
	    RECT 522.3000 5.2500 533.7000 6.7500 ;
	    RECT 522.3000 5.1000 524.1000 5.2500 ;
	    RECT 531.9000 5.1000 533.7000 5.2500 ;
      END
   END din[5]
   PIN din[6]
      PORT
         LAYER metal1 ;
	    RECT 1566.6000 707.4000 1567.8000 708.6000 ;
         LAYER metal2 ;
	    RECT 1566.6000 707.4000 1567.8000 708.6000 ;
         LAYER metal3 ;
	    RECT 1566.3000 708.7500 1568.1000 708.9000 ;
	    RECT 1566.3000 707.2500 1572.7500 708.7500 ;
	    RECT 1566.3000 707.1000 1568.1000 707.2500 ;
	    RECT 1571.2500 704.2500 1572.7500 707.2500 ;
      END
   END din[6]
   PIN din[7]
      PORT
         LAYER metal1 ;
	    RECT 844.2000 14.4000 845.4000 15.6000 ;
         LAYER metal2 ;
	    RECT 844.2000 14.4000 845.4000 15.6000 ;
	    RECT 844.3500 -2.5500 845.2500 14.4000 ;
	    RECT 841.9500 -3.4500 845.2500 -2.5500 ;
      END
   END din[7]
   PIN dout[0]
      PORT
         LAYER metal1 ;
	    RECT 1290.6000 1460.4000 1291.8000 1461.6000 ;
         LAYER metal2 ;
	    RECT 1290.7500 1475.5500 1294.0500 1476.4501 ;
	    RECT 1290.7500 1461.6000 1291.6500 1475.5500 ;
	    RECT 1290.6000 1460.4000 1291.8000 1461.6000 ;
      END
   END dout[0]
   PIN dout[1]
      PORT
         LAYER metal1 ;
	    RECT 1537.8000 41.4000 1539.0000 42.6000 ;
         LAYER metal2 ;
	    RECT 1537.8000 41.4000 1539.0000 42.6000 ;
	    RECT 1537.9501 -2.5500 1538.8500 41.4000 ;
	    RECT 1537.9501 -3.4500 1541.2500 -2.5500 ;
      END
   END dout[1]
   PIN dout[2]
      PORT
         LAYER metal1 ;
	    RECT 1093.8000 41.4000 1095.0000 42.6000 ;
         LAYER metal2 ;
	    RECT 1093.8000 41.4000 1095.0000 42.6000 ;
	    RECT 1093.9501 -2.5500 1094.8500 41.4000 ;
	    RECT 1091.5500 -3.4500 1094.8500 -2.5500 ;
      END
   END dout[2]
   PIN dout[3]
      PORT
         LAYER metal1 ;
	    RECT 1552.2001 1181.4000 1553.4000 1182.6000 ;
         LAYER metal2 ;
	    RECT 1552.2001 1187.4000 1553.4000 1188.6000 ;
	    RECT 1552.3500 1182.6000 1553.2500 1187.4000 ;
	    RECT 1552.2001 1181.4000 1553.4000 1182.6000 ;
         LAYER metal3 ;
	    RECT 1551.9000 1188.7500 1553.7001 1188.9000 ;
	    RECT 1551.9000 1187.2500 1572.7500 1188.7500 ;
	    RECT 1551.9000 1187.1000 1553.7001 1187.2500 ;
	    RECT 1571.2500 1184.2500 1572.7500 1187.2500 ;
      END
   END dout[3]
   PIN dout[4]
      PORT
         LAYER metal1 ;
	    RECT 1540.2001 1302.4501 1541.4000 1302.6000 ;
	    RECT 1552.2001 1302.4501 1553.4000 1302.6000 ;
	    RECT 1540.2001 1301.5500 1553.4000 1302.4501 ;
	    RECT 1540.2001 1301.4000 1541.4000 1301.5500 ;
	    RECT 1552.2001 1301.4000 1553.4000 1301.5500 ;
         LAYER metal2 ;
	    RECT 1552.2001 1307.4000 1553.4000 1308.6000 ;
	    RECT 1552.3500 1302.6000 1553.2500 1307.4000 ;
	    RECT 1552.2001 1301.4000 1553.4000 1302.6000 ;
         LAYER metal3 ;
	    RECT 1551.9000 1308.7500 1553.7001 1308.9000 ;
	    RECT 1551.9000 1307.2500 1572.7500 1308.7500 ;
	    RECT 1551.9000 1307.1000 1553.7001 1307.2500 ;
	    RECT 1571.2500 1304.2500 1572.7500 1307.2500 ;
      END
   END dout[4]
   PIN dout[5]
      PORT
         LAYER metal1 ;
	    RECT 1545.0000 1421.4000 1546.2001 1422.6000 ;
         LAYER metal2 ;
	    RECT 1542.7500 1475.5500 1546.0500 1476.4501 ;
	    RECT 1545.1500 1422.6000 1546.0500 1475.5500 ;
	    RECT 1545.0000 1421.4000 1546.2001 1422.6000 ;
      END
   END dout[5]
   PIN dout[6]
      PORT
         LAYER metal1 ;
	    RECT 1542.6000 1460.4000 1543.8000 1461.6000 ;
         LAYER metal2 ;
	    RECT 1535.5500 1470.6000 1536.4501 1476.4501 ;
	    RECT 1535.4000 1469.4000 1536.6000 1470.6000 ;
	    RECT 1542.6000 1469.4000 1543.8000 1470.6000 ;
	    RECT 1542.7500 1461.6000 1543.6500 1469.4000 ;
	    RECT 1542.6000 1460.4000 1543.8000 1461.6000 ;
         LAYER metal3 ;
	    RECT 1535.1000 1470.7500 1536.9000 1470.9000 ;
	    RECT 1542.3000 1470.7500 1544.1000 1470.9000 ;
	    RECT 1535.1000 1469.2500 1544.1000 1470.7500 ;
	    RECT 1535.1000 1469.1000 1536.9000 1469.2500 ;
	    RECT 1542.3000 1469.1000 1544.1000 1469.2500 ;
      END
   END dout[6]
   PIN dout[7]
      PORT
         LAYER metal1 ;
	    RECT 1461.0000 41.4000 1462.2001 42.6000 ;
         LAYER metal2 ;
	    RECT 1461.0000 41.4000 1462.2001 42.6000 ;
	    RECT 1461.1500 -2.5500 1462.0500 41.4000 ;
	    RECT 1458.7500 -3.4500 1462.0500 -2.5500 ;
      END
   END dout[7]
   OBS
         LAYER metal1 ;
	    RECT 1.2000 1470.6000 1569.0000 1472.4000 ;
	    RECT 126.6000 1460.7001 127.8000 1469.7001 ;
	    RECT 131.4000 1463.7001 132.6000 1469.7001 ;
	    RECT 136.2000 1464.9000 137.4000 1469.7001 ;
	    RECT 138.6000 1465.5000 139.8000 1469.7001 ;
	    RECT 141.0000 1465.5000 142.2000 1469.7001 ;
	    RECT 143.4000 1465.5000 144.6000 1469.7001 ;
	    RECT 145.8000 1466.7001 147.0000 1469.7001 ;
	    RECT 148.2000 1465.5000 149.4000 1469.7001 ;
	    RECT 150.6000 1466.7001 151.8000 1469.7001 ;
	    RECT 153.0000 1465.5000 154.2000 1469.7001 ;
	    RECT 155.4000 1465.5000 156.6000 1469.7001 ;
	    RECT 157.8000 1465.5000 159.0000 1469.7001 ;
	    RECT 160.2000 1465.5000 161.4000 1469.7001 ;
	    RECT 133.5000 1463.7001 137.4000 1464.9000 ;
	    RECT 162.6000 1464.9000 163.8000 1469.7001 ;
	    RECT 142.5000 1463.7001 149.4000 1464.6000 ;
	    RECT 133.5000 1462.8000 134.7000 1463.7001 ;
	    RECT 130.2000 1461.6000 134.7000 1462.8000 ;
	    RECT 126.6000 1459.5000 139.8000 1460.7001 ;
	    RECT 142.5000 1460.1000 143.7000 1463.7001 ;
	    RECT 148.2000 1463.4000 149.4000 1463.7001 ;
	    RECT 150.6000 1463.4000 151.8000 1464.6000 ;
	    RECT 152.7000 1463.4000 153.0000 1464.6000 ;
	    RECT 157.5000 1463.4000 159.0000 1464.6000 ;
	    RECT 162.6000 1463.7001 166.2000 1464.9000 ;
	    RECT 167.4000 1463.7001 168.6000 1469.7001 ;
	    RECT 145.8000 1462.5000 147.0000 1462.8000 ;
	    RECT 148.2000 1462.2001 149.4000 1462.5000 ;
	    RECT 145.8000 1460.4000 147.0000 1461.6000 ;
	    RECT 148.2000 1461.3000 154.8000 1462.2001 ;
	    RECT 153.6000 1461.0000 154.8000 1461.3000 ;
	    RECT 126.6000 1451.1000 127.8000 1459.5000 ;
	    RECT 140.7000 1458.9000 143.7000 1460.1000 ;
	    RECT 149.4000 1458.9000 154.2000 1460.1000 ;
	    RECT 157.8000 1459.2001 159.0000 1463.4000 ;
	    RECT 165.0000 1462.8000 166.2000 1463.7001 ;
	    RECT 165.0000 1461.9000 167.7000 1462.8000 ;
	    RECT 166.5000 1460.1000 167.7000 1461.9000 ;
	    RECT 172.2000 1461.9000 173.4000 1469.7001 ;
	    RECT 174.6000 1464.0000 175.8000 1469.7001 ;
	    RECT 177.0000 1466.7001 178.2000 1469.7001 ;
	    RECT 191.4000 1466.7001 192.6000 1469.7001 ;
	    RECT 191.4000 1465.5000 192.6000 1465.8000 ;
	    RECT 177.0000 1464.4501 178.2000 1464.6000 ;
	    RECT 191.4000 1464.4501 192.6000 1464.6000 ;
	    RECT 174.6000 1462.8000 176.1000 1464.0000 ;
	    RECT 177.0000 1463.5500 192.6000 1464.4501 ;
	    RECT 177.0000 1463.4000 178.2000 1463.5500 ;
	    RECT 191.4000 1463.4000 192.6000 1463.5500 ;
	    RECT 172.2000 1461.0000 174.0000 1461.9000 ;
	    RECT 166.5000 1458.9000 172.2000 1460.1000 ;
	    RECT 128.7000 1458.0000 129.9000 1458.3000 ;
	    RECT 128.7000 1457.1000 135.3000 1458.0000 ;
	    RECT 136.2000 1457.4000 137.4000 1458.6000 ;
	    RECT 162.6000 1458.0000 163.8000 1458.9000 ;
	    RECT 173.1000 1458.0000 174.0000 1461.0000 ;
	    RECT 138.3000 1457.1000 163.8000 1458.0000 ;
	    RECT 172.8000 1457.1000 174.0000 1458.0000 ;
	    RECT 170.7000 1456.2001 171.9000 1456.5000 ;
	    RECT 131.4000 1454.4000 132.6000 1455.6000 ;
	    RECT 133.5000 1455.3000 171.9000 1456.2001 ;
	    RECT 136.5000 1455.0000 137.7000 1455.3000 ;
	    RECT 172.8000 1454.4000 173.7000 1457.1000 ;
	    RECT 174.9000 1456.2001 176.1000 1462.8000 ;
	    RECT 193.8000 1462.5000 195.0000 1469.7001 ;
	    RECT 225.0000 1463.7001 226.2000 1469.7001 ;
	    RECT 227.4000 1464.0000 228.6000 1469.7001 ;
	    RECT 229.8000 1464.9000 231.0000 1469.7001 ;
	    RECT 232.2000 1464.0000 233.4000 1469.7001 ;
	    RECT 227.4000 1463.7001 233.4000 1464.0000 ;
	    RECT 252.3000 1464.6000 253.5000 1469.7001 ;
	    RECT 252.3000 1463.7001 255.0000 1464.6000 ;
	    RECT 256.2000 1463.7001 257.4000 1469.7001 ;
	    RECT 268.2000 1466.7001 269.4000 1469.7001 ;
	    RECT 268.2000 1465.5000 269.4000 1465.8000 ;
	    RECT 225.3000 1462.5000 226.2000 1463.7001 ;
	    RECT 227.7000 1463.1000 233.1000 1463.7001 ;
	    RECT 193.8000 1461.4501 195.0000 1461.6000 ;
	    RECT 222.6000 1461.4501 223.8000 1461.6000 ;
	    RECT 193.8000 1460.5500 223.8000 1461.4501 ;
	    RECT 193.8000 1460.4000 195.0000 1460.5500 ;
	    RECT 222.6000 1460.4000 223.8000 1460.5500 ;
	    RECT 225.0000 1460.4000 226.2000 1461.6000 ;
	    RECT 227.1000 1460.4000 228.9000 1461.6000 ;
	    RECT 231.0000 1460.7001 231.3000 1462.2001 ;
	    RECT 232.2000 1460.4000 233.4000 1461.6000 ;
	    RECT 141.0000 1454.1000 142.2000 1454.4000 ;
	    RECT 134.1000 1453.5000 142.2000 1454.1000 ;
	    RECT 132.9000 1453.2001 142.2000 1453.5000 ;
	    RECT 143.7000 1453.5000 156.6000 1454.4000 ;
	    RECT 129.0000 1452.0000 131.4000 1453.2001 ;
	    RECT 132.9000 1452.3000 135.0000 1453.2001 ;
	    RECT 143.7000 1452.3000 144.6000 1453.5000 ;
	    RECT 155.4000 1453.2001 156.6000 1453.5000 ;
	    RECT 160.2000 1453.5000 173.7000 1454.4000 ;
	    RECT 174.6000 1455.0000 176.1000 1456.2001 ;
	    RECT 174.6000 1453.5000 175.8000 1455.0000 ;
	    RECT 160.2000 1453.2001 161.4000 1453.5000 ;
	    RECT 130.5000 1451.4000 131.4000 1452.0000 ;
	    RECT 135.9000 1451.4000 144.6000 1452.3000 ;
	    RECT 145.5000 1451.4000 149.4000 1452.6000 ;
	    RECT 126.6000 1450.2001 129.6000 1451.1000 ;
	    RECT 130.5000 1450.2001 136.8000 1451.4000 ;
	    RECT 128.7000 1449.3000 129.6000 1450.2001 ;
	    RECT 126.6000 1443.3000 127.8000 1449.3000 ;
	    RECT 128.7000 1448.4000 130.2000 1449.3000 ;
	    RECT 129.0000 1443.3000 130.2000 1448.4000 ;
	    RECT 131.4000 1442.4000 132.6000 1449.3000 ;
	    RECT 133.8000 1443.3000 135.0000 1450.2001 ;
	    RECT 136.2000 1443.3000 137.4000 1449.3000 ;
	    RECT 138.6000 1443.3000 139.8000 1447.5000 ;
	    RECT 141.0000 1443.3000 142.2000 1447.5000 ;
	    RECT 143.4000 1443.3000 144.6000 1450.5000 ;
	    RECT 145.8000 1443.3000 147.0000 1449.3000 ;
	    RECT 148.2000 1443.3000 149.4000 1450.5000 ;
	    RECT 150.6000 1443.3000 151.8000 1449.3000 ;
	    RECT 153.0000 1443.3000 154.2000 1452.6000 ;
	    RECT 165.0000 1451.4000 168.9000 1452.6000 ;
	    RECT 157.8000 1450.2001 164.1000 1451.4000 ;
	    RECT 155.4000 1443.3000 156.6000 1447.5000 ;
	    RECT 157.8000 1443.3000 159.0000 1447.5000 ;
	    RECT 160.2000 1443.3000 161.4000 1447.5000 ;
	    RECT 162.6000 1443.3000 163.8000 1449.3000 ;
	    RECT 165.0000 1443.3000 166.2000 1451.4000 ;
	    RECT 172.8000 1451.1000 173.7000 1453.5000 ;
	    RECT 174.6000 1452.4501 175.8000 1452.6000 ;
	    RECT 177.0000 1452.4501 178.2000 1452.6000 ;
	    RECT 174.6000 1451.5500 178.2000 1452.4501 ;
	    RECT 174.6000 1451.4000 175.8000 1451.5500 ;
	    RECT 177.0000 1451.4000 178.2000 1451.5500 ;
	    RECT 169.8000 1450.2001 173.7000 1451.1000 ;
	    RECT 167.4000 1443.3000 168.6000 1449.3000 ;
	    RECT 169.8000 1443.3000 171.0000 1450.2001 ;
	    RECT 172.2000 1443.3000 173.4000 1449.3000 ;
	    RECT 174.6000 1443.3000 175.8000 1450.5000 ;
	    RECT 177.0000 1443.3000 178.2000 1449.3000 ;
	    RECT 191.4000 1443.3000 192.6000 1449.3000 ;
	    RECT 193.8000 1443.3000 195.0000 1459.5000 ;
	    RECT 225.0000 1454.4000 226.2000 1455.6000 ;
	    RECT 228.0000 1455.3000 228.9000 1460.4000 ;
	    RECT 229.8000 1459.5000 231.0000 1459.8000 ;
	    RECT 253.8000 1459.5000 255.0000 1463.7001 ;
	    RECT 268.2000 1463.4000 269.4000 1464.6000 ;
	    RECT 256.2000 1462.5000 257.4000 1462.8000 ;
	    RECT 270.6000 1462.5000 271.8000 1469.7001 ;
	    RECT 297.0000 1463.7001 298.2000 1469.7001 ;
	    RECT 299.4000 1464.0000 300.6000 1469.7001 ;
	    RECT 301.8000 1464.9000 303.0000 1469.7001 ;
	    RECT 304.2000 1464.0000 305.4000 1469.7001 ;
	    RECT 299.4000 1463.7001 305.4000 1464.0000 ;
	    RECT 297.3000 1462.5000 298.2000 1463.7001 ;
	    RECT 299.7000 1463.1000 305.1000 1463.7001 ;
	    RECT 256.2000 1460.4000 257.4000 1461.6000 ;
	    RECT 270.6000 1461.4501 271.8000 1461.6000 ;
	    RECT 294.6000 1461.4501 295.8000 1461.6000 ;
	    RECT 270.6000 1460.5500 295.8000 1461.4501 ;
	    RECT 270.6000 1460.4000 271.8000 1460.5500 ;
	    RECT 294.6000 1460.4000 295.8000 1460.5500 ;
	    RECT 297.0000 1460.4000 298.2000 1461.6000 ;
	    RECT 299.1000 1460.4000 300.9000 1461.6000 ;
	    RECT 303.0000 1460.7001 303.3000 1462.2001 ;
	    RECT 304.2000 1461.4501 305.4000 1461.6000 ;
	    RECT 385.8000 1461.4501 387.0000 1461.6000 ;
	    RECT 304.2000 1460.5500 387.0000 1461.4501 ;
	    RECT 304.2000 1460.4000 305.4000 1460.5500 ;
	    RECT 385.8000 1460.4000 387.0000 1460.5500 ;
	    RECT 436.2000 1460.7001 437.4000 1469.7001 ;
	    RECT 441.0000 1463.7001 442.2000 1469.7001 ;
	    RECT 445.8000 1464.9000 447.0000 1469.7001 ;
	    RECT 448.2000 1465.5000 449.4000 1469.7001 ;
	    RECT 450.6000 1465.5000 451.8000 1469.7001 ;
	    RECT 453.0000 1465.5000 454.2000 1469.7001 ;
	    RECT 455.4000 1466.7001 456.6000 1469.7001 ;
	    RECT 457.8000 1465.5000 459.0000 1469.7001 ;
	    RECT 460.2000 1466.7001 461.4000 1469.7001 ;
	    RECT 462.6000 1465.5000 463.8000 1469.7001 ;
	    RECT 465.0000 1465.5000 466.2000 1469.7001 ;
	    RECT 467.4000 1465.5000 468.6000 1469.7001 ;
	    RECT 469.8000 1465.5000 471.0000 1469.7001 ;
	    RECT 443.1000 1463.7001 447.0000 1464.9000 ;
	    RECT 472.2000 1464.9000 473.4000 1469.7001 ;
	    RECT 452.1000 1463.7001 459.0000 1464.6000 ;
	    RECT 443.1000 1462.8000 444.3000 1463.7001 ;
	    RECT 439.8000 1461.6000 444.3000 1462.8000 ;
	    RECT 229.8000 1457.4000 231.0000 1458.6000 ;
	    RECT 253.8000 1458.4501 255.0000 1458.6000 ;
	    RECT 265.8000 1458.4501 267.0000 1458.6000 ;
	    RECT 253.8000 1457.5500 267.0000 1458.4501 ;
	    RECT 253.8000 1457.4000 255.0000 1457.5500 ;
	    RECT 265.8000 1457.4000 267.0000 1457.5500 ;
	    RECT 228.0000 1454.4000 229.5000 1455.3000 ;
	    RECT 226.2000 1452.6000 227.1000 1453.5000 ;
	    RECT 226.2000 1451.4000 227.4000 1452.6000 ;
	    RECT 225.9000 1443.3000 227.1000 1449.3000 ;
	    RECT 228.3000 1443.3000 229.5000 1454.4000 ;
	    RECT 232.2000 1443.3000 233.4000 1455.3000 ;
	    RECT 251.4000 1454.4000 252.6000 1455.6000 ;
	    RECT 251.4000 1453.2001 252.6000 1453.5000 ;
	    RECT 251.4000 1443.3000 252.6000 1449.3000 ;
	    RECT 253.8000 1443.3000 255.0000 1456.5000 ;
	    RECT 256.2000 1443.3000 257.4000 1449.3000 ;
	    RECT 268.2000 1443.3000 269.4000 1449.3000 ;
	    RECT 270.6000 1443.3000 271.8000 1459.5000 ;
	    RECT 292.2000 1458.4501 293.4000 1458.6000 ;
	    RECT 297.1500 1458.4501 298.0500 1460.4000 ;
	    RECT 292.2000 1457.5500 298.0500 1458.4501 ;
	    RECT 292.2000 1457.4000 293.4000 1457.5500 ;
	    RECT 297.0000 1454.4000 298.2000 1455.6000 ;
	    RECT 300.0000 1455.3000 300.9000 1460.4000 ;
	    RECT 301.8000 1459.5000 303.0000 1459.8000 ;
	    RECT 436.2000 1459.5000 449.4000 1460.7001 ;
	    RECT 452.1000 1460.1000 453.3000 1463.7001 ;
	    RECT 457.8000 1463.4000 459.0000 1463.7001 ;
	    RECT 460.2000 1463.4000 461.4000 1464.6000 ;
	    RECT 462.3000 1463.4000 462.6000 1464.6000 ;
	    RECT 467.1000 1463.4000 468.6000 1464.6000 ;
	    RECT 472.2000 1463.7001 475.8000 1464.9000 ;
	    RECT 477.0000 1463.7001 478.2000 1469.7001 ;
	    RECT 455.4000 1462.5000 456.6000 1462.8000 ;
	    RECT 457.8000 1462.2001 459.0000 1462.5000 ;
	    RECT 455.4000 1460.4000 456.6000 1461.6000 ;
	    RECT 457.8000 1461.3000 464.4000 1462.2001 ;
	    RECT 463.2000 1461.0000 464.4000 1461.3000 ;
	    RECT 301.8000 1457.4000 303.0000 1458.6000 ;
	    RECT 300.0000 1454.4000 301.5000 1455.3000 ;
	    RECT 298.2000 1452.6000 299.1000 1453.5000 ;
	    RECT 298.2000 1451.4000 299.4000 1452.6000 ;
	    RECT 297.9000 1443.3000 299.1000 1449.3000 ;
	    RECT 300.3000 1443.3000 301.5000 1454.4000 ;
	    RECT 304.2000 1443.3000 305.4000 1455.3000 ;
	    RECT 436.2000 1451.1000 437.4000 1459.5000 ;
	    RECT 450.3000 1458.9000 453.3000 1460.1000 ;
	    RECT 459.0000 1458.9000 463.8000 1460.1000 ;
	    RECT 467.4000 1459.2001 468.6000 1463.4000 ;
	    RECT 474.6000 1462.8000 475.8000 1463.7001 ;
	    RECT 474.6000 1461.9000 477.3000 1462.8000 ;
	    RECT 476.1000 1460.1000 477.3000 1461.9000 ;
	    RECT 481.8000 1461.9000 483.0000 1469.7001 ;
	    RECT 484.2000 1464.0000 485.4000 1469.7001 ;
	    RECT 486.6000 1466.7001 487.8000 1469.7001 ;
	    RECT 506.7000 1464.6000 507.9000 1469.7001 ;
	    RECT 484.2000 1462.8000 485.7000 1464.0000 ;
	    RECT 506.7000 1463.7001 509.4000 1464.6000 ;
	    RECT 510.6000 1463.7001 511.8000 1469.7001 ;
	    RECT 537.0000 1463.7001 538.2000 1469.7001 ;
	    RECT 539.4000 1464.0000 540.6000 1469.7001 ;
	    RECT 541.8000 1464.9000 543.0000 1469.7001 ;
	    RECT 544.2000 1464.0000 545.4000 1469.7001 ;
	    RECT 539.4000 1463.7001 545.4000 1464.0000 ;
	    RECT 481.8000 1461.0000 483.6000 1461.9000 ;
	    RECT 476.1000 1458.9000 481.8000 1460.1000 ;
	    RECT 438.3000 1458.0000 439.5000 1458.3000 ;
	    RECT 438.3000 1457.1000 444.9000 1458.0000 ;
	    RECT 445.8000 1457.4000 447.0000 1458.6000 ;
	    RECT 472.2000 1458.0000 473.4000 1458.9000 ;
	    RECT 482.7000 1458.0000 483.6000 1461.0000 ;
	    RECT 447.9000 1457.1000 473.4000 1458.0000 ;
	    RECT 482.4000 1457.1000 483.6000 1458.0000 ;
	    RECT 480.3000 1456.2001 481.5000 1456.5000 ;
	    RECT 441.0000 1454.4000 442.2000 1455.6000 ;
	    RECT 443.1000 1455.3000 481.5000 1456.2001 ;
	    RECT 446.1000 1455.0000 447.3000 1455.3000 ;
	    RECT 482.4000 1454.4000 483.3000 1457.1000 ;
	    RECT 484.5000 1456.2001 485.7000 1462.8000 ;
	    RECT 508.2000 1459.5000 509.4000 1463.7001 ;
	    RECT 510.6000 1462.5000 511.8000 1462.8000 ;
	    RECT 537.3000 1462.5000 538.2000 1463.7001 ;
	    RECT 539.7000 1463.1000 545.1000 1463.7001 ;
	    RECT 510.6000 1460.4000 511.8000 1461.6000 ;
	    RECT 537.0000 1460.4000 538.2000 1461.6000 ;
	    RECT 539.1000 1460.4000 540.9000 1461.6000 ;
	    RECT 543.0000 1460.7001 543.3000 1462.2001 ;
	    RECT 544.2000 1460.4000 545.4000 1461.6000 ;
	    RECT 678.6000 1460.7001 679.8000 1469.7001 ;
	    RECT 683.4000 1463.7001 684.6000 1469.7001 ;
	    RECT 688.2000 1464.9000 689.4000 1469.7001 ;
	    RECT 690.6000 1465.5000 691.8000 1469.7001 ;
	    RECT 693.0000 1465.5000 694.2000 1469.7001 ;
	    RECT 695.4000 1465.5000 696.6000 1469.7001 ;
	    RECT 697.8000 1466.7001 699.0000 1469.7001 ;
	    RECT 700.2000 1465.5000 701.4000 1469.7001 ;
	    RECT 702.6000 1466.7001 703.8000 1469.7001 ;
	    RECT 705.0000 1465.5000 706.2000 1469.7001 ;
	    RECT 707.4000 1465.5000 708.6000 1469.7001 ;
	    RECT 709.8000 1465.5000 711.0000 1469.7001 ;
	    RECT 712.2000 1465.5000 713.4000 1469.7001 ;
	    RECT 685.5000 1463.7001 689.4000 1464.9000 ;
	    RECT 714.6000 1464.9000 715.8000 1469.7001 ;
	    RECT 694.5000 1463.7001 701.4000 1464.6000 ;
	    RECT 685.5000 1462.8000 686.7000 1463.7001 ;
	    RECT 682.2000 1461.6000 686.7000 1462.8000 ;
	    RECT 508.2000 1458.4501 509.4000 1458.6000 ;
	    RECT 508.2000 1457.5500 538.0500 1458.4501 ;
	    RECT 508.2000 1457.4000 509.4000 1457.5500 ;
	    RECT 450.6000 1454.1000 451.8000 1454.4000 ;
	    RECT 443.7000 1453.5000 451.8000 1454.1000 ;
	    RECT 442.5000 1453.2001 451.8000 1453.5000 ;
	    RECT 453.3000 1453.5000 466.2000 1454.4000 ;
	    RECT 438.6000 1452.0000 441.0000 1453.2001 ;
	    RECT 442.5000 1452.3000 444.6000 1453.2001 ;
	    RECT 453.3000 1452.3000 454.2000 1453.5000 ;
	    RECT 465.0000 1453.2001 466.2000 1453.5000 ;
	    RECT 469.8000 1453.5000 483.3000 1454.4000 ;
	    RECT 484.2000 1455.0000 485.7000 1456.2001 ;
	    RECT 484.2000 1453.5000 485.4000 1455.0000 ;
	    RECT 505.8000 1454.4000 507.0000 1455.6000 ;
	    RECT 469.8000 1453.2001 471.0000 1453.5000 ;
	    RECT 440.1000 1451.4000 441.0000 1452.0000 ;
	    RECT 445.5000 1451.4000 454.2000 1452.3000 ;
	    RECT 455.1000 1451.4000 459.0000 1452.6000 ;
	    RECT 436.2000 1450.2001 439.2000 1451.1000 ;
	    RECT 440.1000 1450.2001 446.4000 1451.4000 ;
	    RECT 438.3000 1449.3000 439.2000 1450.2001 ;
	    RECT 436.2000 1443.3000 437.4000 1449.3000 ;
	    RECT 438.3000 1448.4000 439.8000 1449.3000 ;
	    RECT 438.6000 1443.3000 439.8000 1448.4000 ;
	    RECT 441.0000 1442.4000 442.2000 1449.3000 ;
	    RECT 443.4000 1443.3000 444.6000 1450.2001 ;
	    RECT 445.8000 1443.3000 447.0000 1449.3000 ;
	    RECT 448.2000 1443.3000 449.4000 1447.5000 ;
	    RECT 450.6000 1443.3000 451.8000 1447.5000 ;
	    RECT 453.0000 1443.3000 454.2000 1450.5000 ;
	    RECT 455.4000 1443.3000 456.6000 1449.3000 ;
	    RECT 457.8000 1443.3000 459.0000 1450.5000 ;
	    RECT 460.2000 1443.3000 461.4000 1449.3000 ;
	    RECT 462.6000 1443.3000 463.8000 1452.6000 ;
	    RECT 474.6000 1451.4000 478.5000 1452.6000 ;
	    RECT 467.4000 1450.2001 473.7000 1451.4000 ;
	    RECT 465.0000 1443.3000 466.2000 1447.5000 ;
	    RECT 467.4000 1443.3000 468.6000 1447.5000 ;
	    RECT 469.8000 1443.3000 471.0000 1447.5000 ;
	    RECT 472.2000 1443.3000 473.4000 1449.3000 ;
	    RECT 474.6000 1443.3000 475.8000 1451.4000 ;
	    RECT 482.4000 1451.1000 483.3000 1453.5000 ;
	    RECT 505.8000 1453.2001 507.0000 1453.5000 ;
	    RECT 484.2000 1452.4501 485.4000 1452.6000 ;
	    RECT 491.4000 1452.4501 492.6000 1452.6000 ;
	    RECT 484.2000 1451.5500 492.6000 1452.4501 ;
	    RECT 484.2000 1451.4000 485.4000 1451.5500 ;
	    RECT 491.4000 1451.4000 492.6000 1451.5500 ;
	    RECT 479.4000 1450.2001 483.3000 1451.1000 ;
	    RECT 477.0000 1443.3000 478.2000 1449.3000 ;
	    RECT 479.4000 1443.3000 480.6000 1450.2001 ;
	    RECT 481.8000 1443.3000 483.0000 1449.3000 ;
	    RECT 484.2000 1443.3000 485.4000 1450.5000 ;
	    RECT 486.6000 1443.3000 487.8000 1449.3000 ;
	    RECT 505.8000 1443.3000 507.0000 1449.3000 ;
	    RECT 508.2000 1443.3000 509.4000 1456.5000 ;
	    RECT 537.1500 1455.6000 538.0500 1457.5500 ;
	    RECT 537.0000 1454.4000 538.2000 1455.6000 ;
	    RECT 540.0000 1455.3000 540.9000 1460.4000 ;
	    RECT 541.8000 1459.5000 543.0000 1459.8000 ;
	    RECT 678.6000 1459.5000 691.8000 1460.7001 ;
	    RECT 694.5000 1460.1000 695.7000 1463.7001 ;
	    RECT 700.2000 1463.4000 701.4000 1463.7001 ;
	    RECT 702.6000 1463.4000 703.8000 1464.6000 ;
	    RECT 704.7000 1463.4000 705.0000 1464.6000 ;
	    RECT 709.5000 1463.4000 711.0000 1464.6000 ;
	    RECT 714.6000 1463.7001 718.2000 1464.9000 ;
	    RECT 719.4000 1463.7001 720.6000 1469.7001 ;
	    RECT 697.8000 1462.5000 699.0000 1462.8000 ;
	    RECT 700.2000 1462.2001 701.4000 1462.5000 ;
	    RECT 697.8000 1460.4000 699.0000 1461.6000 ;
	    RECT 700.2000 1461.3000 706.8000 1462.2001 ;
	    RECT 705.6000 1461.0000 706.8000 1461.3000 ;
	    RECT 541.8000 1458.4501 543.0000 1458.6000 ;
	    RECT 611.4000 1458.4501 612.6000 1458.6000 ;
	    RECT 541.8000 1457.5500 612.6000 1458.4501 ;
	    RECT 541.8000 1457.4000 543.0000 1457.5500 ;
	    RECT 611.4000 1457.4000 612.6000 1457.5500 ;
	    RECT 540.0000 1454.4000 541.5000 1455.3000 ;
	    RECT 538.2000 1452.6000 539.1000 1453.5000 ;
	    RECT 538.2000 1451.4000 539.4000 1452.6000 ;
	    RECT 510.6000 1443.3000 511.8000 1449.3000 ;
	    RECT 537.9000 1443.3000 539.1000 1449.3000 ;
	    RECT 540.3000 1443.3000 541.5000 1454.4000 ;
	    RECT 544.2000 1443.3000 545.4000 1455.3000 ;
	    RECT 678.6000 1451.1000 679.8000 1459.5000 ;
	    RECT 692.7000 1458.9000 695.7000 1460.1000 ;
	    RECT 701.4000 1458.9000 706.2000 1460.1000 ;
	    RECT 709.8000 1459.2001 711.0000 1463.4000 ;
	    RECT 717.0000 1462.8000 718.2000 1463.7001 ;
	    RECT 717.0000 1461.9000 719.7000 1462.8000 ;
	    RECT 718.5000 1460.1000 719.7000 1461.9000 ;
	    RECT 724.2000 1461.9000 725.4000 1469.7001 ;
	    RECT 726.6000 1464.0000 727.8000 1469.7001 ;
	    RECT 729.0000 1466.7001 730.2000 1469.7001 ;
	    RECT 853.8000 1466.7001 855.0000 1469.7001 ;
	    RECT 856.2000 1464.0000 857.4000 1469.7001 ;
	    RECT 726.6000 1462.8000 728.1000 1464.0000 ;
	    RECT 724.2000 1461.0000 726.0000 1461.9000 ;
	    RECT 718.5000 1458.9000 724.2000 1460.1000 ;
	    RECT 680.7000 1458.0000 681.9000 1458.3000 ;
	    RECT 680.7000 1457.1000 687.3000 1458.0000 ;
	    RECT 688.2000 1457.4000 689.4000 1458.6000 ;
	    RECT 714.6000 1458.0000 715.8000 1458.9000 ;
	    RECT 725.1000 1458.0000 726.0000 1461.0000 ;
	    RECT 690.3000 1457.1000 715.8000 1458.0000 ;
	    RECT 724.8000 1457.1000 726.0000 1458.0000 ;
	    RECT 722.7000 1456.2001 723.9000 1456.5000 ;
	    RECT 683.4000 1454.4000 684.6000 1455.6000 ;
	    RECT 685.5000 1455.3000 723.9000 1456.2001 ;
	    RECT 688.5000 1455.0000 689.7000 1455.3000 ;
	    RECT 724.8000 1454.4000 725.7000 1457.1000 ;
	    RECT 726.9000 1456.2001 728.1000 1462.8000 ;
	    RECT 693.0000 1454.1000 694.2000 1454.4000 ;
	    RECT 686.1000 1453.5000 694.2000 1454.1000 ;
	    RECT 684.9000 1453.2001 694.2000 1453.5000 ;
	    RECT 695.7000 1453.5000 708.6000 1454.4000 ;
	    RECT 681.0000 1452.0000 683.4000 1453.2001 ;
	    RECT 684.9000 1452.3000 687.0000 1453.2001 ;
	    RECT 695.7000 1452.3000 696.6000 1453.5000 ;
	    RECT 707.4000 1453.2001 708.6000 1453.5000 ;
	    RECT 712.2000 1453.5000 725.7000 1454.4000 ;
	    RECT 726.6000 1455.0000 728.1000 1456.2001 ;
	    RECT 855.9000 1462.8000 857.4000 1464.0000 ;
	    RECT 855.9000 1456.2001 857.1000 1462.8000 ;
	    RECT 858.6000 1461.9000 859.8000 1469.7001 ;
	    RECT 863.4000 1463.7001 864.6000 1469.7001 ;
	    RECT 868.2000 1464.9000 869.4000 1469.7001 ;
	    RECT 870.6000 1465.5000 871.8000 1469.7001 ;
	    RECT 873.0000 1465.5000 874.2000 1469.7001 ;
	    RECT 875.4000 1465.5000 876.6000 1469.7001 ;
	    RECT 877.8000 1465.5000 879.0000 1469.7001 ;
	    RECT 880.2000 1466.7001 881.4000 1469.7001 ;
	    RECT 882.6000 1465.5000 883.8000 1469.7001 ;
	    RECT 885.0000 1466.7001 886.2000 1469.7001 ;
	    RECT 887.4000 1465.5000 888.6000 1469.7001 ;
	    RECT 889.8000 1465.5000 891.0000 1469.7001 ;
	    RECT 892.2000 1465.5000 893.4000 1469.7001 ;
	    RECT 865.8000 1463.7001 869.4000 1464.9000 ;
	    RECT 894.6000 1464.9000 895.8000 1469.7001 ;
	    RECT 865.8000 1462.8000 867.0000 1463.7001 ;
	    RECT 858.0000 1461.0000 859.8000 1461.9000 ;
	    RECT 864.3000 1461.9000 867.0000 1462.8000 ;
	    RECT 873.0000 1463.4000 874.5000 1464.6000 ;
	    RECT 879.0000 1463.4000 879.3000 1464.6000 ;
	    RECT 880.2000 1463.4000 881.4000 1464.6000 ;
	    RECT 882.6000 1463.7001 889.5000 1464.6000 ;
	    RECT 894.6000 1463.7001 898.5000 1464.9000 ;
	    RECT 899.4000 1463.7001 900.6000 1469.7001 ;
	    RECT 882.6000 1463.4000 883.8000 1463.7001 ;
	    RECT 858.0000 1458.0000 858.9000 1461.0000 ;
	    RECT 864.3000 1460.1000 865.5000 1461.9000 ;
	    RECT 859.8000 1458.9000 865.5000 1460.1000 ;
	    RECT 873.0000 1459.2001 874.2000 1463.4000 ;
	    RECT 885.0000 1462.5000 886.2000 1462.8000 ;
	    RECT 882.6000 1462.2001 883.8000 1462.5000 ;
	    RECT 877.2000 1461.3000 883.8000 1462.2001 ;
	    RECT 877.2000 1461.0000 878.4000 1461.3000 ;
	    RECT 885.0000 1460.4000 886.2000 1461.6000 ;
	    RECT 888.3000 1460.1000 889.5000 1463.7001 ;
	    RECT 897.3000 1462.8000 898.5000 1463.7001 ;
	    RECT 897.3000 1461.6000 901.8000 1462.8000 ;
	    RECT 904.2000 1460.7001 905.4000 1469.7001 ;
	    RECT 935.4000 1463.7001 936.6000 1469.7001 ;
	    RECT 937.8000 1464.0000 939.0000 1469.7001 ;
	    RECT 940.2000 1464.9000 941.4000 1469.7001 ;
	    RECT 942.6000 1464.0000 943.8000 1469.7001 ;
	    RECT 1069.8000 1466.7001 1071.0000 1469.7001 ;
	    RECT 1072.2001 1464.0000 1073.4000 1469.7001 ;
	    RECT 937.8000 1463.7001 943.8000 1464.0000 ;
	    RECT 935.7000 1462.5000 936.6000 1463.7001 ;
	    RECT 938.1000 1463.1000 943.5000 1463.7001 ;
	    RECT 1071.9000 1462.8000 1073.4000 1464.0000 ;
	    RECT 877.8000 1458.9000 882.6000 1460.1000 ;
	    RECT 888.3000 1458.9000 891.3000 1460.1000 ;
	    RECT 892.2000 1459.5000 905.4000 1460.7001 ;
	    RECT 906.6000 1461.4501 907.8000 1461.6000 ;
	    RECT 935.4000 1461.4501 936.6000 1461.6000 ;
	    RECT 906.6000 1460.5500 936.6000 1461.4501 ;
	    RECT 906.6000 1460.4000 907.8000 1460.5500 ;
	    RECT 935.4000 1460.4000 936.6000 1460.5500 ;
	    RECT 937.5000 1460.4000 939.3000 1461.6000 ;
	    RECT 941.4000 1460.7001 941.7000 1462.2001 ;
	    RECT 942.6000 1460.4000 943.8000 1461.6000 ;
	    RECT 868.2000 1458.0000 869.4000 1458.9000 ;
	    RECT 858.0000 1457.1000 859.2000 1458.0000 ;
	    RECT 868.2000 1457.1000 893.7000 1458.0000 ;
	    RECT 894.6000 1457.4000 895.8000 1458.6000 ;
	    RECT 902.1000 1458.0000 903.3000 1458.3000 ;
	    RECT 896.7000 1457.1000 903.3000 1458.0000 ;
	    RECT 855.9000 1455.0000 857.4000 1456.2001 ;
	    RECT 726.6000 1453.5000 727.8000 1455.0000 ;
	    RECT 856.2000 1453.5000 857.4000 1455.0000 ;
	    RECT 858.3000 1454.4000 859.2000 1457.1000 ;
	    RECT 860.1000 1456.2001 861.3000 1456.5000 ;
	    RECT 860.1000 1455.3000 898.5000 1456.2001 ;
	    RECT 894.3000 1455.0000 895.5000 1455.3000 ;
	    RECT 899.4000 1454.4000 900.6000 1455.6000 ;
	    RECT 858.3000 1453.5000 871.8000 1454.4000 ;
	    RECT 712.2000 1453.2001 713.4000 1453.5000 ;
	    RECT 682.5000 1451.4000 683.4000 1452.0000 ;
	    RECT 687.9000 1451.4000 696.6000 1452.3000 ;
	    RECT 697.5000 1451.4000 701.4000 1452.6000 ;
	    RECT 678.6000 1450.2001 681.6000 1451.1000 ;
	    RECT 682.5000 1450.2001 688.8000 1451.4000 ;
	    RECT 680.7000 1449.3000 681.6000 1450.2001 ;
	    RECT 678.6000 1443.3000 679.8000 1449.3000 ;
	    RECT 680.7000 1448.4000 682.2000 1449.3000 ;
	    RECT 681.0000 1443.3000 682.2000 1448.4000 ;
	    RECT 683.4000 1442.4000 684.6000 1449.3000 ;
	    RECT 685.8000 1443.3000 687.0000 1450.2001 ;
	    RECT 688.2000 1443.3000 689.4000 1449.3000 ;
	    RECT 690.6000 1443.3000 691.8000 1447.5000 ;
	    RECT 693.0000 1443.3000 694.2000 1447.5000 ;
	    RECT 695.4000 1443.3000 696.6000 1450.5000 ;
	    RECT 697.8000 1443.3000 699.0000 1449.3000 ;
	    RECT 700.2000 1443.3000 701.4000 1450.5000 ;
	    RECT 702.6000 1443.3000 703.8000 1449.3000 ;
	    RECT 705.0000 1443.3000 706.2000 1452.6000 ;
	    RECT 717.0000 1451.4000 720.9000 1452.6000 ;
	    RECT 709.8000 1450.2001 716.1000 1451.4000 ;
	    RECT 707.4000 1443.3000 708.6000 1447.5000 ;
	    RECT 709.8000 1443.3000 711.0000 1447.5000 ;
	    RECT 712.2000 1443.3000 713.4000 1447.5000 ;
	    RECT 714.6000 1443.3000 715.8000 1449.3000 ;
	    RECT 717.0000 1443.3000 718.2000 1451.4000 ;
	    RECT 724.8000 1451.1000 725.7000 1453.5000 ;
	    RECT 726.6000 1451.4000 727.8000 1452.6000 ;
	    RECT 856.2000 1451.4000 857.4000 1452.6000 ;
	    RECT 721.8000 1450.2001 725.7000 1451.1000 ;
	    RECT 858.3000 1451.1000 859.2000 1453.5000 ;
	    RECT 870.6000 1453.2001 871.8000 1453.5000 ;
	    RECT 875.4000 1453.5000 888.3000 1454.4000 ;
	    RECT 875.4000 1453.2001 876.6000 1453.5000 ;
	    RECT 863.1000 1451.4000 867.0000 1452.6000 ;
	    RECT 719.4000 1443.3000 720.6000 1449.3000 ;
	    RECT 721.8000 1443.3000 723.0000 1450.2001 ;
	    RECT 724.2000 1443.3000 725.4000 1449.3000 ;
	    RECT 726.6000 1443.3000 727.8000 1450.5000 ;
	    RECT 729.0000 1443.3000 730.2000 1449.3000 ;
	    RECT 853.8000 1443.3000 855.0000 1449.3000 ;
	    RECT 856.2000 1443.3000 857.4000 1450.5000 ;
	    RECT 858.3000 1450.2001 862.2000 1451.1000 ;
	    RECT 858.6000 1443.3000 859.8000 1449.3000 ;
	    RECT 861.0000 1443.3000 862.2000 1450.2001 ;
	    RECT 863.4000 1443.3000 864.6000 1449.3000 ;
	    RECT 865.8000 1443.3000 867.0000 1451.4000 ;
	    RECT 867.9000 1450.2001 874.2000 1451.4000 ;
	    RECT 868.2000 1443.3000 869.4000 1449.3000 ;
	    RECT 870.6000 1443.3000 871.8000 1447.5000 ;
	    RECT 873.0000 1443.3000 874.2000 1447.5000 ;
	    RECT 875.4000 1443.3000 876.6000 1447.5000 ;
	    RECT 877.8000 1443.3000 879.0000 1452.6000 ;
	    RECT 882.6000 1451.4000 886.5000 1452.6000 ;
	    RECT 887.4000 1452.3000 888.3000 1453.5000 ;
	    RECT 889.8000 1454.1000 891.0000 1454.4000 ;
	    RECT 889.8000 1453.5000 897.9000 1454.1000 ;
	    RECT 889.8000 1453.2001 899.1000 1453.5000 ;
	    RECT 897.0000 1452.3000 899.1000 1453.2001 ;
	    RECT 887.4000 1451.4000 896.1000 1452.3000 ;
	    RECT 900.6000 1452.0000 903.0000 1453.2001 ;
	    RECT 900.6000 1451.4000 901.5000 1452.0000 ;
	    RECT 880.2000 1443.3000 881.4000 1449.3000 ;
	    RECT 882.6000 1443.3000 883.8000 1450.5000 ;
	    RECT 885.0000 1443.3000 886.2000 1449.3000 ;
	    RECT 887.4000 1443.3000 888.6000 1450.5000 ;
	    RECT 895.2000 1450.2001 901.5000 1451.4000 ;
	    RECT 904.2000 1451.1000 905.4000 1459.5000 ;
	    RECT 935.4000 1454.4000 936.6000 1455.6000 ;
	    RECT 938.4000 1455.3000 939.3000 1460.4000 ;
	    RECT 940.2000 1459.5000 941.4000 1459.8000 ;
	    RECT 940.2000 1457.4000 941.4000 1458.6000 ;
	    RECT 1071.9000 1456.2001 1073.1000 1462.8000 ;
	    RECT 1074.6000 1461.9000 1075.8000 1469.7001 ;
	    RECT 1079.4000 1463.7001 1080.6000 1469.7001 ;
	    RECT 1084.2001 1464.9000 1085.4000 1469.7001 ;
	    RECT 1086.6000 1465.5000 1087.8000 1469.7001 ;
	    RECT 1089.0000 1465.5000 1090.2001 1469.7001 ;
	    RECT 1091.4000 1465.5000 1092.6000 1469.7001 ;
	    RECT 1093.8000 1465.5000 1095.0000 1469.7001 ;
	    RECT 1096.2001 1466.7001 1097.4000 1469.7001 ;
	    RECT 1098.6000 1465.5000 1099.8000 1469.7001 ;
	    RECT 1101.0000 1466.7001 1102.2001 1469.7001 ;
	    RECT 1103.4000 1465.5000 1104.6000 1469.7001 ;
	    RECT 1105.8000 1465.5000 1107.0000 1469.7001 ;
	    RECT 1108.2001 1465.5000 1109.4000 1469.7001 ;
	    RECT 1081.8000 1463.7001 1085.4000 1464.9000 ;
	    RECT 1110.6000 1464.9000 1111.8000 1469.7001 ;
	    RECT 1081.8000 1462.8000 1083.0000 1463.7001 ;
	    RECT 1074.0000 1461.0000 1075.8000 1461.9000 ;
	    RECT 1080.3000 1461.9000 1083.0000 1462.8000 ;
	    RECT 1089.0000 1463.4000 1090.5000 1464.6000 ;
	    RECT 1095.0000 1463.4000 1095.3000 1464.6000 ;
	    RECT 1096.2001 1463.4000 1097.4000 1464.6000 ;
	    RECT 1098.6000 1463.7001 1105.5000 1464.6000 ;
	    RECT 1110.6000 1463.7001 1114.5000 1464.9000 ;
	    RECT 1115.4000 1463.7001 1116.6000 1469.7001 ;
	    RECT 1098.6000 1463.4000 1099.8000 1463.7001 ;
	    RECT 1074.0000 1458.0000 1074.9000 1461.0000 ;
	    RECT 1080.3000 1460.1000 1081.5000 1461.9000 ;
	    RECT 1075.8000 1458.9000 1081.5000 1460.1000 ;
	    RECT 1089.0000 1459.2001 1090.2001 1463.4000 ;
	    RECT 1101.0000 1462.5000 1102.2001 1462.8000 ;
	    RECT 1098.6000 1462.2001 1099.8000 1462.5000 ;
	    RECT 1093.2001 1461.3000 1099.8000 1462.2001 ;
	    RECT 1093.2001 1461.0000 1094.4000 1461.3000 ;
	    RECT 1101.0000 1460.4000 1102.2001 1461.6000 ;
	    RECT 1104.3000 1460.1000 1105.5000 1463.7001 ;
	    RECT 1113.3000 1462.8000 1114.5000 1463.7001 ;
	    RECT 1113.3000 1461.6000 1117.8000 1462.8000 ;
	    RECT 1120.2001 1460.7001 1121.4000 1469.7001 ;
	    RECT 1146.6000 1463.7001 1147.8000 1469.7001 ;
	    RECT 1150.5000 1464.6000 1151.7001 1469.7001 ;
	    RECT 1149.0000 1463.7001 1151.7001 1464.6000 ;
	    RECT 1177.8000 1463.7001 1179.0000 1469.7001 ;
	    RECT 1180.2001 1464.0000 1181.4000 1469.7001 ;
	    RECT 1182.6000 1464.9000 1183.8000 1469.7001 ;
	    RECT 1185.0000 1464.0000 1186.2001 1469.7001 ;
	    RECT 1180.2001 1463.7001 1186.2001 1464.0000 ;
	    RECT 1146.6000 1462.5000 1147.8000 1462.8000 ;
	    RECT 1093.8000 1458.9000 1098.6000 1460.1000 ;
	    RECT 1104.3000 1458.9000 1107.3000 1460.1000 ;
	    RECT 1108.2001 1459.5000 1121.4000 1460.7001 ;
	    RECT 1146.6000 1460.4000 1147.8000 1461.6000 ;
	    RECT 1149.0000 1459.5000 1150.2001 1463.7001 ;
	    RECT 1178.1000 1462.5000 1179.0000 1463.7001 ;
	    RECT 1180.5000 1463.1000 1185.9000 1463.7001 ;
	    RECT 1197.0000 1462.5000 1198.2001 1469.7001 ;
	    RECT 1199.4000 1466.7001 1200.6000 1469.7001 ;
	    RECT 1199.4000 1465.5000 1200.6000 1465.8000 ;
	    RECT 1199.4000 1463.4000 1200.6000 1464.6000 ;
	    RECT 1252.2001 1463.7001 1253.4000 1469.7001 ;
	    RECT 1254.6000 1462.8000 1255.8000 1469.7001 ;
	    RECT 1257.0000 1463.7001 1258.2001 1469.7001 ;
	    RECT 1259.4000 1462.8000 1260.6000 1469.7001 ;
	    RECT 1261.8000 1463.7001 1263.0000 1469.7001 ;
	    RECT 1264.2001 1462.8000 1265.4000 1469.7001 ;
	    RECT 1266.6000 1463.7001 1267.8000 1469.7001 ;
	    RECT 1269.0000 1462.8000 1270.2001 1469.7001 ;
	    RECT 1271.4000 1463.7001 1272.6000 1469.7001 ;
	    RECT 1177.8000 1460.4000 1179.0000 1461.6000 ;
	    RECT 1179.9000 1460.4000 1181.7001 1461.6000 ;
	    RECT 1183.8000 1460.7001 1184.1000 1462.2001 ;
	    RECT 1254.6000 1461.6000 1257.3000 1462.8000 ;
	    RECT 1259.4000 1461.6000 1262.7001 1462.8000 ;
	    RECT 1264.2001 1461.6000 1267.5000 1462.8000 ;
	    RECT 1269.0000 1461.6000 1272.6000 1462.8000 ;
	    RECT 1290.6000 1462.5000 1291.8000 1469.7001 ;
	    RECT 1293.0000 1463.7001 1294.2001 1469.7001 ;
	    RECT 1295.4000 1462.8000 1296.6000 1469.7001 ;
	    RECT 1314.6000 1463.7001 1315.8000 1469.7001 ;
	    RECT 1318.5000 1464.6000 1319.7001 1469.7001 ;
	    RECT 1333.8000 1466.7001 1335.0000 1469.7001 ;
	    RECT 1333.8000 1465.5000 1335.0000 1465.8000 ;
	    RECT 1317.0000 1463.7001 1319.7001 1464.6000 ;
	    RECT 1185.0000 1460.4000 1186.2001 1461.6000 ;
	    RECT 1197.0000 1461.4501 1198.2001 1461.6000 ;
	    RECT 1187.5500 1460.5500 1198.2001 1461.4501 ;
	    RECT 1084.2001 1458.0000 1085.4000 1458.9000 ;
	    RECT 1074.0000 1457.1000 1075.2001 1458.0000 ;
	    RECT 1084.2001 1457.1000 1109.7001 1458.0000 ;
	    RECT 1110.6000 1457.4000 1111.8000 1458.6000 ;
	    RECT 1118.1000 1458.0000 1119.3000 1458.3000 ;
	    RECT 1112.7001 1457.1000 1119.3000 1458.0000 ;
	    RECT 938.4000 1454.4000 939.9000 1455.3000 ;
	    RECT 936.6000 1452.6000 937.5000 1453.5000 ;
	    RECT 936.6000 1451.4000 937.8000 1452.6000 ;
	    RECT 902.4000 1450.2001 905.4000 1451.1000 ;
	    RECT 889.8000 1443.3000 891.0000 1447.5000 ;
	    RECT 892.2000 1443.3000 893.4000 1447.5000 ;
	    RECT 894.6000 1443.3000 895.8000 1449.3000 ;
	    RECT 897.0000 1443.3000 898.2000 1450.2001 ;
	    RECT 902.4000 1449.3000 903.3000 1450.2001 ;
	    RECT 899.4000 1442.4000 900.6000 1449.3000 ;
	    RECT 901.8000 1448.4000 903.3000 1449.3000 ;
	    RECT 901.8000 1443.3000 903.0000 1448.4000 ;
	    RECT 904.2000 1443.3000 905.4000 1449.3000 ;
	    RECT 936.3000 1443.3000 937.5000 1449.3000 ;
	    RECT 938.7000 1443.3000 939.9000 1454.4000 ;
	    RECT 942.6000 1443.3000 943.8000 1455.3000 ;
	    RECT 1071.9000 1455.0000 1073.4000 1456.2001 ;
	    RECT 1072.2001 1453.5000 1073.4000 1455.0000 ;
	    RECT 1074.3000 1454.4000 1075.2001 1457.1000 ;
	    RECT 1076.1000 1456.2001 1077.3000 1456.5000 ;
	    RECT 1076.1000 1455.3000 1114.5000 1456.2001 ;
	    RECT 1110.3000 1455.0000 1111.5000 1455.3000 ;
	    RECT 1115.4000 1454.4000 1116.6000 1455.6000 ;
	    RECT 1074.3000 1453.5000 1087.8000 1454.4000 ;
	    RECT 1069.8000 1452.4501 1071.0000 1452.6000 ;
	    RECT 1072.2001 1452.4501 1073.4000 1452.6000 ;
	    RECT 1069.8000 1451.5500 1073.4000 1452.4501 ;
	    RECT 1069.8000 1451.4000 1071.0000 1451.5500 ;
	    RECT 1072.2001 1451.4000 1073.4000 1451.5500 ;
	    RECT 1074.3000 1451.1000 1075.2001 1453.5000 ;
	    RECT 1086.6000 1453.2001 1087.8000 1453.5000 ;
	    RECT 1091.4000 1453.5000 1104.3000 1454.4000 ;
	    RECT 1091.4000 1453.2001 1092.6000 1453.5000 ;
	    RECT 1079.1000 1451.4000 1083.0000 1452.6000 ;
	    RECT 1069.8000 1443.3000 1071.0000 1449.3000 ;
	    RECT 1072.2001 1443.3000 1073.4000 1450.5000 ;
	    RECT 1074.3000 1450.2001 1078.2001 1451.1000 ;
	    RECT 1074.6000 1443.3000 1075.8000 1449.3000 ;
	    RECT 1077.0000 1443.3000 1078.2001 1450.2001 ;
	    RECT 1079.4000 1443.3000 1080.6000 1449.3000 ;
	    RECT 1081.8000 1443.3000 1083.0000 1451.4000 ;
	    RECT 1083.9000 1450.2001 1090.2001 1451.4000 ;
	    RECT 1084.2001 1443.3000 1085.4000 1449.3000 ;
	    RECT 1086.6000 1443.3000 1087.8000 1447.5000 ;
	    RECT 1089.0000 1443.3000 1090.2001 1447.5000 ;
	    RECT 1091.4000 1443.3000 1092.6000 1447.5000 ;
	    RECT 1093.8000 1443.3000 1095.0000 1452.6000 ;
	    RECT 1098.6000 1451.4000 1102.5000 1452.6000 ;
	    RECT 1103.4000 1452.3000 1104.3000 1453.5000 ;
	    RECT 1105.8000 1454.1000 1107.0000 1454.4000 ;
	    RECT 1105.8000 1453.5000 1113.9000 1454.1000 ;
	    RECT 1105.8000 1453.2001 1115.1000 1453.5000 ;
	    RECT 1113.0000 1452.3000 1115.1000 1453.2001 ;
	    RECT 1103.4000 1451.4000 1112.1000 1452.3000 ;
	    RECT 1116.6000 1452.0000 1119.0000 1453.2001 ;
	    RECT 1116.6000 1451.4000 1117.5000 1452.0000 ;
	    RECT 1096.2001 1443.3000 1097.4000 1449.3000 ;
	    RECT 1098.6000 1443.3000 1099.8000 1450.5000 ;
	    RECT 1101.0000 1443.3000 1102.2001 1449.3000 ;
	    RECT 1103.4000 1443.3000 1104.6000 1450.5000 ;
	    RECT 1111.2001 1450.2001 1117.5000 1451.4000 ;
	    RECT 1120.2001 1451.1000 1121.4000 1459.5000 ;
	    RECT 1149.0000 1458.4501 1150.2001 1458.6000 ;
	    RECT 1149.0000 1457.5500 1178.8500 1458.4501 ;
	    RECT 1149.0000 1457.4000 1150.2001 1457.5500 ;
	    RECT 1118.4000 1450.2001 1121.4000 1451.1000 ;
	    RECT 1105.8000 1443.3000 1107.0000 1447.5000 ;
	    RECT 1108.2001 1443.3000 1109.4000 1447.5000 ;
	    RECT 1110.6000 1443.3000 1111.8000 1449.3000 ;
	    RECT 1113.0000 1443.3000 1114.2001 1450.2001 ;
	    RECT 1118.4000 1449.3000 1119.3000 1450.2001 ;
	    RECT 1115.4000 1442.4000 1116.6000 1449.3000 ;
	    RECT 1117.8000 1448.4000 1119.3000 1449.3000 ;
	    RECT 1117.8000 1443.3000 1119.0000 1448.4000 ;
	    RECT 1120.2001 1443.3000 1121.4000 1449.3000 ;
	    RECT 1146.6000 1443.3000 1147.8000 1449.3000 ;
	    RECT 1149.0000 1443.3000 1150.2001 1456.5000 ;
	    RECT 1177.9501 1455.6000 1178.8500 1457.5500 ;
	    RECT 1177.8000 1454.4000 1179.0000 1455.6000 ;
	    RECT 1180.8000 1455.3000 1181.7001 1460.4000 ;
	    RECT 1182.6000 1459.5000 1183.8000 1459.8000 ;
	    RECT 1182.6000 1458.4501 1183.8000 1458.6000 ;
	    RECT 1187.5500 1458.4501 1188.4501 1460.5500 ;
	    RECT 1197.0000 1460.4000 1198.2001 1460.5500 ;
	    RECT 1252.2001 1460.4000 1253.4000 1461.6000 ;
	    RECT 1256.1000 1460.7001 1257.3000 1461.6000 ;
	    RECT 1261.5000 1460.7001 1262.7001 1461.6000 ;
	    RECT 1266.3000 1460.7001 1267.5000 1461.6000 ;
	    RECT 1254.3000 1459.5000 1254.9000 1460.7001 ;
	    RECT 1256.1000 1459.5000 1260.0000 1460.7001 ;
	    RECT 1261.5000 1459.5000 1265.1000 1460.7001 ;
	    RECT 1266.3000 1459.5000 1270.2001 1460.7001 ;
	    RECT 1271.4000 1459.5000 1272.6000 1461.6000 ;
	    RECT 1293.3000 1461.9000 1296.6000 1462.8000 ;
	    RECT 1314.6000 1462.5000 1315.8000 1462.8000 ;
	    RECT 1182.6000 1457.5500 1188.4501 1458.4501 ;
	    RECT 1182.6000 1457.4000 1183.8000 1457.5500 ;
	    RECT 1180.8000 1454.4000 1182.3000 1455.3000 ;
	    RECT 1151.4000 1453.2001 1152.6000 1453.5000 ;
	    RECT 1179.0000 1452.6000 1179.9000 1453.5000 ;
	    RECT 1179.0000 1451.4000 1180.2001 1452.6000 ;
	    RECT 1151.4000 1443.3000 1152.6000 1449.3000 ;
	    RECT 1178.7001 1443.3000 1179.9000 1449.3000 ;
	    RECT 1181.1000 1443.3000 1182.3000 1454.4000 ;
	    RECT 1185.0000 1443.3000 1186.2001 1455.3000 ;
	    RECT 1197.0000 1443.3000 1198.2001 1459.5000 ;
	    RECT 1256.1000 1457.4000 1257.3000 1459.5000 ;
	    RECT 1261.5000 1457.4000 1262.7001 1459.5000 ;
	    RECT 1266.3000 1457.4000 1267.5000 1459.5000 ;
	    RECT 1290.6000 1458.6000 1291.8000 1459.5000 ;
	    RECT 1271.4000 1458.4501 1272.6000 1458.6000 ;
	    RECT 1285.8000 1458.4501 1287.0000 1458.6000 ;
	    RECT 1271.4000 1457.5500 1287.0000 1458.4501 ;
	    RECT 1271.4000 1457.4000 1272.6000 1457.5500 ;
	    RECT 1285.8000 1457.4000 1287.0000 1457.5500 ;
	    RECT 1254.6000 1456.2001 1257.3000 1457.4000 ;
	    RECT 1259.4000 1456.2001 1262.7001 1457.4000 ;
	    RECT 1264.2001 1456.2001 1267.5000 1457.4000 ;
	    RECT 1269.0000 1456.5000 1270.5000 1457.4000 ;
	    RECT 1269.0000 1456.2001 1272.6000 1456.5000 ;
	    RECT 1199.4000 1443.3000 1200.6000 1449.3000 ;
	    RECT 1252.2001 1443.3000 1253.4000 1455.3000 ;
	    RECT 1254.6000 1443.3000 1255.8000 1456.2001 ;
	    RECT 1257.0000 1443.3000 1258.2001 1455.3000 ;
	    RECT 1259.4000 1443.3000 1260.6000 1456.2001 ;
	    RECT 1261.8000 1443.3000 1263.0000 1455.3000 ;
	    RECT 1264.2001 1443.3000 1265.4000 1456.2001 ;
	    RECT 1266.6000 1443.3000 1267.8000 1455.3000 ;
	    RECT 1269.0000 1443.3000 1270.2001 1456.2001 ;
	    RECT 1290.6000 1455.3000 1291.5000 1458.6000 ;
	    RECT 1293.3000 1457.4000 1294.2001 1461.9000 ;
	    RECT 1314.6000 1460.4000 1315.8000 1461.6000 ;
	    RECT 1295.4000 1459.5000 1296.6000 1459.8000 ;
	    RECT 1317.0000 1459.5000 1318.2001 1463.7001 ;
	    RECT 1333.8000 1463.4000 1335.0000 1464.6000 ;
	    RECT 1336.2001 1462.5000 1337.4000 1469.7001 ;
	    RECT 1336.2001 1461.4501 1337.4000 1461.6000 ;
	    RECT 1374.6000 1461.4501 1375.8000 1461.6000 ;
	    RECT 1336.2001 1460.5500 1375.8000 1461.4501 ;
	    RECT 1336.2001 1460.4000 1337.4000 1460.5500 ;
	    RECT 1374.6000 1460.4000 1375.8000 1460.5500 ;
	    RECT 1468.2001 1460.7001 1469.4000 1469.7001 ;
	    RECT 1473.0000 1463.7001 1474.2001 1469.7001 ;
	    RECT 1477.8000 1464.9000 1479.0000 1469.7001 ;
	    RECT 1480.2001 1465.5000 1481.4000 1469.7001 ;
	    RECT 1482.6000 1465.5000 1483.8000 1469.7001 ;
	    RECT 1485.0000 1465.5000 1486.2001 1469.7001 ;
	    RECT 1487.4000 1466.7001 1488.6000 1469.7001 ;
	    RECT 1489.8000 1465.5000 1491.0000 1469.7001 ;
	    RECT 1492.2001 1466.7001 1493.4000 1469.7001 ;
	    RECT 1494.6000 1465.5000 1495.8000 1469.7001 ;
	    RECT 1497.0000 1465.5000 1498.2001 1469.7001 ;
	    RECT 1499.4000 1465.5000 1500.6000 1469.7001 ;
	    RECT 1501.8000 1465.5000 1503.0000 1469.7001 ;
	    RECT 1475.1000 1463.7001 1479.0000 1464.9000 ;
	    RECT 1504.2001 1464.9000 1505.4000 1469.7001 ;
	    RECT 1484.1000 1463.7001 1491.0000 1464.6000 ;
	    RECT 1475.1000 1462.8000 1476.3000 1463.7001 ;
	    RECT 1471.8000 1461.6000 1476.3000 1462.8000 ;
	    RECT 1468.2001 1459.5000 1481.4000 1460.7001 ;
	    RECT 1484.1000 1460.1000 1485.3000 1463.7001 ;
	    RECT 1489.8000 1463.4000 1491.0000 1463.7001 ;
	    RECT 1492.2001 1463.4000 1493.4000 1464.6000 ;
	    RECT 1494.3000 1463.4000 1494.6000 1464.6000 ;
	    RECT 1499.1000 1463.4000 1500.6000 1464.6000 ;
	    RECT 1504.2001 1463.7001 1507.8000 1464.9000 ;
	    RECT 1509.0000 1463.7001 1510.2001 1469.7001 ;
	    RECT 1487.4000 1462.5000 1488.6000 1462.8000 ;
	    RECT 1489.8000 1462.2001 1491.0000 1462.5000 ;
	    RECT 1487.4000 1460.4000 1488.6000 1461.6000 ;
	    RECT 1489.8000 1461.3000 1496.4000 1462.2001 ;
	    RECT 1495.2001 1461.0000 1496.4000 1461.3000 ;
	    RECT 1295.4000 1458.4501 1296.6000 1458.6000 ;
	    RECT 1312.2001 1458.4501 1313.4000 1458.6000 ;
	    RECT 1295.4000 1457.5500 1313.4000 1458.4501 ;
	    RECT 1295.4000 1457.4000 1296.6000 1457.5500 ;
	    RECT 1312.2001 1457.4000 1313.4000 1457.5500 ;
	    RECT 1317.0000 1458.4501 1318.2001 1458.6000 ;
	    RECT 1331.4000 1458.4501 1332.6000 1458.6000 ;
	    RECT 1317.0000 1457.5500 1332.6000 1458.4501 ;
	    RECT 1317.0000 1457.4000 1318.2001 1457.5500 ;
	    RECT 1331.4000 1457.4000 1332.6000 1457.5500 ;
	    RECT 1292.4000 1456.2001 1294.2001 1457.4000 ;
	    RECT 1293.3000 1455.3000 1294.2001 1456.2001 ;
	    RECT 1271.4000 1443.3000 1272.6000 1455.3000 ;
	    RECT 1290.6000 1443.3000 1291.8000 1455.3000 ;
	    RECT 1293.3000 1454.4000 1296.6000 1455.3000 ;
	    RECT 1293.0000 1443.3000 1294.2001 1453.5000 ;
	    RECT 1295.4000 1443.3000 1296.6000 1454.4000 ;
	    RECT 1314.6000 1443.3000 1315.8000 1449.3000 ;
	    RECT 1317.0000 1443.3000 1318.2001 1456.5000 ;
	    RECT 1319.4000 1453.2001 1320.6000 1453.5000 ;
	    RECT 1319.4000 1443.3000 1320.6000 1449.3000 ;
	    RECT 1333.8000 1443.3000 1335.0000 1449.3000 ;
	    RECT 1336.2001 1443.3000 1337.4000 1459.5000 ;
	    RECT 1468.2001 1451.1000 1469.4000 1459.5000 ;
	    RECT 1482.3000 1458.9000 1485.3000 1460.1000 ;
	    RECT 1491.0000 1458.9000 1495.8000 1460.1000 ;
	    RECT 1499.4000 1459.2001 1500.6000 1463.4000 ;
	    RECT 1506.6000 1462.8000 1507.8000 1463.7001 ;
	    RECT 1506.6000 1461.9000 1509.3000 1462.8000 ;
	    RECT 1508.1000 1460.1000 1509.3000 1461.9000 ;
	    RECT 1513.8000 1461.9000 1515.0000 1469.7001 ;
	    RECT 1516.2001 1464.0000 1517.4000 1469.7001 ;
	    RECT 1518.6000 1466.7001 1519.8000 1469.7001 ;
	    RECT 1516.2001 1462.8000 1517.7001 1464.0000 ;
	    RECT 1513.8000 1461.0000 1515.6000 1461.9000 ;
	    RECT 1508.1000 1458.9000 1513.8000 1460.1000 ;
	    RECT 1470.3000 1458.0000 1471.5000 1458.3000 ;
	    RECT 1470.3000 1457.1000 1476.9000 1458.0000 ;
	    RECT 1477.8000 1457.4000 1479.0000 1458.6000 ;
	    RECT 1504.2001 1458.0000 1505.4000 1458.9000 ;
	    RECT 1514.7001 1458.0000 1515.6000 1461.0000 ;
	    RECT 1479.9000 1457.1000 1505.4000 1458.0000 ;
	    RECT 1514.4000 1457.1000 1515.6000 1458.0000 ;
	    RECT 1512.3000 1456.2001 1513.5000 1456.5000 ;
	    RECT 1473.0000 1454.4000 1474.2001 1455.6000 ;
	    RECT 1475.1000 1455.3000 1513.5000 1456.2001 ;
	    RECT 1478.1000 1455.0000 1479.3000 1455.3000 ;
	    RECT 1514.4000 1454.4000 1515.3000 1457.1000 ;
	    RECT 1516.5000 1456.2001 1517.7001 1462.8000 ;
	    RECT 1537.8000 1462.8000 1539.0000 1469.7001 ;
	    RECT 1540.2001 1463.7001 1541.4000 1469.7001 ;
	    RECT 1537.8000 1461.9000 1541.1000 1462.8000 ;
	    RECT 1542.6000 1462.5000 1543.8000 1469.7001 ;
	    RECT 1562.7001 1464.6000 1563.9000 1469.7001 ;
	    RECT 1562.7001 1463.7001 1565.4000 1464.6000 ;
	    RECT 1566.6000 1463.7001 1567.8000 1469.7001 ;
	    RECT 1537.8000 1459.5000 1539.0000 1459.8000 ;
	    RECT 1523.4000 1458.4501 1524.6000 1458.6000 ;
	    RECT 1537.8000 1458.4501 1539.0000 1458.6000 ;
	    RECT 1523.4000 1457.5500 1539.0000 1458.4501 ;
	    RECT 1523.4000 1457.4000 1524.6000 1457.5500 ;
	    RECT 1537.8000 1457.4000 1539.0000 1457.5500 ;
	    RECT 1540.2001 1457.4000 1541.1000 1461.9000 ;
	    RECT 1564.2001 1459.5000 1565.4000 1463.7001 ;
	    RECT 1566.6000 1462.5000 1567.8000 1462.8000 ;
	    RECT 1566.6000 1460.4000 1567.8000 1461.6000 ;
	    RECT 1542.6000 1458.6000 1543.8000 1459.5000 ;
	    RECT 1482.6000 1454.1000 1483.8000 1454.4000 ;
	    RECT 1475.7001 1453.5000 1483.8000 1454.1000 ;
	    RECT 1474.5000 1453.2001 1483.8000 1453.5000 ;
	    RECT 1485.3000 1453.5000 1498.2001 1454.4000 ;
	    RECT 1470.6000 1452.0000 1473.0000 1453.2001 ;
	    RECT 1474.5000 1452.3000 1476.6000 1453.2001 ;
	    RECT 1485.3000 1452.3000 1486.2001 1453.5000 ;
	    RECT 1497.0000 1453.2001 1498.2001 1453.5000 ;
	    RECT 1501.8000 1453.5000 1515.3000 1454.4000 ;
	    RECT 1516.2001 1455.0000 1517.7001 1456.2001 ;
	    RECT 1540.2001 1456.2001 1542.0000 1457.4000 ;
	    RECT 1540.2001 1455.3000 1541.1000 1456.2001 ;
	    RECT 1542.9000 1455.3000 1543.8000 1458.6000 ;
	    RECT 1564.2001 1457.4000 1565.4000 1458.6000 ;
	    RECT 1516.2001 1453.5000 1517.4000 1455.0000 ;
	    RECT 1537.8000 1454.4000 1541.1000 1455.3000 ;
	    RECT 1501.8000 1453.2001 1503.0000 1453.5000 ;
	    RECT 1472.1000 1451.4000 1473.0000 1452.0000 ;
	    RECT 1477.5000 1451.4000 1486.2001 1452.3000 ;
	    RECT 1487.1000 1451.4000 1491.0000 1452.6000 ;
	    RECT 1468.2001 1450.2001 1471.2001 1451.1000 ;
	    RECT 1472.1000 1450.2001 1478.4000 1451.4000 ;
	    RECT 1470.3000 1449.3000 1471.2001 1450.2001 ;
	    RECT 1468.2001 1443.3000 1469.4000 1449.3000 ;
	    RECT 1470.3000 1448.4000 1471.8000 1449.3000 ;
	    RECT 1470.6000 1443.3000 1471.8000 1448.4000 ;
	    RECT 1473.0000 1442.4000 1474.2001 1449.3000 ;
	    RECT 1475.4000 1443.3000 1476.6000 1450.2001 ;
	    RECT 1477.8000 1443.3000 1479.0000 1449.3000 ;
	    RECT 1480.2001 1443.3000 1481.4000 1447.5000 ;
	    RECT 1482.6000 1443.3000 1483.8000 1447.5000 ;
	    RECT 1485.0000 1443.3000 1486.2001 1450.5000 ;
	    RECT 1487.4000 1443.3000 1488.6000 1449.3000 ;
	    RECT 1489.8000 1443.3000 1491.0000 1450.5000 ;
	    RECT 1492.2001 1443.3000 1493.4000 1449.3000 ;
	    RECT 1494.6000 1443.3000 1495.8000 1452.6000 ;
	    RECT 1506.6000 1451.4000 1510.5000 1452.6000 ;
	    RECT 1499.4000 1450.2001 1505.7001 1451.4000 ;
	    RECT 1497.0000 1443.3000 1498.2001 1447.5000 ;
	    RECT 1499.4000 1443.3000 1500.6000 1447.5000 ;
	    RECT 1501.8000 1443.3000 1503.0000 1447.5000 ;
	    RECT 1504.2001 1443.3000 1505.4000 1449.3000 ;
	    RECT 1506.6000 1443.3000 1507.8000 1451.4000 ;
	    RECT 1514.4000 1451.1000 1515.3000 1453.5000 ;
	    RECT 1516.2001 1452.4501 1517.4000 1452.6000 ;
	    RECT 1523.4000 1452.4501 1524.6000 1452.6000 ;
	    RECT 1516.2001 1451.5500 1524.6000 1452.4501 ;
	    RECT 1516.2001 1451.4000 1517.4000 1451.5500 ;
	    RECT 1523.4000 1451.4000 1524.6000 1451.5500 ;
	    RECT 1511.4000 1450.2001 1515.3000 1451.1000 ;
	    RECT 1509.0000 1443.3000 1510.2001 1449.3000 ;
	    RECT 1511.4000 1443.3000 1512.6000 1450.2001 ;
	    RECT 1513.8000 1443.3000 1515.0000 1449.3000 ;
	    RECT 1516.2001 1443.3000 1517.4000 1450.5000 ;
	    RECT 1518.6000 1443.3000 1519.8000 1449.3000 ;
	    RECT 1537.8000 1443.3000 1539.0000 1454.4000 ;
	    RECT 1540.2001 1443.3000 1541.4000 1453.5000 ;
	    RECT 1542.6000 1443.3000 1543.8000 1455.3000 ;
	    RECT 1557.0000 1455.4501 1558.2001 1455.6000 ;
	    RECT 1561.8000 1455.4501 1563.0000 1455.6000 ;
	    RECT 1557.0000 1454.5500 1563.0000 1455.4501 ;
	    RECT 1557.0000 1454.4000 1558.2001 1454.5500 ;
	    RECT 1561.8000 1454.4000 1563.0000 1454.5500 ;
	    RECT 1561.8000 1453.2001 1563.0000 1453.5000 ;
	    RECT 1561.8000 1443.3000 1563.0000 1449.3000 ;
	    RECT 1564.2001 1443.3000 1565.4000 1456.5000 ;
	    RECT 1566.6000 1443.3000 1567.8000 1449.3000 ;
	    RECT 1.2000 1440.6000 1569.0000 1442.4000 ;
	    RECT 124.2000 1433.7001 125.4000 1439.7001 ;
	    RECT 126.6000 1434.6000 127.8000 1439.7001 ;
	    RECT 126.3000 1433.7001 127.8000 1434.6000 ;
	    RECT 129.0000 1433.7001 130.2000 1440.6000 ;
	    RECT 126.3000 1432.8000 127.2000 1433.7001 ;
	    RECT 131.4000 1432.8000 132.6000 1439.7001 ;
	    RECT 133.8000 1433.7001 135.0000 1439.7001 ;
	    RECT 136.2000 1435.5000 137.4000 1439.7001 ;
	    RECT 138.6000 1435.5000 139.8000 1439.7001 ;
	    RECT 124.2000 1431.9000 127.2000 1432.8000 ;
	    RECT 124.2000 1423.5000 125.4000 1431.9000 ;
	    RECT 128.1000 1431.6000 134.4000 1432.8000 ;
	    RECT 141.0000 1432.5000 142.2000 1439.7001 ;
	    RECT 143.4000 1433.7001 144.6000 1439.7001 ;
	    RECT 145.8000 1432.5000 147.0000 1439.7001 ;
	    RECT 148.2000 1433.7001 149.4000 1439.7001 ;
	    RECT 128.1000 1431.0000 129.0000 1431.6000 ;
	    RECT 126.6000 1429.8000 129.0000 1431.0000 ;
	    RECT 133.5000 1430.7001 142.2000 1431.6000 ;
	    RECT 130.5000 1429.8000 132.6000 1430.7001 ;
	    RECT 130.5000 1429.5000 139.8000 1429.8000 ;
	    RECT 131.7000 1428.9000 139.8000 1429.5000 ;
	    RECT 138.6000 1428.6000 139.8000 1428.9000 ;
	    RECT 141.3000 1429.5000 142.2000 1430.7001 ;
	    RECT 143.1000 1430.4000 147.0000 1431.6000 ;
	    RECT 150.6000 1430.4000 151.8000 1439.7001 ;
	    RECT 153.0000 1435.5000 154.2000 1439.7001 ;
	    RECT 155.4000 1435.5000 156.6000 1439.7001 ;
	    RECT 157.8000 1435.5000 159.0000 1439.7001 ;
	    RECT 160.2000 1433.7001 161.4000 1439.7001 ;
	    RECT 155.4000 1431.6000 161.7000 1432.8000 ;
	    RECT 162.6000 1431.6000 163.8000 1439.7001 ;
	    RECT 165.0000 1433.7001 166.2000 1439.7001 ;
	    RECT 167.4000 1432.8000 168.6000 1439.7001 ;
	    RECT 169.8000 1433.7001 171.0000 1439.7001 ;
	    RECT 167.4000 1431.9000 171.3000 1432.8000 ;
	    RECT 172.2000 1432.5000 173.4000 1439.7001 ;
	    RECT 174.6000 1433.7001 175.8000 1439.7001 ;
	    RECT 306.6000 1433.7001 307.8000 1439.7001 ;
	    RECT 309.0000 1432.5000 310.2000 1439.7001 ;
	    RECT 311.4000 1433.7001 312.6000 1439.7001 ;
	    RECT 313.8000 1432.8000 315.0000 1439.7001 ;
	    RECT 316.2000 1433.7001 317.4000 1439.7001 ;
	    RECT 162.6000 1430.4000 166.5000 1431.6000 ;
	    RECT 153.0000 1429.5000 154.2000 1429.8000 ;
	    RECT 141.3000 1428.6000 154.2000 1429.5000 ;
	    RECT 157.8000 1429.5000 159.0000 1429.8000 ;
	    RECT 170.4000 1429.5000 171.3000 1431.9000 ;
	    RECT 311.1000 1431.9000 315.0000 1432.8000 ;
	    RECT 172.2000 1430.4000 173.4000 1431.6000 ;
	    RECT 237.0000 1431.4501 238.2000 1431.6000 ;
	    RECT 268.2000 1431.4501 269.4000 1431.6000 ;
	    RECT 280.2000 1431.4501 281.4000 1431.6000 ;
	    RECT 309.0000 1431.4501 310.2000 1431.6000 ;
	    RECT 237.0000 1430.5500 310.2000 1431.4501 ;
	    RECT 237.0000 1430.4000 238.2000 1430.5500 ;
	    RECT 268.2000 1430.4000 269.4000 1430.5500 ;
	    RECT 280.2000 1430.4000 281.4000 1430.5500 ;
	    RECT 309.0000 1430.4000 310.2000 1430.5500 ;
	    RECT 311.1000 1429.5000 312.0000 1431.9000 ;
	    RECT 318.6000 1431.6000 319.8000 1439.7001 ;
	    RECT 321.0000 1433.7001 322.2000 1439.7001 ;
	    RECT 323.4000 1435.5000 324.6000 1439.7001 ;
	    RECT 325.8000 1435.5000 327.0000 1439.7001 ;
	    RECT 328.2000 1435.5000 329.4000 1439.7001 ;
	    RECT 320.7000 1431.6000 327.0000 1432.8000 ;
	    RECT 315.9000 1430.4000 319.8000 1431.6000 ;
	    RECT 330.6000 1430.4000 331.8000 1439.7001 ;
	    RECT 333.0000 1433.7001 334.2000 1439.7001 ;
	    RECT 335.4000 1432.5000 336.6000 1439.7001 ;
	    RECT 337.8000 1433.7001 339.0000 1439.7001 ;
	    RECT 340.2000 1432.5000 341.4000 1439.7001 ;
	    RECT 342.6000 1435.5000 343.8000 1439.7001 ;
	    RECT 345.0000 1435.5000 346.2000 1439.7001 ;
	    RECT 347.4000 1433.7001 348.6000 1439.7001 ;
	    RECT 349.8000 1432.8000 351.0000 1439.7001 ;
	    RECT 352.2000 1433.7001 353.4000 1440.6000 ;
	    RECT 354.6000 1434.6000 355.8000 1439.7001 ;
	    RECT 354.6000 1433.7001 356.1000 1434.6000 ;
	    RECT 357.0000 1433.7001 358.2000 1439.7001 ;
	    RECT 376.2000 1433.7001 377.4000 1439.7001 ;
	    RECT 355.2000 1432.8000 356.1000 1433.7001 ;
	    RECT 348.0000 1431.6000 354.3000 1432.8000 ;
	    RECT 355.2000 1431.9000 358.2000 1432.8000 ;
	    RECT 335.4000 1430.4000 339.3000 1431.6000 ;
	    RECT 340.2000 1430.7001 348.9000 1431.6000 ;
	    RECT 353.4000 1431.0000 354.3000 1431.6000 ;
	    RECT 323.4000 1429.5000 324.6000 1429.8000 ;
	    RECT 157.8000 1428.6000 171.3000 1429.5000 ;
	    RECT 129.0000 1427.4000 130.2000 1428.6000 ;
	    RECT 134.1000 1427.7001 135.3000 1428.0000 ;
	    RECT 131.1000 1426.8000 169.5000 1427.7001 ;
	    RECT 168.3000 1426.5000 169.5000 1426.8000 ;
	    RECT 170.4000 1425.9000 171.3000 1428.6000 ;
	    RECT 172.2000 1428.0000 173.4000 1429.5000 ;
	    RECT 309.0000 1428.0000 310.2000 1429.5000 ;
	    RECT 172.2000 1426.8000 173.7000 1428.0000 ;
	    RECT 126.3000 1425.0000 132.9000 1425.9000 ;
	    RECT 126.3000 1424.7001 127.5000 1425.0000 ;
	    RECT 133.8000 1424.4000 135.0000 1425.6000 ;
	    RECT 135.9000 1425.0000 161.4000 1425.9000 ;
	    RECT 170.4000 1425.0000 171.6000 1425.9000 ;
	    RECT 160.2000 1424.1000 161.4000 1425.0000 ;
	    RECT 124.2000 1422.3000 137.4000 1423.5000 ;
	    RECT 138.3000 1422.9000 141.3000 1424.1000 ;
	    RECT 147.0000 1422.9000 151.8000 1424.1000 ;
	    RECT 124.2000 1413.3000 125.4000 1422.3000 ;
	    RECT 127.8000 1420.2001 132.3000 1421.4000 ;
	    RECT 131.1000 1419.3000 132.3000 1420.2001 ;
	    RECT 140.1000 1419.3000 141.3000 1422.9000 ;
	    RECT 143.4000 1421.4000 144.6000 1422.6000 ;
	    RECT 151.2000 1421.7001 152.4000 1422.0000 ;
	    RECT 145.8000 1420.8000 152.4000 1421.7001 ;
	    RECT 145.8000 1420.5000 147.0000 1420.8000 ;
	    RECT 143.4000 1420.2001 144.6000 1420.5000 ;
	    RECT 155.4000 1419.6000 156.6000 1423.8000 ;
	    RECT 164.1000 1422.9000 169.8000 1424.1000 ;
	    RECT 164.1000 1421.1000 165.3000 1422.9000 ;
	    RECT 170.7000 1422.0000 171.6000 1425.0000 ;
	    RECT 145.8000 1419.3000 147.0000 1419.6000 ;
	    RECT 129.0000 1413.3000 130.2000 1419.3000 ;
	    RECT 131.1000 1418.1000 135.0000 1419.3000 ;
	    RECT 140.1000 1418.4000 147.0000 1419.3000 ;
	    RECT 148.2000 1418.4000 149.4000 1419.6000 ;
	    RECT 150.3000 1418.4000 150.6000 1419.6000 ;
	    RECT 155.1000 1418.4000 156.6000 1419.6000 ;
	    RECT 162.6000 1420.2001 165.3000 1421.1000 ;
	    RECT 169.8000 1421.1000 171.6000 1422.0000 ;
	    RECT 162.6000 1419.3000 163.8000 1420.2001 ;
	    RECT 133.8000 1413.3000 135.0000 1418.1000 ;
	    RECT 160.2000 1418.1000 163.8000 1419.3000 ;
	    RECT 136.2000 1413.3000 137.4000 1417.5000 ;
	    RECT 138.6000 1413.3000 139.8000 1417.5000 ;
	    RECT 141.0000 1413.3000 142.2000 1417.5000 ;
	    RECT 143.4000 1413.3000 144.6000 1416.3000 ;
	    RECT 145.8000 1413.3000 147.0000 1417.5000 ;
	    RECT 148.2000 1413.3000 149.4000 1416.3000 ;
	    RECT 150.6000 1413.3000 151.8000 1417.5000 ;
	    RECT 153.0000 1413.3000 154.2000 1417.5000 ;
	    RECT 155.4000 1413.3000 156.6000 1417.5000 ;
	    RECT 157.8000 1413.3000 159.0000 1417.5000 ;
	    RECT 160.2000 1413.3000 161.4000 1418.1000 ;
	    RECT 165.0000 1413.3000 166.2000 1419.3000 ;
	    RECT 169.8000 1413.3000 171.0000 1421.1000 ;
	    RECT 172.5000 1420.2001 173.7000 1426.8000 ;
	    RECT 172.2000 1419.0000 173.7000 1420.2001 ;
	    RECT 308.7000 1426.8000 310.2000 1428.0000 ;
	    RECT 311.1000 1428.6000 324.6000 1429.5000 ;
	    RECT 328.2000 1429.5000 329.4000 1429.8000 ;
	    RECT 340.2000 1429.5000 341.1000 1430.7001 ;
	    RECT 349.8000 1429.8000 351.9000 1430.7001 ;
	    RECT 353.4000 1429.8000 355.8000 1431.0000 ;
	    RECT 328.2000 1428.6000 341.1000 1429.5000 ;
	    RECT 342.6000 1429.5000 351.9000 1429.8000 ;
	    RECT 342.6000 1428.9000 350.7000 1429.5000 ;
	    RECT 342.6000 1428.6000 343.8000 1428.9000 ;
	    RECT 308.7000 1420.2001 309.9000 1426.8000 ;
	    RECT 311.1000 1425.9000 312.0000 1428.6000 ;
	    RECT 347.1000 1427.7001 348.3000 1428.0000 ;
	    RECT 312.9000 1426.8000 351.3000 1427.7001 ;
	    RECT 352.2000 1427.4000 353.4000 1428.6000 ;
	    RECT 312.9000 1426.5000 314.1000 1426.8000 ;
	    RECT 310.8000 1425.0000 312.0000 1425.9000 ;
	    RECT 321.0000 1425.0000 346.5000 1425.9000 ;
	    RECT 310.8000 1422.0000 311.7000 1425.0000 ;
	    RECT 321.0000 1424.1000 322.2000 1425.0000 ;
	    RECT 347.4000 1424.4000 348.6000 1425.6000 ;
	    RECT 349.5000 1425.0000 356.1000 1425.9000 ;
	    RECT 354.9000 1424.7001 356.1000 1425.0000 ;
	    RECT 312.6000 1422.9000 318.3000 1424.1000 ;
	    RECT 310.8000 1421.1000 312.6000 1422.0000 ;
	    RECT 308.7000 1419.0000 310.2000 1420.2001 ;
	    RECT 172.2000 1413.3000 173.4000 1419.0000 ;
	    RECT 174.6000 1413.3000 175.8000 1416.3000 ;
	    RECT 306.6000 1413.3000 307.8000 1416.3000 ;
	    RECT 309.0000 1413.3000 310.2000 1419.0000 ;
	    RECT 311.4000 1413.3000 312.6000 1421.1000 ;
	    RECT 317.1000 1421.1000 318.3000 1422.9000 ;
	    RECT 317.1000 1420.2001 319.8000 1421.1000 ;
	    RECT 318.6000 1419.3000 319.8000 1420.2001 ;
	    RECT 325.8000 1419.6000 327.0000 1423.8000 ;
	    RECT 330.6000 1422.9000 335.4000 1424.1000 ;
	    RECT 341.1000 1422.9000 344.1000 1424.1000 ;
	    RECT 357.0000 1423.5000 358.2000 1431.9000 ;
	    RECT 376.2000 1429.5000 377.4000 1429.8000 ;
	    RECT 376.2000 1427.4000 377.4000 1428.6000 ;
	    RECT 378.6000 1426.5000 379.8000 1439.7001 ;
	    RECT 381.0000 1433.7001 382.2000 1439.7001 ;
	    RECT 408.3000 1433.7001 409.5000 1439.7001 ;
	    RECT 408.6000 1430.4000 409.8000 1431.6000 ;
	    RECT 408.6000 1429.5000 409.5000 1430.4000 ;
	    RECT 410.7000 1428.6000 411.9000 1439.7001 ;
	    RECT 407.4000 1427.4000 408.6000 1428.6000 ;
	    RECT 410.4000 1427.7001 411.9000 1428.6000 ;
	    RECT 414.6000 1427.7001 415.8000 1439.7001 ;
	    RECT 426.6000 1433.7001 427.8000 1439.7001 ;
	    RECT 378.6000 1425.4501 379.8000 1425.6000 ;
	    RECT 407.5500 1425.4501 408.4500 1427.4000 ;
	    RECT 378.6000 1424.5500 408.4500 1425.4501 ;
	    RECT 378.6000 1424.4000 379.8000 1424.5500 ;
	    RECT 330.0000 1421.7001 331.2000 1422.0000 ;
	    RECT 330.0000 1420.8000 336.6000 1421.7001 ;
	    RECT 337.8000 1421.4000 339.0000 1422.6000 ;
	    RECT 335.4000 1420.5000 336.6000 1420.8000 ;
	    RECT 337.8000 1420.2001 339.0000 1420.5000 ;
	    RECT 316.2000 1413.3000 317.4000 1419.3000 ;
	    RECT 318.6000 1418.1000 322.2000 1419.3000 ;
	    RECT 325.8000 1418.4000 327.3000 1419.6000 ;
	    RECT 331.8000 1418.4000 332.1000 1419.6000 ;
	    RECT 333.0000 1418.4000 334.2000 1419.6000 ;
	    RECT 335.4000 1419.3000 336.6000 1419.6000 ;
	    RECT 341.1000 1419.3000 342.3000 1422.9000 ;
	    RECT 345.0000 1422.3000 358.2000 1423.5000 ;
	    RECT 350.1000 1420.2001 354.6000 1421.4000 ;
	    RECT 350.1000 1419.3000 351.3000 1420.2001 ;
	    RECT 335.4000 1418.4000 342.3000 1419.3000 ;
	    RECT 321.0000 1413.3000 322.2000 1418.1000 ;
	    RECT 347.4000 1418.1000 351.3000 1419.3000 ;
	    RECT 323.4000 1413.3000 324.6000 1417.5000 ;
	    RECT 325.8000 1413.3000 327.0000 1417.5000 ;
	    RECT 328.2000 1413.3000 329.4000 1417.5000 ;
	    RECT 330.6000 1413.3000 331.8000 1417.5000 ;
	    RECT 333.0000 1413.3000 334.2000 1416.3000 ;
	    RECT 335.4000 1413.3000 336.6000 1417.5000 ;
	    RECT 337.8000 1413.3000 339.0000 1416.3000 ;
	    RECT 340.2000 1413.3000 341.4000 1417.5000 ;
	    RECT 342.6000 1413.3000 343.8000 1417.5000 ;
	    RECT 345.0000 1413.3000 346.2000 1417.5000 ;
	    RECT 347.4000 1413.3000 348.6000 1418.1000 ;
	    RECT 352.2000 1413.3000 353.4000 1419.3000 ;
	    RECT 357.0000 1413.3000 358.2000 1422.3000 ;
	    RECT 378.6000 1419.3000 379.8000 1423.5000 ;
	    RECT 410.4000 1422.6000 411.3000 1427.7001 ;
	    RECT 412.2000 1425.4501 413.4000 1425.6000 ;
	    RECT 412.2000 1424.5500 418.0500 1425.4501 ;
	    RECT 412.2000 1424.4000 413.4000 1424.5500 ;
	    RECT 412.2000 1423.2001 413.4000 1423.5000 ;
	    RECT 381.0000 1422.4501 382.2000 1422.6000 ;
	    RECT 385.8000 1422.4501 387.0000 1422.6000 ;
	    RECT 381.0000 1421.5500 387.0000 1422.4501 ;
	    RECT 381.0000 1421.4000 382.2000 1421.5500 ;
	    RECT 385.8000 1421.4000 387.0000 1421.5500 ;
	    RECT 407.4000 1421.4000 408.6000 1422.6000 ;
	    RECT 409.5000 1421.4000 411.3000 1422.6000 ;
	    RECT 413.4000 1420.8000 413.7000 1422.3000 ;
	    RECT 414.6000 1421.4000 415.8000 1422.6000 ;
	    RECT 417.1500 1422.4501 418.0500 1424.5500 ;
	    RECT 429.0000 1423.5000 430.2000 1439.7001 ;
	    RECT 460.2000 1427.7001 461.4000 1439.7001 ;
	    RECT 464.1000 1428.6000 465.3000 1439.7001 ;
	    RECT 466.5000 1433.7001 467.7000 1439.7001 ;
	    RECT 486.6000 1433.7001 487.8000 1439.7001 ;
	    RECT 466.2000 1430.4000 467.4000 1431.6000 ;
	    RECT 466.5000 1429.5000 467.4000 1430.4000 ;
	    RECT 464.1000 1427.7001 465.6000 1428.6000 ;
	    RECT 457.8000 1425.4501 459.0000 1425.6000 ;
	    RECT 462.6000 1425.4501 463.8000 1425.6000 ;
	    RECT 457.8000 1424.5500 463.8000 1425.4501 ;
	    RECT 457.8000 1424.4000 459.0000 1424.5500 ;
	    RECT 462.6000 1424.4000 463.8000 1424.5500 ;
	    RECT 462.6000 1423.2001 463.8000 1423.5000 ;
	    RECT 464.7000 1422.6000 465.6000 1427.7001 ;
	    RECT 467.4000 1427.4000 468.6000 1428.6000 ;
	    RECT 467.5500 1425.4501 468.4500 1427.4000 ;
	    RECT 489.0000 1426.5000 490.2000 1439.7001 ;
	    RECT 491.4000 1433.7001 492.6000 1439.7001 ;
	    RECT 508.2000 1439.4000 509.4000 1440.6000 ;
	    RECT 541.8000 1439.4000 543.0000 1440.6000 ;
	    RECT 491.4000 1429.5000 492.6000 1429.8000 ;
	    RECT 491.4000 1427.4000 492.6000 1428.6000 ;
	    RECT 561.0000 1426.8000 562.2000 1439.7001 ;
	    RECT 563.4000 1427.7001 564.6000 1439.7001 ;
	    RECT 567.3000 1433.7001 569.1000 1439.7001 ;
	    RECT 571.8000 1433.7001 573.0000 1439.7001 ;
	    RECT 574.2000 1433.7001 575.4000 1439.7001 ;
	    RECT 576.6000 1433.7001 577.8000 1439.7001 ;
	    RECT 580.8000 1434.6000 582.0000 1439.7001 ;
	    RECT 580.8000 1433.7001 583.8000 1434.6000 ;
	    RECT 568.2000 1432.5000 569.4000 1433.7001 ;
	    RECT 574.5000 1432.8000 575.4000 1433.7001 ;
	    RECT 573.3000 1431.9000 578.7000 1432.8000 ;
	    RECT 582.6000 1432.5000 583.8000 1433.7001 ;
	    RECT 573.3000 1431.6000 574.5000 1431.9000 ;
	    RECT 577.5000 1431.6000 578.7000 1431.9000 ;
	    RECT 567.0000 1429.8000 569.1000 1431.0000 ;
	    RECT 568.2000 1428.3000 569.1000 1429.8000 ;
	    RECT 571.5000 1429.5000 574.8000 1430.4000 ;
	    RECT 571.5000 1429.2001 572.7000 1429.5000 ;
	    RECT 568.2000 1427.4000 571.8000 1428.3000 ;
	    RECT 561.0000 1426.5000 567.3000 1426.8000 ;
	    RECT 563.1000 1425.9000 567.3000 1426.5000 ;
	    RECT 566.1000 1425.6000 567.3000 1425.9000 ;
	    RECT 489.0000 1425.4501 490.2000 1425.6000 ;
	    RECT 467.5500 1424.5500 490.2000 1425.4501 ;
	    RECT 489.0000 1424.4000 490.2000 1424.5500 ;
	    RECT 561.0000 1424.4000 562.2000 1425.6000 ;
	    RECT 563.7000 1424.7001 564.9000 1425.0000 ;
	    RECT 563.7000 1423.8000 569.4000 1424.7001 ;
	    RECT 568.2000 1423.5000 569.4000 1423.8000 ;
	    RECT 429.0000 1422.4501 430.2000 1422.6000 ;
	    RECT 417.1500 1421.5500 430.2000 1422.4501 ;
	    RECT 429.0000 1421.4000 430.2000 1421.5500 ;
	    RECT 460.2000 1421.4000 461.4000 1422.6000 ;
	    RECT 462.3000 1420.8000 462.6000 1422.3000 ;
	    RECT 464.7000 1421.4000 466.5000 1422.6000 ;
	    RECT 467.4000 1422.4501 468.6000 1422.6000 ;
	    RECT 472.2000 1422.4501 473.4000 1422.6000 ;
	    RECT 467.4000 1421.5500 473.4000 1422.4501 ;
	    RECT 467.4000 1421.4000 468.6000 1421.5500 ;
	    RECT 472.2000 1421.4000 473.4000 1421.5500 ;
	    RECT 474.6000 1422.4501 475.8000 1422.6000 ;
	    RECT 479.4000 1422.4501 480.6000 1422.6000 ;
	    RECT 486.6000 1422.4501 487.8000 1422.6000 ;
	    RECT 474.6000 1421.5500 487.8000 1422.4501 ;
	    RECT 474.6000 1421.4000 475.8000 1421.5500 ;
	    RECT 479.4000 1421.4000 480.6000 1421.5500 ;
	    RECT 486.6000 1421.4000 487.8000 1421.5500 ;
	    RECT 381.0000 1420.2001 382.2000 1420.5000 ;
	    RECT 407.7000 1419.3000 408.6000 1420.5000 ;
	    RECT 410.1000 1419.3000 415.5000 1419.9000 ;
	    RECT 377.1000 1418.4000 379.8000 1419.3000 ;
	    RECT 377.1000 1413.3000 378.3000 1418.4000 ;
	    RECT 381.0000 1413.3000 382.2000 1419.3000 ;
	    RECT 407.4000 1413.3000 408.6000 1419.3000 ;
	    RECT 409.8000 1419.0000 415.8000 1419.3000 ;
	    RECT 409.8000 1413.3000 411.0000 1419.0000 ;
	    RECT 412.2000 1413.3000 413.4000 1418.1000 ;
	    RECT 414.6000 1413.3000 415.8000 1419.0000 ;
	    RECT 426.6000 1418.4000 427.8000 1419.6000 ;
	    RECT 426.6000 1417.2001 427.8000 1417.5000 ;
	    RECT 426.6000 1413.3000 427.8000 1416.3000 ;
	    RECT 429.0000 1413.3000 430.2000 1420.5000 ;
	    RECT 460.5000 1419.3000 465.9000 1419.9000 ;
	    RECT 467.4000 1419.3000 468.3000 1420.5000 ;
	    RECT 486.6000 1420.2001 487.8000 1420.5000 ;
	    RECT 489.0000 1419.3000 490.2000 1423.5000 ;
	    RECT 561.0000 1420.8000 562.2000 1423.5000 ;
	    RECT 570.9000 1422.6000 571.8000 1427.4000 ;
	    RECT 573.9000 1427.7001 574.8000 1429.5000 ;
	    RECT 575.7000 1429.5000 576.9000 1429.8000 ;
	    RECT 582.6000 1429.5000 583.8000 1429.8000 ;
	    RECT 575.7000 1428.6000 583.8000 1429.5000 ;
	    RECT 585.0000 1428.0000 586.2000 1439.7001 ;
	    RECT 573.9000 1427.1000 581.1000 1427.7001 ;
	    RECT 587.4000 1427.1000 588.6000 1439.7001 ;
	    RECT 606.6000 1427.7001 607.8000 1439.7001 ;
	    RECT 610.5000 1428.9000 611.7000 1439.7001 ;
	    RECT 609.0000 1427.7001 611.7000 1428.9000 ;
	    RECT 573.9000 1426.8000 588.6000 1427.1000 ;
	    RECT 579.9000 1426.5000 588.6000 1426.8000 ;
	    RECT 580.2000 1426.2001 588.6000 1426.5000 ;
	    RECT 577.8000 1424.4000 579.0000 1425.6000 ;
	    RECT 579.9000 1424.4000 585.3000 1425.3000 ;
	    RECT 584.1000 1424.1000 585.3000 1424.4000 ;
	    RECT 609.3000 1423.5000 610.2000 1427.7001 ;
	    RECT 611.4000 1426.5000 612.6000 1426.8000 ;
	    RECT 611.4000 1425.4501 612.6000 1425.6000 ;
	    RECT 613.8000 1425.4501 615.0000 1425.6000 ;
	    RECT 611.4000 1424.5500 615.0000 1425.4501 ;
	    RECT 611.4000 1424.4000 612.6000 1424.5500 ;
	    RECT 613.8000 1424.4000 615.0000 1424.5500 ;
	    RECT 623.4000 1423.5000 624.6000 1439.7001 ;
	    RECT 625.8000 1433.7001 627.0000 1439.7001 ;
	    RECT 650.7000 1433.7001 651.9000 1439.7001 ;
	    RECT 651.0000 1430.4000 652.2000 1431.6000 ;
	    RECT 651.0000 1429.5000 651.9000 1430.4000 ;
	    RECT 653.1000 1428.6000 654.3000 1439.7001 ;
	    RECT 649.8000 1427.4000 651.0000 1428.6000 ;
	    RECT 652.8000 1427.7001 654.3000 1428.6000 ;
	    RECT 657.0000 1427.7001 658.2000 1439.7001 ;
	    RECT 659.4000 1428.4501 660.6000 1428.6000 ;
	    RECT 676.2000 1428.4501 677.4000 1428.6000 ;
	    RECT 581.7000 1422.6000 582.9000 1422.9000 ;
	    RECT 652.8000 1422.6000 653.7000 1427.7001 ;
	    RECT 659.4000 1427.5500 677.4000 1428.4501 ;
	    RECT 659.4000 1427.4000 660.6000 1427.5500 ;
	    RECT 676.2000 1427.4000 677.4000 1427.5500 ;
	    RECT 654.6000 1425.4501 655.8000 1425.6000 ;
	    RECT 654.6000 1424.5500 660.4500 1425.4501 ;
	    RECT 654.6000 1424.4000 655.8000 1424.5500 ;
	    RECT 654.6000 1423.2001 655.8000 1423.5000 ;
	    RECT 570.9000 1421.7001 584.1000 1422.6000 ;
	    RECT 571.5000 1421.4000 572.7000 1421.7001 ;
	    RECT 561.0000 1419.9000 566.7000 1420.8000 ;
	    RECT 460.2000 1419.0000 466.2000 1419.3000 ;
	    RECT 460.2000 1413.3000 461.4000 1419.0000 ;
	    RECT 462.6000 1413.3000 463.8000 1418.1000 ;
	    RECT 465.0000 1413.3000 466.2000 1419.0000 ;
	    RECT 467.4000 1413.3000 468.6000 1419.3000 ;
	    RECT 486.6000 1413.3000 487.8000 1419.3000 ;
	    RECT 489.0000 1418.4000 491.7000 1419.3000 ;
	    RECT 490.5000 1413.3000 491.7000 1418.4000 ;
	    RECT 561.0000 1413.3000 562.2000 1419.9000 ;
	    RECT 565.5000 1419.6000 566.7000 1419.9000 ;
	    RECT 563.4000 1413.3000 564.6000 1419.0000 ;
	    RECT 580.2000 1418.4000 581.1000 1421.7001 ;
	    RECT 585.0000 1421.4000 586.2000 1422.6000 ;
	    RECT 587.1000 1421.4000 587.4000 1422.6000 ;
	    RECT 589.8000 1422.4501 591.0000 1422.6000 ;
	    RECT 609.0000 1422.4501 610.2000 1422.6000 ;
	    RECT 589.8000 1421.5500 610.2000 1422.4501 ;
	    RECT 589.8000 1421.4000 591.0000 1421.5500 ;
	    RECT 609.0000 1421.4000 610.2000 1421.5500 ;
	    RECT 611.4000 1422.4501 612.6000 1422.6000 ;
	    RECT 623.4000 1422.4501 624.6000 1422.6000 ;
	    RECT 611.4000 1421.5500 624.6000 1422.4501 ;
	    RECT 611.4000 1421.4000 612.6000 1421.5500 ;
	    RECT 623.4000 1421.4000 624.6000 1421.5500 ;
	    RECT 649.8000 1421.4000 651.0000 1422.6000 ;
	    RECT 651.9000 1421.4000 653.7000 1422.6000 ;
	    RECT 655.8000 1420.8000 656.1000 1422.3000 ;
	    RECT 657.0000 1421.4000 658.2000 1422.6000 ;
	    RECT 659.5500 1422.4501 660.4500 1424.5500 ;
	    RECT 678.6000 1423.5000 679.8000 1439.7001 ;
	    RECT 681.0000 1433.7001 682.2000 1439.7001 ;
	    RECT 700.2000 1433.7001 701.4000 1439.7001 ;
	    RECT 702.6000 1426.5000 703.8000 1439.7001 ;
	    RECT 705.0000 1433.7001 706.2000 1439.7001 ;
	    RECT 829.8000 1433.7001 831.0000 1439.7001 ;
	    RECT 832.2000 1434.6000 833.4000 1439.7001 ;
	    RECT 831.9000 1433.7001 833.4000 1434.6000 ;
	    RECT 834.6000 1433.7001 835.8000 1440.6000 ;
	    RECT 831.9000 1432.8000 832.8000 1433.7001 ;
	    RECT 837.0000 1432.8000 838.2000 1439.7001 ;
	    RECT 839.4000 1433.7001 840.6000 1439.7001 ;
	    RECT 841.8000 1435.5000 843.0000 1439.7001 ;
	    RECT 844.2000 1435.5000 845.4000 1439.7001 ;
	    RECT 829.8000 1431.9000 832.8000 1432.8000 ;
	    RECT 705.0000 1429.5000 706.2000 1429.8000 ;
	    RECT 705.0000 1428.4501 706.2000 1428.6000 ;
	    RECT 762.6000 1428.4501 763.8000 1428.6000 ;
	    RECT 705.0000 1427.5500 763.8000 1428.4501 ;
	    RECT 705.0000 1427.4000 706.2000 1427.5500 ;
	    RECT 762.6000 1427.4000 763.8000 1427.5500 ;
	    RECT 681.0000 1425.4501 682.2000 1425.6000 ;
	    RECT 702.6000 1425.4501 703.8000 1425.6000 ;
	    RECT 681.0000 1424.5500 703.8000 1425.4501 ;
	    RECT 681.0000 1424.4000 682.2000 1424.5500 ;
	    RECT 702.6000 1424.4000 703.8000 1424.5500 ;
	    RECT 829.8000 1423.5000 831.0000 1431.9000 ;
	    RECT 833.7000 1431.6000 840.0000 1432.8000 ;
	    RECT 846.6000 1432.5000 847.8000 1439.7001 ;
	    RECT 849.0000 1433.7001 850.2000 1439.7001 ;
	    RECT 851.4000 1432.5000 852.6000 1439.7001 ;
	    RECT 853.8000 1433.7001 855.0000 1439.7001 ;
	    RECT 833.7000 1431.0000 834.6000 1431.6000 ;
	    RECT 832.2000 1429.8000 834.6000 1431.0000 ;
	    RECT 839.1000 1430.7001 847.8000 1431.6000 ;
	    RECT 836.1000 1429.8000 838.2000 1430.7001 ;
	    RECT 836.1000 1429.5000 845.4000 1429.8000 ;
	    RECT 837.3000 1428.9000 845.4000 1429.5000 ;
	    RECT 844.2000 1428.6000 845.4000 1428.9000 ;
	    RECT 846.9000 1429.5000 847.8000 1430.7001 ;
	    RECT 848.7000 1430.4000 852.6000 1431.6000 ;
	    RECT 856.2000 1430.4000 857.4000 1439.7001 ;
	    RECT 858.6000 1435.5000 859.8000 1439.7001 ;
	    RECT 861.0000 1435.5000 862.2000 1439.7001 ;
	    RECT 863.4000 1435.5000 864.6000 1439.7001 ;
	    RECT 865.8000 1433.7001 867.0000 1439.7001 ;
	    RECT 861.0000 1431.6000 867.3000 1432.8000 ;
	    RECT 868.2000 1431.6000 869.4000 1439.7001 ;
	    RECT 870.6000 1433.7001 871.8000 1439.7001 ;
	    RECT 873.0000 1432.8000 874.2000 1439.7001 ;
	    RECT 875.4000 1433.7001 876.6000 1439.7001 ;
	    RECT 873.0000 1431.9000 876.9000 1432.8000 ;
	    RECT 877.8000 1432.5000 879.0000 1439.7001 ;
	    RECT 880.2000 1433.7001 881.4000 1439.7001 ;
	    RECT 901.8000 1433.7001 903.0000 1439.7001 ;
	    RECT 868.2000 1430.4000 872.1000 1431.6000 ;
	    RECT 858.6000 1429.5000 859.8000 1429.8000 ;
	    RECT 846.9000 1428.6000 859.8000 1429.5000 ;
	    RECT 863.4000 1429.5000 864.6000 1429.8000 ;
	    RECT 876.0000 1429.5000 876.9000 1431.9000 ;
	    RECT 877.8000 1430.4000 879.0000 1431.6000 ;
	    RECT 863.4000 1428.6000 876.9000 1429.5000 ;
	    RECT 834.6000 1427.4000 835.8000 1428.6000 ;
	    RECT 839.7000 1427.7001 840.9000 1428.0000 ;
	    RECT 836.7000 1426.8000 875.1000 1427.7001 ;
	    RECT 873.9000 1426.5000 875.1000 1426.8000 ;
	    RECT 876.0000 1425.9000 876.9000 1428.6000 ;
	    RECT 877.8000 1428.0000 879.0000 1429.5000 ;
	    RECT 877.8000 1426.8000 879.3000 1428.0000 ;
	    RECT 831.9000 1425.0000 838.5000 1425.9000 ;
	    RECT 831.9000 1424.7001 833.1000 1425.0000 ;
	    RECT 839.4000 1424.4000 840.6000 1425.6000 ;
	    RECT 841.5000 1425.0000 867.0000 1425.9000 ;
	    RECT 876.0000 1425.0000 877.2000 1425.9000 ;
	    RECT 865.8000 1424.1000 867.0000 1425.0000 ;
	    RECT 678.6000 1422.4501 679.8000 1422.6000 ;
	    RECT 659.5500 1421.5500 679.8000 1422.4501 ;
	    RECT 678.6000 1421.4000 679.8000 1421.5500 ;
	    RECT 683.4000 1422.4501 684.6000 1422.6000 ;
	    RECT 700.2000 1422.4501 701.4000 1422.6000 ;
	    RECT 683.4000 1421.5500 701.4000 1422.4501 ;
	    RECT 683.4000 1421.4000 684.6000 1421.5500 ;
	    RECT 700.2000 1421.4000 701.4000 1421.5500 ;
	    RECT 577.5000 1418.1000 578.7000 1418.4000 ;
	    RECT 568.2000 1416.3000 569.4000 1417.5000 ;
	    RECT 574.5000 1417.2001 578.7000 1418.1000 ;
	    RECT 580.2000 1417.2001 581.4000 1418.4000 ;
	    RECT 574.5000 1416.3000 575.4000 1417.2001 ;
	    RECT 582.6000 1416.3000 583.8000 1417.5000 ;
	    RECT 567.3000 1415.4000 569.4000 1416.3000 ;
	    RECT 567.3000 1413.3000 569.1000 1415.4000 ;
	    RECT 571.8000 1413.3000 573.0000 1416.3000 ;
	    RECT 574.2000 1413.3000 575.4000 1416.3000 ;
	    RECT 576.6000 1413.3000 578.1000 1416.3000 ;
	    RECT 580.8000 1415.4000 583.8000 1416.3000 ;
	    RECT 580.8000 1413.3000 582.0000 1415.4000 ;
	    RECT 585.0000 1413.3000 586.2000 1419.3000 ;
	    RECT 587.4000 1413.3000 588.6000 1420.5000 ;
	    RECT 606.6000 1418.4000 607.8000 1419.6000 ;
	    RECT 606.6000 1417.2001 607.8000 1417.5000 ;
	    RECT 609.3000 1416.3000 610.2000 1420.5000 ;
	    RECT 606.6000 1413.3000 607.8000 1416.3000 ;
	    RECT 609.0000 1413.3000 610.2000 1416.3000 ;
	    RECT 611.4000 1413.3000 612.6000 1416.3000 ;
	    RECT 623.4000 1413.3000 624.6000 1420.5000 ;
	    RECT 625.8000 1419.4501 627.0000 1419.6000 ;
	    RECT 647.4000 1419.4501 648.6000 1419.6000 ;
	    RECT 625.8000 1418.5500 648.6000 1419.4501 ;
	    RECT 650.1000 1419.3000 651.0000 1420.5000 ;
	    RECT 652.5000 1419.3000 657.9000 1419.9000 ;
	    RECT 625.8000 1418.4000 627.0000 1418.5500 ;
	    RECT 647.4000 1418.4000 648.6000 1418.5500 ;
	    RECT 625.8000 1417.2001 627.0000 1417.5000 ;
	    RECT 625.8000 1413.3000 627.0000 1416.3000 ;
	    RECT 649.8000 1413.3000 651.0000 1419.3000 ;
	    RECT 652.2000 1419.0000 658.2000 1419.3000 ;
	    RECT 652.2000 1413.3000 653.4000 1419.0000 ;
	    RECT 654.6000 1413.3000 655.8000 1418.1000 ;
	    RECT 657.0000 1413.3000 658.2000 1419.0000 ;
	    RECT 678.6000 1413.3000 679.8000 1420.5000 ;
	    RECT 700.2000 1420.2001 701.4000 1420.5000 ;
	    RECT 681.0000 1419.4501 682.2000 1419.6000 ;
	    RECT 697.8000 1419.4501 699.0000 1419.6000 ;
	    RECT 681.0000 1418.5500 699.0000 1419.4501 ;
	    RECT 702.6000 1419.3000 703.8000 1423.5000 ;
	    RECT 829.8000 1422.3000 843.0000 1423.5000 ;
	    RECT 843.9000 1422.9000 846.9000 1424.1000 ;
	    RECT 852.6000 1422.9000 857.4000 1424.1000 ;
	    RECT 681.0000 1418.4000 682.2000 1418.5500 ;
	    RECT 697.8000 1418.4000 699.0000 1418.5500 ;
	    RECT 681.0000 1417.2001 682.2000 1417.5000 ;
	    RECT 681.0000 1413.3000 682.2000 1416.3000 ;
	    RECT 700.2000 1413.3000 701.4000 1419.3000 ;
	    RECT 702.6000 1418.4000 705.3000 1419.3000 ;
	    RECT 704.1000 1413.3000 705.3000 1418.4000 ;
	    RECT 829.8000 1413.3000 831.0000 1422.3000 ;
	    RECT 833.4000 1420.2001 837.9000 1421.4000 ;
	    RECT 836.7000 1419.3000 837.9000 1420.2001 ;
	    RECT 845.7000 1419.3000 846.9000 1422.9000 ;
	    RECT 849.0000 1421.4000 850.2000 1422.6000 ;
	    RECT 856.8000 1421.7001 858.0000 1422.0000 ;
	    RECT 851.4000 1420.8000 858.0000 1421.7001 ;
	    RECT 851.4000 1420.5000 852.6000 1420.8000 ;
	    RECT 849.0000 1420.2001 850.2000 1420.5000 ;
	    RECT 861.0000 1419.6000 862.2000 1423.8000 ;
	    RECT 869.7000 1422.9000 875.4000 1424.1000 ;
	    RECT 869.7000 1421.1000 870.9000 1422.9000 ;
	    RECT 876.3000 1422.0000 877.2000 1425.0000 ;
	    RECT 851.4000 1419.3000 852.6000 1419.6000 ;
	    RECT 834.6000 1413.3000 835.8000 1419.3000 ;
	    RECT 836.7000 1418.1000 840.6000 1419.3000 ;
	    RECT 845.7000 1418.4000 852.6000 1419.3000 ;
	    RECT 853.8000 1418.4000 855.0000 1419.6000 ;
	    RECT 855.9000 1418.4000 856.2000 1419.6000 ;
	    RECT 860.7000 1418.4000 862.2000 1419.6000 ;
	    RECT 868.2000 1420.2001 870.9000 1421.1000 ;
	    RECT 875.4000 1421.1000 877.2000 1422.0000 ;
	    RECT 868.2000 1419.3000 869.4000 1420.2001 ;
	    RECT 839.4000 1413.3000 840.6000 1418.1000 ;
	    RECT 865.8000 1418.1000 869.4000 1419.3000 ;
	    RECT 841.8000 1413.3000 843.0000 1417.5000 ;
	    RECT 844.2000 1413.3000 845.4000 1417.5000 ;
	    RECT 846.6000 1413.3000 847.8000 1417.5000 ;
	    RECT 849.0000 1413.3000 850.2000 1416.3000 ;
	    RECT 851.4000 1413.3000 852.6000 1417.5000 ;
	    RECT 853.8000 1413.3000 855.0000 1416.3000 ;
	    RECT 856.2000 1413.3000 857.4000 1417.5000 ;
	    RECT 858.6000 1413.3000 859.8000 1417.5000 ;
	    RECT 861.0000 1413.3000 862.2000 1417.5000 ;
	    RECT 863.4000 1413.3000 864.6000 1417.5000 ;
	    RECT 865.8000 1413.3000 867.0000 1418.1000 ;
	    RECT 870.6000 1413.3000 871.8000 1419.3000 ;
	    RECT 875.4000 1413.3000 876.6000 1421.1000 ;
	    RECT 878.1000 1420.2001 879.3000 1426.8000 ;
	    RECT 904.2000 1423.5000 905.4000 1439.7001 ;
	    RECT 923.4000 1433.7001 924.6000 1439.7001 ;
	    RECT 925.8000 1426.5000 927.0000 1439.7001 ;
	    RECT 928.2000 1433.7001 929.4000 1439.7001 ;
	    RECT 940.2000 1439.4000 941.4000 1440.6000 ;
	    RECT 1055.4000 1433.7001 1056.6000 1439.7001 ;
	    RECT 1057.8000 1432.5000 1059.0000 1439.7001 ;
	    RECT 1060.2001 1433.7001 1061.4000 1439.7001 ;
	    RECT 1062.6000 1432.8000 1063.8000 1439.7001 ;
	    RECT 1065.0000 1433.7001 1066.2001 1439.7001 ;
	    RECT 1059.9000 1431.9000 1063.8000 1432.8000 ;
	    RECT 1031.4000 1431.4501 1032.6000 1431.6000 ;
	    RECT 1057.8000 1431.4501 1059.0000 1431.6000 ;
	    RECT 1031.4000 1430.5500 1059.0000 1431.4501 ;
	    RECT 1031.4000 1430.4000 1032.6000 1430.5500 ;
	    RECT 1057.8000 1430.4000 1059.0000 1430.5500 ;
	    RECT 928.2000 1429.5000 929.4000 1429.8000 ;
	    RECT 1059.9000 1429.5000 1060.8000 1431.9000 ;
	    RECT 1067.4000 1431.6000 1068.6000 1439.7001 ;
	    RECT 1069.8000 1433.7001 1071.0000 1439.7001 ;
	    RECT 1072.2001 1435.5000 1073.4000 1439.7001 ;
	    RECT 1074.6000 1435.5000 1075.8000 1439.7001 ;
	    RECT 1077.0000 1435.5000 1078.2001 1439.7001 ;
	    RECT 1069.5000 1431.6000 1075.8000 1432.8000 ;
	    RECT 1064.7001 1430.4000 1068.6000 1431.6000 ;
	    RECT 1079.4000 1430.4000 1080.6000 1439.7001 ;
	    RECT 1081.8000 1433.7001 1083.0000 1439.7001 ;
	    RECT 1084.2001 1432.5000 1085.4000 1439.7001 ;
	    RECT 1086.6000 1433.7001 1087.8000 1439.7001 ;
	    RECT 1089.0000 1432.5000 1090.2001 1439.7001 ;
	    RECT 1091.4000 1435.5000 1092.6000 1439.7001 ;
	    RECT 1093.8000 1435.5000 1095.0000 1439.7001 ;
	    RECT 1096.2001 1433.7001 1097.4000 1439.7001 ;
	    RECT 1098.6000 1432.8000 1099.8000 1439.7001 ;
	    RECT 1101.0000 1433.7001 1102.2001 1440.6000 ;
	    RECT 1103.4000 1434.6000 1104.6000 1439.7001 ;
	    RECT 1103.4000 1433.7001 1104.9000 1434.6000 ;
	    RECT 1105.8000 1433.7001 1107.0000 1439.7001 ;
	    RECT 1140.3000 1433.7001 1141.5000 1439.7001 ;
	    RECT 1104.0000 1432.8000 1104.9000 1433.7001 ;
	    RECT 1096.8000 1431.6000 1103.1000 1432.8000 ;
	    RECT 1104.0000 1431.9000 1107.0000 1432.8000 ;
	    RECT 1084.2001 1430.4000 1088.1000 1431.6000 ;
	    RECT 1089.0000 1430.7001 1097.7001 1431.6000 ;
	    RECT 1102.2001 1431.0000 1103.1000 1431.6000 ;
	    RECT 1072.2001 1429.5000 1073.4000 1429.8000 ;
	    RECT 928.2000 1428.4501 929.4000 1428.6000 ;
	    RECT 966.6000 1428.4501 967.8000 1428.6000 ;
	    RECT 928.2000 1427.5500 967.8000 1428.4501 ;
	    RECT 1057.8000 1428.0000 1059.0000 1429.5000 ;
	    RECT 928.2000 1427.4000 929.4000 1427.5500 ;
	    RECT 966.6000 1427.4000 967.8000 1427.5500 ;
	    RECT 1057.5000 1426.8000 1059.0000 1428.0000 ;
	    RECT 1059.9000 1428.6000 1073.4000 1429.5000 ;
	    RECT 1077.0000 1429.5000 1078.2001 1429.8000 ;
	    RECT 1089.0000 1429.5000 1089.9000 1430.7001 ;
	    RECT 1098.6000 1429.8000 1100.7001 1430.7001 ;
	    RECT 1102.2001 1429.8000 1104.6000 1431.0000 ;
	    RECT 1077.0000 1428.6000 1089.9000 1429.5000 ;
	    RECT 1091.4000 1429.5000 1100.7001 1429.8000 ;
	    RECT 1091.4000 1428.9000 1099.5000 1429.5000 ;
	    RECT 1091.4000 1428.6000 1092.6000 1428.9000 ;
	    RECT 925.8000 1425.4501 927.0000 1425.6000 ;
	    RECT 935.4000 1425.4501 936.6000 1425.6000 ;
	    RECT 925.8000 1424.5500 936.6000 1425.4501 ;
	    RECT 925.8000 1424.4000 927.0000 1424.5500 ;
	    RECT 935.4000 1424.4000 936.6000 1424.5500 ;
	    RECT 904.2000 1421.4000 905.4000 1422.6000 ;
	    RECT 906.6000 1422.4501 907.8000 1422.6000 ;
	    RECT 923.4000 1422.4501 924.6000 1422.6000 ;
	    RECT 906.6000 1421.5500 924.6000 1422.4501 ;
	    RECT 906.6000 1421.4000 907.8000 1421.5500 ;
	    RECT 923.4000 1421.4000 924.6000 1421.5500 ;
	    RECT 877.8000 1419.0000 879.3000 1420.2001 ;
	    RECT 882.6000 1419.4501 883.8000 1419.6000 ;
	    RECT 901.8000 1419.4501 903.0000 1419.6000 ;
	    RECT 877.8000 1413.3000 879.0000 1419.0000 ;
	    RECT 882.6000 1418.5500 903.0000 1419.4501 ;
	    RECT 882.6000 1418.4000 883.8000 1418.5500 ;
	    RECT 901.8000 1418.4000 903.0000 1418.5500 ;
	    RECT 901.8000 1417.2001 903.0000 1417.5000 ;
	    RECT 880.2000 1413.3000 881.4000 1416.3000 ;
	    RECT 901.8000 1413.3000 903.0000 1416.3000 ;
	    RECT 904.2000 1413.3000 905.4000 1420.5000 ;
	    RECT 923.4000 1420.2001 924.6000 1420.5000 ;
	    RECT 925.8000 1419.3000 927.0000 1423.5000 ;
	    RECT 1057.5000 1420.2001 1058.7001 1426.8000 ;
	    RECT 1059.9000 1425.9000 1060.8000 1428.6000 ;
	    RECT 1095.9000 1427.7001 1097.1000 1428.0000 ;
	    RECT 1061.7001 1426.8000 1100.1000 1427.7001 ;
	    RECT 1101.0000 1427.4000 1102.2001 1428.6000 ;
	    RECT 1061.7001 1426.5000 1062.9000 1426.8000 ;
	    RECT 1059.6000 1425.0000 1060.8000 1425.9000 ;
	    RECT 1069.8000 1425.0000 1095.3000 1425.9000 ;
	    RECT 1059.6000 1422.0000 1060.5000 1425.0000 ;
	    RECT 1069.8000 1424.1000 1071.0000 1425.0000 ;
	    RECT 1096.2001 1424.4000 1097.4000 1425.6000 ;
	    RECT 1098.3000 1425.0000 1104.9000 1425.9000 ;
	    RECT 1103.7001 1424.7001 1104.9000 1425.0000 ;
	    RECT 1061.4000 1422.9000 1067.1000 1424.1000 ;
	    RECT 1059.6000 1421.1000 1061.4000 1422.0000 ;
	    RECT 923.4000 1413.3000 924.6000 1419.3000 ;
	    RECT 925.8000 1418.4000 928.5000 1419.3000 ;
	    RECT 1057.5000 1419.0000 1059.0000 1420.2001 ;
	    RECT 927.3000 1413.3000 928.5000 1418.4000 ;
	    RECT 1055.4000 1413.3000 1056.6000 1416.3000 ;
	    RECT 1057.8000 1413.3000 1059.0000 1419.0000 ;
	    RECT 1060.2001 1413.3000 1061.4000 1421.1000 ;
	    RECT 1065.9000 1421.1000 1067.1000 1422.9000 ;
	    RECT 1065.9000 1420.2001 1068.6000 1421.1000 ;
	    RECT 1067.4000 1419.3000 1068.6000 1420.2001 ;
	    RECT 1074.6000 1419.6000 1075.8000 1423.8000 ;
	    RECT 1079.4000 1422.9000 1084.2001 1424.1000 ;
	    RECT 1089.9000 1422.9000 1092.9000 1424.1000 ;
	    RECT 1105.8000 1423.5000 1107.0000 1431.9000 ;
	    RECT 1140.6000 1430.4000 1141.8000 1431.6000 ;
	    RECT 1140.6000 1429.5000 1141.5000 1430.4000 ;
	    RECT 1142.7001 1428.6000 1143.9000 1439.7001 ;
	    RECT 1137.0000 1428.4501 1138.2001 1428.6000 ;
	    RECT 1139.4000 1428.4501 1140.6000 1428.6000 ;
	    RECT 1137.0000 1427.5500 1140.6000 1428.4501 ;
	    RECT 1137.0000 1427.4000 1138.2001 1427.5500 ;
	    RECT 1139.4000 1427.4000 1140.6000 1427.5500 ;
	    RECT 1142.4000 1427.7001 1143.9000 1428.6000 ;
	    RECT 1146.6000 1427.7001 1147.8000 1439.7001 ;
	    RECT 1149.0000 1439.4000 1150.2001 1440.6000 ;
	    RECT 1149.0000 1437.4501 1150.2001 1437.6000 ;
	    RECT 1185.0000 1437.4501 1186.2001 1437.6000 ;
	    RECT 1149.0000 1436.5500 1186.2001 1437.4501 ;
	    RECT 1149.0000 1436.4000 1150.2001 1436.5500 ;
	    RECT 1185.0000 1436.4000 1186.2001 1436.5500 ;
	    RECT 1271.4000 1433.7001 1272.6000 1439.7001 ;
	    RECT 1273.8000 1432.5000 1275.0000 1439.7001 ;
	    RECT 1276.2001 1433.7001 1277.4000 1439.7001 ;
	    RECT 1278.6000 1432.8000 1279.8000 1439.7001 ;
	    RECT 1281.0000 1433.7001 1282.2001 1439.7001 ;
	    RECT 1275.9000 1431.9000 1279.8000 1432.8000 ;
	    RECT 1199.4000 1431.4501 1200.6000 1431.6000 ;
	    RECT 1269.0000 1431.4501 1270.2001 1431.6000 ;
	    RECT 1273.8000 1431.4501 1275.0000 1431.6000 ;
	    RECT 1199.4000 1430.5500 1275.0000 1431.4501 ;
	    RECT 1199.4000 1430.4000 1200.6000 1430.5500 ;
	    RECT 1269.0000 1430.4000 1270.2001 1430.5500 ;
	    RECT 1273.8000 1430.4000 1275.0000 1430.5500 ;
	    RECT 1275.9000 1429.5000 1276.8000 1431.9000 ;
	    RECT 1283.4000 1431.6000 1284.6000 1439.7001 ;
	    RECT 1285.8000 1433.7001 1287.0000 1439.7001 ;
	    RECT 1288.2001 1435.5000 1289.4000 1439.7001 ;
	    RECT 1290.6000 1435.5000 1291.8000 1439.7001 ;
	    RECT 1293.0000 1435.5000 1294.2001 1439.7001 ;
	    RECT 1285.5000 1431.6000 1291.8000 1432.8000 ;
	    RECT 1280.7001 1430.4000 1284.6000 1431.6000 ;
	    RECT 1295.4000 1430.4000 1296.6000 1439.7001 ;
	    RECT 1297.8000 1433.7001 1299.0000 1439.7001 ;
	    RECT 1300.2001 1432.5000 1301.4000 1439.7001 ;
	    RECT 1302.6000 1433.7001 1303.8000 1439.7001 ;
	    RECT 1305.0000 1432.5000 1306.2001 1439.7001 ;
	    RECT 1307.4000 1435.5000 1308.6000 1439.7001 ;
	    RECT 1309.8000 1435.5000 1311.0000 1439.7001 ;
	    RECT 1312.2001 1433.7001 1313.4000 1439.7001 ;
	    RECT 1314.6000 1432.8000 1315.8000 1439.7001 ;
	    RECT 1317.0000 1433.7001 1318.2001 1440.6000 ;
	    RECT 1319.4000 1434.6000 1320.6000 1439.7001 ;
	    RECT 1319.4000 1433.7001 1320.9000 1434.6000 ;
	    RECT 1321.8000 1433.7001 1323.0000 1439.7001 ;
	    RECT 1453.8000 1433.7001 1455.0000 1439.7001 ;
	    RECT 1320.0000 1432.8000 1320.9000 1433.7001 ;
	    RECT 1312.8000 1431.6000 1319.1000 1432.8000 ;
	    RECT 1320.0000 1431.9000 1323.0000 1432.8000 ;
	    RECT 1456.2001 1432.5000 1457.4000 1439.7001 ;
	    RECT 1458.6000 1433.7001 1459.8000 1439.7001 ;
	    RECT 1461.0000 1432.8000 1462.2001 1439.7001 ;
	    RECT 1463.4000 1433.7001 1464.6000 1439.7001 ;
	    RECT 1300.2001 1430.4000 1304.1000 1431.6000 ;
	    RECT 1305.0000 1430.7001 1313.7001 1431.6000 ;
	    RECT 1318.2001 1431.0000 1319.1000 1431.6000 ;
	    RECT 1288.2001 1429.5000 1289.4000 1429.8000 ;
	    RECT 1273.8000 1428.0000 1275.0000 1429.5000 ;
	    RECT 1078.8000 1421.7001 1080.0000 1422.0000 ;
	    RECT 1078.8000 1420.8000 1085.4000 1421.7001 ;
	    RECT 1086.6000 1421.4000 1087.8000 1422.6000 ;
	    RECT 1084.2001 1420.5000 1085.4000 1420.8000 ;
	    RECT 1086.6000 1420.2001 1087.8000 1420.5000 ;
	    RECT 1065.0000 1413.3000 1066.2001 1419.3000 ;
	    RECT 1067.4000 1418.1000 1071.0000 1419.3000 ;
	    RECT 1074.6000 1418.4000 1076.1000 1419.6000 ;
	    RECT 1080.6000 1418.4000 1080.9000 1419.6000 ;
	    RECT 1081.8000 1418.4000 1083.0000 1419.6000 ;
	    RECT 1084.2001 1419.3000 1085.4000 1419.6000 ;
	    RECT 1089.9000 1419.3000 1091.1000 1422.9000 ;
	    RECT 1093.8000 1422.3000 1107.0000 1423.5000 ;
	    RECT 1142.4000 1422.6000 1143.3000 1427.7001 ;
	    RECT 1273.5000 1426.8000 1275.0000 1428.0000 ;
	    RECT 1275.9000 1428.6000 1289.4000 1429.5000 ;
	    RECT 1293.0000 1429.5000 1294.2001 1429.8000 ;
	    RECT 1305.0000 1429.5000 1305.9000 1430.7001 ;
	    RECT 1314.6000 1429.8000 1316.7001 1430.7001 ;
	    RECT 1318.2001 1429.8000 1320.6000 1431.0000 ;
	    RECT 1293.0000 1428.6000 1305.9000 1429.5000 ;
	    RECT 1307.4000 1429.5000 1316.7001 1429.8000 ;
	    RECT 1307.4000 1428.9000 1315.5000 1429.5000 ;
	    RECT 1307.4000 1428.6000 1308.6000 1428.9000 ;
	    RECT 1144.2001 1424.4000 1145.4000 1425.6000 ;
	    RECT 1144.2001 1423.2001 1145.4000 1423.5000 ;
	    RECT 1098.9000 1420.2001 1103.4000 1421.4000 ;
	    RECT 1098.9000 1419.3000 1100.1000 1420.2001 ;
	    RECT 1084.2001 1418.4000 1091.1000 1419.3000 ;
	    RECT 1069.8000 1413.3000 1071.0000 1418.1000 ;
	    RECT 1096.2001 1418.1000 1100.1000 1419.3000 ;
	    RECT 1072.2001 1413.3000 1073.4000 1417.5000 ;
	    RECT 1074.6000 1413.3000 1075.8000 1417.5000 ;
	    RECT 1077.0000 1413.3000 1078.2001 1417.5000 ;
	    RECT 1079.4000 1413.3000 1080.6000 1417.5000 ;
	    RECT 1081.8000 1413.3000 1083.0000 1416.3000 ;
	    RECT 1084.2001 1413.3000 1085.4000 1417.5000 ;
	    RECT 1086.6000 1413.3000 1087.8000 1416.3000 ;
	    RECT 1089.0000 1413.3000 1090.2001 1417.5000 ;
	    RECT 1091.4000 1413.3000 1092.6000 1417.5000 ;
	    RECT 1093.8000 1413.3000 1095.0000 1417.5000 ;
	    RECT 1096.2001 1413.3000 1097.4000 1418.1000 ;
	    RECT 1101.0000 1413.3000 1102.2001 1419.3000 ;
	    RECT 1105.8000 1413.3000 1107.0000 1422.3000 ;
	    RECT 1110.6000 1422.4501 1111.8000 1422.6000 ;
	    RECT 1139.4000 1422.4501 1140.6000 1422.6000 ;
	    RECT 1110.6000 1421.5500 1140.6000 1422.4501 ;
	    RECT 1110.6000 1421.4000 1111.8000 1421.5500 ;
	    RECT 1139.4000 1421.4000 1140.6000 1421.5500 ;
	    RECT 1141.5000 1421.4000 1143.3000 1422.6000 ;
	    RECT 1146.6000 1422.4501 1147.8000 1422.6000 ;
	    RECT 1149.0000 1422.4501 1150.2001 1422.6000 ;
	    RECT 1145.4000 1420.8000 1145.7001 1422.3000 ;
	    RECT 1146.6000 1421.5500 1150.2001 1422.4501 ;
	    RECT 1146.6000 1421.4000 1147.8000 1421.5500 ;
	    RECT 1149.0000 1421.4000 1150.2001 1421.5500 ;
	    RECT 1139.7001 1419.3000 1140.6000 1420.5000 ;
	    RECT 1273.5000 1420.2001 1274.7001 1426.8000 ;
	    RECT 1275.9000 1425.9000 1276.8000 1428.6000 ;
	    RECT 1311.9000 1427.7001 1313.1000 1428.0000 ;
	    RECT 1277.7001 1426.8000 1316.1000 1427.7001 ;
	    RECT 1317.0000 1427.4000 1318.2001 1428.6000 ;
	    RECT 1277.7001 1426.5000 1278.9000 1426.8000 ;
	    RECT 1275.6000 1425.0000 1276.8000 1425.9000 ;
	    RECT 1285.8000 1425.0000 1311.3000 1425.9000 ;
	    RECT 1275.6000 1422.0000 1276.5000 1425.0000 ;
	    RECT 1285.8000 1424.1000 1287.0000 1425.0000 ;
	    RECT 1312.2001 1424.4000 1313.4000 1425.6000 ;
	    RECT 1314.3000 1425.0000 1320.9000 1425.9000 ;
	    RECT 1319.7001 1424.7001 1320.9000 1425.0000 ;
	    RECT 1277.4000 1422.9000 1283.1000 1424.1000 ;
	    RECT 1275.6000 1421.1000 1277.4000 1422.0000 ;
	    RECT 1142.1000 1419.3000 1147.5000 1419.9000 ;
	    RECT 1139.4000 1413.3000 1140.6000 1419.3000 ;
	    RECT 1141.8000 1419.0000 1147.8000 1419.3000 ;
	    RECT 1273.5000 1419.0000 1275.0000 1420.2001 ;
	    RECT 1141.8000 1413.3000 1143.0000 1419.0000 ;
	    RECT 1144.2001 1413.3000 1145.4000 1418.1000 ;
	    RECT 1146.6000 1413.3000 1147.8000 1419.0000 ;
	    RECT 1271.4000 1413.3000 1272.6000 1416.3000 ;
	    RECT 1273.8000 1413.3000 1275.0000 1419.0000 ;
	    RECT 1276.2001 1413.3000 1277.4000 1421.1000 ;
	    RECT 1281.9000 1421.1000 1283.1000 1422.9000 ;
	    RECT 1281.9000 1420.2001 1284.6000 1421.1000 ;
	    RECT 1283.4000 1419.3000 1284.6000 1420.2001 ;
	    RECT 1290.6000 1419.6000 1291.8000 1423.8000 ;
	    RECT 1295.4000 1422.9000 1300.2001 1424.1000 ;
	    RECT 1305.9000 1422.9000 1308.9000 1424.1000 ;
	    RECT 1321.8000 1423.5000 1323.0000 1431.9000 ;
	    RECT 1458.3000 1431.9000 1462.2001 1432.8000 ;
	    RECT 1333.8000 1431.4501 1335.0000 1431.6000 ;
	    RECT 1456.2001 1431.4501 1457.4000 1431.6000 ;
	    RECT 1333.8000 1430.5500 1457.4000 1431.4501 ;
	    RECT 1333.8000 1430.4000 1335.0000 1430.5500 ;
	    RECT 1456.2001 1430.4000 1457.4000 1430.5500 ;
	    RECT 1458.3000 1429.5000 1459.2001 1431.9000 ;
	    RECT 1465.8000 1431.6000 1467.0000 1439.7001 ;
	    RECT 1468.2001 1433.7001 1469.4000 1439.7001 ;
	    RECT 1470.6000 1435.5000 1471.8000 1439.7001 ;
	    RECT 1473.0000 1435.5000 1474.2001 1439.7001 ;
	    RECT 1475.4000 1435.5000 1476.6000 1439.7001 ;
	    RECT 1467.9000 1431.6000 1474.2001 1432.8000 ;
	    RECT 1463.1000 1430.4000 1467.0000 1431.6000 ;
	    RECT 1477.8000 1430.4000 1479.0000 1439.7001 ;
	    RECT 1480.2001 1433.7001 1481.4000 1439.7001 ;
	    RECT 1482.6000 1432.5000 1483.8000 1439.7001 ;
	    RECT 1485.0000 1433.7001 1486.2001 1439.7001 ;
	    RECT 1487.4000 1432.5000 1488.6000 1439.7001 ;
	    RECT 1489.8000 1435.5000 1491.0000 1439.7001 ;
	    RECT 1492.2001 1435.5000 1493.4000 1439.7001 ;
	    RECT 1494.6000 1433.7001 1495.8000 1439.7001 ;
	    RECT 1497.0000 1432.8000 1498.2001 1439.7001 ;
	    RECT 1499.4000 1433.7001 1500.6000 1440.6000 ;
	    RECT 1501.8000 1434.6000 1503.0000 1439.7001 ;
	    RECT 1501.8000 1433.7001 1503.3000 1434.6000 ;
	    RECT 1504.2001 1433.7001 1505.4000 1439.7001 ;
	    RECT 1502.4000 1432.8000 1503.3000 1433.7001 ;
	    RECT 1495.2001 1431.6000 1501.5000 1432.8000 ;
	    RECT 1502.4000 1431.9000 1505.4000 1432.8000 ;
	    RECT 1482.6000 1430.4000 1486.5000 1431.6000 ;
	    RECT 1487.4000 1430.7001 1496.1000 1431.6000 ;
	    RECT 1500.6000 1431.0000 1501.5000 1431.6000 ;
	    RECT 1470.6000 1429.5000 1471.8000 1429.8000 ;
	    RECT 1456.2001 1428.0000 1457.4000 1429.5000 ;
	    RECT 1294.8000 1421.7001 1296.0000 1422.0000 ;
	    RECT 1294.8000 1420.8000 1301.4000 1421.7001 ;
	    RECT 1302.6000 1421.4000 1303.8000 1422.6000 ;
	    RECT 1300.2001 1420.5000 1301.4000 1420.8000 ;
	    RECT 1302.6000 1420.2001 1303.8000 1420.5000 ;
	    RECT 1281.0000 1413.3000 1282.2001 1419.3000 ;
	    RECT 1283.4000 1418.1000 1287.0000 1419.3000 ;
	    RECT 1290.6000 1418.4000 1292.1000 1419.6000 ;
	    RECT 1296.6000 1418.4000 1296.9000 1419.6000 ;
	    RECT 1297.8000 1418.4000 1299.0000 1419.6000 ;
	    RECT 1300.2001 1419.3000 1301.4000 1419.6000 ;
	    RECT 1305.9000 1419.3000 1307.1000 1422.9000 ;
	    RECT 1309.8000 1422.3000 1323.0000 1423.5000 ;
	    RECT 1314.9000 1420.2001 1319.4000 1421.4000 ;
	    RECT 1314.9000 1419.3000 1316.1000 1420.2001 ;
	    RECT 1300.2001 1418.4000 1307.1000 1419.3000 ;
	    RECT 1285.8000 1413.3000 1287.0000 1418.1000 ;
	    RECT 1312.2001 1418.1000 1316.1000 1419.3000 ;
	    RECT 1288.2001 1413.3000 1289.4000 1417.5000 ;
	    RECT 1290.6000 1413.3000 1291.8000 1417.5000 ;
	    RECT 1293.0000 1413.3000 1294.2001 1417.5000 ;
	    RECT 1295.4000 1413.3000 1296.6000 1417.5000 ;
	    RECT 1297.8000 1413.3000 1299.0000 1416.3000 ;
	    RECT 1300.2001 1413.3000 1301.4000 1417.5000 ;
	    RECT 1302.6000 1413.3000 1303.8000 1416.3000 ;
	    RECT 1305.0000 1413.3000 1306.2001 1417.5000 ;
	    RECT 1307.4000 1413.3000 1308.6000 1417.5000 ;
	    RECT 1309.8000 1413.3000 1311.0000 1417.5000 ;
	    RECT 1312.2001 1413.3000 1313.4000 1418.1000 ;
	    RECT 1317.0000 1413.3000 1318.2001 1419.3000 ;
	    RECT 1321.8000 1413.3000 1323.0000 1422.3000 ;
	    RECT 1455.9000 1426.8000 1457.4000 1428.0000 ;
	    RECT 1458.3000 1428.6000 1471.8000 1429.5000 ;
	    RECT 1475.4000 1429.5000 1476.6000 1429.8000 ;
	    RECT 1487.4000 1429.5000 1488.3000 1430.7001 ;
	    RECT 1497.0000 1429.8000 1499.1000 1430.7001 ;
	    RECT 1500.6000 1429.8000 1503.0000 1431.0000 ;
	    RECT 1475.4000 1428.6000 1488.3000 1429.5000 ;
	    RECT 1489.8000 1429.5000 1499.1000 1429.8000 ;
	    RECT 1489.8000 1428.9000 1497.9000 1429.5000 ;
	    RECT 1489.8000 1428.6000 1491.0000 1428.9000 ;
	    RECT 1455.9000 1420.2001 1457.1000 1426.8000 ;
	    RECT 1458.3000 1425.9000 1459.2001 1428.6000 ;
	    RECT 1494.3000 1427.7001 1495.5000 1428.0000 ;
	    RECT 1460.1000 1426.8000 1498.5000 1427.7001 ;
	    RECT 1499.4000 1427.4000 1500.6000 1428.6000 ;
	    RECT 1460.1000 1426.5000 1461.3000 1426.8000 ;
	    RECT 1458.0000 1425.0000 1459.2001 1425.9000 ;
	    RECT 1468.2001 1425.0000 1493.7001 1425.9000 ;
	    RECT 1458.0000 1422.0000 1458.9000 1425.0000 ;
	    RECT 1468.2001 1424.1000 1469.4000 1425.0000 ;
	    RECT 1494.6000 1424.4000 1495.8000 1425.6000 ;
	    RECT 1496.7001 1425.0000 1503.3000 1425.9000 ;
	    RECT 1502.1000 1424.7001 1503.3000 1425.0000 ;
	    RECT 1459.8000 1422.9000 1465.5000 1424.1000 ;
	    RECT 1458.0000 1421.1000 1459.8000 1422.0000 ;
	    RECT 1455.9000 1419.0000 1457.4000 1420.2001 ;
	    RECT 1453.8000 1413.3000 1455.0000 1416.3000 ;
	    RECT 1456.2001 1413.3000 1457.4000 1419.0000 ;
	    RECT 1458.6000 1413.3000 1459.8000 1421.1000 ;
	    RECT 1464.3000 1421.1000 1465.5000 1422.9000 ;
	    RECT 1464.3000 1420.2001 1467.0000 1421.1000 ;
	    RECT 1465.8000 1419.3000 1467.0000 1420.2001 ;
	    RECT 1473.0000 1419.6000 1474.2001 1423.8000 ;
	    RECT 1477.8000 1422.9000 1482.6000 1424.1000 ;
	    RECT 1488.3000 1422.9000 1491.3000 1424.1000 ;
	    RECT 1504.2001 1423.5000 1505.4000 1431.9000 ;
	    RECT 1518.6000 1423.5000 1519.8000 1439.7001 ;
	    RECT 1521.0000 1433.7001 1522.2001 1439.7001 ;
	    RECT 1540.2001 1428.6000 1541.4000 1439.7001 ;
	    RECT 1542.6000 1429.5000 1543.8000 1439.7001 ;
	    RECT 1540.2001 1427.7001 1543.5000 1428.6000 ;
	    RECT 1545.0000 1427.7001 1546.2001 1439.7001 ;
	    RECT 1542.6000 1426.8000 1543.5000 1427.7001 ;
	    RECT 1542.6000 1425.6000 1544.4000 1426.8000 ;
	    RECT 1540.2001 1424.4000 1541.4000 1425.6000 ;
	    RECT 1477.2001 1421.7001 1478.4000 1422.0000 ;
	    RECT 1477.2001 1420.8000 1483.8000 1421.7001 ;
	    RECT 1485.0000 1421.4000 1486.2001 1422.6000 ;
	    RECT 1482.6000 1420.5000 1483.8000 1420.8000 ;
	    RECT 1485.0000 1420.2001 1486.2001 1420.5000 ;
	    RECT 1463.4000 1413.3000 1464.6000 1419.3000 ;
	    RECT 1465.8000 1418.1000 1469.4000 1419.3000 ;
	    RECT 1473.0000 1418.4000 1474.5000 1419.6000 ;
	    RECT 1479.0000 1418.4000 1479.3000 1419.6000 ;
	    RECT 1480.2001 1418.4000 1481.4000 1419.6000 ;
	    RECT 1482.6000 1419.3000 1483.8000 1419.6000 ;
	    RECT 1488.3000 1419.3000 1489.5000 1422.9000 ;
	    RECT 1492.2001 1422.3000 1505.4000 1423.5000 ;
	    RECT 1540.2001 1423.2001 1541.4000 1423.5000 ;
	    RECT 1497.3000 1420.2001 1501.8000 1421.4000 ;
	    RECT 1497.3000 1419.3000 1498.5000 1420.2001 ;
	    RECT 1482.6000 1418.4000 1489.5000 1419.3000 ;
	    RECT 1468.2001 1413.3000 1469.4000 1418.1000 ;
	    RECT 1494.6000 1418.1000 1498.5000 1419.3000 ;
	    RECT 1470.6000 1413.3000 1471.8000 1417.5000 ;
	    RECT 1473.0000 1413.3000 1474.2001 1417.5000 ;
	    RECT 1475.4000 1413.3000 1476.6000 1417.5000 ;
	    RECT 1477.8000 1413.3000 1479.0000 1417.5000 ;
	    RECT 1480.2001 1413.3000 1481.4000 1416.3000 ;
	    RECT 1482.6000 1413.3000 1483.8000 1417.5000 ;
	    RECT 1485.0000 1413.3000 1486.2001 1416.3000 ;
	    RECT 1487.4000 1413.3000 1488.6000 1417.5000 ;
	    RECT 1489.8000 1413.3000 1491.0000 1417.5000 ;
	    RECT 1492.2001 1413.3000 1493.4000 1417.5000 ;
	    RECT 1494.6000 1413.3000 1495.8000 1418.1000 ;
	    RECT 1499.4000 1413.3000 1500.6000 1419.3000 ;
	    RECT 1504.2001 1413.3000 1505.4000 1422.3000 ;
	    RECT 1506.6000 1422.4501 1507.8000 1422.6000 ;
	    RECT 1518.6000 1422.4501 1519.8000 1422.6000 ;
	    RECT 1506.6000 1421.5500 1519.8000 1422.4501 ;
	    RECT 1506.6000 1421.4000 1507.8000 1421.5500 ;
	    RECT 1518.6000 1421.4000 1519.8000 1421.5500 ;
	    RECT 1542.6000 1421.1000 1543.5000 1425.6000 ;
	    RECT 1545.3000 1424.4000 1546.2001 1427.7001 ;
	    RECT 1545.0000 1423.5000 1546.2001 1424.4000 ;
	    RECT 1518.6000 1413.3000 1519.8000 1420.5000 ;
	    RECT 1540.2001 1420.2001 1543.5000 1421.1000 ;
	    RECT 1521.0000 1419.4501 1522.2001 1419.6000 ;
	    RECT 1523.4000 1419.4501 1524.6000 1419.6000 ;
	    RECT 1521.0000 1418.5500 1524.6000 1419.4501 ;
	    RECT 1521.0000 1418.4000 1522.2001 1418.5500 ;
	    RECT 1523.4000 1418.4000 1524.6000 1418.5500 ;
	    RECT 1521.0000 1417.2001 1522.2001 1417.5000 ;
	    RECT 1521.0000 1413.3000 1522.2001 1416.3000 ;
	    RECT 1540.2001 1413.3000 1541.4000 1420.2001 ;
	    RECT 1542.6000 1413.3000 1543.8000 1419.3000 ;
	    RECT 1545.0000 1413.3000 1546.2001 1420.5000 ;
	    RECT 1.2000 1410.6000 1569.0000 1412.4000 ;
	    RECT 124.2000 1406.7001 125.4000 1409.7001 ;
	    RECT 126.6000 1404.0000 127.8000 1409.7001 ;
	    RECT 126.3000 1402.8000 127.8000 1404.0000 ;
	    RECT 126.3000 1396.2001 127.5000 1402.8000 ;
	    RECT 129.0000 1401.9000 130.2000 1409.7001 ;
	    RECT 133.8000 1403.7001 135.0000 1409.7001 ;
	    RECT 138.6000 1404.9000 139.8000 1409.7001 ;
	    RECT 141.0000 1405.5000 142.2000 1409.7001 ;
	    RECT 143.4000 1405.5000 144.6000 1409.7001 ;
	    RECT 145.8000 1405.5000 147.0000 1409.7001 ;
	    RECT 148.2000 1405.5000 149.4000 1409.7001 ;
	    RECT 150.6000 1406.7001 151.8000 1409.7001 ;
	    RECT 153.0000 1405.5000 154.2000 1409.7001 ;
	    RECT 155.4000 1406.7001 156.6000 1409.7001 ;
	    RECT 157.8000 1405.5000 159.0000 1409.7001 ;
	    RECT 160.2000 1405.5000 161.4000 1409.7001 ;
	    RECT 162.6000 1405.5000 163.8000 1409.7001 ;
	    RECT 136.2000 1403.7001 139.8000 1404.9000 ;
	    RECT 165.0000 1404.9000 166.2000 1409.7001 ;
	    RECT 136.2000 1402.8000 137.4000 1403.7001 ;
	    RECT 128.4000 1401.0000 130.2000 1401.9000 ;
	    RECT 134.7000 1401.9000 137.4000 1402.8000 ;
	    RECT 143.4000 1403.4000 144.9000 1404.6000 ;
	    RECT 149.4000 1403.4000 149.7000 1404.6000 ;
	    RECT 150.6000 1403.4000 151.8000 1404.6000 ;
	    RECT 153.0000 1403.7001 159.9000 1404.6000 ;
	    RECT 165.0000 1403.7001 168.9000 1404.9000 ;
	    RECT 169.8000 1403.7001 171.0000 1409.7001 ;
	    RECT 153.0000 1403.4000 154.2000 1403.7001 ;
	    RECT 128.4000 1398.0000 129.3000 1401.0000 ;
	    RECT 134.7000 1400.1000 135.9000 1401.9000 ;
	    RECT 130.2000 1398.9000 135.9000 1400.1000 ;
	    RECT 143.4000 1399.2001 144.6000 1403.4000 ;
	    RECT 155.4000 1402.5000 156.6000 1402.8000 ;
	    RECT 153.0000 1402.2001 154.2000 1402.5000 ;
	    RECT 147.6000 1401.3000 154.2000 1402.2001 ;
	    RECT 147.6000 1401.0000 148.8000 1401.3000 ;
	    RECT 155.4000 1400.4000 156.6000 1401.6000 ;
	    RECT 158.7000 1400.1000 159.9000 1403.7001 ;
	    RECT 167.7000 1402.8000 168.9000 1403.7001 ;
	    RECT 167.7000 1401.6000 172.2000 1402.8000 ;
	    RECT 174.6000 1400.7001 175.8000 1409.7001 ;
	    RECT 198.6000 1403.7001 199.8000 1409.7001 ;
	    RECT 201.0000 1404.0000 202.2000 1409.7001 ;
	    RECT 203.4000 1404.9000 204.6000 1409.7001 ;
	    RECT 205.8000 1404.0000 207.0000 1409.7001 ;
	    RECT 201.0000 1403.7001 207.0000 1404.0000 ;
	    RECT 232.2000 1403.7001 233.4000 1409.7001 ;
	    RECT 236.1000 1404.6000 237.3000 1409.7001 ;
	    RECT 234.6000 1403.7001 237.3000 1404.6000 ;
	    RECT 261.0000 1403.7001 262.2000 1409.7001 ;
	    RECT 263.4000 1404.0000 264.6000 1409.7001 ;
	    RECT 265.8000 1404.9000 267.0000 1409.7001 ;
	    RECT 268.2000 1404.0000 269.4000 1409.7001 ;
	    RECT 280.2000 1406.7001 281.4000 1409.7001 ;
	    RECT 280.2000 1405.5000 281.4000 1405.8000 ;
	    RECT 263.4000 1403.7001 269.4000 1404.0000 ;
	    RECT 198.9000 1402.5000 199.8000 1403.7001 ;
	    RECT 201.3000 1403.1000 206.7000 1403.7001 ;
	    RECT 232.2000 1402.5000 233.4000 1402.8000 ;
	    RECT 148.2000 1398.9000 153.0000 1400.1000 ;
	    RECT 158.7000 1398.9000 161.7000 1400.1000 ;
	    RECT 162.6000 1399.5000 175.8000 1400.7001 ;
	    RECT 177.0000 1401.4501 178.2000 1401.6000 ;
	    RECT 198.6000 1401.4501 199.8000 1401.6000 ;
	    RECT 177.0000 1400.5500 199.8000 1401.4501 ;
	    RECT 177.0000 1400.4000 178.2000 1400.5500 ;
	    RECT 198.6000 1400.4000 199.8000 1400.5500 ;
	    RECT 200.7000 1400.4000 202.5000 1401.6000 ;
	    RECT 204.6000 1400.7001 204.9000 1402.2001 ;
	    RECT 205.8000 1401.4501 207.0000 1401.6000 ;
	    RECT 220.2000 1401.4501 221.4000 1401.6000 ;
	    RECT 232.2000 1401.4501 233.4000 1401.6000 ;
	    RECT 205.8000 1400.5500 233.4000 1401.4501 ;
	    RECT 205.8000 1400.4000 207.0000 1400.5500 ;
	    RECT 220.2000 1400.4000 221.4000 1400.5500 ;
	    RECT 232.2000 1400.4000 233.4000 1400.5500 ;
	    RECT 138.6000 1398.0000 139.8000 1398.9000 ;
	    RECT 128.4000 1397.1000 129.6000 1398.0000 ;
	    RECT 138.6000 1397.1000 164.1000 1398.0000 ;
	    RECT 165.0000 1397.4000 166.2000 1398.6000 ;
	    RECT 172.5000 1398.0000 173.7000 1398.3000 ;
	    RECT 167.1000 1397.1000 173.7000 1398.0000 ;
	    RECT 126.3000 1395.0000 127.8000 1396.2001 ;
	    RECT 126.6000 1393.5000 127.8000 1395.0000 ;
	    RECT 128.7000 1394.4000 129.6000 1397.1000 ;
	    RECT 130.5000 1396.2001 131.7000 1396.5000 ;
	    RECT 130.5000 1395.3000 168.9000 1396.2001 ;
	    RECT 164.7000 1395.0000 165.9000 1395.3000 ;
	    RECT 169.8000 1394.4000 171.0000 1395.6000 ;
	    RECT 128.7000 1393.5000 142.2000 1394.4000 ;
	    RECT 126.6000 1391.4000 127.8000 1392.6000 ;
	    RECT 128.7000 1391.1000 129.6000 1393.5000 ;
	    RECT 141.0000 1393.2001 142.2000 1393.5000 ;
	    RECT 145.8000 1393.5000 158.7000 1394.4000 ;
	    RECT 145.8000 1393.2001 147.0000 1393.5000 ;
	    RECT 133.5000 1391.4000 137.4000 1392.6000 ;
	    RECT 124.2000 1383.3000 125.4000 1389.3000 ;
	    RECT 126.6000 1383.3000 127.8000 1390.5000 ;
	    RECT 128.7000 1390.2001 132.6000 1391.1000 ;
	    RECT 129.0000 1383.3000 130.2000 1389.3000 ;
	    RECT 131.4000 1383.3000 132.6000 1390.2001 ;
	    RECT 133.8000 1383.3000 135.0000 1389.3000 ;
	    RECT 136.2000 1383.3000 137.4000 1391.4000 ;
	    RECT 138.3000 1390.2001 144.6000 1391.4000 ;
	    RECT 138.6000 1383.3000 139.8000 1389.3000 ;
	    RECT 141.0000 1383.3000 142.2000 1387.5000 ;
	    RECT 143.4000 1383.3000 144.6000 1387.5000 ;
	    RECT 145.8000 1383.3000 147.0000 1387.5000 ;
	    RECT 148.2000 1383.3000 149.4000 1392.6000 ;
	    RECT 153.0000 1391.4000 156.9000 1392.6000 ;
	    RECT 157.8000 1392.3000 158.7000 1393.5000 ;
	    RECT 160.2000 1394.1000 161.4000 1394.4000 ;
	    RECT 160.2000 1393.5000 168.3000 1394.1000 ;
	    RECT 160.2000 1393.2001 169.5000 1393.5000 ;
	    RECT 167.4000 1392.3000 169.5000 1393.2001 ;
	    RECT 157.8000 1391.4000 166.5000 1392.3000 ;
	    RECT 171.0000 1392.0000 173.4000 1393.2001 ;
	    RECT 171.0000 1391.4000 171.9000 1392.0000 ;
	    RECT 150.6000 1383.3000 151.8000 1389.3000 ;
	    RECT 153.0000 1383.3000 154.2000 1390.5000 ;
	    RECT 155.4000 1383.3000 156.6000 1389.3000 ;
	    RECT 157.8000 1383.3000 159.0000 1390.5000 ;
	    RECT 165.6000 1390.2001 171.9000 1391.4000 ;
	    RECT 174.6000 1391.1000 175.8000 1399.5000 ;
	    RECT 198.6000 1394.4000 199.8000 1395.6000 ;
	    RECT 201.6000 1395.3000 202.5000 1400.4000 ;
	    RECT 203.4000 1399.5000 204.6000 1399.8000 ;
	    RECT 234.6000 1399.5000 235.8000 1403.7001 ;
	    RECT 261.3000 1402.5000 262.2000 1403.7001 ;
	    RECT 263.7000 1403.1000 269.1000 1403.7001 ;
	    RECT 280.2000 1403.4000 281.4000 1404.6000 ;
	    RECT 282.6000 1402.5000 283.8000 1409.7001 ;
	    RECT 297.0000 1402.5000 298.2000 1409.7001 ;
	    RECT 299.4000 1406.7001 300.6000 1409.7001 ;
	    RECT 299.4000 1405.5000 300.6000 1405.8000 ;
	    RECT 299.4000 1404.4501 300.6000 1404.6000 ;
	    RECT 311.4000 1404.4501 312.6000 1404.6000 ;
	    RECT 299.4000 1403.5500 312.6000 1404.4501 ;
	    RECT 299.4000 1403.4000 300.6000 1403.5500 ;
	    RECT 311.4000 1403.4000 312.6000 1403.5500 ;
	    RECT 313.8000 1402.5000 315.0000 1409.7001 ;
	    RECT 316.2000 1406.7001 317.4000 1409.7001 ;
	    RECT 330.6000 1406.7001 331.8000 1409.7001 ;
	    RECT 316.2000 1405.5000 317.4000 1405.8000 ;
	    RECT 330.6000 1405.5000 331.8000 1405.8000 ;
	    RECT 316.2000 1403.4000 317.4000 1404.6000 ;
	    RECT 330.6000 1403.4000 331.8000 1404.6000 ;
	    RECT 333.0000 1402.5000 334.2000 1409.7001 ;
	    RECT 340.2000 1407.4501 341.4000 1407.6000 ;
	    RECT 347.4000 1407.4501 348.6000 1407.6000 ;
	    RECT 340.2000 1406.5500 348.6000 1407.4501 ;
	    RECT 465.0000 1406.7001 466.2000 1409.7001 ;
	    RECT 340.2000 1406.4000 341.4000 1406.5500 ;
	    RECT 347.4000 1406.4000 348.6000 1406.5500 ;
	    RECT 467.4000 1404.0000 468.6000 1409.7001 ;
	    RECT 467.1000 1402.8000 468.6000 1404.0000 ;
	    RECT 261.0000 1400.4000 262.2000 1401.6000 ;
	    RECT 263.1000 1400.4000 264.9000 1401.6000 ;
	    RECT 267.0000 1400.7001 267.3000 1402.2001 ;
	    RECT 268.2000 1401.4501 269.4000 1401.6000 ;
	    RECT 270.6000 1401.4501 271.8000 1401.6000 ;
	    RECT 268.2000 1400.5500 271.8000 1401.4501 ;
	    RECT 268.2000 1400.4000 269.4000 1400.5500 ;
	    RECT 270.6000 1400.4000 271.8000 1400.5500 ;
	    RECT 282.6000 1400.4000 283.8000 1401.6000 ;
	    RECT 285.0000 1401.4501 286.2000 1401.6000 ;
	    RECT 297.0000 1401.4501 298.2000 1401.6000 ;
	    RECT 285.0000 1400.5500 298.2000 1401.4501 ;
	    RECT 285.0000 1400.4000 286.2000 1400.5500 ;
	    RECT 297.0000 1400.4000 298.2000 1400.5500 ;
	    RECT 313.8000 1400.4000 315.0000 1401.6000 ;
	    RECT 333.0000 1401.4501 334.2000 1401.6000 ;
	    RECT 457.8000 1401.4501 459.0000 1401.6000 ;
	    RECT 333.0000 1400.5500 459.0000 1401.4501 ;
	    RECT 333.0000 1400.4000 334.2000 1400.5500 ;
	    RECT 457.8000 1400.4000 459.0000 1400.5500 ;
	    RECT 203.4000 1397.4000 204.6000 1398.6000 ;
	    RECT 234.6000 1398.4501 235.8000 1398.6000 ;
	    RECT 234.6000 1397.5500 262.0500 1398.4501 ;
	    RECT 234.6000 1397.4000 235.8000 1397.5500 ;
	    RECT 201.6000 1394.4000 203.1000 1395.3000 ;
	    RECT 199.8000 1392.6000 200.7000 1393.5000 ;
	    RECT 199.8000 1391.4000 201.0000 1392.6000 ;
	    RECT 172.8000 1390.2001 175.8000 1391.1000 ;
	    RECT 160.2000 1383.3000 161.4000 1387.5000 ;
	    RECT 162.6000 1383.3000 163.8000 1387.5000 ;
	    RECT 165.0000 1383.3000 166.2000 1389.3000 ;
	    RECT 167.4000 1383.3000 168.6000 1390.2001 ;
	    RECT 172.8000 1389.3000 173.7000 1390.2001 ;
	    RECT 169.8000 1382.4000 171.0000 1389.3000 ;
	    RECT 172.2000 1388.4000 173.7000 1389.3000 ;
	    RECT 172.2000 1383.3000 173.4000 1388.4000 ;
	    RECT 174.6000 1383.3000 175.8000 1389.3000 ;
	    RECT 199.5000 1383.3000 200.7000 1389.3000 ;
	    RECT 201.9000 1383.3000 203.1000 1394.4000 ;
	    RECT 205.8000 1383.3000 207.0000 1395.3000 ;
	    RECT 232.2000 1383.3000 233.4000 1389.3000 ;
	    RECT 234.6000 1383.3000 235.8000 1396.5000 ;
	    RECT 261.1500 1395.6000 262.0500 1397.5500 ;
	    RECT 237.0000 1394.4000 238.2000 1395.6000 ;
	    RECT 261.0000 1394.4000 262.2000 1395.6000 ;
	    RECT 264.0000 1395.3000 264.9000 1400.4000 ;
	    RECT 265.8000 1399.5000 267.0000 1399.8000 ;
	    RECT 265.8000 1397.4000 267.0000 1398.6000 ;
	    RECT 264.0000 1394.4000 265.5000 1395.3000 ;
	    RECT 237.0000 1393.2001 238.2000 1393.5000 ;
	    RECT 262.2000 1392.6000 263.1000 1393.5000 ;
	    RECT 262.2000 1391.4000 263.4000 1392.6000 ;
	    RECT 237.0000 1383.3000 238.2000 1389.3000 ;
	    RECT 261.9000 1383.3000 263.1000 1389.3000 ;
	    RECT 264.3000 1383.3000 265.5000 1394.4000 ;
	    RECT 268.2000 1383.3000 269.4000 1395.3000 ;
	    RECT 280.2000 1383.3000 281.4000 1389.3000 ;
	    RECT 282.6000 1383.3000 283.8000 1399.5000 ;
	    RECT 297.0000 1383.3000 298.2000 1399.5000 ;
	    RECT 299.4000 1383.3000 300.6000 1389.3000 ;
	    RECT 313.8000 1383.3000 315.0000 1399.5000 ;
	    RECT 316.2000 1383.3000 317.4000 1389.3000 ;
	    RECT 330.6000 1383.3000 331.8000 1389.3000 ;
	    RECT 333.0000 1383.3000 334.2000 1399.5000 ;
	    RECT 467.1000 1396.2001 468.3000 1402.8000 ;
	    RECT 469.8000 1401.9000 471.0000 1409.7001 ;
	    RECT 474.6000 1403.7001 475.8000 1409.7001 ;
	    RECT 479.4000 1404.9000 480.6000 1409.7001 ;
	    RECT 481.8000 1405.5000 483.0000 1409.7001 ;
	    RECT 484.2000 1405.5000 485.4000 1409.7001 ;
	    RECT 486.6000 1405.5000 487.8000 1409.7001 ;
	    RECT 489.0000 1405.5000 490.2000 1409.7001 ;
	    RECT 491.4000 1406.7001 492.6000 1409.7001 ;
	    RECT 493.8000 1405.5000 495.0000 1409.7001 ;
	    RECT 496.2000 1406.7001 497.4000 1409.7001 ;
	    RECT 498.6000 1405.5000 499.8000 1409.7001 ;
	    RECT 501.0000 1405.5000 502.2000 1409.7001 ;
	    RECT 503.4000 1405.5000 504.6000 1409.7001 ;
	    RECT 477.0000 1403.7001 480.6000 1404.9000 ;
	    RECT 505.8000 1404.9000 507.0000 1409.7001 ;
	    RECT 477.0000 1402.8000 478.2000 1403.7001 ;
	    RECT 469.2000 1401.0000 471.0000 1401.9000 ;
	    RECT 475.5000 1401.9000 478.2000 1402.8000 ;
	    RECT 484.2000 1403.4000 485.7000 1404.6000 ;
	    RECT 490.2000 1403.4000 490.5000 1404.6000 ;
	    RECT 491.4000 1403.4000 492.6000 1404.6000 ;
	    RECT 493.8000 1403.7001 500.7000 1404.6000 ;
	    RECT 505.8000 1403.7001 509.7000 1404.9000 ;
	    RECT 510.6000 1403.7001 511.8000 1409.7001 ;
	    RECT 493.8000 1403.4000 495.0000 1403.7001 ;
	    RECT 469.2000 1398.0000 470.1000 1401.0000 ;
	    RECT 475.5000 1400.1000 476.7000 1401.9000 ;
	    RECT 471.0000 1398.9000 476.7000 1400.1000 ;
	    RECT 484.2000 1399.2001 485.4000 1403.4000 ;
	    RECT 496.2000 1402.5000 497.4000 1402.8000 ;
	    RECT 493.8000 1402.2001 495.0000 1402.5000 ;
	    RECT 488.4000 1401.3000 495.0000 1402.2001 ;
	    RECT 488.4000 1401.0000 489.6000 1401.3000 ;
	    RECT 496.2000 1400.4000 497.4000 1401.6000 ;
	    RECT 499.5000 1400.1000 500.7000 1403.7001 ;
	    RECT 508.5000 1402.8000 509.7000 1403.7001 ;
	    RECT 508.5000 1401.6000 513.0000 1402.8000 ;
	    RECT 515.4000 1400.7001 516.6000 1409.7001 ;
	    RECT 585.0000 1407.4501 586.2000 1407.6000 ;
	    RECT 645.0000 1407.4501 646.2000 1407.6000 ;
	    RECT 585.0000 1406.5500 646.2000 1407.4501 ;
	    RECT 585.0000 1406.4000 586.2000 1406.5500 ;
	    RECT 645.0000 1406.4000 646.2000 1406.5500 ;
	    RECT 489.0000 1398.9000 493.8000 1400.1000 ;
	    RECT 499.5000 1398.9000 502.5000 1400.1000 ;
	    RECT 503.4000 1399.5000 516.6000 1400.7001 ;
	    RECT 479.4000 1398.0000 480.6000 1398.9000 ;
	    RECT 469.2000 1397.1000 470.4000 1398.0000 ;
	    RECT 479.4000 1397.1000 504.9000 1398.0000 ;
	    RECT 505.8000 1397.4000 507.0000 1398.6000 ;
	    RECT 513.3000 1398.0000 514.5000 1398.3000 ;
	    RECT 507.9000 1397.1000 514.5000 1398.0000 ;
	    RECT 467.1000 1395.0000 468.6000 1396.2001 ;
	    RECT 467.4000 1393.5000 468.6000 1395.0000 ;
	    RECT 469.5000 1394.4000 470.4000 1397.1000 ;
	    RECT 471.3000 1396.2001 472.5000 1396.5000 ;
	    RECT 471.3000 1395.3000 509.7000 1396.2001 ;
	    RECT 505.5000 1395.0000 506.7000 1395.3000 ;
	    RECT 510.6000 1394.4000 511.8000 1395.6000 ;
	    RECT 469.5000 1393.5000 483.0000 1394.4000 ;
	    RECT 455.4000 1392.4501 456.6000 1392.6000 ;
	    RECT 467.4000 1392.4501 468.6000 1392.6000 ;
	    RECT 455.4000 1391.5500 468.6000 1392.4501 ;
	    RECT 455.4000 1391.4000 456.6000 1391.5500 ;
	    RECT 467.4000 1391.4000 468.6000 1391.5500 ;
	    RECT 469.5000 1391.1000 470.4000 1393.5000 ;
	    RECT 481.8000 1393.2001 483.0000 1393.5000 ;
	    RECT 486.6000 1393.5000 499.5000 1394.4000 ;
	    RECT 486.6000 1393.2001 487.8000 1393.5000 ;
	    RECT 474.3000 1391.4000 478.2000 1392.6000 ;
	    RECT 465.0000 1383.3000 466.2000 1389.3000 ;
	    RECT 467.4000 1383.3000 468.6000 1390.5000 ;
	    RECT 469.5000 1390.2001 473.4000 1391.1000 ;
	    RECT 469.8000 1383.3000 471.0000 1389.3000 ;
	    RECT 472.2000 1383.3000 473.4000 1390.2001 ;
	    RECT 474.6000 1383.3000 475.8000 1389.3000 ;
	    RECT 477.0000 1383.3000 478.2000 1391.4000 ;
	    RECT 479.1000 1390.2001 485.4000 1391.4000 ;
	    RECT 479.4000 1383.3000 480.6000 1389.3000 ;
	    RECT 481.8000 1383.3000 483.0000 1387.5000 ;
	    RECT 484.2000 1383.3000 485.4000 1387.5000 ;
	    RECT 486.6000 1383.3000 487.8000 1387.5000 ;
	    RECT 489.0000 1383.3000 490.2000 1392.6000 ;
	    RECT 493.8000 1391.4000 497.7000 1392.6000 ;
	    RECT 498.6000 1392.3000 499.5000 1393.5000 ;
	    RECT 501.0000 1394.1000 502.2000 1394.4000 ;
	    RECT 501.0000 1393.5000 509.1000 1394.1000 ;
	    RECT 501.0000 1393.2001 510.3000 1393.5000 ;
	    RECT 508.2000 1392.3000 510.3000 1393.2001 ;
	    RECT 498.6000 1391.4000 507.3000 1392.3000 ;
	    RECT 511.8000 1392.0000 514.2000 1393.2001 ;
	    RECT 511.8000 1391.4000 512.7000 1392.0000 ;
	    RECT 491.4000 1383.3000 492.6000 1389.3000 ;
	    RECT 493.8000 1383.3000 495.0000 1390.5000 ;
	    RECT 496.2000 1383.3000 497.4000 1389.3000 ;
	    RECT 498.6000 1383.3000 499.8000 1390.5000 ;
	    RECT 506.4000 1390.2001 512.7000 1391.4000 ;
	    RECT 515.4000 1391.1000 516.6000 1399.5000 ;
	    RECT 513.6000 1390.2001 516.6000 1391.1000 ;
	    RECT 647.4000 1400.7001 648.6000 1409.7001 ;
	    RECT 652.2000 1403.7001 653.4000 1409.7001 ;
	    RECT 657.0000 1404.9000 658.2000 1409.7001 ;
	    RECT 659.4000 1405.5000 660.6000 1409.7001 ;
	    RECT 661.8000 1405.5000 663.0000 1409.7001 ;
	    RECT 664.2000 1405.5000 665.4000 1409.7001 ;
	    RECT 666.6000 1406.7001 667.8000 1409.7001 ;
	    RECT 669.0000 1405.5000 670.2000 1409.7001 ;
	    RECT 671.4000 1406.7001 672.6000 1409.7001 ;
	    RECT 673.8000 1405.5000 675.0000 1409.7001 ;
	    RECT 676.2000 1405.5000 677.4000 1409.7001 ;
	    RECT 678.6000 1405.5000 679.8000 1409.7001 ;
	    RECT 681.0000 1405.5000 682.2000 1409.7001 ;
	    RECT 654.3000 1403.7001 658.2000 1404.9000 ;
	    RECT 683.4000 1404.9000 684.6000 1409.7001 ;
	    RECT 663.3000 1403.7001 670.2000 1404.6000 ;
	    RECT 654.3000 1402.8000 655.5000 1403.7001 ;
	    RECT 651.0000 1401.6000 655.5000 1402.8000 ;
	    RECT 647.4000 1399.5000 660.6000 1400.7001 ;
	    RECT 663.3000 1400.1000 664.5000 1403.7001 ;
	    RECT 669.0000 1403.4000 670.2000 1403.7001 ;
	    RECT 671.4000 1403.4000 672.6000 1404.6000 ;
	    RECT 673.5000 1403.4000 673.8000 1404.6000 ;
	    RECT 678.3000 1403.4000 679.8000 1404.6000 ;
	    RECT 683.4000 1403.7001 687.0000 1404.9000 ;
	    RECT 688.2000 1403.7001 689.4000 1409.7001 ;
	    RECT 666.6000 1402.5000 667.8000 1402.8000 ;
	    RECT 669.0000 1402.2001 670.2000 1402.5000 ;
	    RECT 666.6000 1400.4000 667.8000 1401.6000 ;
	    RECT 669.0000 1401.3000 675.6000 1402.2001 ;
	    RECT 674.4000 1401.0000 675.6000 1401.3000 ;
	    RECT 647.4000 1391.1000 648.6000 1399.5000 ;
	    RECT 661.5000 1398.9000 664.5000 1400.1000 ;
	    RECT 670.2000 1398.9000 675.0000 1400.1000 ;
	    RECT 678.6000 1399.2001 679.8000 1403.4000 ;
	    RECT 685.8000 1402.8000 687.0000 1403.7001 ;
	    RECT 685.8000 1401.9000 688.5000 1402.8000 ;
	    RECT 687.3000 1400.1000 688.5000 1401.9000 ;
	    RECT 693.0000 1401.9000 694.2000 1409.7001 ;
	    RECT 695.4000 1404.0000 696.6000 1409.7001 ;
	    RECT 697.8000 1406.7001 699.0000 1409.7001 ;
	    RECT 695.4000 1402.8000 696.9000 1404.0000 ;
	    RECT 724.2000 1403.7001 725.4000 1409.7001 ;
	    RECT 726.6000 1404.0000 727.8000 1409.7001 ;
	    RECT 729.0000 1404.9000 730.2000 1409.7001 ;
	    RECT 731.4000 1404.0000 732.6000 1409.7001 ;
	    RECT 726.6000 1403.7001 732.6000 1404.0000 ;
	    RECT 693.0000 1401.0000 694.8000 1401.9000 ;
	    RECT 687.3000 1398.9000 693.0000 1400.1000 ;
	    RECT 649.5000 1398.0000 650.7000 1398.3000 ;
	    RECT 649.5000 1397.1000 656.1000 1398.0000 ;
	    RECT 657.0000 1397.4000 658.2000 1398.6000 ;
	    RECT 683.4000 1398.0000 684.6000 1398.9000 ;
	    RECT 693.9000 1398.0000 694.8000 1401.0000 ;
	    RECT 659.1000 1397.1000 684.6000 1398.0000 ;
	    RECT 693.6000 1397.1000 694.8000 1398.0000 ;
	    RECT 691.5000 1396.2001 692.7000 1396.5000 ;
	    RECT 649.8000 1395.4501 651.0000 1395.6000 ;
	    RECT 652.2000 1395.4501 653.4000 1395.6000 ;
	    RECT 649.8000 1394.5500 653.4000 1395.4501 ;
	    RECT 654.3000 1395.3000 692.7000 1396.2001 ;
	    RECT 657.3000 1395.0000 658.5000 1395.3000 ;
	    RECT 649.8000 1394.4000 651.0000 1394.5500 ;
	    RECT 652.2000 1394.4000 653.4000 1394.5500 ;
	    RECT 693.6000 1394.4000 694.5000 1397.1000 ;
	    RECT 695.7000 1396.2001 696.9000 1402.8000 ;
	    RECT 724.5000 1402.5000 725.4000 1403.7001 ;
	    RECT 726.9000 1403.1000 732.3000 1403.7001 ;
	    RECT 743.4000 1402.5000 744.6000 1409.7001 ;
	    RECT 745.8000 1406.7001 747.0000 1409.7001 ;
	    RECT 745.8000 1405.5000 747.0000 1405.8000 ;
	    RECT 745.8000 1404.4501 747.0000 1404.6000 ;
	    RECT 755.4000 1404.4501 756.6000 1404.6000 ;
	    RECT 745.8000 1403.5500 756.6000 1404.4501 ;
	    RECT 745.8000 1403.4000 747.0000 1403.5500 ;
	    RECT 755.4000 1403.4000 756.6000 1403.5500 ;
	    RECT 760.2000 1402.5000 761.4000 1409.7001 ;
	    RECT 762.6000 1406.7001 763.8000 1409.7001 ;
	    RECT 762.6000 1405.5000 763.8000 1405.8000 ;
	    RECT 762.6000 1404.4501 763.8000 1404.6000 ;
	    RECT 882.6000 1404.4501 883.8000 1404.6000 ;
	    RECT 762.6000 1403.5500 883.8000 1404.4501 ;
	    RECT 762.6000 1403.4000 763.8000 1403.5500 ;
	    RECT 882.6000 1403.4000 883.8000 1403.5500 ;
	    RECT 724.2000 1400.4000 725.4000 1401.6000 ;
	    RECT 726.3000 1400.4000 728.1000 1401.6000 ;
	    RECT 730.2000 1400.7001 730.5000 1402.2001 ;
	    RECT 731.4000 1401.4501 732.6000 1401.6000 ;
	    RECT 741.0000 1401.4501 742.2000 1401.6000 ;
	    RECT 731.4000 1400.5500 742.2000 1401.4501 ;
	    RECT 731.4000 1400.4000 732.6000 1400.5500 ;
	    RECT 741.0000 1400.4000 742.2000 1400.5500 ;
	    RECT 743.4000 1400.4000 744.6000 1401.6000 ;
	    RECT 760.2000 1401.4501 761.4000 1401.6000 ;
	    RECT 803.4000 1401.4501 804.6000 1401.6000 ;
	    RECT 760.2000 1400.5500 804.6000 1401.4501 ;
	    RECT 760.2000 1400.4000 761.4000 1400.5500 ;
	    RECT 803.4000 1400.4000 804.6000 1400.5500 ;
	    RECT 894.6000 1400.7001 895.8000 1409.7001 ;
	    RECT 899.4000 1403.7001 900.6000 1409.7001 ;
	    RECT 904.2000 1404.9000 905.4000 1409.7001 ;
	    RECT 906.6000 1405.5000 907.8000 1409.7001 ;
	    RECT 909.0000 1405.5000 910.2000 1409.7001 ;
	    RECT 911.4000 1405.5000 912.6000 1409.7001 ;
	    RECT 913.8000 1406.7001 915.0000 1409.7001 ;
	    RECT 916.2000 1405.5000 917.4000 1409.7001 ;
	    RECT 918.6000 1406.7001 919.8000 1409.7001 ;
	    RECT 921.0000 1405.5000 922.2000 1409.7001 ;
	    RECT 923.4000 1405.5000 924.6000 1409.7001 ;
	    RECT 925.8000 1405.5000 927.0000 1409.7001 ;
	    RECT 928.2000 1405.5000 929.4000 1409.7001 ;
	    RECT 901.5000 1403.7001 905.4000 1404.9000 ;
	    RECT 930.6000 1404.9000 931.8000 1409.7001 ;
	    RECT 910.5000 1403.7001 917.4000 1404.6000 ;
	    RECT 901.5000 1402.8000 902.7000 1403.7001 ;
	    RECT 898.2000 1401.6000 902.7000 1402.8000 ;
	    RECT 661.8000 1394.1000 663.0000 1394.4000 ;
	    RECT 654.9000 1393.5000 663.0000 1394.1000 ;
	    RECT 653.7000 1393.2001 663.0000 1393.5000 ;
	    RECT 664.5000 1393.5000 677.4000 1394.4000 ;
	    RECT 649.8000 1392.0000 652.2000 1393.2001 ;
	    RECT 653.7000 1392.3000 655.8000 1393.2001 ;
	    RECT 664.5000 1392.3000 665.4000 1393.5000 ;
	    RECT 676.2000 1393.2001 677.4000 1393.5000 ;
	    RECT 681.0000 1393.5000 694.5000 1394.4000 ;
	    RECT 695.4000 1395.0000 696.9000 1396.2001 ;
	    RECT 695.4000 1393.5000 696.6000 1395.0000 ;
	    RECT 724.2000 1394.4000 725.4000 1395.6000 ;
	    RECT 727.2000 1395.3000 728.1000 1400.4000 ;
	    RECT 729.0000 1399.5000 730.2000 1399.8000 ;
	    RECT 894.6000 1399.5000 907.8000 1400.7001 ;
	    RECT 910.5000 1400.1000 911.7000 1403.7001 ;
	    RECT 916.2000 1403.4000 917.4000 1403.7001 ;
	    RECT 918.6000 1403.4000 919.8000 1404.6000 ;
	    RECT 920.7000 1403.4000 921.0000 1404.6000 ;
	    RECT 925.5000 1403.4000 927.0000 1404.6000 ;
	    RECT 930.6000 1403.7001 934.2000 1404.9000 ;
	    RECT 935.4000 1403.7001 936.6000 1409.7001 ;
	    RECT 913.8000 1402.5000 915.0000 1402.8000 ;
	    RECT 916.2000 1402.2001 917.4000 1402.5000 ;
	    RECT 913.8000 1400.4000 915.0000 1401.6000 ;
	    RECT 916.2000 1401.3000 922.8000 1402.2001 ;
	    RECT 921.6000 1401.0000 922.8000 1401.3000 ;
	    RECT 729.0000 1397.4000 730.2000 1398.6000 ;
	    RECT 727.2000 1394.4000 728.7000 1395.3000 ;
	    RECT 681.0000 1393.2001 682.2000 1393.5000 ;
	    RECT 651.3000 1391.4000 652.2000 1392.0000 ;
	    RECT 656.7000 1391.4000 665.4000 1392.3000 ;
	    RECT 666.3000 1391.4000 670.2000 1392.6000 ;
	    RECT 647.4000 1390.2001 650.4000 1391.1000 ;
	    RECT 651.3000 1390.2001 657.6000 1391.4000 ;
	    RECT 501.0000 1383.3000 502.2000 1387.5000 ;
	    RECT 503.4000 1383.3000 504.6000 1387.5000 ;
	    RECT 505.8000 1383.3000 507.0000 1389.3000 ;
	    RECT 508.2000 1383.3000 509.4000 1390.2001 ;
	    RECT 513.6000 1389.3000 514.5000 1390.2001 ;
	    RECT 649.5000 1389.3000 650.4000 1390.2001 ;
	    RECT 510.6000 1382.4000 511.8000 1389.3000 ;
	    RECT 513.0000 1388.4000 514.5000 1389.3000 ;
	    RECT 513.0000 1383.3000 514.2000 1388.4000 ;
	    RECT 515.4000 1383.3000 516.6000 1389.3000 ;
	    RECT 647.4000 1383.3000 648.6000 1389.3000 ;
	    RECT 649.5000 1388.4000 651.0000 1389.3000 ;
	    RECT 649.8000 1383.3000 651.0000 1388.4000 ;
	    RECT 652.2000 1382.4000 653.4000 1389.3000 ;
	    RECT 654.6000 1383.3000 655.8000 1390.2001 ;
	    RECT 657.0000 1383.3000 658.2000 1389.3000 ;
	    RECT 659.4000 1383.3000 660.6000 1387.5000 ;
	    RECT 661.8000 1383.3000 663.0000 1387.5000 ;
	    RECT 664.2000 1383.3000 665.4000 1390.5000 ;
	    RECT 666.6000 1383.3000 667.8000 1389.3000 ;
	    RECT 669.0000 1383.3000 670.2000 1390.5000 ;
	    RECT 671.4000 1383.3000 672.6000 1389.3000 ;
	    RECT 673.8000 1383.3000 675.0000 1392.6000 ;
	    RECT 685.8000 1391.4000 689.7000 1392.6000 ;
	    RECT 678.6000 1390.2001 684.9000 1391.4000 ;
	    RECT 676.2000 1383.3000 677.4000 1387.5000 ;
	    RECT 678.6000 1383.3000 679.8000 1387.5000 ;
	    RECT 681.0000 1383.3000 682.2000 1387.5000 ;
	    RECT 683.4000 1383.3000 684.6000 1389.3000 ;
	    RECT 685.8000 1383.3000 687.0000 1391.4000 ;
	    RECT 693.6000 1391.1000 694.5000 1393.5000 ;
	    RECT 725.4000 1392.6000 726.3000 1393.5000 ;
	    RECT 695.4000 1391.4000 696.6000 1392.6000 ;
	    RECT 725.4000 1391.4000 726.6000 1392.6000 ;
	    RECT 690.6000 1390.2001 694.5000 1391.1000 ;
	    RECT 688.2000 1383.3000 689.4000 1389.3000 ;
	    RECT 690.6000 1383.3000 691.8000 1390.2001 ;
	    RECT 693.0000 1383.3000 694.2000 1389.3000 ;
	    RECT 695.4000 1383.3000 696.6000 1390.5000 ;
	    RECT 697.8000 1383.3000 699.0000 1389.3000 ;
	    RECT 725.1000 1383.3000 726.3000 1389.3000 ;
	    RECT 727.5000 1383.3000 728.7000 1394.4000 ;
	    RECT 731.4000 1383.3000 732.6000 1395.3000 ;
	    RECT 743.4000 1383.3000 744.6000 1399.5000 ;
	    RECT 745.8000 1383.3000 747.0000 1389.3000 ;
	    RECT 760.2000 1383.3000 761.4000 1399.5000 ;
	    RECT 894.6000 1391.1000 895.8000 1399.5000 ;
	    RECT 908.7000 1398.9000 911.7000 1400.1000 ;
	    RECT 917.4000 1398.9000 922.2000 1400.1000 ;
	    RECT 925.8000 1399.2001 927.0000 1403.4000 ;
	    RECT 933.0000 1402.8000 934.2000 1403.7001 ;
	    RECT 933.0000 1401.9000 935.7000 1402.8000 ;
	    RECT 934.5000 1400.1000 935.7000 1401.9000 ;
	    RECT 940.2000 1401.9000 941.4000 1409.7001 ;
	    RECT 942.6000 1404.0000 943.8000 1409.7001 ;
	    RECT 945.0000 1406.7001 946.2000 1409.7001 ;
	    RECT 969.0000 1404.0000 970.2000 1409.7001 ;
	    RECT 971.4000 1404.9000 972.6000 1409.7001 ;
	    RECT 973.8000 1404.0000 975.0000 1409.7001 ;
	    RECT 942.6000 1402.8000 944.1000 1404.0000 ;
	    RECT 969.0000 1403.7001 975.0000 1404.0000 ;
	    RECT 976.2000 1403.7001 977.4000 1409.7001 ;
	    RECT 969.3000 1403.1000 974.7000 1403.7001 ;
	    RECT 940.2000 1401.0000 942.0000 1401.9000 ;
	    RECT 934.5000 1398.9000 940.2000 1400.1000 ;
	    RECT 896.7000 1398.0000 897.9000 1398.3000 ;
	    RECT 896.7000 1397.1000 903.3000 1398.0000 ;
	    RECT 904.2000 1397.4000 905.4000 1398.6000 ;
	    RECT 930.6000 1398.0000 931.8000 1398.9000 ;
	    RECT 941.1000 1398.0000 942.0000 1401.0000 ;
	    RECT 906.3000 1397.1000 931.8000 1398.0000 ;
	    RECT 940.8000 1397.1000 942.0000 1398.0000 ;
	    RECT 938.7000 1396.2001 939.9000 1396.5000 ;
	    RECT 899.4000 1394.4000 900.6000 1395.6000 ;
	    RECT 901.5000 1395.3000 939.9000 1396.2001 ;
	    RECT 904.5000 1395.0000 905.7000 1395.3000 ;
	    RECT 940.8000 1394.4000 941.7000 1397.1000 ;
	    RECT 942.9000 1396.2001 944.1000 1402.8000 ;
	    RECT 976.2000 1402.5000 977.1000 1403.7001 ;
	    RECT 990.6000 1402.5000 991.8000 1409.7001 ;
	    RECT 993.0000 1406.7001 994.2000 1409.7001 ;
	    RECT 993.0000 1405.5000 994.2000 1405.8000 ;
	    RECT 1013.1000 1404.6000 1014.3000 1409.7001 ;
	    RECT 993.0000 1403.4000 994.2000 1404.6000 ;
	    RECT 1013.1000 1403.7001 1015.8000 1404.6000 ;
	    RECT 1017.0000 1403.7001 1018.2000 1409.7001 ;
	    RECT 1031.4000 1406.7001 1032.6000 1409.7001 ;
	    RECT 1031.4000 1405.5000 1032.6000 1405.8000 ;
	    RECT 969.0000 1400.4000 970.2000 1401.6000 ;
	    RECT 971.1000 1400.7001 971.4000 1402.2001 ;
	    RECT 973.5000 1400.4000 975.3000 1401.6000 ;
	    RECT 976.2000 1400.4000 977.4000 1401.6000 ;
	    RECT 981.0000 1401.4501 982.2000 1401.6000 ;
	    RECT 990.6000 1401.4501 991.8000 1401.6000 ;
	    RECT 981.0000 1400.5500 991.8000 1401.4501 ;
	    RECT 981.0000 1400.4000 982.2000 1400.5500 ;
	    RECT 990.6000 1400.4000 991.8000 1400.5500 ;
	    RECT 971.4000 1399.5000 972.6000 1399.8000 ;
	    RECT 954.6000 1398.4501 955.8000 1398.6000 ;
	    RECT 971.4000 1398.4501 972.6000 1398.6000 ;
	    RECT 954.6000 1397.5500 972.6000 1398.4501 ;
	    RECT 954.6000 1397.4000 955.8000 1397.5500 ;
	    RECT 971.4000 1397.4000 972.6000 1397.5500 ;
	    RECT 909.0000 1394.1000 910.2000 1394.4000 ;
	    RECT 902.1000 1393.5000 910.2000 1394.1000 ;
	    RECT 900.9000 1393.2001 910.2000 1393.5000 ;
	    RECT 911.7000 1393.5000 924.6000 1394.4000 ;
	    RECT 897.0000 1392.0000 899.4000 1393.2001 ;
	    RECT 900.9000 1392.3000 903.0000 1393.2001 ;
	    RECT 911.7000 1392.3000 912.6000 1393.5000 ;
	    RECT 923.4000 1393.2001 924.6000 1393.5000 ;
	    RECT 928.2000 1393.5000 941.7000 1394.4000 ;
	    RECT 942.6000 1395.0000 944.1000 1396.2001 ;
	    RECT 973.5000 1395.3000 974.4000 1400.4000 ;
	    RECT 1014.6000 1399.5000 1015.8000 1403.7001 ;
	    RECT 1031.4000 1403.4000 1032.6000 1404.6000 ;
	    RECT 1017.0000 1402.5000 1018.2000 1402.8000 ;
	    RECT 1033.8000 1402.5000 1035.0000 1409.7001 ;
	    RECT 1057.8000 1403.7001 1059.0000 1409.7001 ;
	    RECT 1060.2001 1404.0000 1061.4000 1409.7001 ;
	    RECT 1062.6000 1404.9000 1063.8000 1409.7001 ;
	    RECT 1065.0000 1404.0000 1066.2001 1409.7001 ;
	    RECT 1060.2001 1403.7001 1066.2001 1404.0000 ;
	    RECT 1084.2001 1403.7001 1085.4000 1409.7001 ;
	    RECT 1088.1000 1404.6000 1089.3000 1409.7001 ;
	    RECT 1101.0000 1406.7001 1102.2001 1409.7001 ;
	    RECT 1101.0000 1405.5000 1102.2001 1405.8000 ;
	    RECT 1086.6000 1403.7001 1089.3000 1404.6000 ;
	    RECT 1091.4000 1404.4501 1092.6000 1404.6000 ;
	    RECT 1101.0000 1404.4501 1102.2001 1404.6000 ;
	    RECT 1058.1000 1402.5000 1059.0000 1403.7001 ;
	    RECT 1060.5000 1403.1000 1065.9000 1403.7001 ;
	    RECT 1084.2001 1402.5000 1085.4000 1402.8000 ;
	    RECT 1017.0000 1401.4501 1018.2000 1401.6000 ;
	    RECT 1019.4000 1401.4501 1020.6000 1401.6000 ;
	    RECT 1031.4000 1401.4501 1032.6000 1401.6000 ;
	    RECT 1017.0000 1400.5500 1032.6000 1401.4501 ;
	    RECT 1017.0000 1400.4000 1018.2000 1400.5500 ;
	    RECT 1019.4000 1400.4000 1020.6000 1400.5500 ;
	    RECT 1031.4000 1400.4000 1032.6000 1400.5500 ;
	    RECT 1033.8000 1401.4501 1035.0000 1401.6000 ;
	    RECT 1055.4000 1401.4501 1056.6000 1401.6000 ;
	    RECT 1033.8000 1400.5500 1056.6000 1401.4501 ;
	    RECT 1033.8000 1400.4000 1035.0000 1400.5500 ;
	    RECT 1055.4000 1400.4000 1056.6000 1400.5500 ;
	    RECT 1057.8000 1400.4000 1059.0000 1401.6000 ;
	    RECT 1059.9000 1400.4000 1061.7001 1401.6000 ;
	    RECT 1063.8000 1400.7001 1064.1000 1402.2001 ;
	    RECT 1065.0000 1401.4501 1066.2001 1401.6000 ;
	    RECT 1067.4000 1401.4501 1068.6000 1401.6000 ;
	    RECT 1065.0000 1400.5500 1068.6000 1401.4501 ;
	    RECT 1065.0000 1400.4000 1066.2001 1400.5500 ;
	    RECT 1067.4000 1400.4000 1068.6000 1400.5500 ;
	    RECT 1084.2001 1400.4000 1085.4000 1401.6000 ;
	    RECT 942.6000 1393.5000 943.8000 1395.0000 ;
	    RECT 928.2000 1393.2001 929.4000 1393.5000 ;
	    RECT 898.5000 1391.4000 899.4000 1392.0000 ;
	    RECT 903.9000 1391.4000 912.6000 1392.3000 ;
	    RECT 913.5000 1391.4000 917.4000 1392.6000 ;
	    RECT 894.6000 1390.2001 897.6000 1391.1000 ;
	    RECT 898.5000 1390.2001 904.8000 1391.4000 ;
	    RECT 896.7000 1389.3000 897.6000 1390.2001 ;
	    RECT 762.6000 1383.3000 763.8000 1389.3000 ;
	    RECT 894.6000 1383.3000 895.8000 1389.3000 ;
	    RECT 896.7000 1388.4000 898.2000 1389.3000 ;
	    RECT 897.0000 1383.3000 898.2000 1388.4000 ;
	    RECT 899.4000 1382.4000 900.6000 1389.3000 ;
	    RECT 901.8000 1383.3000 903.0000 1390.2001 ;
	    RECT 904.2000 1383.3000 905.4000 1389.3000 ;
	    RECT 906.6000 1383.3000 907.8000 1387.5000 ;
	    RECT 909.0000 1383.3000 910.2000 1387.5000 ;
	    RECT 911.4000 1383.3000 912.6000 1390.5000 ;
	    RECT 913.8000 1383.3000 915.0000 1389.3000 ;
	    RECT 916.2000 1383.3000 917.4000 1390.5000 ;
	    RECT 918.6000 1383.3000 919.8000 1389.3000 ;
	    RECT 921.0000 1383.3000 922.2000 1392.6000 ;
	    RECT 933.0000 1391.4000 936.9000 1392.6000 ;
	    RECT 925.8000 1390.2001 932.1000 1391.4000 ;
	    RECT 923.4000 1383.3000 924.6000 1387.5000 ;
	    RECT 925.8000 1383.3000 927.0000 1387.5000 ;
	    RECT 928.2000 1383.3000 929.4000 1387.5000 ;
	    RECT 930.6000 1383.3000 931.8000 1389.3000 ;
	    RECT 933.0000 1383.3000 934.2000 1391.4000 ;
	    RECT 940.8000 1391.1000 941.7000 1393.5000 ;
	    RECT 942.6000 1391.4000 943.8000 1392.6000 ;
	    RECT 937.8000 1390.2001 941.7000 1391.1000 ;
	    RECT 935.4000 1383.3000 936.6000 1389.3000 ;
	    RECT 937.8000 1383.3000 939.0000 1390.2001 ;
	    RECT 940.2000 1383.3000 941.4000 1389.3000 ;
	    RECT 942.6000 1383.3000 943.8000 1390.5000 ;
	    RECT 945.0000 1383.3000 946.2000 1389.3000 ;
	    RECT 969.0000 1383.3000 970.2000 1395.3000 ;
	    RECT 972.9000 1394.4000 974.4000 1395.3000 ;
	    RECT 976.2000 1394.4000 977.4000 1395.6000 ;
	    RECT 972.9000 1383.3000 974.1000 1394.4000 ;
	    RECT 975.3000 1392.6000 976.2000 1393.5000 ;
	    RECT 975.0000 1391.4000 976.2000 1392.6000 ;
	    RECT 975.3000 1383.3000 976.5000 1389.3000 ;
	    RECT 990.6000 1383.3000 991.8000 1399.5000 ;
	    RECT 993.0000 1398.4501 994.2000 1398.6000 ;
	    RECT 1014.6000 1398.4501 1015.8000 1398.6000 ;
	    RECT 993.0000 1397.5500 1015.8000 1398.4501 ;
	    RECT 993.0000 1397.4000 994.2000 1397.5500 ;
	    RECT 1014.6000 1397.4000 1015.8000 1397.5500 ;
	    RECT 1012.2000 1394.4000 1013.4000 1395.6000 ;
	    RECT 1012.2000 1393.2001 1013.4000 1393.5000 ;
	    RECT 993.0000 1383.3000 994.2000 1389.3000 ;
	    RECT 1012.2000 1383.3000 1013.4000 1389.3000 ;
	    RECT 1014.6000 1383.3000 1015.8000 1396.5000 ;
	    RECT 1017.0000 1383.3000 1018.2000 1389.3000 ;
	    RECT 1031.4000 1383.3000 1032.6000 1389.3000 ;
	    RECT 1033.8000 1383.3000 1035.0000 1399.5000 ;
	    RECT 1057.8000 1394.4000 1059.0000 1395.6000 ;
	    RECT 1060.8000 1395.3000 1061.7001 1400.4000 ;
	    RECT 1062.6000 1399.5000 1063.8000 1399.8000 ;
	    RECT 1086.6000 1399.5000 1087.8000 1403.7001 ;
	    RECT 1091.4000 1403.5500 1102.2001 1404.4501 ;
	    RECT 1091.4000 1403.4000 1092.6000 1403.5500 ;
	    RECT 1101.0000 1403.4000 1102.2001 1403.5500 ;
	    RECT 1103.4000 1402.5000 1104.6000 1409.7001 ;
	    RECT 1123.5000 1404.6000 1124.7001 1409.7001 ;
	    RECT 1123.5000 1403.7001 1126.2001 1404.6000 ;
	    RECT 1127.4000 1403.7001 1128.6000 1409.7001 ;
	    RECT 1261.8000 1406.7001 1263.0000 1409.7001 ;
	    RECT 1264.2001 1404.0000 1265.4000 1409.7001 ;
	    RECT 1103.4000 1401.4501 1104.6000 1401.6000 ;
	    RECT 1122.6000 1401.4501 1123.8000 1401.6000 ;
	    RECT 1103.4000 1400.5500 1123.8000 1401.4501 ;
	    RECT 1103.4000 1400.4000 1104.6000 1400.5500 ;
	    RECT 1122.6000 1400.4000 1123.8000 1400.5500 ;
	    RECT 1125.0000 1399.5000 1126.2001 1403.7001 ;
	    RECT 1263.9000 1402.8000 1265.4000 1404.0000 ;
	    RECT 1127.4000 1402.5000 1128.6000 1402.8000 ;
	    RECT 1127.4000 1400.4000 1128.6000 1401.6000 ;
	    RECT 1062.6000 1397.4000 1063.8000 1398.6000 ;
	    RECT 1065.0000 1398.4501 1066.2001 1398.6000 ;
	    RECT 1086.6000 1398.4501 1087.8000 1398.6000 ;
	    RECT 1065.0000 1397.5500 1087.8000 1398.4501 ;
	    RECT 1065.0000 1397.4000 1066.2001 1397.5500 ;
	    RECT 1086.6000 1397.4000 1087.8000 1397.5500 ;
	    RECT 1060.8000 1394.4000 1062.3000 1395.3000 ;
	    RECT 1059.0000 1392.6000 1059.9000 1393.5000 ;
	    RECT 1059.0000 1391.4000 1060.2001 1392.6000 ;
	    RECT 1058.7001 1383.3000 1059.9000 1389.3000 ;
	    RECT 1061.1000 1383.3000 1062.3000 1394.4000 ;
	    RECT 1065.0000 1383.3000 1066.2001 1395.3000 ;
	    RECT 1084.2001 1383.3000 1085.4000 1389.3000 ;
	    RECT 1086.6000 1383.3000 1087.8000 1396.5000 ;
	    RECT 1089.0000 1394.4000 1090.2001 1395.6000 ;
	    RECT 1089.0000 1393.2001 1090.2001 1393.5000 ;
	    RECT 1089.0000 1383.3000 1090.2001 1389.3000 ;
	    RECT 1101.0000 1383.3000 1102.2001 1389.3000 ;
	    RECT 1103.4000 1383.3000 1104.6000 1399.5000 ;
	    RECT 1125.0000 1398.4501 1126.2001 1398.6000 ;
	    RECT 1137.0000 1398.4501 1138.2001 1398.6000 ;
	    RECT 1125.0000 1397.5500 1138.2001 1398.4501 ;
	    RECT 1125.0000 1397.4000 1126.2001 1397.5500 ;
	    RECT 1137.0000 1397.4000 1138.2001 1397.5500 ;
	    RECT 1120.2001 1395.4501 1121.4000 1395.6000 ;
	    RECT 1122.6000 1395.4501 1123.8000 1395.6000 ;
	    RECT 1120.2001 1394.5500 1123.8000 1395.4501 ;
	    RECT 1120.2001 1394.4000 1121.4000 1394.5500 ;
	    RECT 1122.6000 1394.4000 1123.8000 1394.5500 ;
	    RECT 1122.6000 1393.2001 1123.8000 1393.5000 ;
	    RECT 1122.6000 1383.3000 1123.8000 1389.3000 ;
	    RECT 1125.0000 1383.3000 1126.2001 1396.5000 ;
	    RECT 1263.9000 1396.2001 1265.1000 1402.8000 ;
	    RECT 1266.6000 1401.9000 1267.8000 1409.7001 ;
	    RECT 1271.4000 1403.7001 1272.6000 1409.7001 ;
	    RECT 1276.2001 1404.9000 1277.4000 1409.7001 ;
	    RECT 1278.6000 1405.5000 1279.8000 1409.7001 ;
	    RECT 1281.0000 1405.5000 1282.2001 1409.7001 ;
	    RECT 1283.4000 1405.5000 1284.6000 1409.7001 ;
	    RECT 1285.8000 1405.5000 1287.0000 1409.7001 ;
	    RECT 1288.2001 1406.7001 1289.4000 1409.7001 ;
	    RECT 1290.6000 1405.5000 1291.8000 1409.7001 ;
	    RECT 1293.0000 1406.7001 1294.2001 1409.7001 ;
	    RECT 1295.4000 1405.5000 1296.6000 1409.7001 ;
	    RECT 1297.8000 1405.5000 1299.0000 1409.7001 ;
	    RECT 1300.2001 1405.5000 1301.4000 1409.7001 ;
	    RECT 1273.8000 1403.7001 1277.4000 1404.9000 ;
	    RECT 1302.6000 1404.9000 1303.8000 1409.7001 ;
	    RECT 1273.8000 1402.8000 1275.0000 1403.7001 ;
	    RECT 1266.0000 1401.0000 1267.8000 1401.9000 ;
	    RECT 1272.3000 1401.9000 1275.0000 1402.8000 ;
	    RECT 1281.0000 1403.4000 1282.5000 1404.6000 ;
	    RECT 1287.0000 1403.4000 1287.3000 1404.6000 ;
	    RECT 1288.2001 1403.4000 1289.4000 1404.6000 ;
	    RECT 1290.6000 1403.7001 1297.5000 1404.6000 ;
	    RECT 1302.6000 1403.7001 1306.5000 1404.9000 ;
	    RECT 1307.4000 1403.7001 1308.6000 1409.7001 ;
	    RECT 1290.6000 1403.4000 1291.8000 1403.7001 ;
	    RECT 1266.0000 1398.0000 1266.9000 1401.0000 ;
	    RECT 1272.3000 1400.1000 1273.5000 1401.9000 ;
	    RECT 1267.8000 1398.9000 1273.5000 1400.1000 ;
	    RECT 1281.0000 1399.2001 1282.2001 1403.4000 ;
	    RECT 1293.0000 1402.5000 1294.2001 1402.8000 ;
	    RECT 1290.6000 1402.2001 1291.8000 1402.5000 ;
	    RECT 1285.2001 1401.3000 1291.8000 1402.2001 ;
	    RECT 1285.2001 1401.0000 1286.4000 1401.3000 ;
	    RECT 1293.0000 1400.4000 1294.2001 1401.6000 ;
	    RECT 1296.3000 1400.1000 1297.5000 1403.7001 ;
	    RECT 1305.3000 1402.8000 1306.5000 1403.7001 ;
	    RECT 1305.3000 1401.6000 1309.8000 1402.8000 ;
	    RECT 1312.2001 1400.7001 1313.4000 1409.7001 ;
	    RECT 1338.6000 1404.0000 1339.8000 1409.7001 ;
	    RECT 1341.0000 1404.9000 1342.2001 1409.7001 ;
	    RECT 1343.4000 1404.0000 1344.6000 1409.7001 ;
	    RECT 1338.6000 1403.7001 1344.6000 1404.0000 ;
	    RECT 1345.8000 1403.7001 1347.0000 1409.7001 ;
	    RECT 1377.0000 1404.0000 1378.2001 1409.7001 ;
	    RECT 1379.4000 1404.9000 1380.6000 1409.7001 ;
	    RECT 1381.8000 1404.0000 1383.0000 1409.7001 ;
	    RECT 1377.0000 1403.7001 1383.0000 1404.0000 ;
	    RECT 1384.2001 1403.7001 1385.4000 1409.7001 ;
	    RECT 1338.9000 1403.1000 1344.3000 1403.7001 ;
	    RECT 1345.8000 1402.5000 1346.7001 1403.7001 ;
	    RECT 1377.3000 1403.1000 1382.7001 1403.7001 ;
	    RECT 1384.2001 1402.5000 1385.1000 1403.7001 ;
	    RECT 1285.8000 1398.9000 1290.6000 1400.1000 ;
	    RECT 1296.3000 1398.9000 1299.3000 1400.1000 ;
	    RECT 1300.2001 1399.5000 1313.4000 1400.7001 ;
	    RECT 1314.6000 1401.4501 1315.8000 1401.6000 ;
	    RECT 1338.6000 1401.4501 1339.8000 1401.6000 ;
	    RECT 1314.6000 1400.5500 1339.8000 1401.4501 ;
	    RECT 1340.7001 1400.7001 1341.0000 1402.2001 ;
	    RECT 1314.6000 1400.4000 1315.8000 1400.5500 ;
	    RECT 1338.6000 1400.4000 1339.8000 1400.5500 ;
	    RECT 1343.1000 1400.4000 1344.9000 1401.6000 ;
	    RECT 1345.8000 1401.4501 1347.0000 1401.6000 ;
	    RECT 1348.2001 1401.4501 1349.4000 1401.6000 ;
	    RECT 1345.8000 1400.5500 1349.4000 1401.4501 ;
	    RECT 1345.8000 1400.4000 1347.0000 1400.5500 ;
	    RECT 1348.2001 1400.4000 1349.4000 1400.5500 ;
	    RECT 1377.0000 1400.4000 1378.2001 1401.6000 ;
	    RECT 1379.1000 1400.7001 1379.4000 1402.2001 ;
	    RECT 1381.5000 1400.4000 1383.3000 1401.6000 ;
	    RECT 1384.2001 1401.4501 1385.4000 1401.6000 ;
	    RECT 1485.0000 1401.4501 1486.2001 1401.6000 ;
	    RECT 1384.2001 1400.5500 1486.2001 1401.4501 ;
	    RECT 1384.2001 1400.4000 1385.4000 1400.5500 ;
	    RECT 1485.0000 1400.4000 1486.2001 1400.5500 ;
	    RECT 1511.4000 1400.7001 1512.6000 1409.7001 ;
	    RECT 1516.2001 1403.7001 1517.4000 1409.7001 ;
	    RECT 1521.0000 1404.9000 1522.2001 1409.7001 ;
	    RECT 1523.4000 1405.5000 1524.6000 1409.7001 ;
	    RECT 1525.8000 1405.5000 1527.0000 1409.7001 ;
	    RECT 1528.2001 1405.5000 1529.4000 1409.7001 ;
	    RECT 1530.6000 1406.7001 1531.8000 1409.7001 ;
	    RECT 1533.0000 1405.5000 1534.2001 1409.7001 ;
	    RECT 1535.4000 1406.7001 1536.6000 1409.7001 ;
	    RECT 1537.8000 1405.5000 1539.0000 1409.7001 ;
	    RECT 1540.2001 1405.5000 1541.4000 1409.7001 ;
	    RECT 1542.6000 1405.5000 1543.8000 1409.7001 ;
	    RECT 1545.0000 1405.5000 1546.2001 1409.7001 ;
	    RECT 1518.3000 1403.7001 1522.2001 1404.9000 ;
	    RECT 1547.4000 1404.9000 1548.6000 1409.7001 ;
	    RECT 1527.3000 1403.7001 1534.2001 1404.6000 ;
	    RECT 1518.3000 1402.8000 1519.5000 1403.7001 ;
	    RECT 1515.0000 1401.6000 1519.5000 1402.8000 ;
	    RECT 1341.0000 1399.5000 1342.2001 1399.8000 ;
	    RECT 1276.2001 1398.0000 1277.4000 1398.9000 ;
	    RECT 1266.0000 1397.1000 1267.2001 1398.0000 ;
	    RECT 1276.2001 1397.1000 1301.7001 1398.0000 ;
	    RECT 1302.6000 1397.4000 1303.8000 1398.6000 ;
	    RECT 1310.1000 1398.0000 1311.3000 1398.3000 ;
	    RECT 1304.7001 1397.1000 1311.3000 1398.0000 ;
	    RECT 1263.9000 1395.0000 1265.4000 1396.2001 ;
	    RECT 1264.2001 1393.5000 1265.4000 1395.0000 ;
	    RECT 1266.3000 1394.4000 1267.2001 1397.1000 ;
	    RECT 1268.1000 1396.2001 1269.3000 1396.5000 ;
	    RECT 1268.1000 1395.3000 1306.5000 1396.2001 ;
	    RECT 1302.3000 1395.0000 1303.5000 1395.3000 ;
	    RECT 1307.4000 1394.4000 1308.6000 1395.6000 ;
	    RECT 1266.3000 1393.5000 1279.8000 1394.4000 ;
	    RECT 1127.4000 1392.4501 1128.6000 1392.6000 ;
	    RECT 1264.2001 1392.4501 1265.4000 1392.6000 ;
	    RECT 1127.4000 1391.5500 1265.4000 1392.4501 ;
	    RECT 1127.4000 1391.4000 1128.6000 1391.5500 ;
	    RECT 1264.2001 1391.4000 1265.4000 1391.5500 ;
	    RECT 1266.3000 1391.1000 1267.2001 1393.5000 ;
	    RECT 1278.6000 1393.2001 1279.8000 1393.5000 ;
	    RECT 1283.4000 1393.5000 1296.3000 1394.4000 ;
	    RECT 1283.4000 1393.2001 1284.6000 1393.5000 ;
	    RECT 1271.1000 1391.4000 1275.0000 1392.6000 ;
	    RECT 1127.4000 1383.3000 1128.6000 1389.3000 ;
	    RECT 1261.8000 1383.3000 1263.0000 1389.3000 ;
	    RECT 1264.2001 1383.3000 1265.4000 1390.5000 ;
	    RECT 1266.3000 1390.2001 1270.2001 1391.1000 ;
	    RECT 1266.6000 1383.3000 1267.8000 1389.3000 ;
	    RECT 1269.0000 1383.3000 1270.2001 1390.2001 ;
	    RECT 1271.4000 1383.3000 1272.6000 1389.3000 ;
	    RECT 1273.8000 1383.3000 1275.0000 1391.4000 ;
	    RECT 1275.9000 1390.2001 1282.2001 1391.4000 ;
	    RECT 1276.2001 1383.3000 1277.4000 1389.3000 ;
	    RECT 1278.6000 1383.3000 1279.8000 1387.5000 ;
	    RECT 1281.0000 1383.3000 1282.2001 1387.5000 ;
	    RECT 1283.4000 1383.3000 1284.6000 1387.5000 ;
	    RECT 1285.8000 1383.3000 1287.0000 1392.6000 ;
	    RECT 1290.6000 1391.4000 1294.5000 1392.6000 ;
	    RECT 1295.4000 1392.3000 1296.3000 1393.5000 ;
	    RECT 1297.8000 1394.1000 1299.0000 1394.4000 ;
	    RECT 1297.8000 1393.5000 1305.9000 1394.1000 ;
	    RECT 1297.8000 1393.2001 1307.1000 1393.5000 ;
	    RECT 1305.0000 1392.3000 1307.1000 1393.2001 ;
	    RECT 1295.4000 1391.4000 1304.1000 1392.3000 ;
	    RECT 1308.6000 1392.0000 1311.0000 1393.2001 ;
	    RECT 1308.6000 1391.4000 1309.5000 1392.0000 ;
	    RECT 1288.2001 1383.3000 1289.4000 1389.3000 ;
	    RECT 1290.6000 1383.3000 1291.8000 1390.5000 ;
	    RECT 1293.0000 1383.3000 1294.2001 1389.3000 ;
	    RECT 1295.4000 1383.3000 1296.6000 1390.5000 ;
	    RECT 1303.2001 1390.2001 1309.5000 1391.4000 ;
	    RECT 1312.2001 1391.1000 1313.4000 1399.5000 ;
	    RECT 1341.0000 1397.4000 1342.2001 1398.6000 ;
	    RECT 1343.1000 1395.3000 1344.0000 1400.4000 ;
	    RECT 1379.4000 1399.5000 1380.6000 1399.8000 ;
	    RECT 1374.6000 1398.4501 1375.8000 1398.6000 ;
	    RECT 1379.4000 1398.4501 1380.6000 1398.6000 ;
	    RECT 1374.6000 1397.5500 1380.6000 1398.4501 ;
	    RECT 1374.6000 1397.4000 1375.8000 1397.5500 ;
	    RECT 1379.4000 1397.4000 1380.6000 1397.5500 ;
	    RECT 1310.4000 1390.2001 1313.4000 1391.1000 ;
	    RECT 1297.8000 1383.3000 1299.0000 1387.5000 ;
	    RECT 1300.2001 1383.3000 1301.4000 1387.5000 ;
	    RECT 1302.6000 1383.3000 1303.8000 1389.3000 ;
	    RECT 1305.0000 1383.3000 1306.2001 1390.2001 ;
	    RECT 1310.4000 1389.3000 1311.3000 1390.2001 ;
	    RECT 1307.4000 1382.4000 1308.6000 1389.3000 ;
	    RECT 1309.8000 1388.4000 1311.3000 1389.3000 ;
	    RECT 1309.8000 1383.3000 1311.0000 1388.4000 ;
	    RECT 1312.2001 1383.3000 1313.4000 1389.3000 ;
	    RECT 1338.6000 1383.3000 1339.8000 1395.3000 ;
	    RECT 1342.5000 1394.4000 1344.0000 1395.3000 ;
	    RECT 1345.8000 1394.4000 1347.0000 1395.6000 ;
	    RECT 1381.5000 1395.3000 1382.4000 1400.4000 ;
	    RECT 1511.4000 1399.5000 1524.6000 1400.7001 ;
	    RECT 1527.3000 1400.1000 1528.5000 1403.7001 ;
	    RECT 1533.0000 1403.4000 1534.2001 1403.7001 ;
	    RECT 1535.4000 1403.4000 1536.6000 1404.6000 ;
	    RECT 1537.5000 1403.4000 1537.8000 1404.6000 ;
	    RECT 1542.3000 1403.4000 1543.8000 1404.6000 ;
	    RECT 1547.4000 1403.7001 1551.0000 1404.9000 ;
	    RECT 1552.2001 1403.7001 1553.4000 1409.7001 ;
	    RECT 1530.6000 1402.5000 1531.8000 1402.8000 ;
	    RECT 1533.0000 1402.2001 1534.2001 1402.5000 ;
	    RECT 1530.6000 1400.4000 1531.8000 1401.6000 ;
	    RECT 1533.0000 1401.3000 1539.6000 1402.2001 ;
	    RECT 1538.4000 1401.0000 1539.6000 1401.3000 ;
	    RECT 1342.5000 1383.3000 1343.7001 1394.4000 ;
	    RECT 1344.9000 1392.6000 1345.8000 1393.5000 ;
	    RECT 1344.6000 1391.4000 1345.8000 1392.6000 ;
	    RECT 1344.9000 1383.3000 1346.1000 1389.3000 ;
	    RECT 1377.0000 1383.3000 1378.2001 1395.3000 ;
	    RECT 1380.9000 1394.4000 1382.4000 1395.3000 ;
	    RECT 1384.2001 1394.4000 1385.4000 1395.6000 ;
	    RECT 1380.9000 1383.3000 1382.1000 1394.4000 ;
	    RECT 1383.3000 1392.6000 1384.2001 1393.5000 ;
	    RECT 1383.0000 1391.4000 1384.2001 1392.6000 ;
	    RECT 1511.4000 1391.1000 1512.6000 1399.5000 ;
	    RECT 1525.5000 1398.9000 1528.5000 1400.1000 ;
	    RECT 1534.2001 1398.9000 1539.0000 1400.1000 ;
	    RECT 1542.6000 1399.2001 1543.8000 1403.4000 ;
	    RECT 1549.8000 1402.8000 1551.0000 1403.7001 ;
	    RECT 1549.8000 1401.9000 1552.5000 1402.8000 ;
	    RECT 1551.3000 1400.1000 1552.5000 1401.9000 ;
	    RECT 1557.0000 1401.9000 1558.2001 1409.7001 ;
	    RECT 1559.4000 1404.0000 1560.6000 1409.7001 ;
	    RECT 1561.8000 1406.7001 1563.0000 1409.7001 ;
	    RECT 1559.4000 1402.8000 1560.9000 1404.0000 ;
	    RECT 1557.0000 1401.0000 1558.8000 1401.9000 ;
	    RECT 1551.3000 1398.9000 1557.0000 1400.1000 ;
	    RECT 1513.5000 1398.0000 1514.7001 1398.3000 ;
	    RECT 1513.5000 1397.1000 1520.1000 1398.0000 ;
	    RECT 1521.0000 1397.4000 1522.2001 1398.6000 ;
	    RECT 1547.4000 1398.0000 1548.6000 1398.9000 ;
	    RECT 1557.9000 1398.0000 1558.8000 1401.0000 ;
	    RECT 1523.1000 1397.1000 1548.6000 1398.0000 ;
	    RECT 1557.6000 1397.1000 1558.8000 1398.0000 ;
	    RECT 1555.5000 1396.2001 1556.7001 1396.5000 ;
	    RECT 1516.2001 1394.4000 1517.4000 1395.6000 ;
	    RECT 1518.3000 1395.3000 1556.7001 1396.2001 ;
	    RECT 1521.3000 1395.0000 1522.5000 1395.3000 ;
	    RECT 1557.6000 1394.4000 1558.5000 1397.1000 ;
	    RECT 1559.7001 1396.2001 1560.9000 1402.8000 ;
	    RECT 1525.8000 1394.1000 1527.0000 1394.4000 ;
	    RECT 1518.9000 1393.5000 1527.0000 1394.1000 ;
	    RECT 1517.7001 1393.2001 1527.0000 1393.5000 ;
	    RECT 1528.5000 1393.5000 1541.4000 1394.4000 ;
	    RECT 1513.8000 1392.0000 1516.2001 1393.2001 ;
	    RECT 1517.7001 1392.3000 1519.8000 1393.2001 ;
	    RECT 1528.5000 1392.3000 1529.4000 1393.5000 ;
	    RECT 1540.2001 1393.2001 1541.4000 1393.5000 ;
	    RECT 1545.0000 1393.5000 1558.5000 1394.4000 ;
	    RECT 1559.4000 1395.0000 1560.9000 1396.2001 ;
	    RECT 1559.4000 1393.5000 1560.6000 1395.0000 ;
	    RECT 1545.0000 1393.2001 1546.2001 1393.5000 ;
	    RECT 1515.3000 1391.4000 1516.2001 1392.0000 ;
	    RECT 1520.7001 1391.4000 1529.4000 1392.3000 ;
	    RECT 1530.3000 1391.4000 1534.2001 1392.6000 ;
	    RECT 1511.4000 1390.2001 1514.4000 1391.1000 ;
	    RECT 1515.3000 1390.2001 1521.6000 1391.4000 ;
	    RECT 1513.5000 1389.3000 1514.4000 1390.2001 ;
	    RECT 1383.3000 1383.3000 1384.5000 1389.3000 ;
	    RECT 1451.4000 1386.4501 1452.6000 1386.6000 ;
	    RECT 1506.6000 1386.4501 1507.8000 1386.6000 ;
	    RECT 1451.4000 1385.5500 1507.8000 1386.4501 ;
	    RECT 1451.4000 1385.4000 1452.6000 1385.5500 ;
	    RECT 1506.6000 1385.4000 1507.8000 1385.5500 ;
	    RECT 1511.4000 1383.3000 1512.6000 1389.3000 ;
	    RECT 1513.5000 1388.4000 1515.0000 1389.3000 ;
	    RECT 1513.8000 1383.3000 1515.0000 1388.4000 ;
	    RECT 1516.2001 1382.4000 1517.4000 1389.3000 ;
	    RECT 1518.6000 1383.3000 1519.8000 1390.2001 ;
	    RECT 1521.0000 1383.3000 1522.2001 1389.3000 ;
	    RECT 1523.4000 1383.3000 1524.6000 1387.5000 ;
	    RECT 1525.8000 1383.3000 1527.0000 1387.5000 ;
	    RECT 1528.2001 1383.3000 1529.4000 1390.5000 ;
	    RECT 1530.6000 1383.3000 1531.8000 1389.3000 ;
	    RECT 1533.0000 1383.3000 1534.2001 1390.5000 ;
	    RECT 1535.4000 1383.3000 1536.6000 1389.3000 ;
	    RECT 1537.8000 1383.3000 1539.0000 1392.6000 ;
	    RECT 1549.8000 1391.4000 1553.7001 1392.6000 ;
	    RECT 1542.6000 1390.2001 1548.9000 1391.4000 ;
	    RECT 1540.2001 1383.3000 1541.4000 1387.5000 ;
	    RECT 1542.6000 1383.3000 1543.8000 1387.5000 ;
	    RECT 1545.0000 1383.3000 1546.2001 1387.5000 ;
	    RECT 1547.4000 1383.3000 1548.6000 1389.3000 ;
	    RECT 1549.8000 1383.3000 1551.0000 1391.4000 ;
	    RECT 1557.6000 1391.1000 1558.5000 1393.5000 ;
	    RECT 1559.4000 1391.4000 1560.6000 1392.6000 ;
	    RECT 1554.6000 1390.2001 1558.5000 1391.1000 ;
	    RECT 1552.2001 1383.3000 1553.4000 1389.3000 ;
	    RECT 1554.6000 1383.3000 1555.8000 1390.2001 ;
	    RECT 1557.0000 1383.3000 1558.2001 1389.3000 ;
	    RECT 1559.4000 1383.3000 1560.6000 1390.5000 ;
	    RECT 1561.8000 1383.3000 1563.0000 1389.3000 ;
	    RECT 1.2000 1380.6000 1569.0000 1382.4000 ;
	    RECT 126.6000 1373.7001 127.8000 1379.7001 ;
	    RECT 129.0000 1374.6000 130.2000 1379.7001 ;
	    RECT 128.7000 1373.7001 130.2000 1374.6000 ;
	    RECT 131.4000 1373.7001 132.6000 1380.6000 ;
	    RECT 128.7000 1372.8000 129.6000 1373.7001 ;
	    RECT 133.8000 1372.8000 135.0000 1379.7001 ;
	    RECT 136.2000 1373.7001 137.4000 1379.7001 ;
	    RECT 138.6000 1375.5000 139.8000 1379.7001 ;
	    RECT 141.0000 1375.5000 142.2000 1379.7001 ;
	    RECT 126.6000 1371.9000 129.6000 1372.8000 ;
	    RECT 126.6000 1363.5000 127.8000 1371.9000 ;
	    RECT 130.5000 1371.6000 136.8000 1372.8000 ;
	    RECT 143.4000 1372.5000 144.6000 1379.7001 ;
	    RECT 145.8000 1373.7001 147.0000 1379.7001 ;
	    RECT 148.2000 1372.5000 149.4000 1379.7001 ;
	    RECT 150.6000 1373.7001 151.8000 1379.7001 ;
	    RECT 130.5000 1371.0000 131.4000 1371.6000 ;
	    RECT 129.0000 1369.8000 131.4000 1371.0000 ;
	    RECT 135.9000 1370.7001 144.6000 1371.6000 ;
	    RECT 132.9000 1369.8000 135.0000 1370.7001 ;
	    RECT 132.9000 1369.5000 142.2000 1369.8000 ;
	    RECT 134.1000 1368.9000 142.2000 1369.5000 ;
	    RECT 141.0000 1368.6000 142.2000 1368.9000 ;
	    RECT 143.7000 1369.5000 144.6000 1370.7001 ;
	    RECT 145.5000 1370.4000 149.4000 1371.6000 ;
	    RECT 153.0000 1370.4000 154.2000 1379.7001 ;
	    RECT 155.4000 1375.5000 156.6000 1379.7001 ;
	    RECT 157.8000 1375.5000 159.0000 1379.7001 ;
	    RECT 160.2000 1375.5000 161.4000 1379.7001 ;
	    RECT 162.6000 1373.7001 163.8000 1379.7001 ;
	    RECT 157.8000 1371.6000 164.1000 1372.8000 ;
	    RECT 165.0000 1371.6000 166.2000 1379.7001 ;
	    RECT 167.4000 1373.7001 168.6000 1379.7001 ;
	    RECT 169.8000 1372.8000 171.0000 1379.7001 ;
	    RECT 172.2000 1373.7001 173.4000 1379.7001 ;
	    RECT 169.8000 1371.9000 173.7000 1372.8000 ;
	    RECT 174.6000 1372.5000 175.8000 1379.7001 ;
	    RECT 177.0000 1373.7001 178.2000 1379.7001 ;
	    RECT 191.4000 1373.7001 192.6000 1379.7001 ;
	    RECT 165.0000 1370.4000 168.9000 1371.6000 ;
	    RECT 155.4000 1369.5000 156.6000 1369.8000 ;
	    RECT 143.7000 1368.6000 156.6000 1369.5000 ;
	    RECT 160.2000 1369.5000 161.4000 1369.8000 ;
	    RECT 172.8000 1369.5000 173.7000 1371.9000 ;
	    RECT 174.6000 1371.4501 175.8000 1371.6000 ;
	    RECT 179.4000 1371.4501 180.6000 1371.6000 ;
	    RECT 174.6000 1370.5500 180.6000 1371.4501 ;
	    RECT 174.6000 1370.4000 175.8000 1370.5500 ;
	    RECT 179.4000 1370.4000 180.6000 1370.5500 ;
	    RECT 160.2000 1368.6000 173.7000 1369.5000 ;
	    RECT 131.4000 1367.4000 132.6000 1368.6000 ;
	    RECT 136.5000 1367.7001 137.7000 1368.0000 ;
	    RECT 133.5000 1366.8000 171.9000 1367.7001 ;
	    RECT 170.7000 1366.5000 171.9000 1366.8000 ;
	    RECT 172.8000 1365.9000 173.7000 1368.6000 ;
	    RECT 174.6000 1368.0000 175.8000 1369.5000 ;
	    RECT 174.6000 1366.8000 176.1000 1368.0000 ;
	    RECT 128.7000 1365.0000 135.3000 1365.9000 ;
	    RECT 128.7000 1364.7001 129.9000 1365.0000 ;
	    RECT 136.2000 1364.4000 137.4000 1365.6000 ;
	    RECT 138.3000 1365.0000 163.8000 1365.9000 ;
	    RECT 172.8000 1365.0000 174.0000 1365.9000 ;
	    RECT 162.6000 1364.1000 163.8000 1365.0000 ;
	    RECT 126.6000 1362.3000 139.8000 1363.5000 ;
	    RECT 140.7000 1362.9000 143.7000 1364.1000 ;
	    RECT 149.4000 1362.9000 154.2000 1364.1000 ;
	    RECT 126.6000 1353.3000 127.8000 1362.3000 ;
	    RECT 130.2000 1360.2001 134.7000 1361.4000 ;
	    RECT 133.5000 1359.3000 134.7000 1360.2001 ;
	    RECT 142.5000 1359.3000 143.7000 1362.9000 ;
	    RECT 145.8000 1361.4000 147.0000 1362.6000 ;
	    RECT 153.6000 1361.7001 154.8000 1362.0000 ;
	    RECT 148.2000 1360.8000 154.8000 1361.7001 ;
	    RECT 148.2000 1360.5000 149.4000 1360.8000 ;
	    RECT 145.8000 1360.2001 147.0000 1360.5000 ;
	    RECT 157.8000 1359.6000 159.0000 1363.8000 ;
	    RECT 166.5000 1362.9000 172.2000 1364.1000 ;
	    RECT 166.5000 1361.1000 167.7000 1362.9000 ;
	    RECT 173.1000 1362.0000 174.0000 1365.0000 ;
	    RECT 148.2000 1359.3000 149.4000 1359.6000 ;
	    RECT 131.4000 1353.3000 132.6000 1359.3000 ;
	    RECT 133.5000 1358.1000 137.4000 1359.3000 ;
	    RECT 142.5000 1358.4000 149.4000 1359.3000 ;
	    RECT 150.6000 1358.4000 151.8000 1359.6000 ;
	    RECT 152.7000 1358.4000 153.0000 1359.6000 ;
	    RECT 157.5000 1358.4000 159.0000 1359.6000 ;
	    RECT 165.0000 1360.2001 167.7000 1361.1000 ;
	    RECT 172.2000 1361.1000 174.0000 1362.0000 ;
	    RECT 165.0000 1359.3000 166.2000 1360.2001 ;
	    RECT 136.2000 1353.3000 137.4000 1358.1000 ;
	    RECT 162.6000 1358.1000 166.2000 1359.3000 ;
	    RECT 138.6000 1353.3000 139.8000 1357.5000 ;
	    RECT 141.0000 1353.3000 142.2000 1357.5000 ;
	    RECT 143.4000 1353.3000 144.6000 1357.5000 ;
	    RECT 145.8000 1353.3000 147.0000 1356.3000 ;
	    RECT 148.2000 1353.3000 149.4000 1357.5000 ;
	    RECT 150.6000 1353.3000 151.8000 1356.3000 ;
	    RECT 153.0000 1353.3000 154.2000 1357.5000 ;
	    RECT 155.4000 1353.3000 156.6000 1357.5000 ;
	    RECT 157.8000 1353.3000 159.0000 1357.5000 ;
	    RECT 160.2000 1353.3000 161.4000 1357.5000 ;
	    RECT 162.6000 1353.3000 163.8000 1358.1000 ;
	    RECT 167.4000 1353.3000 168.6000 1359.3000 ;
	    RECT 172.2000 1353.3000 173.4000 1361.1000 ;
	    RECT 174.9000 1360.2001 176.1000 1366.8000 ;
	    RECT 193.8000 1363.5000 195.0000 1379.7001 ;
	    RECT 220.2000 1373.7001 221.4000 1379.7001 ;
	    RECT 222.6000 1366.5000 223.8000 1379.7001 ;
	    RECT 225.0000 1373.7001 226.2000 1379.7001 ;
	    RECT 349.8000 1373.7001 351.0000 1379.7001 ;
	    RECT 352.2000 1374.6000 353.4000 1379.7001 ;
	    RECT 351.9000 1373.7001 353.4000 1374.6000 ;
	    RECT 354.6000 1373.7001 355.8000 1380.6000 ;
	    RECT 351.9000 1372.8000 352.8000 1373.7001 ;
	    RECT 357.0000 1372.8000 358.2000 1379.7001 ;
	    RECT 359.4000 1373.7001 360.6000 1379.7001 ;
	    RECT 361.8000 1375.5000 363.0000 1379.7001 ;
	    RECT 364.2000 1375.5000 365.4000 1379.7001 ;
	    RECT 349.8000 1371.9000 352.8000 1372.8000 ;
	    RECT 225.0000 1369.5000 226.2000 1369.8000 ;
	    RECT 225.0000 1368.4501 226.2000 1368.6000 ;
	    RECT 244.2000 1368.4501 245.4000 1368.6000 ;
	    RECT 225.0000 1367.5500 245.4000 1368.4501 ;
	    RECT 225.0000 1367.4000 226.2000 1367.5500 ;
	    RECT 244.2000 1367.4000 245.4000 1367.5500 ;
	    RECT 222.6000 1365.4501 223.8000 1365.6000 ;
	    RECT 225.0000 1365.4501 226.2000 1365.6000 ;
	    RECT 222.6000 1364.5500 226.2000 1365.4501 ;
	    RECT 222.6000 1364.4000 223.8000 1364.5500 ;
	    RECT 225.0000 1364.4000 226.2000 1364.5500 ;
	    RECT 349.8000 1363.5000 351.0000 1371.9000 ;
	    RECT 353.7000 1371.6000 360.0000 1372.8000 ;
	    RECT 366.6000 1372.5000 367.8000 1379.7001 ;
	    RECT 369.0000 1373.7001 370.2000 1379.7001 ;
	    RECT 371.4000 1372.5000 372.6000 1379.7001 ;
	    RECT 373.8000 1373.7001 375.0000 1379.7001 ;
	    RECT 353.7000 1371.0000 354.6000 1371.6000 ;
	    RECT 352.2000 1369.8000 354.6000 1371.0000 ;
	    RECT 359.1000 1370.7001 367.8000 1371.6000 ;
	    RECT 356.1000 1369.8000 358.2000 1370.7001 ;
	    RECT 356.1000 1369.5000 365.4000 1369.8000 ;
	    RECT 357.3000 1368.9000 365.4000 1369.5000 ;
	    RECT 364.2000 1368.6000 365.4000 1368.9000 ;
	    RECT 366.9000 1369.5000 367.8000 1370.7001 ;
	    RECT 368.7000 1370.4000 372.6000 1371.6000 ;
	    RECT 376.2000 1370.4000 377.4000 1379.7001 ;
	    RECT 378.6000 1375.5000 379.8000 1379.7001 ;
	    RECT 381.0000 1375.5000 382.2000 1379.7001 ;
	    RECT 383.4000 1375.5000 384.6000 1379.7001 ;
	    RECT 385.8000 1373.7001 387.0000 1379.7001 ;
	    RECT 381.0000 1371.6000 387.3000 1372.8000 ;
	    RECT 388.2000 1371.6000 389.4000 1379.7001 ;
	    RECT 390.6000 1373.7001 391.8000 1379.7001 ;
	    RECT 393.0000 1372.8000 394.2000 1379.7001 ;
	    RECT 395.4000 1373.7001 396.6000 1379.7001 ;
	    RECT 393.0000 1371.9000 396.9000 1372.8000 ;
	    RECT 397.8000 1372.5000 399.0000 1379.7001 ;
	    RECT 400.2000 1373.7001 401.4000 1379.7001 ;
	    RECT 388.2000 1370.4000 392.1000 1371.6000 ;
	    RECT 378.6000 1369.5000 379.8000 1369.8000 ;
	    RECT 366.9000 1368.6000 379.8000 1369.5000 ;
	    RECT 383.4000 1369.5000 384.6000 1369.8000 ;
	    RECT 396.0000 1369.5000 396.9000 1371.9000 ;
	    RECT 397.8000 1370.4000 399.0000 1371.6000 ;
	    RECT 383.4000 1368.6000 396.9000 1369.5000 ;
	    RECT 354.6000 1367.4000 355.8000 1368.6000 ;
	    RECT 359.7000 1367.7001 360.9000 1368.0000 ;
	    RECT 356.7000 1366.8000 395.1000 1367.7001 ;
	    RECT 393.9000 1366.5000 395.1000 1366.8000 ;
	    RECT 396.0000 1365.9000 396.9000 1368.6000 ;
	    RECT 397.8000 1368.0000 399.0000 1369.5000 ;
	    RECT 397.8000 1366.8000 399.3000 1368.0000 ;
	    RECT 351.9000 1365.0000 358.5000 1365.9000 ;
	    RECT 351.9000 1364.7001 353.1000 1365.0000 ;
	    RECT 359.4000 1364.4000 360.6000 1365.6000 ;
	    RECT 361.5000 1365.0000 387.0000 1365.9000 ;
	    RECT 396.0000 1365.0000 397.2000 1365.9000 ;
	    RECT 385.8000 1364.1000 387.0000 1365.0000 ;
	    RECT 193.8000 1362.4501 195.0000 1362.6000 ;
	    RECT 196.2000 1362.4501 197.4000 1362.6000 ;
	    RECT 193.8000 1361.5500 197.4000 1362.4501 ;
	    RECT 193.8000 1361.4000 195.0000 1361.5500 ;
	    RECT 196.2000 1361.4000 197.4000 1361.5500 ;
	    RECT 220.2000 1361.4000 221.4000 1362.6000 ;
	    RECT 174.6000 1359.0000 176.1000 1360.2001 ;
	    RECT 189.0000 1359.4501 190.2000 1359.6000 ;
	    RECT 191.4000 1359.4501 192.6000 1359.6000 ;
	    RECT 174.6000 1353.3000 175.8000 1359.0000 ;
	    RECT 189.0000 1358.5500 192.6000 1359.4501 ;
	    RECT 189.0000 1358.4000 190.2000 1358.5500 ;
	    RECT 191.4000 1358.4000 192.6000 1358.5500 ;
	    RECT 191.4000 1357.2001 192.6000 1357.5000 ;
	    RECT 177.0000 1353.3000 178.2000 1356.3000 ;
	    RECT 191.4000 1353.3000 192.6000 1356.3000 ;
	    RECT 193.8000 1353.3000 195.0000 1360.5000 ;
	    RECT 220.2000 1360.2001 221.4000 1360.5000 ;
	    RECT 222.6000 1359.3000 223.8000 1363.5000 ;
	    RECT 349.8000 1362.3000 363.0000 1363.5000 ;
	    RECT 363.9000 1362.9000 366.9000 1364.1000 ;
	    RECT 372.6000 1362.9000 377.4000 1364.1000 ;
	    RECT 220.2000 1353.3000 221.4000 1359.3000 ;
	    RECT 222.6000 1358.4000 225.3000 1359.3000 ;
	    RECT 224.1000 1353.3000 225.3000 1358.4000 ;
	    RECT 349.8000 1353.3000 351.0000 1362.3000 ;
	    RECT 353.4000 1360.2001 357.9000 1361.4000 ;
	    RECT 356.7000 1359.3000 357.9000 1360.2001 ;
	    RECT 365.7000 1359.3000 366.9000 1362.9000 ;
	    RECT 369.0000 1361.4000 370.2000 1362.6000 ;
	    RECT 376.8000 1361.7001 378.0000 1362.0000 ;
	    RECT 371.4000 1360.8000 378.0000 1361.7001 ;
	    RECT 371.4000 1360.5000 372.6000 1360.8000 ;
	    RECT 369.0000 1360.2001 370.2000 1360.5000 ;
	    RECT 381.0000 1359.6000 382.2000 1363.8000 ;
	    RECT 389.7000 1362.9000 395.4000 1364.1000 ;
	    RECT 389.7000 1361.1000 390.9000 1362.9000 ;
	    RECT 396.3000 1362.0000 397.2000 1365.0000 ;
	    RECT 371.4000 1359.3000 372.6000 1359.6000 ;
	    RECT 354.6000 1353.3000 355.8000 1359.3000 ;
	    RECT 356.7000 1358.1000 360.6000 1359.3000 ;
	    RECT 365.7000 1358.4000 372.6000 1359.3000 ;
	    RECT 373.8000 1358.4000 375.0000 1359.6000 ;
	    RECT 375.9000 1358.4000 376.2000 1359.6000 ;
	    RECT 380.7000 1358.4000 382.2000 1359.6000 ;
	    RECT 388.2000 1360.2001 390.9000 1361.1000 ;
	    RECT 395.4000 1361.1000 397.2000 1362.0000 ;
	    RECT 388.2000 1359.3000 389.4000 1360.2001 ;
	    RECT 359.4000 1353.3000 360.6000 1358.1000 ;
	    RECT 385.8000 1358.1000 389.4000 1359.3000 ;
	    RECT 361.8000 1353.3000 363.0000 1357.5000 ;
	    RECT 364.2000 1353.3000 365.4000 1357.5000 ;
	    RECT 366.6000 1353.3000 367.8000 1357.5000 ;
	    RECT 369.0000 1353.3000 370.2000 1356.3000 ;
	    RECT 371.4000 1353.3000 372.6000 1357.5000 ;
	    RECT 373.8000 1353.3000 375.0000 1356.3000 ;
	    RECT 376.2000 1353.3000 377.4000 1357.5000 ;
	    RECT 378.6000 1353.3000 379.8000 1357.5000 ;
	    RECT 381.0000 1353.3000 382.2000 1357.5000 ;
	    RECT 383.4000 1353.3000 384.6000 1357.5000 ;
	    RECT 385.8000 1353.3000 387.0000 1358.1000 ;
	    RECT 390.6000 1353.3000 391.8000 1359.3000 ;
	    RECT 395.4000 1353.3000 396.6000 1361.1000 ;
	    RECT 398.1000 1360.2001 399.3000 1366.8000 ;
	    RECT 414.6000 1363.5000 415.8000 1379.7001 ;
	    RECT 417.0000 1373.7001 418.2000 1379.7001 ;
	    RECT 431.4000 1363.5000 432.6000 1379.7001 ;
	    RECT 433.8000 1373.7001 435.0000 1379.7001 ;
	    RECT 460.2000 1373.7001 461.4000 1379.7001 ;
	    RECT 460.2000 1369.5000 461.4000 1369.8000 ;
	    RECT 460.2000 1367.4000 461.4000 1368.6000 ;
	    RECT 462.6000 1366.5000 463.8000 1379.7001 ;
	    RECT 465.0000 1373.7001 466.2000 1379.7001 ;
	    RECT 489.9000 1373.7001 491.1000 1379.7001 ;
	    RECT 490.2000 1370.4000 491.4000 1371.6000 ;
	    RECT 490.2000 1369.5000 491.1000 1370.4000 ;
	    RECT 492.3000 1368.6000 493.5000 1379.7001 ;
	    RECT 489.0000 1367.4000 490.2000 1368.6000 ;
	    RECT 492.0000 1367.7001 493.5000 1368.6000 ;
	    RECT 496.2000 1367.7001 497.4000 1379.7001 ;
	    RECT 508.2000 1373.7001 509.4000 1379.7001 ;
	    RECT 462.6000 1365.4501 463.8000 1365.6000 ;
	    RECT 489.1500 1365.4501 490.0500 1367.4000 ;
	    RECT 462.6000 1364.5500 490.0500 1365.4501 ;
	    RECT 462.6000 1364.4000 463.8000 1364.5500 ;
	    RECT 400.2000 1362.4501 401.4000 1362.6000 ;
	    RECT 414.6000 1362.4501 415.8000 1362.6000 ;
	    RECT 429.0000 1362.4501 430.2000 1362.6000 ;
	    RECT 400.2000 1361.5500 430.2000 1362.4501 ;
	    RECT 400.2000 1361.4000 401.4000 1361.5500 ;
	    RECT 414.6000 1361.4000 415.8000 1361.5500 ;
	    RECT 429.0000 1361.4000 430.2000 1361.5500 ;
	    RECT 431.4000 1362.4501 432.6000 1362.6000 ;
	    RECT 457.8000 1362.4501 459.0000 1362.6000 ;
	    RECT 431.4000 1361.5500 459.0000 1362.4501 ;
	    RECT 431.4000 1361.4000 432.6000 1361.5500 ;
	    RECT 457.8000 1361.4000 459.0000 1361.5500 ;
	    RECT 397.8000 1359.0000 399.3000 1360.2001 ;
	    RECT 397.8000 1353.3000 399.0000 1359.0000 ;
	    RECT 400.2000 1353.3000 401.4000 1356.3000 ;
	    RECT 414.6000 1353.3000 415.8000 1360.5000 ;
	    RECT 417.0000 1358.4000 418.2000 1359.6000 ;
	    RECT 417.0000 1357.2001 418.2000 1357.5000 ;
	    RECT 417.0000 1353.3000 418.2000 1356.3000 ;
	    RECT 431.4000 1353.3000 432.6000 1360.5000 ;
	    RECT 433.8000 1359.4501 435.0000 1359.6000 ;
	    RECT 457.8000 1359.4501 459.0000 1359.6000 ;
	    RECT 433.8000 1358.5500 459.0000 1359.4501 ;
	    RECT 462.6000 1359.3000 463.8000 1363.5000 ;
	    RECT 492.0000 1362.6000 492.9000 1367.7001 ;
	    RECT 493.8000 1364.4000 495.0000 1365.6000 ;
	    RECT 510.6000 1363.5000 511.8000 1379.7001 ;
	    RECT 637.8000 1373.7001 639.0000 1379.7001 ;
	    RECT 640.2000 1372.5000 641.4000 1379.7001 ;
	    RECT 642.6000 1373.7001 643.8000 1379.7001 ;
	    RECT 645.0000 1372.8000 646.2000 1379.7001 ;
	    RECT 647.4000 1373.7001 648.6000 1379.7001 ;
	    RECT 642.3000 1371.9000 646.2000 1372.8000 ;
	    RECT 633.0000 1371.4501 634.2000 1371.6000 ;
	    RECT 640.2000 1371.4501 641.4000 1371.6000 ;
	    RECT 633.0000 1370.5500 641.4000 1371.4501 ;
	    RECT 633.0000 1370.4000 634.2000 1370.5500 ;
	    RECT 640.2000 1370.4000 641.4000 1370.5500 ;
	    RECT 642.3000 1369.5000 643.2000 1371.9000 ;
	    RECT 649.8000 1371.6000 651.0000 1379.7001 ;
	    RECT 652.2000 1373.7001 653.4000 1379.7001 ;
	    RECT 654.6000 1375.5000 655.8000 1379.7001 ;
	    RECT 657.0000 1375.5000 658.2000 1379.7001 ;
	    RECT 659.4000 1375.5000 660.6000 1379.7001 ;
	    RECT 651.9000 1371.6000 658.2000 1372.8000 ;
	    RECT 647.1000 1370.4000 651.0000 1371.6000 ;
	    RECT 661.8000 1370.4000 663.0000 1379.7001 ;
	    RECT 664.2000 1373.7001 665.4000 1379.7001 ;
	    RECT 666.6000 1372.5000 667.8000 1379.7001 ;
	    RECT 669.0000 1373.7001 670.2000 1379.7001 ;
	    RECT 671.4000 1372.5000 672.6000 1379.7001 ;
	    RECT 673.8000 1375.5000 675.0000 1379.7001 ;
	    RECT 676.2000 1375.5000 677.4000 1379.7001 ;
	    RECT 678.6000 1373.7001 679.8000 1379.7001 ;
	    RECT 681.0000 1372.8000 682.2000 1379.7001 ;
	    RECT 683.4000 1373.7001 684.6000 1380.6000 ;
	    RECT 685.8000 1374.6000 687.0000 1379.7001 ;
	    RECT 685.8000 1373.7001 687.3000 1374.6000 ;
	    RECT 688.2000 1373.7001 689.4000 1379.7001 ;
	    RECT 714.6000 1373.7001 715.8000 1379.7001 ;
	    RECT 686.4000 1372.8000 687.3000 1373.7001 ;
	    RECT 679.2000 1371.6000 685.5000 1372.8000 ;
	    RECT 686.4000 1371.9000 689.4000 1372.8000 ;
	    RECT 666.6000 1370.4000 670.5000 1371.6000 ;
	    RECT 671.4000 1370.7001 680.1000 1371.6000 ;
	    RECT 684.6000 1371.0000 685.5000 1371.6000 ;
	    RECT 654.6000 1369.5000 655.8000 1369.8000 ;
	    RECT 640.2000 1368.0000 641.4000 1369.5000 ;
	    RECT 639.9000 1366.8000 641.4000 1368.0000 ;
	    RECT 642.3000 1368.6000 655.8000 1369.5000 ;
	    RECT 659.4000 1369.5000 660.6000 1369.8000 ;
	    RECT 671.4000 1369.5000 672.3000 1370.7001 ;
	    RECT 681.0000 1369.8000 683.1000 1370.7001 ;
	    RECT 684.6000 1369.8000 687.0000 1371.0000 ;
	    RECT 659.4000 1368.6000 672.3000 1369.5000 ;
	    RECT 673.8000 1369.5000 683.1000 1369.8000 ;
	    RECT 673.8000 1368.9000 681.9000 1369.5000 ;
	    RECT 673.8000 1368.6000 675.0000 1368.9000 ;
	    RECT 493.8000 1363.2001 495.0000 1363.5000 ;
	    RECT 465.0000 1362.4501 466.2000 1362.6000 ;
	    RECT 479.4000 1362.4501 480.6000 1362.6000 ;
	    RECT 465.0000 1361.5500 480.6000 1362.4501 ;
	    RECT 465.0000 1361.4000 466.2000 1361.5500 ;
	    RECT 479.4000 1361.4000 480.6000 1361.5500 ;
	    RECT 489.0000 1361.4000 490.2000 1362.6000 ;
	    RECT 491.1000 1361.4000 492.9000 1362.6000 ;
	    RECT 495.0000 1360.8000 495.3000 1362.3000 ;
	    RECT 496.2000 1361.4000 497.4000 1362.6000 ;
	    RECT 510.6000 1362.4501 511.8000 1362.6000 ;
	    RECT 575.4000 1362.4501 576.6000 1362.6000 ;
	    RECT 637.8000 1362.4501 639.0000 1362.6000 ;
	    RECT 510.6000 1361.5500 639.0000 1362.4501 ;
	    RECT 510.6000 1361.4000 511.8000 1361.5500 ;
	    RECT 575.4000 1361.4000 576.6000 1361.5500 ;
	    RECT 637.8000 1361.4000 639.0000 1361.5500 ;
	    RECT 465.0000 1360.2001 466.2000 1360.5000 ;
	    RECT 489.3000 1359.3000 490.2000 1360.5000 ;
	    RECT 491.7000 1359.3000 497.1000 1359.9000 ;
	    RECT 433.8000 1358.4000 435.0000 1358.5500 ;
	    RECT 457.8000 1358.4000 459.0000 1358.5500 ;
	    RECT 461.1000 1358.4000 463.8000 1359.3000 ;
	    RECT 433.8000 1357.2001 435.0000 1357.5000 ;
	    RECT 433.8000 1353.3000 435.0000 1356.3000 ;
	    RECT 461.1000 1353.3000 462.3000 1358.4000 ;
	    RECT 465.0000 1353.3000 466.2000 1359.3000 ;
	    RECT 489.0000 1353.3000 490.2000 1359.3000 ;
	    RECT 491.4000 1359.0000 497.4000 1359.3000 ;
	    RECT 491.4000 1353.3000 492.6000 1359.0000 ;
	    RECT 493.8000 1353.3000 495.0000 1358.1000 ;
	    RECT 496.2000 1353.3000 497.4000 1359.0000 ;
	    RECT 508.2000 1358.4000 509.4000 1359.6000 ;
	    RECT 508.2000 1357.2001 509.4000 1357.5000 ;
	    RECT 508.2000 1353.3000 509.4000 1356.3000 ;
	    RECT 510.6000 1353.3000 511.8000 1360.5000 ;
	    RECT 639.9000 1360.2001 641.1000 1366.8000 ;
	    RECT 642.3000 1365.9000 643.2000 1368.6000 ;
	    RECT 678.3000 1367.7001 679.5000 1368.0000 ;
	    RECT 644.1000 1366.8000 682.5000 1367.7001 ;
	    RECT 683.4000 1367.4000 684.6000 1368.6000 ;
	    RECT 644.1000 1366.5000 645.3000 1366.8000 ;
	    RECT 642.0000 1365.0000 643.2000 1365.9000 ;
	    RECT 652.2000 1365.0000 677.7000 1365.9000 ;
	    RECT 642.0000 1362.0000 642.9000 1365.0000 ;
	    RECT 652.2000 1364.1000 653.4000 1365.0000 ;
	    RECT 678.6000 1364.4000 679.8000 1365.6000 ;
	    RECT 680.7000 1365.0000 687.3000 1365.9000 ;
	    RECT 686.1000 1364.7001 687.3000 1365.0000 ;
	    RECT 643.8000 1362.9000 649.5000 1364.1000 ;
	    RECT 642.0000 1361.1000 643.8000 1362.0000 ;
	    RECT 639.9000 1359.0000 641.4000 1360.2001 ;
	    RECT 637.8000 1353.3000 639.0000 1356.3000 ;
	    RECT 640.2000 1353.3000 641.4000 1359.0000 ;
	    RECT 642.6000 1353.3000 643.8000 1361.1000 ;
	    RECT 648.3000 1361.1000 649.5000 1362.9000 ;
	    RECT 648.3000 1360.2001 651.0000 1361.1000 ;
	    RECT 649.8000 1359.3000 651.0000 1360.2001 ;
	    RECT 657.0000 1359.6000 658.2000 1363.8000 ;
	    RECT 661.8000 1362.9000 666.6000 1364.1000 ;
	    RECT 672.3000 1362.9000 675.3000 1364.1000 ;
	    RECT 688.2000 1363.5000 689.4000 1371.9000 ;
	    RECT 714.6000 1369.5000 715.8000 1369.8000 ;
	    RECT 697.8000 1368.4501 699.0000 1368.6000 ;
	    RECT 714.6000 1368.4501 715.8000 1368.6000 ;
	    RECT 697.8000 1367.5500 715.8000 1368.4501 ;
	    RECT 697.8000 1367.4000 699.0000 1367.5500 ;
	    RECT 714.6000 1367.4000 715.8000 1367.5500 ;
	    RECT 717.0000 1366.5000 718.2000 1379.7001 ;
	    RECT 719.4000 1373.7001 720.6000 1379.7001 ;
	    RECT 741.0000 1377.4501 742.2000 1377.6000 ;
	    RECT 743.5500 1377.4501 744.4500 1380.6000 ;
	    RECT 741.0000 1376.5500 744.4500 1377.4501 ;
	    RECT 741.0000 1376.4000 742.2000 1376.5500 ;
	    RECT 846.6000 1373.7001 847.8000 1379.7001 ;
	    RECT 849.0000 1372.5000 850.2000 1379.7001 ;
	    RECT 851.4000 1373.7001 852.6000 1379.7001 ;
	    RECT 853.8000 1372.8000 855.0000 1379.7001 ;
	    RECT 856.2000 1373.7001 857.4000 1379.7001 ;
	    RECT 851.1000 1371.9000 855.0000 1372.8000 ;
	    RECT 825.0000 1371.4501 826.2000 1371.6000 ;
	    RECT 849.0000 1371.4501 850.2000 1371.6000 ;
	    RECT 825.0000 1370.5500 850.2000 1371.4501 ;
	    RECT 825.0000 1370.4000 826.2000 1370.5500 ;
	    RECT 849.0000 1370.4000 850.2000 1370.5500 ;
	    RECT 851.1000 1369.5000 852.0000 1371.9000 ;
	    RECT 858.6000 1371.6000 859.8000 1379.7001 ;
	    RECT 861.0000 1373.7001 862.2000 1379.7001 ;
	    RECT 863.4000 1375.5000 864.6000 1379.7001 ;
	    RECT 865.8000 1375.5000 867.0000 1379.7001 ;
	    RECT 868.2000 1375.5000 869.4000 1379.7001 ;
	    RECT 860.7000 1371.6000 867.0000 1372.8000 ;
	    RECT 855.9000 1370.4000 859.8000 1371.6000 ;
	    RECT 870.6000 1370.4000 871.8000 1379.7001 ;
	    RECT 873.0000 1373.7001 874.2000 1379.7001 ;
	    RECT 875.4000 1372.5000 876.6000 1379.7001 ;
	    RECT 877.8000 1373.7001 879.0000 1379.7001 ;
	    RECT 880.2000 1372.5000 881.4000 1379.7001 ;
	    RECT 882.6000 1375.5000 883.8000 1379.7001 ;
	    RECT 885.0000 1375.5000 886.2000 1379.7001 ;
	    RECT 887.4000 1373.7001 888.6000 1379.7001 ;
	    RECT 889.8000 1372.8000 891.0000 1379.7001 ;
	    RECT 892.2000 1373.7001 893.4000 1380.6000 ;
	    RECT 894.6000 1374.6000 895.8000 1379.7001 ;
	    RECT 894.6000 1373.7001 896.1000 1374.6000 ;
	    RECT 897.0000 1373.7001 898.2000 1379.7001 ;
	    RECT 921.0000 1373.7001 922.2000 1379.7001 ;
	    RECT 895.2000 1372.8000 896.1000 1373.7001 ;
	    RECT 888.0000 1371.6000 894.3000 1372.8000 ;
	    RECT 895.2000 1371.9000 898.2000 1372.8000 ;
	    RECT 875.4000 1370.4000 879.3000 1371.6000 ;
	    RECT 880.2000 1370.7001 888.9000 1371.6000 ;
	    RECT 893.4000 1371.0000 894.3000 1371.6000 ;
	    RECT 863.4000 1369.5000 864.6000 1369.8000 ;
	    RECT 849.0000 1368.0000 850.2000 1369.5000 ;
	    RECT 848.7000 1366.8000 850.2000 1368.0000 ;
	    RECT 851.1000 1368.6000 864.6000 1369.5000 ;
	    RECT 868.2000 1369.5000 869.4000 1369.8000 ;
	    RECT 880.2000 1369.5000 881.1000 1370.7001 ;
	    RECT 889.8000 1369.8000 891.9000 1370.7001 ;
	    RECT 893.4000 1369.8000 895.8000 1371.0000 ;
	    RECT 868.2000 1368.6000 881.1000 1369.5000 ;
	    RECT 882.6000 1369.5000 891.9000 1369.8000 ;
	    RECT 882.6000 1368.9000 890.7000 1369.5000 ;
	    RECT 882.6000 1368.6000 883.8000 1368.9000 ;
	    RECT 717.0000 1365.4501 718.2000 1365.6000 ;
	    RECT 724.2000 1365.4501 725.4000 1365.6000 ;
	    RECT 717.0000 1364.5500 725.4000 1365.4501 ;
	    RECT 717.0000 1364.4000 718.2000 1364.5500 ;
	    RECT 724.2000 1364.4000 725.4000 1364.5500 ;
	    RECT 661.2000 1361.7001 662.4000 1362.0000 ;
	    RECT 661.2000 1360.8000 667.8000 1361.7001 ;
	    RECT 669.0000 1361.4000 670.2000 1362.6000 ;
	    RECT 666.6000 1360.5000 667.8000 1360.8000 ;
	    RECT 669.0000 1360.2001 670.2000 1360.5000 ;
	    RECT 647.4000 1353.3000 648.6000 1359.3000 ;
	    RECT 649.8000 1358.1000 653.4000 1359.3000 ;
	    RECT 657.0000 1358.4000 658.5000 1359.6000 ;
	    RECT 663.0000 1358.4000 663.3000 1359.6000 ;
	    RECT 664.2000 1358.4000 665.4000 1359.6000 ;
	    RECT 666.6000 1359.3000 667.8000 1359.6000 ;
	    RECT 672.3000 1359.3000 673.5000 1362.9000 ;
	    RECT 676.2000 1362.3000 689.4000 1363.5000 ;
	    RECT 681.3000 1360.2001 685.8000 1361.4000 ;
	    RECT 681.3000 1359.3000 682.5000 1360.2001 ;
	    RECT 666.6000 1358.4000 673.5000 1359.3000 ;
	    RECT 652.2000 1353.3000 653.4000 1358.1000 ;
	    RECT 678.6000 1358.1000 682.5000 1359.3000 ;
	    RECT 654.6000 1353.3000 655.8000 1357.5000 ;
	    RECT 657.0000 1353.3000 658.2000 1357.5000 ;
	    RECT 659.4000 1353.3000 660.6000 1357.5000 ;
	    RECT 661.8000 1353.3000 663.0000 1357.5000 ;
	    RECT 664.2000 1353.3000 665.4000 1356.3000 ;
	    RECT 666.6000 1353.3000 667.8000 1357.5000 ;
	    RECT 669.0000 1353.3000 670.2000 1356.3000 ;
	    RECT 671.4000 1353.3000 672.6000 1357.5000 ;
	    RECT 673.8000 1353.3000 675.0000 1357.5000 ;
	    RECT 676.2000 1353.3000 677.4000 1357.5000 ;
	    RECT 678.6000 1353.3000 679.8000 1358.1000 ;
	    RECT 683.4000 1353.3000 684.6000 1359.3000 ;
	    RECT 688.2000 1353.3000 689.4000 1362.3000 ;
	    RECT 717.0000 1359.3000 718.2000 1363.5000 ;
	    RECT 719.4000 1361.4000 720.6000 1362.6000 ;
	    RECT 719.4000 1360.2001 720.6000 1360.5000 ;
	    RECT 848.7000 1360.2001 849.9000 1366.8000 ;
	    RECT 851.1000 1365.9000 852.0000 1368.6000 ;
	    RECT 887.1000 1367.7001 888.3000 1368.0000 ;
	    RECT 852.9000 1366.8000 891.3000 1367.7001 ;
	    RECT 892.2000 1367.4000 893.4000 1368.6000 ;
	    RECT 852.9000 1366.5000 854.1000 1366.8000 ;
	    RECT 850.8000 1365.0000 852.0000 1365.9000 ;
	    RECT 861.0000 1365.0000 886.5000 1365.9000 ;
	    RECT 850.8000 1362.0000 851.7000 1365.0000 ;
	    RECT 861.0000 1364.1000 862.2000 1365.0000 ;
	    RECT 887.4000 1364.4000 888.6000 1365.6000 ;
	    RECT 889.5000 1365.0000 896.1000 1365.9000 ;
	    RECT 894.9000 1364.7001 896.1000 1365.0000 ;
	    RECT 852.6000 1362.9000 858.3000 1364.1000 ;
	    RECT 850.8000 1361.1000 852.6000 1362.0000 ;
	    RECT 715.5000 1358.4000 718.2000 1359.3000 ;
	    RECT 715.5000 1353.3000 716.7000 1358.4000 ;
	    RECT 719.4000 1353.3000 720.6000 1359.3000 ;
	    RECT 848.7000 1359.0000 850.2000 1360.2001 ;
	    RECT 846.6000 1353.3000 847.8000 1356.3000 ;
	    RECT 849.0000 1353.3000 850.2000 1359.0000 ;
	    RECT 851.4000 1353.3000 852.6000 1361.1000 ;
	    RECT 857.1000 1361.1000 858.3000 1362.9000 ;
	    RECT 857.1000 1360.2001 859.8000 1361.1000 ;
	    RECT 858.6000 1359.3000 859.8000 1360.2001 ;
	    RECT 865.8000 1359.6000 867.0000 1363.8000 ;
	    RECT 870.6000 1362.9000 875.4000 1364.1000 ;
	    RECT 881.1000 1362.9000 884.1000 1364.1000 ;
	    RECT 897.0000 1363.5000 898.2000 1371.9000 ;
	    RECT 923.4000 1366.5000 924.6000 1379.7001 ;
	    RECT 925.8000 1373.7001 927.0000 1379.7001 ;
	    RECT 940.2000 1373.7001 941.4000 1379.7001 ;
	    RECT 925.8000 1369.5000 927.0000 1369.8000 ;
	    RECT 925.8000 1367.4000 927.0000 1368.6000 ;
	    RECT 921.0000 1365.4501 922.2000 1365.6000 ;
	    RECT 923.4000 1365.4501 924.6000 1365.6000 ;
	    RECT 921.0000 1364.5500 924.6000 1365.4501 ;
	    RECT 921.0000 1364.4000 922.2000 1364.5500 ;
	    RECT 923.4000 1364.4000 924.6000 1364.5500 ;
	    RECT 942.6000 1363.5000 943.8000 1379.7001 ;
	    RECT 957.0000 1373.7001 958.2000 1379.7001 ;
	    RECT 959.4000 1363.5000 960.6000 1379.7001 ;
	    RECT 969.0000 1379.4000 970.2000 1380.6000 ;
	    RECT 978.6000 1373.7001 979.8000 1379.7001 ;
	    RECT 978.6000 1369.5000 979.8000 1369.8000 ;
	    RECT 973.8000 1368.4501 975.0000 1368.6000 ;
	    RECT 978.6000 1368.4501 979.8000 1368.6000 ;
	    RECT 973.8000 1367.5500 979.8000 1368.4501 ;
	    RECT 973.8000 1367.4000 975.0000 1367.5500 ;
	    RECT 978.6000 1367.4000 979.8000 1367.5500 ;
	    RECT 981.0000 1366.5000 982.2000 1379.7001 ;
	    RECT 983.4000 1373.7001 984.6000 1379.7001 ;
	    RECT 1031.4000 1379.4000 1032.6000 1380.6000 ;
	    RECT 1084.2001 1379.4000 1085.4000 1380.6000 ;
	    RECT 1115.4000 1373.7001 1116.6000 1379.7001 ;
	    RECT 1117.8000 1374.6000 1119.0000 1379.7001 ;
	    RECT 1117.5000 1373.7001 1119.0000 1374.6000 ;
	    RECT 1120.2001 1373.7001 1121.4000 1380.6000 ;
	    RECT 1117.5000 1372.8000 1118.4000 1373.7001 ;
	    RECT 1122.6000 1372.8000 1123.8000 1379.7001 ;
	    RECT 1125.0000 1373.7001 1126.2001 1379.7001 ;
	    RECT 1127.4000 1375.5000 1128.6000 1379.7001 ;
	    RECT 1129.8000 1375.5000 1131.0000 1379.7001 ;
	    RECT 1115.4000 1371.9000 1118.4000 1372.8000 ;
	    RECT 981.0000 1365.4501 982.2000 1365.6000 ;
	    RECT 1012.2000 1365.4501 1013.4000 1365.6000 ;
	    RECT 981.0000 1364.5500 1013.4000 1365.4501 ;
	    RECT 981.0000 1364.4000 982.2000 1364.5500 ;
	    RECT 1012.2000 1364.4000 1013.4000 1364.5500 ;
	    RECT 1115.4000 1363.5000 1116.6000 1371.9000 ;
	    RECT 1119.3000 1371.6000 1125.6000 1372.8000 ;
	    RECT 1132.2001 1372.5000 1133.4000 1379.7001 ;
	    RECT 1134.6000 1373.7001 1135.8000 1379.7001 ;
	    RECT 1137.0000 1372.5000 1138.2001 1379.7001 ;
	    RECT 1139.4000 1373.7001 1140.6000 1379.7001 ;
	    RECT 1119.3000 1371.0000 1120.2001 1371.6000 ;
	    RECT 1117.8000 1369.8000 1120.2001 1371.0000 ;
	    RECT 1124.7001 1370.7001 1133.4000 1371.6000 ;
	    RECT 1121.7001 1369.8000 1123.8000 1370.7001 ;
	    RECT 1121.7001 1369.5000 1131.0000 1369.8000 ;
	    RECT 1122.9000 1368.9000 1131.0000 1369.5000 ;
	    RECT 1129.8000 1368.6000 1131.0000 1368.9000 ;
	    RECT 1132.5000 1369.5000 1133.4000 1370.7001 ;
	    RECT 1134.3000 1370.4000 1138.2001 1371.6000 ;
	    RECT 1141.8000 1370.4000 1143.0000 1379.7001 ;
	    RECT 1144.2001 1375.5000 1145.4000 1379.7001 ;
	    RECT 1146.6000 1375.5000 1147.8000 1379.7001 ;
	    RECT 1149.0000 1375.5000 1150.2001 1379.7001 ;
	    RECT 1151.4000 1373.7001 1152.6000 1379.7001 ;
	    RECT 1146.6000 1371.6000 1152.9000 1372.8000 ;
	    RECT 1153.8000 1371.6000 1155.0000 1379.7001 ;
	    RECT 1156.2001 1373.7001 1157.4000 1379.7001 ;
	    RECT 1158.6000 1372.8000 1159.8000 1379.7001 ;
	    RECT 1161.0000 1373.7001 1162.2001 1379.7001 ;
	    RECT 1158.6000 1371.9000 1162.5000 1372.8000 ;
	    RECT 1163.4000 1372.5000 1164.6000 1379.7001 ;
	    RECT 1165.8000 1373.7001 1167.0000 1379.7001 ;
	    RECT 1293.0000 1373.7001 1294.2001 1379.7001 ;
	    RECT 1295.4000 1374.6000 1296.6000 1379.7001 ;
	    RECT 1295.1000 1373.7001 1296.6000 1374.6000 ;
	    RECT 1297.8000 1373.7001 1299.0000 1380.6000 ;
	    RECT 1295.1000 1372.8000 1296.0000 1373.7001 ;
	    RECT 1300.2001 1372.8000 1301.4000 1379.7001 ;
	    RECT 1302.6000 1373.7001 1303.8000 1379.7001 ;
	    RECT 1305.0000 1375.5000 1306.2001 1379.7001 ;
	    RECT 1307.4000 1375.5000 1308.6000 1379.7001 ;
	    RECT 1153.8000 1370.4000 1157.7001 1371.6000 ;
	    RECT 1144.2001 1369.5000 1145.4000 1369.8000 ;
	    RECT 1132.5000 1368.6000 1145.4000 1369.5000 ;
	    RECT 1149.0000 1369.5000 1150.2001 1369.8000 ;
	    RECT 1161.6000 1369.5000 1162.5000 1371.9000 ;
	    RECT 1293.0000 1371.9000 1296.0000 1372.8000 ;
	    RECT 1163.4000 1371.4501 1164.6000 1371.6000 ;
	    RECT 1235.4000 1371.4501 1236.6000 1371.6000 ;
	    RECT 1163.4000 1370.5500 1236.6000 1371.4501 ;
	    RECT 1163.4000 1370.4000 1164.6000 1370.5500 ;
	    RECT 1235.4000 1370.4000 1236.6000 1370.5500 ;
	    RECT 1149.0000 1368.6000 1162.5000 1369.5000 ;
	    RECT 1120.2001 1367.4000 1121.4000 1368.6000 ;
	    RECT 1125.3000 1367.7001 1126.5000 1368.0000 ;
	    RECT 1122.3000 1366.8000 1160.7001 1367.7001 ;
	    RECT 1159.5000 1366.5000 1160.7001 1366.8000 ;
	    RECT 1161.6000 1365.9000 1162.5000 1368.6000 ;
	    RECT 1163.4000 1368.0000 1164.6000 1369.5000 ;
	    RECT 1163.4000 1366.8000 1164.9000 1368.0000 ;
	    RECT 1117.5000 1365.0000 1124.1000 1365.9000 ;
	    RECT 1117.5000 1364.7001 1118.7001 1365.0000 ;
	    RECT 1125.0000 1364.4000 1126.2001 1365.6000 ;
	    RECT 1127.1000 1365.0000 1152.6000 1365.9000 ;
	    RECT 1161.6000 1365.0000 1162.8000 1365.9000 ;
	    RECT 1151.4000 1364.1000 1152.6000 1365.0000 ;
	    RECT 870.0000 1361.7001 871.2000 1362.0000 ;
	    RECT 870.0000 1360.8000 876.6000 1361.7001 ;
	    RECT 877.8000 1361.4000 879.0000 1362.6000 ;
	    RECT 875.4000 1360.5000 876.6000 1360.8000 ;
	    RECT 877.8000 1360.2001 879.0000 1360.5000 ;
	    RECT 856.2000 1353.3000 857.4000 1359.3000 ;
	    RECT 858.6000 1358.1000 862.2000 1359.3000 ;
	    RECT 865.8000 1358.4000 867.3000 1359.6000 ;
	    RECT 871.8000 1358.4000 872.1000 1359.6000 ;
	    RECT 873.0000 1358.4000 874.2000 1359.6000 ;
	    RECT 875.4000 1359.3000 876.6000 1359.6000 ;
	    RECT 881.1000 1359.3000 882.3000 1362.9000 ;
	    RECT 885.0000 1362.3000 898.2000 1363.5000 ;
	    RECT 890.1000 1360.2001 894.6000 1361.4000 ;
	    RECT 890.1000 1359.3000 891.3000 1360.2001 ;
	    RECT 875.4000 1358.4000 882.3000 1359.3000 ;
	    RECT 861.0000 1353.3000 862.2000 1358.1000 ;
	    RECT 887.4000 1358.1000 891.3000 1359.3000 ;
	    RECT 863.4000 1353.3000 864.6000 1357.5000 ;
	    RECT 865.8000 1353.3000 867.0000 1357.5000 ;
	    RECT 868.2000 1353.3000 869.4000 1357.5000 ;
	    RECT 870.6000 1353.3000 871.8000 1357.5000 ;
	    RECT 873.0000 1353.3000 874.2000 1356.3000 ;
	    RECT 875.4000 1353.3000 876.6000 1357.5000 ;
	    RECT 877.8000 1353.3000 879.0000 1356.3000 ;
	    RECT 880.2000 1353.3000 881.4000 1357.5000 ;
	    RECT 882.6000 1353.3000 883.8000 1357.5000 ;
	    RECT 885.0000 1353.3000 886.2000 1357.5000 ;
	    RECT 887.4000 1353.3000 888.6000 1358.1000 ;
	    RECT 892.2000 1353.3000 893.4000 1359.3000 ;
	    RECT 897.0000 1353.3000 898.2000 1362.3000 ;
	    RECT 909.0000 1362.4501 910.2000 1362.6000 ;
	    RECT 921.0000 1362.4501 922.2000 1362.6000 ;
	    RECT 909.0000 1361.5500 922.2000 1362.4501 ;
	    RECT 909.0000 1361.4000 910.2000 1361.5500 ;
	    RECT 921.0000 1361.4000 922.2000 1361.5500 ;
	    RECT 921.0000 1360.2001 922.2000 1360.5000 ;
	    RECT 923.4000 1359.3000 924.6000 1363.5000 ;
	    RECT 942.6000 1362.4501 943.8000 1362.6000 ;
	    RECT 954.6000 1362.4501 955.8000 1362.6000 ;
	    RECT 942.6000 1361.5500 955.8000 1362.4501 ;
	    RECT 942.6000 1361.4000 943.8000 1361.5500 ;
	    RECT 954.6000 1361.4000 955.8000 1361.5500 ;
	    RECT 959.4000 1362.4501 960.6000 1362.6000 ;
	    RECT 961.8000 1362.4501 963.0000 1362.6000 ;
	    RECT 959.4000 1361.5500 963.0000 1362.4501 ;
	    RECT 959.4000 1361.4000 960.6000 1361.5500 ;
	    RECT 961.8000 1361.4000 963.0000 1361.5500 ;
	    RECT 921.0000 1353.3000 922.2000 1359.3000 ;
	    RECT 923.4000 1358.4000 926.1000 1359.3000 ;
	    RECT 940.2000 1358.4000 941.4000 1359.6000 ;
	    RECT 924.9000 1353.3000 926.1000 1358.4000 ;
	    RECT 940.2000 1357.2001 941.4000 1357.5000 ;
	    RECT 940.2000 1353.3000 941.4000 1356.3000 ;
	    RECT 942.6000 1353.3000 943.8000 1360.5000 ;
	    RECT 957.0000 1358.4000 958.2000 1359.6000 ;
	    RECT 957.0000 1357.2001 958.2000 1357.5000 ;
	    RECT 957.0000 1353.3000 958.2000 1356.3000 ;
	    RECT 959.4000 1353.3000 960.6000 1360.5000 ;
	    RECT 981.0000 1359.3000 982.2000 1363.5000 ;
	    RECT 983.4000 1361.4000 984.6000 1362.6000 ;
	    RECT 1115.4000 1362.3000 1128.6000 1363.5000 ;
	    RECT 1129.5000 1362.9000 1132.5000 1364.1000 ;
	    RECT 1138.2001 1362.9000 1143.0000 1364.1000 ;
	    RECT 983.4000 1360.2001 984.6000 1360.5000 ;
	    RECT 979.5000 1358.4000 982.2000 1359.3000 ;
	    RECT 979.5000 1353.3000 980.7000 1358.4000 ;
	    RECT 983.4000 1353.3000 984.6000 1359.3000 ;
	    RECT 1115.4000 1353.3000 1116.6000 1362.3000 ;
	    RECT 1119.0000 1360.2001 1123.5000 1361.4000 ;
	    RECT 1122.3000 1359.3000 1123.5000 1360.2001 ;
	    RECT 1131.3000 1359.3000 1132.5000 1362.9000 ;
	    RECT 1134.6000 1361.4000 1135.8000 1362.6000 ;
	    RECT 1142.4000 1361.7001 1143.6000 1362.0000 ;
	    RECT 1137.0000 1360.8000 1143.6000 1361.7001 ;
	    RECT 1137.0000 1360.5000 1138.2001 1360.8000 ;
	    RECT 1134.6000 1360.2001 1135.8000 1360.5000 ;
	    RECT 1146.6000 1359.6000 1147.8000 1363.8000 ;
	    RECT 1155.3000 1362.9000 1161.0000 1364.1000 ;
	    RECT 1155.3000 1361.1000 1156.5000 1362.9000 ;
	    RECT 1161.9000 1362.0000 1162.8000 1365.0000 ;
	    RECT 1137.0000 1359.3000 1138.2001 1359.6000 ;
	    RECT 1120.2001 1353.3000 1121.4000 1359.3000 ;
	    RECT 1122.3000 1358.1000 1126.2001 1359.3000 ;
	    RECT 1131.3000 1358.4000 1138.2001 1359.3000 ;
	    RECT 1139.4000 1358.4000 1140.6000 1359.6000 ;
	    RECT 1141.5000 1358.4000 1141.8000 1359.6000 ;
	    RECT 1146.3000 1358.4000 1147.8000 1359.6000 ;
	    RECT 1153.8000 1360.2001 1156.5000 1361.1000 ;
	    RECT 1161.0000 1361.1000 1162.8000 1362.0000 ;
	    RECT 1153.8000 1359.3000 1155.0000 1360.2001 ;
	    RECT 1125.0000 1353.3000 1126.2001 1358.1000 ;
	    RECT 1151.4000 1358.1000 1155.0000 1359.3000 ;
	    RECT 1127.4000 1353.3000 1128.6000 1357.5000 ;
	    RECT 1129.8000 1353.3000 1131.0000 1357.5000 ;
	    RECT 1132.2001 1353.3000 1133.4000 1357.5000 ;
	    RECT 1134.6000 1353.3000 1135.8000 1356.3000 ;
	    RECT 1137.0000 1353.3000 1138.2001 1357.5000 ;
	    RECT 1139.4000 1353.3000 1140.6000 1356.3000 ;
	    RECT 1141.8000 1353.3000 1143.0000 1357.5000 ;
	    RECT 1144.2001 1353.3000 1145.4000 1357.5000 ;
	    RECT 1146.6000 1353.3000 1147.8000 1357.5000 ;
	    RECT 1149.0000 1353.3000 1150.2001 1357.5000 ;
	    RECT 1151.4000 1353.3000 1152.6000 1358.1000 ;
	    RECT 1156.2001 1353.3000 1157.4000 1359.3000 ;
	    RECT 1161.0000 1353.3000 1162.2001 1361.1000 ;
	    RECT 1163.7001 1360.2001 1164.9000 1366.8000 ;
	    RECT 1163.4000 1359.0000 1164.9000 1360.2001 ;
	    RECT 1293.0000 1363.5000 1294.2001 1371.9000 ;
	    RECT 1296.9000 1371.6000 1303.2001 1372.8000 ;
	    RECT 1309.8000 1372.5000 1311.0000 1379.7001 ;
	    RECT 1312.2001 1373.7001 1313.4000 1379.7001 ;
	    RECT 1314.6000 1372.5000 1315.8000 1379.7001 ;
	    RECT 1317.0000 1373.7001 1318.2001 1379.7001 ;
	    RECT 1296.9000 1371.0000 1297.8000 1371.6000 ;
	    RECT 1295.4000 1369.8000 1297.8000 1371.0000 ;
	    RECT 1302.3000 1370.7001 1311.0000 1371.6000 ;
	    RECT 1299.3000 1369.8000 1301.4000 1370.7001 ;
	    RECT 1299.3000 1369.5000 1308.6000 1369.8000 ;
	    RECT 1300.5000 1368.9000 1308.6000 1369.5000 ;
	    RECT 1307.4000 1368.6000 1308.6000 1368.9000 ;
	    RECT 1310.1000 1369.5000 1311.0000 1370.7001 ;
	    RECT 1311.9000 1370.4000 1315.8000 1371.6000 ;
	    RECT 1319.4000 1370.4000 1320.6000 1379.7001 ;
	    RECT 1321.8000 1375.5000 1323.0000 1379.7001 ;
	    RECT 1324.2001 1375.5000 1325.4000 1379.7001 ;
	    RECT 1326.6000 1375.5000 1327.8000 1379.7001 ;
	    RECT 1329.0000 1373.7001 1330.2001 1379.7001 ;
	    RECT 1324.2001 1371.6000 1330.5000 1372.8000 ;
	    RECT 1331.4000 1371.6000 1332.6000 1379.7001 ;
	    RECT 1333.8000 1373.7001 1335.0000 1379.7001 ;
	    RECT 1336.2001 1372.8000 1337.4000 1379.7001 ;
	    RECT 1338.6000 1373.7001 1339.8000 1379.7001 ;
	    RECT 1336.2001 1371.9000 1340.1000 1372.8000 ;
	    RECT 1341.0000 1372.5000 1342.2001 1379.7001 ;
	    RECT 1343.4000 1373.7001 1344.6000 1379.7001 ;
	    RECT 1377.0000 1379.4000 1378.2001 1380.6000 ;
	    RECT 1475.4000 1373.7001 1476.6000 1379.7001 ;
	    RECT 1477.8000 1374.6000 1479.0000 1379.7001 ;
	    RECT 1477.5000 1373.7001 1479.0000 1374.6000 ;
	    RECT 1480.2001 1373.7001 1481.4000 1380.6000 ;
	    RECT 1477.5000 1372.8000 1478.4000 1373.7001 ;
	    RECT 1482.6000 1372.8000 1483.8000 1379.7001 ;
	    RECT 1485.0000 1373.7001 1486.2001 1379.7001 ;
	    RECT 1487.4000 1375.5000 1488.6000 1379.7001 ;
	    RECT 1489.8000 1375.5000 1491.0000 1379.7001 ;
	    RECT 1331.4000 1370.4000 1335.3000 1371.6000 ;
	    RECT 1321.8000 1369.5000 1323.0000 1369.8000 ;
	    RECT 1310.1000 1368.6000 1323.0000 1369.5000 ;
	    RECT 1326.6000 1369.5000 1327.8000 1369.8000 ;
	    RECT 1339.2001 1369.5000 1340.1000 1371.9000 ;
	    RECT 1475.4000 1371.9000 1478.4000 1372.8000 ;
	    RECT 1341.0000 1371.4501 1342.2001 1371.6000 ;
	    RECT 1345.8000 1371.4501 1347.0000 1371.6000 ;
	    RECT 1341.0000 1370.5500 1347.0000 1371.4501 ;
	    RECT 1341.0000 1370.4000 1342.2001 1370.5500 ;
	    RECT 1345.8000 1370.4000 1347.0000 1370.5500 ;
	    RECT 1326.6000 1368.6000 1340.1000 1369.5000 ;
	    RECT 1297.8000 1367.4000 1299.0000 1368.6000 ;
	    RECT 1302.9000 1367.7001 1304.1000 1368.0000 ;
	    RECT 1299.9000 1366.8000 1338.3000 1367.7001 ;
	    RECT 1337.1000 1366.5000 1338.3000 1366.8000 ;
	    RECT 1339.2001 1365.9000 1340.1000 1368.6000 ;
	    RECT 1341.0000 1368.0000 1342.2001 1369.5000 ;
	    RECT 1341.0000 1366.8000 1342.5000 1368.0000 ;
	    RECT 1295.1000 1365.0000 1301.7001 1365.9000 ;
	    RECT 1295.1000 1364.7001 1296.3000 1365.0000 ;
	    RECT 1302.6000 1364.4000 1303.8000 1365.6000 ;
	    RECT 1304.7001 1365.0000 1330.2001 1365.9000 ;
	    RECT 1339.2001 1365.0000 1340.4000 1365.9000 ;
	    RECT 1329.0000 1364.1000 1330.2001 1365.0000 ;
	    RECT 1293.0000 1362.3000 1306.2001 1363.5000 ;
	    RECT 1307.1000 1362.9000 1310.1000 1364.1000 ;
	    RECT 1315.8000 1362.9000 1320.6000 1364.1000 ;
	    RECT 1163.4000 1353.3000 1164.6000 1359.0000 ;
	    RECT 1165.8000 1353.3000 1167.0000 1356.3000 ;
	    RECT 1293.0000 1353.3000 1294.2001 1362.3000 ;
	    RECT 1296.6000 1360.2001 1301.1000 1361.4000 ;
	    RECT 1299.9000 1359.3000 1301.1000 1360.2001 ;
	    RECT 1308.9000 1359.3000 1310.1000 1362.9000 ;
	    RECT 1312.2001 1361.4000 1313.4000 1362.6000 ;
	    RECT 1320.0000 1361.7001 1321.2001 1362.0000 ;
	    RECT 1314.6000 1360.8000 1321.2001 1361.7001 ;
	    RECT 1314.6000 1360.5000 1315.8000 1360.8000 ;
	    RECT 1312.2001 1360.2001 1313.4000 1360.5000 ;
	    RECT 1324.2001 1359.6000 1325.4000 1363.8000 ;
	    RECT 1332.9000 1362.9000 1338.6000 1364.1000 ;
	    RECT 1332.9000 1361.1000 1334.1000 1362.9000 ;
	    RECT 1339.5000 1362.0000 1340.4000 1365.0000 ;
	    RECT 1314.6000 1359.3000 1315.8000 1359.6000 ;
	    RECT 1297.8000 1353.3000 1299.0000 1359.3000 ;
	    RECT 1299.9000 1358.1000 1303.8000 1359.3000 ;
	    RECT 1308.9000 1358.4000 1315.8000 1359.3000 ;
	    RECT 1317.0000 1358.4000 1318.2001 1359.6000 ;
	    RECT 1319.1000 1358.4000 1319.4000 1359.6000 ;
	    RECT 1323.9000 1358.4000 1325.4000 1359.6000 ;
	    RECT 1331.4000 1360.2001 1334.1000 1361.1000 ;
	    RECT 1338.6000 1361.1000 1340.4000 1362.0000 ;
	    RECT 1331.4000 1359.3000 1332.6000 1360.2001 ;
	    RECT 1302.6000 1353.3000 1303.8000 1358.1000 ;
	    RECT 1329.0000 1358.1000 1332.6000 1359.3000 ;
	    RECT 1305.0000 1353.3000 1306.2001 1357.5000 ;
	    RECT 1307.4000 1353.3000 1308.6000 1357.5000 ;
	    RECT 1309.8000 1353.3000 1311.0000 1357.5000 ;
	    RECT 1312.2001 1353.3000 1313.4000 1356.3000 ;
	    RECT 1314.6000 1353.3000 1315.8000 1357.5000 ;
	    RECT 1317.0000 1353.3000 1318.2001 1356.3000 ;
	    RECT 1319.4000 1353.3000 1320.6000 1357.5000 ;
	    RECT 1321.8000 1353.3000 1323.0000 1357.5000 ;
	    RECT 1324.2001 1353.3000 1325.4000 1357.5000 ;
	    RECT 1326.6000 1353.3000 1327.8000 1357.5000 ;
	    RECT 1329.0000 1353.3000 1330.2001 1358.1000 ;
	    RECT 1333.8000 1353.3000 1335.0000 1359.3000 ;
	    RECT 1338.6000 1353.3000 1339.8000 1361.1000 ;
	    RECT 1341.3000 1360.2001 1342.5000 1366.8000 ;
	    RECT 1341.0000 1359.0000 1342.5000 1360.2001 ;
	    RECT 1475.4000 1363.5000 1476.6000 1371.9000 ;
	    RECT 1479.3000 1371.6000 1485.6000 1372.8000 ;
	    RECT 1492.2001 1372.5000 1493.4000 1379.7001 ;
	    RECT 1494.6000 1373.7001 1495.8000 1379.7001 ;
	    RECT 1497.0000 1372.5000 1498.2001 1379.7001 ;
	    RECT 1499.4000 1373.7001 1500.6000 1379.7001 ;
	    RECT 1479.3000 1371.0000 1480.2001 1371.6000 ;
	    RECT 1477.8000 1369.8000 1480.2001 1371.0000 ;
	    RECT 1484.7001 1370.7001 1493.4000 1371.6000 ;
	    RECT 1481.7001 1369.8000 1483.8000 1370.7001 ;
	    RECT 1481.7001 1369.5000 1491.0000 1369.8000 ;
	    RECT 1482.9000 1368.9000 1491.0000 1369.5000 ;
	    RECT 1489.8000 1368.6000 1491.0000 1368.9000 ;
	    RECT 1492.5000 1369.5000 1493.4000 1370.7001 ;
	    RECT 1494.3000 1370.4000 1498.2001 1371.6000 ;
	    RECT 1501.8000 1370.4000 1503.0000 1379.7001 ;
	    RECT 1504.2001 1375.5000 1505.4000 1379.7001 ;
	    RECT 1506.6000 1375.5000 1507.8000 1379.7001 ;
	    RECT 1509.0000 1375.5000 1510.2001 1379.7001 ;
	    RECT 1511.4000 1373.7001 1512.6000 1379.7001 ;
	    RECT 1506.6000 1371.6000 1512.9000 1372.8000 ;
	    RECT 1513.8000 1371.6000 1515.0000 1379.7001 ;
	    RECT 1516.2001 1373.7001 1517.4000 1379.7001 ;
	    RECT 1518.6000 1372.8000 1519.8000 1379.7001 ;
	    RECT 1521.0000 1373.7001 1522.2001 1379.7001 ;
	    RECT 1518.6000 1371.9000 1522.5000 1372.8000 ;
	    RECT 1523.4000 1372.5000 1524.6000 1379.7001 ;
	    RECT 1525.8000 1373.7001 1527.0000 1379.7001 ;
	    RECT 1549.8000 1373.7001 1551.0000 1379.7001 ;
	    RECT 1552.2001 1374.3000 1553.4000 1379.7001 ;
	    RECT 1550.1000 1373.4000 1551.0000 1373.7001 ;
	    RECT 1554.6000 1373.7001 1555.8000 1379.7001 ;
	    RECT 1557.0000 1373.7001 1558.2001 1379.7001 ;
	    RECT 1554.6000 1373.4000 1555.5000 1373.7001 ;
	    RECT 1550.1000 1372.5000 1555.5000 1373.4000 ;
	    RECT 1513.8000 1370.4000 1517.7001 1371.6000 ;
	    RECT 1504.2001 1369.5000 1505.4000 1369.8000 ;
	    RECT 1492.5000 1368.6000 1505.4000 1369.5000 ;
	    RECT 1509.0000 1369.5000 1510.2001 1369.8000 ;
	    RECT 1521.6000 1369.5000 1522.5000 1371.9000 ;
	    RECT 1523.4000 1370.4000 1524.6000 1371.6000 ;
	    RECT 1550.1000 1369.5000 1551.0000 1372.5000 ;
	    RECT 1552.2001 1371.4501 1553.4000 1371.6000 ;
	    RECT 1559.4000 1371.4501 1560.6000 1371.6000 ;
	    RECT 1552.2001 1370.5500 1560.6000 1371.4501 ;
	    RECT 1552.2001 1370.4000 1553.4000 1370.5500 ;
	    RECT 1559.4000 1370.4000 1560.6000 1370.5500 ;
	    RECT 1509.0000 1368.6000 1522.5000 1369.5000 ;
	    RECT 1480.2001 1367.4000 1481.4000 1368.6000 ;
	    RECT 1485.3000 1367.7001 1486.5000 1368.0000 ;
	    RECT 1482.3000 1366.8000 1520.7001 1367.7001 ;
	    RECT 1519.5000 1366.5000 1520.7001 1366.8000 ;
	    RECT 1521.6000 1365.9000 1522.5000 1368.6000 ;
	    RECT 1523.4000 1368.0000 1524.6000 1369.5000 ;
	    RECT 1552.2001 1369.2001 1553.4000 1369.5000 ;
	    RECT 1545.0000 1368.4501 1546.2001 1368.6000 ;
	    RECT 1549.8000 1368.4501 1551.0000 1368.6000 ;
	    RECT 1523.4000 1366.8000 1524.9000 1368.0000 ;
	    RECT 1545.0000 1367.5500 1551.0000 1368.4501 ;
	    RECT 1545.0000 1367.4000 1546.2001 1367.5500 ;
	    RECT 1549.8000 1367.4000 1551.0000 1367.5500 ;
	    RECT 1557.0000 1368.4501 1558.2001 1368.6000 ;
	    RECT 1561.8000 1368.4501 1563.0000 1368.6000 ;
	    RECT 1557.0000 1367.5500 1563.0000 1368.4501 ;
	    RECT 1557.0000 1367.4000 1558.2001 1367.5500 ;
	    RECT 1561.8000 1367.4000 1563.0000 1367.5500 ;
	    RECT 1477.5000 1365.0000 1484.1000 1365.9000 ;
	    RECT 1477.5000 1364.7001 1478.7001 1365.0000 ;
	    RECT 1485.0000 1364.4000 1486.2001 1365.6000 ;
	    RECT 1487.1000 1365.0000 1512.6000 1365.9000 ;
	    RECT 1521.6000 1365.0000 1522.8000 1365.9000 ;
	    RECT 1511.4000 1364.1000 1512.6000 1365.0000 ;
	    RECT 1475.4000 1362.3000 1488.6000 1363.5000 ;
	    RECT 1489.5000 1362.9000 1492.5000 1364.1000 ;
	    RECT 1498.2001 1362.9000 1503.0000 1364.1000 ;
	    RECT 1341.0000 1353.3000 1342.2001 1359.0000 ;
	    RECT 1343.4000 1353.3000 1344.6000 1356.3000 ;
	    RECT 1475.4000 1353.3000 1476.6000 1362.3000 ;
	    RECT 1479.0000 1360.2001 1483.5000 1361.4000 ;
	    RECT 1482.3000 1359.3000 1483.5000 1360.2001 ;
	    RECT 1491.3000 1359.3000 1492.5000 1362.9000 ;
	    RECT 1494.6000 1361.4000 1495.8000 1362.6000 ;
	    RECT 1502.4000 1361.7001 1503.6000 1362.0000 ;
	    RECT 1497.0000 1360.8000 1503.6000 1361.7001 ;
	    RECT 1497.0000 1360.5000 1498.2001 1360.8000 ;
	    RECT 1494.6000 1360.2001 1495.8000 1360.5000 ;
	    RECT 1506.6000 1359.6000 1507.8000 1363.8000 ;
	    RECT 1515.3000 1362.9000 1521.0000 1364.1000 ;
	    RECT 1515.3000 1361.1000 1516.5000 1362.9000 ;
	    RECT 1521.9000 1362.0000 1522.8000 1365.0000 ;
	    RECT 1497.0000 1359.3000 1498.2001 1359.6000 ;
	    RECT 1480.2001 1353.3000 1481.4000 1359.3000 ;
	    RECT 1482.3000 1358.1000 1486.2001 1359.3000 ;
	    RECT 1491.3000 1358.4000 1498.2001 1359.3000 ;
	    RECT 1499.4000 1358.4000 1500.6000 1359.6000 ;
	    RECT 1501.5000 1358.4000 1501.8000 1359.6000 ;
	    RECT 1506.3000 1358.4000 1507.8000 1359.6000 ;
	    RECT 1513.8000 1360.2001 1516.5000 1361.1000 ;
	    RECT 1521.0000 1361.1000 1522.8000 1362.0000 ;
	    RECT 1513.8000 1359.3000 1515.0000 1360.2001 ;
	    RECT 1485.0000 1353.3000 1486.2001 1358.1000 ;
	    RECT 1511.4000 1358.1000 1515.0000 1359.3000 ;
	    RECT 1487.4000 1353.3000 1488.6000 1357.5000 ;
	    RECT 1489.8000 1353.3000 1491.0000 1357.5000 ;
	    RECT 1492.2001 1353.3000 1493.4000 1357.5000 ;
	    RECT 1494.6000 1353.3000 1495.8000 1356.3000 ;
	    RECT 1497.0000 1353.3000 1498.2001 1357.5000 ;
	    RECT 1499.4000 1353.3000 1500.6000 1356.3000 ;
	    RECT 1501.8000 1353.3000 1503.0000 1357.5000 ;
	    RECT 1504.2001 1353.3000 1505.4000 1357.5000 ;
	    RECT 1506.6000 1353.3000 1507.8000 1357.5000 ;
	    RECT 1509.0000 1353.3000 1510.2001 1357.5000 ;
	    RECT 1511.4000 1353.3000 1512.6000 1358.1000 ;
	    RECT 1516.2001 1353.3000 1517.4000 1359.3000 ;
	    RECT 1521.0000 1353.3000 1522.2001 1361.1000 ;
	    RECT 1523.7001 1360.2001 1524.9000 1366.8000 ;
	    RECT 1550.1000 1362.6000 1551.0000 1366.5000 ;
	    RECT 1557.0000 1366.2001 1558.2001 1366.5000 ;
	    RECT 1553.4000 1364.4000 1553.7001 1365.6000 ;
	    RECT 1554.6000 1364.4000 1555.8000 1365.6000 ;
	    RECT 1550.1000 1362.3000 1552.5000 1362.6000 ;
	    RECT 1550.1000 1361.7001 1552.8000 1362.3000 ;
	    RECT 1523.4000 1359.0000 1524.9000 1360.2001 ;
	    RECT 1523.4000 1353.3000 1524.6000 1359.0000 ;
	    RECT 1525.8000 1353.3000 1527.0000 1356.3000 ;
	    RECT 1551.6000 1353.3000 1552.8000 1361.7001 ;
	    RECT 1557.0000 1353.3000 1558.2001 1362.3000 ;
	    RECT 1.2000 1350.6000 1569.0000 1352.4000 ;
	    RECT 126.6000 1346.7001 127.8000 1349.7001 ;
	    RECT 129.0000 1344.0000 130.2000 1349.7001 ;
	    RECT 128.7000 1342.8000 130.2000 1344.0000 ;
	    RECT 128.7000 1336.2001 129.9000 1342.8000 ;
	    RECT 131.4000 1341.9000 132.6000 1349.7001 ;
	    RECT 136.2000 1343.7001 137.4000 1349.7001 ;
	    RECT 141.0000 1344.9000 142.2000 1349.7001 ;
	    RECT 143.4000 1345.5000 144.6000 1349.7001 ;
	    RECT 145.8000 1345.5000 147.0000 1349.7001 ;
	    RECT 148.2000 1345.5000 149.4000 1349.7001 ;
	    RECT 150.6000 1345.5000 151.8000 1349.7001 ;
	    RECT 153.0000 1346.7001 154.2000 1349.7001 ;
	    RECT 155.4000 1345.5000 156.6000 1349.7001 ;
	    RECT 157.8000 1346.7001 159.0000 1349.7001 ;
	    RECT 160.2000 1345.5000 161.4000 1349.7001 ;
	    RECT 162.6000 1345.5000 163.8000 1349.7001 ;
	    RECT 165.0000 1345.5000 166.2000 1349.7001 ;
	    RECT 138.6000 1343.7001 142.2000 1344.9000 ;
	    RECT 167.4000 1344.9000 168.6000 1349.7001 ;
	    RECT 138.6000 1342.8000 139.8000 1343.7001 ;
	    RECT 130.8000 1341.0000 132.6000 1341.9000 ;
	    RECT 137.1000 1341.9000 139.8000 1342.8000 ;
	    RECT 145.8000 1343.4000 147.3000 1344.6000 ;
	    RECT 151.8000 1343.4000 152.1000 1344.6000 ;
	    RECT 153.0000 1343.4000 154.2000 1344.6000 ;
	    RECT 155.4000 1343.7001 162.3000 1344.6000 ;
	    RECT 167.4000 1343.7001 171.3000 1344.9000 ;
	    RECT 172.2000 1343.7001 173.4000 1349.7001 ;
	    RECT 155.4000 1343.4000 156.6000 1343.7001 ;
	    RECT 130.8000 1338.0000 131.7000 1341.0000 ;
	    RECT 137.1000 1340.1000 138.3000 1341.9000 ;
	    RECT 132.6000 1338.9000 138.3000 1340.1000 ;
	    RECT 145.8000 1339.2001 147.0000 1343.4000 ;
	    RECT 157.8000 1342.5000 159.0000 1342.8000 ;
	    RECT 155.4000 1342.2001 156.6000 1342.5000 ;
	    RECT 150.0000 1341.3000 156.6000 1342.2001 ;
	    RECT 150.0000 1341.0000 151.2000 1341.3000 ;
	    RECT 157.8000 1340.4000 159.0000 1341.6000 ;
	    RECT 161.1000 1340.1000 162.3000 1343.7001 ;
	    RECT 170.1000 1342.8000 171.3000 1343.7001 ;
	    RECT 170.1000 1341.6000 174.6000 1342.8000 ;
	    RECT 177.0000 1340.7001 178.2000 1349.7001 ;
	    RECT 191.4000 1346.7001 192.6000 1349.7001 ;
	    RECT 191.4000 1345.5000 192.6000 1345.8000 ;
	    RECT 179.4000 1344.4501 180.6000 1344.6000 ;
	    RECT 191.4000 1344.4501 192.6000 1344.6000 ;
	    RECT 179.4000 1343.5500 192.6000 1344.4501 ;
	    RECT 179.4000 1343.4000 180.6000 1343.5500 ;
	    RECT 191.4000 1343.4000 192.6000 1343.5500 ;
	    RECT 193.8000 1342.5000 195.0000 1349.7001 ;
	    RECT 325.8000 1346.7001 327.0000 1349.7001 ;
	    RECT 328.2000 1344.0000 329.4000 1349.7001 ;
	    RECT 327.9000 1342.8000 329.4000 1344.0000 ;
	    RECT 150.6000 1338.9000 155.4000 1340.1000 ;
	    RECT 161.1000 1338.9000 164.1000 1340.1000 ;
	    RECT 165.0000 1339.5000 178.2000 1340.7001 ;
	    RECT 181.8000 1341.4501 183.0000 1341.6000 ;
	    RECT 193.8000 1341.4501 195.0000 1341.6000 ;
	    RECT 181.8000 1340.5500 195.0000 1341.4501 ;
	    RECT 181.8000 1340.4000 183.0000 1340.5500 ;
	    RECT 193.8000 1340.4000 195.0000 1340.5500 ;
	    RECT 141.0000 1338.0000 142.2000 1338.9000 ;
	    RECT 130.8000 1337.1000 132.0000 1338.0000 ;
	    RECT 141.0000 1337.1000 166.5000 1338.0000 ;
	    RECT 167.4000 1337.4000 168.6000 1338.6000 ;
	    RECT 174.9000 1338.0000 176.1000 1338.3000 ;
	    RECT 169.5000 1337.1000 176.1000 1338.0000 ;
	    RECT 128.7000 1335.0000 130.2000 1336.2001 ;
	    RECT 129.0000 1333.5000 130.2000 1335.0000 ;
	    RECT 131.1000 1334.4000 132.0000 1337.1000 ;
	    RECT 132.9000 1336.2001 134.1000 1336.5000 ;
	    RECT 132.9000 1335.3000 171.3000 1336.2001 ;
	    RECT 167.1000 1335.0000 168.3000 1335.3000 ;
	    RECT 172.2000 1334.4000 173.4000 1335.6000 ;
	    RECT 131.1000 1333.5000 144.6000 1334.4000 ;
	    RECT 126.6000 1332.4501 127.8000 1332.6000 ;
	    RECT 129.0000 1332.4501 130.2000 1332.6000 ;
	    RECT 126.6000 1331.5500 130.2000 1332.4501 ;
	    RECT 126.6000 1331.4000 127.8000 1331.5500 ;
	    RECT 129.0000 1331.4000 130.2000 1331.5500 ;
	    RECT 131.1000 1331.1000 132.0000 1333.5000 ;
	    RECT 143.4000 1333.2001 144.6000 1333.5000 ;
	    RECT 148.2000 1333.5000 161.1000 1334.4000 ;
	    RECT 148.2000 1333.2001 149.4000 1333.5000 ;
	    RECT 135.9000 1331.4000 139.8000 1332.6000 ;
	    RECT 126.6000 1323.3000 127.8000 1329.3000 ;
	    RECT 129.0000 1323.3000 130.2000 1330.5000 ;
	    RECT 131.1000 1330.2001 135.0000 1331.1000 ;
	    RECT 131.4000 1323.3000 132.6000 1329.3000 ;
	    RECT 133.8000 1323.3000 135.0000 1330.2001 ;
	    RECT 136.2000 1323.3000 137.4000 1329.3000 ;
	    RECT 138.6000 1323.3000 139.8000 1331.4000 ;
	    RECT 140.7000 1330.2001 147.0000 1331.4000 ;
	    RECT 141.0000 1323.3000 142.2000 1329.3000 ;
	    RECT 143.4000 1323.3000 144.6000 1327.5000 ;
	    RECT 145.8000 1323.3000 147.0000 1327.5000 ;
	    RECT 148.2000 1323.3000 149.4000 1327.5000 ;
	    RECT 150.6000 1323.3000 151.8000 1332.6000 ;
	    RECT 155.4000 1331.4000 159.3000 1332.6000 ;
	    RECT 160.2000 1332.3000 161.1000 1333.5000 ;
	    RECT 162.6000 1334.1000 163.8000 1334.4000 ;
	    RECT 162.6000 1333.5000 170.7000 1334.1000 ;
	    RECT 162.6000 1333.2001 171.9000 1333.5000 ;
	    RECT 169.8000 1332.3000 171.9000 1333.2001 ;
	    RECT 160.2000 1331.4000 168.9000 1332.3000 ;
	    RECT 173.4000 1332.0000 175.8000 1333.2001 ;
	    RECT 173.4000 1331.4000 174.3000 1332.0000 ;
	    RECT 153.0000 1323.3000 154.2000 1329.3000 ;
	    RECT 155.4000 1323.3000 156.6000 1330.5000 ;
	    RECT 157.8000 1323.3000 159.0000 1329.3000 ;
	    RECT 160.2000 1323.3000 161.4000 1330.5000 ;
	    RECT 168.0000 1330.2001 174.3000 1331.4000 ;
	    RECT 177.0000 1331.1000 178.2000 1339.5000 ;
	    RECT 175.2000 1330.2001 178.2000 1331.1000 ;
	    RECT 162.6000 1323.3000 163.8000 1327.5000 ;
	    RECT 165.0000 1323.3000 166.2000 1327.5000 ;
	    RECT 167.4000 1323.3000 168.6000 1329.3000 ;
	    RECT 169.8000 1323.3000 171.0000 1330.2001 ;
	    RECT 175.2000 1329.3000 176.1000 1330.2001 ;
	    RECT 172.2000 1322.4000 173.4000 1329.3000 ;
	    RECT 174.6000 1328.4000 176.1000 1329.3000 ;
	    RECT 174.6000 1323.3000 175.8000 1328.4000 ;
	    RECT 177.0000 1323.3000 178.2000 1329.3000 ;
	    RECT 191.4000 1323.3000 192.6000 1329.3000 ;
	    RECT 193.8000 1323.3000 195.0000 1339.5000 ;
	    RECT 327.9000 1336.2001 329.1000 1342.8000 ;
	    RECT 330.6000 1341.9000 331.8000 1349.7001 ;
	    RECT 335.4000 1343.7001 336.6000 1349.7001 ;
	    RECT 340.2000 1344.9000 341.4000 1349.7001 ;
	    RECT 342.6000 1345.5000 343.8000 1349.7001 ;
	    RECT 345.0000 1345.5000 346.2000 1349.7001 ;
	    RECT 347.4000 1345.5000 348.6000 1349.7001 ;
	    RECT 349.8000 1345.5000 351.0000 1349.7001 ;
	    RECT 352.2000 1346.7001 353.4000 1349.7001 ;
	    RECT 354.6000 1345.5000 355.8000 1349.7001 ;
	    RECT 357.0000 1346.7001 358.2000 1349.7001 ;
	    RECT 359.4000 1345.5000 360.6000 1349.7001 ;
	    RECT 361.8000 1345.5000 363.0000 1349.7001 ;
	    RECT 364.2000 1345.5000 365.4000 1349.7001 ;
	    RECT 337.8000 1343.7001 341.4000 1344.9000 ;
	    RECT 366.6000 1344.9000 367.8000 1349.7001 ;
	    RECT 337.8000 1342.8000 339.0000 1343.7001 ;
	    RECT 330.0000 1341.0000 331.8000 1341.9000 ;
	    RECT 336.3000 1341.9000 339.0000 1342.8000 ;
	    RECT 345.0000 1343.4000 346.5000 1344.6000 ;
	    RECT 351.0000 1343.4000 351.3000 1344.6000 ;
	    RECT 352.2000 1343.4000 353.4000 1344.6000 ;
	    RECT 354.6000 1343.7001 361.5000 1344.6000 ;
	    RECT 366.6000 1343.7001 370.5000 1344.9000 ;
	    RECT 371.4000 1343.7001 372.6000 1349.7001 ;
	    RECT 354.6000 1343.4000 355.8000 1343.7001 ;
	    RECT 330.0000 1338.0000 330.9000 1341.0000 ;
	    RECT 336.3000 1340.1000 337.5000 1341.9000 ;
	    RECT 331.8000 1338.9000 337.5000 1340.1000 ;
	    RECT 345.0000 1339.2001 346.2000 1343.4000 ;
	    RECT 357.0000 1342.5000 358.2000 1342.8000 ;
	    RECT 354.6000 1342.2001 355.8000 1342.5000 ;
	    RECT 349.2000 1341.3000 355.8000 1342.2001 ;
	    RECT 349.2000 1341.0000 350.4000 1341.3000 ;
	    RECT 357.0000 1340.4000 358.2000 1341.6000 ;
	    RECT 360.3000 1340.1000 361.5000 1343.7001 ;
	    RECT 369.3000 1342.8000 370.5000 1343.7001 ;
	    RECT 369.3000 1341.6000 373.8000 1342.8000 ;
	    RECT 376.2000 1340.7001 377.4000 1349.7001 ;
	    RECT 510.6000 1346.7001 511.8000 1349.7001 ;
	    RECT 513.0000 1344.0000 514.2000 1349.7001 ;
	    RECT 349.8000 1338.9000 354.6000 1340.1000 ;
	    RECT 360.3000 1338.9000 363.3000 1340.1000 ;
	    RECT 364.2000 1339.5000 377.4000 1340.7001 ;
	    RECT 340.2000 1338.0000 341.4000 1338.9000 ;
	    RECT 330.0000 1337.1000 331.2000 1338.0000 ;
	    RECT 340.2000 1337.1000 365.7000 1338.0000 ;
	    RECT 366.6000 1337.4000 367.8000 1338.6000 ;
	    RECT 374.1000 1338.0000 375.3000 1338.3000 ;
	    RECT 368.7000 1337.1000 375.3000 1338.0000 ;
	    RECT 327.9000 1335.0000 329.4000 1336.2001 ;
	    RECT 328.2000 1333.5000 329.4000 1335.0000 ;
	    RECT 330.3000 1334.4000 331.2000 1337.1000 ;
	    RECT 332.1000 1336.2001 333.3000 1336.5000 ;
	    RECT 332.1000 1335.3000 370.5000 1336.2001 ;
	    RECT 366.3000 1335.0000 367.5000 1335.3000 ;
	    RECT 371.4000 1334.4000 372.6000 1335.6000 ;
	    RECT 330.3000 1333.5000 343.8000 1334.4000 ;
	    RECT 244.2000 1332.4501 245.4000 1332.6000 ;
	    RECT 263.4000 1332.4501 264.6000 1332.6000 ;
	    RECT 328.2000 1332.4501 329.4000 1332.6000 ;
	    RECT 244.2000 1331.5500 329.4000 1332.4501 ;
	    RECT 244.2000 1331.4000 245.4000 1331.5500 ;
	    RECT 263.4000 1331.4000 264.6000 1331.5500 ;
	    RECT 328.2000 1331.4000 329.4000 1331.5500 ;
	    RECT 330.3000 1331.1000 331.2000 1333.5000 ;
	    RECT 342.6000 1333.2001 343.8000 1333.5000 ;
	    RECT 347.4000 1333.5000 360.3000 1334.4000 ;
	    RECT 347.4000 1333.2001 348.6000 1333.5000 ;
	    RECT 335.1000 1331.4000 339.0000 1332.6000 ;
	    RECT 325.8000 1323.3000 327.0000 1329.3000 ;
	    RECT 328.2000 1323.3000 329.4000 1330.5000 ;
	    RECT 330.3000 1330.2001 334.2000 1331.1000 ;
	    RECT 330.6000 1323.3000 331.8000 1329.3000 ;
	    RECT 333.0000 1323.3000 334.2000 1330.2001 ;
	    RECT 335.4000 1323.3000 336.6000 1329.3000 ;
	    RECT 337.8000 1323.3000 339.0000 1331.4000 ;
	    RECT 339.9000 1330.2001 346.2000 1331.4000 ;
	    RECT 340.2000 1323.3000 341.4000 1329.3000 ;
	    RECT 342.6000 1323.3000 343.8000 1327.5000 ;
	    RECT 345.0000 1323.3000 346.2000 1327.5000 ;
	    RECT 347.4000 1323.3000 348.6000 1327.5000 ;
	    RECT 349.8000 1323.3000 351.0000 1332.6000 ;
	    RECT 354.6000 1331.4000 358.5000 1332.6000 ;
	    RECT 359.4000 1332.3000 360.3000 1333.5000 ;
	    RECT 361.8000 1334.1000 363.0000 1334.4000 ;
	    RECT 361.8000 1333.5000 369.9000 1334.1000 ;
	    RECT 361.8000 1333.2001 371.1000 1333.5000 ;
	    RECT 369.0000 1332.3000 371.1000 1333.2001 ;
	    RECT 359.4000 1331.4000 368.1000 1332.3000 ;
	    RECT 372.6000 1332.0000 375.0000 1333.2001 ;
	    RECT 372.6000 1331.4000 373.5000 1332.0000 ;
	    RECT 352.2000 1323.3000 353.4000 1329.3000 ;
	    RECT 354.6000 1323.3000 355.8000 1330.5000 ;
	    RECT 357.0000 1323.3000 358.2000 1329.3000 ;
	    RECT 359.4000 1323.3000 360.6000 1330.5000 ;
	    RECT 367.2000 1330.2001 373.5000 1331.4000 ;
	    RECT 376.2000 1331.1000 377.4000 1339.5000 ;
	    RECT 512.7000 1342.8000 514.2000 1344.0000 ;
	    RECT 512.7000 1336.2001 513.9000 1342.8000 ;
	    RECT 515.4000 1341.9000 516.6000 1349.7001 ;
	    RECT 520.2000 1343.7001 521.4000 1349.7001 ;
	    RECT 525.0000 1344.9000 526.2000 1349.7001 ;
	    RECT 527.4000 1345.5000 528.6000 1349.7001 ;
	    RECT 529.8000 1345.5000 531.0000 1349.7001 ;
	    RECT 532.2000 1345.5000 533.4000 1349.7001 ;
	    RECT 534.6000 1345.5000 535.8000 1349.7001 ;
	    RECT 537.0000 1346.7001 538.2000 1349.7001 ;
	    RECT 539.4000 1345.5000 540.6000 1349.7001 ;
	    RECT 541.8000 1346.7001 543.0000 1349.7001 ;
	    RECT 544.2000 1345.5000 545.4000 1349.7001 ;
	    RECT 546.6000 1345.5000 547.8000 1349.7001 ;
	    RECT 549.0000 1345.5000 550.2000 1349.7001 ;
	    RECT 522.6000 1343.7001 526.2000 1344.9000 ;
	    RECT 551.4000 1344.9000 552.6000 1349.7001 ;
	    RECT 522.6000 1342.8000 523.8000 1343.7001 ;
	    RECT 514.8000 1341.0000 516.6000 1341.9000 ;
	    RECT 521.1000 1341.9000 523.8000 1342.8000 ;
	    RECT 529.8000 1343.4000 531.3000 1344.6000 ;
	    RECT 535.8000 1343.4000 536.1000 1344.6000 ;
	    RECT 537.0000 1343.4000 538.2000 1344.6000 ;
	    RECT 539.4000 1343.7001 546.3000 1344.6000 ;
	    RECT 551.4000 1343.7001 555.3000 1344.9000 ;
	    RECT 556.2000 1343.7001 557.4000 1349.7001 ;
	    RECT 539.4000 1343.4000 540.6000 1343.7001 ;
	    RECT 514.8000 1338.0000 515.7000 1341.0000 ;
	    RECT 521.1000 1340.1000 522.3000 1341.9000 ;
	    RECT 516.6000 1338.9000 522.3000 1340.1000 ;
	    RECT 529.8000 1339.2001 531.0000 1343.4000 ;
	    RECT 541.8000 1342.5000 543.0000 1342.8000 ;
	    RECT 539.4000 1342.2001 540.6000 1342.5000 ;
	    RECT 534.0000 1341.3000 540.6000 1342.2001 ;
	    RECT 534.0000 1341.0000 535.2000 1341.3000 ;
	    RECT 541.8000 1340.4000 543.0000 1341.6000 ;
	    RECT 545.1000 1340.1000 546.3000 1343.7001 ;
	    RECT 554.1000 1342.8000 555.3000 1343.7001 ;
	    RECT 554.1000 1341.6000 558.6000 1342.8000 ;
	    RECT 561.0000 1340.7001 562.2000 1349.7001 ;
	    RECT 652.2000 1347.4501 653.4000 1347.6000 ;
	    RECT 659.4000 1347.4501 660.6000 1347.6000 ;
	    RECT 678.6000 1347.4501 679.8000 1347.6000 ;
	    RECT 652.2000 1346.5500 679.8000 1347.4501 ;
	    RECT 652.2000 1346.4000 653.4000 1346.5500 ;
	    RECT 659.4000 1346.4000 660.6000 1346.5500 ;
	    RECT 678.6000 1346.4000 679.8000 1346.5500 ;
	    RECT 534.6000 1338.9000 539.4000 1340.1000 ;
	    RECT 545.1000 1338.9000 548.1000 1340.1000 ;
	    RECT 549.0000 1339.5000 562.2000 1340.7001 ;
	    RECT 525.0000 1338.0000 526.2000 1338.9000 ;
	    RECT 514.8000 1337.1000 516.0000 1338.0000 ;
	    RECT 525.0000 1337.1000 550.5000 1338.0000 ;
	    RECT 551.4000 1337.4000 552.6000 1338.6000 ;
	    RECT 558.9000 1338.0000 560.1000 1338.3000 ;
	    RECT 553.5000 1337.1000 560.1000 1338.0000 ;
	    RECT 512.7000 1335.0000 514.2000 1336.2001 ;
	    RECT 513.0000 1333.5000 514.2000 1335.0000 ;
	    RECT 515.1000 1334.4000 516.0000 1337.1000 ;
	    RECT 516.9000 1336.2001 518.1000 1336.5000 ;
	    RECT 516.9000 1335.3000 555.3000 1336.2001 ;
	    RECT 551.1000 1335.0000 552.3000 1335.3000 ;
	    RECT 556.2000 1334.4000 557.4000 1335.6000 ;
	    RECT 515.1000 1333.5000 528.6000 1334.4000 ;
	    RECT 429.0000 1332.4501 430.2000 1332.6000 ;
	    RECT 457.8000 1332.4501 459.0000 1332.6000 ;
	    RECT 513.0000 1332.4501 514.2000 1332.6000 ;
	    RECT 429.0000 1331.5500 514.2000 1332.4501 ;
	    RECT 429.0000 1331.4000 430.2000 1331.5500 ;
	    RECT 457.8000 1331.4000 459.0000 1331.5500 ;
	    RECT 513.0000 1331.4000 514.2000 1331.5500 ;
	    RECT 374.4000 1330.2001 377.4000 1331.1000 ;
	    RECT 515.1000 1331.1000 516.0000 1333.5000 ;
	    RECT 527.4000 1333.2001 528.6000 1333.5000 ;
	    RECT 532.2000 1333.5000 545.1000 1334.4000 ;
	    RECT 532.2000 1333.2001 533.4000 1333.5000 ;
	    RECT 519.9000 1331.4000 523.8000 1332.6000 ;
	    RECT 361.8000 1323.3000 363.0000 1327.5000 ;
	    RECT 364.2000 1323.3000 365.4000 1327.5000 ;
	    RECT 366.6000 1323.3000 367.8000 1329.3000 ;
	    RECT 369.0000 1323.3000 370.2000 1330.2001 ;
	    RECT 374.4000 1329.3000 375.3000 1330.2001 ;
	    RECT 371.4000 1322.4000 372.6000 1329.3000 ;
	    RECT 373.8000 1328.4000 375.3000 1329.3000 ;
	    RECT 373.8000 1323.3000 375.0000 1328.4000 ;
	    RECT 376.2000 1323.3000 377.4000 1329.3000 ;
	    RECT 510.6000 1323.3000 511.8000 1329.3000 ;
	    RECT 513.0000 1323.3000 514.2000 1330.5000 ;
	    RECT 515.1000 1330.2001 519.0000 1331.1000 ;
	    RECT 515.4000 1323.3000 516.6000 1329.3000 ;
	    RECT 517.8000 1323.3000 519.0000 1330.2001 ;
	    RECT 520.2000 1323.3000 521.4000 1329.3000 ;
	    RECT 522.6000 1323.3000 523.8000 1331.4000 ;
	    RECT 524.7000 1330.2001 531.0000 1331.4000 ;
	    RECT 525.0000 1323.3000 526.2000 1329.3000 ;
	    RECT 527.4000 1323.3000 528.6000 1327.5000 ;
	    RECT 529.8000 1323.3000 531.0000 1327.5000 ;
	    RECT 532.2000 1323.3000 533.4000 1327.5000 ;
	    RECT 534.6000 1323.3000 535.8000 1332.6000 ;
	    RECT 539.4000 1331.4000 543.3000 1332.6000 ;
	    RECT 544.2000 1332.3000 545.1000 1333.5000 ;
	    RECT 546.6000 1334.1000 547.8000 1334.4000 ;
	    RECT 546.6000 1333.5000 554.7000 1334.1000 ;
	    RECT 546.6000 1333.2001 555.9000 1333.5000 ;
	    RECT 553.8000 1332.3000 555.9000 1333.2001 ;
	    RECT 544.2000 1331.4000 552.9000 1332.3000 ;
	    RECT 557.4000 1332.0000 559.8000 1333.2001 ;
	    RECT 557.4000 1331.4000 558.3000 1332.0000 ;
	    RECT 537.0000 1323.3000 538.2000 1329.3000 ;
	    RECT 539.4000 1323.3000 540.6000 1330.5000 ;
	    RECT 541.8000 1323.3000 543.0000 1329.3000 ;
	    RECT 544.2000 1323.3000 545.4000 1330.5000 ;
	    RECT 552.0000 1330.2001 558.3000 1331.4000 ;
	    RECT 561.0000 1331.1000 562.2000 1339.5000 ;
	    RECT 559.2000 1330.2001 562.2000 1331.1000 ;
	    RECT 695.4000 1340.7001 696.6000 1349.7001 ;
	    RECT 700.2000 1343.7001 701.4000 1349.7001 ;
	    RECT 705.0000 1344.9000 706.2000 1349.7001 ;
	    RECT 707.4000 1345.5000 708.6000 1349.7001 ;
	    RECT 709.8000 1345.5000 711.0000 1349.7001 ;
	    RECT 712.2000 1345.5000 713.4000 1349.7001 ;
	    RECT 714.6000 1346.7001 715.8000 1349.7001 ;
	    RECT 717.0000 1345.5000 718.2000 1349.7001 ;
	    RECT 719.4000 1346.7001 720.6000 1349.7001 ;
	    RECT 721.8000 1345.5000 723.0000 1349.7001 ;
	    RECT 724.2000 1345.5000 725.4000 1349.7001 ;
	    RECT 726.6000 1345.5000 727.8000 1349.7001 ;
	    RECT 729.0000 1345.5000 730.2000 1349.7001 ;
	    RECT 702.3000 1343.7001 706.2000 1344.9000 ;
	    RECT 731.4000 1344.9000 732.6000 1349.7001 ;
	    RECT 711.3000 1343.7001 718.2000 1344.6000 ;
	    RECT 702.3000 1342.8000 703.5000 1343.7001 ;
	    RECT 699.0000 1341.6000 703.5000 1342.8000 ;
	    RECT 695.4000 1339.5000 708.6000 1340.7001 ;
	    RECT 711.3000 1340.1000 712.5000 1343.7001 ;
	    RECT 717.0000 1343.4000 718.2000 1343.7001 ;
	    RECT 719.4000 1343.4000 720.6000 1344.6000 ;
	    RECT 721.5000 1343.4000 721.8000 1344.6000 ;
	    RECT 726.3000 1343.4000 727.8000 1344.6000 ;
	    RECT 731.4000 1343.7001 735.0000 1344.9000 ;
	    RECT 736.2000 1343.7001 737.4000 1349.7001 ;
	    RECT 714.6000 1342.5000 715.8000 1342.8000 ;
	    RECT 717.0000 1342.2001 718.2000 1342.5000 ;
	    RECT 714.6000 1340.4000 715.8000 1341.6000 ;
	    RECT 717.0000 1341.3000 723.6000 1342.2001 ;
	    RECT 722.4000 1341.0000 723.6000 1341.3000 ;
	    RECT 695.4000 1331.1000 696.6000 1339.5000 ;
	    RECT 709.5000 1338.9000 712.5000 1340.1000 ;
	    RECT 718.2000 1338.9000 723.0000 1340.1000 ;
	    RECT 726.6000 1339.2001 727.8000 1343.4000 ;
	    RECT 733.8000 1342.8000 735.0000 1343.7001 ;
	    RECT 733.8000 1341.9000 736.5000 1342.8000 ;
	    RECT 735.3000 1340.1000 736.5000 1341.9000 ;
	    RECT 741.0000 1341.9000 742.2000 1349.7001 ;
	    RECT 743.4000 1344.0000 744.6000 1349.7001 ;
	    RECT 745.8000 1346.7001 747.0000 1349.7001 ;
	    RECT 760.2000 1346.7001 761.4000 1349.7001 ;
	    RECT 760.2000 1345.5000 761.4000 1345.8000 ;
	    RECT 750.6000 1344.4501 751.8000 1344.6000 ;
	    RECT 760.2000 1344.4501 761.4000 1344.6000 ;
	    RECT 743.4000 1342.8000 744.9000 1344.0000 ;
	    RECT 750.6000 1343.5500 761.4000 1344.4501 ;
	    RECT 750.6000 1343.4000 751.8000 1343.5500 ;
	    RECT 760.2000 1343.4000 761.4000 1343.5500 ;
	    RECT 741.0000 1341.0000 742.8000 1341.9000 ;
	    RECT 735.3000 1338.9000 741.0000 1340.1000 ;
	    RECT 697.5000 1338.0000 698.7000 1338.3000 ;
	    RECT 697.5000 1337.1000 704.1000 1338.0000 ;
	    RECT 705.0000 1337.4000 706.2000 1338.6000 ;
	    RECT 731.4000 1338.0000 732.6000 1338.9000 ;
	    RECT 741.9000 1338.0000 742.8000 1341.0000 ;
	    RECT 707.1000 1337.1000 732.6000 1338.0000 ;
	    RECT 741.6000 1337.1000 742.8000 1338.0000 ;
	    RECT 739.5000 1336.2001 740.7000 1336.5000 ;
	    RECT 700.2000 1334.4000 701.4000 1335.6000 ;
	    RECT 702.3000 1335.3000 740.7000 1336.2001 ;
	    RECT 705.3000 1335.0000 706.5000 1335.3000 ;
	    RECT 741.6000 1334.4000 742.5000 1337.1000 ;
	    RECT 743.7000 1336.2001 744.9000 1342.8000 ;
	    RECT 762.6000 1342.5000 763.8000 1349.7001 ;
	    RECT 897.0000 1346.7001 898.2000 1349.7001 ;
	    RECT 839.4000 1344.4501 840.6000 1344.6000 ;
	    RECT 880.2000 1344.4501 881.4000 1344.6000 ;
	    RECT 839.4000 1343.5500 881.4000 1344.4501 ;
	    RECT 899.4000 1344.0000 900.6000 1349.7001 ;
	    RECT 839.4000 1343.4000 840.6000 1343.5500 ;
	    RECT 880.2000 1343.4000 881.4000 1343.5500 ;
	    RECT 899.1000 1342.8000 900.6000 1344.0000 ;
	    RECT 762.6000 1341.4501 763.8000 1341.6000 ;
	    RECT 817.8000 1341.4501 819.0000 1341.6000 ;
	    RECT 762.6000 1340.5500 819.0000 1341.4501 ;
	    RECT 762.6000 1340.4000 763.8000 1340.5500 ;
	    RECT 817.8000 1340.4000 819.0000 1340.5500 ;
	    RECT 709.8000 1334.1000 711.0000 1334.4000 ;
	    RECT 702.9000 1333.5000 711.0000 1334.1000 ;
	    RECT 701.7000 1333.2001 711.0000 1333.5000 ;
	    RECT 712.5000 1333.5000 725.4000 1334.4000 ;
	    RECT 697.8000 1332.0000 700.2000 1333.2001 ;
	    RECT 701.7000 1332.3000 703.8000 1333.2001 ;
	    RECT 712.5000 1332.3000 713.4000 1333.5000 ;
	    RECT 724.2000 1333.2001 725.4000 1333.5000 ;
	    RECT 729.0000 1333.5000 742.5000 1334.4000 ;
	    RECT 743.4000 1335.0000 744.9000 1336.2001 ;
	    RECT 743.4000 1333.5000 744.6000 1335.0000 ;
	    RECT 729.0000 1333.2001 730.2000 1333.5000 ;
	    RECT 699.3000 1331.4000 700.2000 1332.0000 ;
	    RECT 704.7000 1331.4000 713.4000 1332.3000 ;
	    RECT 714.3000 1331.4000 718.2000 1332.6000 ;
	    RECT 695.4000 1330.2001 698.4000 1331.1000 ;
	    RECT 699.3000 1330.2001 705.6000 1331.4000 ;
	    RECT 546.6000 1323.3000 547.8000 1327.5000 ;
	    RECT 549.0000 1323.3000 550.2000 1327.5000 ;
	    RECT 551.4000 1323.3000 552.6000 1329.3000 ;
	    RECT 553.8000 1323.3000 555.0000 1330.2001 ;
	    RECT 559.2000 1329.3000 560.1000 1330.2001 ;
	    RECT 697.5000 1329.3000 698.4000 1330.2001 ;
	    RECT 556.2000 1322.4000 557.4000 1329.3000 ;
	    RECT 558.6000 1328.4000 560.1000 1329.3000 ;
	    RECT 558.6000 1323.3000 559.8000 1328.4000 ;
	    RECT 561.0000 1323.3000 562.2000 1329.3000 ;
	    RECT 695.4000 1323.3000 696.6000 1329.3000 ;
	    RECT 697.5000 1328.4000 699.0000 1329.3000 ;
	    RECT 697.8000 1323.3000 699.0000 1328.4000 ;
	    RECT 700.2000 1322.4000 701.4000 1329.3000 ;
	    RECT 702.6000 1323.3000 703.8000 1330.2001 ;
	    RECT 705.0000 1323.3000 706.2000 1329.3000 ;
	    RECT 707.4000 1323.3000 708.6000 1327.5000 ;
	    RECT 709.8000 1323.3000 711.0000 1327.5000 ;
	    RECT 712.2000 1323.3000 713.4000 1330.5000 ;
	    RECT 714.6000 1323.3000 715.8000 1329.3000 ;
	    RECT 717.0000 1323.3000 718.2000 1330.5000 ;
	    RECT 719.4000 1323.3000 720.6000 1329.3000 ;
	    RECT 721.8000 1323.3000 723.0000 1332.6000 ;
	    RECT 733.8000 1331.4000 737.7000 1332.6000 ;
	    RECT 726.6000 1330.2001 732.9000 1331.4000 ;
	    RECT 724.2000 1323.3000 725.4000 1327.5000 ;
	    RECT 726.6000 1323.3000 727.8000 1327.5000 ;
	    RECT 729.0000 1323.3000 730.2000 1327.5000 ;
	    RECT 731.4000 1323.3000 732.6000 1329.3000 ;
	    RECT 733.8000 1323.3000 735.0000 1331.4000 ;
	    RECT 741.6000 1331.1000 742.5000 1333.5000 ;
	    RECT 743.4000 1331.4000 744.6000 1332.6000 ;
	    RECT 738.6000 1330.2001 742.5000 1331.1000 ;
	    RECT 736.2000 1323.3000 737.4000 1329.3000 ;
	    RECT 738.6000 1323.3000 739.8000 1330.2001 ;
	    RECT 741.0000 1323.3000 742.2000 1329.3000 ;
	    RECT 743.4000 1323.3000 744.6000 1330.5000 ;
	    RECT 745.8000 1323.3000 747.0000 1329.3000 ;
	    RECT 760.2000 1323.3000 761.4000 1329.3000 ;
	    RECT 762.6000 1323.3000 763.8000 1339.5000 ;
	    RECT 899.1000 1336.2001 900.3000 1342.8000 ;
	    RECT 901.8000 1341.9000 903.0000 1349.7001 ;
	    RECT 906.6000 1343.7001 907.8000 1349.7001 ;
	    RECT 911.4000 1344.9000 912.6000 1349.7001 ;
	    RECT 913.8000 1345.5000 915.0000 1349.7001 ;
	    RECT 916.2000 1345.5000 917.4000 1349.7001 ;
	    RECT 918.6000 1345.5000 919.8000 1349.7001 ;
	    RECT 921.0000 1345.5000 922.2000 1349.7001 ;
	    RECT 923.4000 1346.7001 924.6000 1349.7001 ;
	    RECT 925.8000 1345.5000 927.0000 1349.7001 ;
	    RECT 928.2000 1346.7001 929.4000 1349.7001 ;
	    RECT 930.6000 1345.5000 931.8000 1349.7001 ;
	    RECT 933.0000 1345.5000 934.2000 1349.7001 ;
	    RECT 935.4000 1345.5000 936.6000 1349.7001 ;
	    RECT 909.0000 1343.7001 912.6000 1344.9000 ;
	    RECT 937.8000 1344.9000 939.0000 1349.7001 ;
	    RECT 909.0000 1342.8000 910.2000 1343.7001 ;
	    RECT 901.2000 1341.0000 903.0000 1341.9000 ;
	    RECT 907.5000 1341.9000 910.2000 1342.8000 ;
	    RECT 916.2000 1343.4000 917.7000 1344.6000 ;
	    RECT 922.2000 1343.4000 922.5000 1344.6000 ;
	    RECT 923.4000 1343.4000 924.6000 1344.6000 ;
	    RECT 925.8000 1343.7001 932.7000 1344.6000 ;
	    RECT 937.8000 1343.7001 941.7000 1344.9000 ;
	    RECT 942.6000 1343.7001 943.8000 1349.7001 ;
	    RECT 925.8000 1343.4000 927.0000 1343.7001 ;
	    RECT 901.2000 1338.0000 902.1000 1341.0000 ;
	    RECT 907.5000 1340.1000 908.7000 1341.9000 ;
	    RECT 903.0000 1338.9000 908.7000 1340.1000 ;
	    RECT 916.2000 1339.2001 917.4000 1343.4000 ;
	    RECT 928.2000 1342.5000 929.4000 1342.8000 ;
	    RECT 925.8000 1342.2001 927.0000 1342.5000 ;
	    RECT 920.4000 1341.3000 927.0000 1342.2001 ;
	    RECT 920.4000 1341.0000 921.6000 1341.3000 ;
	    RECT 928.2000 1340.4000 929.4000 1341.6000 ;
	    RECT 931.5000 1340.1000 932.7000 1343.7001 ;
	    RECT 940.5000 1342.8000 941.7000 1343.7001 ;
	    RECT 940.5000 1341.6000 945.0000 1342.8000 ;
	    RECT 947.4000 1340.7001 948.6000 1349.7001 ;
	    RECT 971.4000 1343.7001 972.6000 1349.7001 ;
	    RECT 973.8000 1344.0000 975.0000 1349.7001 ;
	    RECT 976.2000 1344.9000 977.4000 1349.7001 ;
	    RECT 978.6000 1344.0000 979.8000 1349.7001 ;
	    RECT 993.0000 1346.7001 994.2000 1349.7001 ;
	    RECT 993.0000 1345.5000 994.2000 1345.8000 ;
	    RECT 973.8000 1343.7001 979.8000 1344.0000 ;
	    RECT 983.4000 1344.4501 984.6000 1344.6000 ;
	    RECT 993.0000 1344.4501 994.2000 1344.6000 ;
	    RECT 971.7000 1342.5000 972.6000 1343.7001 ;
	    RECT 974.1000 1343.1000 979.5000 1343.7001 ;
	    RECT 983.4000 1343.5500 994.2000 1344.4501 ;
	    RECT 983.4000 1343.4000 984.6000 1343.5500 ;
	    RECT 993.0000 1343.4000 994.2000 1343.5500 ;
	    RECT 995.4000 1342.5000 996.6000 1349.7001 ;
	    RECT 1019.4000 1344.0000 1020.6000 1349.7001 ;
	    RECT 1021.8000 1344.9000 1023.0000 1349.7001 ;
	    RECT 1024.2001 1344.0000 1025.4000 1349.7001 ;
	    RECT 1019.4000 1343.7001 1025.4000 1344.0000 ;
	    RECT 1026.6000 1343.7001 1027.8000 1349.7001 ;
	    RECT 1031.4000 1344.4501 1032.6000 1344.6000 ;
	    RECT 1019.7000 1343.1000 1025.1000 1343.7001 ;
	    RECT 1026.6000 1342.5000 1027.5000 1343.7001 ;
	    RECT 1031.4000 1343.5500 1044.4501 1344.4501 ;
	    RECT 1045.8000 1343.7001 1047.0000 1349.7001 ;
	    RECT 1049.7001 1344.6000 1050.9000 1349.7001 ;
	    RECT 1182.6000 1346.7001 1183.8000 1349.7001 ;
	    RECT 1048.2001 1343.7001 1050.9000 1344.6000 ;
	    RECT 1185.0000 1344.0000 1186.2001 1349.7001 ;
	    RECT 1031.4000 1343.4000 1032.6000 1343.5500 ;
	    RECT 921.0000 1338.9000 925.8000 1340.1000 ;
	    RECT 931.5000 1338.9000 934.5000 1340.1000 ;
	    RECT 935.4000 1339.5000 948.6000 1340.7001 ;
	    RECT 949.8000 1341.4501 951.0000 1341.6000 ;
	    RECT 971.4000 1341.4501 972.6000 1341.6000 ;
	    RECT 949.8000 1340.5500 972.6000 1341.4501 ;
	    RECT 949.8000 1340.4000 951.0000 1340.5500 ;
	    RECT 971.4000 1340.4000 972.6000 1340.5500 ;
	    RECT 973.5000 1340.4000 975.3000 1341.6000 ;
	    RECT 977.4000 1340.7001 977.7000 1342.2001 ;
	    RECT 978.6000 1340.4000 979.8000 1341.6000 ;
	    RECT 995.4000 1341.4501 996.6000 1341.6000 ;
	    RECT 981.1500 1340.5500 996.6000 1341.4501 ;
	    RECT 911.4000 1338.0000 912.6000 1338.9000 ;
	    RECT 901.2000 1337.1000 902.4000 1338.0000 ;
	    RECT 911.4000 1337.1000 936.9000 1338.0000 ;
	    RECT 937.8000 1337.4000 939.0000 1338.6000 ;
	    RECT 945.3000 1338.0000 946.5000 1338.3000 ;
	    RECT 939.9000 1337.1000 946.5000 1338.0000 ;
	    RECT 899.1000 1335.0000 900.6000 1336.2001 ;
	    RECT 899.4000 1333.5000 900.6000 1335.0000 ;
	    RECT 901.5000 1334.4000 902.4000 1337.1000 ;
	    RECT 903.3000 1336.2001 904.5000 1336.5000 ;
	    RECT 903.3000 1335.3000 941.7000 1336.2001 ;
	    RECT 942.6000 1335.4501 943.8000 1335.6000 ;
	    RECT 945.0000 1335.4501 946.2000 1335.6000 ;
	    RECT 937.5000 1335.0000 938.7000 1335.3000 ;
	    RECT 942.6000 1334.5500 946.2000 1335.4501 ;
	    RECT 942.6000 1334.4000 943.8000 1334.5500 ;
	    RECT 945.0000 1334.4000 946.2000 1334.5500 ;
	    RECT 901.5000 1333.5000 915.0000 1334.4000 ;
	    RECT 899.4000 1331.4000 900.6000 1332.6000 ;
	    RECT 901.5000 1331.1000 902.4000 1333.5000 ;
	    RECT 913.8000 1333.2001 915.0000 1333.5000 ;
	    RECT 918.6000 1333.5000 931.5000 1334.4000 ;
	    RECT 918.6000 1333.2001 919.8000 1333.5000 ;
	    RECT 906.3000 1331.4000 910.2000 1332.6000 ;
	    RECT 897.0000 1323.3000 898.2000 1329.3000 ;
	    RECT 899.4000 1323.3000 900.6000 1330.5000 ;
	    RECT 901.5000 1330.2001 905.4000 1331.1000 ;
	    RECT 901.8000 1323.3000 903.0000 1329.3000 ;
	    RECT 904.2000 1323.3000 905.4000 1330.2001 ;
	    RECT 906.6000 1323.3000 907.8000 1329.3000 ;
	    RECT 909.0000 1323.3000 910.2000 1331.4000 ;
	    RECT 911.1000 1330.2001 917.4000 1331.4000 ;
	    RECT 911.4000 1323.3000 912.6000 1329.3000 ;
	    RECT 913.8000 1323.3000 915.0000 1327.5000 ;
	    RECT 916.2000 1323.3000 917.4000 1327.5000 ;
	    RECT 918.6000 1323.3000 919.8000 1327.5000 ;
	    RECT 921.0000 1323.3000 922.2000 1332.6000 ;
	    RECT 925.8000 1331.4000 929.7000 1332.6000 ;
	    RECT 930.6000 1332.3000 931.5000 1333.5000 ;
	    RECT 933.0000 1334.1000 934.2000 1334.4000 ;
	    RECT 933.0000 1333.5000 941.1000 1334.1000 ;
	    RECT 933.0000 1333.2001 942.3000 1333.5000 ;
	    RECT 940.2000 1332.3000 942.3000 1333.2001 ;
	    RECT 930.6000 1331.4000 939.3000 1332.3000 ;
	    RECT 943.8000 1332.0000 946.2000 1333.2001 ;
	    RECT 943.8000 1331.4000 944.7000 1332.0000 ;
	    RECT 923.4000 1323.3000 924.6000 1329.3000 ;
	    RECT 925.8000 1323.3000 927.0000 1330.5000 ;
	    RECT 928.2000 1323.3000 929.4000 1329.3000 ;
	    RECT 930.6000 1323.3000 931.8000 1330.5000 ;
	    RECT 938.4000 1330.2001 944.7000 1331.4000 ;
	    RECT 947.4000 1331.1000 948.6000 1339.5000 ;
	    RECT 971.4000 1334.4000 972.6000 1335.6000 ;
	    RECT 974.4000 1335.3000 975.3000 1340.4000 ;
	    RECT 976.2000 1339.5000 977.4000 1339.8000 ;
	    RECT 976.2000 1338.4501 977.4000 1338.6000 ;
	    RECT 981.1500 1338.4501 982.0500 1340.5500 ;
	    RECT 995.4000 1340.4000 996.6000 1340.5500 ;
	    RECT 1019.4000 1340.4000 1020.6000 1341.6000 ;
	    RECT 1021.5000 1340.7001 1021.8000 1342.2001 ;
	    RECT 1023.9000 1340.4000 1025.7001 1341.6000 ;
	    RECT 1026.6000 1341.4501 1027.8000 1341.6000 ;
	    RECT 1041.0000 1341.4501 1042.2001 1341.6000 ;
	    RECT 1026.6000 1340.5500 1042.2001 1341.4501 ;
	    RECT 1043.5500 1341.4501 1044.4501 1343.5500 ;
	    RECT 1045.8000 1342.5000 1047.0000 1342.8000 ;
	    RECT 1045.8000 1341.4501 1047.0000 1341.6000 ;
	    RECT 1043.5500 1340.5500 1047.0000 1341.4501 ;
	    RECT 1026.6000 1340.4000 1027.8000 1340.5500 ;
	    RECT 1041.0000 1340.4000 1042.2001 1340.5500 ;
	    RECT 1045.8000 1340.4000 1047.0000 1340.5500 ;
	    RECT 1021.8000 1339.5000 1023.0000 1339.8000 ;
	    RECT 976.2000 1337.5500 982.0500 1338.4501 ;
	    RECT 976.2000 1337.4000 977.4000 1337.5500 ;
	    RECT 974.4000 1334.4000 975.9000 1335.3000 ;
	    RECT 972.6000 1332.6000 973.5000 1333.5000 ;
	    RECT 972.6000 1331.4000 973.8000 1332.6000 ;
	    RECT 945.6000 1330.2001 948.6000 1331.1000 ;
	    RECT 933.0000 1323.3000 934.2000 1327.5000 ;
	    RECT 935.4000 1323.3000 936.6000 1327.5000 ;
	    RECT 937.8000 1323.3000 939.0000 1329.3000 ;
	    RECT 940.2000 1323.3000 941.4000 1330.2001 ;
	    RECT 945.6000 1329.3000 946.5000 1330.2001 ;
	    RECT 942.6000 1322.4000 943.8000 1329.3000 ;
	    RECT 945.0000 1328.4000 946.5000 1329.3000 ;
	    RECT 945.0000 1323.3000 946.2000 1328.4000 ;
	    RECT 947.4000 1323.3000 948.6000 1329.3000 ;
	    RECT 972.3000 1323.3000 973.5000 1329.3000 ;
	    RECT 974.7000 1323.3000 975.9000 1334.4000 ;
	    RECT 978.6000 1323.3000 979.8000 1335.3000 ;
	    RECT 993.0000 1323.3000 994.2000 1329.3000 ;
	    RECT 995.4000 1323.3000 996.6000 1339.5000 ;
	    RECT 1021.8000 1337.4000 1023.0000 1338.6000 ;
	    RECT 1023.9000 1335.3000 1024.8000 1340.4000 ;
	    RECT 1048.2001 1339.5000 1049.4000 1343.7001 ;
	    RECT 1184.7001 1342.8000 1186.2001 1344.0000 ;
	    RECT 1048.2001 1338.4501 1049.4000 1338.6000 ;
	    RECT 1026.7500 1337.5500 1049.4000 1338.4501 ;
	    RECT 1026.7500 1335.6000 1027.6500 1337.5500 ;
	    RECT 1048.2001 1337.4000 1049.4000 1337.5500 ;
	    RECT 1019.4000 1323.3000 1020.6000 1335.3000 ;
	    RECT 1023.3000 1334.4000 1024.8000 1335.3000 ;
	    RECT 1026.6000 1334.4000 1027.8000 1335.6000 ;
	    RECT 1023.3000 1323.3000 1024.5000 1334.4000 ;
	    RECT 1025.7001 1332.6000 1026.6000 1333.5000 ;
	    RECT 1025.4000 1331.4000 1026.6000 1332.6000 ;
	    RECT 1025.7001 1323.3000 1026.9000 1329.3000 ;
	    RECT 1045.8000 1323.3000 1047.0000 1329.3000 ;
	    RECT 1048.2001 1323.3000 1049.4000 1336.5000 ;
	    RECT 1184.7001 1336.2001 1185.9000 1342.8000 ;
	    RECT 1187.4000 1341.9000 1188.6000 1349.7001 ;
	    RECT 1192.2001 1343.7001 1193.4000 1349.7001 ;
	    RECT 1197.0000 1344.9000 1198.2001 1349.7001 ;
	    RECT 1199.4000 1345.5000 1200.6000 1349.7001 ;
	    RECT 1201.8000 1345.5000 1203.0000 1349.7001 ;
	    RECT 1204.2001 1345.5000 1205.4000 1349.7001 ;
	    RECT 1206.6000 1345.5000 1207.8000 1349.7001 ;
	    RECT 1209.0000 1346.7001 1210.2001 1349.7001 ;
	    RECT 1211.4000 1345.5000 1212.6000 1349.7001 ;
	    RECT 1213.8000 1346.7001 1215.0000 1349.7001 ;
	    RECT 1216.2001 1345.5000 1217.4000 1349.7001 ;
	    RECT 1218.6000 1345.5000 1219.8000 1349.7001 ;
	    RECT 1221.0000 1345.5000 1222.2001 1349.7001 ;
	    RECT 1194.6000 1343.7001 1198.2001 1344.9000 ;
	    RECT 1223.4000 1344.9000 1224.6000 1349.7001 ;
	    RECT 1194.6000 1342.8000 1195.8000 1343.7001 ;
	    RECT 1186.8000 1341.0000 1188.6000 1341.9000 ;
	    RECT 1193.1000 1341.9000 1195.8000 1342.8000 ;
	    RECT 1201.8000 1343.4000 1203.3000 1344.6000 ;
	    RECT 1207.8000 1343.4000 1208.1000 1344.6000 ;
	    RECT 1209.0000 1343.4000 1210.2001 1344.6000 ;
	    RECT 1211.4000 1343.7001 1218.3000 1344.6000 ;
	    RECT 1223.4000 1343.7001 1227.3000 1344.9000 ;
	    RECT 1228.2001 1343.7001 1229.4000 1349.7001 ;
	    RECT 1211.4000 1343.4000 1212.6000 1343.7001 ;
	    RECT 1186.8000 1338.0000 1187.7001 1341.0000 ;
	    RECT 1193.1000 1340.1000 1194.3000 1341.9000 ;
	    RECT 1188.6000 1338.9000 1194.3000 1340.1000 ;
	    RECT 1201.8000 1339.2001 1203.0000 1343.4000 ;
	    RECT 1213.8000 1342.5000 1215.0000 1342.8000 ;
	    RECT 1211.4000 1342.2001 1212.6000 1342.5000 ;
	    RECT 1206.0000 1341.3000 1212.6000 1342.2001 ;
	    RECT 1206.0000 1341.0000 1207.2001 1341.3000 ;
	    RECT 1213.8000 1340.4000 1215.0000 1341.6000 ;
	    RECT 1217.1000 1340.1000 1218.3000 1343.7001 ;
	    RECT 1226.1000 1342.8000 1227.3000 1343.7001 ;
	    RECT 1226.1000 1341.6000 1230.6000 1342.8000 ;
	    RECT 1233.0000 1340.7001 1234.2001 1349.7001 ;
	    RECT 1247.4000 1346.7001 1248.6000 1349.7001 ;
	    RECT 1247.4000 1345.5000 1248.6000 1345.8000 ;
	    RECT 1235.4000 1344.4501 1236.6000 1344.6000 ;
	    RECT 1247.4000 1344.4501 1248.6000 1344.6000 ;
	    RECT 1235.4000 1343.5500 1248.6000 1344.4501 ;
	    RECT 1235.4000 1343.4000 1236.6000 1343.5500 ;
	    RECT 1247.4000 1343.4000 1248.6000 1343.5500 ;
	    RECT 1249.8000 1342.5000 1251.0000 1349.7001 ;
	    RECT 1273.8000 1344.0000 1275.0000 1349.7001 ;
	    RECT 1276.2001 1344.9000 1277.4000 1349.7001 ;
	    RECT 1278.6000 1344.0000 1279.8000 1349.7001 ;
	    RECT 1273.8000 1343.7001 1279.8000 1344.0000 ;
	    RECT 1281.0000 1343.7001 1282.2001 1349.7001 ;
	    RECT 1274.1000 1343.1000 1279.5000 1343.7001 ;
	    RECT 1281.0000 1342.5000 1281.9000 1343.7001 ;
	    RECT 1293.0000 1342.5000 1294.2001 1349.7001 ;
	    RECT 1295.4000 1346.7001 1296.6000 1349.7001 ;
	    RECT 1309.8000 1346.7001 1311.0000 1349.7001 ;
	    RECT 1295.4000 1345.5000 1296.6000 1345.8000 ;
	    RECT 1309.8000 1345.5000 1311.0000 1345.8000 ;
	    RECT 1295.4000 1343.4000 1296.6000 1344.6000 ;
	    RECT 1300.2001 1344.4501 1301.4000 1344.6000 ;
	    RECT 1309.8000 1344.4501 1311.0000 1344.6000 ;
	    RECT 1300.2001 1343.5500 1311.0000 1344.4501 ;
	    RECT 1300.2001 1343.4000 1301.4000 1343.5500 ;
	    RECT 1309.8000 1343.4000 1311.0000 1343.5500 ;
	    RECT 1312.2001 1342.5000 1313.4000 1349.7001 ;
	    RECT 1336.2001 1344.0000 1337.4000 1349.7001 ;
	    RECT 1338.6000 1344.9000 1339.8000 1349.7001 ;
	    RECT 1341.0000 1344.0000 1342.2001 1349.7001 ;
	    RECT 1336.2001 1343.7001 1342.2001 1344.0000 ;
	    RECT 1343.4000 1343.7001 1344.6000 1349.7001 ;
	    RECT 1370.7001 1344.6000 1371.9000 1349.7001 ;
	    RECT 1370.7001 1343.7001 1373.4000 1344.6000 ;
	    RECT 1374.6000 1343.7001 1375.8000 1349.7001 ;
	    RECT 1394.7001 1344.6000 1395.9000 1349.7001 ;
	    RECT 1394.7001 1343.7001 1397.4000 1344.6000 ;
	    RECT 1398.6000 1343.7001 1399.8000 1349.7001 ;
	    RECT 1417.8000 1343.7001 1419.0000 1349.7001 ;
	    RECT 1421.7001 1344.6000 1422.9000 1349.7001 ;
	    RECT 1420.2001 1343.7001 1422.9000 1344.6000 ;
	    RECT 1446.6000 1343.7001 1447.8000 1349.7001 ;
	    RECT 1449.0000 1344.0000 1450.2001 1349.7001 ;
	    RECT 1451.4000 1344.9000 1452.6000 1349.7001 ;
	    RECT 1453.8000 1344.0000 1455.0000 1349.7001 ;
	    RECT 1449.0000 1343.7001 1455.0000 1344.0000 ;
	    RECT 1477.8000 1343.7001 1479.0000 1349.7001 ;
	    RECT 1480.2001 1344.0000 1481.4000 1349.7001 ;
	    RECT 1482.6000 1344.9000 1483.8000 1349.7001 ;
	    RECT 1485.0000 1344.0000 1486.2001 1349.7001 ;
	    RECT 1480.2001 1343.7001 1486.2001 1344.0000 ;
	    RECT 1336.5000 1343.1000 1341.9000 1343.7001 ;
	    RECT 1343.4000 1342.5000 1344.3000 1343.7001 ;
	    RECT 1206.6000 1338.9000 1211.4000 1340.1000 ;
	    RECT 1217.1000 1338.9000 1220.1000 1340.1000 ;
	    RECT 1221.0000 1339.5000 1234.2001 1340.7001 ;
	    RECT 1249.8000 1341.4501 1251.0000 1341.6000 ;
	    RECT 1249.8000 1340.5500 1272.4501 1341.4501 ;
	    RECT 1249.8000 1340.4000 1251.0000 1340.5500 ;
	    RECT 1197.0000 1338.0000 1198.2001 1338.9000 ;
	    RECT 1186.8000 1337.1000 1188.0000 1338.0000 ;
	    RECT 1197.0000 1337.1000 1222.5000 1338.0000 ;
	    RECT 1223.4000 1337.4000 1224.6000 1338.6000 ;
	    RECT 1230.9000 1338.0000 1232.1000 1338.3000 ;
	    RECT 1225.5000 1337.1000 1232.1000 1338.0000 ;
	    RECT 1050.6000 1335.4501 1051.8000 1335.6000 ;
	    RECT 1074.6000 1335.4501 1075.8000 1335.6000 ;
	    RECT 1050.6000 1334.5500 1075.8000 1335.4501 ;
	    RECT 1184.7001 1335.0000 1186.2001 1336.2001 ;
	    RECT 1050.6000 1334.4000 1051.8000 1334.5500 ;
	    RECT 1074.6000 1334.4000 1075.8000 1334.5500 ;
	    RECT 1185.0000 1333.5000 1186.2001 1335.0000 ;
	    RECT 1187.1000 1334.4000 1188.0000 1337.1000 ;
	    RECT 1188.9000 1336.2001 1190.1000 1336.5000 ;
	    RECT 1188.9000 1335.3000 1227.3000 1336.2001 ;
	    RECT 1223.1000 1335.0000 1224.3000 1335.3000 ;
	    RECT 1228.2001 1334.4000 1229.4000 1335.6000 ;
	    RECT 1187.1000 1333.5000 1200.6000 1334.4000 ;
	    RECT 1050.6000 1333.2001 1051.8000 1333.5000 ;
	    RECT 1125.0000 1332.4501 1126.2001 1332.6000 ;
	    RECT 1185.0000 1332.4501 1186.2001 1332.6000 ;
	    RECT 1125.0000 1331.5500 1186.2001 1332.4501 ;
	    RECT 1125.0000 1331.4000 1126.2001 1331.5500 ;
	    RECT 1185.0000 1331.4000 1186.2001 1331.5500 ;
	    RECT 1187.1000 1331.1000 1188.0000 1333.5000 ;
	    RECT 1199.4000 1333.2001 1200.6000 1333.5000 ;
	    RECT 1204.2001 1333.5000 1217.1000 1334.4000 ;
	    RECT 1204.2001 1333.2001 1205.4000 1333.5000 ;
	    RECT 1191.9000 1331.4000 1195.8000 1332.6000 ;
	    RECT 1050.6000 1323.3000 1051.8000 1329.3000 ;
	    RECT 1182.6000 1323.3000 1183.8000 1329.3000 ;
	    RECT 1185.0000 1323.3000 1186.2001 1330.5000 ;
	    RECT 1187.1000 1330.2001 1191.0000 1331.1000 ;
	    RECT 1187.4000 1323.3000 1188.6000 1329.3000 ;
	    RECT 1189.8000 1323.3000 1191.0000 1330.2001 ;
	    RECT 1192.2001 1323.3000 1193.4000 1329.3000 ;
	    RECT 1194.6000 1323.3000 1195.8000 1331.4000 ;
	    RECT 1196.7001 1330.2001 1203.0000 1331.4000 ;
	    RECT 1197.0000 1323.3000 1198.2001 1329.3000 ;
	    RECT 1199.4000 1323.3000 1200.6000 1327.5000 ;
	    RECT 1201.8000 1323.3000 1203.0000 1327.5000 ;
	    RECT 1204.2001 1323.3000 1205.4000 1327.5000 ;
	    RECT 1206.6000 1323.3000 1207.8000 1332.6000 ;
	    RECT 1211.4000 1331.4000 1215.3000 1332.6000 ;
	    RECT 1216.2001 1332.3000 1217.1000 1333.5000 ;
	    RECT 1218.6000 1334.1000 1219.8000 1334.4000 ;
	    RECT 1218.6000 1333.5000 1226.7001 1334.1000 ;
	    RECT 1218.6000 1333.2001 1227.9000 1333.5000 ;
	    RECT 1225.8000 1332.3000 1227.9000 1333.2001 ;
	    RECT 1216.2001 1331.4000 1224.9000 1332.3000 ;
	    RECT 1229.4000 1332.0000 1231.8000 1333.2001 ;
	    RECT 1229.4000 1331.4000 1230.3000 1332.0000 ;
	    RECT 1209.0000 1323.3000 1210.2001 1329.3000 ;
	    RECT 1211.4000 1323.3000 1212.6000 1330.5000 ;
	    RECT 1213.8000 1323.3000 1215.0000 1329.3000 ;
	    RECT 1216.2001 1323.3000 1217.4000 1330.5000 ;
	    RECT 1224.0000 1330.2001 1230.3000 1331.4000 ;
	    RECT 1233.0000 1331.1000 1234.2001 1339.5000 ;
	    RECT 1231.2001 1330.2001 1234.2001 1331.1000 ;
	    RECT 1218.6000 1323.3000 1219.8000 1327.5000 ;
	    RECT 1221.0000 1323.3000 1222.2001 1327.5000 ;
	    RECT 1223.4000 1323.3000 1224.6000 1329.3000 ;
	    RECT 1225.8000 1323.3000 1227.0000 1330.2001 ;
	    RECT 1231.2001 1329.3000 1232.1000 1330.2001 ;
	    RECT 1228.2001 1322.4000 1229.4000 1329.3000 ;
	    RECT 1230.6000 1328.4000 1232.1000 1329.3000 ;
	    RECT 1230.6000 1323.3000 1231.8000 1328.4000 ;
	    RECT 1233.0000 1323.3000 1234.2001 1329.3000 ;
	    RECT 1247.4000 1323.3000 1248.6000 1329.3000 ;
	    RECT 1249.8000 1323.3000 1251.0000 1339.5000 ;
	    RECT 1271.5500 1338.4501 1272.4501 1340.5500 ;
	    RECT 1273.8000 1340.4000 1275.0000 1341.6000 ;
	    RECT 1275.9000 1340.7001 1276.2001 1342.2001 ;
	    RECT 1278.3000 1340.4000 1280.1000 1341.6000 ;
	    RECT 1281.0000 1340.4000 1282.2001 1341.6000 ;
	    RECT 1293.0000 1341.4501 1294.2001 1341.6000 ;
	    RECT 1309.8000 1341.4501 1311.0000 1341.6000 ;
	    RECT 1293.0000 1340.5500 1311.0000 1341.4501 ;
	    RECT 1293.0000 1340.4000 1294.2001 1340.5500 ;
	    RECT 1309.8000 1340.4000 1311.0000 1340.5500 ;
	    RECT 1312.2001 1341.4501 1313.4000 1341.6000 ;
	    RECT 1312.2001 1340.5500 1327.6500 1341.4501 ;
	    RECT 1312.2001 1340.4000 1313.4000 1340.5500 ;
	    RECT 1276.2001 1339.5000 1277.4000 1339.8000 ;
	    RECT 1276.2001 1338.4501 1277.4000 1338.6000 ;
	    RECT 1271.5500 1337.5500 1277.4000 1338.4501 ;
	    RECT 1276.2001 1337.4000 1277.4000 1337.5500 ;
	    RECT 1278.3000 1335.3000 1279.2001 1340.4000 ;
	    RECT 1273.8000 1323.3000 1275.0000 1335.3000 ;
	    RECT 1277.7001 1334.4000 1279.2001 1335.3000 ;
	    RECT 1281.0000 1335.4501 1282.2001 1335.6000 ;
	    RECT 1283.4000 1335.4501 1284.6000 1335.6000 ;
	    RECT 1281.0000 1334.5500 1284.6000 1335.4501 ;
	    RECT 1281.0000 1334.4000 1282.2001 1334.5500 ;
	    RECT 1283.4000 1334.4000 1284.6000 1334.5500 ;
	    RECT 1277.7001 1323.3000 1278.9000 1334.4000 ;
	    RECT 1280.1000 1332.6000 1281.0000 1333.5000 ;
	    RECT 1279.8000 1331.4000 1281.0000 1332.6000 ;
	    RECT 1280.1000 1323.3000 1281.3000 1329.3000 ;
	    RECT 1293.0000 1323.3000 1294.2001 1339.5000 ;
	    RECT 1295.4000 1323.3000 1296.6000 1329.3000 ;
	    RECT 1309.8000 1323.3000 1311.0000 1329.3000 ;
	    RECT 1312.2001 1323.3000 1313.4000 1339.5000 ;
	    RECT 1326.7500 1338.4501 1327.6500 1340.5500 ;
	    RECT 1336.2001 1340.4000 1337.4000 1341.6000 ;
	    RECT 1338.3000 1340.7001 1338.6000 1342.2001 ;
	    RECT 1340.7001 1340.4000 1342.5000 1341.6000 ;
	    RECT 1343.4000 1340.4000 1344.6000 1341.6000 ;
	    RECT 1338.6000 1339.5000 1339.8000 1339.8000 ;
	    RECT 1338.6000 1338.4501 1339.8000 1338.6000 ;
	    RECT 1326.7500 1337.5500 1339.8000 1338.4501 ;
	    RECT 1338.6000 1337.4000 1339.8000 1337.5500 ;
	    RECT 1340.7001 1335.3000 1341.6000 1340.4000 ;
	    RECT 1372.2001 1339.5000 1373.4000 1343.7001 ;
	    RECT 1374.6000 1342.5000 1375.8000 1342.8000 ;
	    RECT 1374.6000 1341.4501 1375.8000 1341.6000 ;
	    RECT 1377.0000 1341.4501 1378.2001 1341.6000 ;
	    RECT 1374.6000 1340.5500 1378.2001 1341.4501 ;
	    RECT 1374.6000 1340.4000 1375.8000 1340.5500 ;
	    RECT 1377.0000 1340.4000 1378.2001 1340.5500 ;
	    RECT 1396.2001 1339.5000 1397.4000 1343.7001 ;
	    RECT 1398.6000 1342.5000 1399.8000 1342.8000 ;
	    RECT 1417.8000 1342.5000 1419.0000 1342.8000 ;
	    RECT 1398.6000 1341.4501 1399.8000 1341.6000 ;
	    RECT 1408.2001 1341.4501 1409.4000 1341.6000 ;
	    RECT 1398.6000 1340.5500 1409.4000 1341.4501 ;
	    RECT 1398.6000 1340.4000 1399.8000 1340.5500 ;
	    RECT 1408.2001 1340.4000 1409.4000 1340.5500 ;
	    RECT 1417.8000 1340.4000 1419.0000 1341.6000 ;
	    RECT 1420.2001 1339.5000 1421.4000 1343.7001 ;
	    RECT 1446.9000 1342.5000 1447.8000 1343.7001 ;
	    RECT 1449.3000 1343.1000 1454.7001 1343.7001 ;
	    RECT 1478.1000 1342.5000 1479.0000 1343.7001 ;
	    RECT 1480.5000 1343.1000 1485.9000 1343.7001 ;
	    RECT 1499.4000 1342.5000 1500.6000 1349.7001 ;
	    RECT 1501.8000 1346.7001 1503.0000 1349.7001 ;
	    RECT 1516.2001 1346.7001 1517.4000 1349.7001 ;
	    RECT 1501.8000 1345.5000 1503.0000 1345.8000 ;
	    RECT 1516.2001 1345.5000 1517.4000 1345.8000 ;
	    RECT 1501.8000 1344.4501 1503.0000 1344.6000 ;
	    RECT 1513.8000 1344.4501 1515.0000 1344.6000 ;
	    RECT 1501.8000 1343.5500 1515.0000 1344.4501 ;
	    RECT 1501.8000 1343.4000 1503.0000 1343.5500 ;
	    RECT 1513.8000 1343.4000 1515.0000 1343.5500 ;
	    RECT 1516.2001 1343.4000 1517.4000 1344.6000 ;
	    RECT 1518.6000 1342.5000 1519.8000 1349.7001 ;
	    RECT 1542.6000 1343.7001 1543.8000 1349.7001 ;
	    RECT 1545.0000 1344.0000 1546.2001 1349.7001 ;
	    RECT 1547.4000 1344.9000 1548.6000 1349.7001 ;
	    RECT 1549.8000 1344.0000 1551.0000 1349.7001 ;
	    RECT 1545.0000 1343.7001 1551.0000 1344.0000 ;
	    RECT 1542.9000 1342.5000 1543.8000 1343.7001 ;
	    RECT 1545.3000 1343.1000 1550.7001 1343.7001 ;
	    RECT 1446.6000 1340.4000 1447.8000 1341.6000 ;
	    RECT 1448.7001 1340.4000 1450.5000 1341.6000 ;
	    RECT 1452.6000 1340.7001 1452.9000 1342.2001 ;
	    RECT 1453.8000 1340.4000 1455.0000 1341.6000 ;
	    RECT 1477.8000 1340.4000 1479.0000 1341.6000 ;
	    RECT 1479.9000 1340.4000 1481.7001 1341.6000 ;
	    RECT 1483.8000 1340.7001 1484.1000 1342.2001 ;
	    RECT 1485.0000 1340.4000 1486.2001 1341.6000 ;
	    RECT 1499.4000 1341.4501 1500.6000 1341.6000 ;
	    RECT 1487.5500 1340.5500 1500.6000 1341.4501 ;
	    RECT 1348.2001 1338.4501 1349.4000 1338.6000 ;
	    RECT 1343.5500 1337.5500 1349.4000 1338.4501 ;
	    RECT 1343.5500 1335.6000 1344.4501 1337.5500 ;
	    RECT 1348.2001 1337.4000 1349.4000 1337.5500 ;
	    RECT 1350.6000 1338.4501 1351.8000 1338.6000 ;
	    RECT 1372.2001 1338.4501 1373.4000 1338.6000 ;
	    RECT 1350.6000 1337.5500 1373.4000 1338.4501 ;
	    RECT 1350.6000 1337.4000 1351.8000 1337.5500 ;
	    RECT 1372.2001 1337.4000 1373.4000 1337.5500 ;
	    RECT 1384.2001 1338.4501 1385.4000 1338.6000 ;
	    RECT 1396.2001 1338.4501 1397.4000 1338.6000 ;
	    RECT 1384.2001 1337.5500 1397.4000 1338.4501 ;
	    RECT 1384.2001 1337.4000 1385.4000 1337.5500 ;
	    RECT 1396.2001 1337.4000 1397.4000 1337.5500 ;
	    RECT 1398.6000 1338.4501 1399.8000 1338.6000 ;
	    RECT 1420.2001 1338.4501 1421.4000 1338.6000 ;
	    RECT 1398.6000 1337.5500 1421.4000 1338.4501 ;
	    RECT 1398.6000 1337.4000 1399.8000 1337.5500 ;
	    RECT 1420.2001 1337.4000 1421.4000 1337.5500 ;
	    RECT 1336.2001 1323.3000 1337.4000 1335.3000 ;
	    RECT 1340.1000 1334.4000 1341.6000 1335.3000 ;
	    RECT 1343.4000 1334.4000 1344.6000 1335.6000 ;
	    RECT 1345.8000 1335.4501 1347.0000 1335.6000 ;
	    RECT 1369.8000 1335.4501 1371.0000 1335.6000 ;
	    RECT 1345.8000 1334.5500 1371.0000 1335.4501 ;
	    RECT 1345.8000 1334.4000 1347.0000 1334.5500 ;
	    RECT 1369.8000 1334.4000 1371.0000 1334.5500 ;
	    RECT 1340.1000 1323.3000 1341.3000 1334.4000 ;
	    RECT 1342.5000 1332.6000 1343.4000 1333.5000 ;
	    RECT 1369.8000 1333.2001 1371.0000 1333.5000 ;
	    RECT 1342.2001 1331.4000 1343.4000 1332.6000 ;
	    RECT 1342.5000 1323.3000 1343.7001 1329.3000 ;
	    RECT 1369.8000 1323.3000 1371.0000 1329.3000 ;
	    RECT 1372.2001 1323.3000 1373.4000 1336.5000 ;
	    RECT 1377.0000 1335.4501 1378.2001 1335.6000 ;
	    RECT 1393.8000 1335.4501 1395.0000 1335.6000 ;
	    RECT 1377.0000 1334.5500 1395.0000 1335.4501 ;
	    RECT 1377.0000 1334.4000 1378.2001 1334.5500 ;
	    RECT 1393.8000 1334.4000 1395.0000 1334.5500 ;
	    RECT 1393.8000 1333.2001 1395.0000 1333.5000 ;
	    RECT 1374.6000 1323.3000 1375.8000 1329.3000 ;
	    RECT 1393.8000 1323.3000 1395.0000 1329.3000 ;
	    RECT 1396.2001 1323.3000 1397.4000 1336.5000 ;
	    RECT 1398.6000 1323.3000 1399.8000 1329.3000 ;
	    RECT 1417.8000 1323.3000 1419.0000 1329.3000 ;
	    RECT 1420.2001 1323.3000 1421.4000 1336.5000 ;
	    RECT 1422.6000 1335.4501 1423.8000 1335.6000 ;
	    RECT 1444.2001 1335.4501 1445.4000 1335.6000 ;
	    RECT 1422.6000 1334.5500 1445.4000 1335.4501 ;
	    RECT 1422.6000 1334.4000 1423.8000 1334.5500 ;
	    RECT 1444.2001 1334.4000 1445.4000 1334.5500 ;
	    RECT 1446.6000 1334.4000 1447.8000 1335.6000 ;
	    RECT 1449.6000 1335.3000 1450.5000 1340.4000 ;
	    RECT 1451.4000 1339.5000 1452.6000 1339.8000 ;
	    RECT 1451.4000 1337.4000 1452.6000 1338.6000 ;
	    RECT 1473.0000 1335.4501 1474.2001 1335.6000 ;
	    RECT 1477.8000 1335.4501 1479.0000 1335.6000 ;
	    RECT 1449.6000 1334.4000 1451.1000 1335.3000 ;
	    RECT 1422.6000 1333.2001 1423.8000 1333.5000 ;
	    RECT 1447.8000 1332.6000 1448.7001 1333.5000 ;
	    RECT 1447.8000 1331.4000 1449.0000 1332.6000 ;
	    RECT 1422.6000 1323.3000 1423.8000 1329.3000 ;
	    RECT 1447.5000 1323.3000 1448.7001 1329.3000 ;
	    RECT 1449.9000 1323.3000 1451.1000 1334.4000 ;
	    RECT 1453.8000 1323.3000 1455.0000 1335.3000 ;
	    RECT 1473.0000 1334.5500 1479.0000 1335.4501 ;
	    RECT 1473.0000 1334.4000 1474.2001 1334.5500 ;
	    RECT 1477.8000 1334.4000 1479.0000 1334.5500 ;
	    RECT 1480.8000 1335.3000 1481.7001 1340.4000 ;
	    RECT 1482.6000 1339.5000 1483.8000 1339.8000 ;
	    RECT 1482.6000 1338.4501 1483.8000 1338.6000 ;
	    RECT 1487.5500 1338.4501 1488.4501 1340.5500 ;
	    RECT 1499.4000 1340.4000 1500.6000 1340.5500 ;
	    RECT 1518.6000 1341.4501 1519.8000 1341.6000 ;
	    RECT 1540.2001 1341.4501 1541.4000 1341.6000 ;
	    RECT 1518.6000 1340.5500 1541.4000 1341.4501 ;
	    RECT 1518.6000 1340.4000 1519.8000 1340.5500 ;
	    RECT 1540.2001 1340.4000 1541.4000 1340.5500 ;
	    RECT 1542.6000 1340.4000 1543.8000 1341.6000 ;
	    RECT 1544.7001 1340.4000 1546.5000 1341.6000 ;
	    RECT 1548.6000 1340.7001 1548.9000 1342.2001 ;
	    RECT 1549.8000 1340.4000 1551.0000 1341.6000 ;
	    RECT 1482.6000 1337.5500 1488.4501 1338.4501 ;
	    RECT 1482.6000 1337.4000 1483.8000 1337.5500 ;
	    RECT 1480.8000 1334.4000 1482.3000 1335.3000 ;
	    RECT 1479.0000 1332.6000 1479.9000 1333.5000 ;
	    RECT 1479.0000 1331.4000 1480.2001 1332.6000 ;
	    RECT 1478.7001 1323.3000 1479.9000 1329.3000 ;
	    RECT 1481.1000 1323.3000 1482.3000 1334.4000 ;
	    RECT 1485.0000 1323.3000 1486.2001 1335.3000 ;
	    RECT 1499.4000 1323.3000 1500.6000 1339.5000 ;
	    RECT 1501.8000 1323.3000 1503.0000 1329.3000 ;
	    RECT 1516.2001 1323.3000 1517.4000 1329.3000 ;
	    RECT 1518.6000 1323.3000 1519.8000 1339.5000 ;
	    RECT 1540.2001 1335.4501 1541.4000 1335.6000 ;
	    RECT 1542.6000 1335.4501 1543.8000 1335.6000 ;
	    RECT 1540.2001 1334.5500 1543.8000 1335.4501 ;
	    RECT 1540.2001 1334.4000 1541.4000 1334.5500 ;
	    RECT 1542.6000 1334.4000 1543.8000 1334.5500 ;
	    RECT 1545.6000 1335.3000 1546.5000 1340.4000 ;
	    RECT 1547.4000 1339.5000 1548.6000 1339.8000 ;
	    RECT 1547.4000 1337.4000 1548.6000 1338.6000 ;
	    RECT 1545.6000 1334.4000 1547.1000 1335.3000 ;
	    RECT 1543.8000 1332.6000 1544.7001 1333.5000 ;
	    RECT 1543.8000 1331.4000 1545.0000 1332.6000 ;
	    RECT 1543.5000 1323.3000 1544.7001 1329.3000 ;
	    RECT 1545.9000 1323.3000 1547.1000 1334.4000 ;
	    RECT 1549.8000 1323.3000 1551.0000 1335.3000 ;
	    RECT 1.2000 1320.6000 1569.0000 1322.4000 ;
	    RECT 18.6000 1313.7001 19.8000 1319.7001 ;
	    RECT 21.0000 1306.5000 22.2000 1319.7001 ;
	    RECT 23.4000 1313.7001 24.6000 1319.7001 ;
	    RECT 50.7000 1313.7001 51.9000 1319.7001 ;
	    RECT 51.0000 1310.4000 52.2000 1311.6000 ;
	    RECT 23.4000 1309.5000 24.6000 1309.8000 ;
	    RECT 51.0000 1309.5000 51.9000 1310.4000 ;
	    RECT 53.1000 1308.6000 54.3000 1319.7001 ;
	    RECT 23.4000 1307.4000 24.6000 1308.6000 ;
	    RECT 49.8000 1307.4000 51.0000 1308.6000 ;
	    RECT 52.8000 1307.7001 54.3000 1308.6000 ;
	    RECT 57.0000 1307.7001 58.2000 1319.7001 ;
	    RECT 81.0000 1307.7001 82.2000 1319.7001 ;
	    RECT 84.9000 1308.6000 86.1000 1319.7001 ;
	    RECT 87.3000 1313.7001 88.5000 1319.7001 ;
	    RECT 107.4000 1313.7001 108.6000 1319.7001 ;
	    RECT 87.0000 1310.4000 88.2000 1311.6000 ;
	    RECT 87.3000 1309.5000 88.2000 1310.4000 ;
	    RECT 84.9000 1307.7001 86.4000 1308.6000 ;
	    RECT 21.0000 1305.4501 22.2000 1305.6000 ;
	    RECT 49.9500 1305.4501 50.8500 1307.4000 ;
	    RECT 21.0000 1304.5500 50.8500 1305.4501 ;
	    RECT 21.0000 1304.4000 22.2000 1304.5500 ;
	    RECT 18.6000 1301.4000 19.8000 1302.6000 ;
	    RECT 18.6000 1300.2001 19.8000 1300.5000 ;
	    RECT 21.0000 1299.3000 22.2000 1303.5000 ;
	    RECT 52.8000 1302.6000 53.7000 1307.7001 ;
	    RECT 54.6000 1304.4000 55.8000 1305.6000 ;
	    RECT 83.4000 1304.4000 84.6000 1305.6000 ;
	    RECT 54.6000 1303.2001 55.8000 1303.5000 ;
	    RECT 83.4000 1303.2001 84.6000 1303.5000 ;
	    RECT 85.5000 1302.6000 86.4000 1307.7001 ;
	    RECT 88.2000 1307.4000 89.4000 1308.6000 ;
	    RECT 88.3500 1305.4501 89.2500 1307.4000 ;
	    RECT 109.8000 1306.5000 111.0000 1319.7001 ;
	    RECT 112.2000 1313.7001 113.4000 1319.7001 ;
	    RECT 126.6000 1313.7001 127.8000 1319.7001 ;
	    RECT 112.2000 1309.5000 113.4000 1309.8000 ;
	    RECT 112.2000 1308.4501 113.4000 1308.6000 ;
	    RECT 114.6000 1308.4501 115.8000 1308.6000 ;
	    RECT 112.2000 1307.5500 115.8000 1308.4501 ;
	    RECT 112.2000 1307.4000 113.4000 1307.5500 ;
	    RECT 114.6000 1307.4000 115.8000 1307.5500 ;
	    RECT 109.8000 1305.4501 111.0000 1305.6000 ;
	    RECT 88.3500 1304.5500 111.0000 1305.4501 ;
	    RECT 109.8000 1304.4000 111.0000 1304.5500 ;
	    RECT 129.0000 1303.5000 130.2000 1319.7001 ;
	    RECT 153.0000 1307.7001 154.2000 1319.7001 ;
	    RECT 156.9000 1308.6000 158.1000 1319.7001 ;
	    RECT 159.3000 1313.7001 160.5000 1319.7001 ;
	    RECT 179.4000 1313.7001 180.6000 1319.7001 ;
	    RECT 159.0000 1310.4000 160.2000 1311.6000 ;
	    RECT 159.3000 1309.5000 160.2000 1310.4000 ;
	    RECT 179.4000 1309.5000 180.6000 1309.8000 ;
	    RECT 156.9000 1307.7001 158.4000 1308.6000 ;
	    RECT 155.4000 1305.4501 156.6000 1305.6000 ;
	    RECT 150.7500 1304.5500 156.6000 1305.4501 ;
	    RECT 49.8000 1301.4000 51.0000 1302.6000 ;
	    RECT 51.9000 1301.4000 53.7000 1302.6000 ;
	    RECT 57.0000 1302.4501 58.2000 1302.6000 ;
	    RECT 81.0000 1302.4501 82.2000 1302.6000 ;
	    RECT 55.8000 1300.8000 56.1000 1302.3000 ;
	    RECT 57.0000 1301.5500 82.2000 1302.4501 ;
	    RECT 57.0000 1301.4000 58.2000 1301.5500 ;
	    RECT 81.0000 1301.4000 82.2000 1301.5500 ;
	    RECT 83.1000 1300.8000 83.4000 1302.3000 ;
	    RECT 85.5000 1301.4000 87.3000 1302.6000 ;
	    RECT 88.2000 1302.4501 89.4000 1302.6000 ;
	    RECT 105.0000 1302.4501 106.2000 1302.6000 ;
	    RECT 88.2000 1301.5500 106.2000 1302.4501 ;
	    RECT 88.2000 1301.4000 89.4000 1301.5500 ;
	    RECT 105.0000 1301.4000 106.2000 1301.5500 ;
	    RECT 107.4000 1301.4000 108.6000 1302.6000 ;
	    RECT 50.1000 1299.3000 51.0000 1300.5000 ;
	    RECT 52.5000 1299.3000 57.9000 1299.9000 ;
	    RECT 81.3000 1299.3000 86.7000 1299.9000 ;
	    RECT 88.2000 1299.3000 89.1000 1300.5000 ;
	    RECT 107.4000 1300.2001 108.6000 1300.5000 ;
	    RECT 109.8000 1299.3000 111.0000 1303.5000 ;
	    RECT 129.0000 1302.4501 130.2000 1302.6000 ;
	    RECT 150.7500 1302.4501 151.6500 1304.5500 ;
	    RECT 155.4000 1304.4000 156.6000 1304.5500 ;
	    RECT 155.4000 1303.2001 156.6000 1303.5000 ;
	    RECT 157.5000 1302.6000 158.4000 1307.7001 ;
	    RECT 160.2000 1308.4501 161.4000 1308.6000 ;
	    RECT 162.6000 1308.4501 163.8000 1308.6000 ;
	    RECT 160.2000 1307.5500 163.8000 1308.4501 ;
	    RECT 160.2000 1307.4000 161.4000 1307.5500 ;
	    RECT 162.6000 1307.4000 163.8000 1307.5500 ;
	    RECT 179.4000 1307.4000 180.6000 1308.6000 ;
	    RECT 181.8000 1306.5000 183.0000 1319.7001 ;
	    RECT 184.2000 1313.7001 185.4000 1319.7001 ;
	    RECT 196.2000 1313.7001 197.4000 1319.7001 ;
	    RECT 181.8000 1305.4501 183.0000 1305.6000 ;
	    RECT 196.2000 1305.4501 197.4000 1305.6000 ;
	    RECT 181.8000 1304.5500 197.4000 1305.4501 ;
	    RECT 181.8000 1304.4000 183.0000 1304.5500 ;
	    RECT 196.2000 1304.4000 197.4000 1304.5500 ;
	    RECT 198.6000 1303.5000 199.8000 1319.7001 ;
	    RECT 233.1000 1313.7001 234.3000 1319.7001 ;
	    RECT 233.4000 1310.4000 234.6000 1311.6000 ;
	    RECT 233.4000 1309.5000 234.3000 1310.4000 ;
	    RECT 235.5000 1308.6000 236.7000 1319.7001 ;
	    RECT 232.2000 1307.4000 233.4000 1308.6000 ;
	    RECT 235.2000 1307.7001 236.7000 1308.6000 ;
	    RECT 239.4000 1307.7001 240.6000 1319.7001 ;
	    RECT 253.8000 1313.7001 255.0000 1319.7001 ;
	    RECT 129.0000 1301.5500 151.6500 1302.4501 ;
	    RECT 129.0000 1301.4000 130.2000 1301.5500 ;
	    RECT 153.0000 1301.4000 154.2000 1302.6000 ;
	    RECT 155.1000 1300.8000 155.4000 1302.3000 ;
	    RECT 157.5000 1301.4000 159.3000 1302.6000 ;
	    RECT 160.2000 1301.4000 161.4000 1302.6000 ;
	    RECT 18.6000 1293.3000 19.8000 1299.3000 ;
	    RECT 21.0000 1298.4000 23.7000 1299.3000 ;
	    RECT 22.5000 1293.3000 23.7000 1298.4000 ;
	    RECT 49.8000 1293.3000 51.0000 1299.3000 ;
	    RECT 52.2000 1299.0000 58.2000 1299.3000 ;
	    RECT 52.2000 1293.3000 53.4000 1299.0000 ;
	    RECT 54.6000 1293.3000 55.8000 1298.1000 ;
	    RECT 57.0000 1293.3000 58.2000 1299.0000 ;
	    RECT 81.0000 1299.0000 87.0000 1299.3000 ;
	    RECT 81.0000 1293.3000 82.2000 1299.0000 ;
	    RECT 83.4000 1293.3000 84.6000 1298.1000 ;
	    RECT 85.8000 1293.3000 87.0000 1299.0000 ;
	    RECT 88.2000 1293.3000 89.4000 1299.3000 ;
	    RECT 107.4000 1293.3000 108.6000 1299.3000 ;
	    RECT 109.8000 1298.4000 112.5000 1299.3000 ;
	    RECT 126.6000 1298.4000 127.8000 1299.6000 ;
	    RECT 111.3000 1293.3000 112.5000 1298.4000 ;
	    RECT 126.6000 1297.2001 127.8000 1297.5000 ;
	    RECT 126.6000 1293.3000 127.8000 1296.3000 ;
	    RECT 129.0000 1293.3000 130.2000 1300.5000 ;
	    RECT 153.3000 1299.3000 158.7000 1299.9000 ;
	    RECT 160.2000 1299.3000 161.1000 1300.5000 ;
	    RECT 181.8000 1299.3000 183.0000 1303.5000 ;
	    RECT 235.2000 1302.6000 236.1000 1307.7001 ;
	    RECT 237.0000 1304.4000 238.2000 1305.6000 ;
	    RECT 256.2000 1303.5000 257.4000 1319.7001 ;
	    RECT 280.2000 1307.7001 281.4000 1319.7001 ;
	    RECT 284.1000 1308.6000 285.3000 1319.7001 ;
	    RECT 286.5000 1313.7001 287.7000 1319.7001 ;
	    RECT 333.0000 1317.4501 334.2000 1317.6000 ;
	    RECT 349.8000 1317.4501 351.0000 1317.6000 ;
	    RECT 373.8000 1317.4501 375.0000 1317.6000 ;
	    RECT 333.0000 1316.5500 375.0000 1317.4501 ;
	    RECT 333.0000 1316.4000 334.2000 1316.5500 ;
	    RECT 349.8000 1316.4000 351.0000 1316.5500 ;
	    RECT 373.8000 1316.4000 375.0000 1316.5500 ;
	    RECT 419.4000 1313.7001 420.6000 1319.7001 ;
	    RECT 421.8000 1312.5000 423.0000 1319.7001 ;
	    RECT 424.2000 1313.7001 425.4000 1319.7001 ;
	    RECT 426.6000 1312.8000 427.8000 1319.7001 ;
	    RECT 429.0000 1313.7001 430.2000 1319.7001 ;
	    RECT 423.9000 1311.9000 427.8000 1312.8000 ;
	    RECT 286.2000 1310.4000 287.4000 1311.6000 ;
	    RECT 381.0000 1311.4501 382.2000 1311.6000 ;
	    RECT 421.8000 1311.4501 423.0000 1311.6000 ;
	    RECT 381.0000 1310.5500 423.0000 1311.4501 ;
	    RECT 381.0000 1310.4000 382.2000 1310.5500 ;
	    RECT 421.8000 1310.4000 423.0000 1310.5500 ;
	    RECT 286.5000 1309.5000 287.4000 1310.4000 ;
	    RECT 423.9000 1309.5000 424.8000 1311.9000 ;
	    RECT 431.4000 1311.6000 432.6000 1319.7001 ;
	    RECT 433.8000 1313.7001 435.0000 1319.7001 ;
	    RECT 436.2000 1315.5000 437.4000 1319.7001 ;
	    RECT 438.6000 1315.5000 439.8000 1319.7001 ;
	    RECT 441.0000 1315.5000 442.2000 1319.7001 ;
	    RECT 433.5000 1311.6000 439.8000 1312.8000 ;
	    RECT 428.7000 1310.4000 432.6000 1311.6000 ;
	    RECT 443.4000 1310.4000 444.6000 1319.7001 ;
	    RECT 445.8000 1313.7001 447.0000 1319.7001 ;
	    RECT 448.2000 1312.5000 449.4000 1319.7001 ;
	    RECT 450.6000 1313.7001 451.8000 1319.7001 ;
	    RECT 453.0000 1312.5000 454.2000 1319.7001 ;
	    RECT 455.4000 1315.5000 456.6000 1319.7001 ;
	    RECT 457.8000 1315.5000 459.0000 1319.7001 ;
	    RECT 460.2000 1313.7001 461.4000 1319.7001 ;
	    RECT 462.6000 1312.8000 463.8000 1319.7001 ;
	    RECT 465.0000 1313.7001 466.2000 1320.6000 ;
	    RECT 467.4000 1314.6000 468.6000 1319.7001 ;
	    RECT 467.4000 1313.7001 468.9000 1314.6000 ;
	    RECT 469.8000 1313.7001 471.0000 1319.7001 ;
	    RECT 489.0000 1313.7001 490.2000 1319.7001 ;
	    RECT 468.0000 1312.8000 468.9000 1313.7001 ;
	    RECT 460.8000 1311.6000 467.1000 1312.8000 ;
	    RECT 468.0000 1311.9000 471.0000 1312.8000 ;
	    RECT 448.2000 1310.4000 452.1000 1311.6000 ;
	    RECT 453.0000 1310.7001 461.7000 1311.6000 ;
	    RECT 466.2000 1311.0000 467.1000 1311.6000 ;
	    RECT 436.2000 1309.5000 437.4000 1309.8000 ;
	    RECT 284.1000 1307.7001 285.6000 1308.6000 ;
	    RECT 282.6000 1305.4501 283.8000 1305.6000 ;
	    RECT 277.9500 1304.5500 283.8000 1305.4501 ;
	    RECT 237.0000 1303.2001 238.2000 1303.5000 ;
	    RECT 184.2000 1301.4000 185.4000 1302.6000 ;
	    RECT 198.6000 1302.4501 199.8000 1302.6000 ;
	    RECT 229.8000 1302.4501 231.0000 1302.6000 ;
	    RECT 198.6000 1301.5500 231.0000 1302.4501 ;
	    RECT 198.6000 1301.4000 199.8000 1301.5500 ;
	    RECT 229.8000 1301.4000 231.0000 1301.5500 ;
	    RECT 232.2000 1301.4000 233.4000 1302.6000 ;
	    RECT 234.3000 1301.4000 236.1000 1302.6000 ;
	    RECT 238.2000 1300.8000 238.5000 1302.3000 ;
	    RECT 239.4000 1301.4000 240.6000 1302.6000 ;
	    RECT 256.2000 1302.4501 257.4000 1302.6000 ;
	    RECT 277.9500 1302.4501 278.8500 1304.5500 ;
	    RECT 282.6000 1304.4000 283.8000 1304.5500 ;
	    RECT 282.6000 1303.2001 283.8000 1303.5000 ;
	    RECT 284.7000 1302.6000 285.6000 1307.7001 ;
	    RECT 287.4000 1307.4000 288.6000 1308.6000 ;
	    RECT 421.8000 1308.0000 423.0000 1309.5000 ;
	    RECT 421.5000 1306.8000 423.0000 1308.0000 ;
	    RECT 423.9000 1308.6000 437.4000 1309.5000 ;
	    RECT 441.0000 1309.5000 442.2000 1309.8000 ;
	    RECT 453.0000 1309.5000 453.9000 1310.7001 ;
	    RECT 462.6000 1309.8000 464.7000 1310.7001 ;
	    RECT 466.2000 1309.8000 468.6000 1311.0000 ;
	    RECT 441.0000 1308.6000 453.9000 1309.5000 ;
	    RECT 455.4000 1309.5000 464.7000 1309.8000 ;
	    RECT 455.4000 1308.9000 463.5000 1309.5000 ;
	    RECT 455.4000 1308.6000 456.6000 1308.9000 ;
	    RECT 256.2000 1301.5500 278.8500 1302.4501 ;
	    RECT 256.2000 1301.4000 257.4000 1301.5500 ;
	    RECT 280.2000 1301.4000 281.4000 1302.6000 ;
	    RECT 282.3000 1300.8000 282.6000 1302.3000 ;
	    RECT 284.7000 1301.4000 286.5000 1302.6000 ;
	    RECT 287.4000 1302.4501 288.6000 1302.6000 ;
	    RECT 357.0000 1302.4501 358.2000 1302.6000 ;
	    RECT 287.4000 1301.5500 358.2000 1302.4501 ;
	    RECT 287.4000 1301.4000 288.6000 1301.5500 ;
	    RECT 357.0000 1301.4000 358.2000 1301.5500 ;
	    RECT 184.2000 1300.2001 185.4000 1300.5000 ;
	    RECT 153.0000 1299.0000 159.0000 1299.3000 ;
	    RECT 153.0000 1293.3000 154.2000 1299.0000 ;
	    RECT 155.4000 1293.3000 156.6000 1298.1000 ;
	    RECT 157.8000 1293.3000 159.0000 1299.0000 ;
	    RECT 160.2000 1293.3000 161.4000 1299.3000 ;
	    RECT 180.3000 1298.4000 183.0000 1299.3000 ;
	    RECT 180.3000 1293.3000 181.5000 1298.4000 ;
	    RECT 184.2000 1293.3000 185.4000 1299.3000 ;
	    RECT 196.2000 1298.4000 197.4000 1299.6000 ;
	    RECT 196.2000 1297.2001 197.4000 1297.5000 ;
	    RECT 196.2000 1293.3000 197.4000 1296.3000 ;
	    RECT 198.6000 1293.3000 199.8000 1300.5000 ;
	    RECT 232.5000 1299.3000 233.4000 1300.5000 ;
	    RECT 234.9000 1299.3000 240.3000 1299.9000 ;
	    RECT 244.2000 1299.4501 245.4000 1299.6000 ;
	    RECT 253.8000 1299.4501 255.0000 1299.6000 ;
	    RECT 232.2000 1293.3000 233.4000 1299.3000 ;
	    RECT 234.6000 1299.0000 240.6000 1299.3000 ;
	    RECT 234.6000 1293.3000 235.8000 1299.0000 ;
	    RECT 237.0000 1293.3000 238.2000 1298.1000 ;
	    RECT 239.4000 1293.3000 240.6000 1299.0000 ;
	    RECT 244.2000 1298.5500 255.0000 1299.4501 ;
	    RECT 244.2000 1298.4000 245.4000 1298.5500 ;
	    RECT 253.8000 1298.4000 255.0000 1298.5500 ;
	    RECT 253.8000 1297.2001 255.0000 1297.5000 ;
	    RECT 253.8000 1293.3000 255.0000 1296.3000 ;
	    RECT 256.2000 1293.3000 257.4000 1300.5000 ;
	    RECT 280.5000 1299.3000 285.9000 1299.9000 ;
	    RECT 287.4000 1299.3000 288.3000 1300.5000 ;
	    RECT 421.5000 1300.2001 422.7000 1306.8000 ;
	    RECT 423.9000 1305.9000 424.8000 1308.6000 ;
	    RECT 459.9000 1307.7001 461.1000 1308.0000 ;
	    RECT 425.7000 1306.8000 464.1000 1307.7001 ;
	    RECT 465.0000 1307.4000 466.2000 1308.6000 ;
	    RECT 425.7000 1306.5000 426.9000 1306.8000 ;
	    RECT 423.6000 1305.0000 424.8000 1305.9000 ;
	    RECT 433.8000 1305.0000 459.3000 1305.9000 ;
	    RECT 423.6000 1302.0000 424.5000 1305.0000 ;
	    RECT 433.8000 1304.1000 435.0000 1305.0000 ;
	    RECT 460.2000 1304.4000 461.4000 1305.6000 ;
	    RECT 462.3000 1305.0000 468.9000 1305.9000 ;
	    RECT 467.7000 1304.7001 468.9000 1305.0000 ;
	    RECT 425.4000 1302.9000 431.1000 1304.1000 ;
	    RECT 423.6000 1301.1000 425.4000 1302.0000 ;
	    RECT 280.2000 1299.0000 286.2000 1299.3000 ;
	    RECT 280.2000 1293.3000 281.4000 1299.0000 ;
	    RECT 282.6000 1293.3000 283.8000 1298.1000 ;
	    RECT 285.0000 1293.3000 286.2000 1299.0000 ;
	    RECT 287.4000 1293.3000 288.6000 1299.3000 ;
	    RECT 421.5000 1299.0000 423.0000 1300.2001 ;
	    RECT 419.4000 1293.3000 420.6000 1296.3000 ;
	    RECT 421.8000 1293.3000 423.0000 1299.0000 ;
	    RECT 424.2000 1293.3000 425.4000 1301.1000 ;
	    RECT 429.9000 1301.1000 431.1000 1302.9000 ;
	    RECT 429.9000 1300.2001 432.6000 1301.1000 ;
	    RECT 431.4000 1299.3000 432.6000 1300.2001 ;
	    RECT 438.6000 1299.6000 439.8000 1303.8000 ;
	    RECT 443.4000 1302.9000 448.2000 1304.1000 ;
	    RECT 453.9000 1302.9000 456.9000 1304.1000 ;
	    RECT 469.8000 1303.5000 471.0000 1311.9000 ;
	    RECT 491.4000 1306.5000 492.6000 1319.7001 ;
	    RECT 493.8000 1313.7001 495.0000 1319.7001 ;
	    RECT 618.6000 1313.7001 619.8000 1319.7001 ;
	    RECT 621.0000 1312.5000 622.2000 1319.7001 ;
	    RECT 623.4000 1313.7001 624.6000 1319.7001 ;
	    RECT 625.8000 1312.8000 627.0000 1319.7001 ;
	    RECT 628.2000 1313.7001 629.4000 1319.7001 ;
	    RECT 623.1000 1311.9000 627.0000 1312.8000 ;
	    RECT 580.2000 1311.4501 581.4000 1311.6000 ;
	    RECT 621.0000 1311.4501 622.2000 1311.6000 ;
	    RECT 580.2000 1310.5500 622.2000 1311.4501 ;
	    RECT 580.2000 1310.4000 581.4000 1310.5500 ;
	    RECT 621.0000 1310.4000 622.2000 1310.5500 ;
	    RECT 493.8000 1309.5000 495.0000 1309.8000 ;
	    RECT 623.1000 1309.5000 624.0000 1311.9000 ;
	    RECT 630.6000 1311.6000 631.8000 1319.7001 ;
	    RECT 633.0000 1313.7001 634.2000 1319.7001 ;
	    RECT 635.4000 1315.5000 636.6000 1319.7001 ;
	    RECT 637.8000 1315.5000 639.0000 1319.7001 ;
	    RECT 640.2000 1315.5000 641.4000 1319.7001 ;
	    RECT 632.7000 1311.6000 639.0000 1312.8000 ;
	    RECT 627.9000 1310.4000 631.8000 1311.6000 ;
	    RECT 642.6000 1310.4000 643.8000 1319.7001 ;
	    RECT 645.0000 1313.7001 646.2000 1319.7001 ;
	    RECT 647.4000 1312.5000 648.6000 1319.7001 ;
	    RECT 649.8000 1313.7001 651.0000 1319.7001 ;
	    RECT 652.2000 1312.5000 653.4000 1319.7001 ;
	    RECT 654.6000 1315.5000 655.8000 1319.7001 ;
	    RECT 657.0000 1315.5000 658.2000 1319.7001 ;
	    RECT 659.4000 1313.7001 660.6000 1319.7001 ;
	    RECT 661.8000 1312.8000 663.0000 1319.7001 ;
	    RECT 664.2000 1313.7001 665.4000 1320.6000 ;
	    RECT 666.6000 1314.6000 667.8000 1319.7001 ;
	    RECT 666.6000 1313.7001 668.1000 1314.6000 ;
	    RECT 669.0000 1313.7001 670.2000 1319.7001 ;
	    RECT 688.2000 1313.7001 689.4000 1319.7001 ;
	    RECT 667.2000 1312.8000 668.1000 1313.7001 ;
	    RECT 660.0000 1311.6000 666.3000 1312.8000 ;
	    RECT 667.2000 1311.9000 670.2000 1312.8000 ;
	    RECT 647.4000 1310.4000 651.3000 1311.6000 ;
	    RECT 652.2000 1310.7001 660.9000 1311.6000 ;
	    RECT 665.4000 1311.0000 666.3000 1311.6000 ;
	    RECT 635.4000 1309.5000 636.6000 1309.8000 ;
	    RECT 493.8000 1308.4501 495.0000 1308.6000 ;
	    RECT 618.6000 1308.4501 619.8000 1308.6000 ;
	    RECT 493.8000 1307.5500 619.8000 1308.4501 ;
	    RECT 621.0000 1308.0000 622.2000 1309.5000 ;
	    RECT 493.8000 1307.4000 495.0000 1307.5500 ;
	    RECT 618.6000 1307.4000 619.8000 1307.5500 ;
	    RECT 620.7000 1306.8000 622.2000 1308.0000 ;
	    RECT 623.1000 1308.6000 636.6000 1309.5000 ;
	    RECT 640.2000 1309.5000 641.4000 1309.8000 ;
	    RECT 652.2000 1309.5000 653.1000 1310.7001 ;
	    RECT 661.8000 1309.8000 663.9000 1310.7001 ;
	    RECT 665.4000 1309.8000 667.8000 1311.0000 ;
	    RECT 640.2000 1308.6000 653.1000 1309.5000 ;
	    RECT 654.6000 1309.5000 663.9000 1309.8000 ;
	    RECT 654.6000 1308.9000 662.7000 1309.5000 ;
	    RECT 654.6000 1308.6000 655.8000 1308.9000 ;
	    RECT 472.2000 1305.4501 473.4000 1305.6000 ;
	    RECT 491.4000 1305.4501 492.6000 1305.6000 ;
	    RECT 472.2000 1304.5500 492.6000 1305.4501 ;
	    RECT 472.2000 1304.4000 473.4000 1304.5500 ;
	    RECT 491.4000 1304.4000 492.6000 1304.5500 ;
	    RECT 442.8000 1301.7001 444.0000 1302.0000 ;
	    RECT 442.8000 1300.8000 449.4000 1301.7001 ;
	    RECT 450.6000 1301.4000 451.8000 1302.6000 ;
	    RECT 448.2000 1300.5000 449.4000 1300.8000 ;
	    RECT 450.6000 1300.2001 451.8000 1300.5000 ;
	    RECT 429.0000 1293.3000 430.2000 1299.3000 ;
	    RECT 431.4000 1298.1000 435.0000 1299.3000 ;
	    RECT 438.6000 1298.4000 440.1000 1299.6000 ;
	    RECT 444.6000 1298.4000 444.9000 1299.6000 ;
	    RECT 445.8000 1298.4000 447.0000 1299.6000 ;
	    RECT 448.2000 1299.3000 449.4000 1299.6000 ;
	    RECT 453.9000 1299.3000 455.1000 1302.9000 ;
	    RECT 457.8000 1302.3000 471.0000 1303.5000 ;
	    RECT 462.9000 1300.2001 467.4000 1301.4000 ;
	    RECT 462.9000 1299.3000 464.1000 1300.2001 ;
	    RECT 448.2000 1298.4000 455.1000 1299.3000 ;
	    RECT 433.8000 1293.3000 435.0000 1298.1000 ;
	    RECT 460.2000 1298.1000 464.1000 1299.3000 ;
	    RECT 436.2000 1293.3000 437.4000 1297.5000 ;
	    RECT 438.6000 1293.3000 439.8000 1297.5000 ;
	    RECT 441.0000 1293.3000 442.2000 1297.5000 ;
	    RECT 443.4000 1293.3000 444.6000 1297.5000 ;
	    RECT 445.8000 1293.3000 447.0000 1296.3000 ;
	    RECT 448.2000 1293.3000 449.4000 1297.5000 ;
	    RECT 450.6000 1293.3000 451.8000 1296.3000 ;
	    RECT 453.0000 1293.3000 454.2000 1297.5000 ;
	    RECT 455.4000 1293.3000 456.6000 1297.5000 ;
	    RECT 457.8000 1293.3000 459.0000 1297.5000 ;
	    RECT 460.2000 1293.3000 461.4000 1298.1000 ;
	    RECT 465.0000 1293.3000 466.2000 1299.3000 ;
	    RECT 469.8000 1293.3000 471.0000 1302.3000 ;
	    RECT 479.4000 1302.4501 480.6000 1302.6000 ;
	    RECT 489.0000 1302.4501 490.2000 1302.6000 ;
	    RECT 479.4000 1301.5500 490.2000 1302.4501 ;
	    RECT 479.4000 1301.4000 480.6000 1301.5500 ;
	    RECT 489.0000 1301.4000 490.2000 1301.5500 ;
	    RECT 489.0000 1300.2001 490.2000 1300.5000 ;
	    RECT 491.4000 1299.3000 492.6000 1303.5000 ;
	    RECT 620.7000 1300.2001 621.9000 1306.8000 ;
	    RECT 623.1000 1305.9000 624.0000 1308.6000 ;
	    RECT 659.1000 1307.7001 660.3000 1308.0000 ;
	    RECT 624.9000 1306.8000 663.3000 1307.7001 ;
	    RECT 664.2000 1307.4000 665.4000 1308.6000 ;
	    RECT 624.9000 1306.5000 626.1000 1306.8000 ;
	    RECT 622.8000 1305.0000 624.0000 1305.9000 ;
	    RECT 633.0000 1305.0000 658.5000 1305.9000 ;
	    RECT 622.8000 1302.0000 623.7000 1305.0000 ;
	    RECT 633.0000 1304.1000 634.2000 1305.0000 ;
	    RECT 659.4000 1304.4000 660.6000 1305.6000 ;
	    RECT 661.5000 1305.0000 668.1000 1305.9000 ;
	    RECT 666.9000 1304.7001 668.1000 1305.0000 ;
	    RECT 624.6000 1302.9000 630.3000 1304.1000 ;
	    RECT 622.8000 1301.1000 624.6000 1302.0000 ;
	    RECT 489.0000 1293.3000 490.2000 1299.3000 ;
	    RECT 491.4000 1298.4000 494.1000 1299.3000 ;
	    RECT 620.7000 1299.0000 622.2000 1300.2001 ;
	    RECT 492.9000 1293.3000 494.1000 1298.4000 ;
	    RECT 618.6000 1293.3000 619.8000 1296.3000 ;
	    RECT 621.0000 1293.3000 622.2000 1299.0000 ;
	    RECT 623.4000 1293.3000 624.6000 1301.1000 ;
	    RECT 629.1000 1301.1000 630.3000 1302.9000 ;
	    RECT 629.1000 1300.2001 631.8000 1301.1000 ;
	    RECT 630.6000 1299.3000 631.8000 1300.2001 ;
	    RECT 637.8000 1299.6000 639.0000 1303.8000 ;
	    RECT 642.6000 1302.9000 647.4000 1304.1000 ;
	    RECT 653.1000 1302.9000 656.1000 1304.1000 ;
	    RECT 669.0000 1303.5000 670.2000 1311.9000 ;
	    RECT 690.6000 1303.5000 691.8000 1319.7001 ;
	    RECT 714.6000 1317.4501 715.8000 1317.6000 ;
	    RECT 729.0000 1317.4501 730.2000 1317.6000 ;
	    RECT 714.6000 1316.5500 730.2000 1317.4501 ;
	    RECT 714.6000 1316.4000 715.8000 1316.5500 ;
	    RECT 729.0000 1316.4000 730.2000 1316.5500 ;
	    RECT 743.4000 1307.7001 744.6000 1319.7001 ;
	    RECT 745.8000 1306.8000 747.0000 1319.7001 ;
	    RECT 748.2000 1307.7001 749.4000 1319.7001 ;
	    RECT 750.6000 1306.8000 751.8000 1319.7001 ;
	    RECT 753.0000 1307.7001 754.2000 1319.7001 ;
	    RECT 755.4000 1306.8000 756.6000 1319.7001 ;
	    RECT 757.8000 1307.7001 759.0000 1319.7001 ;
	    RECT 760.2000 1306.8000 761.4000 1319.7001 ;
	    RECT 762.6000 1307.7001 763.8000 1319.7001 ;
	    RECT 774.6000 1313.7001 775.8000 1319.7001 ;
	    RECT 743.4000 1306.5000 747.0000 1306.8000 ;
	    RECT 745.5000 1305.6000 747.0000 1306.5000 ;
	    RECT 748.5000 1305.6000 751.8000 1306.8000 ;
	    RECT 753.3000 1305.6000 756.6000 1306.8000 ;
	    RECT 758.7000 1305.6000 761.4000 1306.8000 ;
	    RECT 702.6000 1305.4501 703.8000 1305.6000 ;
	    RECT 719.4000 1305.4501 720.6000 1305.6000 ;
	    RECT 743.4000 1305.4501 744.6000 1305.6000 ;
	    RECT 702.6000 1304.5500 744.6000 1305.4501 ;
	    RECT 702.6000 1304.4000 703.8000 1304.5500 ;
	    RECT 719.4000 1304.4000 720.6000 1304.5500 ;
	    RECT 743.4000 1304.4000 744.6000 1304.5500 ;
	    RECT 748.5000 1303.5000 749.7000 1305.6000 ;
	    RECT 753.3000 1303.5000 754.5000 1305.6000 ;
	    RECT 758.7000 1303.5000 759.9000 1305.6000 ;
	    RECT 777.0000 1303.5000 778.2000 1319.7001 ;
	    RECT 808.2000 1307.7001 809.4000 1319.7001 ;
	    RECT 812.1000 1307.7001 815.1000 1319.7001 ;
	    RECT 817.8000 1307.7001 819.0000 1319.7001 ;
	    RECT 837.0000 1313.7001 838.2000 1319.7001 ;
	    RECT 837.0000 1309.5000 838.2000 1309.8000 ;
	    RECT 820.2000 1308.4501 821.4000 1308.6000 ;
	    RECT 832.2000 1308.4501 833.4000 1308.6000 ;
	    RECT 810.6000 1304.4000 811.8000 1305.6000 ;
	    RECT 808.2000 1303.5000 809.4000 1303.8000 ;
	    RECT 813.3000 1303.5000 814.2000 1307.7001 ;
	    RECT 820.2000 1307.5500 833.4000 1308.4501 ;
	    RECT 820.2000 1307.4000 821.4000 1307.5500 ;
	    RECT 832.2000 1307.4000 833.4000 1307.5500 ;
	    RECT 834.6000 1308.4501 835.8000 1308.6000 ;
	    RECT 837.0000 1308.4501 838.2000 1308.6000 ;
	    RECT 834.6000 1307.5500 838.2000 1308.4501 ;
	    RECT 834.6000 1307.4000 835.8000 1307.5500 ;
	    RECT 837.0000 1307.4000 838.2000 1307.5500 ;
	    RECT 839.4000 1306.5000 840.6000 1319.7001 ;
	    RECT 841.8000 1313.7001 843.0000 1319.7001 ;
	    RECT 861.9000 1308.9000 863.1000 1319.7001 ;
	    RECT 861.9000 1307.7001 864.6000 1308.9000 ;
	    RECT 865.8000 1307.7001 867.0000 1319.7001 ;
	    RECT 925.8000 1307.7001 927.0000 1319.7001 ;
	    RECT 861.0000 1306.5000 862.2000 1306.8000 ;
	    RECT 815.4000 1305.4501 816.6000 1305.6000 ;
	    RECT 829.8000 1305.4501 831.0000 1305.6000 ;
	    RECT 815.4000 1304.5500 831.0000 1305.4501 ;
	    RECT 815.4000 1304.4000 816.6000 1304.5500 ;
	    RECT 829.8000 1304.4000 831.0000 1304.5500 ;
	    RECT 839.4000 1304.4000 840.6000 1305.6000 ;
	    RECT 861.0000 1304.4000 862.2000 1305.6000 ;
	    RECT 863.4000 1303.5000 864.3000 1307.7001 ;
	    RECT 928.2000 1306.8000 929.4000 1319.7001 ;
	    RECT 930.6000 1307.7001 931.8000 1319.7001 ;
	    RECT 933.0000 1306.8000 934.2000 1319.7001 ;
	    RECT 935.4000 1307.7001 936.6000 1319.7001 ;
	    RECT 937.8000 1306.8000 939.0000 1319.7001 ;
	    RECT 940.2000 1307.7001 941.4000 1319.7001 ;
	    RECT 942.6000 1306.8000 943.8000 1319.7001 ;
	    RECT 945.0000 1307.7001 946.2000 1319.7001 ;
	    RECT 964.2000 1313.7001 965.4000 1319.7001 ;
	    RECT 964.2000 1309.5000 965.4000 1309.8000 ;
	    RECT 964.2000 1307.4000 965.4000 1308.6000 ;
	    RECT 925.8000 1306.5000 929.4000 1306.8000 ;
	    RECT 927.9000 1305.6000 929.4000 1306.5000 ;
	    RECT 930.9000 1305.6000 934.2000 1306.8000 ;
	    RECT 935.7000 1305.6000 939.0000 1306.8000 ;
	    RECT 941.1000 1305.6000 943.8000 1306.8000 ;
	    RECT 966.6000 1306.5000 967.8000 1319.7001 ;
	    RECT 969.0000 1313.7001 970.2000 1319.7001 ;
	    RECT 911.4000 1305.4501 912.6000 1305.6000 ;
	    RECT 923.4000 1305.4501 924.6000 1305.6000 ;
	    RECT 925.8000 1305.4501 927.0000 1305.6000 ;
	    RECT 911.4000 1304.5500 927.0000 1305.4501 ;
	    RECT 911.4000 1304.4000 912.6000 1304.5500 ;
	    RECT 923.4000 1304.4000 924.6000 1304.5500 ;
	    RECT 925.8000 1304.4000 927.0000 1304.5500 ;
	    RECT 930.9000 1303.5000 932.1000 1305.6000 ;
	    RECT 935.7000 1303.5000 936.9000 1305.6000 ;
	    RECT 941.1000 1303.5000 942.3000 1305.6000 ;
	    RECT 966.6000 1305.4501 967.8000 1305.6000 ;
	    RECT 971.4000 1305.4501 972.6000 1305.6000 ;
	    RECT 966.6000 1304.5500 972.6000 1305.4501 ;
	    RECT 966.6000 1304.4000 967.8000 1304.5500 ;
	    RECT 971.4000 1304.4000 972.6000 1304.5500 ;
	    RECT 983.4000 1303.5000 984.6000 1319.7001 ;
	    RECT 985.8000 1313.7001 987.0000 1319.7001 ;
	    RECT 1013.1000 1313.7001 1014.3000 1319.7001 ;
	    RECT 1013.4000 1310.4000 1014.6000 1311.6000 ;
	    RECT 1013.4000 1309.5000 1014.3000 1310.4000 ;
	    RECT 1015.5000 1308.6000 1016.7000 1319.7001 ;
	    RECT 1012.2000 1307.4000 1013.4000 1308.6000 ;
	    RECT 1015.2000 1307.7001 1016.7000 1308.6000 ;
	    RECT 1019.4000 1307.7001 1020.6000 1319.7001 ;
	    RECT 1024.2001 1319.4000 1025.4000 1320.6000 ;
	    RECT 642.0000 1301.7001 643.2000 1302.0000 ;
	    RECT 642.0000 1300.8000 648.6000 1301.7001 ;
	    RECT 649.8000 1301.4000 651.0000 1302.6000 ;
	    RECT 647.4000 1300.5000 648.6000 1300.8000 ;
	    RECT 649.8000 1300.2001 651.0000 1300.5000 ;
	    RECT 628.2000 1293.3000 629.4000 1299.3000 ;
	    RECT 630.6000 1298.1000 634.2000 1299.3000 ;
	    RECT 637.8000 1298.4000 639.3000 1299.6000 ;
	    RECT 643.8000 1298.4000 644.1000 1299.6000 ;
	    RECT 645.0000 1298.4000 646.2000 1299.6000 ;
	    RECT 647.4000 1299.3000 648.6000 1299.6000 ;
	    RECT 653.1000 1299.3000 654.3000 1302.9000 ;
	    RECT 657.0000 1302.3000 670.2000 1303.5000 ;
	    RECT 662.1000 1300.2001 666.6000 1301.4000 ;
	    RECT 662.1000 1299.3000 663.3000 1300.2001 ;
	    RECT 647.4000 1298.4000 654.3000 1299.3000 ;
	    RECT 633.0000 1293.3000 634.2000 1298.1000 ;
	    RECT 659.4000 1298.1000 663.3000 1299.3000 ;
	    RECT 635.4000 1293.3000 636.6000 1297.5000 ;
	    RECT 637.8000 1293.3000 639.0000 1297.5000 ;
	    RECT 640.2000 1293.3000 641.4000 1297.5000 ;
	    RECT 642.6000 1293.3000 643.8000 1297.5000 ;
	    RECT 645.0000 1293.3000 646.2000 1296.3000 ;
	    RECT 647.4000 1293.3000 648.6000 1297.5000 ;
	    RECT 649.8000 1293.3000 651.0000 1296.3000 ;
	    RECT 652.2000 1293.3000 653.4000 1297.5000 ;
	    RECT 654.6000 1293.3000 655.8000 1297.5000 ;
	    RECT 657.0000 1293.3000 658.2000 1297.5000 ;
	    RECT 659.4000 1293.3000 660.6000 1298.1000 ;
	    RECT 664.2000 1293.3000 665.4000 1299.3000 ;
	    RECT 669.0000 1293.3000 670.2000 1302.3000 ;
	    RECT 690.6000 1302.4501 691.8000 1302.6000 ;
	    RECT 724.2000 1302.4501 725.4000 1302.6000 ;
	    RECT 690.6000 1301.5500 725.4000 1302.4501 ;
	    RECT 690.6000 1301.4000 691.8000 1301.5500 ;
	    RECT 724.2000 1301.4000 725.4000 1301.5500 ;
	    RECT 743.4000 1301.4000 744.6000 1303.5000 ;
	    RECT 745.8000 1302.3000 749.7000 1303.5000 ;
	    RECT 750.9000 1302.3000 754.5000 1303.5000 ;
	    RECT 756.0000 1302.3000 759.9000 1303.5000 ;
	    RECT 761.1000 1302.3000 761.7000 1303.5000 ;
	    RECT 810.6000 1303.2001 811.8000 1303.5000 ;
	    RECT 815.4000 1303.2001 816.6000 1303.5000 ;
	    RECT 777.0000 1302.4501 778.2000 1302.6000 ;
	    RECT 808.2000 1302.4501 809.4000 1302.6000 ;
	    RECT 748.5000 1301.4000 749.7000 1302.3000 ;
	    RECT 753.3000 1301.4000 754.5000 1302.3000 ;
	    RECT 758.7000 1301.4000 759.9000 1302.3000 ;
	    RECT 777.0000 1301.5500 809.4000 1302.4501 ;
	    RECT 777.0000 1301.4000 778.2000 1301.5500 ;
	    RECT 808.2000 1301.4000 809.4000 1301.5500 ;
	    RECT 810.6000 1301.4000 812.1000 1302.3000 ;
	    RECT 813.0000 1301.4000 814.2000 1302.6000 ;
	    RECT 676.2000 1299.4501 677.4000 1299.6000 ;
	    RECT 688.2000 1299.4501 689.4000 1299.6000 ;
	    RECT 676.2000 1298.5500 689.4000 1299.4501 ;
	    RECT 676.2000 1298.4000 677.4000 1298.5500 ;
	    RECT 688.2000 1298.4000 689.4000 1298.5500 ;
	    RECT 688.2000 1297.2001 689.4000 1297.5000 ;
	    RECT 688.2000 1293.3000 689.4000 1296.3000 ;
	    RECT 690.6000 1293.3000 691.8000 1300.5000 ;
	    RECT 743.4000 1300.2001 747.0000 1301.4000 ;
	    RECT 748.5000 1300.2001 751.8000 1301.4000 ;
	    RECT 753.3000 1300.2001 756.6000 1301.4000 ;
	    RECT 758.7000 1300.2001 761.4000 1301.4000 ;
	    RECT 743.4000 1293.3000 744.6000 1299.3000 ;
	    RECT 745.8000 1293.3000 747.0000 1300.2001 ;
	    RECT 748.2000 1293.3000 749.4000 1299.3000 ;
	    RECT 750.6000 1293.3000 751.8000 1300.2001 ;
	    RECT 753.0000 1293.3000 754.2000 1299.3000 ;
	    RECT 755.4000 1293.3000 756.6000 1300.2001 ;
	    RECT 757.8000 1293.3000 759.0000 1299.3000 ;
	    RECT 760.2000 1293.3000 761.4000 1300.2001 ;
	    RECT 765.0000 1299.4501 766.2000 1299.6000 ;
	    RECT 774.6000 1299.4501 775.8000 1299.6000 ;
	    RECT 762.6000 1293.3000 763.8000 1299.3000 ;
	    RECT 765.0000 1298.5500 775.8000 1299.4501 ;
	    RECT 765.0000 1298.4000 766.2000 1298.5500 ;
	    RECT 774.6000 1298.4000 775.8000 1298.5500 ;
	    RECT 774.6000 1297.2001 775.8000 1297.5000 ;
	    RECT 774.6000 1293.3000 775.8000 1296.3000 ;
	    RECT 777.0000 1293.3000 778.2000 1300.5000 ;
	    RECT 810.6000 1299.3000 811.5000 1301.4000 ;
	    RECT 816.6000 1300.8000 816.9000 1302.3000 ;
	    RECT 817.8000 1301.4000 819.0000 1302.6000 ;
	    RECT 813.3000 1299.3000 818.7000 1299.9000 ;
	    RECT 839.4000 1299.3000 840.6000 1303.5000 ;
	    RECT 841.8000 1302.4501 843.0000 1302.6000 ;
	    RECT 863.4000 1302.4501 864.6000 1302.6000 ;
	    RECT 841.8000 1301.5500 864.6000 1302.4501 ;
	    RECT 841.8000 1301.4000 843.0000 1301.5500 ;
	    RECT 863.4000 1301.4000 864.6000 1301.5500 ;
	    RECT 925.8000 1301.4000 927.0000 1303.5000 ;
	    RECT 928.2000 1302.3000 932.1000 1303.5000 ;
	    RECT 933.3000 1302.3000 936.9000 1303.5000 ;
	    RECT 938.4000 1302.3000 942.3000 1303.5000 ;
	    RECT 943.5000 1302.3000 944.1000 1303.5000 ;
	    RECT 945.0000 1302.4501 946.2000 1302.6000 ;
	    RECT 947.4000 1302.4501 948.6000 1302.6000 ;
	    RECT 930.9000 1301.4000 932.1000 1302.3000 ;
	    RECT 935.7000 1301.4000 936.9000 1302.3000 ;
	    RECT 941.1000 1301.4000 942.3000 1302.3000 ;
	    RECT 945.0000 1301.5500 948.6000 1302.4501 ;
	    RECT 945.0000 1301.4000 946.2000 1301.5500 ;
	    RECT 947.4000 1301.4000 948.6000 1301.5500 ;
	    RECT 841.8000 1300.2001 843.0000 1300.5000 ;
	    RECT 808.2000 1294.2001 809.4000 1299.3000 ;
	    RECT 810.6000 1295.1000 811.8000 1299.3000 ;
	    RECT 813.0000 1299.0000 819.0000 1299.3000 ;
	    RECT 813.0000 1294.2001 814.2000 1299.0000 ;
	    RECT 808.2000 1293.3000 814.2000 1294.2001 ;
	    RECT 815.4000 1293.3000 816.6000 1298.1000 ;
	    RECT 817.8000 1293.3000 819.0000 1299.0000 ;
	    RECT 837.9000 1298.4000 840.6000 1299.3000 ;
	    RECT 837.9000 1293.3000 839.1000 1298.4000 ;
	    RECT 841.8000 1293.3000 843.0000 1299.3000 ;
	    RECT 863.4000 1296.3000 864.3000 1300.5000 ;
	    RECT 925.8000 1300.2001 929.4000 1301.4000 ;
	    RECT 930.9000 1300.2001 934.2000 1301.4000 ;
	    RECT 935.7000 1300.2001 939.0000 1301.4000 ;
	    RECT 941.1000 1300.2001 943.8000 1301.4000 ;
	    RECT 865.8000 1298.4000 867.0000 1299.6000 ;
	    RECT 865.8000 1297.2001 867.0000 1297.5000 ;
	    RECT 861.0000 1293.3000 862.2000 1296.3000 ;
	    RECT 863.4000 1293.3000 864.6000 1296.3000 ;
	    RECT 865.8000 1293.3000 867.0000 1296.3000 ;
	    RECT 925.8000 1293.3000 927.0000 1299.3000 ;
	    RECT 928.2000 1293.3000 929.4000 1300.2001 ;
	    RECT 930.6000 1293.3000 931.8000 1299.3000 ;
	    RECT 933.0000 1293.3000 934.2000 1300.2001 ;
	    RECT 935.4000 1293.3000 936.6000 1299.3000 ;
	    RECT 937.8000 1293.3000 939.0000 1300.2001 ;
	    RECT 940.2000 1293.3000 941.4000 1299.3000 ;
	    RECT 942.6000 1293.3000 943.8000 1300.2001 ;
	    RECT 966.6000 1299.3000 967.8000 1303.5000 ;
	    RECT 1015.2000 1302.6000 1016.1000 1307.7001 ;
	    RECT 1017.0000 1305.4501 1018.2000 1305.6000 ;
	    RECT 1017.0000 1304.5500 1025.2500 1305.4501 ;
	    RECT 1017.0000 1304.4000 1018.2000 1304.5500 ;
	    RECT 1017.0000 1303.2001 1018.2000 1303.5000 ;
	    RECT 969.0000 1301.4000 970.2000 1302.6000 ;
	    RECT 983.4000 1302.4501 984.6000 1302.6000 ;
	    RECT 993.0000 1302.4501 994.2000 1302.6000 ;
	    RECT 983.4000 1301.5500 994.2000 1302.4501 ;
	    RECT 983.4000 1301.4000 984.6000 1301.5500 ;
	    RECT 993.0000 1301.4000 994.2000 1301.5500 ;
	    RECT 1012.2000 1301.4000 1013.4000 1302.6000 ;
	    RECT 1014.3000 1301.4000 1016.1000 1302.6000 ;
	    RECT 1018.2000 1300.8000 1018.5000 1302.3000 ;
	    RECT 1019.4000 1301.4000 1020.6000 1302.6000 ;
	    RECT 1024.3500 1302.4501 1025.2500 1304.5500 ;
	    RECT 1031.4000 1303.5000 1032.6000 1319.7001 ;
	    RECT 1033.8000 1313.7001 1035.0000 1319.7001 ;
	    RECT 1045.8000 1303.5000 1047.0000 1319.7001 ;
	    RECT 1048.2001 1313.7001 1049.4000 1319.7001 ;
	    RECT 1180.2001 1313.7001 1181.4000 1319.7001 ;
	    RECT 1182.6000 1312.5000 1183.8000 1319.7001 ;
	    RECT 1185.0000 1313.7001 1186.2001 1319.7001 ;
	    RECT 1187.4000 1312.8000 1188.6000 1319.7001 ;
	    RECT 1189.8000 1313.7001 1191.0000 1319.7001 ;
	    RECT 1184.7001 1311.9000 1188.6000 1312.8000 ;
	    RECT 1048.2001 1311.4501 1049.4000 1311.6000 ;
	    RECT 1182.6000 1311.4501 1183.8000 1311.6000 ;
	    RECT 1048.2001 1310.5500 1183.8000 1311.4501 ;
	    RECT 1048.2001 1310.4000 1049.4000 1310.5500 ;
	    RECT 1182.6000 1310.4000 1183.8000 1310.5500 ;
	    RECT 1184.7001 1309.5000 1185.6000 1311.9000 ;
	    RECT 1192.2001 1311.6000 1193.4000 1319.7001 ;
	    RECT 1194.6000 1313.7001 1195.8000 1319.7001 ;
	    RECT 1197.0000 1315.5000 1198.2001 1319.7001 ;
	    RECT 1199.4000 1315.5000 1200.6000 1319.7001 ;
	    RECT 1201.8000 1315.5000 1203.0000 1319.7001 ;
	    RECT 1194.3000 1311.6000 1200.6000 1312.8000 ;
	    RECT 1189.5000 1310.4000 1193.4000 1311.6000 ;
	    RECT 1204.2001 1310.4000 1205.4000 1319.7001 ;
	    RECT 1206.6000 1313.7001 1207.8000 1319.7001 ;
	    RECT 1209.0000 1312.5000 1210.2001 1319.7001 ;
	    RECT 1211.4000 1313.7001 1212.6000 1319.7001 ;
	    RECT 1213.8000 1312.5000 1215.0000 1319.7001 ;
	    RECT 1216.2001 1315.5000 1217.4000 1319.7001 ;
	    RECT 1218.6000 1315.5000 1219.8000 1319.7001 ;
	    RECT 1221.0000 1313.7001 1222.2001 1319.7001 ;
	    RECT 1223.4000 1312.8000 1224.6000 1319.7001 ;
	    RECT 1225.8000 1313.7001 1227.0000 1320.6000 ;
	    RECT 1228.2001 1314.6000 1229.4000 1319.7001 ;
	    RECT 1228.2001 1313.7001 1229.7001 1314.6000 ;
	    RECT 1230.6000 1313.7001 1231.8000 1319.7001 ;
	    RECT 1249.8000 1313.7001 1251.0000 1319.7001 ;
	    RECT 1228.8000 1312.8000 1229.7001 1313.7001 ;
	    RECT 1221.6000 1311.6000 1227.9000 1312.8000 ;
	    RECT 1228.8000 1311.9000 1231.8000 1312.8000 ;
	    RECT 1209.0000 1310.4000 1212.9000 1311.6000 ;
	    RECT 1213.8000 1310.7001 1222.5000 1311.6000 ;
	    RECT 1227.0000 1311.0000 1227.9000 1311.6000 ;
	    RECT 1197.0000 1309.5000 1198.2001 1309.8000 ;
	    RECT 1182.6000 1308.0000 1183.8000 1309.5000 ;
	    RECT 1182.3000 1306.8000 1183.8000 1308.0000 ;
	    RECT 1184.7001 1308.6000 1198.2001 1309.5000 ;
	    RECT 1201.8000 1309.5000 1203.0000 1309.8000 ;
	    RECT 1213.8000 1309.5000 1214.7001 1310.7001 ;
	    RECT 1223.4000 1309.8000 1225.5000 1310.7001 ;
	    RECT 1227.0000 1309.8000 1229.4000 1311.0000 ;
	    RECT 1201.8000 1308.6000 1214.7001 1309.5000 ;
	    RECT 1216.2001 1309.5000 1225.5000 1309.8000 ;
	    RECT 1216.2001 1308.9000 1224.3000 1309.5000 ;
	    RECT 1216.2001 1308.6000 1217.4000 1308.9000 ;
	    RECT 1031.4000 1302.4501 1032.6000 1302.6000 ;
	    RECT 1024.3500 1301.5500 1032.6000 1302.4501 ;
	    RECT 1031.4000 1301.4000 1032.6000 1301.5500 ;
	    RECT 1045.8000 1301.4000 1047.0000 1302.6000 ;
	    RECT 969.0000 1300.2001 970.2000 1300.5000 ;
	    RECT 945.0000 1293.3000 946.2000 1299.3000 ;
	    RECT 965.1000 1298.4000 967.8000 1299.3000 ;
	    RECT 965.1000 1293.3000 966.3000 1298.4000 ;
	    RECT 969.0000 1293.3000 970.2000 1299.3000 ;
	    RECT 983.4000 1293.3000 984.6000 1300.5000 ;
	    RECT 985.8000 1299.4501 987.0000 1299.6000 ;
	    RECT 1005.0000 1299.4501 1006.2000 1299.6000 ;
	    RECT 985.8000 1298.5500 1006.2000 1299.4501 ;
	    RECT 1012.5000 1299.3000 1013.4000 1300.5000 ;
	    RECT 1014.9000 1299.3000 1020.3000 1299.9000 ;
	    RECT 985.8000 1298.4000 987.0000 1298.5500 ;
	    RECT 1005.0000 1298.4000 1006.2000 1298.5500 ;
	    RECT 985.8000 1297.2001 987.0000 1297.5000 ;
	    RECT 985.8000 1293.3000 987.0000 1296.3000 ;
	    RECT 1012.2000 1293.3000 1013.4000 1299.3000 ;
	    RECT 1014.6000 1299.0000 1020.6000 1299.3000 ;
	    RECT 1014.6000 1293.3000 1015.8000 1299.0000 ;
	    RECT 1017.0000 1293.3000 1018.2000 1298.1000 ;
	    RECT 1019.4000 1293.3000 1020.6000 1299.0000 ;
	    RECT 1031.4000 1293.3000 1032.6000 1300.5000 ;
	    RECT 1033.8000 1299.4501 1035.0000 1299.6000 ;
	    RECT 1041.0000 1299.4501 1042.2001 1299.6000 ;
	    RECT 1033.8000 1298.5500 1042.2001 1299.4501 ;
	    RECT 1033.8000 1298.4000 1035.0000 1298.5500 ;
	    RECT 1041.0000 1298.4000 1042.2001 1298.5500 ;
	    RECT 1033.8000 1297.2001 1035.0000 1297.5000 ;
	    RECT 1033.8000 1293.3000 1035.0000 1296.3000 ;
	    RECT 1045.8000 1293.3000 1047.0000 1300.5000 ;
	    RECT 1182.3000 1300.2001 1183.5000 1306.8000 ;
	    RECT 1184.7001 1305.9000 1185.6000 1308.6000 ;
	    RECT 1220.7001 1307.7001 1221.9000 1308.0000 ;
	    RECT 1186.5000 1306.8000 1224.9000 1307.7001 ;
	    RECT 1225.8000 1307.4000 1227.0000 1308.6000 ;
	    RECT 1186.5000 1306.5000 1187.7001 1306.8000 ;
	    RECT 1184.4000 1305.0000 1185.6000 1305.9000 ;
	    RECT 1194.6000 1305.0000 1220.1000 1305.9000 ;
	    RECT 1184.4000 1302.0000 1185.3000 1305.0000 ;
	    RECT 1194.6000 1304.1000 1195.8000 1305.0000 ;
	    RECT 1221.0000 1304.4000 1222.2001 1305.6000 ;
	    RECT 1223.1000 1305.0000 1229.7001 1305.9000 ;
	    RECT 1228.5000 1304.7001 1229.7001 1305.0000 ;
	    RECT 1186.2001 1302.9000 1191.9000 1304.1000 ;
	    RECT 1184.4000 1301.1000 1186.2001 1302.0000 ;
	    RECT 1048.2001 1298.4000 1049.4000 1299.6000 ;
	    RECT 1182.3000 1299.0000 1183.8000 1300.2001 ;
	    RECT 1048.2001 1297.2001 1049.4000 1297.5000 ;
	    RECT 1072.2001 1296.4501 1073.4000 1296.6000 ;
	    RECT 1177.8000 1296.4501 1179.0000 1296.6000 ;
	    RECT 1048.2001 1293.3000 1049.4000 1296.3000 ;
	    RECT 1072.2001 1295.5500 1179.0000 1296.4501 ;
	    RECT 1072.2001 1295.4000 1073.4000 1295.5500 ;
	    RECT 1177.8000 1295.4000 1179.0000 1295.5500 ;
	    RECT 1180.2001 1293.3000 1181.4000 1296.3000 ;
	    RECT 1182.6000 1293.3000 1183.8000 1299.0000 ;
	    RECT 1185.0000 1293.3000 1186.2001 1301.1000 ;
	    RECT 1190.7001 1301.1000 1191.9000 1302.9000 ;
	    RECT 1190.7001 1300.2001 1193.4000 1301.1000 ;
	    RECT 1192.2001 1299.3000 1193.4000 1300.2001 ;
	    RECT 1199.4000 1299.6000 1200.6000 1303.8000 ;
	    RECT 1204.2001 1302.9000 1209.0000 1304.1000 ;
	    RECT 1214.7001 1302.9000 1217.7001 1304.1000 ;
	    RECT 1230.6000 1303.5000 1231.8000 1311.9000 ;
	    RECT 1252.2001 1306.5000 1253.4000 1319.7001 ;
	    RECT 1254.6000 1313.7001 1255.8000 1319.7001 ;
	    RECT 1276.2001 1319.4000 1277.4000 1320.6000 ;
	    RECT 1254.6000 1309.5000 1255.8000 1309.8000 ;
	    RECT 1254.6000 1308.4501 1255.8000 1308.6000 ;
	    RECT 1269.0000 1308.4501 1270.2001 1308.6000 ;
	    RECT 1254.6000 1307.5500 1270.2001 1308.4501 ;
	    RECT 1278.6000 1307.7001 1279.8000 1319.7001 ;
	    RECT 1282.5000 1308.6000 1283.7001 1319.7001 ;
	    RECT 1284.9000 1313.7001 1286.1000 1319.7001 ;
	    RECT 1300.2001 1313.7001 1301.4000 1319.7001 ;
	    RECT 1284.6000 1310.4000 1285.8000 1311.6000 ;
	    RECT 1284.9000 1309.5000 1285.8000 1310.4000 ;
	    RECT 1282.5000 1307.7001 1284.0000 1308.6000 ;
	    RECT 1254.6000 1307.4000 1255.8000 1307.5500 ;
	    RECT 1269.0000 1307.4000 1270.2001 1307.5500 ;
	    RECT 1252.2001 1305.4501 1253.4000 1305.6000 ;
	    RECT 1278.6000 1305.4501 1279.8000 1305.6000 ;
	    RECT 1252.2001 1304.5500 1279.8000 1305.4501 ;
	    RECT 1252.2001 1304.4000 1253.4000 1304.5500 ;
	    RECT 1278.6000 1304.4000 1279.8000 1304.5500 ;
	    RECT 1281.0000 1304.4000 1282.2001 1305.6000 ;
	    RECT 1203.6000 1301.7001 1204.8000 1302.0000 ;
	    RECT 1203.6000 1300.8000 1210.2001 1301.7001 ;
	    RECT 1211.4000 1301.4000 1212.6000 1302.6000 ;
	    RECT 1209.0000 1300.5000 1210.2001 1300.8000 ;
	    RECT 1211.4000 1300.2001 1212.6000 1300.5000 ;
	    RECT 1189.8000 1293.3000 1191.0000 1299.3000 ;
	    RECT 1192.2001 1298.1000 1195.8000 1299.3000 ;
	    RECT 1199.4000 1298.4000 1200.9000 1299.6000 ;
	    RECT 1205.4000 1298.4000 1205.7001 1299.6000 ;
	    RECT 1206.6000 1298.4000 1207.8000 1299.6000 ;
	    RECT 1209.0000 1299.3000 1210.2001 1299.6000 ;
	    RECT 1214.7001 1299.3000 1215.9000 1302.9000 ;
	    RECT 1218.6000 1302.3000 1231.8000 1303.5000 ;
	    RECT 1223.7001 1300.2001 1228.2001 1301.4000 ;
	    RECT 1223.7001 1299.3000 1224.9000 1300.2001 ;
	    RECT 1209.0000 1298.4000 1215.9000 1299.3000 ;
	    RECT 1194.6000 1293.3000 1195.8000 1298.1000 ;
	    RECT 1221.0000 1298.1000 1224.9000 1299.3000 ;
	    RECT 1197.0000 1293.3000 1198.2001 1297.5000 ;
	    RECT 1199.4000 1293.3000 1200.6000 1297.5000 ;
	    RECT 1201.8000 1293.3000 1203.0000 1297.5000 ;
	    RECT 1204.2001 1293.3000 1205.4000 1297.5000 ;
	    RECT 1206.6000 1293.3000 1207.8000 1296.3000 ;
	    RECT 1209.0000 1293.3000 1210.2001 1297.5000 ;
	    RECT 1211.4000 1293.3000 1212.6000 1296.3000 ;
	    RECT 1213.8000 1293.3000 1215.0000 1297.5000 ;
	    RECT 1216.2001 1293.3000 1217.4000 1297.5000 ;
	    RECT 1218.6000 1293.3000 1219.8000 1297.5000 ;
	    RECT 1221.0000 1293.3000 1222.2001 1298.1000 ;
	    RECT 1225.8000 1293.3000 1227.0000 1299.3000 ;
	    RECT 1230.6000 1293.3000 1231.8000 1302.3000 ;
	    RECT 1233.0000 1302.4501 1234.2001 1302.6000 ;
	    RECT 1249.8000 1302.4501 1251.0000 1302.6000 ;
	    RECT 1233.0000 1301.5500 1251.0000 1302.4501 ;
	    RECT 1233.0000 1301.4000 1234.2001 1301.5500 ;
	    RECT 1249.8000 1301.4000 1251.0000 1301.5500 ;
	    RECT 1249.8000 1300.2001 1251.0000 1300.5000 ;
	    RECT 1252.2001 1299.3000 1253.4000 1303.5000 ;
	    RECT 1281.0000 1303.2001 1282.2001 1303.5000 ;
	    RECT 1283.1000 1302.6000 1284.0000 1307.7001 ;
	    RECT 1285.8000 1307.4000 1287.0000 1308.6000 ;
	    RECT 1302.6000 1303.5000 1303.8000 1319.7001 ;
	    RECT 1326.6000 1307.7001 1327.8000 1319.7001 ;
	    RECT 1330.5000 1308.6000 1331.7001 1319.7001 ;
	    RECT 1332.9000 1313.7001 1334.1000 1319.7001 ;
	    RECT 1336.2001 1319.4000 1337.4000 1320.6000 ;
	    RECT 1465.8000 1313.7001 1467.0000 1319.7001 ;
	    RECT 1468.2001 1314.6000 1469.4000 1319.7001 ;
	    RECT 1467.9000 1313.7001 1469.4000 1314.6000 ;
	    RECT 1470.6000 1313.7001 1471.8000 1320.6000 ;
	    RECT 1467.9000 1312.8000 1468.8000 1313.7001 ;
	    RECT 1473.0000 1312.8000 1474.2001 1319.7001 ;
	    RECT 1475.4000 1313.7001 1476.6000 1319.7001 ;
	    RECT 1477.8000 1315.5000 1479.0000 1319.7001 ;
	    RECT 1480.2001 1315.5000 1481.4000 1319.7001 ;
	    RECT 1465.8000 1311.9000 1468.8000 1312.8000 ;
	    RECT 1332.6000 1310.4000 1333.8000 1311.6000 ;
	    RECT 1332.9000 1309.5000 1333.8000 1310.4000 ;
	    RECT 1330.5000 1307.7001 1332.0000 1308.6000 ;
	    RECT 1329.0000 1305.4501 1330.2001 1305.6000 ;
	    RECT 1324.3500 1304.5500 1330.2001 1305.4501 ;
	    RECT 1276.2001 1302.4501 1277.4000 1302.6000 ;
	    RECT 1278.6000 1302.4501 1279.8000 1302.6000 ;
	    RECT 1276.2001 1301.5500 1279.8000 1302.4501 ;
	    RECT 1276.2001 1301.4000 1277.4000 1301.5500 ;
	    RECT 1278.6000 1301.4000 1279.8000 1301.5500 ;
	    RECT 1280.7001 1300.8000 1281.0000 1302.3000 ;
	    RECT 1283.1000 1301.4000 1284.9000 1302.6000 ;
	    RECT 1285.8000 1302.4501 1287.0000 1302.6000 ;
	    RECT 1297.8000 1302.4501 1299.0000 1302.6000 ;
	    RECT 1285.8000 1301.5500 1299.0000 1302.4501 ;
	    RECT 1285.8000 1301.4000 1287.0000 1301.5500 ;
	    RECT 1297.8000 1301.4000 1299.0000 1301.5500 ;
	    RECT 1302.6000 1302.4501 1303.8000 1302.6000 ;
	    RECT 1324.3500 1302.4501 1325.2500 1304.5500 ;
	    RECT 1329.0000 1304.4000 1330.2001 1304.5500 ;
	    RECT 1329.0000 1303.2001 1330.2001 1303.5000 ;
	    RECT 1331.1000 1302.6000 1332.0000 1307.7001 ;
	    RECT 1333.8000 1308.4501 1335.0000 1308.6000 ;
	    RECT 1350.6000 1308.4501 1351.8000 1308.6000 ;
	    RECT 1333.8000 1307.5500 1351.8000 1308.4501 ;
	    RECT 1333.8000 1307.4000 1335.0000 1307.5500 ;
	    RECT 1350.6000 1307.4000 1351.8000 1307.5500 ;
	    RECT 1465.8000 1303.5000 1467.0000 1311.9000 ;
	    RECT 1469.7001 1311.6000 1476.0000 1312.8000 ;
	    RECT 1482.6000 1312.5000 1483.8000 1319.7001 ;
	    RECT 1485.0000 1313.7001 1486.2001 1319.7001 ;
	    RECT 1487.4000 1312.5000 1488.6000 1319.7001 ;
	    RECT 1489.8000 1313.7001 1491.0000 1319.7001 ;
	    RECT 1469.7001 1311.0000 1470.6000 1311.6000 ;
	    RECT 1468.2001 1309.8000 1470.6000 1311.0000 ;
	    RECT 1475.1000 1310.7001 1483.8000 1311.6000 ;
	    RECT 1472.1000 1309.8000 1474.2001 1310.7001 ;
	    RECT 1472.1000 1309.5000 1481.4000 1309.8000 ;
	    RECT 1473.3000 1308.9000 1481.4000 1309.5000 ;
	    RECT 1480.2001 1308.6000 1481.4000 1308.9000 ;
	    RECT 1482.9000 1309.5000 1483.8000 1310.7001 ;
	    RECT 1484.7001 1310.4000 1488.6000 1311.6000 ;
	    RECT 1492.2001 1310.4000 1493.4000 1319.7001 ;
	    RECT 1494.6000 1315.5000 1495.8000 1319.7001 ;
	    RECT 1497.0000 1315.5000 1498.2001 1319.7001 ;
	    RECT 1499.4000 1315.5000 1500.6000 1319.7001 ;
	    RECT 1501.8000 1313.7001 1503.0000 1319.7001 ;
	    RECT 1497.0000 1311.6000 1503.3000 1312.8000 ;
	    RECT 1504.2001 1311.6000 1505.4000 1319.7001 ;
	    RECT 1506.6000 1313.7001 1507.8000 1319.7001 ;
	    RECT 1509.0000 1312.8000 1510.2001 1319.7001 ;
	    RECT 1511.4000 1313.7001 1512.6000 1319.7001 ;
	    RECT 1509.0000 1311.9000 1512.9000 1312.8000 ;
	    RECT 1513.8000 1312.5000 1515.0000 1319.7001 ;
	    RECT 1516.2001 1313.7001 1517.4000 1319.7001 ;
	    RECT 1504.2001 1310.4000 1508.1000 1311.6000 ;
	    RECT 1494.6000 1309.5000 1495.8000 1309.8000 ;
	    RECT 1482.9000 1308.6000 1495.8000 1309.5000 ;
	    RECT 1499.4000 1309.5000 1500.6000 1309.8000 ;
	    RECT 1512.0000 1309.5000 1512.9000 1311.9000 ;
	    RECT 1513.8000 1310.4000 1515.0000 1311.6000 ;
	    RECT 1499.4000 1308.6000 1512.9000 1309.5000 ;
	    RECT 1470.6000 1307.4000 1471.8000 1308.6000 ;
	    RECT 1475.7001 1307.7001 1476.9000 1308.0000 ;
	    RECT 1472.7001 1306.8000 1511.1000 1307.7001 ;
	    RECT 1509.9000 1306.5000 1511.1000 1306.8000 ;
	    RECT 1512.0000 1305.9000 1512.9000 1308.6000 ;
	    RECT 1513.8000 1308.0000 1515.0000 1309.5000 ;
	    RECT 1535.4000 1308.6000 1536.6000 1319.7001 ;
	    RECT 1537.8000 1309.5000 1539.0000 1319.7001 ;
	    RECT 1513.8000 1306.8000 1515.3000 1308.0000 ;
	    RECT 1535.4000 1307.7001 1538.7001 1308.6000 ;
	    RECT 1540.2001 1307.7001 1541.4000 1319.7001 ;
	    RECT 1547.4000 1319.4000 1548.6000 1320.6000 ;
	    RECT 1552.2001 1313.7001 1553.4000 1319.7001 ;
	    RECT 1467.9000 1305.0000 1474.5000 1305.9000 ;
	    RECT 1467.9000 1304.7001 1469.1000 1305.0000 ;
	    RECT 1475.4000 1304.4000 1476.6000 1305.6000 ;
	    RECT 1477.5000 1305.0000 1503.0000 1305.9000 ;
	    RECT 1512.0000 1305.0000 1513.2001 1305.9000 ;
	    RECT 1501.8000 1304.1000 1503.0000 1305.0000 ;
	    RECT 1302.6000 1301.5500 1325.2500 1302.4501 ;
	    RECT 1302.6000 1301.4000 1303.8000 1301.5500 ;
	    RECT 1326.6000 1301.4000 1327.8000 1302.6000 ;
	    RECT 1328.7001 1300.8000 1329.0000 1302.3000 ;
	    RECT 1331.1000 1301.4000 1332.9000 1302.6000 ;
	    RECT 1333.8000 1302.4501 1335.0000 1302.6000 ;
	    RECT 1463.4000 1302.4501 1464.6000 1302.6000 ;
	    RECT 1333.8000 1301.5500 1464.6000 1302.4501 ;
	    RECT 1333.8000 1301.4000 1335.0000 1301.5500 ;
	    RECT 1463.4000 1301.4000 1464.6000 1301.5500 ;
	    RECT 1465.8000 1302.3000 1479.0000 1303.5000 ;
	    RECT 1479.9000 1302.9000 1482.9000 1304.1000 ;
	    RECT 1488.6000 1302.9000 1493.4000 1304.1000 ;
	    RECT 1278.9000 1299.3000 1284.3000 1299.9000 ;
	    RECT 1285.8000 1299.3000 1286.7001 1300.5000 ;
	    RECT 1249.8000 1293.3000 1251.0000 1299.3000 ;
	    RECT 1252.2001 1298.4000 1254.9000 1299.3000 ;
	    RECT 1253.7001 1293.3000 1254.9000 1298.4000 ;
	    RECT 1278.6000 1299.0000 1284.6000 1299.3000 ;
	    RECT 1278.6000 1293.3000 1279.8000 1299.0000 ;
	    RECT 1281.0000 1293.3000 1282.2001 1298.1000 ;
	    RECT 1283.4000 1293.3000 1284.6000 1299.0000 ;
	    RECT 1285.8000 1293.3000 1287.0000 1299.3000 ;
	    RECT 1300.2001 1298.4000 1301.4000 1299.6000 ;
	    RECT 1300.2001 1297.2001 1301.4000 1297.5000 ;
	    RECT 1300.2001 1293.3000 1301.4000 1296.3000 ;
	    RECT 1302.6000 1293.3000 1303.8000 1300.5000 ;
	    RECT 1326.9000 1299.3000 1332.3000 1299.9000 ;
	    RECT 1333.8000 1299.3000 1334.7001 1300.5000 ;
	    RECT 1326.6000 1299.0000 1332.6000 1299.3000 ;
	    RECT 1326.6000 1293.3000 1327.8000 1299.0000 ;
	    RECT 1329.0000 1293.3000 1330.2001 1298.1000 ;
	    RECT 1331.4000 1293.3000 1332.6000 1299.0000 ;
	    RECT 1333.8000 1293.3000 1335.0000 1299.3000 ;
	    RECT 1465.8000 1293.3000 1467.0000 1302.3000 ;
	    RECT 1469.4000 1300.2001 1473.9000 1301.4000 ;
	    RECT 1472.7001 1299.3000 1473.9000 1300.2001 ;
	    RECT 1481.7001 1299.3000 1482.9000 1302.9000 ;
	    RECT 1485.0000 1301.4000 1486.2001 1302.6000 ;
	    RECT 1492.8000 1301.7001 1494.0000 1302.0000 ;
	    RECT 1487.4000 1300.8000 1494.0000 1301.7001 ;
	    RECT 1487.4000 1300.5000 1488.6000 1300.8000 ;
	    RECT 1485.0000 1300.2001 1486.2001 1300.5000 ;
	    RECT 1497.0000 1299.6000 1498.2001 1303.8000 ;
	    RECT 1505.7001 1302.9000 1511.4000 1304.1000 ;
	    RECT 1505.7001 1301.1000 1506.9000 1302.9000 ;
	    RECT 1512.3000 1302.0000 1513.2001 1305.0000 ;
	    RECT 1487.4000 1299.3000 1488.6000 1299.6000 ;
	    RECT 1470.6000 1293.3000 1471.8000 1299.3000 ;
	    RECT 1472.7001 1298.1000 1476.6000 1299.3000 ;
	    RECT 1481.7001 1298.4000 1488.6000 1299.3000 ;
	    RECT 1489.8000 1298.4000 1491.0000 1299.6000 ;
	    RECT 1491.9000 1298.4000 1492.2001 1299.6000 ;
	    RECT 1496.7001 1298.4000 1498.2001 1299.6000 ;
	    RECT 1504.2001 1300.2001 1506.9000 1301.1000 ;
	    RECT 1511.4000 1301.1000 1513.2001 1302.0000 ;
	    RECT 1504.2001 1299.3000 1505.4000 1300.2001 ;
	    RECT 1475.4000 1293.3000 1476.6000 1298.1000 ;
	    RECT 1501.8000 1298.1000 1505.4000 1299.3000 ;
	    RECT 1477.8000 1293.3000 1479.0000 1297.5000 ;
	    RECT 1480.2001 1293.3000 1481.4000 1297.5000 ;
	    RECT 1482.6000 1293.3000 1483.8000 1297.5000 ;
	    RECT 1485.0000 1293.3000 1486.2001 1296.3000 ;
	    RECT 1487.4000 1293.3000 1488.6000 1297.5000 ;
	    RECT 1489.8000 1293.3000 1491.0000 1296.3000 ;
	    RECT 1492.2001 1293.3000 1493.4000 1297.5000 ;
	    RECT 1494.6000 1293.3000 1495.8000 1297.5000 ;
	    RECT 1497.0000 1293.3000 1498.2001 1297.5000 ;
	    RECT 1499.4000 1293.3000 1500.6000 1297.5000 ;
	    RECT 1501.8000 1293.3000 1503.0000 1298.1000 ;
	    RECT 1506.6000 1293.3000 1507.8000 1299.3000 ;
	    RECT 1511.4000 1293.3000 1512.6000 1301.1000 ;
	    RECT 1514.1000 1300.2001 1515.3000 1306.8000 ;
	    RECT 1537.8000 1306.8000 1538.7001 1307.7001 ;
	    RECT 1537.8000 1305.6000 1539.6000 1306.8000 ;
	    RECT 1516.2001 1305.4501 1517.4000 1305.6000 ;
	    RECT 1535.4000 1305.4501 1536.6000 1305.6000 ;
	    RECT 1516.2001 1304.5500 1536.6000 1305.4501 ;
	    RECT 1516.2001 1304.4000 1517.4000 1304.5500 ;
	    RECT 1535.4000 1304.4000 1536.6000 1304.5500 ;
	    RECT 1535.4000 1303.2001 1536.6000 1303.5000 ;
	    RECT 1537.8000 1301.1000 1538.7001 1305.6000 ;
	    RECT 1540.5000 1304.4000 1541.4000 1307.7001 ;
	    RECT 1540.2001 1303.5000 1541.4000 1304.4000 ;
	    RECT 1554.6000 1303.5000 1555.8000 1319.7001 ;
	    RECT 1554.6000 1301.4000 1555.8000 1302.6000 ;
	    RECT 1513.8000 1299.0000 1515.3000 1300.2001 ;
	    RECT 1535.4000 1300.2001 1538.7001 1301.1000 ;
	    RECT 1513.8000 1293.3000 1515.0000 1299.0000 ;
	    RECT 1516.2001 1293.3000 1517.4000 1296.3000 ;
	    RECT 1535.4000 1293.3000 1536.6000 1300.2001 ;
	    RECT 1537.8000 1293.3000 1539.0000 1299.3000 ;
	    RECT 1540.2001 1293.3000 1541.4000 1300.5000 ;
	    RECT 1552.2001 1298.4000 1553.4000 1299.6000 ;
	    RECT 1552.2001 1297.2001 1553.4000 1297.5000 ;
	    RECT 1552.2001 1293.3000 1553.4000 1296.3000 ;
	    RECT 1554.6000 1293.3000 1555.8000 1300.5000 ;
	    RECT 1.2000 1290.6000 1569.0000 1292.4000 ;
	    RECT 25.8000 1284.0000 27.0000 1289.7001 ;
	    RECT 28.2000 1284.9000 29.4000 1289.7001 ;
	    RECT 30.6000 1284.0000 31.8000 1289.7001 ;
	    RECT 25.8000 1283.7001 31.8000 1284.0000 ;
	    RECT 33.0000 1283.7001 34.2000 1289.7001 ;
	    RECT 26.1000 1283.1000 31.5000 1283.7001 ;
	    RECT 33.0000 1282.5000 33.9000 1283.7001 ;
	    RECT 45.0000 1282.5000 46.2000 1289.7001 ;
	    RECT 47.4000 1286.7001 48.6000 1289.7001 ;
	    RECT 47.4000 1285.5000 48.6000 1285.8000 ;
	    RECT 47.4000 1284.4501 48.6000 1284.6000 ;
	    RECT 57.0000 1284.4501 58.2000 1284.6000 ;
	    RECT 47.4000 1283.5500 58.2000 1284.4501 ;
	    RECT 47.4000 1283.4000 48.6000 1283.5500 ;
	    RECT 57.0000 1283.4000 58.2000 1283.5500 ;
	    RECT 59.4000 1282.5000 60.6000 1289.7001 ;
	    RECT 61.8000 1286.7001 63.0000 1289.7001 ;
	    RECT 61.8000 1285.5000 63.0000 1285.8000 ;
	    RECT 61.8000 1284.4501 63.0000 1284.6000 ;
	    RECT 76.2000 1284.4501 77.4000 1284.6000 ;
	    RECT 61.8000 1283.5500 77.4000 1284.4501 ;
	    RECT 85.8000 1283.7001 87.0000 1289.7001 ;
	    RECT 88.2000 1284.0000 89.4000 1289.7001 ;
	    RECT 90.6000 1284.9000 91.8000 1289.7001 ;
	    RECT 93.0000 1284.0000 94.2000 1289.7001 ;
	    RECT 88.2000 1283.7001 94.2000 1284.0000 ;
	    RECT 112.2000 1283.7001 113.4000 1289.7001 ;
	    RECT 116.1000 1284.6000 117.3000 1289.7001 ;
	    RECT 249.0000 1286.7001 250.2000 1289.7001 ;
	    RECT 114.6000 1283.7001 117.3000 1284.6000 ;
	    RECT 251.4000 1284.0000 252.6000 1289.7001 ;
	    RECT 61.8000 1283.4000 63.0000 1283.5500 ;
	    RECT 76.2000 1283.4000 77.4000 1283.5500 ;
	    RECT 86.1000 1282.5000 87.0000 1283.7001 ;
	    RECT 88.5000 1283.1000 93.9000 1283.7001 ;
	    RECT 112.2000 1282.5000 113.4000 1282.8000 ;
	    RECT 18.6000 1281.4501 19.8000 1281.6000 ;
	    RECT 25.8000 1281.4501 27.0000 1281.6000 ;
	    RECT 18.6000 1280.5500 27.0000 1281.4501 ;
	    RECT 27.9000 1280.7001 28.2000 1282.2001 ;
	    RECT 18.6000 1280.4000 19.8000 1280.5500 ;
	    RECT 25.8000 1280.4000 27.0000 1280.5500 ;
	    RECT 30.3000 1280.4000 32.1000 1281.6000 ;
	    RECT 33.0000 1280.4000 34.2000 1281.6000 ;
	    RECT 35.4000 1281.4501 36.6000 1281.6000 ;
	    RECT 45.0000 1281.4501 46.2000 1281.6000 ;
	    RECT 35.4000 1280.5500 46.2000 1281.4501 ;
	    RECT 35.4000 1280.4000 36.6000 1280.5500 ;
	    RECT 45.0000 1280.4000 46.2000 1280.5500 ;
	    RECT 54.6000 1281.4501 55.8000 1281.6000 ;
	    RECT 59.4000 1281.4501 60.6000 1281.6000 ;
	    RECT 54.6000 1280.5500 60.6000 1281.4501 ;
	    RECT 54.6000 1280.4000 55.8000 1280.5500 ;
	    RECT 59.4000 1280.4000 60.6000 1280.5500 ;
	    RECT 83.4000 1281.4501 84.6000 1281.6000 ;
	    RECT 85.8000 1281.4501 87.0000 1281.6000 ;
	    RECT 83.4000 1280.5500 87.0000 1281.4501 ;
	    RECT 83.4000 1280.4000 84.6000 1280.5500 ;
	    RECT 85.8000 1280.4000 87.0000 1280.5500 ;
	    RECT 87.9000 1280.4000 89.7000 1281.6000 ;
	    RECT 91.8000 1280.7001 92.1000 1282.2001 ;
	    RECT 93.0000 1281.4501 94.2000 1281.6000 ;
	    RECT 107.4000 1281.4501 108.6000 1281.6000 ;
	    RECT 112.2000 1281.4501 113.4000 1281.6000 ;
	    RECT 93.0000 1280.5500 113.4000 1281.4501 ;
	    RECT 93.0000 1280.4000 94.2000 1280.5500 ;
	    RECT 107.4000 1280.4000 108.6000 1280.5500 ;
	    RECT 112.2000 1280.4000 113.4000 1280.5500 ;
	    RECT 28.2000 1279.5000 29.4000 1279.8000 ;
	    RECT 28.2000 1277.4000 29.4000 1278.6000 ;
	    RECT 30.3000 1275.3000 31.2000 1280.4000 ;
	    RECT 25.8000 1263.3000 27.0000 1275.3000 ;
	    RECT 29.7000 1274.4000 31.2000 1275.3000 ;
	    RECT 33.0000 1275.4501 34.2000 1275.6000 ;
	    RECT 35.4000 1275.4501 36.6000 1275.6000 ;
	    RECT 33.0000 1274.5500 36.6000 1275.4501 ;
	    RECT 33.0000 1274.4000 34.2000 1274.5500 ;
	    RECT 35.4000 1274.4000 36.6000 1274.5500 ;
	    RECT 29.7000 1263.3000 30.9000 1274.4000 ;
	    RECT 32.1000 1272.6000 33.0000 1273.5000 ;
	    RECT 31.8000 1271.4000 33.0000 1272.6000 ;
	    RECT 32.1000 1263.3000 33.3000 1269.3000 ;
	    RECT 45.0000 1263.3000 46.2000 1279.5000 ;
	    RECT 47.4000 1263.3000 48.6000 1269.3000 ;
	    RECT 59.4000 1263.3000 60.6000 1279.5000 ;
	    RECT 85.8000 1274.4000 87.0000 1275.6000 ;
	    RECT 88.8000 1275.3000 89.7000 1280.4000 ;
	    RECT 90.6000 1279.5000 91.8000 1279.8000 ;
	    RECT 114.6000 1279.5000 115.8000 1283.7001 ;
	    RECT 251.1000 1282.8000 252.6000 1284.0000 ;
	    RECT 90.6000 1278.4501 91.8000 1278.6000 ;
	    RECT 93.0000 1278.4501 94.2000 1278.6000 ;
	    RECT 90.6000 1277.5500 94.2000 1278.4501 ;
	    RECT 90.6000 1277.4000 91.8000 1277.5500 ;
	    RECT 93.0000 1277.4000 94.2000 1277.5500 ;
	    RECT 95.4000 1278.4501 96.6000 1278.6000 ;
	    RECT 114.6000 1278.4501 115.8000 1278.6000 ;
	    RECT 95.4000 1277.5500 115.8000 1278.4501 ;
	    RECT 95.4000 1277.4000 96.6000 1277.5500 ;
	    RECT 114.6000 1277.4000 115.8000 1277.5500 ;
	    RECT 88.8000 1274.4000 90.3000 1275.3000 ;
	    RECT 87.0000 1272.6000 87.9000 1273.5000 ;
	    RECT 87.0000 1271.4000 88.2000 1272.6000 ;
	    RECT 61.8000 1263.3000 63.0000 1269.3000 ;
	    RECT 86.7000 1263.3000 87.9000 1269.3000 ;
	    RECT 89.1000 1263.3000 90.3000 1274.4000 ;
	    RECT 93.0000 1263.3000 94.2000 1275.3000 ;
	    RECT 112.2000 1263.3000 113.4000 1269.3000 ;
	    RECT 114.6000 1263.3000 115.8000 1276.5000 ;
	    RECT 251.1000 1276.2001 252.3000 1282.8000 ;
	    RECT 253.8000 1281.9000 255.0000 1289.7001 ;
	    RECT 258.6000 1283.7001 259.8000 1289.7001 ;
	    RECT 263.4000 1284.9000 264.6000 1289.7001 ;
	    RECT 265.8000 1285.5000 267.0000 1289.7001 ;
	    RECT 268.2000 1285.5000 269.4000 1289.7001 ;
	    RECT 270.6000 1285.5000 271.8000 1289.7001 ;
	    RECT 273.0000 1285.5000 274.2000 1289.7001 ;
	    RECT 275.4000 1286.7001 276.6000 1289.7001 ;
	    RECT 277.8000 1285.5000 279.0000 1289.7001 ;
	    RECT 280.2000 1286.7001 281.4000 1289.7001 ;
	    RECT 282.6000 1285.5000 283.8000 1289.7001 ;
	    RECT 285.0000 1285.5000 286.2000 1289.7001 ;
	    RECT 287.4000 1285.5000 288.6000 1289.7001 ;
	    RECT 261.0000 1283.7001 264.6000 1284.9000 ;
	    RECT 289.8000 1284.9000 291.0000 1289.7001 ;
	    RECT 261.0000 1282.8000 262.2000 1283.7001 ;
	    RECT 253.2000 1281.0000 255.0000 1281.9000 ;
	    RECT 259.5000 1281.9000 262.2000 1282.8000 ;
	    RECT 268.2000 1283.4000 269.7000 1284.6000 ;
	    RECT 274.2000 1283.4000 274.5000 1284.6000 ;
	    RECT 275.4000 1283.4000 276.6000 1284.6000 ;
	    RECT 277.8000 1283.7001 284.7000 1284.6000 ;
	    RECT 289.8000 1283.7001 293.7000 1284.9000 ;
	    RECT 294.6000 1283.7001 295.8000 1289.7001 ;
	    RECT 277.8000 1283.4000 279.0000 1283.7001 ;
	    RECT 253.2000 1278.0000 254.1000 1281.0000 ;
	    RECT 259.5000 1280.1000 260.7000 1281.9000 ;
	    RECT 255.0000 1278.9000 260.7000 1280.1000 ;
	    RECT 268.2000 1279.2001 269.4000 1283.4000 ;
	    RECT 280.2000 1282.5000 281.4000 1282.8000 ;
	    RECT 277.8000 1282.2001 279.0000 1282.5000 ;
	    RECT 272.4000 1281.3000 279.0000 1282.2001 ;
	    RECT 272.4000 1281.0000 273.6000 1281.3000 ;
	    RECT 280.2000 1280.4000 281.4000 1281.6000 ;
	    RECT 283.5000 1280.1000 284.7000 1283.7001 ;
	    RECT 292.5000 1282.8000 293.7000 1283.7001 ;
	    RECT 292.5000 1281.6000 297.0000 1282.8000 ;
	    RECT 299.4000 1280.7001 300.6000 1289.7001 ;
	    RECT 311.4000 1286.7001 312.6000 1289.7001 ;
	    RECT 311.4000 1285.5000 312.6000 1285.8000 ;
	    RECT 311.4000 1283.4000 312.6000 1284.6000 ;
	    RECT 313.8000 1282.5000 315.0000 1289.7001 ;
	    RECT 325.8000 1282.5000 327.0000 1289.7001 ;
	    RECT 328.2000 1286.7001 329.4000 1289.7001 ;
	    RECT 328.2000 1285.5000 329.4000 1285.8000 ;
	    RECT 328.2000 1283.4000 329.4000 1284.6000 ;
	    RECT 354.6000 1283.7001 355.8000 1289.7001 ;
	    RECT 357.0000 1284.0000 358.2000 1289.7001 ;
	    RECT 359.4000 1284.9000 360.6000 1289.7001 ;
	    RECT 361.8000 1284.0000 363.0000 1289.7001 ;
	    RECT 357.0000 1283.7001 363.0000 1284.0000 ;
	    RECT 385.8000 1284.0000 387.0000 1289.7001 ;
	    RECT 388.2000 1284.9000 389.4000 1289.7001 ;
	    RECT 390.6000 1284.0000 391.8000 1289.7001 ;
	    RECT 385.8000 1283.7001 391.8000 1284.0000 ;
	    RECT 393.0000 1283.7001 394.2000 1289.7001 ;
	    RECT 354.9000 1282.5000 355.8000 1283.7001 ;
	    RECT 357.3000 1283.1000 362.7000 1283.7001 ;
	    RECT 386.1000 1283.1000 391.5000 1283.7001 ;
	    RECT 393.0000 1282.5000 393.9000 1283.7001 ;
	    RECT 407.4000 1282.5000 408.6000 1289.7001 ;
	    RECT 409.8000 1286.7001 411.0000 1289.7001 ;
	    RECT 409.8000 1285.5000 411.0000 1285.8000 ;
	    RECT 429.9000 1284.6000 431.1000 1289.7001 ;
	    RECT 409.8000 1284.4501 411.0000 1284.6000 ;
	    RECT 414.6000 1284.4501 415.8000 1284.6000 ;
	    RECT 409.8000 1283.5500 415.8000 1284.4501 ;
	    RECT 429.9000 1283.7001 432.6000 1284.6000 ;
	    RECT 433.8000 1283.7001 435.0000 1289.7001 ;
	    RECT 465.0000 1284.0000 466.2000 1289.7001 ;
	    RECT 467.4000 1284.9000 468.6000 1289.7001 ;
	    RECT 469.8000 1284.0000 471.0000 1289.7001 ;
	    RECT 465.0000 1283.7001 471.0000 1284.0000 ;
	    RECT 472.2000 1283.7001 473.4000 1289.7001 ;
	    RECT 409.8000 1283.4000 411.0000 1283.5500 ;
	    RECT 414.6000 1283.4000 415.8000 1283.5500 ;
	    RECT 273.0000 1278.9000 277.8000 1280.1000 ;
	    RECT 283.5000 1278.9000 286.5000 1280.1000 ;
	    RECT 287.4000 1279.5000 300.6000 1280.7001 ;
	    RECT 313.8000 1281.4501 315.0000 1281.6000 ;
	    RECT 323.4000 1281.4501 324.6000 1281.6000 ;
	    RECT 313.8000 1280.5500 324.6000 1281.4501 ;
	    RECT 313.8000 1280.4000 315.0000 1280.5500 ;
	    RECT 323.4000 1280.4000 324.6000 1280.5500 ;
	    RECT 325.8000 1280.4000 327.0000 1281.6000 ;
	    RECT 354.6000 1280.4000 355.8000 1281.6000 ;
	    RECT 356.7000 1280.4000 358.5000 1281.6000 ;
	    RECT 360.6000 1280.7001 360.9000 1282.2001 ;
	    RECT 361.8000 1281.4501 363.0000 1281.6000 ;
	    RECT 383.4000 1281.4501 384.6000 1281.6000 ;
	    RECT 385.8000 1281.4501 387.0000 1281.6000 ;
	    RECT 361.8000 1280.5500 387.0000 1281.4501 ;
	    RECT 387.9000 1280.7001 388.2000 1282.2001 ;
	    RECT 361.8000 1280.4000 363.0000 1280.5500 ;
	    RECT 383.4000 1280.4000 384.6000 1280.5500 ;
	    RECT 385.8000 1280.4000 387.0000 1280.5500 ;
	    RECT 390.3000 1280.4000 392.1000 1281.6000 ;
	    RECT 393.0000 1281.4501 394.2000 1281.6000 ;
	    RECT 405.0000 1281.4501 406.2000 1281.6000 ;
	    RECT 393.0000 1280.5500 406.2000 1281.4501 ;
	    RECT 393.0000 1280.4000 394.2000 1280.5500 ;
	    RECT 405.0000 1280.4000 406.2000 1280.5500 ;
	    RECT 407.4000 1281.4501 408.6000 1281.6000 ;
	    RECT 412.2000 1281.4501 413.4000 1281.6000 ;
	    RECT 407.4000 1280.5500 413.4000 1281.4501 ;
	    RECT 407.4000 1280.4000 408.6000 1280.5500 ;
	    RECT 412.2000 1280.4000 413.4000 1280.5500 ;
	    RECT 263.4000 1278.0000 264.6000 1278.9000 ;
	    RECT 253.2000 1277.1000 254.4000 1278.0000 ;
	    RECT 263.4000 1277.1000 288.9000 1278.0000 ;
	    RECT 289.8000 1277.4000 291.0000 1278.6000 ;
	    RECT 297.3000 1278.0000 298.5000 1278.3000 ;
	    RECT 291.9000 1277.1000 298.5000 1278.0000 ;
	    RECT 117.0000 1275.4501 118.2000 1275.6000 ;
	    RECT 196.2000 1275.4501 197.4000 1275.6000 ;
	    RECT 117.0000 1274.5500 197.4000 1275.4501 ;
	    RECT 251.1000 1275.0000 252.6000 1276.2001 ;
	    RECT 117.0000 1274.4000 118.2000 1274.5500 ;
	    RECT 196.2000 1274.4000 197.4000 1274.5500 ;
	    RECT 251.4000 1273.5000 252.6000 1275.0000 ;
	    RECT 253.5000 1274.4000 254.4000 1277.1000 ;
	    RECT 255.3000 1276.2001 256.5000 1276.5000 ;
	    RECT 255.3000 1275.3000 293.7000 1276.2001 ;
	    RECT 289.5000 1275.0000 290.7000 1275.3000 ;
	    RECT 294.6000 1274.4000 295.8000 1275.6000 ;
	    RECT 253.5000 1273.5000 267.0000 1274.4000 ;
	    RECT 117.0000 1273.2001 118.2000 1273.5000 ;
	    RECT 196.2000 1272.4501 197.4000 1272.6000 ;
	    RECT 213.0000 1272.4501 214.2000 1272.6000 ;
	    RECT 251.4000 1272.4501 252.6000 1272.6000 ;
	    RECT 196.2000 1271.5500 252.6000 1272.4501 ;
	    RECT 196.2000 1271.4000 197.4000 1271.5500 ;
	    RECT 213.0000 1271.4000 214.2000 1271.5500 ;
	    RECT 251.4000 1271.4000 252.6000 1271.5500 ;
	    RECT 253.5000 1271.1000 254.4000 1273.5000 ;
	    RECT 265.8000 1273.2001 267.0000 1273.5000 ;
	    RECT 270.6000 1273.5000 283.5000 1274.4000 ;
	    RECT 270.6000 1273.2001 271.8000 1273.5000 ;
	    RECT 258.3000 1271.4000 262.2000 1272.6000 ;
	    RECT 117.0000 1263.3000 118.2000 1269.3000 ;
	    RECT 249.0000 1263.3000 250.2000 1269.3000 ;
	    RECT 251.4000 1263.3000 252.6000 1270.5000 ;
	    RECT 253.5000 1270.2001 257.4000 1271.1000 ;
	    RECT 253.8000 1263.3000 255.0000 1269.3000 ;
	    RECT 256.2000 1263.3000 257.4000 1270.2001 ;
	    RECT 258.6000 1263.3000 259.8000 1269.3000 ;
	    RECT 261.0000 1263.3000 262.2000 1271.4000 ;
	    RECT 263.1000 1270.2001 269.4000 1271.4000 ;
	    RECT 263.4000 1263.3000 264.6000 1269.3000 ;
	    RECT 265.8000 1263.3000 267.0000 1267.5000 ;
	    RECT 268.2000 1263.3000 269.4000 1267.5000 ;
	    RECT 270.6000 1263.3000 271.8000 1267.5000 ;
	    RECT 273.0000 1263.3000 274.2000 1272.6000 ;
	    RECT 277.8000 1271.4000 281.7000 1272.6000 ;
	    RECT 282.6000 1272.3000 283.5000 1273.5000 ;
	    RECT 285.0000 1274.1000 286.2000 1274.4000 ;
	    RECT 285.0000 1273.5000 293.1000 1274.1000 ;
	    RECT 285.0000 1273.2001 294.3000 1273.5000 ;
	    RECT 292.2000 1272.3000 294.3000 1273.2001 ;
	    RECT 282.6000 1271.4000 291.3000 1272.3000 ;
	    RECT 295.8000 1272.0000 298.2000 1273.2001 ;
	    RECT 295.8000 1271.4000 296.7000 1272.0000 ;
	    RECT 275.4000 1263.3000 276.6000 1269.3000 ;
	    RECT 277.8000 1263.3000 279.0000 1270.5000 ;
	    RECT 280.2000 1263.3000 281.4000 1269.3000 ;
	    RECT 282.6000 1263.3000 283.8000 1270.5000 ;
	    RECT 290.4000 1270.2001 296.7000 1271.4000 ;
	    RECT 299.4000 1271.1000 300.6000 1279.5000 ;
	    RECT 297.6000 1270.2001 300.6000 1271.1000 ;
	    RECT 285.0000 1263.3000 286.2000 1267.5000 ;
	    RECT 287.4000 1263.3000 288.6000 1267.5000 ;
	    RECT 289.8000 1263.3000 291.0000 1269.3000 ;
	    RECT 292.2000 1263.3000 293.4000 1270.2001 ;
	    RECT 297.6000 1269.3000 298.5000 1270.2001 ;
	    RECT 294.6000 1262.4000 295.8000 1269.3000 ;
	    RECT 297.0000 1268.4000 298.5000 1269.3000 ;
	    RECT 297.0000 1263.3000 298.2000 1268.4000 ;
	    RECT 299.4000 1263.3000 300.6000 1269.3000 ;
	    RECT 311.4000 1263.3000 312.6000 1269.3000 ;
	    RECT 313.8000 1263.3000 315.0000 1279.5000 ;
	    RECT 325.8000 1263.3000 327.0000 1279.5000 ;
	    RECT 337.8000 1275.4501 339.0000 1275.6000 ;
	    RECT 354.6000 1275.4501 355.8000 1275.6000 ;
	    RECT 337.8000 1274.5500 355.8000 1275.4501 ;
	    RECT 337.8000 1274.4000 339.0000 1274.5500 ;
	    RECT 354.6000 1274.4000 355.8000 1274.5500 ;
	    RECT 357.6000 1275.3000 358.5000 1280.4000 ;
	    RECT 359.4000 1279.5000 360.6000 1279.8000 ;
	    RECT 388.2000 1279.5000 389.4000 1279.8000 ;
	    RECT 359.4000 1277.4000 360.6000 1278.6000 ;
	    RECT 378.6000 1278.4501 379.8000 1278.6000 ;
	    RECT 388.2000 1278.4501 389.4000 1278.6000 ;
	    RECT 378.6000 1277.5500 389.4000 1278.4501 ;
	    RECT 378.6000 1277.4000 379.8000 1277.5500 ;
	    RECT 388.2000 1277.4000 389.4000 1277.5500 ;
	    RECT 390.3000 1275.3000 391.2000 1280.4000 ;
	    RECT 431.4000 1279.5000 432.6000 1283.7001 ;
	    RECT 465.3000 1283.1000 470.7000 1283.7001 ;
	    RECT 433.8000 1282.5000 435.0000 1282.8000 ;
	    RECT 472.2000 1282.5000 473.1000 1283.7001 ;
	    RECT 541.8000 1283.1000 543.0000 1289.7001 ;
	    RECT 544.2000 1284.0000 545.4000 1289.7001 ;
	    RECT 548.1000 1287.6000 549.9000 1289.7001 ;
	    RECT 548.1000 1286.7001 550.2000 1287.6000 ;
	    RECT 552.6000 1286.7001 553.8000 1289.7001 ;
	    RECT 555.0000 1286.7001 556.2000 1289.7001 ;
	    RECT 557.4000 1286.7001 558.9000 1289.7001 ;
	    RECT 561.6000 1287.6000 562.8000 1289.7001 ;
	    RECT 561.6000 1286.7001 564.6000 1287.6000 ;
	    RECT 549.0000 1285.5000 550.2000 1286.7001 ;
	    RECT 555.3000 1285.8000 556.2000 1286.7001 ;
	    RECT 555.3000 1284.9000 559.5000 1285.8000 ;
	    RECT 558.3000 1284.6000 559.5000 1284.9000 ;
	    RECT 561.0000 1284.6000 562.2000 1285.8000 ;
	    RECT 563.4000 1285.5000 564.6000 1286.7001 ;
	    RECT 546.3000 1283.1000 547.5000 1283.4000 ;
	    RECT 541.8000 1282.2001 547.5000 1283.1000 ;
	    RECT 433.8000 1281.4501 435.0000 1281.6000 ;
	    RECT 453.0000 1281.4501 454.2000 1281.6000 ;
	    RECT 433.8000 1280.5500 454.2000 1281.4501 ;
	    RECT 433.8000 1280.4000 435.0000 1280.5500 ;
	    RECT 453.0000 1280.4000 454.2000 1280.5500 ;
	    RECT 465.0000 1280.4000 466.2000 1281.6000 ;
	    RECT 467.1000 1280.7001 467.4000 1282.2001 ;
	    RECT 469.5000 1280.4000 471.3000 1281.6000 ;
	    RECT 472.2000 1281.4501 473.4000 1281.6000 ;
	    RECT 539.4000 1281.4501 540.6000 1281.6000 ;
	    RECT 472.2000 1280.5500 540.6000 1281.4501 ;
	    RECT 472.2000 1280.4000 473.4000 1280.5500 ;
	    RECT 539.4000 1280.4000 540.6000 1280.5500 ;
	    RECT 467.4000 1279.5000 468.6000 1279.8000 ;
	    RECT 357.6000 1274.4000 359.1000 1275.3000 ;
	    RECT 355.8000 1272.6000 356.7000 1273.5000 ;
	    RECT 355.8000 1271.4000 357.0000 1272.6000 ;
	    RECT 328.2000 1263.3000 329.4000 1269.3000 ;
	    RECT 355.5000 1263.3000 356.7000 1269.3000 ;
	    RECT 357.9000 1263.3000 359.1000 1274.4000 ;
	    RECT 361.8000 1263.3000 363.0000 1275.3000 ;
	    RECT 385.8000 1263.3000 387.0000 1275.3000 ;
	    RECT 389.7000 1274.4000 391.2000 1275.3000 ;
	    RECT 393.0000 1275.4501 394.2000 1275.6000 ;
	    RECT 395.4000 1275.4501 396.6000 1275.6000 ;
	    RECT 393.0000 1274.5500 396.6000 1275.4501 ;
	    RECT 393.0000 1274.4000 394.2000 1274.5500 ;
	    RECT 395.4000 1274.4000 396.6000 1274.5500 ;
	    RECT 389.7000 1263.3000 390.9000 1274.4000 ;
	    RECT 392.1000 1272.6000 393.0000 1273.5000 ;
	    RECT 391.8000 1271.4000 393.0000 1272.6000 ;
	    RECT 392.1000 1263.3000 393.3000 1269.3000 ;
	    RECT 407.4000 1263.3000 408.6000 1279.5000 ;
	    RECT 409.8000 1278.4501 411.0000 1278.6000 ;
	    RECT 431.4000 1278.4501 432.6000 1278.6000 ;
	    RECT 409.8000 1277.5500 432.6000 1278.4501 ;
	    RECT 409.8000 1277.4000 411.0000 1277.5500 ;
	    RECT 431.4000 1277.4000 432.6000 1277.5500 ;
	    RECT 467.4000 1277.4000 468.6000 1278.6000 ;
	    RECT 414.6000 1275.4501 415.8000 1275.6000 ;
	    RECT 429.0000 1275.4501 430.2000 1275.6000 ;
	    RECT 414.6000 1274.5500 430.2000 1275.4501 ;
	    RECT 414.6000 1274.4000 415.8000 1274.5500 ;
	    RECT 429.0000 1274.4000 430.2000 1274.5500 ;
	    RECT 429.0000 1273.2001 430.2000 1273.5000 ;
	    RECT 409.8000 1263.3000 411.0000 1269.3000 ;
	    RECT 429.0000 1263.3000 430.2000 1269.3000 ;
	    RECT 431.4000 1263.3000 432.6000 1276.5000 ;
	    RECT 469.5000 1275.3000 470.4000 1280.4000 ;
	    RECT 541.8000 1279.5000 543.0000 1282.2001 ;
	    RECT 552.3000 1281.3000 553.5000 1281.6000 ;
	    RECT 561.0000 1281.3000 561.9000 1284.6000 ;
	    RECT 565.8000 1283.7001 567.0000 1289.7001 ;
	    RECT 568.2000 1282.5000 569.4000 1289.7001 ;
	    RECT 580.2000 1286.7001 581.4000 1289.7001 ;
	    RECT 580.2000 1285.5000 581.4000 1285.8000 ;
	    RECT 580.2000 1283.4000 581.4000 1284.6000 ;
	    RECT 582.6000 1282.5000 583.8000 1289.7001 ;
	    RECT 609.0000 1284.0000 610.2000 1289.7001 ;
	    RECT 611.4000 1284.9000 612.6000 1289.7001 ;
	    RECT 613.8000 1284.0000 615.0000 1289.7001 ;
	    RECT 609.0000 1283.7001 615.0000 1284.0000 ;
	    RECT 616.2000 1283.7001 617.4000 1289.7001 ;
	    RECT 636.3000 1284.6000 637.5000 1289.7001 ;
	    RECT 636.3000 1283.7001 639.0000 1284.6000 ;
	    RECT 640.2000 1283.7001 641.4000 1289.7001 ;
	    RECT 652.2000 1286.7001 653.4000 1289.7001 ;
	    RECT 652.2000 1285.5000 653.4000 1285.8000 ;
	    RECT 642.6000 1284.4501 643.8000 1284.6000 ;
	    RECT 652.2000 1284.4501 653.4000 1284.6000 ;
	    RECT 609.3000 1283.1000 614.7000 1283.7001 ;
	    RECT 616.2000 1282.5000 617.1000 1283.7001 ;
	    RECT 551.7000 1280.4000 564.9000 1281.3000 ;
	    RECT 565.8000 1280.4000 567.0000 1281.6000 ;
	    RECT 567.9000 1280.4000 568.2000 1281.6000 ;
	    RECT 582.6000 1281.4501 583.8000 1281.6000 ;
	    RECT 582.6000 1280.5500 607.6500 1281.4501 ;
	    RECT 582.6000 1280.4000 583.8000 1280.5500 ;
	    RECT 549.0000 1279.2001 550.2000 1279.5000 ;
	    RECT 532.2000 1278.4501 533.4000 1278.6000 ;
	    RECT 541.8000 1278.4501 543.0000 1278.6000 ;
	    RECT 532.2000 1277.5500 543.0000 1278.4501 ;
	    RECT 544.5000 1278.3000 550.2000 1279.2001 ;
	    RECT 544.5000 1278.0000 545.7000 1278.3000 ;
	    RECT 532.2000 1277.4000 533.4000 1277.5500 ;
	    RECT 541.8000 1277.4000 543.0000 1277.5500 ;
	    RECT 546.9000 1277.1000 548.1000 1277.4000 ;
	    RECT 543.9000 1276.5000 548.1000 1277.1000 ;
	    RECT 541.8000 1276.2001 548.1000 1276.5000 ;
	    RECT 433.8000 1263.3000 435.0000 1269.3000 ;
	    RECT 465.0000 1263.3000 466.2000 1275.3000 ;
	    RECT 468.9000 1274.4000 470.4000 1275.3000 ;
	    RECT 472.2000 1274.4000 473.4000 1275.6000 ;
	    RECT 468.9000 1263.3000 470.1000 1274.4000 ;
	    RECT 471.3000 1272.6000 472.2000 1273.5000 ;
	    RECT 471.0000 1271.4000 472.2000 1272.6000 ;
	    RECT 471.3000 1263.3000 472.5000 1269.3000 ;
	    RECT 541.8000 1263.3000 543.0000 1276.2001 ;
	    RECT 551.7000 1275.6000 552.6000 1280.4000 ;
	    RECT 562.5000 1280.1000 563.7000 1280.4000 ;
	    RECT 564.9000 1278.6000 566.1000 1278.9000 ;
	    RECT 558.6000 1277.4000 559.8000 1278.6000 ;
	    RECT 560.7000 1277.7001 566.1000 1278.6000 ;
	    RECT 561.0000 1276.5000 569.4000 1276.8000 ;
	    RECT 560.7000 1276.2001 569.4000 1276.5000 ;
	    RECT 544.2000 1263.3000 545.4000 1275.3000 ;
	    RECT 549.0000 1274.7001 552.6000 1275.6000 ;
	    RECT 554.7000 1275.9000 569.4000 1276.2001 ;
	    RECT 554.7000 1275.3000 561.9000 1275.9000 ;
	    RECT 549.0000 1273.2001 549.9000 1274.7001 ;
	    RECT 547.8000 1272.0000 549.9000 1273.2001 ;
	    RECT 552.3000 1273.5000 553.5000 1273.8000 ;
	    RECT 554.7000 1273.5000 555.6000 1275.3000 ;
	    RECT 552.3000 1272.6000 555.6000 1273.5000 ;
	    RECT 556.5000 1273.5000 564.6000 1274.4000 ;
	    RECT 556.5000 1273.2001 557.7000 1273.5000 ;
	    RECT 563.4000 1273.2001 564.6000 1273.5000 ;
	    RECT 554.1000 1271.1000 555.3000 1271.4000 ;
	    RECT 558.3000 1271.1000 559.5000 1271.4000 ;
	    RECT 549.0000 1269.3000 550.2000 1270.5000 ;
	    RECT 554.1000 1270.2001 559.5000 1271.1000 ;
	    RECT 555.3000 1269.3000 556.2000 1270.2001 ;
	    RECT 563.4000 1269.3000 564.6000 1270.5000 ;
	    RECT 548.1000 1263.3000 549.9000 1269.3000 ;
	    RECT 552.6000 1263.3000 553.8000 1269.3000 ;
	    RECT 555.0000 1263.3000 556.2000 1269.3000 ;
	    RECT 557.4000 1263.3000 558.6000 1269.3000 ;
	    RECT 561.6000 1268.4000 564.6000 1269.3000 ;
	    RECT 561.6000 1263.3000 562.8000 1268.4000 ;
	    RECT 565.8000 1263.3000 567.0000 1275.0000 ;
	    RECT 568.2000 1263.3000 569.4000 1275.9000 ;
	    RECT 580.2000 1263.3000 581.4000 1269.3000 ;
	    RECT 582.6000 1263.3000 583.8000 1279.5000 ;
	    RECT 606.7500 1278.4501 607.6500 1280.5500 ;
	    RECT 609.0000 1280.4000 610.2000 1281.6000 ;
	    RECT 611.1000 1280.7001 611.4000 1282.2001 ;
	    RECT 613.5000 1280.4000 615.3000 1281.6000 ;
	    RECT 616.2000 1281.4501 617.4000 1281.6000 ;
	    RECT 635.4000 1281.4501 636.6000 1281.6000 ;
	    RECT 616.2000 1280.5500 636.6000 1281.4501 ;
	    RECT 616.2000 1280.4000 617.4000 1280.5500 ;
	    RECT 635.4000 1280.4000 636.6000 1280.5500 ;
	    RECT 611.4000 1279.5000 612.6000 1279.8000 ;
	    RECT 611.4000 1278.4501 612.6000 1278.6000 ;
	    RECT 606.7500 1277.5500 612.6000 1278.4501 ;
	    RECT 611.4000 1277.4000 612.6000 1277.5500 ;
	    RECT 613.5000 1275.3000 614.4000 1280.4000 ;
	    RECT 637.8000 1279.5000 639.0000 1283.7001 ;
	    RECT 642.6000 1283.5500 653.4000 1284.4501 ;
	    RECT 642.6000 1283.4000 643.8000 1283.5500 ;
	    RECT 652.2000 1283.4000 653.4000 1283.5500 ;
	    RECT 640.2000 1282.5000 641.4000 1282.8000 ;
	    RECT 654.6000 1282.5000 655.8000 1289.7001 ;
	    RECT 688.2000 1284.0000 689.4000 1289.7001 ;
	    RECT 690.6000 1284.9000 691.8000 1289.7001 ;
	    RECT 693.0000 1284.0000 694.2000 1289.7001 ;
	    RECT 688.2000 1283.7001 694.2000 1284.0000 ;
	    RECT 695.4000 1283.7001 696.6000 1289.7001 ;
	    RECT 721.8000 1284.0000 723.0000 1289.7001 ;
	    RECT 724.2000 1284.9000 725.4000 1289.7001 ;
	    RECT 726.6000 1284.0000 727.8000 1289.7001 ;
	    RECT 721.8000 1283.7001 727.8000 1284.0000 ;
	    RECT 729.0000 1283.7001 730.2000 1289.7001 ;
	    RECT 749.1000 1284.6000 750.3000 1289.7001 ;
	    RECT 749.1000 1283.7001 751.8000 1284.6000 ;
	    RECT 753.0000 1283.7001 754.2000 1289.7001 ;
	    RECT 810.6000 1284.4501 811.8000 1284.6000 ;
	    RECT 885.0000 1284.4501 886.2000 1284.6000 ;
	    RECT 688.5000 1283.1000 693.9000 1283.7001 ;
	    RECT 695.4000 1282.5000 696.3000 1283.7001 ;
	    RECT 722.1000 1283.1000 727.5000 1283.7001 ;
	    RECT 729.0000 1282.5000 729.9000 1283.7001 ;
	    RECT 640.2000 1281.4501 641.4000 1281.6000 ;
	    RECT 652.2000 1281.4501 653.4000 1281.6000 ;
	    RECT 640.2000 1280.5500 653.4000 1281.4501 ;
	    RECT 640.2000 1280.4000 641.4000 1280.5500 ;
	    RECT 652.2000 1280.4000 653.4000 1280.5500 ;
	    RECT 654.6000 1281.4501 655.8000 1281.6000 ;
	    RECT 654.6000 1280.5500 686.8500 1281.4501 ;
	    RECT 654.6000 1280.4000 655.8000 1280.5500 ;
	    RECT 637.8000 1278.4501 639.0000 1278.6000 ;
	    RECT 616.3500 1277.5500 639.0000 1278.4501 ;
	    RECT 616.3500 1275.6000 617.2500 1277.5500 ;
	    RECT 637.8000 1277.4000 639.0000 1277.5500 ;
	    RECT 609.0000 1263.3000 610.2000 1275.3000 ;
	    RECT 612.9000 1274.4000 614.4000 1275.3000 ;
	    RECT 616.2000 1274.4000 617.4000 1275.6000 ;
	    RECT 618.6000 1275.4501 619.8000 1275.6000 ;
	    RECT 635.4000 1275.4501 636.6000 1275.6000 ;
	    RECT 618.6000 1274.5500 636.6000 1275.4501 ;
	    RECT 618.6000 1274.4000 619.8000 1274.5500 ;
	    RECT 635.4000 1274.4000 636.6000 1274.5500 ;
	    RECT 612.9000 1263.3000 614.1000 1274.4000 ;
	    RECT 615.3000 1272.6000 616.2000 1273.5000 ;
	    RECT 635.4000 1273.2001 636.6000 1273.5000 ;
	    RECT 615.0000 1271.4000 616.2000 1272.6000 ;
	    RECT 615.3000 1263.3000 616.5000 1269.3000 ;
	    RECT 635.4000 1263.3000 636.6000 1269.3000 ;
	    RECT 637.8000 1263.3000 639.0000 1276.5000 ;
	    RECT 640.2000 1263.3000 641.4000 1269.3000 ;
	    RECT 652.2000 1263.3000 653.4000 1269.3000 ;
	    RECT 654.6000 1263.3000 655.8000 1279.5000 ;
	    RECT 685.9500 1278.4501 686.8500 1280.5500 ;
	    RECT 688.2000 1280.4000 689.4000 1281.6000 ;
	    RECT 690.3000 1280.7001 690.6000 1282.2001 ;
	    RECT 692.7000 1280.4000 694.5000 1281.6000 ;
	    RECT 695.4000 1280.4000 696.6000 1281.6000 ;
	    RECT 700.2000 1281.4501 701.4000 1281.6000 ;
	    RECT 721.8000 1281.4501 723.0000 1281.6000 ;
	    RECT 700.2000 1280.5500 723.0000 1281.4501 ;
	    RECT 723.9000 1280.7001 724.2000 1282.2001 ;
	    RECT 700.2000 1280.4000 701.4000 1280.5500 ;
	    RECT 721.8000 1280.4000 723.0000 1280.5500 ;
	    RECT 726.3000 1280.4000 728.1000 1281.6000 ;
	    RECT 729.0000 1280.4000 730.2000 1281.6000 ;
	    RECT 690.6000 1279.5000 691.8000 1279.8000 ;
	    RECT 690.6000 1278.4501 691.8000 1278.6000 ;
	    RECT 685.9500 1277.5500 691.8000 1278.4501 ;
	    RECT 690.6000 1277.4000 691.8000 1277.5500 ;
	    RECT 692.7000 1275.3000 693.6000 1280.4000 ;
	    RECT 724.2000 1279.5000 725.4000 1279.8000 ;
	    RECT 724.2000 1277.4000 725.4000 1278.6000 ;
	    RECT 688.2000 1263.3000 689.4000 1275.3000 ;
	    RECT 692.1000 1274.4000 693.6000 1275.3000 ;
	    RECT 695.4000 1274.4000 696.6000 1275.6000 ;
	    RECT 726.3000 1275.3000 727.2000 1280.4000 ;
	    RECT 750.6000 1279.5000 751.8000 1283.7001 ;
	    RECT 810.6000 1283.5500 886.2000 1284.4501 ;
	    RECT 810.6000 1283.4000 811.8000 1283.5500 ;
	    RECT 885.0000 1283.4000 886.2000 1283.5500 ;
	    RECT 753.0000 1282.5000 754.2000 1282.8000 ;
	    RECT 753.0000 1280.4000 754.2000 1281.6000 ;
	    RECT 887.4000 1280.7001 888.6000 1289.7001 ;
	    RECT 892.2000 1283.7001 893.4000 1289.7001 ;
	    RECT 897.0000 1284.9000 898.2000 1289.7001 ;
	    RECT 899.4000 1285.5000 900.6000 1289.7001 ;
	    RECT 901.8000 1285.5000 903.0000 1289.7001 ;
	    RECT 904.2000 1285.5000 905.4000 1289.7001 ;
	    RECT 906.6000 1286.7001 907.8000 1289.7001 ;
	    RECT 909.0000 1285.5000 910.2000 1289.7001 ;
	    RECT 911.4000 1286.7001 912.6000 1289.7001 ;
	    RECT 913.8000 1285.5000 915.0000 1289.7001 ;
	    RECT 916.2000 1285.5000 917.4000 1289.7001 ;
	    RECT 918.6000 1285.5000 919.8000 1289.7001 ;
	    RECT 921.0000 1285.5000 922.2000 1289.7001 ;
	    RECT 894.3000 1283.7001 898.2000 1284.9000 ;
	    RECT 923.4000 1284.9000 924.6000 1289.7001 ;
	    RECT 903.3000 1283.7001 910.2000 1284.6000 ;
	    RECT 894.3000 1282.8000 895.5000 1283.7001 ;
	    RECT 891.0000 1281.6000 895.5000 1282.8000 ;
	    RECT 887.4000 1279.5000 900.6000 1280.7001 ;
	    RECT 903.3000 1280.1000 904.5000 1283.7001 ;
	    RECT 909.0000 1283.4000 910.2000 1283.7001 ;
	    RECT 911.4000 1283.4000 912.6000 1284.6000 ;
	    RECT 913.5000 1283.4000 913.8000 1284.6000 ;
	    RECT 918.3000 1283.4000 919.8000 1284.6000 ;
	    RECT 923.4000 1283.7001 927.0000 1284.9000 ;
	    RECT 928.2000 1283.7001 929.4000 1289.7001 ;
	    RECT 906.6000 1282.5000 907.8000 1282.8000 ;
	    RECT 909.0000 1282.2001 910.2000 1282.5000 ;
	    RECT 906.6000 1280.4000 907.8000 1281.6000 ;
	    RECT 909.0000 1281.3000 915.6000 1282.2001 ;
	    RECT 914.4000 1281.0000 915.6000 1281.3000 ;
	    RECT 729.0000 1278.4501 730.2000 1278.6000 ;
	    RECT 750.6000 1278.4501 751.8000 1278.6000 ;
	    RECT 729.0000 1277.5500 751.8000 1278.4501 ;
	    RECT 729.0000 1277.4000 730.2000 1277.5500 ;
	    RECT 750.6000 1277.4000 751.8000 1277.5500 ;
	    RECT 837.0000 1278.4501 838.2000 1278.6000 ;
	    RECT 882.6000 1278.4501 883.8000 1278.6000 ;
	    RECT 837.0000 1277.5500 883.8000 1278.4501 ;
	    RECT 837.0000 1277.4000 838.2000 1277.5500 ;
	    RECT 882.6000 1277.4000 883.8000 1277.5500 ;
	    RECT 692.1000 1263.3000 693.3000 1274.4000 ;
	    RECT 694.5000 1272.6000 695.4000 1273.5000 ;
	    RECT 694.2000 1271.4000 695.4000 1272.6000 ;
	    RECT 694.5000 1263.3000 695.7000 1269.3000 ;
	    RECT 721.8000 1263.3000 723.0000 1275.3000 ;
	    RECT 725.7000 1274.4000 727.2000 1275.3000 ;
	    RECT 729.0000 1275.4501 730.2000 1275.6000 ;
	    RECT 738.6000 1275.4501 739.8000 1275.6000 ;
	    RECT 729.0000 1274.5500 739.8000 1275.4501 ;
	    RECT 729.0000 1274.4000 730.2000 1274.5500 ;
	    RECT 738.6000 1274.4000 739.8000 1274.5500 ;
	    RECT 741.0000 1275.4501 742.2000 1275.6000 ;
	    RECT 748.2000 1275.4501 749.4000 1275.6000 ;
	    RECT 741.0000 1274.5500 749.4000 1275.4501 ;
	    RECT 741.0000 1274.4000 742.2000 1274.5500 ;
	    RECT 748.2000 1274.4000 749.4000 1274.5500 ;
	    RECT 725.7000 1263.3000 726.9000 1274.4000 ;
	    RECT 728.1000 1272.6000 729.0000 1273.5000 ;
	    RECT 748.2000 1273.2001 749.4000 1273.5000 ;
	    RECT 727.8000 1271.4000 729.0000 1272.6000 ;
	    RECT 728.1000 1263.3000 729.3000 1269.3000 ;
	    RECT 748.2000 1263.3000 749.4000 1269.3000 ;
	    RECT 750.6000 1263.3000 751.8000 1276.5000 ;
	    RECT 753.0000 1272.4501 754.2000 1272.6000 ;
	    RECT 882.6000 1272.4501 883.8000 1272.6000 ;
	    RECT 753.0000 1271.5500 883.8000 1272.4501 ;
	    RECT 753.0000 1271.4000 754.2000 1271.5500 ;
	    RECT 882.6000 1271.4000 883.8000 1271.5500 ;
	    RECT 887.4000 1271.1000 888.6000 1279.5000 ;
	    RECT 901.5000 1278.9000 904.5000 1280.1000 ;
	    RECT 910.2000 1278.9000 915.0000 1280.1000 ;
	    RECT 918.6000 1279.2001 919.8000 1283.4000 ;
	    RECT 925.8000 1282.8000 927.0000 1283.7001 ;
	    RECT 925.8000 1281.9000 928.5000 1282.8000 ;
	    RECT 927.3000 1280.1000 928.5000 1281.9000 ;
	    RECT 933.0000 1281.9000 934.2000 1289.7001 ;
	    RECT 935.4000 1284.0000 936.6000 1289.7001 ;
	    RECT 937.8000 1286.7001 939.0000 1289.7001 ;
	    RECT 935.4000 1282.8000 936.9000 1284.0000 ;
	    RECT 933.0000 1281.0000 934.8000 1281.9000 ;
	    RECT 927.3000 1278.9000 933.0000 1280.1000 ;
	    RECT 889.5000 1278.0000 890.7000 1278.3000 ;
	    RECT 889.5000 1277.1000 896.1000 1278.0000 ;
	    RECT 897.0000 1277.4000 898.2000 1278.6000 ;
	    RECT 923.4000 1278.0000 924.6000 1278.9000 ;
	    RECT 933.9000 1278.0000 934.8000 1281.0000 ;
	    RECT 899.1000 1277.1000 924.6000 1278.0000 ;
	    RECT 933.6000 1277.1000 934.8000 1278.0000 ;
	    RECT 931.5000 1276.2001 932.7000 1276.5000 ;
	    RECT 892.2000 1274.4000 893.4000 1275.6000 ;
	    RECT 894.3000 1275.3000 932.7000 1276.2001 ;
	    RECT 897.3000 1275.0000 898.5000 1275.3000 ;
	    RECT 933.6000 1274.4000 934.5000 1277.1000 ;
	    RECT 935.7000 1276.2001 936.9000 1282.8000 ;
	    RECT 949.8000 1282.5000 951.0000 1289.7001 ;
	    RECT 952.2000 1286.7001 953.4000 1289.7001 ;
	    RECT 983.4000 1288.8000 989.4000 1289.7001 ;
	    RECT 952.2000 1285.5000 953.4000 1285.8000 ;
	    RECT 952.2000 1284.4501 953.4000 1284.6000 ;
	    RECT 969.0000 1284.4501 970.2000 1284.6000 ;
	    RECT 973.8000 1284.4501 975.0000 1284.6000 ;
	    RECT 952.2000 1283.5500 975.0000 1284.4501 ;
	    RECT 983.4000 1283.7001 984.6000 1288.8000 ;
	    RECT 985.8000 1283.7001 987.0000 1287.9000 ;
	    RECT 988.2000 1284.0000 989.4000 1288.8000 ;
	    RECT 990.6000 1284.9000 991.8000 1289.7001 ;
	    RECT 993.0000 1284.0000 994.2000 1289.7001 ;
	    RECT 1012.2000 1286.7001 1013.4000 1289.7001 ;
	    RECT 1014.6000 1286.7001 1015.8000 1289.7001 ;
	    RECT 1017.0000 1286.7001 1018.2000 1289.7001 ;
	    RECT 988.2000 1283.7001 994.2000 1284.0000 ;
	    RECT 952.2000 1283.4000 953.4000 1283.5500 ;
	    RECT 969.0000 1283.4000 970.2000 1283.5500 ;
	    RECT 973.8000 1283.4000 975.0000 1283.5500 ;
	    RECT 985.8000 1281.6000 986.7000 1283.7001 ;
	    RECT 988.5000 1283.1000 993.9000 1283.7001 ;
	    RECT 1014.6000 1282.5000 1015.5000 1286.7001 ;
	    RECT 1017.0000 1285.5000 1018.2000 1285.8000 ;
	    RECT 1017.0000 1284.4501 1018.2000 1284.6000 ;
	    RECT 1033.8000 1284.4501 1035.0000 1284.6000 ;
	    RECT 1017.0000 1283.5500 1035.0000 1284.4501 ;
	    RECT 1048.2001 1284.0000 1049.4000 1289.7001 ;
	    RECT 1050.6000 1284.9000 1051.8000 1289.7001 ;
	    RECT 1053.0000 1288.8000 1059.0000 1289.7001 ;
	    RECT 1053.0000 1284.0000 1054.2001 1288.8000 ;
	    RECT 1048.2001 1283.7001 1054.2001 1284.0000 ;
	    RECT 1055.4000 1283.7001 1056.6000 1287.9000 ;
	    RECT 1057.8000 1283.7001 1059.0000 1288.8000 ;
	    RECT 1017.0000 1283.4000 1018.2000 1283.5500 ;
	    RECT 1033.8000 1283.4000 1035.0000 1283.5500 ;
	    RECT 1048.5000 1283.1000 1053.9000 1283.7001 ;
	    RECT 949.8000 1281.4501 951.0000 1281.6000 ;
	    RECT 957.0000 1281.4501 958.2000 1281.6000 ;
	    RECT 949.8000 1280.5500 958.2000 1281.4501 ;
	    RECT 949.8000 1280.4000 951.0000 1280.5500 ;
	    RECT 957.0000 1280.4000 958.2000 1280.5500 ;
	    RECT 978.6000 1281.4501 979.8000 1281.6000 ;
	    RECT 983.4000 1281.4501 984.6000 1281.6000 ;
	    RECT 978.6000 1280.5500 984.6000 1281.4501 ;
	    RECT 985.8000 1280.7001 987.3000 1281.6000 ;
	    RECT 978.6000 1280.4000 979.8000 1280.5500 ;
	    RECT 983.4000 1280.4000 984.6000 1280.5500 ;
	    RECT 988.2000 1280.4000 989.4000 1281.6000 ;
	    RECT 991.8000 1280.7001 992.1000 1282.2001 ;
	    RECT 993.0000 1280.4000 994.2000 1281.6000 ;
	    RECT 995.4000 1281.4501 996.6000 1281.6000 ;
	    RECT 1014.6000 1281.4501 1015.8000 1281.6000 ;
	    RECT 995.4000 1280.5500 1015.8000 1281.4501 ;
	    RECT 995.4000 1280.4000 996.6000 1280.5500 ;
	    RECT 1014.6000 1280.4000 1015.8000 1280.5500 ;
	    RECT 1045.8000 1281.4501 1047.0000 1281.6000 ;
	    RECT 1048.2001 1281.4501 1049.4000 1281.6000 ;
	    RECT 1045.8000 1280.5500 1049.4000 1281.4501 ;
	    RECT 1050.3000 1280.7001 1050.6000 1282.2001 ;
	    RECT 1055.7001 1281.6000 1056.6000 1283.7001 ;
	    RECT 1072.2001 1282.5000 1073.4000 1289.7001 ;
	    RECT 1074.6000 1286.7001 1075.8000 1289.7001 ;
	    RECT 1081.8000 1287.4501 1083.0000 1287.6000 ;
	    RECT 1108.2001 1287.4501 1109.4000 1287.6000 ;
	    RECT 1206.6000 1287.4501 1207.8000 1287.6000 ;
	    RECT 1081.8000 1286.5500 1207.8000 1287.4501 ;
	    RECT 1081.8000 1286.4000 1083.0000 1286.5500 ;
	    RECT 1108.2001 1286.4000 1109.4000 1286.5500 ;
	    RECT 1206.6000 1286.4000 1207.8000 1286.5500 ;
	    RECT 1074.6000 1285.5000 1075.8000 1285.8000 ;
	    RECT 1074.6000 1283.4000 1075.8000 1284.6000 ;
	    RECT 1045.8000 1280.4000 1047.0000 1280.5500 ;
	    RECT 1048.2001 1280.4000 1049.4000 1280.5500 ;
	    RECT 1053.0000 1280.4000 1054.2001 1281.6000 ;
	    RECT 1055.1000 1280.7001 1056.6000 1281.6000 ;
	    RECT 1057.8000 1281.4501 1059.0000 1281.6000 ;
	    RECT 1072.2001 1281.4501 1073.4000 1281.6000 ;
	    RECT 1057.8000 1280.5500 1073.4000 1281.4501 ;
	    RECT 1057.8000 1280.4000 1059.0000 1280.5500 ;
	    RECT 1072.2001 1280.4000 1073.4000 1280.5500 ;
	    RECT 1209.0000 1280.7001 1210.2001 1289.7001 ;
	    RECT 1213.8000 1283.7001 1215.0000 1289.7001 ;
	    RECT 1218.6000 1284.9000 1219.8000 1289.7001 ;
	    RECT 1221.0000 1285.5000 1222.2001 1289.7001 ;
	    RECT 1223.4000 1285.5000 1224.6000 1289.7001 ;
	    RECT 1225.8000 1285.5000 1227.0000 1289.7001 ;
	    RECT 1228.2001 1286.7001 1229.4000 1289.7001 ;
	    RECT 1230.6000 1285.5000 1231.8000 1289.7001 ;
	    RECT 1233.0000 1286.7001 1234.2001 1289.7001 ;
	    RECT 1235.4000 1285.5000 1236.6000 1289.7001 ;
	    RECT 1237.8000 1285.5000 1239.0000 1289.7001 ;
	    RECT 1240.2001 1285.5000 1241.4000 1289.7001 ;
	    RECT 1242.6000 1285.5000 1243.8000 1289.7001 ;
	    RECT 1215.9000 1283.7001 1219.8000 1284.9000 ;
	    RECT 1245.0000 1284.9000 1246.2001 1289.7001 ;
	    RECT 1224.9000 1283.7001 1231.8000 1284.6000 ;
	    RECT 1215.9000 1282.8000 1217.1000 1283.7001 ;
	    RECT 1212.6000 1281.6000 1217.1000 1282.8000 ;
	    RECT 985.8000 1279.5000 987.0000 1279.8000 ;
	    RECT 990.6000 1279.5000 991.8000 1279.8000 ;
	    RECT 1050.6000 1279.5000 1051.8000 1279.8000 ;
	    RECT 1055.4000 1279.5000 1056.6000 1279.8000 ;
	    RECT 1209.0000 1279.5000 1222.2001 1280.7001 ;
	    RECT 1224.9000 1280.1000 1226.1000 1283.7001 ;
	    RECT 1230.6000 1283.4000 1231.8000 1283.7001 ;
	    RECT 1233.0000 1283.4000 1234.2001 1284.6000 ;
	    RECT 1235.1000 1283.4000 1235.4000 1284.6000 ;
	    RECT 1239.9000 1283.4000 1241.4000 1284.6000 ;
	    RECT 1245.0000 1283.7001 1248.6000 1284.9000 ;
	    RECT 1249.8000 1283.7001 1251.0000 1289.7001 ;
	    RECT 1228.2001 1282.5000 1229.4000 1282.8000 ;
	    RECT 1230.6000 1282.2001 1231.8000 1282.5000 ;
	    RECT 1228.2001 1280.4000 1229.4000 1281.6000 ;
	    RECT 1230.6000 1281.3000 1237.2001 1282.2001 ;
	    RECT 1236.0000 1281.0000 1237.2001 1281.3000 ;
	    RECT 901.8000 1274.1000 903.0000 1274.4000 ;
	    RECT 894.9000 1273.5000 903.0000 1274.1000 ;
	    RECT 893.7000 1273.2001 903.0000 1273.5000 ;
	    RECT 904.5000 1273.5000 917.4000 1274.4000 ;
	    RECT 889.8000 1272.0000 892.2000 1273.2001 ;
	    RECT 893.7000 1272.3000 895.8000 1273.2001 ;
	    RECT 904.5000 1272.3000 905.4000 1273.5000 ;
	    RECT 916.2000 1273.2001 917.4000 1273.5000 ;
	    RECT 921.0000 1273.5000 934.5000 1274.4000 ;
	    RECT 935.4000 1275.0000 936.9000 1276.2001 ;
	    RECT 935.4000 1273.5000 936.6000 1275.0000 ;
	    RECT 921.0000 1273.2001 922.2000 1273.5000 ;
	    RECT 891.3000 1271.4000 892.2000 1272.0000 ;
	    RECT 896.7000 1271.4000 905.4000 1272.3000 ;
	    RECT 906.3000 1271.4000 910.2000 1272.6000 ;
	    RECT 887.4000 1270.2001 890.4000 1271.1000 ;
	    RECT 891.3000 1270.2001 897.6000 1271.4000 ;
	    RECT 889.5000 1269.3000 890.4000 1270.2001 ;
	    RECT 753.0000 1263.3000 754.2000 1269.3000 ;
	    RECT 813.0000 1266.4501 814.2000 1266.6000 ;
	    RECT 885.0000 1266.4501 886.2000 1266.6000 ;
	    RECT 813.0000 1265.5500 886.2000 1266.4501 ;
	    RECT 813.0000 1265.4000 814.2000 1265.5500 ;
	    RECT 885.0000 1265.4000 886.2000 1265.5500 ;
	    RECT 887.4000 1263.3000 888.6000 1269.3000 ;
	    RECT 889.5000 1268.4000 891.0000 1269.3000 ;
	    RECT 889.8000 1263.3000 891.0000 1268.4000 ;
	    RECT 892.2000 1262.4000 893.4000 1269.3000 ;
	    RECT 894.6000 1263.3000 895.8000 1270.2001 ;
	    RECT 897.0000 1263.3000 898.2000 1269.3000 ;
	    RECT 899.4000 1263.3000 900.6000 1267.5000 ;
	    RECT 901.8000 1263.3000 903.0000 1267.5000 ;
	    RECT 904.2000 1263.3000 905.4000 1270.5000 ;
	    RECT 906.6000 1263.3000 907.8000 1269.3000 ;
	    RECT 909.0000 1263.3000 910.2000 1270.5000 ;
	    RECT 911.4000 1263.3000 912.6000 1269.3000 ;
	    RECT 913.8000 1263.3000 915.0000 1272.6000 ;
	    RECT 925.8000 1271.4000 929.7000 1272.6000 ;
	    RECT 918.6000 1270.2001 924.9000 1271.4000 ;
	    RECT 916.2000 1263.3000 917.4000 1267.5000 ;
	    RECT 918.6000 1263.3000 919.8000 1267.5000 ;
	    RECT 921.0000 1263.3000 922.2000 1267.5000 ;
	    RECT 923.4000 1263.3000 924.6000 1269.3000 ;
	    RECT 925.8000 1263.3000 927.0000 1271.4000 ;
	    RECT 933.6000 1271.1000 934.5000 1273.5000 ;
	    RECT 935.4000 1271.4000 936.6000 1272.6000 ;
	    RECT 930.6000 1270.2001 934.5000 1271.1000 ;
	    RECT 928.2000 1263.3000 929.4000 1269.3000 ;
	    RECT 930.6000 1263.3000 931.8000 1270.2001 ;
	    RECT 933.0000 1263.3000 934.2000 1269.3000 ;
	    RECT 935.4000 1263.3000 936.6000 1270.5000 ;
	    RECT 937.8000 1263.3000 939.0000 1269.3000 ;
	    RECT 949.8000 1263.3000 951.0000 1279.5000 ;
	    RECT 983.4000 1279.2001 984.6000 1279.5000 ;
	    RECT 985.8000 1277.4000 987.0000 1278.6000 ;
	    RECT 988.5000 1275.3000 989.4000 1279.5000 ;
	    RECT 990.6000 1278.4501 991.8000 1278.6000 ;
	    RECT 997.8000 1278.4501 999.0000 1278.6000 ;
	    RECT 990.6000 1277.5500 999.0000 1278.4501 ;
	    RECT 990.6000 1277.4000 991.8000 1277.5500 ;
	    RECT 997.8000 1277.4000 999.0000 1277.5500 ;
	    RECT 1012.2000 1277.4000 1013.4000 1278.6000 ;
	    RECT 1012.2000 1276.2001 1013.4000 1276.5000 ;
	    RECT 1014.6000 1275.3000 1015.5000 1279.5000 ;
	    RECT 1050.6000 1277.4000 1051.8000 1278.6000 ;
	    RECT 1053.0000 1275.3000 1053.9000 1279.5000 ;
	    RECT 1057.8000 1279.2001 1059.0000 1279.5000 ;
	    RECT 1055.4000 1277.4000 1056.6000 1278.6000 ;
	    RECT 952.2000 1263.3000 953.4000 1269.3000 ;
	    RECT 983.4000 1263.3000 984.6000 1275.3000 ;
	    RECT 987.3000 1263.3000 990.3000 1275.3000 ;
	    RECT 993.0000 1263.3000 994.2000 1275.3000 ;
	    RECT 1013.1000 1274.1000 1015.8000 1275.3000 ;
	    RECT 1013.1000 1263.3000 1014.3000 1274.1000 ;
	    RECT 1017.0000 1263.3000 1018.2000 1275.3000 ;
	    RECT 1048.2001 1263.3000 1049.4000 1275.3000 ;
	    RECT 1052.1000 1263.3000 1055.1000 1275.3000 ;
	    RECT 1057.8000 1263.3000 1059.0000 1275.3000 ;
	    RECT 1072.2001 1263.3000 1073.4000 1279.5000 ;
	    RECT 1084.2001 1272.4501 1085.4000 1272.6000 ;
	    RECT 1168.2001 1272.4501 1169.4000 1272.6000 ;
	    RECT 1084.2001 1271.5500 1169.4000 1272.4501 ;
	    RECT 1084.2001 1271.4000 1085.4000 1271.5500 ;
	    RECT 1168.2001 1271.4000 1169.4000 1271.5500 ;
	    RECT 1209.0000 1271.1000 1210.2001 1279.5000 ;
	    RECT 1223.1000 1278.9000 1226.1000 1280.1000 ;
	    RECT 1231.8000 1278.9000 1236.6000 1280.1000 ;
	    RECT 1240.2001 1279.2001 1241.4000 1283.4000 ;
	    RECT 1247.4000 1282.8000 1248.6000 1283.7001 ;
	    RECT 1247.4000 1281.9000 1250.1000 1282.8000 ;
	    RECT 1248.9000 1280.1000 1250.1000 1281.9000 ;
	    RECT 1254.6000 1281.9000 1255.8000 1289.7001 ;
	    RECT 1257.0000 1284.0000 1258.2001 1289.7001 ;
	    RECT 1259.4000 1286.7001 1260.6000 1289.7001 ;
	    RECT 1273.8000 1286.7001 1275.0000 1289.7001 ;
	    RECT 1273.8000 1285.5000 1275.0000 1285.8000 ;
	    RECT 1257.0000 1282.8000 1258.5000 1284.0000 ;
	    RECT 1273.8000 1283.4000 1275.0000 1284.6000 ;
	    RECT 1254.6000 1281.0000 1256.4000 1281.9000 ;
	    RECT 1248.9000 1278.9000 1254.6000 1280.1000 ;
	    RECT 1211.1000 1278.0000 1212.3000 1278.3000 ;
	    RECT 1211.1000 1277.1000 1217.7001 1278.0000 ;
	    RECT 1218.6000 1277.4000 1219.8000 1278.6000 ;
	    RECT 1245.0000 1278.0000 1246.2001 1278.9000 ;
	    RECT 1255.5000 1278.0000 1256.4000 1281.0000 ;
	    RECT 1220.7001 1277.1000 1246.2001 1278.0000 ;
	    RECT 1255.2001 1277.1000 1256.4000 1278.0000 ;
	    RECT 1253.1000 1276.2001 1254.3000 1276.5000 ;
	    RECT 1213.8000 1274.4000 1215.0000 1275.6000 ;
	    RECT 1215.9000 1275.3000 1254.3000 1276.2001 ;
	    RECT 1218.9000 1275.0000 1220.1000 1275.3000 ;
	    RECT 1255.2001 1274.4000 1256.1000 1277.1000 ;
	    RECT 1257.3000 1276.2001 1258.5000 1282.8000 ;
	    RECT 1276.2001 1282.5000 1277.4000 1289.7001 ;
	    RECT 1296.3000 1284.6000 1297.5000 1289.7001 ;
	    RECT 1296.3000 1283.7001 1299.0000 1284.6000 ;
	    RECT 1300.2001 1283.7001 1301.4000 1289.7001 ;
	    RECT 1432.2001 1286.7001 1433.4000 1289.7001 ;
	    RECT 1434.6000 1284.0000 1435.8000 1289.7001 ;
	    RECT 1276.2001 1281.4501 1277.4000 1281.6000 ;
	    RECT 1281.0000 1281.4501 1282.2001 1281.6000 ;
	    RECT 1276.2001 1280.5500 1282.2001 1281.4501 ;
	    RECT 1276.2001 1280.4000 1277.4000 1280.5500 ;
	    RECT 1281.0000 1280.4000 1282.2001 1280.5500 ;
	    RECT 1297.8000 1279.5000 1299.0000 1283.7001 ;
	    RECT 1434.3000 1282.8000 1435.8000 1284.0000 ;
	    RECT 1300.2001 1282.5000 1301.4000 1282.8000 ;
	    RECT 1300.2001 1281.4501 1301.4000 1281.6000 ;
	    RECT 1326.6000 1281.4501 1327.8000 1281.6000 ;
	    RECT 1300.2001 1280.5500 1327.8000 1281.4501 ;
	    RECT 1300.2001 1280.4000 1301.4000 1280.5500 ;
	    RECT 1326.6000 1280.4000 1327.8000 1280.5500 ;
	    RECT 1223.4000 1274.1000 1224.6000 1274.4000 ;
	    RECT 1216.5000 1273.5000 1224.6000 1274.1000 ;
	    RECT 1215.3000 1273.2001 1224.6000 1273.5000 ;
	    RECT 1226.1000 1273.5000 1239.0000 1274.4000 ;
	    RECT 1211.4000 1272.0000 1213.8000 1273.2001 ;
	    RECT 1215.3000 1272.3000 1217.4000 1273.2001 ;
	    RECT 1226.1000 1272.3000 1227.0000 1273.5000 ;
	    RECT 1237.8000 1273.2001 1239.0000 1273.5000 ;
	    RECT 1242.6000 1273.5000 1256.1000 1274.4000 ;
	    RECT 1257.0000 1275.0000 1258.5000 1276.2001 ;
	    RECT 1257.0000 1273.5000 1258.2001 1275.0000 ;
	    RECT 1242.6000 1273.2001 1243.8000 1273.5000 ;
	    RECT 1212.9000 1271.4000 1213.8000 1272.0000 ;
	    RECT 1218.3000 1271.4000 1227.0000 1272.3000 ;
	    RECT 1227.9000 1271.4000 1231.8000 1272.6000 ;
	    RECT 1209.0000 1270.2001 1212.0000 1271.1000 ;
	    RECT 1212.9000 1270.2001 1219.2001 1271.4000 ;
	    RECT 1211.1000 1269.3000 1212.0000 1270.2001 ;
	    RECT 1074.6000 1263.3000 1075.8000 1269.3000 ;
	    RECT 1209.0000 1263.3000 1210.2001 1269.3000 ;
	    RECT 1211.1000 1268.4000 1212.6000 1269.3000 ;
	    RECT 1211.4000 1263.3000 1212.6000 1268.4000 ;
	    RECT 1213.8000 1262.4000 1215.0000 1269.3000 ;
	    RECT 1216.2001 1263.3000 1217.4000 1270.2001 ;
	    RECT 1218.6000 1263.3000 1219.8000 1269.3000 ;
	    RECT 1221.0000 1263.3000 1222.2001 1267.5000 ;
	    RECT 1223.4000 1263.3000 1224.6000 1267.5000 ;
	    RECT 1225.8000 1263.3000 1227.0000 1270.5000 ;
	    RECT 1228.2001 1263.3000 1229.4000 1269.3000 ;
	    RECT 1230.6000 1263.3000 1231.8000 1270.5000 ;
	    RECT 1233.0000 1263.3000 1234.2001 1269.3000 ;
	    RECT 1235.4000 1263.3000 1236.6000 1272.6000 ;
	    RECT 1247.4000 1271.4000 1251.3000 1272.6000 ;
	    RECT 1240.2001 1270.2001 1246.5000 1271.4000 ;
	    RECT 1237.8000 1263.3000 1239.0000 1267.5000 ;
	    RECT 1240.2001 1263.3000 1241.4000 1267.5000 ;
	    RECT 1242.6000 1263.3000 1243.8000 1267.5000 ;
	    RECT 1245.0000 1263.3000 1246.2001 1269.3000 ;
	    RECT 1247.4000 1263.3000 1248.6000 1271.4000 ;
	    RECT 1255.2001 1271.1000 1256.1000 1273.5000 ;
	    RECT 1257.0000 1271.4000 1258.2001 1272.6000 ;
	    RECT 1252.2001 1270.2001 1256.1000 1271.1000 ;
	    RECT 1249.8000 1263.3000 1251.0000 1269.3000 ;
	    RECT 1252.2001 1263.3000 1253.4000 1270.2001 ;
	    RECT 1254.6000 1263.3000 1255.8000 1269.3000 ;
	    RECT 1257.0000 1263.3000 1258.2001 1270.5000 ;
	    RECT 1259.4000 1263.3000 1260.6000 1269.3000 ;
	    RECT 1273.8000 1263.3000 1275.0000 1269.3000 ;
	    RECT 1276.2001 1263.3000 1277.4000 1279.5000 ;
	    RECT 1283.4000 1278.4501 1284.6000 1278.6000 ;
	    RECT 1297.8000 1278.4501 1299.0000 1278.6000 ;
	    RECT 1283.4000 1277.5500 1299.0000 1278.4501 ;
	    RECT 1283.4000 1277.4000 1284.6000 1277.5500 ;
	    RECT 1297.8000 1277.4000 1299.0000 1277.5500 ;
	    RECT 1295.4000 1274.4000 1296.6000 1275.6000 ;
	    RECT 1295.4000 1273.2001 1296.6000 1273.5000 ;
	    RECT 1295.4000 1263.3000 1296.6000 1269.3000 ;
	    RECT 1297.8000 1263.3000 1299.0000 1276.5000 ;
	    RECT 1434.3000 1276.2001 1435.5000 1282.8000 ;
	    RECT 1437.0000 1281.9000 1438.2001 1289.7001 ;
	    RECT 1441.8000 1283.7001 1443.0000 1289.7001 ;
	    RECT 1446.6000 1284.9000 1447.8000 1289.7001 ;
	    RECT 1449.0000 1285.5000 1450.2001 1289.7001 ;
	    RECT 1451.4000 1285.5000 1452.6000 1289.7001 ;
	    RECT 1453.8000 1285.5000 1455.0000 1289.7001 ;
	    RECT 1456.2001 1285.5000 1457.4000 1289.7001 ;
	    RECT 1458.6000 1286.7001 1459.8000 1289.7001 ;
	    RECT 1461.0000 1285.5000 1462.2001 1289.7001 ;
	    RECT 1463.4000 1286.7001 1464.6000 1289.7001 ;
	    RECT 1465.8000 1285.5000 1467.0000 1289.7001 ;
	    RECT 1468.2001 1285.5000 1469.4000 1289.7001 ;
	    RECT 1470.6000 1285.5000 1471.8000 1289.7001 ;
	    RECT 1444.2001 1283.7001 1447.8000 1284.9000 ;
	    RECT 1473.0000 1284.9000 1474.2001 1289.7001 ;
	    RECT 1444.2001 1282.8000 1445.4000 1283.7001 ;
	    RECT 1436.4000 1281.0000 1438.2001 1281.9000 ;
	    RECT 1442.7001 1281.9000 1445.4000 1282.8000 ;
	    RECT 1451.4000 1283.4000 1452.9000 1284.6000 ;
	    RECT 1457.4000 1283.4000 1457.7001 1284.6000 ;
	    RECT 1458.6000 1283.4000 1459.8000 1284.6000 ;
	    RECT 1461.0000 1283.7001 1467.9000 1284.6000 ;
	    RECT 1473.0000 1283.7001 1476.9000 1284.9000 ;
	    RECT 1477.8000 1283.7001 1479.0000 1289.7001 ;
	    RECT 1461.0000 1283.4000 1462.2001 1283.7001 ;
	    RECT 1436.4000 1278.0000 1437.3000 1281.0000 ;
	    RECT 1442.7001 1280.1000 1443.9000 1281.9000 ;
	    RECT 1438.2001 1278.9000 1443.9000 1280.1000 ;
	    RECT 1451.4000 1279.2001 1452.6000 1283.4000 ;
	    RECT 1463.4000 1282.5000 1464.6000 1282.8000 ;
	    RECT 1461.0000 1282.2001 1462.2001 1282.5000 ;
	    RECT 1455.6000 1281.3000 1462.2001 1282.2001 ;
	    RECT 1455.6000 1281.0000 1456.8000 1281.3000 ;
	    RECT 1463.4000 1280.4000 1464.6000 1281.6000 ;
	    RECT 1466.7001 1280.1000 1467.9000 1283.7001 ;
	    RECT 1475.7001 1282.8000 1476.9000 1283.7001 ;
	    RECT 1475.7001 1281.6000 1480.2001 1282.8000 ;
	    RECT 1482.6000 1280.7001 1483.8000 1289.7001 ;
	    RECT 1497.0000 1282.5000 1498.2001 1289.7001 ;
	    RECT 1499.4000 1286.7001 1500.6000 1289.7001 ;
	    RECT 1499.4000 1285.5000 1500.6000 1285.8000 ;
	    RECT 1519.5000 1284.6000 1520.7001 1289.7001 ;
	    RECT 1499.4000 1284.4501 1500.6000 1284.6000 ;
	    RECT 1509.0000 1284.4501 1510.2001 1284.6000 ;
	    RECT 1513.8000 1284.4501 1515.0000 1284.6000 ;
	    RECT 1499.4000 1283.5500 1515.0000 1284.4501 ;
	    RECT 1519.5000 1283.7001 1522.2001 1284.6000 ;
	    RECT 1523.4000 1283.7001 1524.6000 1289.7001 ;
	    RECT 1543.5000 1284.6000 1544.7001 1289.7001 ;
	    RECT 1543.5000 1283.7001 1546.2001 1284.6000 ;
	    RECT 1547.4000 1283.7001 1548.6000 1289.7001 ;
	    RECT 1499.4000 1283.4000 1500.6000 1283.5500 ;
	    RECT 1509.0000 1283.4000 1510.2001 1283.5500 ;
	    RECT 1513.8000 1283.4000 1515.0000 1283.5500 ;
	    RECT 1456.2001 1278.9000 1461.0000 1280.1000 ;
	    RECT 1466.7001 1278.9000 1469.7001 1280.1000 ;
	    RECT 1470.6000 1279.5000 1483.8000 1280.7001 ;
	    RECT 1485.0000 1281.4501 1486.2001 1281.6000 ;
	    RECT 1497.0000 1281.4501 1498.2001 1281.6000 ;
	    RECT 1485.0000 1280.5500 1498.2001 1281.4501 ;
	    RECT 1485.0000 1280.4000 1486.2001 1280.5500 ;
	    RECT 1497.0000 1280.4000 1498.2001 1280.5500 ;
	    RECT 1521.0000 1279.5000 1522.2001 1283.7001 ;
	    RECT 1523.4000 1282.5000 1524.6000 1282.8000 ;
	    RECT 1523.4000 1280.4000 1524.6000 1281.6000 ;
	    RECT 1545.0000 1279.5000 1546.2001 1283.7001 ;
	    RECT 1547.4000 1282.5000 1548.6000 1282.8000 ;
	    RECT 1547.4000 1280.4000 1548.6000 1281.6000 ;
	    RECT 1446.6000 1278.0000 1447.8000 1278.9000 ;
	    RECT 1436.4000 1277.1000 1437.6000 1278.0000 ;
	    RECT 1446.6000 1277.1000 1472.1000 1278.0000 ;
	    RECT 1473.0000 1277.4000 1474.2001 1278.6000 ;
	    RECT 1480.5000 1278.0000 1481.7001 1278.3000 ;
	    RECT 1475.1000 1277.1000 1481.7001 1278.0000 ;
	    RECT 1434.3000 1275.0000 1435.8000 1276.2001 ;
	    RECT 1434.6000 1273.5000 1435.8000 1275.0000 ;
	    RECT 1436.7001 1274.4000 1437.6000 1277.1000 ;
	    RECT 1438.5000 1276.2001 1439.7001 1276.5000 ;
	    RECT 1438.5000 1275.3000 1476.9000 1276.2001 ;
	    RECT 1472.7001 1275.0000 1473.9000 1275.3000 ;
	    RECT 1477.8000 1274.4000 1479.0000 1275.6000 ;
	    RECT 1436.7001 1273.5000 1450.2001 1274.4000 ;
	    RECT 1302.6000 1272.4501 1303.8000 1272.6000 ;
	    RECT 1434.6000 1272.4501 1435.8000 1272.6000 ;
	    RECT 1302.6000 1271.5500 1435.8000 1272.4501 ;
	    RECT 1302.6000 1271.4000 1303.8000 1271.5500 ;
	    RECT 1434.6000 1271.4000 1435.8000 1271.5500 ;
	    RECT 1436.7001 1271.1000 1437.6000 1273.5000 ;
	    RECT 1449.0000 1273.2001 1450.2001 1273.5000 ;
	    RECT 1453.8000 1273.5000 1466.7001 1274.4000 ;
	    RECT 1453.8000 1273.2001 1455.0000 1273.5000 ;
	    RECT 1441.5000 1271.4000 1445.4000 1272.6000 ;
	    RECT 1300.2001 1263.3000 1301.4000 1269.3000 ;
	    RECT 1432.2001 1263.3000 1433.4000 1269.3000 ;
	    RECT 1434.6000 1263.3000 1435.8000 1270.5000 ;
	    RECT 1436.7001 1270.2001 1440.6000 1271.1000 ;
	    RECT 1437.0000 1263.3000 1438.2001 1269.3000 ;
	    RECT 1439.4000 1263.3000 1440.6000 1270.2001 ;
	    RECT 1441.8000 1263.3000 1443.0000 1269.3000 ;
	    RECT 1444.2001 1263.3000 1445.4000 1271.4000 ;
	    RECT 1446.3000 1270.2001 1452.6000 1271.4000 ;
	    RECT 1446.6000 1263.3000 1447.8000 1269.3000 ;
	    RECT 1449.0000 1263.3000 1450.2001 1267.5000 ;
	    RECT 1451.4000 1263.3000 1452.6000 1267.5000 ;
	    RECT 1453.8000 1263.3000 1455.0000 1267.5000 ;
	    RECT 1456.2001 1263.3000 1457.4000 1272.6000 ;
	    RECT 1461.0000 1271.4000 1464.9000 1272.6000 ;
	    RECT 1465.8000 1272.3000 1466.7001 1273.5000 ;
	    RECT 1468.2001 1274.1000 1469.4000 1274.4000 ;
	    RECT 1468.2001 1273.5000 1476.3000 1274.1000 ;
	    RECT 1468.2001 1273.2001 1477.5000 1273.5000 ;
	    RECT 1475.4000 1272.3000 1477.5000 1273.2001 ;
	    RECT 1465.8000 1271.4000 1474.5000 1272.3000 ;
	    RECT 1479.0000 1272.0000 1481.4000 1273.2001 ;
	    RECT 1479.0000 1271.4000 1479.9000 1272.0000 ;
	    RECT 1458.6000 1263.3000 1459.8000 1269.3000 ;
	    RECT 1461.0000 1263.3000 1462.2001 1270.5000 ;
	    RECT 1463.4000 1263.3000 1464.6000 1269.3000 ;
	    RECT 1465.8000 1263.3000 1467.0000 1270.5000 ;
	    RECT 1473.6000 1270.2001 1479.9000 1271.4000 ;
	    RECT 1482.6000 1271.1000 1483.8000 1279.5000 ;
	    RECT 1480.8000 1270.2001 1483.8000 1271.1000 ;
	    RECT 1468.2001 1263.3000 1469.4000 1267.5000 ;
	    RECT 1470.6000 1263.3000 1471.8000 1267.5000 ;
	    RECT 1473.0000 1263.3000 1474.2001 1269.3000 ;
	    RECT 1475.4000 1263.3000 1476.6000 1270.2001 ;
	    RECT 1480.8000 1269.3000 1481.7001 1270.2001 ;
	    RECT 1477.8000 1262.4000 1479.0000 1269.3000 ;
	    RECT 1480.2001 1268.4000 1481.7001 1269.3000 ;
	    RECT 1480.2001 1263.3000 1481.4000 1268.4000 ;
	    RECT 1482.6000 1263.3000 1483.8000 1269.3000 ;
	    RECT 1497.0000 1263.3000 1498.2001 1279.5000 ;
	    RECT 1501.8000 1278.4501 1503.0000 1278.6000 ;
	    RECT 1521.0000 1278.4501 1522.2001 1278.6000 ;
	    RECT 1501.8000 1277.5500 1522.2001 1278.4501 ;
	    RECT 1501.8000 1277.4000 1503.0000 1277.5500 ;
	    RECT 1521.0000 1277.4000 1522.2001 1277.5500 ;
	    RECT 1540.2001 1278.4501 1541.4000 1278.6000 ;
	    RECT 1545.0000 1278.4501 1546.2001 1278.6000 ;
	    RECT 1540.2001 1277.5500 1546.2001 1278.4501 ;
	    RECT 1540.2001 1277.4000 1541.4000 1277.5500 ;
	    RECT 1545.0000 1277.4000 1546.2001 1277.5500 ;
	    RECT 1509.0000 1275.4501 1510.2001 1275.6000 ;
	    RECT 1518.6000 1275.4501 1519.8000 1275.6000 ;
	    RECT 1509.0000 1274.5500 1519.8000 1275.4501 ;
	    RECT 1509.0000 1274.4000 1510.2001 1274.5500 ;
	    RECT 1518.6000 1274.4000 1519.8000 1274.5500 ;
	    RECT 1518.6000 1273.2001 1519.8000 1273.5000 ;
	    RECT 1499.4000 1263.3000 1500.6000 1269.3000 ;
	    RECT 1518.6000 1263.3000 1519.8000 1269.3000 ;
	    RECT 1521.0000 1263.3000 1522.2001 1276.5000 ;
	    RECT 1537.8000 1275.4501 1539.0000 1275.6000 ;
	    RECT 1542.6000 1275.4501 1543.8000 1275.6000 ;
	    RECT 1537.8000 1274.5500 1543.8000 1275.4501 ;
	    RECT 1537.8000 1274.4000 1539.0000 1274.5500 ;
	    RECT 1542.6000 1274.4000 1543.8000 1274.5500 ;
	    RECT 1542.6000 1273.2001 1543.8000 1273.5000 ;
	    RECT 1523.4000 1263.3000 1524.6000 1269.3000 ;
	    RECT 1542.6000 1263.3000 1543.8000 1269.3000 ;
	    RECT 1545.0000 1263.3000 1546.2001 1276.5000 ;
	    RECT 1547.4000 1263.3000 1548.6000 1269.3000 ;
	    RECT 1.2000 1260.6000 1569.0000 1262.4000 ;
	    RECT 126.6000 1253.7001 127.8000 1259.7001 ;
	    RECT 129.0000 1254.6000 130.2000 1259.7001 ;
	    RECT 128.7000 1253.7001 130.2000 1254.6000 ;
	    RECT 131.4000 1253.7001 132.6000 1260.6000 ;
	    RECT 128.7000 1252.8000 129.6000 1253.7001 ;
	    RECT 133.8000 1252.8000 135.0000 1259.7001 ;
	    RECT 136.2000 1253.7001 137.4000 1259.7001 ;
	    RECT 138.6000 1255.5000 139.8000 1259.7001 ;
	    RECT 141.0000 1255.5000 142.2000 1259.7001 ;
	    RECT 126.6000 1251.9000 129.6000 1252.8000 ;
	    RECT 33.0000 1248.4501 34.2000 1248.6000 ;
	    RECT 124.2000 1248.4501 125.4000 1248.6000 ;
	    RECT 33.0000 1247.5500 125.4000 1248.4501 ;
	    RECT 33.0000 1247.4000 34.2000 1247.5500 ;
	    RECT 124.2000 1247.4000 125.4000 1247.5500 ;
	    RECT 126.6000 1243.5000 127.8000 1251.9000 ;
	    RECT 130.5000 1251.6000 136.8000 1252.8000 ;
	    RECT 143.4000 1252.5000 144.6000 1259.7001 ;
	    RECT 145.8000 1253.7001 147.0000 1259.7001 ;
	    RECT 148.2000 1252.5000 149.4000 1259.7001 ;
	    RECT 150.6000 1253.7001 151.8000 1259.7001 ;
	    RECT 130.5000 1251.0000 131.4000 1251.6000 ;
	    RECT 129.0000 1249.8000 131.4000 1251.0000 ;
	    RECT 135.9000 1250.7001 144.6000 1251.6000 ;
	    RECT 132.9000 1249.8000 135.0000 1250.7001 ;
	    RECT 132.9000 1249.5000 142.2000 1249.8000 ;
	    RECT 134.1000 1248.9000 142.2000 1249.5000 ;
	    RECT 141.0000 1248.6000 142.2000 1248.9000 ;
	    RECT 143.7000 1249.5000 144.6000 1250.7001 ;
	    RECT 145.5000 1250.4000 149.4000 1251.6000 ;
	    RECT 153.0000 1250.4000 154.2000 1259.7001 ;
	    RECT 155.4000 1255.5000 156.6000 1259.7001 ;
	    RECT 157.8000 1255.5000 159.0000 1259.7001 ;
	    RECT 160.2000 1255.5000 161.4000 1259.7001 ;
	    RECT 162.6000 1253.7001 163.8000 1259.7001 ;
	    RECT 157.8000 1251.6000 164.1000 1252.8000 ;
	    RECT 165.0000 1251.6000 166.2000 1259.7001 ;
	    RECT 167.4000 1253.7001 168.6000 1259.7001 ;
	    RECT 169.8000 1252.8000 171.0000 1259.7001 ;
	    RECT 172.2000 1253.7001 173.4000 1259.7001 ;
	    RECT 169.8000 1251.9000 173.7000 1252.8000 ;
	    RECT 174.6000 1252.5000 175.8000 1259.7001 ;
	    RECT 177.0000 1253.7001 178.2000 1259.7001 ;
	    RECT 189.0000 1253.7001 190.2000 1259.7001 ;
	    RECT 165.0000 1250.4000 168.9000 1251.6000 ;
	    RECT 155.4000 1249.5000 156.6000 1249.8000 ;
	    RECT 143.7000 1248.6000 156.6000 1249.5000 ;
	    RECT 160.2000 1249.5000 161.4000 1249.8000 ;
	    RECT 172.8000 1249.5000 173.7000 1251.9000 ;
	    RECT 174.6000 1250.4000 175.8000 1251.6000 ;
	    RECT 160.2000 1248.6000 173.7000 1249.5000 ;
	    RECT 131.4000 1247.4000 132.6000 1248.6000 ;
	    RECT 136.5000 1247.7001 137.7000 1248.0000 ;
	    RECT 133.5000 1246.8000 171.9000 1247.7001 ;
	    RECT 170.7000 1246.5000 171.9000 1246.8000 ;
	    RECT 172.8000 1245.9000 173.7000 1248.6000 ;
	    RECT 174.6000 1248.0000 175.8000 1249.5000 ;
	    RECT 174.6000 1246.8000 176.1000 1248.0000 ;
	    RECT 128.7000 1245.0000 135.3000 1245.9000 ;
	    RECT 128.7000 1244.7001 129.9000 1245.0000 ;
	    RECT 136.2000 1244.4000 137.4000 1245.6000 ;
	    RECT 138.3000 1245.0000 163.8000 1245.9000 ;
	    RECT 172.8000 1245.0000 174.0000 1245.9000 ;
	    RECT 162.6000 1244.1000 163.8000 1245.0000 ;
	    RECT 126.6000 1242.3000 139.8000 1243.5000 ;
	    RECT 140.7000 1242.9000 143.7000 1244.1000 ;
	    RECT 149.4000 1242.9000 154.2000 1244.1000 ;
	    RECT 126.6000 1233.3000 127.8000 1242.3000 ;
	    RECT 130.2000 1240.2001 134.7000 1241.4000 ;
	    RECT 133.5000 1239.3000 134.7000 1240.2001 ;
	    RECT 142.5000 1239.3000 143.7000 1242.9000 ;
	    RECT 145.8000 1241.4000 147.0000 1242.6000 ;
	    RECT 153.6000 1241.7001 154.8000 1242.0000 ;
	    RECT 148.2000 1240.8000 154.8000 1241.7001 ;
	    RECT 148.2000 1240.5000 149.4000 1240.8000 ;
	    RECT 145.8000 1240.2001 147.0000 1240.5000 ;
	    RECT 157.8000 1239.6000 159.0000 1243.8000 ;
	    RECT 166.5000 1242.9000 172.2000 1244.1000 ;
	    RECT 166.5000 1241.1000 167.7000 1242.9000 ;
	    RECT 173.1000 1242.0000 174.0000 1245.0000 ;
	    RECT 148.2000 1239.3000 149.4000 1239.6000 ;
	    RECT 131.4000 1233.3000 132.6000 1239.3000 ;
	    RECT 133.5000 1238.1000 137.4000 1239.3000 ;
	    RECT 142.5000 1238.4000 149.4000 1239.3000 ;
	    RECT 150.6000 1238.4000 151.8000 1239.6000 ;
	    RECT 152.7000 1238.4000 153.0000 1239.6000 ;
	    RECT 157.5000 1238.4000 159.0000 1239.6000 ;
	    RECT 165.0000 1240.2001 167.7000 1241.1000 ;
	    RECT 172.2000 1241.1000 174.0000 1242.0000 ;
	    RECT 165.0000 1239.3000 166.2000 1240.2001 ;
	    RECT 136.2000 1233.3000 137.4000 1238.1000 ;
	    RECT 162.6000 1238.1000 166.2000 1239.3000 ;
	    RECT 138.6000 1233.3000 139.8000 1237.5000 ;
	    RECT 141.0000 1233.3000 142.2000 1237.5000 ;
	    RECT 143.4000 1233.3000 144.6000 1237.5000 ;
	    RECT 145.8000 1233.3000 147.0000 1236.3000 ;
	    RECT 148.2000 1233.3000 149.4000 1237.5000 ;
	    RECT 150.6000 1233.3000 151.8000 1236.3000 ;
	    RECT 153.0000 1233.3000 154.2000 1237.5000 ;
	    RECT 155.4000 1233.3000 156.6000 1237.5000 ;
	    RECT 157.8000 1233.3000 159.0000 1237.5000 ;
	    RECT 160.2000 1233.3000 161.4000 1237.5000 ;
	    RECT 162.6000 1233.3000 163.8000 1238.1000 ;
	    RECT 167.4000 1233.3000 168.6000 1239.3000 ;
	    RECT 172.2000 1233.3000 173.4000 1241.1000 ;
	    RECT 174.9000 1240.2001 176.1000 1246.8000 ;
	    RECT 191.4000 1243.5000 192.6000 1259.7001 ;
	    RECT 323.4000 1253.7001 324.6000 1259.7001 ;
	    RECT 325.8000 1252.5000 327.0000 1259.7001 ;
	    RECT 328.2000 1253.7001 329.4000 1259.7001 ;
	    RECT 330.6000 1252.8000 331.8000 1259.7001 ;
	    RECT 333.0000 1253.7001 334.2000 1259.7001 ;
	    RECT 327.9000 1251.9000 331.8000 1252.8000 ;
	    RECT 311.4000 1251.4501 312.6000 1251.6000 ;
	    RECT 325.8000 1251.4501 327.0000 1251.6000 ;
	    RECT 311.4000 1250.5500 327.0000 1251.4501 ;
	    RECT 311.4000 1250.4000 312.6000 1250.5500 ;
	    RECT 325.8000 1250.4000 327.0000 1250.5500 ;
	    RECT 327.9000 1249.5000 328.8000 1251.9000 ;
	    RECT 335.4000 1251.6000 336.6000 1259.7001 ;
	    RECT 337.8000 1253.7001 339.0000 1259.7001 ;
	    RECT 340.2000 1255.5000 341.4000 1259.7001 ;
	    RECT 342.6000 1255.5000 343.8000 1259.7001 ;
	    RECT 345.0000 1255.5000 346.2000 1259.7001 ;
	    RECT 337.5000 1251.6000 343.8000 1252.8000 ;
	    RECT 332.7000 1250.4000 336.6000 1251.6000 ;
	    RECT 347.4000 1250.4000 348.6000 1259.7001 ;
	    RECT 349.8000 1253.7001 351.0000 1259.7001 ;
	    RECT 352.2000 1252.5000 353.4000 1259.7001 ;
	    RECT 354.6000 1253.7001 355.8000 1259.7001 ;
	    RECT 357.0000 1252.5000 358.2000 1259.7001 ;
	    RECT 359.4000 1255.5000 360.6000 1259.7001 ;
	    RECT 361.8000 1255.5000 363.0000 1259.7001 ;
	    RECT 364.2000 1253.7001 365.4000 1259.7001 ;
	    RECT 366.6000 1252.8000 367.8000 1259.7001 ;
	    RECT 369.0000 1253.7001 370.2000 1260.6000 ;
	    RECT 371.4000 1254.6000 372.6000 1259.7001 ;
	    RECT 371.4000 1253.7001 372.9000 1254.6000 ;
	    RECT 373.8000 1253.7001 375.0000 1259.7001 ;
	    RECT 372.0000 1252.8000 372.9000 1253.7001 ;
	    RECT 364.8000 1251.6000 371.1000 1252.8000 ;
	    RECT 372.0000 1251.9000 375.0000 1252.8000 ;
	    RECT 352.2000 1250.4000 356.1000 1251.6000 ;
	    RECT 357.0000 1250.7001 365.7000 1251.6000 ;
	    RECT 370.2000 1251.0000 371.1000 1251.6000 ;
	    RECT 340.2000 1249.5000 341.4000 1249.8000 ;
	    RECT 325.8000 1248.0000 327.0000 1249.5000 ;
	    RECT 325.5000 1246.8000 327.0000 1248.0000 ;
	    RECT 327.9000 1248.6000 341.4000 1249.5000 ;
	    RECT 345.0000 1249.5000 346.2000 1249.8000 ;
	    RECT 357.0000 1249.5000 357.9000 1250.7001 ;
	    RECT 366.6000 1249.8000 368.7000 1250.7001 ;
	    RECT 370.2000 1249.8000 372.6000 1251.0000 ;
	    RECT 345.0000 1248.6000 357.9000 1249.5000 ;
	    RECT 359.4000 1249.5000 368.7000 1249.8000 ;
	    RECT 359.4000 1248.9000 367.5000 1249.5000 ;
	    RECT 359.4000 1248.6000 360.6000 1248.9000 ;
	    RECT 191.4000 1242.4501 192.6000 1242.6000 ;
	    RECT 253.8000 1242.4501 255.0000 1242.6000 ;
	    RECT 191.4000 1241.5500 255.0000 1242.4501 ;
	    RECT 191.4000 1241.4000 192.6000 1241.5500 ;
	    RECT 253.8000 1241.4000 255.0000 1241.5500 ;
	    RECT 174.6000 1239.0000 176.1000 1240.2001 ;
	    RECT 179.4000 1239.4501 180.6000 1239.6000 ;
	    RECT 189.0000 1239.4501 190.2000 1239.6000 ;
	    RECT 174.6000 1233.3000 175.8000 1239.0000 ;
	    RECT 179.4000 1238.5500 190.2000 1239.4501 ;
	    RECT 179.4000 1238.4000 180.6000 1238.5500 ;
	    RECT 189.0000 1238.4000 190.2000 1238.5500 ;
	    RECT 189.0000 1237.2001 190.2000 1237.5000 ;
	    RECT 177.0000 1233.3000 178.2000 1236.3000 ;
	    RECT 189.0000 1233.3000 190.2000 1236.3000 ;
	    RECT 191.4000 1233.3000 192.6000 1240.5000 ;
	    RECT 325.5000 1240.2001 326.7000 1246.8000 ;
	    RECT 327.9000 1245.9000 328.8000 1248.6000 ;
	    RECT 363.9000 1247.7001 365.1000 1248.0000 ;
	    RECT 329.7000 1246.8000 368.1000 1247.7001 ;
	    RECT 369.0000 1247.4000 370.2000 1248.6000 ;
	    RECT 329.7000 1246.5000 330.9000 1246.8000 ;
	    RECT 327.6000 1245.0000 328.8000 1245.9000 ;
	    RECT 337.8000 1245.0000 363.3000 1245.9000 ;
	    RECT 327.6000 1242.0000 328.5000 1245.0000 ;
	    RECT 337.8000 1244.1000 339.0000 1245.0000 ;
	    RECT 364.2000 1244.4000 365.4000 1245.6000 ;
	    RECT 366.3000 1245.0000 372.9000 1245.9000 ;
	    RECT 371.7000 1244.7001 372.9000 1245.0000 ;
	    RECT 329.4000 1242.9000 335.1000 1244.1000 ;
	    RECT 327.6000 1241.1000 329.4000 1242.0000 ;
	    RECT 325.5000 1239.0000 327.0000 1240.2001 ;
	    RECT 323.4000 1233.3000 324.6000 1236.3000 ;
	    RECT 325.8000 1233.3000 327.0000 1239.0000 ;
	    RECT 328.2000 1233.3000 329.4000 1241.1000 ;
	    RECT 333.9000 1241.1000 335.1000 1242.9000 ;
	    RECT 333.9000 1240.2001 336.6000 1241.1000 ;
	    RECT 335.4000 1239.3000 336.6000 1240.2001 ;
	    RECT 342.6000 1239.6000 343.8000 1243.8000 ;
	    RECT 347.4000 1242.9000 352.2000 1244.1000 ;
	    RECT 357.9000 1242.9000 360.9000 1244.1000 ;
	    RECT 373.8000 1243.5000 375.0000 1251.9000 ;
	    RECT 397.8000 1248.6000 399.0000 1259.7001 ;
	    RECT 400.2000 1249.5000 401.4000 1259.7001 ;
	    RECT 402.6000 1248.6000 403.8000 1259.7001 ;
	    RECT 397.8000 1247.7001 403.8000 1248.6000 ;
	    RECT 405.0000 1247.7001 406.2000 1259.7001 ;
	    RECT 419.4000 1253.7001 420.6000 1259.7001 ;
	    RECT 405.0000 1246.5000 405.9000 1247.7001 ;
	    RECT 393.0000 1245.4501 394.2000 1245.6000 ;
	    RECT 397.8000 1245.4501 399.0000 1245.6000 ;
	    RECT 393.0000 1244.5500 399.0000 1245.4501 ;
	    RECT 399.9000 1244.7001 400.2000 1246.2001 ;
	    RECT 402.6000 1244.7001 404.1000 1245.6000 ;
	    RECT 405.0000 1245.4501 406.2000 1245.6000 ;
	    RECT 419.4000 1245.4501 420.6000 1245.6000 ;
	    RECT 393.0000 1244.4000 394.2000 1244.5500 ;
	    RECT 397.8000 1244.4000 399.0000 1244.5500 ;
	    RECT 400.2000 1243.5000 401.4000 1243.8000 ;
	    RECT 346.8000 1241.7001 348.0000 1242.0000 ;
	    RECT 346.8000 1240.8000 353.4000 1241.7001 ;
	    RECT 354.6000 1241.4000 355.8000 1242.6000 ;
	    RECT 352.2000 1240.5000 353.4000 1240.8000 ;
	    RECT 354.6000 1240.2001 355.8000 1240.5000 ;
	    RECT 333.0000 1233.3000 334.2000 1239.3000 ;
	    RECT 335.4000 1238.1000 339.0000 1239.3000 ;
	    RECT 342.6000 1238.4000 344.1000 1239.6000 ;
	    RECT 348.6000 1238.4000 348.9000 1239.6000 ;
	    RECT 349.8000 1238.4000 351.0000 1239.6000 ;
	    RECT 352.2000 1239.3000 353.4000 1239.6000 ;
	    RECT 357.9000 1239.3000 359.1000 1242.9000 ;
	    RECT 361.8000 1242.3000 375.0000 1243.5000 ;
	    RECT 366.9000 1240.2001 371.4000 1241.4000 ;
	    RECT 366.9000 1239.3000 368.1000 1240.2001 ;
	    RECT 352.2000 1238.4000 359.1000 1239.3000 ;
	    RECT 337.8000 1233.3000 339.0000 1238.1000 ;
	    RECT 364.2000 1238.1000 368.1000 1239.3000 ;
	    RECT 340.2000 1233.3000 341.4000 1237.5000 ;
	    RECT 342.6000 1233.3000 343.8000 1237.5000 ;
	    RECT 345.0000 1233.3000 346.2000 1237.5000 ;
	    RECT 347.4000 1233.3000 348.6000 1237.5000 ;
	    RECT 349.8000 1233.3000 351.0000 1236.3000 ;
	    RECT 352.2000 1233.3000 353.4000 1237.5000 ;
	    RECT 354.6000 1233.3000 355.8000 1236.3000 ;
	    RECT 357.0000 1233.3000 358.2000 1237.5000 ;
	    RECT 359.4000 1233.3000 360.6000 1237.5000 ;
	    RECT 361.8000 1233.3000 363.0000 1237.5000 ;
	    RECT 364.2000 1233.3000 365.4000 1238.1000 ;
	    RECT 369.0000 1233.3000 370.2000 1239.3000 ;
	    RECT 373.8000 1233.3000 375.0000 1242.3000 ;
	    RECT 400.2000 1241.4000 401.4000 1242.6000 ;
	    RECT 402.6000 1239.3000 403.5000 1244.7001 ;
	    RECT 405.0000 1244.5500 420.6000 1245.4501 ;
	    RECT 405.0000 1244.4000 406.2000 1244.5500 ;
	    RECT 419.4000 1244.4000 420.6000 1244.5500 ;
	    RECT 421.8000 1243.5000 423.0000 1259.7001 ;
	    RECT 453.0000 1247.7001 454.2000 1259.7001 ;
	    RECT 456.9000 1248.6000 458.1000 1259.7001 ;
	    RECT 459.3000 1253.7001 460.5000 1259.7001 ;
	    RECT 479.4000 1253.7001 480.6000 1259.7001 ;
	    RECT 459.0000 1250.4000 460.2000 1251.6000 ;
	    RECT 459.3000 1249.5000 460.2000 1250.4000 ;
	    RECT 479.4000 1249.5000 480.6000 1249.8000 ;
	    RECT 456.9000 1247.7001 458.4000 1248.6000 ;
	    RECT 455.4000 1245.4501 456.6000 1245.6000 ;
	    RECT 450.7500 1244.5500 456.6000 1245.4501 ;
	    RECT 421.8000 1242.4501 423.0000 1242.6000 ;
	    RECT 450.7500 1242.4501 451.6500 1244.5500 ;
	    RECT 455.4000 1244.4000 456.6000 1244.5500 ;
	    RECT 455.4000 1243.2001 456.6000 1243.5000 ;
	    RECT 457.5000 1242.6000 458.4000 1247.7001 ;
	    RECT 460.2000 1247.4000 461.4000 1248.6000 ;
	    RECT 479.4000 1247.4000 480.6000 1248.6000 ;
	    RECT 460.3500 1245.4501 461.2500 1247.4000 ;
	    RECT 481.8000 1246.5000 483.0000 1259.7001 ;
	    RECT 484.2000 1253.7001 485.4000 1259.7001 ;
	    RECT 611.4000 1253.7001 612.6000 1259.7001 ;
	    RECT 613.8000 1252.5000 615.0000 1259.7001 ;
	    RECT 616.2000 1253.7001 617.4000 1259.7001 ;
	    RECT 618.6000 1252.8000 619.8000 1259.7001 ;
	    RECT 621.0000 1253.7001 622.2000 1259.7001 ;
	    RECT 615.9000 1251.9000 619.8000 1252.8000 ;
	    RECT 613.8000 1250.4000 615.0000 1251.6000 ;
	    RECT 615.9000 1249.5000 616.8000 1251.9000 ;
	    RECT 623.4000 1251.6000 624.6000 1259.7001 ;
	    RECT 625.8000 1253.7001 627.0000 1259.7001 ;
	    RECT 628.2000 1255.5000 629.4000 1259.7001 ;
	    RECT 630.6000 1255.5000 631.8000 1259.7001 ;
	    RECT 633.0000 1255.5000 634.2000 1259.7001 ;
	    RECT 625.5000 1251.6000 631.8000 1252.8000 ;
	    RECT 620.7000 1250.4000 624.6000 1251.6000 ;
	    RECT 635.4000 1250.4000 636.6000 1259.7001 ;
	    RECT 637.8000 1253.7001 639.0000 1259.7001 ;
	    RECT 640.2000 1252.5000 641.4000 1259.7001 ;
	    RECT 642.6000 1253.7001 643.8000 1259.7001 ;
	    RECT 645.0000 1252.5000 646.2000 1259.7001 ;
	    RECT 647.4000 1255.5000 648.6000 1259.7001 ;
	    RECT 649.8000 1255.5000 651.0000 1259.7001 ;
	    RECT 652.2000 1253.7001 653.4000 1259.7001 ;
	    RECT 654.6000 1252.8000 655.8000 1259.7001 ;
	    RECT 657.0000 1253.7001 658.2000 1260.6000 ;
	    RECT 659.4000 1254.6000 660.6000 1259.7001 ;
	    RECT 659.4000 1253.7001 660.9000 1254.6000 ;
	    RECT 661.8000 1253.7001 663.0000 1259.7001 ;
	    RECT 693.9000 1253.7001 695.1000 1259.7001 ;
	    RECT 660.0000 1252.8000 660.9000 1253.7001 ;
	    RECT 652.8000 1251.6000 659.1000 1252.8000 ;
	    RECT 660.0000 1251.9000 663.0000 1252.8000 ;
	    RECT 640.2000 1250.4000 644.1000 1251.6000 ;
	    RECT 645.0000 1250.7001 653.7000 1251.6000 ;
	    RECT 658.2000 1251.0000 659.1000 1251.6000 ;
	    RECT 628.2000 1249.5000 629.4000 1249.8000 ;
	    RECT 613.8000 1248.0000 615.0000 1249.5000 ;
	    RECT 613.5000 1246.8000 615.0000 1248.0000 ;
	    RECT 615.9000 1248.6000 629.4000 1249.5000 ;
	    RECT 633.0000 1249.5000 634.2000 1249.8000 ;
	    RECT 645.0000 1249.5000 645.9000 1250.7001 ;
	    RECT 654.6000 1249.8000 656.7000 1250.7001 ;
	    RECT 658.2000 1249.8000 660.6000 1251.0000 ;
	    RECT 633.0000 1248.6000 645.9000 1249.5000 ;
	    RECT 647.4000 1249.5000 656.7000 1249.8000 ;
	    RECT 647.4000 1248.9000 655.5000 1249.5000 ;
	    RECT 647.4000 1248.6000 648.6000 1248.9000 ;
	    RECT 481.8000 1245.4501 483.0000 1245.6000 ;
	    RECT 460.3500 1244.5500 483.0000 1245.4501 ;
	    RECT 481.8000 1244.4000 483.0000 1244.5500 ;
	    RECT 421.8000 1241.5500 451.6500 1242.4501 ;
	    RECT 421.8000 1241.4000 423.0000 1241.5500 ;
	    RECT 453.0000 1241.4000 454.2000 1242.6000 ;
	    RECT 455.1000 1240.8000 455.4000 1242.3000 ;
	    RECT 457.5000 1241.4000 459.3000 1242.6000 ;
	    RECT 460.2000 1242.4501 461.4000 1242.6000 ;
	    RECT 479.4000 1242.4501 480.6000 1242.6000 ;
	    RECT 460.2000 1241.5500 480.6000 1242.4501 ;
	    RECT 460.2000 1241.4000 461.4000 1241.5500 ;
	    RECT 479.4000 1241.4000 480.6000 1241.5500 ;
	    RECT 405.0000 1239.4501 406.2000 1239.6000 ;
	    RECT 407.4000 1239.4501 408.6000 1239.6000 ;
	    RECT 417.0000 1239.4501 418.2000 1239.6000 ;
	    RECT 398.7000 1233.3000 399.9000 1239.3000 ;
	    RECT 402.6000 1233.3000 403.8000 1239.3000 ;
	    RECT 405.0000 1238.5500 418.2000 1239.4501 ;
	    RECT 405.0000 1238.4000 406.2000 1238.5500 ;
	    RECT 407.4000 1238.4000 408.6000 1238.5500 ;
	    RECT 417.0000 1238.4000 418.2000 1238.5500 ;
	    RECT 419.4000 1238.4000 420.6000 1239.6000 ;
	    RECT 404.7000 1237.2001 405.9000 1237.5000 ;
	    RECT 419.4000 1237.2001 420.6000 1237.5000 ;
	    RECT 405.0000 1233.3000 406.2000 1236.3000 ;
	    RECT 419.4000 1233.3000 420.6000 1236.3000 ;
	    RECT 421.8000 1233.3000 423.0000 1240.5000 ;
	    RECT 453.3000 1239.3000 458.7000 1239.9000 ;
	    RECT 460.2000 1239.3000 461.1000 1240.5000 ;
	    RECT 481.8000 1239.3000 483.0000 1243.5000 ;
	    RECT 484.2000 1242.4501 485.4000 1242.6000 ;
	    RECT 611.4000 1242.4501 612.6000 1242.6000 ;
	    RECT 484.2000 1241.5500 612.6000 1242.4501 ;
	    RECT 484.2000 1241.4000 485.4000 1241.5500 ;
	    RECT 611.4000 1241.4000 612.6000 1241.5500 ;
	    RECT 484.2000 1240.2001 485.4000 1240.5000 ;
	    RECT 613.5000 1240.2001 614.7000 1246.8000 ;
	    RECT 615.9000 1245.9000 616.8000 1248.6000 ;
	    RECT 651.9000 1247.7001 653.1000 1248.0000 ;
	    RECT 617.7000 1246.8000 656.1000 1247.7001 ;
	    RECT 657.0000 1247.4000 658.2000 1248.6000 ;
	    RECT 617.7000 1246.5000 618.9000 1246.8000 ;
	    RECT 615.6000 1245.0000 616.8000 1245.9000 ;
	    RECT 625.8000 1245.0000 651.3000 1245.9000 ;
	    RECT 615.6000 1242.0000 616.5000 1245.0000 ;
	    RECT 625.8000 1244.1000 627.0000 1245.0000 ;
	    RECT 652.2000 1244.4000 653.4000 1245.6000 ;
	    RECT 654.3000 1245.0000 660.9000 1245.9000 ;
	    RECT 659.7000 1244.7001 660.9000 1245.0000 ;
	    RECT 617.4000 1242.9000 623.1000 1244.1000 ;
	    RECT 615.6000 1241.1000 617.4000 1242.0000 ;
	    RECT 453.0000 1239.0000 459.0000 1239.3000 ;
	    RECT 453.0000 1233.3000 454.2000 1239.0000 ;
	    RECT 455.4000 1233.3000 456.6000 1238.1000 ;
	    RECT 457.8000 1233.3000 459.0000 1239.0000 ;
	    RECT 460.2000 1233.3000 461.4000 1239.3000 ;
	    RECT 480.3000 1238.4000 483.0000 1239.3000 ;
	    RECT 480.3000 1233.3000 481.5000 1238.4000 ;
	    RECT 484.2000 1233.3000 485.4000 1239.3000 ;
	    RECT 613.5000 1239.0000 615.0000 1240.2001 ;
	    RECT 611.4000 1233.3000 612.6000 1236.3000 ;
	    RECT 613.8000 1233.3000 615.0000 1239.0000 ;
	    RECT 616.2000 1233.3000 617.4000 1241.1000 ;
	    RECT 621.9000 1241.1000 623.1000 1242.9000 ;
	    RECT 621.9000 1240.2001 624.6000 1241.1000 ;
	    RECT 623.4000 1239.3000 624.6000 1240.2001 ;
	    RECT 630.6000 1239.6000 631.8000 1243.8000 ;
	    RECT 635.4000 1242.9000 640.2000 1244.1000 ;
	    RECT 645.9000 1242.9000 648.9000 1244.1000 ;
	    RECT 661.8000 1243.5000 663.0000 1251.9000 ;
	    RECT 694.2000 1250.4000 695.4000 1251.6000 ;
	    RECT 694.2000 1249.5000 695.1000 1250.4000 ;
	    RECT 696.3000 1248.6000 697.5000 1259.7001 ;
	    RECT 690.6000 1248.4501 691.8000 1248.6000 ;
	    RECT 693.0000 1248.4501 694.2000 1248.6000 ;
	    RECT 690.6000 1247.5500 694.2000 1248.4501 ;
	    RECT 690.6000 1247.4000 691.8000 1247.5500 ;
	    RECT 693.0000 1247.4000 694.2000 1247.5500 ;
	    RECT 696.0000 1247.7001 697.5000 1248.6000 ;
	    RECT 700.2000 1247.7001 701.4000 1259.7001 ;
	    RECT 719.4000 1253.7001 720.6000 1259.7001 ;
	    RECT 634.8000 1241.7001 636.0000 1242.0000 ;
	    RECT 634.8000 1240.8000 641.4000 1241.7001 ;
	    RECT 642.6000 1241.4000 643.8000 1242.6000 ;
	    RECT 640.2000 1240.5000 641.4000 1240.8000 ;
	    RECT 642.6000 1240.2001 643.8000 1240.5000 ;
	    RECT 621.0000 1233.3000 622.2000 1239.3000 ;
	    RECT 623.4000 1238.1000 627.0000 1239.3000 ;
	    RECT 630.6000 1238.4000 632.1000 1239.6000 ;
	    RECT 636.6000 1238.4000 636.9000 1239.6000 ;
	    RECT 637.8000 1238.4000 639.0000 1239.6000 ;
	    RECT 640.2000 1239.3000 641.4000 1239.6000 ;
	    RECT 645.9000 1239.3000 647.1000 1242.9000 ;
	    RECT 649.8000 1242.3000 663.0000 1243.5000 ;
	    RECT 696.0000 1242.6000 696.9000 1247.7001 ;
	    RECT 721.8000 1246.5000 723.0000 1259.7001 ;
	    RECT 724.2000 1253.7001 725.4000 1259.7001 ;
	    RECT 724.2000 1249.5000 725.4000 1249.8000 ;
	    RECT 724.2000 1248.4501 725.4000 1248.6000 ;
	    RECT 731.4000 1248.4501 732.6000 1248.6000 ;
	    RECT 724.2000 1247.5500 732.6000 1248.4501 ;
	    RECT 748.2000 1247.7001 749.4000 1259.7001 ;
	    RECT 752.1000 1248.6000 753.3000 1259.7001 ;
	    RECT 754.5000 1253.7001 755.7000 1259.7001 ;
	    RECT 754.2000 1250.4000 755.4000 1251.6000 ;
	    RECT 754.5000 1249.5000 755.4000 1250.4000 ;
	    RECT 752.1000 1247.7001 753.6000 1248.6000 ;
	    RECT 724.2000 1247.4000 725.4000 1247.5500 ;
	    RECT 731.4000 1247.4000 732.6000 1247.5500 ;
	    RECT 697.8000 1244.4000 699.0000 1245.6000 ;
	    RECT 700.2000 1245.4501 701.4000 1245.6000 ;
	    RECT 721.8000 1245.4501 723.0000 1245.6000 ;
	    RECT 745.8000 1245.4501 747.0000 1245.6000 ;
	    RECT 700.2000 1244.5500 703.6500 1245.4501 ;
	    RECT 700.2000 1244.4000 701.4000 1244.5500 ;
	    RECT 697.8000 1243.2001 699.0000 1243.5000 ;
	    RECT 654.9000 1240.2001 659.4000 1241.4000 ;
	    RECT 654.9000 1239.3000 656.1000 1240.2001 ;
	    RECT 640.2000 1238.4000 647.1000 1239.3000 ;
	    RECT 625.8000 1233.3000 627.0000 1238.1000 ;
	    RECT 652.2000 1238.1000 656.1000 1239.3000 ;
	    RECT 628.2000 1233.3000 629.4000 1237.5000 ;
	    RECT 630.6000 1233.3000 631.8000 1237.5000 ;
	    RECT 633.0000 1233.3000 634.2000 1237.5000 ;
	    RECT 635.4000 1233.3000 636.6000 1237.5000 ;
	    RECT 637.8000 1233.3000 639.0000 1236.3000 ;
	    RECT 640.2000 1233.3000 641.4000 1237.5000 ;
	    RECT 642.6000 1233.3000 643.8000 1236.3000 ;
	    RECT 645.0000 1233.3000 646.2000 1237.5000 ;
	    RECT 647.4000 1233.3000 648.6000 1237.5000 ;
	    RECT 649.8000 1233.3000 651.0000 1237.5000 ;
	    RECT 652.2000 1233.3000 653.4000 1238.1000 ;
	    RECT 657.0000 1233.3000 658.2000 1239.3000 ;
	    RECT 661.8000 1233.3000 663.0000 1242.3000 ;
	    RECT 693.0000 1241.4000 694.2000 1242.6000 ;
	    RECT 695.1000 1241.4000 696.9000 1242.6000 ;
	    RECT 699.0000 1240.8000 699.3000 1242.3000 ;
	    RECT 700.2000 1241.4000 701.4000 1242.6000 ;
	    RECT 702.7500 1242.4501 703.6500 1244.5500 ;
	    RECT 721.8000 1244.5500 747.0000 1245.4501 ;
	    RECT 721.8000 1244.4000 723.0000 1244.5500 ;
	    RECT 745.8000 1244.4000 747.0000 1244.5500 ;
	    RECT 750.6000 1244.4000 751.8000 1245.6000 ;
	    RECT 719.4000 1242.4501 720.6000 1242.6000 ;
	    RECT 702.7500 1241.5500 720.6000 1242.4501 ;
	    RECT 719.4000 1241.4000 720.6000 1241.5500 ;
	    RECT 693.3000 1239.3000 694.2000 1240.5000 ;
	    RECT 719.4000 1240.2001 720.6000 1240.5000 ;
	    RECT 695.7000 1239.3000 701.1000 1239.9000 ;
	    RECT 721.8000 1239.3000 723.0000 1243.5000 ;
	    RECT 750.6000 1243.2001 751.8000 1243.5000 ;
	    RECT 752.7000 1242.6000 753.6000 1247.7001 ;
	    RECT 755.4000 1247.4000 756.6000 1248.6000 ;
	    RECT 769.8000 1243.5000 771.0000 1259.7001 ;
	    RECT 772.2000 1253.7001 773.4000 1259.7001 ;
	    RECT 803.4000 1247.7001 804.6000 1259.7001 ;
	    RECT 807.3000 1247.7001 810.3000 1259.7001 ;
	    RECT 813.0000 1247.7001 814.2000 1259.7001 ;
	    RECT 832.2000 1247.7001 833.4000 1259.7001 ;
	    RECT 836.1000 1248.9000 837.3000 1259.7001 ;
	    RECT 834.6000 1247.7001 837.3000 1248.9000 ;
	    RECT 868.2000 1247.7001 869.4000 1259.7001 ;
	    RECT 872.1000 1247.7001 875.1000 1259.7001 ;
	    RECT 877.8000 1247.7001 879.0000 1259.7001 ;
	    RECT 805.8000 1244.4000 807.0000 1245.6000 ;
	    RECT 803.4000 1243.5000 804.6000 1243.8000 ;
	    RECT 808.5000 1243.5000 809.4000 1247.7001 ;
	    RECT 810.6000 1245.4501 811.8000 1245.6000 ;
	    RECT 813.0000 1245.4501 814.2000 1245.6000 ;
	    RECT 810.6000 1244.5500 814.2000 1245.4501 ;
	    RECT 810.6000 1244.4000 811.8000 1244.5500 ;
	    RECT 813.0000 1244.4000 814.2000 1244.5500 ;
	    RECT 834.9000 1243.5000 835.8000 1247.7001 ;
	    RECT 837.0000 1246.5000 838.2000 1246.8000 ;
	    RECT 837.0000 1245.4501 838.2000 1245.6000 ;
	    RECT 865.8000 1245.4501 867.0000 1245.6000 ;
	    RECT 837.0000 1244.5500 867.0000 1245.4501 ;
	    RECT 837.0000 1244.4000 838.2000 1244.5500 ;
	    RECT 865.8000 1244.4000 867.0000 1244.5500 ;
	    RECT 870.6000 1244.4000 871.8000 1245.6000 ;
	    RECT 868.2000 1243.5000 869.4000 1243.8000 ;
	    RECT 873.3000 1243.5000 874.2000 1247.7001 ;
	    RECT 875.4000 1244.4000 876.6000 1245.6000 ;
	    RECT 877.8000 1245.4501 879.0000 1245.6000 ;
	    RECT 877.8000 1244.5500 881.2500 1245.4501 ;
	    RECT 877.8000 1244.4000 879.0000 1244.5500 ;
	    RECT 805.8000 1243.2001 807.0000 1243.5000 ;
	    RECT 810.6000 1243.2001 811.8000 1243.5000 ;
	    RECT 870.6000 1243.2001 871.8000 1243.5000 ;
	    RECT 875.4000 1243.2001 876.6000 1243.5000 ;
	    RECT 741.0000 1242.4501 742.2000 1242.6000 ;
	    RECT 748.2000 1242.4501 749.4000 1242.6000 ;
	    RECT 741.0000 1241.5500 749.4000 1242.4501 ;
	    RECT 741.0000 1241.4000 742.2000 1241.5500 ;
	    RECT 748.2000 1241.4000 749.4000 1241.5500 ;
	    RECT 750.3000 1240.8000 750.6000 1242.3000 ;
	    RECT 752.7000 1241.4000 754.5000 1242.6000 ;
	    RECT 755.4000 1241.4000 756.6000 1242.6000 ;
	    RECT 757.8000 1242.4501 759.0000 1242.6000 ;
	    RECT 769.8000 1242.4501 771.0000 1242.6000 ;
	    RECT 757.8000 1241.5500 771.0000 1242.4501 ;
	    RECT 757.8000 1241.4000 759.0000 1241.5500 ;
	    RECT 769.8000 1241.4000 771.0000 1241.5500 ;
	    RECT 803.4000 1241.4000 804.6000 1242.6000 ;
	    RECT 805.8000 1241.4000 807.3000 1242.3000 ;
	    RECT 808.2000 1241.4000 809.4000 1242.6000 ;
	    RECT 813.0000 1242.4501 814.2000 1242.6000 ;
	    RECT 815.4000 1242.4501 816.6000 1242.6000 ;
	    RECT 748.5000 1239.3000 753.9000 1239.9000 ;
	    RECT 755.4000 1239.3000 756.3000 1240.5000 ;
	    RECT 693.0000 1233.3000 694.2000 1239.3000 ;
	    RECT 695.4000 1239.0000 701.4000 1239.3000 ;
	    RECT 695.4000 1233.3000 696.6000 1239.0000 ;
	    RECT 697.8000 1233.3000 699.0000 1238.1000 ;
	    RECT 700.2000 1233.3000 701.4000 1239.0000 ;
	    RECT 719.4000 1233.3000 720.6000 1239.3000 ;
	    RECT 721.8000 1238.4000 724.5000 1239.3000 ;
	    RECT 723.3000 1233.3000 724.5000 1238.4000 ;
	    RECT 748.2000 1239.0000 754.2000 1239.3000 ;
	    RECT 748.2000 1233.3000 749.4000 1239.0000 ;
	    RECT 750.6000 1233.3000 751.8000 1238.1000 ;
	    RECT 753.0000 1233.3000 754.2000 1239.0000 ;
	    RECT 755.4000 1233.3000 756.6000 1239.3000 ;
	    RECT 769.8000 1233.3000 771.0000 1240.5000 ;
	    RECT 772.2000 1239.4501 773.4000 1239.6000 ;
	    RECT 777.0000 1239.4501 778.2000 1239.6000 ;
	    RECT 772.2000 1238.5500 778.2000 1239.4501 ;
	    RECT 805.8000 1239.3000 806.7000 1241.4000 ;
	    RECT 811.8000 1240.8000 812.1000 1242.3000 ;
	    RECT 813.0000 1241.5500 816.6000 1242.4501 ;
	    RECT 813.0000 1241.4000 814.2000 1241.5500 ;
	    RECT 815.4000 1241.4000 816.6000 1241.5500 ;
	    RECT 834.6000 1241.4000 835.8000 1242.6000 ;
	    RECT 868.2000 1241.4000 869.4000 1242.6000 ;
	    RECT 870.6000 1241.4000 872.1000 1242.3000 ;
	    RECT 873.0000 1241.4000 874.2000 1242.6000 ;
	    RECT 808.5000 1239.3000 813.9000 1239.9000 ;
	    RECT 772.2000 1238.4000 773.4000 1238.5500 ;
	    RECT 777.0000 1238.4000 778.2000 1238.5500 ;
	    RECT 772.2000 1237.2001 773.4000 1237.5000 ;
	    RECT 772.2000 1233.3000 773.4000 1236.3000 ;
	    RECT 803.4000 1234.2001 804.6000 1239.3000 ;
	    RECT 805.8000 1235.1000 807.0000 1239.3000 ;
	    RECT 808.2000 1239.0000 814.2000 1239.3000 ;
	    RECT 808.2000 1234.2001 809.4000 1239.0000 ;
	    RECT 803.4000 1233.3000 809.4000 1234.2001 ;
	    RECT 810.6000 1233.3000 811.8000 1238.1000 ;
	    RECT 813.0000 1233.3000 814.2000 1239.0000 ;
	    RECT 832.2000 1238.4000 833.4000 1239.6000 ;
	    RECT 832.2000 1237.2001 833.4000 1237.5000 ;
	    RECT 834.9000 1236.3000 835.8000 1240.5000 ;
	    RECT 870.6000 1239.3000 871.5000 1241.4000 ;
	    RECT 876.6000 1240.8000 876.9000 1242.3000 ;
	    RECT 877.8000 1241.4000 879.0000 1242.6000 ;
	    RECT 880.3500 1242.4501 881.2500 1244.5500 ;
	    RECT 889.8000 1243.5000 891.0000 1259.7001 ;
	    RECT 892.2000 1253.7001 893.4000 1259.7001 ;
	    RECT 913.8000 1243.5000 915.0000 1259.7001 ;
	    RECT 916.2000 1253.7001 917.4000 1259.7001 ;
	    RECT 947.4000 1247.7001 948.6000 1259.7001 ;
	    RECT 951.3000 1247.7001 954.3000 1259.7001 ;
	    RECT 957.0000 1247.7001 958.2000 1259.7001 ;
	    RECT 985.8000 1259.4000 987.0000 1260.6000 ;
	    RECT 959.4000 1257.4501 960.6000 1257.6000 ;
	    RECT 1055.4000 1257.4501 1056.6000 1257.6000 ;
	    RECT 959.4000 1256.5500 1056.6000 1257.4501 ;
	    RECT 959.4000 1256.4000 960.6000 1256.5500 ;
	    RECT 1055.4000 1256.4000 1056.6000 1256.5500 ;
	    RECT 997.8000 1254.4501 999.0000 1254.6000 ;
	    RECT 1069.8000 1254.4501 1071.0000 1254.6000 ;
	    RECT 997.8000 1253.5500 1071.0000 1254.4501 ;
	    RECT 1081.8000 1253.7001 1083.0000 1259.7001 ;
	    RECT 997.8000 1253.4000 999.0000 1253.5500 ;
	    RECT 1069.8000 1253.4000 1071.0000 1253.5500 ;
	    RECT 1084.2001 1252.5000 1085.4000 1259.7001 ;
	    RECT 1086.6000 1253.7001 1087.8000 1259.7001 ;
	    RECT 1089.0000 1252.8000 1090.2001 1259.7001 ;
	    RECT 1091.4000 1253.7001 1092.6000 1259.7001 ;
	    RECT 1086.3000 1251.9000 1090.2001 1252.8000 ;
	    RECT 1019.4000 1251.4501 1020.6000 1251.6000 ;
	    RECT 1084.2001 1251.4501 1085.4000 1251.6000 ;
	    RECT 1019.4000 1250.5500 1085.4000 1251.4501 ;
	    RECT 1019.4000 1250.4000 1020.6000 1250.5500 ;
	    RECT 1084.2001 1250.4000 1085.4000 1250.5500 ;
	    RECT 1086.3000 1249.5000 1087.2001 1251.9000 ;
	    RECT 1093.8000 1251.6000 1095.0000 1259.7001 ;
	    RECT 1096.2001 1253.7001 1097.4000 1259.7001 ;
	    RECT 1098.6000 1255.5000 1099.8000 1259.7001 ;
	    RECT 1101.0000 1255.5000 1102.2001 1259.7001 ;
	    RECT 1103.4000 1255.5000 1104.6000 1259.7001 ;
	    RECT 1095.9000 1251.6000 1102.2001 1252.8000 ;
	    RECT 1091.1000 1250.4000 1095.0000 1251.6000 ;
	    RECT 1105.8000 1250.4000 1107.0000 1259.7001 ;
	    RECT 1108.2001 1253.7001 1109.4000 1259.7001 ;
	    RECT 1110.6000 1252.5000 1111.8000 1259.7001 ;
	    RECT 1113.0000 1253.7001 1114.2001 1259.7001 ;
	    RECT 1115.4000 1252.5000 1116.6000 1259.7001 ;
	    RECT 1117.8000 1255.5000 1119.0000 1259.7001 ;
	    RECT 1120.2001 1255.5000 1121.4000 1259.7001 ;
	    RECT 1122.6000 1253.7001 1123.8000 1259.7001 ;
	    RECT 1125.0000 1252.8000 1126.2001 1259.7001 ;
	    RECT 1127.4000 1253.7001 1128.6000 1260.6000 ;
	    RECT 1129.8000 1254.6000 1131.0000 1259.7001 ;
	    RECT 1129.8000 1253.7001 1131.3000 1254.6000 ;
	    RECT 1132.2001 1253.7001 1133.4000 1259.7001 ;
	    RECT 1158.6000 1253.7001 1159.8000 1259.7001 ;
	    RECT 1130.4000 1252.8000 1131.3000 1253.7001 ;
	    RECT 1123.2001 1251.6000 1129.5000 1252.8000 ;
	    RECT 1130.4000 1251.9000 1133.4000 1252.8000 ;
	    RECT 1110.6000 1250.4000 1114.5000 1251.6000 ;
	    RECT 1115.4000 1250.7001 1124.1000 1251.6000 ;
	    RECT 1128.6000 1251.0000 1129.5000 1251.6000 ;
	    RECT 1098.6000 1249.5000 1099.8000 1249.8000 ;
	    RECT 1084.2001 1248.0000 1085.4000 1249.5000 ;
	    RECT 949.8000 1244.4000 951.0000 1245.6000 ;
	    RECT 947.4000 1243.5000 948.6000 1243.8000 ;
	    RECT 952.5000 1243.5000 953.4000 1247.7001 ;
	    RECT 1083.9000 1246.8000 1085.4000 1248.0000 ;
	    RECT 1086.3000 1248.6000 1099.8000 1249.5000 ;
	    RECT 1103.4000 1249.5000 1104.6000 1249.8000 ;
	    RECT 1115.4000 1249.5000 1116.3000 1250.7001 ;
	    RECT 1125.0000 1249.8000 1127.1000 1250.7001 ;
	    RECT 1128.6000 1249.8000 1131.0000 1251.0000 ;
	    RECT 1103.4000 1248.6000 1116.3000 1249.5000 ;
	    RECT 1117.8000 1249.5000 1127.1000 1249.8000 ;
	    RECT 1117.8000 1248.9000 1125.9000 1249.5000 ;
	    RECT 1117.8000 1248.6000 1119.0000 1248.9000 ;
	    RECT 954.6000 1244.4000 955.8000 1245.6000 ;
	    RECT 949.8000 1243.2001 951.0000 1243.5000 ;
	    RECT 954.6000 1243.2001 955.8000 1243.5000 ;
	    RECT 889.8000 1242.4501 891.0000 1242.6000 ;
	    RECT 880.3500 1241.5500 891.0000 1242.4501 ;
	    RECT 889.8000 1241.4000 891.0000 1241.5500 ;
	    RECT 892.2000 1242.4501 893.4000 1242.6000 ;
	    RECT 913.8000 1242.4501 915.0000 1242.6000 ;
	    RECT 892.2000 1241.5500 915.0000 1242.4501 ;
	    RECT 892.2000 1241.4000 893.4000 1241.5500 ;
	    RECT 913.8000 1241.4000 915.0000 1241.5500 ;
	    RECT 945.0000 1242.4501 946.2000 1242.6000 ;
	    RECT 947.4000 1242.4501 948.6000 1242.6000 ;
	    RECT 945.0000 1241.5500 948.6000 1242.4501 ;
	    RECT 945.0000 1241.4000 946.2000 1241.5500 ;
	    RECT 947.4000 1241.4000 948.6000 1241.5500 ;
	    RECT 949.8000 1241.4000 951.3000 1242.3000 ;
	    RECT 952.2000 1241.4000 953.4000 1242.6000 ;
	    RECT 873.3000 1239.3000 878.7000 1239.9000 ;
	    RECT 832.2000 1233.3000 833.4000 1236.3000 ;
	    RECT 834.6000 1233.3000 835.8000 1236.3000 ;
	    RECT 837.0000 1233.3000 838.2000 1236.3000 ;
	    RECT 868.2000 1234.2001 869.4000 1239.3000 ;
	    RECT 870.6000 1235.1000 871.8000 1239.3000 ;
	    RECT 873.0000 1239.0000 879.0000 1239.3000 ;
	    RECT 873.0000 1234.2001 874.2000 1239.0000 ;
	    RECT 868.2000 1233.3000 874.2000 1234.2001 ;
	    RECT 875.4000 1233.3000 876.6000 1238.1000 ;
	    RECT 877.8000 1233.3000 879.0000 1239.0000 ;
	    RECT 889.8000 1233.3000 891.0000 1240.5000 ;
	    RECT 892.2000 1239.4501 893.4000 1239.6000 ;
	    RECT 909.0000 1239.4501 910.2000 1239.6000 ;
	    RECT 892.2000 1238.5500 910.2000 1239.4501 ;
	    RECT 892.2000 1238.4000 893.4000 1238.5500 ;
	    RECT 909.0000 1238.4000 910.2000 1238.5500 ;
	    RECT 892.2000 1237.2001 893.4000 1237.5000 ;
	    RECT 892.2000 1233.3000 893.4000 1236.3000 ;
	    RECT 913.8000 1233.3000 915.0000 1240.5000 ;
	    RECT 916.2000 1239.4501 917.4000 1239.6000 ;
	    RECT 935.4000 1239.4501 936.6000 1239.6000 ;
	    RECT 916.2000 1238.5500 936.6000 1239.4501 ;
	    RECT 949.8000 1239.3000 950.7000 1241.4000 ;
	    RECT 955.8000 1240.8000 956.1000 1242.3000 ;
	    RECT 957.0000 1241.4000 958.2000 1242.6000 ;
	    RECT 1083.9000 1240.2001 1085.1000 1246.8000 ;
	    RECT 1086.3000 1245.9000 1087.2001 1248.6000 ;
	    RECT 1122.3000 1247.7001 1123.5000 1248.0000 ;
	    RECT 1088.1000 1246.8000 1126.5000 1247.7001 ;
	    RECT 1127.4000 1247.4000 1128.6000 1248.6000 ;
	    RECT 1088.1000 1246.5000 1089.3000 1246.8000 ;
	    RECT 1086.0000 1245.0000 1087.2001 1245.9000 ;
	    RECT 1096.2001 1245.0000 1121.7001 1245.9000 ;
	    RECT 1086.0000 1242.0000 1086.9000 1245.0000 ;
	    RECT 1096.2001 1244.1000 1097.4000 1245.0000 ;
	    RECT 1122.6000 1244.4000 1123.8000 1245.6000 ;
	    RECT 1124.7001 1245.0000 1131.3000 1245.9000 ;
	    RECT 1130.1000 1244.7001 1131.3000 1245.0000 ;
	    RECT 1087.8000 1242.9000 1093.5000 1244.1000 ;
	    RECT 1086.0000 1241.1000 1087.8000 1242.0000 ;
	    RECT 952.5000 1239.3000 957.9000 1239.9000 ;
	    RECT 916.2000 1238.4000 917.4000 1238.5500 ;
	    RECT 935.4000 1238.4000 936.6000 1238.5500 ;
	    RECT 916.2000 1237.2001 917.4000 1237.5000 ;
	    RECT 916.2000 1233.3000 917.4000 1236.3000 ;
	    RECT 947.4000 1234.2001 948.6000 1239.3000 ;
	    RECT 949.8000 1235.1000 951.0000 1239.3000 ;
	    RECT 952.2000 1239.0000 958.2000 1239.3000 ;
	    RECT 1083.9000 1239.0000 1085.4000 1240.2001 ;
	    RECT 952.2000 1234.2001 953.4000 1239.0000 ;
	    RECT 947.4000 1233.3000 953.4000 1234.2001 ;
	    RECT 954.6000 1233.3000 955.8000 1238.1000 ;
	    RECT 957.0000 1233.3000 958.2000 1239.0000 ;
	    RECT 959.4000 1236.4501 960.6000 1236.6000 ;
	    RECT 1017.0000 1236.4501 1018.2000 1236.6000 ;
	    RECT 959.4000 1235.5500 1018.2000 1236.4501 ;
	    RECT 959.4000 1235.4000 960.6000 1235.5500 ;
	    RECT 1017.0000 1235.4000 1018.2000 1235.5500 ;
	    RECT 1081.8000 1233.3000 1083.0000 1236.3000 ;
	    RECT 1084.2001 1233.3000 1085.4000 1239.0000 ;
	    RECT 1086.6000 1233.3000 1087.8000 1241.1000 ;
	    RECT 1092.3000 1241.1000 1093.5000 1242.9000 ;
	    RECT 1092.3000 1240.2001 1095.0000 1241.1000 ;
	    RECT 1093.8000 1239.3000 1095.0000 1240.2001 ;
	    RECT 1101.0000 1239.6000 1102.2001 1243.8000 ;
	    RECT 1105.8000 1242.9000 1110.6000 1244.1000 ;
	    RECT 1116.3000 1242.9000 1119.3000 1244.1000 ;
	    RECT 1132.2001 1243.5000 1133.4000 1251.9000 ;
	    RECT 1158.6000 1249.5000 1159.8000 1249.8000 ;
	    RECT 1144.2001 1248.4501 1145.4000 1248.6000 ;
	    RECT 1158.6000 1248.4501 1159.8000 1248.6000 ;
	    RECT 1144.2001 1247.5500 1159.8000 1248.4501 ;
	    RECT 1144.2001 1247.4000 1145.4000 1247.5500 ;
	    RECT 1158.6000 1247.4000 1159.8000 1247.5500 ;
	    RECT 1161.0000 1246.5000 1162.2001 1259.7001 ;
	    RECT 1163.4000 1253.7001 1164.6000 1259.7001 ;
	    RECT 1288.2001 1253.7001 1289.4000 1259.7001 ;
	    RECT 1290.6000 1252.5000 1291.8000 1259.7001 ;
	    RECT 1293.0000 1253.7001 1294.2001 1259.7001 ;
	    RECT 1295.4000 1252.8000 1296.6000 1259.7001 ;
	    RECT 1297.8000 1253.7001 1299.0000 1259.7001 ;
	    RECT 1292.7001 1251.9000 1296.6000 1252.8000 ;
	    RECT 1165.8000 1251.4501 1167.0000 1251.6000 ;
	    RECT 1273.8000 1251.4501 1275.0000 1251.6000 ;
	    RECT 1290.6000 1251.4501 1291.8000 1251.6000 ;
	    RECT 1165.8000 1250.5500 1291.8000 1251.4501 ;
	    RECT 1165.8000 1250.4000 1167.0000 1250.5500 ;
	    RECT 1273.8000 1250.4000 1275.0000 1250.5500 ;
	    RECT 1290.6000 1250.4000 1291.8000 1250.5500 ;
	    RECT 1292.7001 1249.5000 1293.6000 1251.9000 ;
	    RECT 1300.2001 1251.6000 1301.4000 1259.7001 ;
	    RECT 1302.6000 1253.7001 1303.8000 1259.7001 ;
	    RECT 1305.0000 1255.5000 1306.2001 1259.7001 ;
	    RECT 1307.4000 1255.5000 1308.6000 1259.7001 ;
	    RECT 1309.8000 1255.5000 1311.0000 1259.7001 ;
	    RECT 1302.3000 1251.6000 1308.6000 1252.8000 ;
	    RECT 1297.5000 1250.4000 1301.4000 1251.6000 ;
	    RECT 1312.2001 1250.4000 1313.4000 1259.7001 ;
	    RECT 1314.6000 1253.7001 1315.8000 1259.7001 ;
	    RECT 1317.0000 1252.5000 1318.2001 1259.7001 ;
	    RECT 1319.4000 1253.7001 1320.6000 1259.7001 ;
	    RECT 1321.8000 1252.5000 1323.0000 1259.7001 ;
	    RECT 1324.2001 1255.5000 1325.4000 1259.7001 ;
	    RECT 1326.6000 1255.5000 1327.8000 1259.7001 ;
	    RECT 1329.0000 1253.7001 1330.2001 1259.7001 ;
	    RECT 1331.4000 1252.8000 1332.6000 1259.7001 ;
	    RECT 1333.8000 1253.7001 1335.0000 1260.6000 ;
	    RECT 1336.2001 1254.6000 1337.4000 1259.7001 ;
	    RECT 1336.2001 1253.7001 1337.7001 1254.6000 ;
	    RECT 1338.6000 1253.7001 1339.8000 1259.7001 ;
	    RECT 1370.7001 1253.7001 1371.9000 1259.7001 ;
	    RECT 1336.8000 1252.8000 1337.7001 1253.7001 ;
	    RECT 1329.6000 1251.6000 1335.9000 1252.8000 ;
	    RECT 1336.8000 1251.9000 1339.8000 1252.8000 ;
	    RECT 1317.0000 1250.4000 1320.9000 1251.6000 ;
	    RECT 1321.8000 1250.7001 1330.5000 1251.6000 ;
	    RECT 1335.0000 1251.0000 1335.9000 1251.6000 ;
	    RECT 1305.0000 1249.5000 1306.2001 1249.8000 ;
	    RECT 1290.6000 1248.0000 1291.8000 1249.5000 ;
	    RECT 1290.3000 1246.8000 1291.8000 1248.0000 ;
	    RECT 1292.7001 1248.6000 1306.2001 1249.5000 ;
	    RECT 1309.8000 1249.5000 1311.0000 1249.8000 ;
	    RECT 1321.8000 1249.5000 1322.7001 1250.7001 ;
	    RECT 1331.4000 1249.8000 1333.5000 1250.7001 ;
	    RECT 1335.0000 1249.8000 1337.4000 1251.0000 ;
	    RECT 1309.8000 1248.6000 1322.7001 1249.5000 ;
	    RECT 1324.2001 1249.5000 1333.5000 1249.8000 ;
	    RECT 1324.2001 1248.9000 1332.3000 1249.5000 ;
	    RECT 1324.2001 1248.6000 1325.4000 1248.9000 ;
	    RECT 1134.6000 1245.4501 1135.8000 1245.6000 ;
	    RECT 1161.0000 1245.4501 1162.2001 1245.6000 ;
	    RECT 1134.6000 1244.5500 1162.2001 1245.4501 ;
	    RECT 1134.6000 1244.4000 1135.8000 1244.5500 ;
	    RECT 1161.0000 1244.4000 1162.2001 1244.5500 ;
	    RECT 1105.2001 1241.7001 1106.4000 1242.0000 ;
	    RECT 1105.2001 1240.8000 1111.8000 1241.7001 ;
	    RECT 1113.0000 1241.4000 1114.2001 1242.6000 ;
	    RECT 1110.6000 1240.5000 1111.8000 1240.8000 ;
	    RECT 1113.0000 1240.2001 1114.2001 1240.5000 ;
	    RECT 1091.4000 1233.3000 1092.6000 1239.3000 ;
	    RECT 1093.8000 1238.1000 1097.4000 1239.3000 ;
	    RECT 1101.0000 1238.4000 1102.5000 1239.6000 ;
	    RECT 1107.0000 1238.4000 1107.3000 1239.6000 ;
	    RECT 1108.2001 1238.4000 1109.4000 1239.6000 ;
	    RECT 1110.6000 1239.3000 1111.8000 1239.6000 ;
	    RECT 1116.3000 1239.3000 1117.5000 1242.9000 ;
	    RECT 1120.2001 1242.3000 1133.4000 1243.5000 ;
	    RECT 1125.3000 1240.2001 1129.8000 1241.4000 ;
	    RECT 1125.3000 1239.3000 1126.5000 1240.2001 ;
	    RECT 1110.6000 1238.4000 1117.5000 1239.3000 ;
	    RECT 1096.2001 1233.3000 1097.4000 1238.1000 ;
	    RECT 1122.6000 1238.1000 1126.5000 1239.3000 ;
	    RECT 1098.6000 1233.3000 1099.8000 1237.5000 ;
	    RECT 1101.0000 1233.3000 1102.2001 1237.5000 ;
	    RECT 1103.4000 1233.3000 1104.6000 1237.5000 ;
	    RECT 1105.8000 1233.3000 1107.0000 1237.5000 ;
	    RECT 1108.2001 1233.3000 1109.4000 1236.3000 ;
	    RECT 1110.6000 1233.3000 1111.8000 1237.5000 ;
	    RECT 1113.0000 1233.3000 1114.2001 1236.3000 ;
	    RECT 1115.4000 1233.3000 1116.6000 1237.5000 ;
	    RECT 1117.8000 1233.3000 1119.0000 1237.5000 ;
	    RECT 1120.2001 1233.3000 1121.4000 1237.5000 ;
	    RECT 1122.6000 1233.3000 1123.8000 1238.1000 ;
	    RECT 1127.4000 1233.3000 1128.6000 1239.3000 ;
	    RECT 1132.2001 1233.3000 1133.4000 1242.3000 ;
	    RECT 1161.0000 1239.3000 1162.2001 1243.5000 ;
	    RECT 1163.4000 1242.4501 1164.6000 1242.6000 ;
	    RECT 1213.8000 1242.4501 1215.0000 1242.6000 ;
	    RECT 1163.4000 1241.5500 1215.0000 1242.4501 ;
	    RECT 1163.4000 1241.4000 1164.6000 1241.5500 ;
	    RECT 1213.8000 1241.4000 1215.0000 1241.5500 ;
	    RECT 1163.4000 1240.2001 1164.6000 1240.5000 ;
	    RECT 1290.3000 1240.2001 1291.5000 1246.8000 ;
	    RECT 1292.7001 1245.9000 1293.6000 1248.6000 ;
	    RECT 1328.7001 1247.7001 1329.9000 1248.0000 ;
	    RECT 1294.5000 1246.8000 1332.9000 1247.7001 ;
	    RECT 1333.8000 1247.4000 1335.0000 1248.6000 ;
	    RECT 1294.5000 1246.5000 1295.7001 1246.8000 ;
	    RECT 1292.4000 1245.0000 1293.6000 1245.9000 ;
	    RECT 1302.6000 1245.0000 1328.1000 1245.9000 ;
	    RECT 1292.4000 1242.0000 1293.3000 1245.0000 ;
	    RECT 1302.6000 1244.1000 1303.8000 1245.0000 ;
	    RECT 1329.0000 1244.4000 1330.2001 1245.6000 ;
	    RECT 1331.1000 1245.0000 1337.7001 1245.9000 ;
	    RECT 1336.5000 1244.7001 1337.7001 1245.0000 ;
	    RECT 1294.2001 1242.9000 1299.9000 1244.1000 ;
	    RECT 1292.4000 1241.1000 1294.2001 1242.0000 ;
	    RECT 1159.5000 1238.4000 1162.2001 1239.3000 ;
	    RECT 1159.5000 1233.3000 1160.7001 1238.4000 ;
	    RECT 1163.4000 1233.3000 1164.6000 1239.3000 ;
	    RECT 1290.3000 1239.0000 1291.8000 1240.2001 ;
	    RECT 1288.2001 1233.3000 1289.4000 1236.3000 ;
	    RECT 1290.6000 1233.3000 1291.8000 1239.0000 ;
	    RECT 1293.0000 1233.3000 1294.2001 1241.1000 ;
	    RECT 1298.7001 1241.1000 1299.9000 1242.9000 ;
	    RECT 1298.7001 1240.2001 1301.4000 1241.1000 ;
	    RECT 1300.2001 1239.3000 1301.4000 1240.2001 ;
	    RECT 1307.4000 1239.6000 1308.6000 1243.8000 ;
	    RECT 1312.2001 1242.9000 1317.0000 1244.1000 ;
	    RECT 1322.7001 1242.9000 1325.7001 1244.1000 ;
	    RECT 1338.6000 1243.5000 1339.8000 1251.9000 ;
	    RECT 1371.0000 1250.4000 1372.2001 1251.6000 ;
	    RECT 1371.0000 1249.5000 1371.9000 1250.4000 ;
	    RECT 1373.1000 1248.6000 1374.3000 1259.7001 ;
	    RECT 1367.4000 1248.4501 1368.6000 1248.6000 ;
	    RECT 1369.8000 1248.4501 1371.0000 1248.6000 ;
	    RECT 1367.4000 1247.5500 1371.0000 1248.4501 ;
	    RECT 1367.4000 1247.4000 1368.6000 1247.5500 ;
	    RECT 1369.8000 1247.4000 1371.0000 1247.5500 ;
	    RECT 1372.8000 1247.7001 1374.3000 1248.6000 ;
	    RECT 1377.0000 1247.7001 1378.2001 1259.7001 ;
	    RECT 1391.4000 1253.7001 1392.6000 1259.7001 ;
	    RECT 1311.6000 1241.7001 1312.8000 1242.0000 ;
	    RECT 1311.6000 1240.8000 1318.2001 1241.7001 ;
	    RECT 1319.4000 1241.4000 1320.6000 1242.6000 ;
	    RECT 1317.0000 1240.5000 1318.2001 1240.8000 ;
	    RECT 1319.4000 1240.2001 1320.6000 1240.5000 ;
	    RECT 1297.8000 1233.3000 1299.0000 1239.3000 ;
	    RECT 1300.2001 1238.1000 1303.8000 1239.3000 ;
	    RECT 1307.4000 1238.4000 1308.9000 1239.6000 ;
	    RECT 1313.4000 1238.4000 1313.7001 1239.6000 ;
	    RECT 1314.6000 1238.4000 1315.8000 1239.6000 ;
	    RECT 1317.0000 1239.3000 1318.2001 1239.6000 ;
	    RECT 1322.7001 1239.3000 1323.9000 1242.9000 ;
	    RECT 1326.6000 1242.3000 1339.8000 1243.5000 ;
	    RECT 1372.8000 1242.6000 1373.7001 1247.7001 ;
	    RECT 1374.6000 1245.4501 1375.8000 1245.6000 ;
	    RECT 1374.6000 1244.5500 1380.4501 1245.4501 ;
	    RECT 1374.6000 1244.4000 1375.8000 1244.5500 ;
	    RECT 1374.6000 1243.2001 1375.8000 1243.5000 ;
	    RECT 1331.7001 1240.2001 1336.2001 1241.4000 ;
	    RECT 1331.7001 1239.3000 1332.9000 1240.2001 ;
	    RECT 1317.0000 1238.4000 1323.9000 1239.3000 ;
	    RECT 1302.6000 1233.3000 1303.8000 1238.1000 ;
	    RECT 1329.0000 1238.1000 1332.9000 1239.3000 ;
	    RECT 1305.0000 1233.3000 1306.2001 1237.5000 ;
	    RECT 1307.4000 1233.3000 1308.6000 1237.5000 ;
	    RECT 1309.8000 1233.3000 1311.0000 1237.5000 ;
	    RECT 1312.2001 1233.3000 1313.4000 1237.5000 ;
	    RECT 1314.6000 1233.3000 1315.8000 1236.3000 ;
	    RECT 1317.0000 1233.3000 1318.2001 1237.5000 ;
	    RECT 1319.4000 1233.3000 1320.6000 1236.3000 ;
	    RECT 1321.8000 1233.3000 1323.0000 1237.5000 ;
	    RECT 1324.2001 1233.3000 1325.4000 1237.5000 ;
	    RECT 1326.6000 1233.3000 1327.8000 1237.5000 ;
	    RECT 1329.0000 1233.3000 1330.2001 1238.1000 ;
	    RECT 1333.8000 1233.3000 1335.0000 1239.3000 ;
	    RECT 1338.6000 1233.3000 1339.8000 1242.3000 ;
	    RECT 1369.8000 1241.4000 1371.0000 1242.6000 ;
	    RECT 1371.9000 1241.4000 1373.7001 1242.6000 ;
	    RECT 1375.8000 1240.8000 1376.1000 1242.3000 ;
	    RECT 1377.0000 1241.4000 1378.2001 1242.6000 ;
	    RECT 1379.5500 1242.4501 1380.4501 1244.5500 ;
	    RECT 1393.8000 1243.5000 1395.0000 1259.7001 ;
	    RECT 1420.2001 1247.7001 1421.4000 1259.7001 ;
	    RECT 1424.1000 1248.6000 1425.3000 1259.7001 ;
	    RECT 1426.5000 1253.7001 1427.7001 1259.7001 ;
	    RECT 1452.3000 1253.7001 1453.5000 1259.7001 ;
	    RECT 1426.2001 1250.4000 1427.4000 1251.6000 ;
	    RECT 1426.5000 1249.5000 1427.4000 1250.4000 ;
	    RECT 1452.6000 1250.4000 1453.8000 1251.6000 ;
	    RECT 1452.6000 1249.5000 1453.5000 1250.4000 ;
	    RECT 1454.7001 1248.6000 1455.9000 1259.7001 ;
	    RECT 1424.1000 1247.7001 1425.6000 1248.6000 ;
	    RECT 1422.6000 1244.4000 1423.8000 1245.6000 ;
	    RECT 1422.6000 1243.2001 1423.8000 1243.5000 ;
	    RECT 1424.7001 1242.6000 1425.6000 1247.7001 ;
	    RECT 1427.4000 1247.4000 1428.6000 1248.6000 ;
	    RECT 1451.4000 1247.4000 1452.6000 1248.6000 ;
	    RECT 1454.4000 1247.7001 1455.9000 1248.6000 ;
	    RECT 1458.6000 1247.7001 1459.8000 1259.7001 ;
	    RECT 1477.8000 1253.7001 1479.0000 1259.7001 ;
	    RECT 1454.4000 1242.6000 1455.3000 1247.7001 ;
	    RECT 1480.2001 1246.5000 1481.4000 1259.7001 ;
	    RECT 1482.6000 1253.7001 1483.8000 1259.7001 ;
	    RECT 1507.5000 1253.7001 1508.7001 1259.7001 ;
	    RECT 1507.8000 1250.4000 1509.0000 1251.6000 ;
	    RECT 1482.6000 1249.5000 1483.8000 1249.8000 ;
	    RECT 1507.8000 1249.5000 1508.7001 1250.4000 ;
	    RECT 1509.9000 1248.6000 1511.1000 1259.7001 ;
	    RECT 1482.6000 1247.4000 1483.8000 1248.6000 ;
	    RECT 1506.6000 1247.4000 1507.8000 1248.6000 ;
	    RECT 1509.6000 1247.7001 1511.1000 1248.6000 ;
	    RECT 1513.8000 1247.7001 1515.0000 1259.7001 ;
	    RECT 1521.0000 1259.4000 1522.2001 1260.6000 ;
	    RECT 1456.2001 1245.4501 1457.4000 1245.6000 ;
	    RECT 1458.6000 1245.4501 1459.8000 1245.6000 ;
	    RECT 1456.2001 1244.5500 1459.8000 1245.4501 ;
	    RECT 1456.2001 1244.4000 1457.4000 1244.5500 ;
	    RECT 1458.6000 1244.4000 1459.8000 1244.5500 ;
	    RECT 1480.2001 1245.4501 1481.4000 1245.6000 ;
	    RECT 1506.7500 1245.4501 1507.6500 1247.4000 ;
	    RECT 1480.2001 1244.5500 1507.6500 1245.4501 ;
	    RECT 1480.2001 1244.4000 1481.4000 1244.5500 ;
	    RECT 1456.2001 1243.2001 1457.4000 1243.5000 ;
	    RECT 1393.8000 1242.4501 1395.0000 1242.6000 ;
	    RECT 1379.5500 1241.5500 1395.0000 1242.4501 ;
	    RECT 1393.8000 1241.4000 1395.0000 1241.5500 ;
	    RECT 1413.0000 1242.4501 1414.2001 1242.6000 ;
	    RECT 1420.2001 1242.4501 1421.4000 1242.6000 ;
	    RECT 1413.0000 1241.5500 1421.4000 1242.4501 ;
	    RECT 1413.0000 1241.4000 1414.2001 1241.5500 ;
	    RECT 1420.2001 1241.4000 1421.4000 1241.5500 ;
	    RECT 1422.3000 1240.8000 1422.6000 1242.3000 ;
	    RECT 1424.7001 1241.4000 1426.5000 1242.6000 ;
	    RECT 1427.4000 1242.4501 1428.6000 1242.6000 ;
	    RECT 1441.8000 1242.4501 1443.0000 1242.6000 ;
	    RECT 1427.4000 1241.5500 1443.0000 1242.4501 ;
	    RECT 1427.4000 1241.4000 1428.6000 1241.5500 ;
	    RECT 1441.8000 1241.4000 1443.0000 1241.5500 ;
	    RECT 1444.2001 1242.4501 1445.4000 1242.6000 ;
	    RECT 1451.4000 1242.4501 1452.6000 1242.6000 ;
	    RECT 1444.2001 1241.5500 1452.6000 1242.4501 ;
	    RECT 1444.2001 1241.4000 1445.4000 1241.5500 ;
	    RECT 1451.4000 1241.4000 1452.6000 1241.5500 ;
	    RECT 1453.5000 1241.4000 1455.3000 1242.6000 ;
	    RECT 1457.4000 1240.8000 1457.7001 1242.3000 ;
	    RECT 1458.6000 1241.4000 1459.8000 1242.6000 ;
	    RECT 1477.8000 1241.4000 1479.0000 1242.6000 ;
	    RECT 1370.1000 1239.3000 1371.0000 1240.5000 ;
	    RECT 1372.5000 1239.3000 1377.9000 1239.9000 ;
	    RECT 1369.8000 1233.3000 1371.0000 1239.3000 ;
	    RECT 1372.2001 1239.0000 1378.2001 1239.3000 ;
	    RECT 1372.2001 1233.3000 1373.4000 1239.0000 ;
	    RECT 1374.6000 1233.3000 1375.8000 1238.1000 ;
	    RECT 1377.0000 1233.3000 1378.2001 1239.0000 ;
	    RECT 1391.4000 1238.4000 1392.6000 1239.6000 ;
	    RECT 1391.4000 1237.2001 1392.6000 1237.5000 ;
	    RECT 1391.4000 1233.3000 1392.6000 1236.3000 ;
	    RECT 1393.8000 1233.3000 1395.0000 1240.5000 ;
	    RECT 1420.5000 1239.3000 1425.9000 1239.9000 ;
	    RECT 1427.4000 1239.3000 1428.3000 1240.5000 ;
	    RECT 1451.7001 1239.3000 1452.6000 1240.5000 ;
	    RECT 1477.8000 1240.2001 1479.0000 1240.5000 ;
	    RECT 1454.1000 1239.3000 1459.5000 1239.9000 ;
	    RECT 1480.2001 1239.3000 1481.4000 1243.5000 ;
	    RECT 1509.6000 1242.6000 1510.5000 1247.7001 ;
	    RECT 1511.4000 1245.4501 1512.6000 1245.6000 ;
	    RECT 1511.4000 1244.5500 1517.2500 1245.4501 ;
	    RECT 1511.4000 1244.4000 1512.6000 1244.5500 ;
	    RECT 1511.4000 1243.2001 1512.6000 1243.5000 ;
	    RECT 1494.6000 1242.4501 1495.8000 1242.6000 ;
	    RECT 1506.6000 1242.4501 1507.8000 1242.6000 ;
	    RECT 1494.6000 1241.5500 1507.8000 1242.4501 ;
	    RECT 1494.6000 1241.4000 1495.8000 1241.5500 ;
	    RECT 1506.6000 1241.4000 1507.8000 1241.5500 ;
	    RECT 1508.7001 1241.4000 1510.5000 1242.6000 ;
	    RECT 1512.6000 1240.8000 1512.9000 1242.3000 ;
	    RECT 1513.8000 1241.4000 1515.0000 1242.6000 ;
	    RECT 1516.3500 1242.4501 1517.2500 1244.5500 ;
	    RECT 1528.2001 1243.5000 1529.4000 1259.7001 ;
	    RECT 1530.6000 1253.7001 1531.8000 1259.7001 ;
	    RECT 1549.8000 1253.7001 1551.0000 1259.7001 ;
	    RECT 1549.8000 1249.5000 1551.0000 1249.8000 ;
	    RECT 1530.6000 1248.4501 1531.8000 1248.6000 ;
	    RECT 1549.8000 1248.4501 1551.0000 1248.6000 ;
	    RECT 1530.6000 1247.5500 1551.0000 1248.4501 ;
	    RECT 1530.6000 1247.4000 1531.8000 1247.5500 ;
	    RECT 1549.8000 1247.4000 1551.0000 1247.5500 ;
	    RECT 1552.2001 1246.5000 1553.4000 1259.7001 ;
	    RECT 1554.6000 1253.7001 1555.8000 1259.7001 ;
	    RECT 1530.6000 1245.4501 1531.8000 1245.6000 ;
	    RECT 1552.2001 1245.4501 1553.4000 1245.6000 ;
	    RECT 1530.6000 1244.5500 1553.4000 1245.4501 ;
	    RECT 1530.6000 1244.4000 1531.8000 1244.5500 ;
	    RECT 1552.2001 1244.4000 1553.4000 1244.5500 ;
	    RECT 1528.2001 1242.4501 1529.4000 1242.6000 ;
	    RECT 1516.3500 1241.5500 1529.4000 1242.4501 ;
	    RECT 1528.2001 1241.4000 1529.4000 1241.5500 ;
	    RECT 1506.9000 1239.3000 1507.8000 1240.5000 ;
	    RECT 1509.3000 1239.3000 1514.7001 1239.9000 ;
	    RECT 1420.2001 1239.0000 1426.2001 1239.3000 ;
	    RECT 1420.2001 1233.3000 1421.4000 1239.0000 ;
	    RECT 1422.6000 1233.3000 1423.8000 1238.1000 ;
	    RECT 1425.0000 1233.3000 1426.2001 1239.0000 ;
	    RECT 1427.4000 1233.3000 1428.6000 1239.3000 ;
	    RECT 1451.4000 1233.3000 1452.6000 1239.3000 ;
	    RECT 1453.8000 1239.0000 1459.8000 1239.3000 ;
	    RECT 1453.8000 1233.3000 1455.0000 1239.0000 ;
	    RECT 1456.2001 1233.3000 1457.4000 1238.1000 ;
	    RECT 1458.6000 1233.3000 1459.8000 1239.0000 ;
	    RECT 1477.8000 1233.3000 1479.0000 1239.3000 ;
	    RECT 1480.2001 1238.4000 1482.9000 1239.3000 ;
	    RECT 1481.7001 1233.3000 1482.9000 1238.4000 ;
	    RECT 1506.6000 1233.3000 1507.8000 1239.3000 ;
	    RECT 1509.0000 1239.0000 1515.0000 1239.3000 ;
	    RECT 1509.0000 1233.3000 1510.2001 1239.0000 ;
	    RECT 1511.4000 1233.3000 1512.6000 1238.1000 ;
	    RECT 1513.8000 1233.3000 1515.0000 1239.0000 ;
	    RECT 1528.2001 1233.3000 1529.4000 1240.5000 ;
	    RECT 1530.6000 1239.4501 1531.8000 1239.6000 ;
	    RECT 1547.4000 1239.4501 1548.6000 1239.6000 ;
	    RECT 1530.6000 1238.5500 1548.6000 1239.4501 ;
	    RECT 1552.2001 1239.3000 1553.4000 1243.5000 ;
	    RECT 1554.6000 1240.2001 1555.8000 1240.5000 ;
	    RECT 1530.6000 1238.4000 1531.8000 1238.5500 ;
	    RECT 1547.4000 1238.4000 1548.6000 1238.5500 ;
	    RECT 1550.7001 1238.4000 1553.4000 1239.3000 ;
	    RECT 1530.6000 1237.2001 1531.8000 1237.5000 ;
	    RECT 1530.6000 1233.3000 1531.8000 1236.3000 ;
	    RECT 1550.7001 1233.3000 1551.9000 1238.4000 ;
	    RECT 1554.6000 1233.3000 1555.8000 1239.3000 ;
	    RECT 1.2000 1230.6000 1569.0000 1232.4000 ;
	    RECT 124.2000 1220.7001 125.4000 1229.7001 ;
	    RECT 129.0000 1223.7001 130.2000 1229.7001 ;
	    RECT 133.8000 1224.9000 135.0000 1229.7001 ;
	    RECT 136.2000 1225.5000 137.4000 1229.7001 ;
	    RECT 138.6000 1225.5000 139.8000 1229.7001 ;
	    RECT 141.0000 1225.5000 142.2000 1229.7001 ;
	    RECT 143.4000 1226.7001 144.6000 1229.7001 ;
	    RECT 145.8000 1225.5000 147.0000 1229.7001 ;
	    RECT 148.2000 1226.7001 149.4000 1229.7001 ;
	    RECT 150.6000 1225.5000 151.8000 1229.7001 ;
	    RECT 153.0000 1225.5000 154.2000 1229.7001 ;
	    RECT 155.4000 1225.5000 156.6000 1229.7001 ;
	    RECT 157.8000 1225.5000 159.0000 1229.7001 ;
	    RECT 131.1000 1223.7001 135.0000 1224.9000 ;
	    RECT 160.2000 1224.9000 161.4000 1229.7001 ;
	    RECT 140.1000 1223.7001 147.0000 1224.6000 ;
	    RECT 131.1000 1222.8000 132.3000 1223.7001 ;
	    RECT 127.8000 1221.6000 132.3000 1222.8000 ;
	    RECT 124.2000 1219.5000 137.4000 1220.7001 ;
	    RECT 140.1000 1220.1000 141.3000 1223.7001 ;
	    RECT 145.8000 1223.4000 147.0000 1223.7001 ;
	    RECT 148.2000 1223.4000 149.4000 1224.6000 ;
	    RECT 150.3000 1223.4000 150.6000 1224.6000 ;
	    RECT 155.1000 1223.4000 156.6000 1224.6000 ;
	    RECT 160.2000 1223.7001 163.8000 1224.9000 ;
	    RECT 165.0000 1223.7001 166.2000 1229.7001 ;
	    RECT 143.4000 1222.5000 144.6000 1222.8000 ;
	    RECT 145.8000 1222.2001 147.0000 1222.5000 ;
	    RECT 143.4000 1220.4000 144.6000 1221.6000 ;
	    RECT 145.8000 1221.3000 152.4000 1222.2001 ;
	    RECT 151.2000 1221.0000 152.4000 1221.3000 ;
	    RECT 124.2000 1211.1000 125.4000 1219.5000 ;
	    RECT 138.3000 1218.9000 141.3000 1220.1000 ;
	    RECT 147.0000 1218.9000 151.8000 1220.1000 ;
	    RECT 155.4000 1219.2001 156.6000 1223.4000 ;
	    RECT 162.6000 1222.8000 163.8000 1223.7001 ;
	    RECT 162.6000 1221.9000 165.3000 1222.8000 ;
	    RECT 164.1000 1220.1000 165.3000 1221.9000 ;
	    RECT 169.8000 1221.9000 171.0000 1229.7001 ;
	    RECT 172.2000 1224.0000 173.4000 1229.7001 ;
	    RECT 174.6000 1226.7001 175.8000 1229.7001 ;
	    RECT 172.2000 1222.8000 173.7000 1224.0000 ;
	    RECT 169.8000 1221.0000 171.6000 1221.9000 ;
	    RECT 164.1000 1218.9000 169.8000 1220.1000 ;
	    RECT 126.3000 1218.0000 127.5000 1218.3000 ;
	    RECT 126.3000 1217.1000 132.9000 1218.0000 ;
	    RECT 133.8000 1217.4000 135.0000 1218.6000 ;
	    RECT 160.2000 1218.0000 161.4000 1218.9000 ;
	    RECT 170.7000 1218.0000 171.6000 1221.0000 ;
	    RECT 135.9000 1217.1000 161.4000 1218.0000 ;
	    RECT 170.4000 1217.1000 171.6000 1218.0000 ;
	    RECT 168.3000 1216.2001 169.5000 1216.5000 ;
	    RECT 129.0000 1214.4000 130.2000 1215.6000 ;
	    RECT 131.1000 1215.3000 169.5000 1216.2001 ;
	    RECT 134.1000 1215.0000 135.3000 1215.3000 ;
	    RECT 170.4000 1214.4000 171.3000 1217.1000 ;
	    RECT 172.5000 1216.2001 173.7000 1222.8000 ;
	    RECT 186.6000 1222.5000 187.8000 1229.7001 ;
	    RECT 189.0000 1226.7001 190.2000 1229.7001 ;
	    RECT 189.0000 1225.5000 190.2000 1225.8000 ;
	    RECT 189.0000 1223.4000 190.2000 1224.6000 ;
	    RECT 210.6000 1222.5000 211.8000 1229.7001 ;
	    RECT 213.0000 1226.7001 214.2000 1229.7001 ;
	    RECT 244.2000 1228.8000 250.2000 1229.7001 ;
	    RECT 213.0000 1225.5000 214.2000 1225.8000 ;
	    RECT 213.0000 1223.4000 214.2000 1224.6000 ;
	    RECT 244.2000 1223.7001 245.4000 1228.8000 ;
	    RECT 246.6000 1223.7001 247.8000 1227.9000 ;
	    RECT 249.0000 1224.0000 250.2000 1228.8000 ;
	    RECT 251.4000 1224.9000 252.6000 1229.7001 ;
	    RECT 253.8000 1224.0000 255.0000 1229.7001 ;
	    RECT 268.2000 1226.7001 269.4000 1229.7001 ;
	    RECT 268.2000 1225.5000 269.4000 1225.8000 ;
	    RECT 249.0000 1223.7001 255.0000 1224.0000 ;
	    RECT 263.4000 1224.4501 264.6000 1224.6000 ;
	    RECT 268.2000 1224.4501 269.4000 1224.6000 ;
	    RECT 246.6000 1221.6000 247.5000 1223.7001 ;
	    RECT 249.3000 1223.1000 254.7000 1223.7001 ;
	    RECT 263.4000 1223.5500 269.4000 1224.4501 ;
	    RECT 263.4000 1223.4000 264.6000 1223.5500 ;
	    RECT 268.2000 1223.4000 269.4000 1223.5500 ;
	    RECT 270.6000 1222.5000 271.8000 1229.7001 ;
	    RECT 282.6000 1222.5000 283.8000 1229.7001 ;
	    RECT 285.0000 1226.7001 286.2000 1229.7001 ;
	    RECT 285.0000 1225.5000 286.2000 1225.8000 ;
	    RECT 305.1000 1224.6000 306.3000 1229.7001 ;
	    RECT 285.0000 1223.4000 286.2000 1224.6000 ;
	    RECT 305.1000 1223.7001 307.8000 1224.6000 ;
	    RECT 309.0000 1223.7001 310.2000 1229.7001 ;
	    RECT 186.6000 1221.4501 187.8000 1221.6000 ;
	    RECT 198.6000 1221.4501 199.8000 1221.6000 ;
	    RECT 186.6000 1220.5500 199.8000 1221.4501 ;
	    RECT 186.6000 1220.4000 187.8000 1220.5500 ;
	    RECT 198.6000 1220.4000 199.8000 1220.5500 ;
	    RECT 210.6000 1221.4501 211.8000 1221.6000 ;
	    RECT 244.2000 1221.4501 245.4000 1221.6000 ;
	    RECT 210.6000 1220.5500 245.4000 1221.4501 ;
	    RECT 246.6000 1220.7001 248.1000 1221.6000 ;
	    RECT 210.6000 1220.4000 211.8000 1220.5500 ;
	    RECT 244.2000 1220.4000 245.4000 1220.5500 ;
	    RECT 249.0000 1220.4000 250.2000 1221.6000 ;
	    RECT 252.6000 1220.7001 252.9000 1222.2001 ;
	    RECT 253.8000 1220.4000 255.0000 1221.6000 ;
	    RECT 256.2000 1221.4501 257.4000 1221.6000 ;
	    RECT 270.6000 1221.4501 271.8000 1221.6000 ;
	    RECT 256.2000 1220.5500 271.8000 1221.4501 ;
	    RECT 256.2000 1220.4000 257.4000 1220.5500 ;
	    RECT 270.6000 1220.4000 271.8000 1220.5500 ;
	    RECT 273.0000 1221.4501 274.2000 1221.6000 ;
	    RECT 282.6000 1221.4501 283.8000 1221.6000 ;
	    RECT 273.0000 1220.5500 283.8000 1221.4501 ;
	    RECT 273.0000 1220.4000 274.2000 1220.5500 ;
	    RECT 282.6000 1220.4000 283.8000 1220.5500 ;
	    RECT 246.6000 1219.5000 247.8000 1219.8000 ;
	    RECT 251.4000 1219.5000 252.6000 1219.8000 ;
	    RECT 306.6000 1219.5000 307.8000 1223.7001 ;
	    RECT 309.0000 1222.5000 310.2000 1222.8000 ;
	    RECT 323.4000 1222.5000 324.6000 1229.7001 ;
	    RECT 325.8000 1226.7001 327.0000 1229.7001 ;
	    RECT 325.8000 1225.5000 327.0000 1225.8000 ;
	    RECT 325.8000 1223.4000 327.0000 1224.6000 ;
	    RECT 345.0000 1223.7001 346.2000 1229.7001 ;
	    RECT 348.9000 1224.6000 350.1000 1229.7001 ;
	    RECT 347.4000 1223.7001 350.1000 1224.6000 ;
	    RECT 345.0000 1222.5000 346.2000 1222.8000 ;
	    RECT 309.0000 1220.4000 310.2000 1221.6000 ;
	    RECT 323.4000 1221.4501 324.6000 1221.6000 ;
	    RECT 330.6000 1221.4501 331.8000 1221.6000 ;
	    RECT 323.4000 1220.5500 331.8000 1221.4501 ;
	    RECT 323.4000 1220.4000 324.6000 1220.5500 ;
	    RECT 330.6000 1220.4000 331.8000 1220.5500 ;
	    RECT 345.0000 1220.4000 346.2000 1221.6000 ;
	    RECT 347.4000 1219.5000 348.6000 1223.7001 ;
	    RECT 364.2000 1222.5000 365.4000 1229.7001 ;
	    RECT 366.6000 1226.7001 367.8000 1229.7001 ;
	    RECT 366.6000 1225.5000 367.8000 1225.8000 ;
	    RECT 366.6000 1224.4501 367.8000 1224.6000 ;
	    RECT 369.0000 1224.4501 370.2000 1224.6000 ;
	    RECT 381.0000 1224.4501 382.2000 1224.6000 ;
	    RECT 366.6000 1223.5500 382.2000 1224.4501 ;
	    RECT 366.6000 1223.4000 367.8000 1223.5500 ;
	    RECT 369.0000 1223.4000 370.2000 1223.5500 ;
	    RECT 381.0000 1223.4000 382.2000 1223.5500 ;
	    RECT 385.8000 1222.8000 387.0000 1229.7001 ;
	    RECT 388.2000 1223.7001 389.4000 1229.7001 ;
	    RECT 385.8000 1221.9000 389.1000 1222.8000 ;
	    RECT 390.6000 1222.5000 391.8000 1229.7001 ;
	    RECT 522.6000 1226.7001 523.8000 1229.7001 ;
	    RECT 525.0000 1224.0000 526.2000 1229.7001 ;
	    RECT 524.7000 1222.8000 526.2000 1224.0000 ;
	    RECT 364.2000 1221.4501 365.4000 1221.6000 ;
	    RECT 378.6000 1221.4501 379.8000 1221.6000 ;
	    RECT 364.2000 1220.5500 379.8000 1221.4501 ;
	    RECT 364.2000 1220.4000 365.4000 1220.5500 ;
	    RECT 378.6000 1220.4000 379.8000 1220.5500 ;
	    RECT 385.8000 1219.5000 387.0000 1219.8000 ;
	    RECT 138.6000 1214.1000 139.8000 1214.4000 ;
	    RECT 131.7000 1213.5000 139.8000 1214.1000 ;
	    RECT 130.5000 1213.2001 139.8000 1213.5000 ;
	    RECT 141.3000 1213.5000 154.2000 1214.4000 ;
	    RECT 126.6000 1212.0000 129.0000 1213.2001 ;
	    RECT 130.5000 1212.3000 132.6000 1213.2001 ;
	    RECT 141.3000 1212.3000 142.2000 1213.5000 ;
	    RECT 153.0000 1213.2001 154.2000 1213.5000 ;
	    RECT 157.8000 1213.5000 171.3000 1214.4000 ;
	    RECT 172.2000 1215.0000 173.7000 1216.2001 ;
	    RECT 172.2000 1213.5000 173.4000 1215.0000 ;
	    RECT 157.8000 1213.2001 159.0000 1213.5000 ;
	    RECT 128.1000 1211.4000 129.0000 1212.0000 ;
	    RECT 133.5000 1211.4000 142.2000 1212.3000 ;
	    RECT 143.1000 1211.4000 147.0000 1212.6000 ;
	    RECT 124.2000 1210.2001 127.2000 1211.1000 ;
	    RECT 128.1000 1210.2001 134.4000 1211.4000 ;
	    RECT 126.3000 1209.3000 127.2000 1210.2001 ;
	    RECT 124.2000 1203.3000 125.4000 1209.3000 ;
	    RECT 126.3000 1208.4000 127.8000 1209.3000 ;
	    RECT 126.6000 1203.3000 127.8000 1208.4000 ;
	    RECT 129.0000 1202.4000 130.2000 1209.3000 ;
	    RECT 131.4000 1203.3000 132.6000 1210.2001 ;
	    RECT 133.8000 1203.3000 135.0000 1209.3000 ;
	    RECT 136.2000 1203.3000 137.4000 1207.5000 ;
	    RECT 138.6000 1203.3000 139.8000 1207.5000 ;
	    RECT 141.0000 1203.3000 142.2000 1210.5000 ;
	    RECT 143.4000 1203.3000 144.6000 1209.3000 ;
	    RECT 145.8000 1203.3000 147.0000 1210.5000 ;
	    RECT 148.2000 1203.3000 149.4000 1209.3000 ;
	    RECT 150.6000 1203.3000 151.8000 1212.6000 ;
	    RECT 162.6000 1211.4000 166.5000 1212.6000 ;
	    RECT 155.4000 1210.2001 161.7000 1211.4000 ;
	    RECT 153.0000 1203.3000 154.2000 1207.5000 ;
	    RECT 155.4000 1203.3000 156.6000 1207.5000 ;
	    RECT 157.8000 1203.3000 159.0000 1207.5000 ;
	    RECT 160.2000 1203.3000 161.4000 1209.3000 ;
	    RECT 162.6000 1203.3000 163.8000 1211.4000 ;
	    RECT 170.4000 1211.1000 171.3000 1213.5000 ;
	    RECT 172.2000 1211.4000 173.4000 1212.6000 ;
	    RECT 167.4000 1210.2001 171.3000 1211.1000 ;
	    RECT 165.0000 1203.3000 166.2000 1209.3000 ;
	    RECT 167.4000 1203.3000 168.6000 1210.2001 ;
	    RECT 169.8000 1203.3000 171.0000 1209.3000 ;
	    RECT 172.2000 1203.3000 173.4000 1210.5000 ;
	    RECT 174.6000 1203.3000 175.8000 1209.3000 ;
	    RECT 186.6000 1203.3000 187.8000 1219.5000 ;
	    RECT 189.0000 1203.3000 190.2000 1209.3000 ;
	    RECT 210.6000 1203.3000 211.8000 1219.5000 ;
	    RECT 244.2000 1219.2001 245.4000 1219.5000 ;
	    RECT 246.6000 1217.4000 247.8000 1218.6000 ;
	    RECT 249.3000 1215.3000 250.2000 1219.5000 ;
	    RECT 251.4000 1217.4000 252.6000 1218.6000 ;
	    RECT 213.0000 1203.3000 214.2000 1209.3000 ;
	    RECT 244.2000 1203.3000 245.4000 1215.3000 ;
	    RECT 248.1000 1203.3000 251.1000 1215.3000 ;
	    RECT 253.8000 1203.3000 255.0000 1215.3000 ;
	    RECT 268.2000 1203.3000 269.4000 1209.3000 ;
	    RECT 270.6000 1203.3000 271.8000 1219.5000 ;
	    RECT 282.6000 1203.3000 283.8000 1219.5000 ;
	    RECT 287.4000 1218.4501 288.6000 1218.6000 ;
	    RECT 306.6000 1218.4501 307.8000 1218.6000 ;
	    RECT 287.4000 1217.5500 307.8000 1218.4501 ;
	    RECT 287.4000 1217.4000 288.6000 1217.5500 ;
	    RECT 306.6000 1217.4000 307.8000 1217.5500 ;
	    RECT 304.2000 1214.4000 305.4000 1215.6000 ;
	    RECT 304.2000 1213.2001 305.4000 1213.5000 ;
	    RECT 285.0000 1203.3000 286.2000 1209.3000 ;
	    RECT 304.2000 1203.3000 305.4000 1209.3000 ;
	    RECT 306.6000 1203.3000 307.8000 1216.5000 ;
	    RECT 309.0000 1203.3000 310.2000 1209.3000 ;
	    RECT 323.4000 1203.3000 324.6000 1219.5000 ;
	    RECT 337.8000 1218.4501 339.0000 1218.6000 ;
	    RECT 347.4000 1218.4501 348.6000 1218.6000 ;
	    RECT 337.8000 1217.5500 348.6000 1218.4501 ;
	    RECT 337.8000 1217.4000 339.0000 1217.5500 ;
	    RECT 347.4000 1217.4000 348.6000 1217.5500 ;
	    RECT 325.8000 1203.3000 327.0000 1209.3000 ;
	    RECT 345.0000 1203.3000 346.2000 1209.3000 ;
	    RECT 347.4000 1203.3000 348.6000 1216.5000 ;
	    RECT 349.8000 1215.4501 351.0000 1215.6000 ;
	    RECT 357.0000 1215.4501 358.2000 1215.6000 ;
	    RECT 349.8000 1214.5500 358.2000 1215.4501 ;
	    RECT 349.8000 1214.4000 351.0000 1214.5500 ;
	    RECT 357.0000 1214.4000 358.2000 1214.5500 ;
	    RECT 349.8000 1213.2001 351.0000 1213.5000 ;
	    RECT 349.8000 1203.3000 351.0000 1209.3000 ;
	    RECT 364.2000 1203.3000 365.4000 1219.5000 ;
	    RECT 385.8000 1217.4000 387.0000 1218.6000 ;
	    RECT 388.2000 1217.4000 389.1000 1221.9000 ;
	    RECT 390.6000 1220.4000 391.8000 1221.6000 ;
	    RECT 390.6000 1218.6000 391.8000 1219.5000 ;
	    RECT 388.2000 1216.2001 390.0000 1217.4000 ;
	    RECT 388.2000 1215.3000 389.1000 1216.2001 ;
	    RECT 390.9000 1215.3000 391.8000 1218.6000 ;
	    RECT 385.8000 1214.4000 389.1000 1215.3000 ;
	    RECT 366.6000 1203.3000 367.8000 1209.3000 ;
	    RECT 385.8000 1203.3000 387.0000 1214.4000 ;
	    RECT 388.2000 1203.3000 389.4000 1213.5000 ;
	    RECT 390.6000 1203.3000 391.8000 1215.3000 ;
	    RECT 524.7000 1216.2001 525.9000 1222.8000 ;
	    RECT 527.4000 1221.9000 528.6000 1229.7001 ;
	    RECT 532.2000 1223.7001 533.4000 1229.7001 ;
	    RECT 537.0000 1224.9000 538.2000 1229.7001 ;
	    RECT 539.4000 1225.5000 540.6000 1229.7001 ;
	    RECT 541.8000 1225.5000 543.0000 1229.7001 ;
	    RECT 544.2000 1225.5000 545.4000 1229.7001 ;
	    RECT 546.6000 1225.5000 547.8000 1229.7001 ;
	    RECT 549.0000 1226.7001 550.2000 1229.7001 ;
	    RECT 551.4000 1225.5000 552.6000 1229.7001 ;
	    RECT 553.8000 1226.7001 555.0000 1229.7001 ;
	    RECT 556.2000 1225.5000 557.4000 1229.7001 ;
	    RECT 558.6000 1225.5000 559.8000 1229.7001 ;
	    RECT 561.0000 1225.5000 562.2000 1229.7001 ;
	    RECT 534.6000 1223.7001 538.2000 1224.9000 ;
	    RECT 563.4000 1224.9000 564.6000 1229.7001 ;
	    RECT 534.6000 1222.8000 535.8000 1223.7001 ;
	    RECT 526.8000 1221.0000 528.6000 1221.9000 ;
	    RECT 533.1000 1221.9000 535.8000 1222.8000 ;
	    RECT 541.8000 1223.4000 543.3000 1224.6000 ;
	    RECT 547.8000 1223.4000 548.1000 1224.6000 ;
	    RECT 549.0000 1223.4000 550.2000 1224.6000 ;
	    RECT 551.4000 1223.7001 558.3000 1224.6000 ;
	    RECT 563.4000 1223.7001 567.3000 1224.9000 ;
	    RECT 568.2000 1223.7001 569.4000 1229.7001 ;
	    RECT 551.4000 1223.4000 552.6000 1223.7001 ;
	    RECT 526.8000 1218.0000 527.7000 1221.0000 ;
	    RECT 533.1000 1220.1000 534.3000 1221.9000 ;
	    RECT 528.6000 1218.9000 534.3000 1220.1000 ;
	    RECT 541.8000 1219.2001 543.0000 1223.4000 ;
	    RECT 553.8000 1222.5000 555.0000 1222.8000 ;
	    RECT 551.4000 1222.2001 552.6000 1222.5000 ;
	    RECT 546.0000 1221.3000 552.6000 1222.2001 ;
	    RECT 546.0000 1221.0000 547.2000 1221.3000 ;
	    RECT 553.8000 1220.4000 555.0000 1221.6000 ;
	    RECT 557.1000 1220.1000 558.3000 1223.7001 ;
	    RECT 566.1000 1222.8000 567.3000 1223.7001 ;
	    RECT 566.1000 1221.6000 570.6000 1222.8000 ;
	    RECT 573.0000 1220.7001 574.2000 1229.7001 ;
	    RECT 597.0000 1223.7001 598.2000 1229.7001 ;
	    RECT 599.4000 1224.0000 600.6000 1229.7001 ;
	    RECT 601.8000 1224.9000 603.0000 1229.7001 ;
	    RECT 604.2000 1224.0000 605.4000 1229.7001 ;
	    RECT 599.4000 1223.7001 605.4000 1224.0000 ;
	    RECT 630.6000 1223.7001 631.8000 1229.7001 ;
	    RECT 634.5000 1224.0000 635.7000 1229.7001 ;
	    RECT 636.9000 1225.2001 638.1000 1229.7001 ;
	    RECT 649.8000 1226.7001 651.0000 1229.7001 ;
	    RECT 649.8000 1225.5000 651.0000 1225.8000 ;
	    RECT 636.9000 1223.7001 639.0000 1225.2001 ;
	    RECT 597.3000 1222.5000 598.2000 1223.7001 ;
	    RECT 599.7000 1223.1000 605.1000 1223.7001 ;
	    RECT 630.9000 1223.4000 631.8000 1223.7001 ;
	    RECT 630.9000 1222.8000 633.6000 1223.4000 ;
	    RECT 630.9000 1222.5000 637.2000 1222.8000 ;
	    RECT 546.6000 1218.9000 551.4000 1220.1000 ;
	    RECT 557.1000 1218.9000 560.1000 1220.1000 ;
	    RECT 561.0000 1219.5000 574.2000 1220.7001 ;
	    RECT 597.0000 1220.4000 598.2000 1221.6000 ;
	    RECT 599.1000 1220.4000 600.9000 1221.6000 ;
	    RECT 603.0000 1220.7001 603.3000 1222.2001 ;
	    RECT 632.7000 1221.9000 637.2000 1222.5000 ;
	    RECT 636.0000 1221.6000 637.2000 1221.9000 ;
	    RECT 604.2000 1220.4000 605.4000 1221.6000 ;
	    RECT 625.8000 1221.4501 627.0000 1221.6000 ;
	    RECT 630.6000 1221.4501 631.8000 1221.6000 ;
	    RECT 625.8000 1220.5500 631.8000 1221.4501 ;
	    RECT 633.6000 1220.7001 634.8000 1221.0000 ;
	    RECT 625.8000 1220.4000 627.0000 1220.5500 ;
	    RECT 630.6000 1220.4000 631.8000 1220.5500 ;
	    RECT 537.0000 1218.0000 538.2000 1218.9000 ;
	    RECT 526.8000 1217.1000 528.0000 1218.0000 ;
	    RECT 537.0000 1217.1000 562.5000 1218.0000 ;
	    RECT 563.4000 1217.4000 564.6000 1218.6000 ;
	    RECT 570.9000 1218.0000 572.1000 1218.3000 ;
	    RECT 565.5000 1217.1000 572.1000 1218.0000 ;
	    RECT 524.7000 1215.0000 526.2000 1216.2001 ;
	    RECT 525.0000 1213.5000 526.2000 1215.0000 ;
	    RECT 527.1000 1214.4000 528.0000 1217.1000 ;
	    RECT 528.9000 1216.2001 530.1000 1216.5000 ;
	    RECT 528.9000 1215.3000 567.3000 1216.2001 ;
	    RECT 563.1000 1215.0000 564.3000 1215.3000 ;
	    RECT 568.2000 1214.4000 569.4000 1215.6000 ;
	    RECT 527.1000 1213.5000 540.6000 1214.4000 ;
	    RECT 419.4000 1212.4501 420.6000 1212.6000 ;
	    RECT 525.0000 1212.4501 526.2000 1212.6000 ;
	    RECT 419.4000 1211.5500 526.2000 1212.4501 ;
	    RECT 419.4000 1211.4000 420.6000 1211.5500 ;
	    RECT 525.0000 1211.4000 526.2000 1211.5500 ;
	    RECT 527.1000 1211.1000 528.0000 1213.5000 ;
	    RECT 539.4000 1213.2001 540.6000 1213.5000 ;
	    RECT 544.2000 1213.5000 557.1000 1214.4000 ;
	    RECT 544.2000 1213.2001 545.4000 1213.5000 ;
	    RECT 531.9000 1211.4000 535.8000 1212.6000 ;
	    RECT 522.6000 1203.3000 523.8000 1209.3000 ;
	    RECT 525.0000 1203.3000 526.2000 1210.5000 ;
	    RECT 527.1000 1210.2001 531.0000 1211.1000 ;
	    RECT 527.4000 1203.3000 528.6000 1209.3000 ;
	    RECT 529.8000 1203.3000 531.0000 1210.2001 ;
	    RECT 532.2000 1203.3000 533.4000 1209.3000 ;
	    RECT 534.6000 1203.3000 535.8000 1211.4000 ;
	    RECT 536.7000 1210.2001 543.0000 1211.4000 ;
	    RECT 537.0000 1203.3000 538.2000 1209.3000 ;
	    RECT 539.4000 1203.3000 540.6000 1207.5000 ;
	    RECT 541.8000 1203.3000 543.0000 1207.5000 ;
	    RECT 544.2000 1203.3000 545.4000 1207.5000 ;
	    RECT 546.6000 1203.3000 547.8000 1212.6000 ;
	    RECT 551.4000 1211.4000 555.3000 1212.6000 ;
	    RECT 556.2000 1212.3000 557.1000 1213.5000 ;
	    RECT 558.6000 1214.1000 559.8000 1214.4000 ;
	    RECT 558.6000 1213.5000 566.7000 1214.1000 ;
	    RECT 558.6000 1213.2001 567.9000 1213.5000 ;
	    RECT 565.8000 1212.3000 567.9000 1213.2001 ;
	    RECT 556.2000 1211.4000 564.9000 1212.3000 ;
	    RECT 569.4000 1212.0000 571.8000 1213.2001 ;
	    RECT 569.4000 1211.4000 570.3000 1212.0000 ;
	    RECT 549.0000 1203.3000 550.2000 1209.3000 ;
	    RECT 551.4000 1203.3000 552.6000 1210.5000 ;
	    RECT 553.8000 1203.3000 555.0000 1209.3000 ;
	    RECT 556.2000 1203.3000 557.4000 1210.5000 ;
	    RECT 564.0000 1210.2001 570.3000 1211.4000 ;
	    RECT 573.0000 1211.1000 574.2000 1219.5000 ;
	    RECT 597.0000 1214.4000 598.2000 1215.6000 ;
	    RECT 600.0000 1215.3000 600.9000 1220.4000 ;
	    RECT 633.3000 1219.8000 634.8000 1220.7001 ;
	    RECT 601.8000 1219.5000 603.0000 1219.8000 ;
	    RECT 633.3000 1219.5000 634.2000 1219.8000 ;
	    RECT 630.6000 1219.2001 631.8000 1219.5000 ;
	    RECT 601.8000 1217.4000 603.0000 1218.6000 ;
	    RECT 633.0000 1217.4000 634.2000 1218.6000 ;
	    RECT 636.0000 1216.5000 636.9000 1221.6000 ;
	    RECT 638.1000 1219.5000 639.0000 1223.7001 ;
	    RECT 649.8000 1223.4000 651.0000 1224.6000 ;
	    RECT 652.2000 1222.5000 653.4000 1229.7001 ;
	    RECT 678.6000 1223.7001 679.8000 1229.7001 ;
	    RECT 682.5000 1224.6000 683.7000 1229.7001 ;
	    RECT 681.0000 1223.7001 683.7000 1224.6000 ;
	    RECT 678.6000 1222.5000 679.8000 1222.8000 ;
	    RECT 652.2000 1221.4501 653.4000 1221.6000 ;
	    RECT 657.0000 1221.4501 658.2000 1221.6000 ;
	    RECT 652.2000 1220.5500 658.2000 1221.4501 ;
	    RECT 652.2000 1220.4000 653.4000 1220.5500 ;
	    RECT 657.0000 1220.4000 658.2000 1220.5500 ;
	    RECT 661.8000 1221.4501 663.0000 1221.6000 ;
	    RECT 678.6000 1221.4501 679.8000 1221.6000 ;
	    RECT 661.8000 1220.5500 679.8000 1221.4501 ;
	    RECT 661.8000 1220.4000 663.0000 1220.5500 ;
	    RECT 678.6000 1220.4000 679.8000 1220.5500 ;
	    RECT 681.0000 1219.5000 682.2000 1223.7001 ;
	    RECT 697.8000 1222.5000 699.0000 1229.7001 ;
	    RECT 700.2000 1226.7001 701.4000 1229.7001 ;
	    RECT 803.4000 1227.4501 804.6000 1227.6000 ;
	    RECT 810.6000 1227.4501 811.8000 1227.6000 ;
	    RECT 803.4000 1226.5500 811.8000 1227.4501 ;
	    RECT 803.4000 1226.4000 804.6000 1226.5500 ;
	    RECT 810.6000 1226.4000 811.8000 1226.5500 ;
	    RECT 700.2000 1225.5000 701.4000 1225.8000 ;
	    RECT 700.2000 1224.4501 701.4000 1224.6000 ;
	    RECT 757.8000 1224.4501 759.0000 1224.6000 ;
	    RECT 825.0000 1224.4501 826.2000 1224.6000 ;
	    RECT 700.2000 1223.5500 826.2000 1224.4501 ;
	    RECT 700.2000 1223.4000 701.4000 1223.5500 ;
	    RECT 757.8000 1223.4000 759.0000 1223.5500 ;
	    RECT 825.0000 1223.4000 826.2000 1223.5500 ;
	    RECT 697.8000 1220.4000 699.0000 1221.6000 ;
	    RECT 827.4000 1220.7001 828.6000 1229.7001 ;
	    RECT 832.2000 1223.7001 833.4000 1229.7001 ;
	    RECT 837.0000 1224.9000 838.2000 1229.7001 ;
	    RECT 839.4000 1225.5000 840.6000 1229.7001 ;
	    RECT 841.8000 1225.5000 843.0000 1229.7001 ;
	    RECT 844.2000 1225.5000 845.4000 1229.7001 ;
	    RECT 846.6000 1226.7001 847.8000 1229.7001 ;
	    RECT 849.0000 1225.5000 850.2000 1229.7001 ;
	    RECT 851.4000 1226.7001 852.6000 1229.7001 ;
	    RECT 853.8000 1225.5000 855.0000 1229.7001 ;
	    RECT 856.2000 1225.5000 857.4000 1229.7001 ;
	    RECT 858.6000 1225.5000 859.8000 1229.7001 ;
	    RECT 861.0000 1225.5000 862.2000 1229.7001 ;
	    RECT 834.3000 1223.7001 838.2000 1224.9000 ;
	    RECT 863.4000 1224.9000 864.6000 1229.7001 ;
	    RECT 843.3000 1223.7001 850.2000 1224.6000 ;
	    RECT 834.3000 1222.8000 835.5000 1223.7001 ;
	    RECT 831.0000 1221.6000 835.5000 1222.8000 ;
	    RECT 827.4000 1219.5000 840.6000 1220.7001 ;
	    RECT 843.3000 1220.1000 844.5000 1223.7001 ;
	    RECT 849.0000 1223.4000 850.2000 1223.7001 ;
	    RECT 851.4000 1223.4000 852.6000 1224.6000 ;
	    RECT 853.5000 1223.4000 853.8000 1224.6000 ;
	    RECT 858.3000 1223.4000 859.8000 1224.6000 ;
	    RECT 863.4000 1223.7001 867.0000 1224.9000 ;
	    RECT 868.2000 1223.7001 869.4000 1229.7001 ;
	    RECT 846.6000 1222.5000 847.8000 1222.8000 ;
	    RECT 849.0000 1222.2001 850.2000 1222.5000 ;
	    RECT 846.6000 1220.4000 847.8000 1221.6000 ;
	    RECT 849.0000 1221.3000 855.6000 1222.2001 ;
	    RECT 854.4000 1221.0000 855.6000 1221.3000 ;
	    RECT 637.8000 1218.4501 639.0000 1218.6000 ;
	    RECT 640.2000 1218.4501 641.4000 1218.6000 ;
	    RECT 637.8000 1217.5500 641.4000 1218.4501 ;
	    RECT 637.8000 1217.4000 639.0000 1217.5500 ;
	    RECT 640.2000 1217.4000 641.4000 1217.5500 ;
	    RECT 633.3000 1215.6000 636.9000 1216.5000 ;
	    RECT 600.0000 1214.4000 601.5000 1215.3000 ;
	    RECT 598.2000 1212.6000 599.1000 1213.5000 ;
	    RECT 598.2000 1211.4000 599.4000 1212.6000 ;
	    RECT 571.2000 1210.2001 574.2000 1211.1000 ;
	    RECT 558.6000 1203.3000 559.8000 1207.5000 ;
	    RECT 561.0000 1203.3000 562.2000 1207.5000 ;
	    RECT 563.4000 1203.3000 564.6000 1209.3000 ;
	    RECT 565.8000 1203.3000 567.0000 1210.2001 ;
	    RECT 571.2000 1209.3000 572.1000 1210.2001 ;
	    RECT 568.2000 1202.4000 569.4000 1209.3000 ;
	    RECT 570.6000 1208.4000 572.1000 1209.3000 ;
	    RECT 570.6000 1203.3000 571.8000 1208.4000 ;
	    RECT 573.0000 1203.3000 574.2000 1209.3000 ;
	    RECT 597.9000 1203.3000 599.1000 1209.3000 ;
	    RECT 600.3000 1203.3000 601.5000 1214.4000 ;
	    RECT 604.2000 1203.3000 605.4000 1215.3000 ;
	    RECT 633.3000 1209.3000 634.2000 1215.6000 ;
	    RECT 638.1000 1215.3000 639.0000 1216.5000 ;
	    RECT 630.6000 1203.3000 631.8000 1209.3000 ;
	    RECT 633.0000 1203.3000 634.2000 1209.3000 ;
	    RECT 635.4000 1203.3000 636.6000 1214.7001 ;
	    RECT 637.8000 1203.3000 639.0000 1215.3000 ;
	    RECT 649.8000 1203.3000 651.0000 1209.3000 ;
	    RECT 652.2000 1203.3000 653.4000 1219.5000 ;
	    RECT 681.0000 1218.4501 682.2000 1218.6000 ;
	    RECT 690.6000 1218.4501 691.8000 1218.6000 ;
	    RECT 681.0000 1217.5500 691.8000 1218.4501 ;
	    RECT 681.0000 1217.4000 682.2000 1217.5500 ;
	    RECT 690.6000 1217.4000 691.8000 1217.5500 ;
	    RECT 678.6000 1203.3000 679.8000 1209.3000 ;
	    RECT 681.0000 1203.3000 682.2000 1216.5000 ;
	    RECT 683.4000 1215.4501 684.6000 1215.6000 ;
	    RECT 693.0000 1215.4501 694.2000 1215.6000 ;
	    RECT 683.4000 1214.5500 694.2000 1215.4501 ;
	    RECT 683.4000 1214.4000 684.6000 1214.5500 ;
	    RECT 693.0000 1214.4000 694.2000 1214.5500 ;
	    RECT 683.4000 1213.2001 684.6000 1213.5000 ;
	    RECT 683.4000 1203.3000 684.6000 1209.3000 ;
	    RECT 697.8000 1203.3000 699.0000 1219.5000 ;
	    RECT 827.4000 1211.1000 828.6000 1219.5000 ;
	    RECT 841.5000 1218.9000 844.5000 1220.1000 ;
	    RECT 850.2000 1218.9000 855.0000 1220.1000 ;
	    RECT 858.6000 1219.2001 859.8000 1223.4000 ;
	    RECT 865.8000 1222.8000 867.0000 1223.7001 ;
	    RECT 865.8000 1221.9000 868.5000 1222.8000 ;
	    RECT 867.3000 1220.1000 868.5000 1221.9000 ;
	    RECT 873.0000 1221.9000 874.2000 1229.7001 ;
	    RECT 875.4000 1224.0000 876.6000 1229.7001 ;
	    RECT 877.8000 1226.7001 879.0000 1229.7001 ;
	    RECT 875.4000 1222.8000 876.9000 1224.0000 ;
	    RECT 904.2000 1223.7001 905.4000 1229.7001 ;
	    RECT 908.1000 1224.6000 909.3000 1229.7001 ;
	    RECT 928.2000 1226.7001 929.4000 1229.7001 ;
	    RECT 930.6000 1226.7001 931.8000 1229.7001 ;
	    RECT 933.0000 1226.7001 934.2000 1229.7001 ;
	    RECT 945.0000 1226.7001 946.2000 1229.7001 ;
	    RECT 906.6000 1223.7001 909.3000 1224.6000 ;
	    RECT 873.0000 1221.0000 874.8000 1221.9000 ;
	    RECT 867.3000 1218.9000 873.0000 1220.1000 ;
	    RECT 829.5000 1218.0000 830.7000 1218.3000 ;
	    RECT 829.5000 1217.1000 836.1000 1218.0000 ;
	    RECT 837.0000 1217.4000 838.2000 1218.6000 ;
	    RECT 863.4000 1218.0000 864.6000 1218.9000 ;
	    RECT 873.9000 1218.0000 874.8000 1221.0000 ;
	    RECT 839.1000 1217.1000 864.6000 1218.0000 ;
	    RECT 873.6000 1217.1000 874.8000 1218.0000 ;
	    RECT 871.5000 1216.2001 872.7000 1216.5000 ;
	    RECT 832.2000 1214.4000 833.4000 1215.6000 ;
	    RECT 834.3000 1215.3000 872.7000 1216.2001 ;
	    RECT 837.3000 1215.0000 838.5000 1215.3000 ;
	    RECT 873.6000 1214.4000 874.5000 1217.1000 ;
	    RECT 875.7000 1216.2001 876.9000 1222.8000 ;
	    RECT 904.2000 1222.5000 905.4000 1222.8000 ;
	    RECT 904.2000 1220.4000 905.4000 1221.6000 ;
	    RECT 906.6000 1219.5000 907.8000 1223.7001 ;
	    RECT 930.6000 1222.5000 931.5000 1226.7001 ;
	    RECT 933.0000 1225.5000 934.2000 1225.8000 ;
	    RECT 945.0000 1225.5000 946.2000 1225.8000 ;
	    RECT 933.0000 1223.4000 934.2000 1224.6000 ;
	    RECT 935.4000 1224.4501 936.6000 1224.6000 ;
	    RECT 945.0000 1224.4501 946.2000 1224.6000 ;
	    RECT 935.4000 1223.5500 946.2000 1224.4501 ;
	    RECT 935.4000 1223.4000 936.6000 1223.5500 ;
	    RECT 945.0000 1223.4000 946.2000 1223.5500 ;
	    RECT 947.4000 1222.5000 948.6000 1229.7001 ;
	    RECT 973.8000 1223.7001 975.0000 1229.7001 ;
	    RECT 976.2000 1224.0000 977.4000 1229.7001 ;
	    RECT 978.6000 1224.9000 979.8000 1229.7001 ;
	    RECT 981.0000 1224.0000 982.2000 1229.7001 ;
	    RECT 976.2000 1223.7001 982.2000 1224.0000 ;
	    RECT 1012.2000 1228.8000 1018.2000 1229.7001 ;
	    RECT 1012.2000 1223.7001 1013.4000 1228.8000 ;
	    RECT 1014.6000 1223.7001 1015.8000 1227.9000 ;
	    RECT 1017.0000 1224.0000 1018.2000 1228.8000 ;
	    RECT 1019.4000 1224.9000 1020.6000 1229.7001 ;
	    RECT 1021.8000 1224.0000 1023.0000 1229.7001 ;
	    RECT 1017.0000 1223.7001 1023.0000 1224.0000 ;
	    RECT 974.1000 1222.5000 975.0000 1223.7001 ;
	    RECT 976.5000 1223.1000 981.9000 1223.7001 ;
	    RECT 928.2000 1221.4501 929.4000 1221.6000 ;
	    RECT 930.6000 1221.4501 931.8000 1221.6000 ;
	    RECT 928.2000 1220.5500 931.8000 1221.4501 ;
	    RECT 928.2000 1220.4000 929.4000 1220.5500 ;
	    RECT 930.6000 1220.4000 931.8000 1220.5500 ;
	    RECT 947.4000 1221.4501 948.6000 1221.6000 ;
	    RECT 971.4000 1221.4501 972.6000 1221.6000 ;
	    RECT 947.4000 1220.5500 972.6000 1221.4501 ;
	    RECT 947.4000 1220.4000 948.6000 1220.5500 ;
	    RECT 971.4000 1220.4000 972.6000 1220.5500 ;
	    RECT 973.8000 1220.4000 975.0000 1221.6000 ;
	    RECT 975.9000 1220.4000 977.7000 1221.6000 ;
	    RECT 979.8000 1220.7001 980.1000 1222.2001 ;
	    RECT 1014.6000 1221.6000 1015.5000 1223.7001 ;
	    RECT 1017.3000 1223.1000 1022.7000 1223.7001 ;
	    RECT 1036.2001 1222.5000 1037.4000 1229.7001 ;
	    RECT 1038.6000 1226.7001 1039.8000 1229.7001 ;
	    RECT 1038.6000 1225.5000 1039.8000 1225.8000 ;
	    RECT 1038.6000 1223.4000 1039.8000 1224.6000 ;
	    RECT 1053.0000 1222.5000 1054.2001 1229.7001 ;
	    RECT 1055.4000 1226.7001 1056.6000 1229.7001 ;
	    RECT 1055.4000 1225.5000 1056.6000 1225.8000 ;
	    RECT 1055.4000 1224.4501 1056.6000 1224.6000 ;
	    RECT 1057.8000 1224.4501 1059.0000 1224.6000 ;
	    RECT 1055.4000 1223.5500 1059.0000 1224.4501 ;
	    RECT 1055.4000 1223.4000 1056.6000 1223.5500 ;
	    RECT 1057.8000 1223.4000 1059.0000 1223.5500 ;
	    RECT 1067.4000 1222.5000 1068.6000 1229.7001 ;
	    RECT 1069.8000 1226.7001 1071.0000 1229.7001 ;
	    RECT 1084.2001 1226.7001 1085.4000 1229.7001 ;
	    RECT 1069.8000 1225.5000 1071.0000 1225.8000 ;
	    RECT 1084.2001 1225.5000 1085.4000 1225.8000 ;
	    RECT 1069.8000 1223.4000 1071.0000 1224.6000 ;
	    RECT 1084.2001 1223.4000 1085.4000 1224.6000 ;
	    RECT 1086.6000 1222.5000 1087.8000 1229.7001 ;
	    RECT 1110.6000 1224.0000 1111.8000 1229.7001 ;
	    RECT 1113.0000 1224.9000 1114.2001 1229.7001 ;
	    RECT 1115.4000 1224.0000 1116.6000 1229.7001 ;
	    RECT 1110.6000 1223.7001 1116.6000 1224.0000 ;
	    RECT 1117.8000 1223.7001 1119.0000 1229.7001 ;
	    RECT 1110.9000 1223.1000 1116.3000 1223.7001 ;
	    RECT 1117.8000 1222.5000 1118.7001 1223.7001 ;
	    RECT 1194.6000 1222.5000 1195.8000 1229.7001 ;
	    RECT 1197.0000 1223.7001 1198.2001 1229.7001 ;
	    RECT 1201.2001 1227.6000 1202.4000 1229.7001 ;
	    RECT 1199.4000 1226.7001 1202.4000 1227.6000 ;
	    RECT 1205.1000 1226.7001 1206.6000 1229.7001 ;
	    RECT 1207.8000 1226.7001 1209.0000 1229.7001 ;
	    RECT 1210.2001 1226.7001 1211.4000 1229.7001 ;
	    RECT 1214.1000 1227.6000 1215.9000 1229.7001 ;
	    RECT 1213.8000 1226.7001 1215.9000 1227.6000 ;
	    RECT 1199.4000 1225.5000 1200.6000 1226.7001 ;
	    RECT 1207.8000 1225.8000 1208.7001 1226.7001 ;
	    RECT 1201.8000 1224.6000 1203.0000 1225.8000 ;
	    RECT 1204.5000 1224.9000 1208.7001 1225.8000 ;
	    RECT 1213.8000 1225.5000 1215.0000 1226.7001 ;
	    RECT 1204.5000 1224.6000 1205.7001 1224.9000 ;
	    RECT 981.0000 1221.4501 982.2000 1221.6000 ;
	    RECT 985.8000 1221.4501 987.0000 1221.6000 ;
	    RECT 981.0000 1220.5500 987.0000 1221.4501 ;
	    RECT 981.0000 1220.4000 982.2000 1220.5500 ;
	    RECT 985.8000 1220.4000 987.0000 1220.5500 ;
	    RECT 1012.2000 1220.4000 1013.4000 1221.6000 ;
	    RECT 1014.6000 1220.7001 1016.1000 1221.6000 ;
	    RECT 1017.0000 1220.4000 1018.2000 1221.6000 ;
	    RECT 1020.6000 1220.7001 1020.9000 1222.2001 ;
	    RECT 1021.8000 1221.4501 1023.0000 1221.6000 ;
	    RECT 1036.2001 1221.4501 1037.4000 1221.6000 ;
	    RECT 1021.8000 1220.5500 1037.4000 1221.4501 ;
	    RECT 1021.8000 1220.4000 1023.0000 1220.5500 ;
	    RECT 1036.2001 1220.4000 1037.4000 1220.5500 ;
	    RECT 1053.0000 1220.4000 1054.2001 1221.6000 ;
	    RECT 1060.2001 1221.4501 1061.4000 1221.6000 ;
	    RECT 1067.4000 1221.4501 1068.6000 1221.6000 ;
	    RECT 1060.2001 1220.5500 1068.6000 1221.4501 ;
	    RECT 1060.2001 1220.4000 1061.4000 1220.5500 ;
	    RECT 1067.4000 1220.4000 1068.6000 1220.5500 ;
	    RECT 1086.6000 1221.4501 1087.8000 1221.6000 ;
	    RECT 1086.6000 1220.5500 1106.8500 1221.4501 ;
	    RECT 1086.6000 1220.4000 1087.8000 1220.5500 ;
	    RECT 906.6000 1218.4501 907.8000 1218.6000 ;
	    RECT 925.8000 1218.4501 927.0000 1218.6000 ;
	    RECT 906.6000 1217.5500 927.0000 1218.4501 ;
	    RECT 906.6000 1217.4000 907.8000 1217.5500 ;
	    RECT 925.8000 1217.4000 927.0000 1217.5500 ;
	    RECT 928.2000 1217.4000 929.4000 1218.6000 ;
	    RECT 841.8000 1214.1000 843.0000 1214.4000 ;
	    RECT 834.9000 1213.5000 843.0000 1214.1000 ;
	    RECT 833.7000 1213.2001 843.0000 1213.5000 ;
	    RECT 844.5000 1213.5000 857.4000 1214.4000 ;
	    RECT 829.8000 1212.0000 832.2000 1213.2001 ;
	    RECT 833.7000 1212.3000 835.8000 1213.2001 ;
	    RECT 844.5000 1212.3000 845.4000 1213.5000 ;
	    RECT 856.2000 1213.2001 857.4000 1213.5000 ;
	    RECT 861.0000 1213.5000 874.5000 1214.4000 ;
	    RECT 875.4000 1215.0000 876.9000 1216.2001 ;
	    RECT 875.4000 1213.5000 876.6000 1215.0000 ;
	    RECT 861.0000 1213.2001 862.2000 1213.5000 ;
	    RECT 831.3000 1211.4000 832.2000 1212.0000 ;
	    RECT 836.7000 1211.4000 845.4000 1212.3000 ;
	    RECT 846.3000 1211.4000 850.2000 1212.6000 ;
	    RECT 827.4000 1210.2001 830.4000 1211.1000 ;
	    RECT 831.3000 1210.2001 837.6000 1211.4000 ;
	    RECT 829.5000 1209.3000 830.4000 1210.2001 ;
	    RECT 700.2000 1203.3000 701.4000 1209.3000 ;
	    RECT 827.4000 1203.3000 828.6000 1209.3000 ;
	    RECT 829.5000 1208.4000 831.0000 1209.3000 ;
	    RECT 829.8000 1203.3000 831.0000 1208.4000 ;
	    RECT 832.2000 1202.4000 833.4000 1209.3000 ;
	    RECT 834.6000 1203.3000 835.8000 1210.2001 ;
	    RECT 837.0000 1203.3000 838.2000 1209.3000 ;
	    RECT 839.4000 1203.3000 840.6000 1207.5000 ;
	    RECT 841.8000 1203.3000 843.0000 1207.5000 ;
	    RECT 844.2000 1203.3000 845.4000 1210.5000 ;
	    RECT 846.6000 1203.3000 847.8000 1209.3000 ;
	    RECT 849.0000 1203.3000 850.2000 1210.5000 ;
	    RECT 851.4000 1203.3000 852.6000 1209.3000 ;
	    RECT 853.8000 1203.3000 855.0000 1212.6000 ;
	    RECT 865.8000 1211.4000 869.7000 1212.6000 ;
	    RECT 858.6000 1210.2001 864.9000 1211.4000 ;
	    RECT 856.2000 1203.3000 857.4000 1207.5000 ;
	    RECT 858.6000 1203.3000 859.8000 1207.5000 ;
	    RECT 861.0000 1203.3000 862.2000 1207.5000 ;
	    RECT 863.4000 1203.3000 864.6000 1209.3000 ;
	    RECT 865.8000 1203.3000 867.0000 1211.4000 ;
	    RECT 873.6000 1211.1000 874.5000 1213.5000 ;
	    RECT 875.4000 1211.4000 876.6000 1212.6000 ;
	    RECT 870.6000 1210.2001 874.5000 1211.1000 ;
	    RECT 868.2000 1203.3000 869.4000 1209.3000 ;
	    RECT 870.6000 1203.3000 871.8000 1210.2001 ;
	    RECT 873.0000 1203.3000 874.2000 1209.3000 ;
	    RECT 875.4000 1203.3000 876.6000 1210.5000 ;
	    RECT 877.8000 1203.3000 879.0000 1209.3000 ;
	    RECT 904.2000 1203.3000 905.4000 1209.3000 ;
	    RECT 906.6000 1203.3000 907.8000 1216.5000 ;
	    RECT 928.2000 1216.2001 929.4000 1216.5000 ;
	    RECT 909.0000 1214.4000 910.2000 1215.6000 ;
	    RECT 930.6000 1215.3000 931.5000 1219.5000 ;
	    RECT 929.1000 1214.1000 931.8000 1215.3000 ;
	    RECT 909.0000 1213.2001 910.2000 1213.5000 ;
	    RECT 909.0000 1203.3000 910.2000 1209.3000 ;
	    RECT 929.1000 1203.3000 930.3000 1214.1000 ;
	    RECT 933.0000 1203.3000 934.2000 1215.3000 ;
	    RECT 945.0000 1203.3000 946.2000 1209.3000 ;
	    RECT 947.4000 1203.3000 948.6000 1219.5000 ;
	    RECT 949.8000 1218.4501 951.0000 1218.6000 ;
	    RECT 959.4000 1218.4501 960.6000 1218.6000 ;
	    RECT 949.8000 1217.5500 960.6000 1218.4501 ;
	    RECT 949.8000 1217.4000 951.0000 1217.5500 ;
	    RECT 959.4000 1217.4000 960.6000 1217.5500 ;
	    RECT 966.6000 1215.4501 967.8000 1215.6000 ;
	    RECT 971.4000 1215.4501 972.6000 1215.6000 ;
	    RECT 966.6000 1214.5500 972.6000 1215.4501 ;
	    RECT 966.6000 1214.4000 967.8000 1214.5500 ;
	    RECT 971.4000 1214.4000 972.6000 1214.5500 ;
	    RECT 973.8000 1214.4000 975.0000 1215.6000 ;
	    RECT 976.8000 1215.3000 977.7000 1220.4000 ;
	    RECT 978.6000 1219.5000 979.8000 1219.8000 ;
	    RECT 1014.6000 1219.5000 1015.8000 1219.8000 ;
	    RECT 1019.4000 1219.5000 1020.6000 1219.8000 ;
	    RECT 1012.2000 1219.2001 1013.4000 1219.5000 ;
	    RECT 978.6000 1217.4000 979.8000 1218.6000 ;
	    RECT 1014.6000 1217.4000 1015.8000 1218.6000 ;
	    RECT 1017.3000 1215.3000 1018.2000 1219.5000 ;
	    RECT 1019.4000 1218.4501 1020.6000 1218.6000 ;
	    RECT 1024.2001 1218.4501 1025.4000 1218.6000 ;
	    RECT 1019.4000 1217.5500 1025.4000 1218.4501 ;
	    RECT 1019.4000 1217.4000 1020.6000 1217.5500 ;
	    RECT 1024.2001 1217.4000 1025.4000 1217.5500 ;
	    RECT 976.8000 1214.4000 978.3000 1215.3000 ;
	    RECT 975.0000 1212.6000 975.9000 1213.5000 ;
	    RECT 975.0000 1211.4000 976.2000 1212.6000 ;
	    RECT 974.7000 1203.3000 975.9000 1209.3000 ;
	    RECT 977.1000 1203.3000 978.3000 1214.4000 ;
	    RECT 981.0000 1203.3000 982.2000 1215.3000 ;
	    RECT 1012.2000 1203.3000 1013.4000 1215.3000 ;
	    RECT 1016.1000 1203.3000 1019.1000 1215.3000 ;
	    RECT 1021.8000 1203.3000 1023.0000 1215.3000 ;
	    RECT 1036.2001 1203.3000 1037.4000 1219.5000 ;
	    RECT 1038.6000 1203.3000 1039.8000 1209.3000 ;
	    RECT 1053.0000 1203.3000 1054.2001 1219.5000 ;
	    RECT 1055.4000 1203.3000 1056.6000 1209.3000 ;
	    RECT 1067.4000 1203.3000 1068.6000 1219.5000 ;
	    RECT 1069.8000 1203.3000 1071.0000 1209.3000 ;
	    RECT 1084.2001 1203.3000 1085.4000 1209.3000 ;
	    RECT 1086.6000 1203.3000 1087.8000 1219.5000 ;
	    RECT 1105.9501 1218.4501 1106.8500 1220.5500 ;
	    RECT 1110.6000 1220.4000 1111.8000 1221.6000 ;
	    RECT 1112.7001 1220.7001 1113.0000 1222.2001 ;
	    RECT 1115.1000 1220.4000 1116.9000 1221.6000 ;
	    RECT 1117.8000 1221.4501 1119.0000 1221.6000 ;
	    RECT 1192.2001 1221.4501 1193.4000 1221.6000 ;
	    RECT 1117.8000 1220.5500 1193.4000 1221.4501 ;
	    RECT 1117.8000 1220.4000 1119.0000 1220.5500 ;
	    RECT 1192.2001 1220.4000 1193.4000 1220.5500 ;
	    RECT 1195.8000 1220.4000 1196.1000 1221.6000 ;
	    RECT 1197.0000 1220.4000 1198.2001 1221.6000 ;
	    RECT 1202.1000 1221.3000 1203.0000 1224.6000 ;
	    RECT 1218.6000 1224.0000 1219.8000 1229.7001 ;
	    RECT 1216.5000 1223.1000 1217.7001 1223.4000 ;
	    RECT 1221.0000 1223.1000 1222.2001 1229.7001 ;
	    RECT 1233.0000 1226.7001 1234.2001 1229.7001 ;
	    RECT 1233.0000 1225.5000 1234.2001 1225.8000 ;
	    RECT 1233.0000 1223.4000 1234.2001 1224.6000 ;
	    RECT 1216.5000 1222.2001 1222.2001 1223.1000 ;
	    RECT 1235.4000 1222.5000 1236.6000 1229.7001 ;
	    RECT 1210.5000 1221.3000 1211.7001 1221.6000 ;
	    RECT 1199.1000 1220.4000 1212.3000 1221.3000 ;
	    RECT 1113.0000 1219.5000 1114.2001 1219.8000 ;
	    RECT 1113.0000 1218.4501 1114.2001 1218.6000 ;
	    RECT 1105.9501 1217.5500 1114.2001 1218.4501 ;
	    RECT 1113.0000 1217.4000 1114.2001 1217.5500 ;
	    RECT 1115.1000 1215.3000 1116.0000 1220.4000 ;
	    RECT 1200.3000 1220.1000 1201.5000 1220.4000 ;
	    RECT 1197.9000 1218.6000 1199.1000 1218.9000 ;
	    RECT 1197.9000 1217.7001 1203.3000 1218.6000 ;
	    RECT 1204.2001 1217.4000 1205.4000 1218.6000 ;
	    RECT 1194.6000 1216.5000 1203.0000 1216.8000 ;
	    RECT 1194.6000 1216.2001 1203.3000 1216.5000 ;
	    RECT 1194.6000 1215.9000 1209.3000 1216.2001 ;
	    RECT 1110.6000 1203.3000 1111.8000 1215.3000 ;
	    RECT 1114.5000 1214.4000 1116.0000 1215.3000 ;
	    RECT 1117.8000 1215.4501 1119.0000 1215.6000 ;
	    RECT 1134.6000 1215.4501 1135.8000 1215.6000 ;
	    RECT 1117.8000 1214.5500 1135.8000 1215.4501 ;
	    RECT 1117.8000 1214.4000 1119.0000 1214.5500 ;
	    RECT 1134.6000 1214.4000 1135.8000 1214.5500 ;
	    RECT 1114.5000 1203.3000 1115.7001 1214.4000 ;
	    RECT 1116.9000 1212.6000 1117.8000 1213.5000 ;
	    RECT 1116.6000 1211.4000 1117.8000 1212.6000 ;
	    RECT 1116.9000 1203.3000 1118.1000 1209.3000 ;
	    RECT 1194.6000 1203.3000 1195.8000 1215.9000 ;
	    RECT 1202.1000 1215.3000 1209.3000 1215.9000 ;
	    RECT 1197.0000 1203.3000 1198.2001 1215.0000 ;
	    RECT 1199.4000 1213.5000 1207.5000 1214.4000 ;
	    RECT 1199.4000 1213.2001 1200.6000 1213.5000 ;
	    RECT 1206.3000 1213.2001 1207.5000 1213.5000 ;
	    RECT 1208.4000 1213.5000 1209.3000 1215.3000 ;
	    RECT 1211.4000 1215.6000 1212.3000 1220.4000 ;
	    RECT 1221.0000 1219.5000 1222.2001 1222.2001 ;
	    RECT 1235.4000 1221.4501 1236.6000 1221.6000 ;
	    RECT 1343.4000 1221.4501 1344.6000 1221.6000 ;
	    RECT 1235.4000 1220.5500 1344.6000 1221.4501 ;
	    RECT 1235.4000 1220.4000 1236.6000 1220.5500 ;
	    RECT 1343.4000 1220.4000 1344.6000 1220.5500 ;
	    RECT 1367.4000 1220.7001 1368.6000 1229.7001 ;
	    RECT 1372.2001 1223.7001 1373.4000 1229.7001 ;
	    RECT 1377.0000 1224.9000 1378.2001 1229.7001 ;
	    RECT 1379.4000 1225.5000 1380.6000 1229.7001 ;
	    RECT 1381.8000 1225.5000 1383.0000 1229.7001 ;
	    RECT 1384.2001 1225.5000 1385.4000 1229.7001 ;
	    RECT 1386.6000 1226.7001 1387.8000 1229.7001 ;
	    RECT 1389.0000 1225.5000 1390.2001 1229.7001 ;
	    RECT 1391.4000 1226.7001 1392.6000 1229.7001 ;
	    RECT 1393.8000 1225.5000 1395.0000 1229.7001 ;
	    RECT 1396.2001 1225.5000 1397.4000 1229.7001 ;
	    RECT 1398.6000 1225.5000 1399.8000 1229.7001 ;
	    RECT 1401.0000 1225.5000 1402.2001 1229.7001 ;
	    RECT 1374.3000 1223.7001 1378.2001 1224.9000 ;
	    RECT 1403.4000 1224.9000 1404.6000 1229.7001 ;
	    RECT 1383.3000 1223.7001 1390.2001 1224.6000 ;
	    RECT 1374.3000 1222.8000 1375.5000 1223.7001 ;
	    RECT 1371.0000 1221.6000 1375.5000 1222.8000 ;
	    RECT 1367.4000 1219.5000 1380.6000 1220.7001 ;
	    RECT 1383.3000 1220.1000 1384.5000 1223.7001 ;
	    RECT 1389.0000 1223.4000 1390.2001 1223.7001 ;
	    RECT 1391.4000 1223.4000 1392.6000 1224.6000 ;
	    RECT 1393.5000 1223.4000 1393.8000 1224.6000 ;
	    RECT 1398.3000 1223.4000 1399.8000 1224.6000 ;
	    RECT 1403.4000 1223.7001 1407.0000 1224.9000 ;
	    RECT 1408.2001 1223.7001 1409.4000 1229.7001 ;
	    RECT 1386.6000 1222.5000 1387.8000 1222.8000 ;
	    RECT 1389.0000 1222.2001 1390.2001 1222.5000 ;
	    RECT 1386.6000 1220.4000 1387.8000 1221.6000 ;
	    RECT 1389.0000 1221.3000 1395.6000 1222.2001 ;
	    RECT 1394.4000 1221.0000 1395.6000 1221.3000 ;
	    RECT 1213.8000 1219.2001 1215.0000 1219.5000 ;
	    RECT 1213.8000 1218.3000 1219.5000 1219.2001 ;
	    RECT 1218.3000 1218.0000 1219.5000 1218.3000 ;
	    RECT 1221.0000 1217.4000 1222.2001 1218.6000 ;
	    RECT 1215.9000 1217.1000 1217.1000 1217.4000 ;
	    RECT 1215.9000 1216.5000 1220.1000 1217.1000 ;
	    RECT 1215.9000 1216.2001 1222.2001 1216.5000 ;
	    RECT 1211.4000 1214.7001 1215.0000 1215.6000 ;
	    RECT 1210.5000 1213.5000 1211.7001 1213.8000 ;
	    RECT 1208.4000 1212.6000 1211.7001 1213.5000 ;
	    RECT 1214.1000 1213.2001 1215.0000 1214.7001 ;
	    RECT 1214.1000 1212.0000 1216.2001 1213.2001 ;
	    RECT 1204.5000 1211.1000 1205.7001 1211.4000 ;
	    RECT 1208.7001 1211.1000 1209.9000 1211.4000 ;
	    RECT 1199.4000 1209.3000 1200.6000 1210.5000 ;
	    RECT 1204.5000 1210.2001 1209.9000 1211.1000 ;
	    RECT 1207.8000 1209.3000 1208.7001 1210.2001 ;
	    RECT 1213.8000 1209.3000 1215.0000 1210.5000 ;
	    RECT 1199.4000 1208.4000 1202.4000 1209.3000 ;
	    RECT 1201.2001 1203.3000 1202.4000 1208.4000 ;
	    RECT 1205.4000 1203.3000 1206.6000 1209.3000 ;
	    RECT 1207.8000 1203.3000 1209.0000 1209.3000 ;
	    RECT 1210.2001 1203.3000 1211.4000 1209.3000 ;
	    RECT 1214.1000 1203.3000 1215.9000 1209.3000 ;
	    RECT 1218.6000 1203.3000 1219.8000 1215.3000 ;
	    RECT 1221.0000 1203.3000 1222.2001 1216.2001 ;
	    RECT 1233.0000 1203.3000 1234.2001 1209.3000 ;
	    RECT 1235.4000 1203.3000 1236.6000 1219.5000 ;
	    RECT 1367.4000 1211.1000 1368.6000 1219.5000 ;
	    RECT 1381.5000 1218.9000 1384.5000 1220.1000 ;
	    RECT 1390.2001 1218.9000 1395.0000 1220.1000 ;
	    RECT 1398.6000 1219.2001 1399.8000 1223.4000 ;
	    RECT 1405.8000 1222.8000 1407.0000 1223.7001 ;
	    RECT 1405.8000 1221.9000 1408.5000 1222.8000 ;
	    RECT 1407.3000 1220.1000 1408.5000 1221.9000 ;
	    RECT 1413.0000 1221.9000 1414.2001 1229.7001 ;
	    RECT 1415.4000 1224.0000 1416.6000 1229.7001 ;
	    RECT 1417.8000 1226.7001 1419.0000 1229.7001 ;
	    RECT 1429.8000 1226.7001 1431.0000 1229.7001 ;
	    RECT 1429.8000 1225.5000 1431.0000 1225.8000 ;
	    RECT 1417.8000 1224.4501 1419.0000 1224.6000 ;
	    RECT 1429.8000 1224.4501 1431.0000 1224.6000 ;
	    RECT 1415.4000 1222.8000 1416.9000 1224.0000 ;
	    RECT 1417.8000 1223.5500 1431.0000 1224.4501 ;
	    RECT 1417.8000 1223.4000 1419.0000 1223.5500 ;
	    RECT 1429.8000 1223.4000 1431.0000 1223.5500 ;
	    RECT 1413.0000 1221.0000 1414.8000 1221.9000 ;
	    RECT 1407.3000 1218.9000 1413.0000 1220.1000 ;
	    RECT 1369.5000 1218.0000 1370.7001 1218.3000 ;
	    RECT 1369.5000 1217.1000 1376.1000 1218.0000 ;
	    RECT 1377.0000 1217.4000 1378.2001 1218.6000 ;
	    RECT 1403.4000 1218.0000 1404.6000 1218.9000 ;
	    RECT 1413.9000 1218.0000 1414.8000 1221.0000 ;
	    RECT 1379.1000 1217.1000 1404.6000 1218.0000 ;
	    RECT 1413.6000 1217.1000 1414.8000 1218.0000 ;
	    RECT 1411.5000 1216.2001 1412.7001 1216.5000 ;
	    RECT 1372.2001 1214.4000 1373.4000 1215.6000 ;
	    RECT 1374.3000 1215.3000 1412.7001 1216.2001 ;
	    RECT 1377.3000 1215.0000 1378.5000 1215.3000 ;
	    RECT 1413.6000 1214.4000 1414.5000 1217.1000 ;
	    RECT 1415.7001 1216.2001 1416.9000 1222.8000 ;
	    RECT 1432.2001 1222.5000 1433.4000 1229.7001 ;
	    RECT 1451.4000 1223.7001 1452.6000 1229.7001 ;
	    RECT 1455.3000 1224.6000 1456.5000 1229.7001 ;
	    RECT 1453.8000 1223.7001 1456.5000 1224.6000 ;
	    RECT 1451.4000 1222.5000 1452.6000 1222.8000 ;
	    RECT 1422.6000 1221.4501 1423.8000 1221.6000 ;
	    RECT 1432.2001 1221.4501 1433.4000 1221.6000 ;
	    RECT 1422.6000 1220.5500 1433.4000 1221.4501 ;
	    RECT 1422.6000 1220.4000 1423.8000 1220.5500 ;
	    RECT 1432.2001 1220.4000 1433.4000 1220.5500 ;
	    RECT 1451.4000 1220.4000 1452.6000 1221.6000 ;
	    RECT 1453.8000 1219.5000 1455.0000 1223.7001 ;
	    RECT 1525.8000 1222.5000 1527.0000 1229.7001 ;
	    RECT 1528.2001 1223.7001 1529.4000 1229.7001 ;
	    RECT 1532.4000 1227.6000 1533.6000 1229.7001 ;
	    RECT 1530.6000 1226.7001 1533.6000 1227.6000 ;
	    RECT 1536.3000 1226.7001 1537.8000 1229.7001 ;
	    RECT 1539.0000 1226.7001 1540.2001 1229.7001 ;
	    RECT 1541.4000 1226.7001 1542.6000 1229.7001 ;
	    RECT 1545.3000 1227.6000 1547.1000 1229.7001 ;
	    RECT 1545.0000 1226.7001 1547.1000 1227.6000 ;
	    RECT 1530.6000 1225.5000 1531.8000 1226.7001 ;
	    RECT 1539.0000 1225.8000 1539.9000 1226.7001 ;
	    RECT 1533.0000 1224.6000 1534.2001 1225.8000 ;
	    RECT 1535.7001 1224.9000 1539.9000 1225.8000 ;
	    RECT 1545.0000 1225.5000 1546.2001 1226.7001 ;
	    RECT 1535.7001 1224.6000 1536.9000 1224.9000 ;
	    RECT 1527.0000 1220.4000 1527.3000 1221.6000 ;
	    RECT 1528.2001 1220.4000 1529.4000 1221.6000 ;
	    RECT 1533.3000 1221.3000 1534.2001 1224.6000 ;
	    RECT 1549.8000 1224.0000 1551.0000 1229.7001 ;
	    RECT 1547.7001 1223.1000 1548.9000 1223.4000 ;
	    RECT 1552.2001 1223.1000 1553.4000 1229.7001 ;
	    RECT 1547.7001 1222.2001 1553.4000 1223.1000 ;
	    RECT 1541.7001 1221.3000 1542.9000 1221.6000 ;
	    RECT 1530.3000 1220.4000 1543.5000 1221.3000 ;
	    RECT 1531.5000 1220.1000 1532.7001 1220.4000 ;
	    RECT 1381.8000 1214.1000 1383.0000 1214.4000 ;
	    RECT 1374.9000 1213.5000 1383.0000 1214.1000 ;
	    RECT 1373.7001 1213.2001 1383.0000 1213.5000 ;
	    RECT 1384.5000 1213.5000 1397.4000 1214.4000 ;
	    RECT 1369.8000 1212.0000 1372.2001 1213.2001 ;
	    RECT 1373.7001 1212.3000 1375.8000 1213.2001 ;
	    RECT 1384.5000 1212.3000 1385.4000 1213.5000 ;
	    RECT 1396.2001 1213.2001 1397.4000 1213.5000 ;
	    RECT 1401.0000 1213.5000 1414.5000 1214.4000 ;
	    RECT 1415.4000 1215.0000 1416.9000 1216.2001 ;
	    RECT 1415.4000 1213.5000 1416.6000 1215.0000 ;
	    RECT 1401.0000 1213.2001 1402.2001 1213.5000 ;
	    RECT 1371.3000 1211.4000 1372.2001 1212.0000 ;
	    RECT 1376.7001 1211.4000 1385.4000 1212.3000 ;
	    RECT 1386.3000 1211.4000 1390.2001 1212.6000 ;
	    RECT 1367.4000 1210.2001 1370.4000 1211.1000 ;
	    RECT 1371.3000 1210.2001 1377.6000 1211.4000 ;
	    RECT 1369.5000 1209.3000 1370.4000 1210.2001 ;
	    RECT 1367.4000 1203.3000 1368.6000 1209.3000 ;
	    RECT 1369.5000 1208.4000 1371.0000 1209.3000 ;
	    RECT 1369.8000 1203.3000 1371.0000 1208.4000 ;
	    RECT 1372.2001 1202.4000 1373.4000 1209.3000 ;
	    RECT 1374.6000 1203.3000 1375.8000 1210.2001 ;
	    RECT 1377.0000 1203.3000 1378.2001 1209.3000 ;
	    RECT 1379.4000 1203.3000 1380.6000 1207.5000 ;
	    RECT 1381.8000 1203.3000 1383.0000 1207.5000 ;
	    RECT 1384.2001 1203.3000 1385.4000 1210.5000 ;
	    RECT 1386.6000 1203.3000 1387.8000 1209.3000 ;
	    RECT 1389.0000 1203.3000 1390.2001 1210.5000 ;
	    RECT 1391.4000 1203.3000 1392.6000 1209.3000 ;
	    RECT 1393.8000 1203.3000 1395.0000 1212.6000 ;
	    RECT 1405.8000 1211.4000 1409.7001 1212.6000 ;
	    RECT 1398.6000 1210.2001 1404.9000 1211.4000 ;
	    RECT 1396.2001 1203.3000 1397.4000 1207.5000 ;
	    RECT 1398.6000 1203.3000 1399.8000 1207.5000 ;
	    RECT 1401.0000 1203.3000 1402.2001 1207.5000 ;
	    RECT 1403.4000 1203.3000 1404.6000 1209.3000 ;
	    RECT 1405.8000 1203.3000 1407.0000 1211.4000 ;
	    RECT 1413.6000 1211.1000 1414.5000 1213.5000 ;
	    RECT 1415.4000 1211.4000 1416.6000 1212.6000 ;
	    RECT 1410.6000 1210.2001 1414.5000 1211.1000 ;
	    RECT 1408.2001 1203.3000 1409.4000 1209.3000 ;
	    RECT 1410.6000 1203.3000 1411.8000 1210.2001 ;
	    RECT 1413.0000 1203.3000 1414.2001 1209.3000 ;
	    RECT 1415.4000 1203.3000 1416.6000 1210.5000 ;
	    RECT 1417.8000 1203.3000 1419.0000 1209.3000 ;
	    RECT 1429.8000 1203.3000 1431.0000 1209.3000 ;
	    RECT 1432.2001 1203.3000 1433.4000 1219.5000 ;
	    RECT 1529.1000 1218.6000 1530.3000 1218.9000 ;
	    RECT 1453.8000 1217.4000 1455.0000 1218.6000 ;
	    RECT 1529.1000 1217.7001 1534.5000 1218.6000 ;
	    RECT 1535.4000 1217.4000 1536.6000 1218.6000 ;
	    RECT 1525.8000 1216.5000 1534.2001 1216.8000 ;
	    RECT 1451.4000 1203.3000 1452.6000 1209.3000 ;
	    RECT 1453.8000 1203.3000 1455.0000 1216.5000 ;
	    RECT 1525.8000 1216.2001 1534.5000 1216.5000 ;
	    RECT 1525.8000 1215.9000 1540.5000 1216.2001 ;
	    RECT 1456.2001 1215.4501 1457.4000 1215.6000 ;
	    RECT 1463.4000 1215.4501 1464.6000 1215.6000 ;
	    RECT 1456.2001 1214.5500 1464.6000 1215.4501 ;
	    RECT 1456.2001 1214.4000 1457.4000 1214.5500 ;
	    RECT 1463.4000 1214.4000 1464.6000 1214.5500 ;
	    RECT 1456.2001 1213.2001 1457.4000 1213.5000 ;
	    RECT 1509.0000 1212.4501 1510.2001 1212.6000 ;
	    RECT 1523.4000 1212.4501 1524.6000 1212.6000 ;
	    RECT 1509.0000 1211.5500 1524.6000 1212.4501 ;
	    RECT 1509.0000 1211.4000 1510.2001 1211.5500 ;
	    RECT 1523.4000 1211.4000 1524.6000 1211.5500 ;
	    RECT 1456.2001 1203.3000 1457.4000 1209.3000 ;
	    RECT 1525.8000 1203.3000 1527.0000 1215.9000 ;
	    RECT 1533.3000 1215.3000 1540.5000 1215.9000 ;
	    RECT 1528.2001 1203.3000 1529.4000 1215.0000 ;
	    RECT 1530.6000 1213.5000 1538.7001 1214.4000 ;
	    RECT 1530.6000 1213.2001 1531.8000 1213.5000 ;
	    RECT 1537.5000 1213.2001 1538.7001 1213.5000 ;
	    RECT 1539.6000 1213.5000 1540.5000 1215.3000 ;
	    RECT 1542.6000 1215.6000 1543.5000 1220.4000 ;
	    RECT 1552.2001 1219.5000 1553.4000 1222.2001 ;
	    RECT 1545.0000 1219.2001 1546.2001 1219.5000 ;
	    RECT 1545.0000 1218.3000 1550.7001 1219.2001 ;
	    RECT 1549.5000 1218.0000 1550.7001 1218.3000 ;
	    RECT 1552.2001 1217.4000 1553.4000 1218.6000 ;
	    RECT 1547.1000 1217.1000 1548.3000 1217.4000 ;
	    RECT 1547.1000 1216.5000 1551.3000 1217.1000 ;
	    RECT 1547.1000 1216.2001 1553.4000 1216.5000 ;
	    RECT 1542.6000 1214.7001 1546.2001 1215.6000 ;
	    RECT 1541.7001 1213.5000 1542.9000 1213.8000 ;
	    RECT 1539.6000 1212.6000 1542.9000 1213.5000 ;
	    RECT 1545.3000 1213.2001 1546.2001 1214.7001 ;
	    RECT 1545.3000 1212.0000 1547.4000 1213.2001 ;
	    RECT 1535.7001 1211.1000 1536.9000 1211.4000 ;
	    RECT 1539.9000 1211.1000 1541.1000 1211.4000 ;
	    RECT 1530.6000 1209.3000 1531.8000 1210.5000 ;
	    RECT 1535.7001 1210.2001 1541.1000 1211.1000 ;
	    RECT 1539.0000 1209.3000 1539.9000 1210.2001 ;
	    RECT 1545.0000 1209.3000 1546.2001 1210.5000 ;
	    RECT 1530.6000 1208.4000 1533.6000 1209.3000 ;
	    RECT 1532.4000 1203.3000 1533.6000 1208.4000 ;
	    RECT 1536.6000 1203.3000 1537.8000 1209.3000 ;
	    RECT 1539.0000 1203.3000 1540.2001 1209.3000 ;
	    RECT 1541.4000 1203.3000 1542.6000 1209.3000 ;
	    RECT 1545.3000 1203.3000 1547.1000 1209.3000 ;
	    RECT 1549.8000 1203.3000 1551.0000 1215.3000 ;
	    RECT 1552.2001 1203.3000 1553.4000 1216.2001 ;
	    RECT 1.2000 1200.6000 1569.0000 1202.4000 ;
	    RECT 18.6000 1187.7001 19.8000 1199.7001 ;
	    RECT 21.0000 1189.5000 22.2000 1199.7001 ;
	    RECT 23.4000 1188.6000 24.6000 1199.7001 ;
	    RECT 21.3000 1187.7001 24.6000 1188.6000 ;
	    RECT 47.4000 1187.7001 48.6000 1199.7001 ;
	    RECT 51.3000 1188.6000 52.5000 1199.7001 ;
	    RECT 53.7000 1193.7001 54.9000 1199.7001 ;
	    RECT 53.4000 1190.4000 54.6000 1191.6000 ;
	    RECT 53.7000 1189.5000 54.6000 1190.4000 ;
	    RECT 73.8000 1188.6000 75.0000 1199.7001 ;
	    RECT 76.2000 1189.5000 77.4000 1199.7001 ;
	    RECT 51.3000 1187.7001 52.8000 1188.6000 ;
	    RECT 18.6000 1184.4000 19.5000 1187.7001 ;
	    RECT 21.3000 1186.8000 22.2000 1187.7001 ;
	    RECT 20.4000 1185.6000 22.2000 1186.8000 ;
	    RECT 18.6000 1183.5000 19.8000 1184.4000 ;
	    RECT 18.6000 1181.4000 19.8000 1182.6000 ;
	    RECT 21.3000 1181.1000 22.2000 1185.6000 ;
	    RECT 23.4000 1184.4000 24.6000 1185.6000 ;
	    RECT 49.8000 1184.4000 51.0000 1185.6000 ;
	    RECT 23.4000 1183.2001 24.6000 1183.5000 ;
	    RECT 49.8000 1183.2001 51.0000 1183.5000 ;
	    RECT 51.9000 1182.6000 52.8000 1187.7001 ;
	    RECT 54.6000 1188.4501 55.8000 1188.6000 ;
	    RECT 59.4000 1188.4501 60.6000 1188.6000 ;
	    RECT 54.6000 1187.5500 60.6000 1188.4501 ;
	    RECT 73.8000 1187.7001 77.1000 1188.6000 ;
	    RECT 78.6000 1187.7001 79.8000 1199.7001 ;
	    RECT 54.6000 1187.4000 55.8000 1187.5500 ;
	    RECT 59.4000 1187.4000 60.6000 1187.5500 ;
	    RECT 76.2000 1186.8000 77.1000 1187.7001 ;
	    RECT 76.2000 1185.6000 78.0000 1186.8000 ;
	    RECT 54.6000 1185.4501 55.8000 1185.6000 ;
	    RECT 73.8000 1185.4501 75.0000 1185.6000 ;
	    RECT 54.6000 1184.5500 75.0000 1185.4501 ;
	    RECT 54.6000 1184.4000 55.8000 1184.5500 ;
	    RECT 73.8000 1184.4000 75.0000 1184.5500 ;
	    RECT 73.8000 1183.2001 75.0000 1183.5000 ;
	    RECT 33.0000 1182.4501 34.2000 1182.6000 ;
	    RECT 47.4000 1182.4501 48.6000 1182.6000 ;
	    RECT 33.0000 1181.5500 48.6000 1182.4501 ;
	    RECT 33.0000 1181.4000 34.2000 1181.5500 ;
	    RECT 47.4000 1181.4000 48.6000 1181.5500 ;
	    RECT 18.6000 1173.3000 19.8000 1180.5000 ;
	    RECT 21.3000 1180.2001 24.6000 1181.1000 ;
	    RECT 49.5000 1180.8000 49.8000 1182.3000 ;
	    RECT 51.9000 1181.4000 53.7000 1182.6000 ;
	    RECT 54.6000 1182.4501 55.8000 1182.6000 ;
	    RECT 71.4000 1182.4501 72.6000 1182.6000 ;
	    RECT 54.6000 1181.5500 72.6000 1182.4501 ;
	    RECT 54.6000 1181.4000 55.8000 1181.5500 ;
	    RECT 71.4000 1181.4000 72.6000 1181.5500 ;
	    RECT 76.2000 1181.1000 77.1000 1185.6000 ;
	    RECT 78.9000 1184.4000 79.8000 1187.7001 ;
	    RECT 78.6000 1183.5000 79.8000 1184.4000 ;
	    RECT 93.0000 1183.5000 94.2000 1199.7001 ;
	    RECT 95.4000 1193.7001 96.6000 1199.7001 ;
	    RECT 114.6000 1193.7001 115.8000 1199.7001 ;
	    RECT 117.0000 1186.5000 118.2000 1199.7001 ;
	    RECT 119.4000 1193.7001 120.6000 1199.7001 ;
	    RECT 237.0000 1197.4501 238.2000 1197.6000 ;
	    RECT 246.6000 1197.4501 247.8000 1197.6000 ;
	    RECT 237.0000 1196.5500 247.8000 1197.4501 ;
	    RECT 237.0000 1196.4000 238.2000 1196.5500 ;
	    RECT 246.6000 1196.4000 247.8000 1196.5500 ;
	    RECT 251.4000 1193.7001 252.6000 1199.7001 ;
	    RECT 253.8000 1194.6000 255.0000 1199.7001 ;
	    RECT 253.5000 1193.7001 255.0000 1194.6000 ;
	    RECT 256.2000 1193.7001 257.4000 1200.6000 ;
	    RECT 253.5000 1192.8000 254.4000 1193.7001 ;
	    RECT 258.6000 1192.8000 259.8000 1199.7001 ;
	    RECT 261.0000 1193.7001 262.2000 1199.7001 ;
	    RECT 263.4000 1195.5000 264.6000 1199.7001 ;
	    RECT 265.8000 1195.5000 267.0000 1199.7001 ;
	    RECT 251.4000 1191.9000 254.4000 1192.8000 ;
	    RECT 119.4000 1189.5000 120.6000 1189.8000 ;
	    RECT 119.4000 1188.4501 120.6000 1188.6000 ;
	    RECT 172.2000 1188.4501 173.4000 1188.6000 ;
	    RECT 119.4000 1187.5500 173.4000 1188.4501 ;
	    RECT 119.4000 1187.4000 120.6000 1187.5500 ;
	    RECT 172.2000 1187.4000 173.4000 1187.5500 ;
	    RECT 95.4000 1185.4501 96.6000 1185.6000 ;
	    RECT 117.0000 1185.4501 118.2000 1185.6000 ;
	    RECT 95.4000 1184.5500 118.2000 1185.4501 ;
	    RECT 95.4000 1184.4000 96.6000 1184.5500 ;
	    RECT 117.0000 1184.4000 118.2000 1184.5500 ;
	    RECT 251.4000 1183.5000 252.6000 1191.9000 ;
	    RECT 255.3000 1191.6000 261.6000 1192.8000 ;
	    RECT 268.2000 1192.5000 269.4000 1199.7001 ;
	    RECT 270.6000 1193.7001 271.8000 1199.7001 ;
	    RECT 273.0000 1192.5000 274.2000 1199.7001 ;
	    RECT 275.4000 1193.7001 276.6000 1199.7001 ;
	    RECT 255.3000 1191.0000 256.2000 1191.6000 ;
	    RECT 253.8000 1189.8000 256.2000 1191.0000 ;
	    RECT 260.7000 1190.7001 269.4000 1191.6000 ;
	    RECT 257.7000 1189.8000 259.8000 1190.7001 ;
	    RECT 257.7000 1189.5000 267.0000 1189.8000 ;
	    RECT 258.9000 1188.9000 267.0000 1189.5000 ;
	    RECT 265.8000 1188.6000 267.0000 1188.9000 ;
	    RECT 268.5000 1189.5000 269.4000 1190.7001 ;
	    RECT 270.3000 1190.4000 274.2000 1191.6000 ;
	    RECT 277.8000 1190.4000 279.0000 1199.7001 ;
	    RECT 280.2000 1195.5000 281.4000 1199.7001 ;
	    RECT 282.6000 1195.5000 283.8000 1199.7001 ;
	    RECT 285.0000 1195.5000 286.2000 1199.7001 ;
	    RECT 287.4000 1193.7001 288.6000 1199.7001 ;
	    RECT 282.6000 1191.6000 288.9000 1192.8000 ;
	    RECT 289.8000 1191.6000 291.0000 1199.7001 ;
	    RECT 292.2000 1193.7001 293.4000 1199.7001 ;
	    RECT 294.6000 1192.8000 295.8000 1199.7001 ;
	    RECT 297.0000 1193.7001 298.2000 1199.7001 ;
	    RECT 294.6000 1191.9000 298.5000 1192.8000 ;
	    RECT 299.4000 1192.5000 300.6000 1199.7001 ;
	    RECT 301.8000 1193.7001 303.0000 1199.7001 ;
	    RECT 304.2000 1197.4501 305.4000 1197.6000 ;
	    RECT 359.4000 1197.4501 360.6000 1197.6000 ;
	    RECT 304.2000 1196.5500 360.6000 1197.4501 ;
	    RECT 304.2000 1196.4000 305.4000 1196.5500 ;
	    RECT 359.4000 1196.4000 360.6000 1196.5500 ;
	    RECT 436.2000 1193.7001 437.4000 1199.7001 ;
	    RECT 438.6000 1192.5000 439.8000 1199.7001 ;
	    RECT 441.0000 1193.7001 442.2000 1199.7001 ;
	    RECT 443.4000 1192.8000 444.6000 1199.7001 ;
	    RECT 445.8000 1193.7001 447.0000 1199.7001 ;
	    RECT 289.8000 1190.4000 293.7000 1191.6000 ;
	    RECT 280.2000 1189.5000 281.4000 1189.8000 ;
	    RECT 268.5000 1188.6000 281.4000 1189.5000 ;
	    RECT 285.0000 1189.5000 286.2000 1189.8000 ;
	    RECT 297.6000 1189.5000 298.5000 1191.9000 ;
	    RECT 440.7000 1191.9000 444.6000 1192.8000 ;
	    RECT 299.4000 1190.4000 300.6000 1191.6000 ;
	    RECT 357.0000 1191.4501 358.2000 1191.6000 ;
	    RECT 438.6000 1191.4501 439.8000 1191.6000 ;
	    RECT 357.0000 1190.5500 439.8000 1191.4501 ;
	    RECT 357.0000 1190.4000 358.2000 1190.5500 ;
	    RECT 438.6000 1190.4000 439.8000 1190.5500 ;
	    RECT 440.7000 1189.5000 441.6000 1191.9000 ;
	    RECT 448.2000 1191.6000 449.4000 1199.7001 ;
	    RECT 450.6000 1193.7001 451.8000 1199.7001 ;
	    RECT 453.0000 1195.5000 454.2000 1199.7001 ;
	    RECT 455.4000 1195.5000 456.6000 1199.7001 ;
	    RECT 457.8000 1195.5000 459.0000 1199.7001 ;
	    RECT 450.3000 1191.6000 456.6000 1192.8000 ;
	    RECT 445.5000 1190.4000 449.4000 1191.6000 ;
	    RECT 460.2000 1190.4000 461.4000 1199.7001 ;
	    RECT 462.6000 1193.7001 463.8000 1199.7001 ;
	    RECT 465.0000 1192.5000 466.2000 1199.7001 ;
	    RECT 467.4000 1193.7001 468.6000 1199.7001 ;
	    RECT 469.8000 1192.5000 471.0000 1199.7001 ;
	    RECT 472.2000 1195.5000 473.4000 1199.7001 ;
	    RECT 474.6000 1195.5000 475.8000 1199.7001 ;
	    RECT 477.0000 1193.7001 478.2000 1199.7001 ;
	    RECT 479.4000 1192.8000 480.6000 1199.7001 ;
	    RECT 481.8000 1193.7001 483.0000 1200.6000 ;
	    RECT 484.2000 1194.6000 485.4000 1199.7001 ;
	    RECT 484.2000 1193.7001 485.7000 1194.6000 ;
	    RECT 486.6000 1193.7001 487.8000 1199.7001 ;
	    RECT 501.0000 1193.7001 502.2000 1199.7001 ;
	    RECT 484.8000 1192.8000 485.7000 1193.7001 ;
	    RECT 477.6000 1191.6000 483.9000 1192.8000 ;
	    RECT 484.8000 1191.9000 487.8000 1192.8000 ;
	    RECT 465.0000 1190.4000 468.9000 1191.6000 ;
	    RECT 469.8000 1190.7001 478.5000 1191.6000 ;
	    RECT 483.0000 1191.0000 483.9000 1191.6000 ;
	    RECT 453.0000 1189.5000 454.2000 1189.8000 ;
	    RECT 285.0000 1188.6000 298.5000 1189.5000 ;
	    RECT 256.2000 1187.4000 257.4000 1188.6000 ;
	    RECT 261.3000 1187.7001 262.5000 1188.0000 ;
	    RECT 258.3000 1186.8000 296.7000 1187.7001 ;
	    RECT 295.5000 1186.5000 296.7000 1186.8000 ;
	    RECT 297.6000 1185.9000 298.5000 1188.6000 ;
	    RECT 299.4000 1188.0000 300.6000 1189.5000 ;
	    RECT 438.6000 1188.0000 439.8000 1189.5000 ;
	    RECT 299.4000 1186.8000 300.9000 1188.0000 ;
	    RECT 253.5000 1185.0000 260.1000 1185.9000 ;
	    RECT 253.5000 1184.7001 254.7000 1185.0000 ;
	    RECT 261.0000 1184.4000 262.2000 1185.6000 ;
	    RECT 263.1000 1185.0000 288.6000 1185.9000 ;
	    RECT 297.6000 1185.0000 298.8000 1185.9000 ;
	    RECT 287.4000 1184.1000 288.6000 1185.0000 ;
	    RECT 78.6000 1182.4501 79.8000 1182.6000 ;
	    RECT 90.6000 1182.4501 91.8000 1182.6000 ;
	    RECT 78.6000 1181.5500 91.8000 1182.4501 ;
	    RECT 78.6000 1181.4000 79.8000 1181.5500 ;
	    RECT 90.6000 1181.4000 91.8000 1181.5500 ;
	    RECT 93.0000 1181.4000 94.2000 1182.6000 ;
	    RECT 114.6000 1181.4000 115.8000 1182.6000 ;
	    RECT 21.0000 1173.3000 22.2000 1179.3000 ;
	    RECT 23.4000 1173.3000 24.6000 1180.2001 ;
	    RECT 47.7000 1179.3000 53.1000 1179.9000 ;
	    RECT 54.6000 1179.3000 55.5000 1180.5000 ;
	    RECT 73.8000 1180.2001 77.1000 1181.1000 ;
	    RECT 47.4000 1179.0000 53.4000 1179.3000 ;
	    RECT 47.4000 1173.3000 48.6000 1179.0000 ;
	    RECT 49.8000 1173.3000 51.0000 1178.1000 ;
	    RECT 52.2000 1173.3000 53.4000 1179.0000 ;
	    RECT 54.6000 1173.3000 55.8000 1179.3000 ;
	    RECT 73.8000 1173.3000 75.0000 1180.2001 ;
	    RECT 76.2000 1173.3000 77.4000 1179.3000 ;
	    RECT 78.6000 1173.3000 79.8000 1180.5000 ;
	    RECT 81.0000 1179.4501 82.2000 1179.6000 ;
	    RECT 90.6000 1179.4501 91.8000 1179.6000 ;
	    RECT 81.0000 1178.5500 91.8000 1179.4501 ;
	    RECT 81.0000 1178.4000 82.2000 1178.5500 ;
	    RECT 90.6000 1178.4000 91.8000 1178.5500 ;
	    RECT 93.0000 1173.3000 94.2000 1180.5000 ;
	    RECT 114.6000 1180.2001 115.8000 1180.5000 ;
	    RECT 95.4000 1179.4501 96.6000 1179.6000 ;
	    RECT 100.2000 1179.4501 101.4000 1179.6000 ;
	    RECT 112.2000 1179.4501 113.4000 1179.6000 ;
	    RECT 95.4000 1178.5500 113.4000 1179.4501 ;
	    RECT 117.0000 1179.3000 118.2000 1183.5000 ;
	    RECT 251.4000 1182.3000 264.6000 1183.5000 ;
	    RECT 265.5000 1182.9000 268.5000 1184.1000 ;
	    RECT 274.2000 1182.9000 279.0000 1184.1000 ;
	    RECT 95.4000 1178.4000 96.6000 1178.5500 ;
	    RECT 100.2000 1178.4000 101.4000 1178.5500 ;
	    RECT 112.2000 1178.4000 113.4000 1178.5500 ;
	    RECT 95.4000 1177.2001 96.6000 1177.5000 ;
	    RECT 95.4000 1173.3000 96.6000 1176.3000 ;
	    RECT 114.6000 1173.3000 115.8000 1179.3000 ;
	    RECT 117.0000 1178.4000 119.7000 1179.3000 ;
	    RECT 118.5000 1173.3000 119.7000 1178.4000 ;
	    RECT 133.8000 1176.4501 135.0000 1176.6000 ;
	    RECT 193.8000 1176.4501 195.0000 1176.6000 ;
	    RECT 133.8000 1175.5500 195.0000 1176.4501 ;
	    RECT 133.8000 1175.4000 135.0000 1175.5500 ;
	    RECT 193.8000 1175.4000 195.0000 1175.5500 ;
	    RECT 251.4000 1173.3000 252.6000 1182.3000 ;
	    RECT 255.0000 1180.2001 259.5000 1181.4000 ;
	    RECT 258.3000 1179.3000 259.5000 1180.2001 ;
	    RECT 267.3000 1179.3000 268.5000 1182.9000 ;
	    RECT 270.6000 1181.4000 271.8000 1182.6000 ;
	    RECT 278.4000 1181.7001 279.6000 1182.0000 ;
	    RECT 273.0000 1180.8000 279.6000 1181.7001 ;
	    RECT 273.0000 1180.5000 274.2000 1180.8000 ;
	    RECT 270.6000 1180.2001 271.8000 1180.5000 ;
	    RECT 282.6000 1179.6000 283.8000 1183.8000 ;
	    RECT 291.3000 1182.9000 297.0000 1184.1000 ;
	    RECT 291.3000 1181.1000 292.5000 1182.9000 ;
	    RECT 297.9000 1182.0000 298.8000 1185.0000 ;
	    RECT 273.0000 1179.3000 274.2000 1179.6000 ;
	    RECT 256.2000 1173.3000 257.4000 1179.3000 ;
	    RECT 258.3000 1178.1000 262.2000 1179.3000 ;
	    RECT 267.3000 1178.4000 274.2000 1179.3000 ;
	    RECT 275.4000 1178.4000 276.6000 1179.6000 ;
	    RECT 277.5000 1178.4000 277.8000 1179.6000 ;
	    RECT 282.3000 1178.4000 283.8000 1179.6000 ;
	    RECT 289.8000 1180.2001 292.5000 1181.1000 ;
	    RECT 297.0000 1181.1000 298.8000 1182.0000 ;
	    RECT 289.8000 1179.3000 291.0000 1180.2001 ;
	    RECT 261.0000 1173.3000 262.2000 1178.1000 ;
	    RECT 287.4000 1178.1000 291.0000 1179.3000 ;
	    RECT 263.4000 1173.3000 264.6000 1177.5000 ;
	    RECT 265.8000 1173.3000 267.0000 1177.5000 ;
	    RECT 268.2000 1173.3000 269.4000 1177.5000 ;
	    RECT 270.6000 1173.3000 271.8000 1176.3000 ;
	    RECT 273.0000 1173.3000 274.2000 1177.5000 ;
	    RECT 275.4000 1173.3000 276.6000 1176.3000 ;
	    RECT 277.8000 1173.3000 279.0000 1177.5000 ;
	    RECT 280.2000 1173.3000 281.4000 1177.5000 ;
	    RECT 282.6000 1173.3000 283.8000 1177.5000 ;
	    RECT 285.0000 1173.3000 286.2000 1177.5000 ;
	    RECT 287.4000 1173.3000 288.6000 1178.1000 ;
	    RECT 292.2000 1173.3000 293.4000 1179.3000 ;
	    RECT 297.0000 1173.3000 298.2000 1181.1000 ;
	    RECT 299.7000 1180.2001 300.9000 1186.8000 ;
	    RECT 438.3000 1186.8000 439.8000 1188.0000 ;
	    RECT 440.7000 1188.6000 454.2000 1189.5000 ;
	    RECT 457.8000 1189.5000 459.0000 1189.8000 ;
	    RECT 469.8000 1189.5000 470.7000 1190.7001 ;
	    RECT 479.4000 1189.8000 481.5000 1190.7001 ;
	    RECT 483.0000 1189.8000 485.4000 1191.0000 ;
	    RECT 457.8000 1188.6000 470.7000 1189.5000 ;
	    RECT 472.2000 1189.5000 481.5000 1189.8000 ;
	    RECT 472.2000 1188.9000 480.3000 1189.5000 ;
	    RECT 472.2000 1188.6000 473.4000 1188.9000 ;
	    RECT 304.2000 1185.4501 305.4000 1185.6000 ;
	    RECT 419.4000 1185.4501 420.6000 1185.6000 ;
	    RECT 304.2000 1184.5500 420.6000 1185.4501 ;
	    RECT 304.2000 1184.4000 305.4000 1184.5500 ;
	    RECT 419.4000 1184.4000 420.6000 1184.5500 ;
	    RECT 299.4000 1179.0000 300.9000 1180.2001 ;
	    RECT 438.3000 1180.2001 439.5000 1186.8000 ;
	    RECT 440.7000 1185.9000 441.6000 1188.6000 ;
	    RECT 476.7000 1187.7001 477.9000 1188.0000 ;
	    RECT 442.5000 1186.8000 480.9000 1187.7001 ;
	    RECT 481.8000 1187.4000 483.0000 1188.6000 ;
	    RECT 442.5000 1186.5000 443.7000 1186.8000 ;
	    RECT 440.4000 1185.0000 441.6000 1185.9000 ;
	    RECT 450.6000 1185.0000 476.1000 1185.9000 ;
	    RECT 440.4000 1182.0000 441.3000 1185.0000 ;
	    RECT 450.6000 1184.1000 451.8000 1185.0000 ;
	    RECT 477.0000 1184.4000 478.2000 1185.6000 ;
	    RECT 479.1000 1185.0000 485.7000 1185.9000 ;
	    RECT 484.5000 1184.7001 485.7000 1185.0000 ;
	    RECT 442.2000 1182.9000 447.9000 1184.1000 ;
	    RECT 440.4000 1181.1000 442.2000 1182.0000 ;
	    RECT 438.3000 1179.0000 439.8000 1180.2001 ;
	    RECT 299.4000 1173.3000 300.6000 1179.0000 ;
	    RECT 301.8000 1173.3000 303.0000 1176.3000 ;
	    RECT 436.2000 1173.3000 437.4000 1176.3000 ;
	    RECT 438.6000 1173.3000 439.8000 1179.0000 ;
	    RECT 441.0000 1173.3000 442.2000 1181.1000 ;
	    RECT 446.7000 1181.1000 447.9000 1182.9000 ;
	    RECT 446.7000 1180.2001 449.4000 1181.1000 ;
	    RECT 448.2000 1179.3000 449.4000 1180.2001 ;
	    RECT 455.4000 1179.6000 456.6000 1183.8000 ;
	    RECT 460.2000 1182.9000 465.0000 1184.1000 ;
	    RECT 470.7000 1182.9000 473.7000 1184.1000 ;
	    RECT 486.6000 1183.5000 487.8000 1191.9000 ;
	    RECT 503.4000 1183.5000 504.6000 1199.7001 ;
	    RECT 522.6000 1193.7001 523.8000 1199.7001 ;
	    RECT 522.6000 1189.5000 523.8000 1189.8000 ;
	    RECT 522.6000 1187.4000 523.8000 1188.6000 ;
	    RECT 525.0000 1186.5000 526.2000 1199.7001 ;
	    RECT 527.4000 1193.7001 528.6000 1199.7001 ;
	    RECT 546.6000 1187.7001 547.8000 1199.7001 ;
	    RECT 550.5000 1188.9000 551.7000 1199.7001 ;
	    RECT 549.0000 1187.7001 551.7000 1188.9000 ;
	    RECT 525.0000 1185.4501 526.2000 1185.6000 ;
	    RECT 544.2000 1185.4501 545.4000 1185.6000 ;
	    RECT 525.0000 1184.5500 545.4000 1185.4501 ;
	    RECT 525.0000 1184.4000 526.2000 1184.5500 ;
	    RECT 544.2000 1184.4000 545.4000 1184.5500 ;
	    RECT 549.3000 1183.5000 550.2000 1187.7001 ;
	    RECT 551.4000 1186.5000 552.6000 1186.8000 ;
	    RECT 551.4000 1184.4000 552.6000 1185.6000 ;
	    RECT 565.8000 1183.5000 567.0000 1199.7001 ;
	    RECT 568.2000 1193.7001 569.4000 1199.7001 ;
	    RECT 601.9500 1197.4501 602.8500 1200.6000 ;
	    RECT 604.2000 1197.4501 605.4000 1197.6000 ;
	    RECT 601.9500 1196.5500 605.4000 1197.4501 ;
	    RECT 604.2000 1196.4000 605.4000 1196.5500 ;
	    RECT 609.0000 1197.4501 610.2000 1197.6000 ;
	    RECT 659.4000 1197.4501 660.6000 1197.6000 ;
	    RECT 609.0000 1196.5500 660.6000 1197.4501 ;
	    RECT 609.0000 1196.4000 610.2000 1196.5500 ;
	    RECT 659.4000 1196.4000 660.6000 1196.5500 ;
	    RECT 700.2000 1193.7001 701.4000 1199.7001 ;
	    RECT 702.6000 1194.6000 703.8000 1199.7001 ;
	    RECT 702.3000 1193.7001 703.8000 1194.6000 ;
	    RECT 705.0000 1193.7001 706.2000 1200.6000 ;
	    RECT 702.3000 1192.8000 703.2000 1193.7001 ;
	    RECT 707.4000 1192.8000 708.6000 1199.7001 ;
	    RECT 709.8000 1193.7001 711.0000 1199.7001 ;
	    RECT 712.2000 1195.5000 713.4000 1199.7001 ;
	    RECT 714.6000 1195.5000 715.8000 1199.7001 ;
	    RECT 700.2000 1191.9000 703.2000 1192.8000 ;
	    RECT 700.2000 1183.5000 701.4000 1191.9000 ;
	    RECT 704.1000 1191.6000 710.4000 1192.8000 ;
	    RECT 717.0000 1192.5000 718.2000 1199.7001 ;
	    RECT 719.4000 1193.7001 720.6000 1199.7001 ;
	    RECT 721.8000 1192.5000 723.0000 1199.7001 ;
	    RECT 724.2000 1193.7001 725.4000 1199.7001 ;
	    RECT 704.1000 1191.0000 705.0000 1191.6000 ;
	    RECT 702.6000 1189.8000 705.0000 1191.0000 ;
	    RECT 709.5000 1190.7001 718.2000 1191.6000 ;
	    RECT 706.5000 1189.8000 708.6000 1190.7001 ;
	    RECT 706.5000 1189.5000 715.8000 1189.8000 ;
	    RECT 707.7000 1188.9000 715.8000 1189.5000 ;
	    RECT 714.6000 1188.6000 715.8000 1188.9000 ;
	    RECT 717.3000 1189.5000 718.2000 1190.7001 ;
	    RECT 719.1000 1190.4000 723.0000 1191.6000 ;
	    RECT 726.6000 1190.4000 727.8000 1199.7001 ;
	    RECT 729.0000 1195.5000 730.2000 1199.7001 ;
	    RECT 731.4000 1195.5000 732.6000 1199.7001 ;
	    RECT 733.8000 1195.5000 735.0000 1199.7001 ;
	    RECT 736.2000 1193.7001 737.4000 1199.7001 ;
	    RECT 731.4000 1191.6000 737.7000 1192.8000 ;
	    RECT 738.6000 1191.6000 739.8000 1199.7001 ;
	    RECT 741.0000 1193.7001 742.2000 1199.7001 ;
	    RECT 743.4000 1192.8000 744.6000 1199.7001 ;
	    RECT 745.8000 1193.7001 747.0000 1199.7001 ;
	    RECT 743.4000 1191.9000 747.3000 1192.8000 ;
	    RECT 748.2000 1192.5000 749.4000 1199.7001 ;
	    RECT 750.6000 1193.7001 751.8000 1199.7001 ;
	    RECT 775.5000 1193.7001 776.7000 1199.7001 ;
	    RECT 738.6000 1190.4000 742.5000 1191.6000 ;
	    RECT 729.0000 1189.5000 730.2000 1189.8000 ;
	    RECT 717.3000 1188.6000 730.2000 1189.5000 ;
	    RECT 733.8000 1189.5000 735.0000 1189.8000 ;
	    RECT 746.4000 1189.5000 747.3000 1191.9000 ;
	    RECT 748.2000 1190.4000 749.4000 1191.6000 ;
	    RECT 775.8000 1190.4000 777.0000 1191.6000 ;
	    RECT 775.8000 1189.5000 776.7000 1190.4000 ;
	    RECT 733.8000 1188.6000 747.3000 1189.5000 ;
	    RECT 705.0000 1187.4000 706.2000 1188.6000 ;
	    RECT 710.1000 1187.7001 711.3000 1188.0000 ;
	    RECT 707.1000 1186.8000 745.5000 1187.7001 ;
	    RECT 744.3000 1186.5000 745.5000 1186.8000 ;
	    RECT 746.4000 1185.9000 747.3000 1188.6000 ;
	    RECT 748.2000 1188.0000 749.4000 1189.5000 ;
	    RECT 777.9000 1188.6000 779.1000 1199.7001 ;
	    RECT 748.2000 1186.8000 749.7000 1188.0000 ;
	    RECT 774.6000 1187.4000 775.8000 1188.6000 ;
	    RECT 777.6000 1187.7001 779.1000 1188.6000 ;
	    RECT 781.8000 1187.7001 783.0000 1199.7001 ;
	    RECT 702.3000 1185.0000 708.9000 1185.9000 ;
	    RECT 702.3000 1184.7001 703.5000 1185.0000 ;
	    RECT 709.8000 1184.4000 711.0000 1185.6000 ;
	    RECT 711.9000 1185.0000 737.4000 1185.9000 ;
	    RECT 746.4000 1185.0000 747.6000 1185.9000 ;
	    RECT 736.2000 1184.1000 737.4000 1185.0000 ;
	    RECT 459.6000 1181.7001 460.8000 1182.0000 ;
	    RECT 459.6000 1180.8000 466.2000 1181.7001 ;
	    RECT 467.4000 1181.4000 468.6000 1182.6000 ;
	    RECT 465.0000 1180.5000 466.2000 1180.8000 ;
	    RECT 467.4000 1180.2001 468.6000 1180.5000 ;
	    RECT 445.8000 1173.3000 447.0000 1179.3000 ;
	    RECT 448.2000 1178.1000 451.8000 1179.3000 ;
	    RECT 455.4000 1178.4000 456.9000 1179.6000 ;
	    RECT 461.4000 1178.4000 461.7000 1179.6000 ;
	    RECT 462.6000 1178.4000 463.8000 1179.6000 ;
	    RECT 465.0000 1179.3000 466.2000 1179.6000 ;
	    RECT 470.7000 1179.3000 471.9000 1182.9000 ;
	    RECT 474.6000 1182.3000 487.8000 1183.5000 ;
	    RECT 479.7000 1180.2001 484.2000 1181.4000 ;
	    RECT 479.7000 1179.3000 480.9000 1180.2001 ;
	    RECT 465.0000 1178.4000 471.9000 1179.3000 ;
	    RECT 450.6000 1173.3000 451.8000 1178.1000 ;
	    RECT 477.0000 1178.1000 480.9000 1179.3000 ;
	    RECT 453.0000 1173.3000 454.2000 1177.5000 ;
	    RECT 455.4000 1173.3000 456.6000 1177.5000 ;
	    RECT 457.8000 1173.3000 459.0000 1177.5000 ;
	    RECT 460.2000 1173.3000 461.4000 1177.5000 ;
	    RECT 462.6000 1173.3000 463.8000 1176.3000 ;
	    RECT 465.0000 1173.3000 466.2000 1177.5000 ;
	    RECT 467.4000 1173.3000 468.6000 1176.3000 ;
	    RECT 469.8000 1173.3000 471.0000 1177.5000 ;
	    RECT 472.2000 1173.3000 473.4000 1177.5000 ;
	    RECT 474.6000 1173.3000 475.8000 1177.5000 ;
	    RECT 477.0000 1173.3000 478.2000 1178.1000 ;
	    RECT 481.8000 1173.3000 483.0000 1179.3000 ;
	    RECT 486.6000 1173.3000 487.8000 1182.3000 ;
	    RECT 503.4000 1182.4501 504.6000 1182.6000 ;
	    RECT 522.6000 1182.4501 523.8000 1182.6000 ;
	    RECT 503.4000 1181.5500 523.8000 1182.4501 ;
	    RECT 503.4000 1181.4000 504.6000 1181.5500 ;
	    RECT 522.6000 1181.4000 523.8000 1181.5500 ;
	    RECT 501.0000 1178.4000 502.2000 1179.6000 ;
	    RECT 501.0000 1177.2001 502.2000 1177.5000 ;
	    RECT 501.0000 1173.3000 502.2000 1176.3000 ;
	    RECT 503.4000 1173.3000 504.6000 1180.5000 ;
	    RECT 525.0000 1179.3000 526.2000 1183.5000 ;
	    RECT 527.4000 1181.4000 528.6000 1182.6000 ;
	    RECT 529.8000 1182.4501 531.0000 1182.6000 ;
	    RECT 549.0000 1182.4501 550.2000 1182.6000 ;
	    RECT 563.4000 1182.4501 564.6000 1182.6000 ;
	    RECT 529.8000 1181.5500 564.6000 1182.4501 ;
	    RECT 529.8000 1181.4000 531.0000 1181.5500 ;
	    RECT 549.0000 1181.4000 550.2000 1181.5500 ;
	    RECT 563.4000 1181.4000 564.6000 1181.5500 ;
	    RECT 565.8000 1182.4501 567.0000 1182.6000 ;
	    RECT 601.8000 1182.4501 603.0000 1182.6000 ;
	    RECT 565.8000 1181.5500 603.0000 1182.4501 ;
	    RECT 565.8000 1181.4000 567.0000 1181.5500 ;
	    RECT 601.8000 1181.4000 603.0000 1181.5500 ;
	    RECT 700.2000 1182.3000 713.4000 1183.5000 ;
	    RECT 714.3000 1182.9000 717.3000 1184.1000 ;
	    RECT 723.0000 1182.9000 727.8000 1184.1000 ;
	    RECT 527.4000 1180.2001 528.6000 1180.5000 ;
	    RECT 523.5000 1178.4000 526.2000 1179.3000 ;
	    RECT 523.5000 1173.3000 524.7000 1178.4000 ;
	    RECT 527.4000 1173.3000 528.6000 1179.3000 ;
	    RECT 546.6000 1178.4000 547.8000 1179.6000 ;
	    RECT 546.6000 1177.2001 547.8000 1177.5000 ;
	    RECT 549.3000 1176.3000 550.2000 1180.5000 ;
	    RECT 546.6000 1173.3000 547.8000 1176.3000 ;
	    RECT 549.0000 1173.3000 550.2000 1176.3000 ;
	    RECT 551.4000 1173.3000 552.6000 1176.3000 ;
	    RECT 565.8000 1173.3000 567.0000 1180.5000 ;
	    RECT 568.2000 1179.4501 569.4000 1179.6000 ;
	    RECT 613.8000 1179.4501 615.0000 1179.6000 ;
	    RECT 633.0000 1179.4501 634.2000 1179.6000 ;
	    RECT 568.2000 1178.5500 634.2000 1179.4501 ;
	    RECT 568.2000 1178.4000 569.4000 1178.5500 ;
	    RECT 613.8000 1178.4000 615.0000 1178.5500 ;
	    RECT 633.0000 1178.4000 634.2000 1178.5500 ;
	    RECT 568.2000 1177.2001 569.4000 1177.5000 ;
	    RECT 568.2000 1173.3000 569.4000 1176.3000 ;
	    RECT 700.2000 1173.3000 701.4000 1182.3000 ;
	    RECT 703.8000 1180.2001 708.3000 1181.4000 ;
	    RECT 707.1000 1179.3000 708.3000 1180.2001 ;
	    RECT 716.1000 1179.3000 717.3000 1182.9000 ;
	    RECT 719.4000 1181.4000 720.6000 1182.6000 ;
	    RECT 727.2000 1181.7001 728.4000 1182.0000 ;
	    RECT 721.8000 1180.8000 728.4000 1181.7001 ;
	    RECT 721.8000 1180.5000 723.0000 1180.8000 ;
	    RECT 719.4000 1180.2001 720.6000 1180.5000 ;
	    RECT 731.4000 1179.6000 732.6000 1183.8000 ;
	    RECT 740.1000 1182.9000 745.8000 1184.1000 ;
	    RECT 740.1000 1181.1000 741.3000 1182.9000 ;
	    RECT 746.7000 1182.0000 747.6000 1185.0000 ;
	    RECT 721.8000 1179.3000 723.0000 1179.6000 ;
	    RECT 705.0000 1173.3000 706.2000 1179.3000 ;
	    RECT 707.1000 1178.1000 711.0000 1179.3000 ;
	    RECT 716.1000 1178.4000 723.0000 1179.3000 ;
	    RECT 724.2000 1178.4000 725.4000 1179.6000 ;
	    RECT 726.3000 1178.4000 726.6000 1179.6000 ;
	    RECT 731.1000 1178.4000 732.6000 1179.6000 ;
	    RECT 738.6000 1180.2001 741.3000 1181.1000 ;
	    RECT 745.8000 1181.1000 747.6000 1182.0000 ;
	    RECT 738.6000 1179.3000 739.8000 1180.2001 ;
	    RECT 709.8000 1173.3000 711.0000 1178.1000 ;
	    RECT 736.2000 1178.1000 739.8000 1179.3000 ;
	    RECT 712.2000 1173.3000 713.4000 1177.5000 ;
	    RECT 714.6000 1173.3000 715.8000 1177.5000 ;
	    RECT 717.0000 1173.3000 718.2000 1177.5000 ;
	    RECT 719.4000 1173.3000 720.6000 1176.3000 ;
	    RECT 721.8000 1173.3000 723.0000 1177.5000 ;
	    RECT 724.2000 1173.3000 725.4000 1176.3000 ;
	    RECT 726.6000 1173.3000 727.8000 1177.5000 ;
	    RECT 729.0000 1173.3000 730.2000 1177.5000 ;
	    RECT 731.4000 1173.3000 732.6000 1177.5000 ;
	    RECT 733.8000 1173.3000 735.0000 1177.5000 ;
	    RECT 736.2000 1173.3000 737.4000 1178.1000 ;
	    RECT 741.0000 1173.3000 742.2000 1179.3000 ;
	    RECT 745.8000 1173.3000 747.0000 1181.1000 ;
	    RECT 748.5000 1180.2001 749.7000 1186.8000 ;
	    RECT 777.6000 1182.6000 778.5000 1187.7001 ;
	    RECT 779.4000 1185.4501 780.6000 1185.6000 ;
	    RECT 779.4000 1184.5500 785.2500 1185.4501 ;
	    RECT 779.4000 1184.4000 780.6000 1184.5500 ;
	    RECT 779.4000 1183.2001 780.6000 1183.5000 ;
	    RECT 772.2000 1182.4501 773.4000 1182.6000 ;
	    RECT 774.6000 1182.4501 775.8000 1182.6000 ;
	    RECT 772.2000 1181.5500 775.8000 1182.4501 ;
	    RECT 772.2000 1181.4000 773.4000 1181.5500 ;
	    RECT 774.6000 1181.4000 775.8000 1181.5500 ;
	    RECT 776.7000 1181.4000 778.5000 1182.6000 ;
	    RECT 780.6000 1180.8000 780.9000 1182.3000 ;
	    RECT 781.8000 1181.4000 783.0000 1182.6000 ;
	    RECT 784.3500 1182.4501 785.2500 1184.5500 ;
	    RECT 796.2000 1183.5000 797.4000 1199.7001 ;
	    RECT 798.6000 1193.7001 799.8000 1199.7001 ;
	    RECT 813.0000 1183.5000 814.2000 1199.7001 ;
	    RECT 815.4000 1193.7001 816.6000 1199.7001 ;
	    RECT 834.6000 1193.7001 835.8000 1199.7001 ;
	    RECT 837.0000 1186.5000 838.2000 1199.7001 ;
	    RECT 839.4000 1193.7001 840.6000 1199.7001 ;
	    RECT 863.4000 1199.4000 864.6000 1200.6000 ;
	    RECT 839.4000 1189.5000 840.6000 1189.8000 ;
	    RECT 839.4000 1187.4000 840.6000 1188.6000 ;
	    RECT 865.8000 1187.7001 867.0000 1199.7001 ;
	    RECT 869.7000 1188.6000 870.9000 1199.7001 ;
	    RECT 872.1000 1193.7001 873.3000 1199.7001 ;
	    RECT 892.2000 1193.7001 893.4000 1199.7001 ;
	    RECT 871.8000 1190.4000 873.0000 1191.6000 ;
	    RECT 872.1000 1189.5000 873.0000 1190.4000 ;
	    RECT 892.2000 1189.5000 893.4000 1189.8000 ;
	    RECT 869.7000 1187.7001 871.2000 1188.6000 ;
	    RECT 837.0000 1185.4501 838.2000 1185.6000 ;
	    RECT 844.2000 1185.4501 845.4000 1185.6000 ;
	    RECT 837.0000 1184.5500 845.4000 1185.4501 ;
	    RECT 837.0000 1184.4000 838.2000 1184.5500 ;
	    RECT 844.2000 1184.4000 845.4000 1184.5500 ;
	    RECT 846.6000 1185.4501 847.8000 1185.6000 ;
	    RECT 868.2000 1185.4501 869.4000 1185.6000 ;
	    RECT 846.6000 1184.5500 869.4000 1185.4501 ;
	    RECT 846.6000 1184.4000 847.8000 1184.5500 ;
	    RECT 868.2000 1184.4000 869.4000 1184.5500 ;
	    RECT 796.2000 1182.4501 797.4000 1182.6000 ;
	    RECT 784.3500 1181.5500 797.4000 1182.4501 ;
	    RECT 796.2000 1181.4000 797.4000 1181.5500 ;
	    RECT 805.8000 1182.4501 807.0000 1182.6000 ;
	    RECT 813.0000 1182.4501 814.2000 1182.6000 ;
	    RECT 805.8000 1181.5500 814.2000 1182.4501 ;
	    RECT 805.8000 1181.4000 807.0000 1181.5500 ;
	    RECT 813.0000 1181.4000 814.2000 1181.5500 ;
	    RECT 832.2000 1182.4501 833.4000 1182.6000 ;
	    RECT 834.6000 1182.4501 835.8000 1182.6000 ;
	    RECT 832.2000 1181.5500 835.8000 1182.4501 ;
	    RECT 832.2000 1181.4000 833.4000 1181.5500 ;
	    RECT 834.6000 1181.4000 835.8000 1181.5500 ;
	    RECT 748.2000 1179.0000 749.7000 1180.2001 ;
	    RECT 774.9000 1179.3000 775.8000 1180.5000 ;
	    RECT 777.3000 1179.3000 782.7000 1179.9000 ;
	    RECT 748.2000 1173.3000 749.4000 1179.0000 ;
	    RECT 750.6000 1173.3000 751.8000 1176.3000 ;
	    RECT 774.6000 1173.3000 775.8000 1179.3000 ;
	    RECT 777.0000 1179.0000 783.0000 1179.3000 ;
	    RECT 777.0000 1173.3000 778.2000 1179.0000 ;
	    RECT 779.4000 1173.3000 780.6000 1178.1000 ;
	    RECT 781.8000 1173.3000 783.0000 1179.0000 ;
	    RECT 796.2000 1173.3000 797.4000 1180.5000 ;
	    RECT 798.6000 1179.4501 799.8000 1179.6000 ;
	    RECT 808.2000 1179.4501 809.4000 1179.6000 ;
	    RECT 798.6000 1178.5500 809.4000 1179.4501 ;
	    RECT 798.6000 1178.4000 799.8000 1178.5500 ;
	    RECT 808.2000 1178.4000 809.4000 1178.5500 ;
	    RECT 798.6000 1177.2001 799.8000 1177.5000 ;
	    RECT 798.6000 1173.3000 799.8000 1176.3000 ;
	    RECT 813.0000 1173.3000 814.2000 1180.5000 ;
	    RECT 834.6000 1180.2001 835.8000 1180.5000 ;
	    RECT 815.4000 1179.4501 816.6000 1179.6000 ;
	    RECT 827.4000 1179.4501 828.6000 1179.6000 ;
	    RECT 815.4000 1178.5500 828.6000 1179.4501 ;
	    RECT 837.0000 1179.3000 838.2000 1183.5000 ;
	    RECT 868.2000 1183.2001 869.4000 1183.5000 ;
	    RECT 870.3000 1182.6000 871.2000 1187.7001 ;
	    RECT 873.0000 1187.4000 874.2000 1188.6000 ;
	    RECT 892.2000 1187.4000 893.4000 1188.6000 ;
	    RECT 894.6000 1186.5000 895.8000 1199.7001 ;
	    RECT 897.0000 1193.7001 898.2000 1199.7001 ;
	    RECT 904.2000 1199.4000 905.4000 1200.6000 ;
	    RECT 924.3000 1188.9000 925.5000 1199.7001 ;
	    RECT 924.3000 1187.7001 927.0000 1188.9000 ;
	    RECT 928.2000 1187.7001 929.4000 1199.7001 ;
	    RECT 959.4000 1187.7001 960.6000 1199.7001 ;
	    RECT 963.3000 1187.7001 966.3000 1199.7001 ;
	    RECT 969.0000 1187.7001 970.2000 1199.7001 ;
	    RECT 923.4000 1186.5000 924.6000 1186.8000 ;
	    RECT 882.6000 1185.4501 883.8000 1185.6000 ;
	    RECT 894.6000 1185.4501 895.8000 1185.6000 ;
	    RECT 904.2000 1185.4501 905.4000 1185.6000 ;
	    RECT 882.6000 1184.5500 895.8000 1185.4501 ;
	    RECT 882.6000 1184.4000 883.8000 1184.5500 ;
	    RECT 894.6000 1184.4000 895.8000 1184.5500 ;
	    RECT 897.1500 1184.5500 905.4000 1185.4501 ;
	    RECT 863.4000 1182.4501 864.6000 1182.6000 ;
	    RECT 865.8000 1182.4501 867.0000 1182.6000 ;
	    RECT 863.4000 1181.5500 867.0000 1182.4501 ;
	    RECT 863.4000 1181.4000 864.6000 1181.5500 ;
	    RECT 865.8000 1181.4000 867.0000 1181.5500 ;
	    RECT 867.9000 1180.8000 868.2000 1182.3000 ;
	    RECT 870.3000 1181.4000 872.1000 1182.6000 ;
	    RECT 873.0000 1182.4501 874.2000 1182.6000 ;
	    RECT 889.8000 1182.4501 891.0000 1182.6000 ;
	    RECT 873.0000 1181.5500 891.0000 1182.4501 ;
	    RECT 873.0000 1181.4000 874.2000 1181.5500 ;
	    RECT 889.8000 1181.4000 891.0000 1181.5500 ;
	    RECT 866.1000 1179.3000 871.5000 1179.9000 ;
	    RECT 873.0000 1179.3000 873.9000 1180.5000 ;
	    RECT 894.6000 1179.3000 895.8000 1183.5000 ;
	    RECT 897.1500 1182.6000 898.0500 1184.5500 ;
	    RECT 904.2000 1184.4000 905.4000 1184.5500 ;
	    RECT 923.4000 1184.4000 924.6000 1185.6000 ;
	    RECT 925.8000 1183.5000 926.7000 1187.7001 ;
	    RECT 961.8000 1184.4000 963.0000 1185.6000 ;
	    RECT 959.4000 1183.5000 960.6000 1183.8000 ;
	    RECT 964.5000 1183.5000 965.4000 1187.7001 ;
	    RECT 966.6000 1184.4000 967.8000 1185.6000 ;
	    RECT 981.0000 1183.5000 982.2000 1199.7001 ;
	    RECT 983.4000 1193.7001 984.6000 1199.7001 ;
	    RECT 995.4000 1183.5000 996.6000 1199.7001 ;
	    RECT 997.8000 1193.7001 999.0000 1199.7001 ;
	    RECT 1009.8000 1193.7001 1011.0000 1199.7001 ;
	    RECT 1012.2000 1183.5000 1013.4000 1199.7001 ;
	    RECT 1043.4000 1188.4501 1044.6000 1188.6000 ;
	    RECT 1079.4000 1188.4501 1080.6000 1188.6000 ;
	    RECT 1043.4000 1187.5500 1080.6000 1188.4501 ;
	    RECT 1043.4000 1187.4000 1044.6000 1187.5500 ;
	    RECT 1079.4000 1187.4000 1080.6000 1187.5500 ;
	    RECT 1081.8000 1187.1000 1083.0000 1199.7001 ;
	    RECT 1084.2001 1188.0000 1085.4000 1199.7001 ;
	    RECT 1088.4000 1194.6000 1089.6000 1199.7001 ;
	    RECT 1086.6000 1193.7001 1089.6000 1194.6000 ;
	    RECT 1092.6000 1193.7001 1093.8000 1199.7001 ;
	    RECT 1095.0000 1193.7001 1096.2001 1199.7001 ;
	    RECT 1097.4000 1193.7001 1098.6000 1199.7001 ;
	    RECT 1101.3000 1193.7001 1103.1000 1199.7001 ;
	    RECT 1086.6000 1192.5000 1087.8000 1193.7001 ;
	    RECT 1095.0000 1192.8000 1095.9000 1193.7001 ;
	    RECT 1091.7001 1191.9000 1097.1000 1192.8000 ;
	    RECT 1101.0000 1192.5000 1102.2001 1193.7001 ;
	    RECT 1091.7001 1191.6000 1092.9000 1191.9000 ;
	    RECT 1095.9000 1191.6000 1097.1000 1191.9000 ;
	    RECT 1086.6000 1189.5000 1087.8000 1189.8000 ;
	    RECT 1093.5000 1189.5000 1094.7001 1189.8000 ;
	    RECT 1086.6000 1188.6000 1094.7001 1189.5000 ;
	    RECT 1095.6000 1189.5000 1098.9000 1190.4000 ;
	    RECT 1095.6000 1187.7001 1096.5000 1189.5000 ;
	    RECT 1097.7001 1189.2001 1098.9000 1189.5000 ;
	    RECT 1101.3000 1189.8000 1103.4000 1191.0000 ;
	    RECT 1101.3000 1188.3000 1102.2001 1189.8000 ;
	    RECT 1089.3000 1187.1000 1096.5000 1187.7001 ;
	    RECT 1081.8000 1186.8000 1096.5000 1187.1000 ;
	    RECT 1098.6000 1187.4000 1102.2001 1188.3000 ;
	    RECT 1105.8000 1187.7001 1107.0000 1199.7001 ;
	    RECT 1081.8000 1186.5000 1090.5000 1186.8000 ;
	    RECT 1081.8000 1186.2001 1090.2001 1186.5000 ;
	    RECT 1091.4000 1185.4501 1092.6000 1185.6000 ;
	    RECT 1093.8000 1185.4501 1095.0000 1185.6000 ;
	    RECT 1085.1000 1184.4000 1090.5000 1185.3000 ;
	    RECT 1091.4000 1184.5500 1095.0000 1185.4501 ;
	    RECT 1091.4000 1184.4000 1092.6000 1184.5500 ;
	    RECT 1093.8000 1184.4000 1095.0000 1184.5500 ;
	    RECT 1085.1000 1184.1000 1086.3000 1184.4000 ;
	    RECT 961.8000 1183.2001 963.0000 1183.5000 ;
	    RECT 966.6000 1183.2001 967.8000 1183.5000 ;
	    RECT 1087.5000 1182.6000 1088.7001 1182.9000 ;
	    RECT 1098.6000 1182.6000 1099.5000 1187.4000 ;
	    RECT 1108.2001 1186.8000 1109.4000 1199.7001 ;
	    RECT 1110.6000 1199.4000 1111.8000 1200.6000 ;
	    RECT 1134.6000 1193.7001 1135.8000 1199.7001 ;
	    RECT 1103.1000 1186.5000 1109.4000 1186.8000 ;
	    RECT 1137.0000 1186.5000 1138.2001 1199.7001 ;
	    RECT 1139.4000 1193.7001 1140.6000 1199.7001 ;
	    RECT 1264.2001 1193.7001 1265.4000 1199.7001 ;
	    RECT 1266.6000 1192.5000 1267.8000 1199.7001 ;
	    RECT 1269.0000 1193.7001 1270.2001 1199.7001 ;
	    RECT 1271.4000 1192.8000 1272.6000 1199.7001 ;
	    RECT 1273.8000 1193.7001 1275.0000 1199.7001 ;
	    RECT 1268.7001 1191.9000 1272.6000 1192.8000 ;
	    RECT 1233.0000 1191.4501 1234.2001 1191.6000 ;
	    RECT 1266.6000 1191.4501 1267.8000 1191.6000 ;
	    RECT 1233.0000 1190.5500 1267.8000 1191.4501 ;
	    RECT 1233.0000 1190.4000 1234.2001 1190.5500 ;
	    RECT 1266.6000 1190.4000 1267.8000 1190.5500 ;
	    RECT 1139.4000 1189.5000 1140.6000 1189.8000 ;
	    RECT 1268.7001 1189.5000 1269.6000 1191.9000 ;
	    RECT 1276.2001 1191.6000 1277.4000 1199.7001 ;
	    RECT 1278.6000 1193.7001 1279.8000 1199.7001 ;
	    RECT 1281.0000 1195.5000 1282.2001 1199.7001 ;
	    RECT 1283.4000 1195.5000 1284.6000 1199.7001 ;
	    RECT 1285.8000 1195.5000 1287.0000 1199.7001 ;
	    RECT 1278.3000 1191.6000 1284.6000 1192.8000 ;
	    RECT 1273.5000 1190.4000 1277.4000 1191.6000 ;
	    RECT 1288.2001 1190.4000 1289.4000 1199.7001 ;
	    RECT 1290.6000 1193.7001 1291.8000 1199.7001 ;
	    RECT 1293.0000 1192.5000 1294.2001 1199.7001 ;
	    RECT 1295.4000 1193.7001 1296.6000 1199.7001 ;
	    RECT 1297.8000 1192.5000 1299.0000 1199.7001 ;
	    RECT 1300.2001 1195.5000 1301.4000 1199.7001 ;
	    RECT 1302.6000 1195.5000 1303.8000 1199.7001 ;
	    RECT 1305.0000 1193.7001 1306.2001 1199.7001 ;
	    RECT 1307.4000 1192.8000 1308.6000 1199.7001 ;
	    RECT 1309.8000 1193.7001 1311.0000 1200.6000 ;
	    RECT 1312.2001 1194.6000 1313.4000 1199.7001 ;
	    RECT 1312.2001 1193.7001 1313.7001 1194.6000 ;
	    RECT 1314.6000 1193.7001 1315.8000 1199.7001 ;
	    RECT 1312.8000 1192.8000 1313.7001 1193.7001 ;
	    RECT 1305.6000 1191.6000 1311.9000 1192.8000 ;
	    RECT 1312.8000 1191.9000 1315.8000 1192.8000 ;
	    RECT 1293.0000 1190.4000 1296.9000 1191.6000 ;
	    RECT 1297.8000 1190.7001 1306.5000 1191.6000 ;
	    RECT 1311.0000 1191.0000 1311.9000 1191.6000 ;
	    RECT 1281.0000 1189.5000 1282.2001 1189.8000 ;
	    RECT 1139.4000 1188.4501 1140.6000 1188.6000 ;
	    RECT 1165.8000 1188.4501 1167.0000 1188.6000 ;
	    RECT 1139.4000 1187.5500 1167.0000 1188.4501 ;
	    RECT 1266.6000 1188.0000 1267.8000 1189.5000 ;
	    RECT 1139.4000 1187.4000 1140.6000 1187.5500 ;
	    RECT 1165.8000 1187.4000 1167.0000 1187.5500 ;
	    RECT 1266.3000 1186.8000 1267.8000 1188.0000 ;
	    RECT 1268.7001 1188.6000 1282.2001 1189.5000 ;
	    RECT 1285.8000 1189.5000 1287.0000 1189.8000 ;
	    RECT 1297.8000 1189.5000 1298.7001 1190.7001 ;
	    RECT 1307.4000 1189.8000 1309.5000 1190.7001 ;
	    RECT 1311.0000 1189.8000 1313.4000 1191.0000 ;
	    RECT 1285.8000 1188.6000 1298.7001 1189.5000 ;
	    RECT 1300.2001 1189.5000 1309.5000 1189.8000 ;
	    RECT 1300.2001 1188.9000 1308.3000 1189.5000 ;
	    RECT 1300.2001 1188.6000 1301.4000 1188.9000 ;
	    RECT 1103.1000 1185.9000 1107.3000 1186.5000 ;
	    RECT 1103.1000 1185.6000 1104.3000 1185.9000 ;
	    RECT 1108.2001 1185.4501 1109.4000 1185.6000 ;
	    RECT 1117.8000 1185.4501 1119.0000 1185.6000 ;
	    RECT 1105.5000 1184.7001 1106.7001 1185.0000 ;
	    RECT 1101.0000 1183.8000 1106.7001 1184.7001 ;
	    RECT 1108.2001 1184.5500 1119.0000 1185.4501 ;
	    RECT 1108.2001 1184.4000 1109.4000 1184.5500 ;
	    RECT 1117.8000 1184.4000 1119.0000 1184.5500 ;
	    RECT 1137.0000 1185.4501 1138.2001 1185.6000 ;
	    RECT 1180.2001 1185.4501 1181.4000 1185.6000 ;
	    RECT 1137.0000 1184.5500 1181.4000 1185.4501 ;
	    RECT 1137.0000 1184.4000 1138.2001 1184.5500 ;
	    RECT 1180.2001 1184.4000 1181.4000 1184.5500 ;
	    RECT 1101.0000 1183.5000 1102.2001 1183.8000 ;
	    RECT 897.0000 1181.4000 898.2000 1182.6000 ;
	    RECT 899.4000 1182.4501 900.6000 1182.6000 ;
	    RECT 925.8000 1182.4501 927.0000 1182.6000 ;
	    RECT 899.4000 1181.5500 927.0000 1182.4501 ;
	    RECT 899.4000 1181.4000 900.6000 1181.5500 ;
	    RECT 925.8000 1181.4000 927.0000 1181.5500 ;
	    RECT 959.4000 1181.4000 960.6000 1182.6000 ;
	    RECT 961.8000 1181.4000 963.3000 1182.3000 ;
	    RECT 964.2000 1181.4000 965.4000 1182.6000 ;
	    RECT 969.0000 1182.4501 970.2000 1182.6000 ;
	    RECT 976.2000 1182.4501 977.4000 1182.6000 ;
	    RECT 897.0000 1180.2001 898.2000 1180.5000 ;
	    RECT 815.4000 1178.4000 816.6000 1178.5500 ;
	    RECT 827.4000 1178.4000 828.6000 1178.5500 ;
	    RECT 815.4000 1177.2001 816.6000 1177.5000 ;
	    RECT 815.4000 1173.3000 816.6000 1176.3000 ;
	    RECT 834.6000 1173.3000 835.8000 1179.3000 ;
	    RECT 837.0000 1178.4000 839.7000 1179.3000 ;
	    RECT 838.5000 1173.3000 839.7000 1178.4000 ;
	    RECT 865.8000 1179.0000 871.8000 1179.3000 ;
	    RECT 865.8000 1173.3000 867.0000 1179.0000 ;
	    RECT 868.2000 1173.3000 869.4000 1178.1000 ;
	    RECT 870.6000 1173.3000 871.8000 1179.0000 ;
	    RECT 873.0000 1173.3000 874.2000 1179.3000 ;
	    RECT 893.1000 1178.4000 895.8000 1179.3000 ;
	    RECT 893.1000 1173.3000 894.3000 1178.4000 ;
	    RECT 897.0000 1173.3000 898.2000 1179.3000 ;
	    RECT 899.4000 1176.4501 900.6000 1176.6000 ;
	    RECT 916.2000 1176.4501 917.4000 1176.6000 ;
	    RECT 899.4000 1175.5500 917.4000 1176.4501 ;
	    RECT 925.8000 1176.3000 926.7000 1180.5000 ;
	    RECT 928.2000 1179.4501 929.4000 1179.6000 ;
	    RECT 933.0000 1179.4501 934.2000 1179.6000 ;
	    RECT 928.2000 1178.5500 934.2000 1179.4501 ;
	    RECT 961.8000 1179.3000 962.7000 1181.4000 ;
	    RECT 967.8000 1180.8000 968.1000 1182.3000 ;
	    RECT 969.0000 1181.5500 977.4000 1182.4501 ;
	    RECT 969.0000 1181.4000 970.2000 1181.5500 ;
	    RECT 976.2000 1181.4000 977.4000 1181.5500 ;
	    RECT 981.0000 1181.4000 982.2000 1182.6000 ;
	    RECT 983.4000 1182.4501 984.6000 1182.6000 ;
	    RECT 995.4000 1182.4501 996.6000 1182.6000 ;
	    RECT 983.4000 1181.5500 996.6000 1182.4501 ;
	    RECT 983.4000 1181.4000 984.6000 1181.5500 ;
	    RECT 995.4000 1181.4000 996.6000 1181.5500 ;
	    RECT 1012.2000 1182.4501 1013.4000 1182.6000 ;
	    RECT 1021.8000 1182.4501 1023.0000 1182.6000 ;
	    RECT 1012.2000 1181.5500 1023.0000 1182.4501 ;
	    RECT 1012.2000 1181.4000 1013.4000 1181.5500 ;
	    RECT 1021.8000 1181.4000 1023.0000 1181.5500 ;
	    RECT 1083.0000 1181.4000 1083.3000 1182.6000 ;
	    RECT 1084.2001 1181.4000 1085.4000 1182.6000 ;
	    RECT 1086.3000 1181.7001 1099.5000 1182.6000 ;
	    RECT 964.5000 1179.3000 969.9000 1179.9000 ;
	    RECT 928.2000 1178.4000 929.4000 1178.5500 ;
	    RECT 933.0000 1178.4000 934.2000 1178.5500 ;
	    RECT 928.2000 1177.2001 929.4000 1177.5000 ;
	    RECT 899.4000 1175.4000 900.6000 1175.5500 ;
	    RECT 916.2000 1175.4000 917.4000 1175.5500 ;
	    RECT 923.4000 1173.3000 924.6000 1176.3000 ;
	    RECT 925.8000 1173.3000 927.0000 1176.3000 ;
	    RECT 928.2000 1173.3000 929.4000 1176.3000 ;
	    RECT 959.4000 1174.2001 960.6000 1179.3000 ;
	    RECT 961.8000 1175.1000 963.0000 1179.3000 ;
	    RECT 964.2000 1179.0000 970.2000 1179.3000 ;
	    RECT 964.2000 1174.2001 965.4000 1179.0000 ;
	    RECT 959.4000 1173.3000 965.4000 1174.2001 ;
	    RECT 966.6000 1173.3000 967.8000 1178.1000 ;
	    RECT 969.0000 1173.3000 970.2000 1179.0000 ;
	    RECT 981.0000 1173.3000 982.2000 1180.5000 ;
	    RECT 983.4000 1178.4000 984.6000 1179.6000 ;
	    RECT 983.4000 1177.2001 984.6000 1177.5000 ;
	    RECT 983.4000 1173.3000 984.6000 1176.3000 ;
	    RECT 995.4000 1173.3000 996.6000 1180.5000 ;
	    RECT 997.8000 1178.4000 999.0000 1179.6000 ;
	    RECT 1000.2000 1179.4501 1001.4000 1179.6000 ;
	    RECT 1009.8000 1179.4501 1011.0000 1179.6000 ;
	    RECT 1000.2000 1178.5500 1011.0000 1179.4501 ;
	    RECT 1000.2000 1178.4000 1001.4000 1178.5500 ;
	    RECT 1009.8000 1178.4000 1011.0000 1178.5500 ;
	    RECT 997.8000 1177.2001 999.0000 1177.5000 ;
	    RECT 1009.8000 1177.2001 1011.0000 1177.5000 ;
	    RECT 997.8000 1173.3000 999.0000 1176.3000 ;
	    RECT 1009.8000 1173.3000 1011.0000 1176.3000 ;
	    RECT 1012.2000 1173.3000 1013.4000 1180.5000 ;
	    RECT 1081.8000 1173.3000 1083.0000 1180.5000 ;
	    RECT 1084.2001 1173.3000 1085.4000 1179.3000 ;
	    RECT 1089.3000 1178.4000 1090.2001 1181.7001 ;
	    RECT 1097.7001 1181.4000 1098.9000 1181.7001 ;
	    RECT 1108.2001 1180.8000 1109.4000 1183.5000 ;
	    RECT 1110.6000 1182.4501 1111.8000 1182.6000 ;
	    RECT 1134.6000 1182.4501 1135.8000 1182.6000 ;
	    RECT 1110.6000 1181.5500 1135.8000 1182.4501 ;
	    RECT 1110.6000 1181.4000 1111.8000 1181.5500 ;
	    RECT 1134.6000 1181.4000 1135.8000 1181.5500 ;
	    RECT 1103.7001 1179.9000 1109.4000 1180.8000 ;
	    RECT 1134.6000 1180.2001 1135.8000 1180.5000 ;
	    RECT 1103.7001 1179.6000 1104.9000 1179.9000 ;
	    RECT 1086.6000 1176.3000 1087.8000 1177.5000 ;
	    RECT 1089.0000 1177.2001 1090.2001 1178.4000 ;
	    RECT 1091.7001 1178.1000 1092.9000 1178.4000 ;
	    RECT 1091.7001 1177.2001 1095.9000 1178.1000 ;
	    RECT 1095.0000 1176.3000 1095.9000 1177.2001 ;
	    RECT 1101.0000 1176.3000 1102.2001 1177.5000 ;
	    RECT 1086.6000 1175.4000 1089.6000 1176.3000 ;
	    RECT 1088.4000 1173.3000 1089.6000 1175.4000 ;
	    RECT 1092.3000 1173.3000 1093.8000 1176.3000 ;
	    RECT 1095.0000 1173.3000 1096.2001 1176.3000 ;
	    RECT 1097.4000 1173.3000 1098.6000 1176.3000 ;
	    RECT 1101.0000 1175.4000 1103.1000 1176.3000 ;
	    RECT 1101.3000 1173.3000 1103.1000 1175.4000 ;
	    RECT 1105.8000 1173.3000 1107.0000 1179.0000 ;
	    RECT 1108.2001 1173.3000 1109.4000 1179.9000 ;
	    RECT 1137.0000 1179.3000 1138.2001 1183.5000 ;
	    RECT 1266.3000 1180.2001 1267.5000 1186.8000 ;
	    RECT 1268.7001 1185.9000 1269.6000 1188.6000 ;
	    RECT 1304.7001 1187.7001 1305.9000 1188.0000 ;
	    RECT 1270.5000 1186.8000 1308.9000 1187.7001 ;
	    RECT 1309.8000 1187.4000 1311.0000 1188.6000 ;
	    RECT 1270.5000 1186.5000 1271.7001 1186.8000 ;
	    RECT 1268.4000 1185.0000 1269.6000 1185.9000 ;
	    RECT 1278.6000 1185.0000 1304.1000 1185.9000 ;
	    RECT 1268.4000 1182.0000 1269.3000 1185.0000 ;
	    RECT 1278.6000 1184.1000 1279.8000 1185.0000 ;
	    RECT 1305.0000 1184.4000 1306.2001 1185.6000 ;
	    RECT 1307.1000 1185.0000 1313.7001 1185.9000 ;
	    RECT 1312.5000 1184.7001 1313.7001 1185.0000 ;
	    RECT 1270.2001 1182.9000 1275.9000 1184.1000 ;
	    RECT 1268.4000 1181.1000 1270.2001 1182.0000 ;
	    RECT 1134.6000 1173.3000 1135.8000 1179.3000 ;
	    RECT 1137.0000 1178.4000 1139.7001 1179.3000 ;
	    RECT 1266.3000 1179.0000 1267.8000 1180.2001 ;
	    RECT 1138.5000 1173.3000 1139.7001 1178.4000 ;
	    RECT 1264.2001 1173.3000 1265.4000 1176.3000 ;
	    RECT 1266.6000 1173.3000 1267.8000 1179.0000 ;
	    RECT 1269.0000 1173.3000 1270.2001 1181.1000 ;
	    RECT 1274.7001 1181.1000 1275.9000 1182.9000 ;
	    RECT 1274.7001 1180.2001 1277.4000 1181.1000 ;
	    RECT 1276.2001 1179.3000 1277.4000 1180.2001 ;
	    RECT 1283.4000 1179.6000 1284.6000 1183.8000 ;
	    RECT 1288.2001 1182.9000 1293.0000 1184.1000 ;
	    RECT 1298.7001 1182.9000 1301.7001 1184.1000 ;
	    RECT 1314.6000 1183.5000 1315.8000 1191.9000 ;
	    RECT 1341.0000 1187.7001 1342.2001 1199.7001 ;
	    RECT 1344.9000 1188.6000 1346.1000 1199.7001 ;
	    RECT 1347.3000 1193.7001 1348.5000 1199.7001 ;
	    RECT 1482.6000 1193.7001 1483.8000 1199.7001 ;
	    RECT 1485.0000 1192.5000 1486.2001 1199.7001 ;
	    RECT 1487.4000 1193.7001 1488.6000 1199.7001 ;
	    RECT 1489.8000 1192.8000 1491.0000 1199.7001 ;
	    RECT 1492.2001 1193.7001 1493.4000 1199.7001 ;
	    RECT 1487.1000 1191.9000 1491.0000 1192.8000 ;
	    RECT 1347.0000 1190.4000 1348.2001 1191.6000 ;
	    RECT 1429.8000 1191.4501 1431.0000 1191.6000 ;
	    RECT 1485.0000 1191.4501 1486.2001 1191.6000 ;
	    RECT 1429.8000 1190.5500 1486.2001 1191.4501 ;
	    RECT 1429.8000 1190.4000 1431.0000 1190.5500 ;
	    RECT 1485.0000 1190.4000 1486.2001 1190.5500 ;
	    RECT 1347.3000 1189.5000 1348.2001 1190.4000 ;
	    RECT 1487.1000 1189.5000 1488.0000 1191.9000 ;
	    RECT 1494.6000 1191.6000 1495.8000 1199.7001 ;
	    RECT 1497.0000 1193.7001 1498.2001 1199.7001 ;
	    RECT 1499.4000 1195.5000 1500.6000 1199.7001 ;
	    RECT 1501.8000 1195.5000 1503.0000 1199.7001 ;
	    RECT 1504.2001 1195.5000 1505.4000 1199.7001 ;
	    RECT 1496.7001 1191.6000 1503.0000 1192.8000 ;
	    RECT 1491.9000 1190.4000 1495.8000 1191.6000 ;
	    RECT 1506.6000 1190.4000 1507.8000 1199.7001 ;
	    RECT 1509.0000 1193.7001 1510.2001 1199.7001 ;
	    RECT 1511.4000 1192.5000 1512.6000 1199.7001 ;
	    RECT 1513.8000 1193.7001 1515.0000 1199.7001 ;
	    RECT 1516.2001 1192.5000 1517.4000 1199.7001 ;
	    RECT 1518.6000 1195.5000 1519.8000 1199.7001 ;
	    RECT 1521.0000 1195.5000 1522.2001 1199.7001 ;
	    RECT 1523.4000 1193.7001 1524.6000 1199.7001 ;
	    RECT 1525.8000 1192.8000 1527.0000 1199.7001 ;
	    RECT 1528.2001 1193.7001 1529.4000 1200.6000 ;
	    RECT 1530.6000 1194.6000 1531.8000 1199.7001 ;
	    RECT 1530.6000 1193.7001 1532.1000 1194.6000 ;
	    RECT 1533.0000 1193.7001 1534.2001 1199.7001 ;
	    RECT 1540.2001 1199.4000 1541.4000 1200.6000 ;
	    RECT 1531.2001 1192.8000 1532.1000 1193.7001 ;
	    RECT 1524.0000 1191.6000 1530.3000 1192.8000 ;
	    RECT 1531.2001 1191.9000 1534.2001 1192.8000 ;
	    RECT 1511.4000 1190.4000 1515.3000 1191.6000 ;
	    RECT 1516.2001 1190.7001 1524.9000 1191.6000 ;
	    RECT 1529.4000 1191.0000 1530.3000 1191.6000 ;
	    RECT 1499.4000 1189.5000 1500.6000 1189.8000 ;
	    RECT 1344.9000 1187.7001 1346.4000 1188.6000 ;
	    RECT 1343.4000 1184.4000 1344.6000 1185.6000 ;
	    RECT 1287.6000 1181.7001 1288.8000 1182.0000 ;
	    RECT 1287.6000 1180.8000 1294.2001 1181.7001 ;
	    RECT 1295.4000 1181.4000 1296.6000 1182.6000 ;
	    RECT 1293.0000 1180.5000 1294.2001 1180.8000 ;
	    RECT 1295.4000 1180.2001 1296.6000 1180.5000 ;
	    RECT 1273.8000 1173.3000 1275.0000 1179.3000 ;
	    RECT 1276.2001 1178.1000 1279.8000 1179.3000 ;
	    RECT 1283.4000 1178.4000 1284.9000 1179.6000 ;
	    RECT 1289.4000 1178.4000 1289.7001 1179.6000 ;
	    RECT 1290.6000 1178.4000 1291.8000 1179.6000 ;
	    RECT 1293.0000 1179.3000 1294.2001 1179.6000 ;
	    RECT 1298.7001 1179.3000 1299.9000 1182.9000 ;
	    RECT 1302.6000 1182.3000 1315.8000 1183.5000 ;
	    RECT 1343.4000 1183.2001 1344.6000 1183.5000 ;
	    RECT 1345.5000 1182.6000 1346.4000 1187.7001 ;
	    RECT 1348.2001 1188.4501 1349.4000 1188.6000 ;
	    RECT 1393.8000 1188.4501 1395.0000 1188.6000 ;
	    RECT 1348.2001 1187.5500 1395.0000 1188.4501 ;
	    RECT 1485.0000 1188.0000 1486.2001 1189.5000 ;
	    RECT 1348.2001 1187.4000 1349.4000 1187.5500 ;
	    RECT 1393.8000 1187.4000 1395.0000 1187.5500 ;
	    RECT 1484.7001 1186.8000 1486.2001 1188.0000 ;
	    RECT 1487.1000 1188.6000 1500.6000 1189.5000 ;
	    RECT 1504.2001 1189.5000 1505.4000 1189.8000 ;
	    RECT 1516.2001 1189.5000 1517.1000 1190.7001 ;
	    RECT 1525.8000 1189.8000 1527.9000 1190.7001 ;
	    RECT 1529.4000 1189.8000 1531.8000 1191.0000 ;
	    RECT 1504.2001 1188.6000 1517.1000 1189.5000 ;
	    RECT 1518.6000 1189.5000 1527.9000 1189.8000 ;
	    RECT 1518.6000 1188.9000 1526.7001 1189.5000 ;
	    RECT 1518.6000 1188.6000 1519.8000 1188.9000 ;
	    RECT 1307.7001 1180.2001 1312.2001 1181.4000 ;
	    RECT 1307.7001 1179.3000 1308.9000 1180.2001 ;
	    RECT 1293.0000 1178.4000 1299.9000 1179.3000 ;
	    RECT 1278.6000 1173.3000 1279.8000 1178.1000 ;
	    RECT 1305.0000 1178.1000 1308.9000 1179.3000 ;
	    RECT 1281.0000 1173.3000 1282.2001 1177.5000 ;
	    RECT 1283.4000 1173.3000 1284.6000 1177.5000 ;
	    RECT 1285.8000 1173.3000 1287.0000 1177.5000 ;
	    RECT 1288.2001 1173.3000 1289.4000 1177.5000 ;
	    RECT 1290.6000 1173.3000 1291.8000 1176.3000 ;
	    RECT 1293.0000 1173.3000 1294.2001 1177.5000 ;
	    RECT 1295.4000 1173.3000 1296.6000 1176.3000 ;
	    RECT 1297.8000 1173.3000 1299.0000 1177.5000 ;
	    RECT 1300.2001 1173.3000 1301.4000 1177.5000 ;
	    RECT 1302.6000 1173.3000 1303.8000 1177.5000 ;
	    RECT 1305.0000 1173.3000 1306.2001 1178.1000 ;
	    RECT 1309.8000 1173.3000 1311.0000 1179.3000 ;
	    RECT 1314.6000 1173.3000 1315.8000 1182.3000 ;
	    RECT 1317.0000 1182.4501 1318.2001 1182.6000 ;
	    RECT 1341.0000 1182.4501 1342.2001 1182.6000 ;
	    RECT 1317.0000 1181.5500 1342.2001 1182.4501 ;
	    RECT 1317.0000 1181.4000 1318.2001 1181.5500 ;
	    RECT 1341.0000 1181.4000 1342.2001 1181.5500 ;
	    RECT 1343.1000 1180.8000 1343.4000 1182.3000 ;
	    RECT 1345.5000 1181.4000 1347.3000 1182.6000 ;
	    RECT 1348.2001 1181.4000 1349.4000 1182.6000 ;
	    RECT 1341.3000 1179.3000 1346.7001 1179.9000 ;
	    RECT 1348.2001 1179.3000 1349.1000 1180.5000 ;
	    RECT 1484.7001 1180.2001 1485.9000 1186.8000 ;
	    RECT 1487.1000 1185.9000 1488.0000 1188.6000 ;
	    RECT 1528.2001 1188.4501 1529.4000 1188.6000 ;
	    RECT 1530.6000 1188.4501 1531.8000 1188.6000 ;
	    RECT 1523.1000 1187.7001 1524.3000 1188.0000 ;
	    RECT 1488.9000 1186.8000 1527.3000 1187.7001 ;
	    RECT 1528.2001 1187.5500 1531.8000 1188.4501 ;
	    RECT 1528.2001 1187.4000 1529.4000 1187.5500 ;
	    RECT 1530.6000 1187.4000 1531.8000 1187.5500 ;
	    RECT 1488.9000 1186.5000 1490.1000 1186.8000 ;
	    RECT 1486.8000 1185.0000 1488.0000 1185.9000 ;
	    RECT 1497.0000 1185.0000 1522.5000 1185.9000 ;
	    RECT 1486.8000 1182.0000 1487.7001 1185.0000 ;
	    RECT 1497.0000 1184.1000 1498.2001 1185.0000 ;
	    RECT 1523.4000 1184.4000 1524.6000 1185.6000 ;
	    RECT 1525.5000 1185.0000 1532.1000 1185.9000 ;
	    RECT 1530.9000 1184.7001 1532.1000 1185.0000 ;
	    RECT 1488.6000 1182.9000 1494.3000 1184.1000 ;
	    RECT 1486.8000 1181.1000 1488.6000 1182.0000 ;
	    RECT 1341.0000 1179.0000 1347.0000 1179.3000 ;
	    RECT 1341.0000 1173.3000 1342.2001 1179.0000 ;
	    RECT 1343.4000 1173.3000 1344.6000 1178.1000 ;
	    RECT 1345.8000 1173.3000 1347.0000 1179.0000 ;
	    RECT 1348.2001 1173.3000 1349.4000 1179.3000 ;
	    RECT 1484.7001 1179.0000 1486.2001 1180.2001 ;
	    RECT 1482.6000 1173.3000 1483.8000 1176.3000 ;
	    RECT 1485.0000 1173.3000 1486.2001 1179.0000 ;
	    RECT 1487.4000 1173.3000 1488.6000 1181.1000 ;
	    RECT 1493.1000 1181.1000 1494.3000 1182.9000 ;
	    RECT 1493.1000 1180.2001 1495.8000 1181.1000 ;
	    RECT 1494.6000 1179.3000 1495.8000 1180.2001 ;
	    RECT 1501.8000 1179.6000 1503.0000 1183.8000 ;
	    RECT 1506.6000 1182.9000 1511.4000 1184.1000 ;
	    RECT 1517.1000 1182.9000 1520.1000 1184.1000 ;
	    RECT 1533.0000 1183.5000 1534.2001 1191.9000 ;
	    RECT 1552.2001 1187.7001 1553.4000 1199.7001 ;
	    RECT 1554.6000 1189.5000 1555.8000 1199.7001 ;
	    RECT 1557.0000 1188.6000 1558.2001 1199.7001 ;
	    RECT 1554.9000 1187.7001 1558.2001 1188.6000 ;
	    RECT 1552.2001 1184.4000 1553.1000 1187.7001 ;
	    RECT 1554.9000 1186.8000 1555.8000 1187.7001 ;
	    RECT 1554.0000 1185.6000 1555.8000 1186.8000 ;
	    RECT 1552.2001 1183.5000 1553.4000 1184.4000 ;
	    RECT 1506.0000 1181.7001 1507.2001 1182.0000 ;
	    RECT 1506.0000 1180.8000 1512.6000 1181.7001 ;
	    RECT 1513.8000 1181.4000 1515.0000 1182.6000 ;
	    RECT 1511.4000 1180.5000 1512.6000 1180.8000 ;
	    RECT 1513.8000 1180.2001 1515.0000 1180.5000 ;
	    RECT 1492.2001 1173.3000 1493.4000 1179.3000 ;
	    RECT 1494.6000 1178.1000 1498.2001 1179.3000 ;
	    RECT 1501.8000 1178.4000 1503.3000 1179.6000 ;
	    RECT 1507.8000 1178.4000 1508.1000 1179.6000 ;
	    RECT 1509.0000 1178.4000 1510.2001 1179.6000 ;
	    RECT 1511.4000 1179.3000 1512.6000 1179.6000 ;
	    RECT 1517.1000 1179.3000 1518.3000 1182.9000 ;
	    RECT 1521.0000 1182.3000 1534.2001 1183.5000 ;
	    RECT 1526.1000 1180.2001 1530.6000 1181.4000 ;
	    RECT 1526.1000 1179.3000 1527.3000 1180.2001 ;
	    RECT 1511.4000 1178.4000 1518.3000 1179.3000 ;
	    RECT 1497.0000 1173.3000 1498.2001 1178.1000 ;
	    RECT 1523.4000 1178.1000 1527.3000 1179.3000 ;
	    RECT 1499.4000 1173.3000 1500.6000 1177.5000 ;
	    RECT 1501.8000 1173.3000 1503.0000 1177.5000 ;
	    RECT 1504.2001 1173.3000 1505.4000 1177.5000 ;
	    RECT 1506.6000 1173.3000 1507.8000 1177.5000 ;
	    RECT 1509.0000 1173.3000 1510.2001 1176.3000 ;
	    RECT 1511.4000 1173.3000 1512.6000 1177.5000 ;
	    RECT 1513.8000 1173.3000 1515.0000 1176.3000 ;
	    RECT 1516.2001 1173.3000 1517.4000 1177.5000 ;
	    RECT 1518.6000 1173.3000 1519.8000 1177.5000 ;
	    RECT 1521.0000 1173.3000 1522.2001 1177.5000 ;
	    RECT 1523.4000 1173.3000 1524.6000 1178.1000 ;
	    RECT 1528.2001 1173.3000 1529.4000 1179.3000 ;
	    RECT 1533.0000 1173.3000 1534.2001 1182.3000 ;
	    RECT 1554.9000 1181.1000 1555.8000 1185.6000 ;
	    RECT 1557.0000 1184.4000 1558.2001 1185.6000 ;
	    RECT 1557.0000 1183.2001 1558.2001 1183.5000 ;
	    RECT 1542.6000 1179.4501 1543.8000 1179.6000 ;
	    RECT 1547.4000 1179.4501 1548.6000 1179.6000 ;
	    RECT 1542.6000 1178.5500 1548.6000 1179.4501 ;
	    RECT 1542.6000 1178.4000 1543.8000 1178.5500 ;
	    RECT 1547.4000 1178.4000 1548.6000 1178.5500 ;
	    RECT 1552.2001 1173.3000 1553.4000 1180.5000 ;
	    RECT 1554.9000 1180.2001 1558.2001 1181.1000 ;
	    RECT 1554.6000 1173.3000 1555.8000 1179.3000 ;
	    RECT 1557.0000 1173.3000 1558.2001 1180.2001 ;
	    RECT 1.2000 1170.6000 1569.0000 1172.4000 ;
	    RECT 13.8000 1166.7001 15.0000 1169.7001 ;
	    RECT 13.8000 1165.5000 15.0000 1165.8000 ;
	    RECT 13.8000 1163.4000 15.0000 1164.6000 ;
	    RECT 16.2000 1162.5000 17.4000 1169.7001 ;
	    RECT 141.0000 1166.7001 142.2000 1169.7001 ;
	    RECT 143.4000 1164.0000 144.6000 1169.7001 ;
	    RECT 143.1000 1162.8000 144.6000 1164.0000 ;
	    RECT 16.2000 1161.4501 17.4000 1161.6000 ;
	    RECT 49.8000 1161.4501 51.0000 1161.6000 ;
	    RECT 16.2000 1160.5500 51.0000 1161.4501 ;
	    RECT 16.2000 1160.4000 17.4000 1160.5500 ;
	    RECT 49.8000 1160.4000 51.0000 1160.5500 ;
	    RECT 13.8000 1143.3000 15.0000 1149.3000 ;
	    RECT 16.2000 1143.3000 17.4000 1159.5000 ;
	    RECT 143.1000 1156.2001 144.3000 1162.8000 ;
	    RECT 145.8000 1161.9000 147.0000 1169.7001 ;
	    RECT 150.6000 1163.7001 151.8000 1169.7001 ;
	    RECT 155.4000 1164.9000 156.6000 1169.7001 ;
	    RECT 157.8000 1165.5000 159.0000 1169.7001 ;
	    RECT 160.2000 1165.5000 161.4000 1169.7001 ;
	    RECT 162.6000 1165.5000 163.8000 1169.7001 ;
	    RECT 165.0000 1165.5000 166.2000 1169.7001 ;
	    RECT 167.4000 1166.7001 168.6000 1169.7001 ;
	    RECT 169.8000 1165.5000 171.0000 1169.7001 ;
	    RECT 172.2000 1166.7001 173.4000 1169.7001 ;
	    RECT 174.6000 1165.5000 175.8000 1169.7001 ;
	    RECT 177.0000 1165.5000 178.2000 1169.7001 ;
	    RECT 179.4000 1165.5000 180.6000 1169.7001 ;
	    RECT 153.0000 1163.7001 156.6000 1164.9000 ;
	    RECT 181.8000 1164.9000 183.0000 1169.7001 ;
	    RECT 153.0000 1162.8000 154.2000 1163.7001 ;
	    RECT 145.2000 1161.0000 147.0000 1161.9000 ;
	    RECT 151.5000 1161.9000 154.2000 1162.8000 ;
	    RECT 160.2000 1163.4000 161.7000 1164.6000 ;
	    RECT 166.2000 1163.4000 166.5000 1164.6000 ;
	    RECT 167.4000 1163.4000 168.6000 1164.6000 ;
	    RECT 169.8000 1163.7001 176.7000 1164.6000 ;
	    RECT 181.8000 1163.7001 185.7000 1164.9000 ;
	    RECT 186.6000 1163.7001 187.8000 1169.7001 ;
	    RECT 169.8000 1163.4000 171.0000 1163.7001 ;
	    RECT 145.2000 1158.0000 146.1000 1161.0000 ;
	    RECT 151.5000 1160.1000 152.7000 1161.9000 ;
	    RECT 147.0000 1158.9000 152.7000 1160.1000 ;
	    RECT 160.2000 1159.2001 161.4000 1163.4000 ;
	    RECT 172.2000 1162.5000 173.4000 1162.8000 ;
	    RECT 169.8000 1162.2001 171.0000 1162.5000 ;
	    RECT 164.4000 1161.3000 171.0000 1162.2001 ;
	    RECT 164.4000 1161.0000 165.6000 1161.3000 ;
	    RECT 172.2000 1160.4000 173.4000 1161.6000 ;
	    RECT 175.5000 1160.1000 176.7000 1163.7001 ;
	    RECT 184.5000 1162.8000 185.7000 1163.7001 ;
	    RECT 184.5000 1161.6000 189.0000 1162.8000 ;
	    RECT 191.4000 1160.7001 192.6000 1169.7001 ;
	    RECT 218.7000 1164.6000 219.9000 1169.7001 ;
	    RECT 218.7000 1163.7001 221.4000 1164.6000 ;
	    RECT 222.6000 1163.7001 223.8000 1169.7001 ;
	    RECT 246.6000 1163.7001 247.8000 1169.7001 ;
	    RECT 249.0000 1164.0000 250.2000 1169.7001 ;
	    RECT 251.4000 1164.9000 252.6000 1169.7001 ;
	    RECT 253.8000 1164.0000 255.0000 1169.7001 ;
	    RECT 249.0000 1163.7001 255.0000 1164.0000 ;
	    RECT 165.0000 1158.9000 169.8000 1160.1000 ;
	    RECT 175.5000 1158.9000 178.5000 1160.1000 ;
	    RECT 179.4000 1159.5000 192.6000 1160.7001 ;
	    RECT 220.2000 1159.5000 221.4000 1163.7001 ;
	    RECT 222.6000 1162.5000 223.8000 1162.8000 ;
	    RECT 246.9000 1162.5000 247.8000 1163.7001 ;
	    RECT 249.3000 1163.1000 254.7000 1163.7001 ;
	    RECT 268.2000 1162.5000 269.4000 1169.7001 ;
	    RECT 270.6000 1166.7001 271.8000 1169.7001 ;
	    RECT 275.4000 1167.4501 276.6000 1167.6000 ;
	    RECT 289.8000 1167.4501 291.0000 1167.6000 ;
	    RECT 275.4000 1166.5500 291.0000 1167.4501 ;
	    RECT 275.4000 1166.4000 276.6000 1166.5500 ;
	    RECT 289.8000 1166.4000 291.0000 1166.5500 ;
	    RECT 270.6000 1165.5000 271.8000 1165.8000 ;
	    RECT 270.6000 1164.4501 271.8000 1164.6000 ;
	    RECT 299.4000 1164.4501 300.6000 1164.6000 ;
	    RECT 270.6000 1163.5500 300.6000 1164.4501 ;
	    RECT 301.8000 1164.0000 303.0000 1169.7001 ;
	    RECT 304.2000 1164.9000 305.4000 1169.7001 ;
	    RECT 306.6000 1168.8000 312.6000 1169.7001 ;
	    RECT 306.6000 1164.0000 307.8000 1168.8000 ;
	    RECT 301.8000 1163.7001 307.8000 1164.0000 ;
	    RECT 309.0000 1163.7001 310.2000 1167.9000 ;
	    RECT 311.4000 1163.7001 312.6000 1168.8000 ;
	    RECT 323.4000 1166.7001 324.6000 1169.7001 ;
	    RECT 323.4000 1165.5000 324.6000 1165.8000 ;
	    RECT 270.6000 1163.4000 271.8000 1163.5500 ;
	    RECT 299.4000 1163.4000 300.6000 1163.5500 ;
	    RECT 302.1000 1163.1000 307.5000 1163.7001 ;
	    RECT 222.6000 1160.4000 223.8000 1161.6000 ;
	    RECT 246.6000 1160.4000 247.8000 1161.6000 ;
	    RECT 248.7000 1160.4000 250.5000 1161.6000 ;
	    RECT 252.6000 1160.7001 252.9000 1162.2001 ;
	    RECT 253.8000 1160.4000 255.0000 1161.6000 ;
	    RECT 268.2000 1161.4501 269.4000 1161.6000 ;
	    RECT 256.3500 1160.5500 269.4000 1161.4501 ;
	    RECT 155.4000 1158.0000 156.6000 1158.9000 ;
	    RECT 145.2000 1157.1000 146.4000 1158.0000 ;
	    RECT 155.4000 1157.1000 180.9000 1158.0000 ;
	    RECT 181.8000 1157.4000 183.0000 1158.6000 ;
	    RECT 189.3000 1158.0000 190.5000 1158.3000 ;
	    RECT 183.9000 1157.1000 190.5000 1158.0000 ;
	    RECT 143.1000 1155.0000 144.6000 1156.2001 ;
	    RECT 143.4000 1153.5000 144.6000 1155.0000 ;
	    RECT 145.5000 1154.4000 146.4000 1157.1000 ;
	    RECT 147.3000 1156.2001 148.5000 1156.5000 ;
	    RECT 147.3000 1155.3000 185.7000 1156.2001 ;
	    RECT 181.5000 1155.0000 182.7000 1155.3000 ;
	    RECT 186.6000 1154.4000 187.8000 1155.6000 ;
	    RECT 145.5000 1153.5000 159.0000 1154.4000 ;
	    RECT 114.6000 1152.4501 115.8000 1152.6000 ;
	    RECT 143.4000 1152.4501 144.6000 1152.6000 ;
	    RECT 114.6000 1151.5500 144.6000 1152.4501 ;
	    RECT 114.6000 1151.4000 115.8000 1151.5500 ;
	    RECT 143.4000 1151.4000 144.6000 1151.5500 ;
	    RECT 145.5000 1151.1000 146.4000 1153.5000 ;
	    RECT 157.8000 1153.2001 159.0000 1153.5000 ;
	    RECT 162.6000 1153.5000 175.5000 1154.4000 ;
	    RECT 162.6000 1153.2001 163.8000 1153.5000 ;
	    RECT 150.3000 1151.4000 154.2000 1152.6000 ;
	    RECT 141.0000 1143.3000 142.2000 1149.3000 ;
	    RECT 143.4000 1143.3000 144.6000 1150.5000 ;
	    RECT 145.5000 1150.2001 149.4000 1151.1000 ;
	    RECT 145.8000 1143.3000 147.0000 1149.3000 ;
	    RECT 148.2000 1143.3000 149.4000 1150.2001 ;
	    RECT 150.6000 1143.3000 151.8000 1149.3000 ;
	    RECT 153.0000 1143.3000 154.2000 1151.4000 ;
	    RECT 155.1000 1150.2001 161.4000 1151.4000 ;
	    RECT 155.4000 1143.3000 156.6000 1149.3000 ;
	    RECT 157.8000 1143.3000 159.0000 1147.5000 ;
	    RECT 160.2000 1143.3000 161.4000 1147.5000 ;
	    RECT 162.6000 1143.3000 163.8000 1147.5000 ;
	    RECT 165.0000 1143.3000 166.2000 1152.6000 ;
	    RECT 169.8000 1151.4000 173.7000 1152.6000 ;
	    RECT 174.6000 1152.3000 175.5000 1153.5000 ;
	    RECT 177.0000 1154.1000 178.2000 1154.4000 ;
	    RECT 177.0000 1153.5000 185.1000 1154.1000 ;
	    RECT 177.0000 1153.2001 186.3000 1153.5000 ;
	    RECT 184.2000 1152.3000 186.3000 1153.2001 ;
	    RECT 174.6000 1151.4000 183.3000 1152.3000 ;
	    RECT 187.8000 1152.0000 190.2000 1153.2001 ;
	    RECT 187.8000 1151.4000 188.7000 1152.0000 ;
	    RECT 167.4000 1143.3000 168.6000 1149.3000 ;
	    RECT 169.8000 1143.3000 171.0000 1150.5000 ;
	    RECT 172.2000 1143.3000 173.4000 1149.3000 ;
	    RECT 174.6000 1143.3000 175.8000 1150.5000 ;
	    RECT 182.4000 1150.2001 188.7000 1151.4000 ;
	    RECT 191.4000 1151.1000 192.6000 1159.5000 ;
	    RECT 220.2000 1158.4501 221.4000 1158.6000 ;
	    RECT 220.2000 1157.5500 247.6500 1158.4501 ;
	    RECT 220.2000 1157.4000 221.4000 1157.5500 ;
	    RECT 196.2000 1155.4501 197.4000 1155.6000 ;
	    RECT 217.8000 1155.4501 219.0000 1155.6000 ;
	    RECT 196.2000 1154.5500 219.0000 1155.4501 ;
	    RECT 196.2000 1154.4000 197.4000 1154.5500 ;
	    RECT 217.8000 1154.4000 219.0000 1154.5500 ;
	    RECT 217.8000 1153.2001 219.0000 1153.5000 ;
	    RECT 189.6000 1150.2001 192.6000 1151.1000 ;
	    RECT 177.0000 1143.3000 178.2000 1147.5000 ;
	    RECT 179.4000 1143.3000 180.6000 1147.5000 ;
	    RECT 181.8000 1143.3000 183.0000 1149.3000 ;
	    RECT 184.2000 1143.3000 185.4000 1150.2001 ;
	    RECT 189.6000 1149.3000 190.5000 1150.2001 ;
	    RECT 186.6000 1142.4000 187.8000 1149.3000 ;
	    RECT 189.0000 1148.4000 190.5000 1149.3000 ;
	    RECT 189.0000 1143.3000 190.2000 1148.4000 ;
	    RECT 191.4000 1143.3000 192.6000 1149.3000 ;
	    RECT 217.8000 1143.3000 219.0000 1149.3000 ;
	    RECT 220.2000 1143.3000 221.4000 1156.5000 ;
	    RECT 246.7500 1155.6000 247.6500 1157.5500 ;
	    RECT 246.6000 1154.4000 247.8000 1155.6000 ;
	    RECT 249.6000 1155.3000 250.5000 1160.4000 ;
	    RECT 251.4000 1159.5000 252.6000 1159.8000 ;
	    RECT 251.4000 1158.4501 252.6000 1158.6000 ;
	    RECT 256.3500 1158.4501 257.2500 1160.5500 ;
	    RECT 268.2000 1160.4000 269.4000 1160.5500 ;
	    RECT 297.0000 1161.4501 298.2000 1161.6000 ;
	    RECT 301.8000 1161.4501 303.0000 1161.6000 ;
	    RECT 297.0000 1160.5500 303.0000 1161.4501 ;
	    RECT 303.9000 1160.7001 304.2000 1162.2001 ;
	    RECT 309.3000 1161.6000 310.2000 1163.7001 ;
	    RECT 323.4000 1163.4000 324.6000 1164.6000 ;
	    RECT 325.8000 1162.5000 327.0000 1169.7001 ;
	    RECT 460.2000 1166.7001 461.4000 1169.7001 ;
	    RECT 462.6000 1164.0000 463.8000 1169.7001 ;
	    RECT 462.3000 1162.8000 463.8000 1164.0000 ;
	    RECT 297.0000 1160.4000 298.2000 1160.5500 ;
	    RECT 301.8000 1160.4000 303.0000 1160.5500 ;
	    RECT 306.6000 1160.4000 307.8000 1161.6000 ;
	    RECT 308.7000 1160.7001 310.2000 1161.6000 ;
	    RECT 311.4000 1161.4501 312.6000 1161.6000 ;
	    RECT 313.8000 1161.4501 315.0000 1161.6000 ;
	    RECT 311.4000 1160.5500 315.0000 1161.4501 ;
	    RECT 311.4000 1160.4000 312.6000 1160.5500 ;
	    RECT 313.8000 1160.4000 315.0000 1160.5500 ;
	    RECT 325.8000 1161.4501 327.0000 1161.6000 ;
	    RECT 364.2000 1161.4501 365.4000 1161.6000 ;
	    RECT 325.8000 1160.5500 365.4000 1161.4501 ;
	    RECT 325.8000 1160.4000 327.0000 1160.5500 ;
	    RECT 364.2000 1160.4000 365.4000 1160.5500 ;
	    RECT 304.2000 1159.5000 305.4000 1159.8000 ;
	    RECT 309.0000 1159.5000 310.2000 1159.8000 ;
	    RECT 251.4000 1157.5500 257.2500 1158.4501 ;
	    RECT 251.4000 1157.4000 252.6000 1157.5500 ;
	    RECT 249.6000 1154.4000 251.1000 1155.3000 ;
	    RECT 247.8000 1152.6000 248.7000 1153.5000 ;
	    RECT 247.8000 1151.4000 249.0000 1152.6000 ;
	    RECT 222.6000 1143.3000 223.8000 1149.3000 ;
	    RECT 247.5000 1143.3000 248.7000 1149.3000 ;
	    RECT 249.9000 1143.3000 251.1000 1154.4000 ;
	    RECT 253.8000 1143.3000 255.0000 1155.3000 ;
	    RECT 256.2000 1146.4501 257.4000 1146.6000 ;
	    RECT 263.4000 1146.4501 264.6000 1146.6000 ;
	    RECT 256.2000 1145.5500 264.6000 1146.4501 ;
	    RECT 256.2000 1145.4000 257.4000 1145.5500 ;
	    RECT 263.4000 1145.4000 264.6000 1145.5500 ;
	    RECT 268.2000 1143.3000 269.4000 1159.5000 ;
	    RECT 275.4000 1158.4501 276.6000 1158.6000 ;
	    RECT 287.4000 1158.4501 288.6000 1158.6000 ;
	    RECT 304.2000 1158.4501 305.4000 1158.6000 ;
	    RECT 275.4000 1157.5500 305.4000 1158.4501 ;
	    RECT 275.4000 1157.4000 276.6000 1157.5500 ;
	    RECT 287.4000 1157.4000 288.6000 1157.5500 ;
	    RECT 304.2000 1157.4000 305.4000 1157.5500 ;
	    RECT 306.6000 1155.3000 307.5000 1159.5000 ;
	    RECT 311.4000 1159.2001 312.6000 1159.5000 ;
	    RECT 309.0000 1157.4000 310.2000 1158.6000 ;
	    RECT 270.6000 1143.3000 271.8000 1149.3000 ;
	    RECT 301.8000 1143.3000 303.0000 1155.3000 ;
	    RECT 305.7000 1143.3000 308.7000 1155.3000 ;
	    RECT 311.4000 1143.3000 312.6000 1155.3000 ;
	    RECT 323.4000 1143.3000 324.6000 1149.3000 ;
	    RECT 325.8000 1143.3000 327.0000 1159.5000 ;
	    RECT 462.3000 1156.2001 463.5000 1162.8000 ;
	    RECT 465.0000 1161.9000 466.2000 1169.7001 ;
	    RECT 469.8000 1163.7001 471.0000 1169.7001 ;
	    RECT 474.6000 1164.9000 475.8000 1169.7001 ;
	    RECT 477.0000 1165.5000 478.2000 1169.7001 ;
	    RECT 479.4000 1165.5000 480.6000 1169.7001 ;
	    RECT 481.8000 1165.5000 483.0000 1169.7001 ;
	    RECT 484.2000 1165.5000 485.4000 1169.7001 ;
	    RECT 486.6000 1166.7001 487.8000 1169.7001 ;
	    RECT 489.0000 1165.5000 490.2000 1169.7001 ;
	    RECT 491.4000 1166.7001 492.6000 1169.7001 ;
	    RECT 493.8000 1165.5000 495.0000 1169.7001 ;
	    RECT 496.2000 1165.5000 497.4000 1169.7001 ;
	    RECT 498.6000 1165.5000 499.8000 1169.7001 ;
	    RECT 472.2000 1163.7001 475.8000 1164.9000 ;
	    RECT 501.0000 1164.9000 502.2000 1169.7001 ;
	    RECT 472.2000 1162.8000 473.4000 1163.7001 ;
	    RECT 464.4000 1161.0000 466.2000 1161.9000 ;
	    RECT 470.7000 1161.9000 473.4000 1162.8000 ;
	    RECT 479.4000 1163.4000 480.9000 1164.6000 ;
	    RECT 485.4000 1163.4000 485.7000 1164.6000 ;
	    RECT 486.6000 1163.4000 487.8000 1164.6000 ;
	    RECT 489.0000 1163.7001 495.9000 1164.6000 ;
	    RECT 501.0000 1163.7001 504.9000 1164.9000 ;
	    RECT 505.8000 1163.7001 507.0000 1169.7001 ;
	    RECT 489.0000 1163.4000 490.2000 1163.7001 ;
	    RECT 464.4000 1158.0000 465.3000 1161.0000 ;
	    RECT 470.7000 1160.1000 471.9000 1161.9000 ;
	    RECT 466.2000 1158.9000 471.9000 1160.1000 ;
	    RECT 479.4000 1159.2001 480.6000 1163.4000 ;
	    RECT 491.4000 1162.5000 492.6000 1162.8000 ;
	    RECT 489.0000 1162.2001 490.2000 1162.5000 ;
	    RECT 483.6000 1161.3000 490.2000 1162.2001 ;
	    RECT 483.6000 1161.0000 484.8000 1161.3000 ;
	    RECT 491.4000 1160.4000 492.6000 1161.6000 ;
	    RECT 494.7000 1160.1000 495.9000 1163.7001 ;
	    RECT 503.7000 1162.8000 504.9000 1163.7001 ;
	    RECT 503.7000 1161.6000 508.2000 1162.8000 ;
	    RECT 510.6000 1160.7001 511.8000 1169.7001 ;
	    RECT 551.4000 1163.7001 552.6000 1169.7001 ;
	    RECT 553.8000 1164.6000 555.3000 1169.7001 ;
	    RECT 558.0000 1164.3000 560.4000 1169.7001 ;
	    RECT 563.1000 1164.6000 564.6000 1169.7001 ;
	    RECT 551.4000 1162.8000 555.3000 1163.7001 ;
	    RECT 554.1000 1162.5000 555.3000 1162.8000 ;
	    RECT 556.2000 1162.2001 558.6000 1163.4000 ;
	    RECT 484.2000 1158.9000 489.0000 1160.1000 ;
	    RECT 494.7000 1158.9000 497.7000 1160.1000 ;
	    RECT 498.6000 1159.5000 511.8000 1160.7001 ;
	    RECT 544.2000 1161.4501 545.4000 1161.6000 ;
	    RECT 551.4000 1161.4501 552.6000 1161.6000 ;
	    RECT 544.2000 1160.5500 552.6000 1161.4501 ;
	    RECT 544.2000 1160.4000 545.4000 1160.5500 ;
	    RECT 551.4000 1160.4000 552.6000 1160.5500 ;
	    RECT 553.5000 1161.3000 553.8000 1161.6000 ;
	    RECT 559.5000 1161.3000 560.4000 1164.3000 ;
	    RECT 565.8000 1163.7001 567.0000 1169.7001 ;
	    RECT 585.0000 1163.7001 586.2000 1169.7001 ;
	    RECT 588.9000 1164.6000 590.1000 1169.7001 ;
	    RECT 587.4000 1163.7001 590.1000 1164.6000 ;
	    RECT 616.2000 1164.0000 617.4000 1169.7001 ;
	    RECT 618.6000 1164.9000 619.8000 1169.7001 ;
	    RECT 621.0000 1164.0000 622.2000 1169.7001 ;
	    RECT 616.2000 1163.7001 622.2000 1164.0000 ;
	    RECT 623.4000 1163.7001 624.6000 1169.7001 ;
	    RECT 561.3000 1162.2001 562.5000 1163.4000 ;
	    RECT 563.4000 1162.8000 567.0000 1163.7001 ;
	    RECT 563.4000 1162.5000 564.6000 1162.8000 ;
	    RECT 585.0000 1162.5000 586.2000 1162.8000 ;
	    RECT 553.5000 1161.0000 554.7000 1161.3000 ;
	    RECT 553.5000 1160.4000 558.0000 1161.0000 ;
	    RECT 553.8000 1160.1000 558.0000 1160.4000 ;
	    RECT 556.8000 1159.8000 558.0000 1160.1000 ;
	    RECT 558.9000 1160.4000 560.4000 1161.3000 ;
	    RECT 561.6000 1161.6000 562.5000 1162.2001 ;
	    RECT 561.6000 1160.4000 562.8000 1161.6000 ;
	    RECT 564.6000 1160.4000 564.9000 1161.6000 ;
	    RECT 565.8000 1160.4000 567.0000 1161.6000 ;
	    RECT 580.2000 1161.4501 581.4000 1161.6000 ;
	    RECT 585.0000 1161.4501 586.2000 1161.6000 ;
	    RECT 580.2000 1160.5500 586.2000 1161.4501 ;
	    RECT 580.2000 1160.4000 581.4000 1160.5500 ;
	    RECT 585.0000 1160.4000 586.2000 1160.5500 ;
	    RECT 558.9000 1159.5000 559.8000 1160.4000 ;
	    RECT 587.4000 1159.5000 588.6000 1163.7001 ;
	    RECT 616.5000 1163.1000 621.9000 1163.7001 ;
	    RECT 623.4000 1162.5000 624.3000 1163.7001 ;
	    RECT 700.2000 1162.5000 701.4000 1169.7001 ;
	    RECT 702.6000 1163.7001 703.8000 1169.7001 ;
	    RECT 706.8000 1167.6000 708.0000 1169.7001 ;
	    RECT 705.0000 1166.7001 708.0000 1167.6000 ;
	    RECT 710.7000 1166.7001 712.2000 1169.7001 ;
	    RECT 713.4000 1166.7001 714.6000 1169.7001 ;
	    RECT 715.8000 1166.7001 717.0000 1169.7001 ;
	    RECT 719.7000 1167.6000 721.5000 1169.7001 ;
	    RECT 719.4000 1166.7001 721.5000 1167.6000 ;
	    RECT 705.0000 1165.5000 706.2000 1166.7001 ;
	    RECT 713.4000 1165.8000 714.3000 1166.7001 ;
	    RECT 707.4000 1164.6000 708.6000 1165.8000 ;
	    RECT 710.1000 1164.9000 714.3000 1165.8000 ;
	    RECT 719.4000 1165.5000 720.6000 1166.7001 ;
	    RECT 710.1000 1164.6000 711.3000 1164.9000 ;
	    RECT 589.8000 1161.4501 591.0000 1161.6000 ;
	    RECT 613.8000 1161.4501 615.0000 1161.6000 ;
	    RECT 616.2000 1161.4501 617.4000 1161.6000 ;
	    RECT 589.8000 1160.5500 617.4000 1161.4501 ;
	    RECT 618.3000 1160.7001 618.6000 1162.2001 ;
	    RECT 589.8000 1160.4000 591.0000 1160.5500 ;
	    RECT 613.8000 1160.4000 615.0000 1160.5500 ;
	    RECT 616.2000 1160.4000 617.4000 1160.5500 ;
	    RECT 620.7000 1160.4000 622.5000 1161.6000 ;
	    RECT 623.4000 1161.4501 624.6000 1161.6000 ;
	    RECT 628.2000 1161.4501 629.4000 1161.6000 ;
	    RECT 623.4000 1160.5500 629.4000 1161.4501 ;
	    RECT 623.4000 1160.4000 624.6000 1160.5500 ;
	    RECT 628.2000 1160.4000 629.4000 1160.5500 ;
	    RECT 701.4000 1160.4000 701.7000 1161.6000 ;
	    RECT 702.6000 1160.4000 703.8000 1161.6000 ;
	    RECT 707.7000 1161.3000 708.6000 1164.6000 ;
	    RECT 724.2000 1164.0000 725.4000 1169.7001 ;
	    RECT 722.1000 1163.1000 723.3000 1163.4000 ;
	    RECT 726.6000 1163.1000 727.8000 1169.7001 ;
	    RECT 745.8000 1163.7001 747.0000 1169.7001 ;
	    RECT 749.7000 1164.6000 750.9000 1169.7001 ;
	    RECT 748.2000 1163.7001 750.9000 1164.6000 ;
	    RECT 722.1000 1162.2001 727.8000 1163.1000 ;
	    RECT 745.8000 1162.5000 747.0000 1162.8000 ;
	    RECT 716.1000 1161.3000 717.3000 1161.6000 ;
	    RECT 704.7000 1160.4000 717.9000 1161.3000 ;
	    RECT 618.6000 1159.5000 619.8000 1159.8000 ;
	    RECT 474.6000 1158.0000 475.8000 1158.9000 ;
	    RECT 464.4000 1157.1000 465.6000 1158.0000 ;
	    RECT 474.6000 1157.1000 500.1000 1158.0000 ;
	    RECT 501.0000 1157.4000 502.2000 1158.6000 ;
	    RECT 508.5000 1158.0000 509.7000 1158.3000 ;
	    RECT 503.1000 1157.1000 509.7000 1158.0000 ;
	    RECT 414.6000 1155.4501 415.8000 1155.6000 ;
	    RECT 460.2000 1155.4501 461.4000 1155.6000 ;
	    RECT 414.6000 1154.5500 461.4000 1155.4501 ;
	    RECT 462.3000 1155.0000 463.8000 1156.2001 ;
	    RECT 414.6000 1154.4000 415.8000 1154.5500 ;
	    RECT 460.2000 1154.4000 461.4000 1154.5500 ;
	    RECT 462.6000 1153.5000 463.8000 1155.0000 ;
	    RECT 464.7000 1154.4000 465.6000 1157.1000 ;
	    RECT 466.5000 1156.2001 467.7000 1156.5000 ;
	    RECT 466.5000 1155.3000 504.9000 1156.2001 ;
	    RECT 500.7000 1155.0000 501.9000 1155.3000 ;
	    RECT 505.8000 1154.4000 507.0000 1155.6000 ;
	    RECT 464.7000 1153.5000 478.2000 1154.4000 ;
	    RECT 364.2000 1152.4501 365.4000 1152.6000 ;
	    RECT 462.6000 1152.4501 463.8000 1152.6000 ;
	    RECT 364.2000 1151.5500 463.8000 1152.4501 ;
	    RECT 364.2000 1151.4000 365.4000 1151.5500 ;
	    RECT 462.6000 1151.4000 463.8000 1151.5500 ;
	    RECT 464.7000 1151.1000 465.6000 1153.5000 ;
	    RECT 477.0000 1153.2001 478.2000 1153.5000 ;
	    RECT 481.8000 1153.5000 494.7000 1154.4000 ;
	    RECT 481.8000 1153.2001 483.0000 1153.5000 ;
	    RECT 469.5000 1151.4000 473.4000 1152.6000 ;
	    RECT 460.2000 1143.3000 461.4000 1149.3000 ;
	    RECT 462.6000 1143.3000 463.8000 1150.5000 ;
	    RECT 464.7000 1150.2001 468.6000 1151.1000 ;
	    RECT 465.0000 1143.3000 466.2000 1149.3000 ;
	    RECT 467.4000 1143.3000 468.6000 1150.2001 ;
	    RECT 469.8000 1143.3000 471.0000 1149.3000 ;
	    RECT 472.2000 1143.3000 473.4000 1151.4000 ;
	    RECT 474.3000 1150.2001 480.6000 1151.4000 ;
	    RECT 474.6000 1143.3000 475.8000 1149.3000 ;
	    RECT 477.0000 1143.3000 478.2000 1147.5000 ;
	    RECT 479.4000 1143.3000 480.6000 1147.5000 ;
	    RECT 481.8000 1143.3000 483.0000 1147.5000 ;
	    RECT 484.2000 1143.3000 485.4000 1152.6000 ;
	    RECT 489.0000 1151.4000 492.9000 1152.6000 ;
	    RECT 493.8000 1152.3000 494.7000 1153.5000 ;
	    RECT 496.2000 1154.1000 497.4000 1154.4000 ;
	    RECT 496.2000 1153.5000 504.3000 1154.1000 ;
	    RECT 496.2000 1153.2001 505.5000 1153.5000 ;
	    RECT 503.4000 1152.3000 505.5000 1153.2001 ;
	    RECT 493.8000 1151.4000 502.5000 1152.3000 ;
	    RECT 507.0000 1152.0000 509.4000 1153.2001 ;
	    RECT 507.0000 1151.4000 507.9000 1152.0000 ;
	    RECT 486.6000 1143.3000 487.8000 1149.3000 ;
	    RECT 489.0000 1143.3000 490.2000 1150.5000 ;
	    RECT 491.4000 1143.3000 492.6000 1149.3000 ;
	    RECT 493.8000 1143.3000 495.0000 1150.5000 ;
	    RECT 501.6000 1150.2001 507.9000 1151.4000 ;
	    RECT 510.6000 1151.1000 511.8000 1159.5000 ;
	    RECT 554.7000 1158.3000 555.9000 1158.6000 ;
	    RECT 558.6000 1158.4501 559.8000 1158.6000 ;
	    RECT 582.6000 1158.4501 583.8000 1158.6000 ;
	    RECT 554.7000 1157.4000 557.1000 1158.3000 ;
	    RECT 558.6000 1157.5500 583.8000 1158.4501 ;
	    RECT 558.6000 1157.4000 559.8000 1157.5500 ;
	    RECT 582.6000 1157.4000 583.8000 1157.5500 ;
	    RECT 585.0000 1158.4501 586.2000 1158.6000 ;
	    RECT 587.4000 1158.4501 588.6000 1158.6000 ;
	    RECT 611.4000 1158.4501 612.6000 1158.6000 ;
	    RECT 585.0000 1157.5500 612.6000 1158.4501 ;
	    RECT 585.0000 1157.4000 586.2000 1157.5500 ;
	    RECT 587.4000 1157.4000 588.6000 1157.5500 ;
	    RECT 611.4000 1157.4000 612.6000 1157.5500 ;
	    RECT 616.2000 1158.4501 617.4000 1158.6000 ;
	    RECT 618.6000 1158.4501 619.8000 1158.6000 ;
	    RECT 616.2000 1157.5500 619.8000 1158.4501 ;
	    RECT 616.2000 1157.4000 617.4000 1157.5500 ;
	    RECT 618.6000 1157.4000 619.8000 1157.5500 ;
	    RECT 555.9000 1157.1000 557.1000 1157.4000 ;
	    RECT 558.9000 1155.3000 559.8000 1156.5000 ;
	    RECT 508.8000 1150.2001 511.8000 1151.1000 ;
	    RECT 551.4000 1154.4000 555.3000 1155.3000 ;
	    RECT 496.2000 1143.3000 497.4000 1147.5000 ;
	    RECT 498.6000 1143.3000 499.8000 1147.5000 ;
	    RECT 501.0000 1143.3000 502.2000 1149.3000 ;
	    RECT 503.4000 1143.3000 504.6000 1150.2001 ;
	    RECT 508.8000 1149.3000 509.7000 1150.2001 ;
	    RECT 505.8000 1142.4000 507.0000 1149.3000 ;
	    RECT 508.2000 1148.4000 509.7000 1149.3000 ;
	    RECT 508.2000 1143.3000 509.4000 1148.4000 ;
	    RECT 510.6000 1143.3000 511.8000 1149.3000 ;
	    RECT 551.4000 1143.3000 552.6000 1154.4000 ;
	    RECT 554.1000 1154.1000 555.3000 1154.4000 ;
	    RECT 553.8000 1143.3000 555.3000 1153.2001 ;
	    RECT 558.0000 1143.3000 560.4000 1155.3000 ;
	    RECT 563.4000 1154.4000 567.0000 1155.3000 ;
	    RECT 563.4000 1154.1000 564.6000 1154.4000 ;
	    RECT 563.1000 1143.3000 564.6000 1153.2001 ;
	    RECT 565.8000 1143.3000 567.0000 1154.4000 ;
	    RECT 585.0000 1143.3000 586.2000 1149.3000 ;
	    RECT 587.4000 1143.3000 588.6000 1156.5000 ;
	    RECT 589.8000 1154.4000 591.0000 1155.6000 ;
	    RECT 620.7000 1155.3000 621.6000 1160.4000 ;
	    RECT 705.9000 1160.1000 707.1000 1160.4000 ;
	    RECT 703.5000 1158.6000 704.7000 1158.9000 ;
	    RECT 703.5000 1157.7001 708.9000 1158.6000 ;
	    RECT 709.8000 1157.4000 711.0000 1158.6000 ;
	    RECT 700.2000 1156.5000 708.6000 1156.8000 ;
	    RECT 700.2000 1156.2001 708.9000 1156.5000 ;
	    RECT 700.2000 1155.9000 714.9000 1156.2001 ;
	    RECT 589.8000 1153.2001 591.0000 1153.5000 ;
	    RECT 589.8000 1143.3000 591.0000 1149.3000 ;
	    RECT 616.2000 1143.3000 617.4000 1155.3000 ;
	    RECT 620.1000 1154.4000 621.6000 1155.3000 ;
	    RECT 623.4000 1154.4000 624.6000 1155.6000 ;
	    RECT 620.1000 1143.3000 621.3000 1154.4000 ;
	    RECT 622.5000 1152.6000 623.4000 1153.5000 ;
	    RECT 622.2000 1151.4000 623.4000 1152.6000 ;
	    RECT 622.5000 1143.3000 623.7000 1149.3000 ;
	    RECT 625.8000 1146.4501 627.0000 1146.6000 ;
	    RECT 693.0000 1146.4501 694.2000 1146.6000 ;
	    RECT 625.8000 1145.5500 694.2000 1146.4501 ;
	    RECT 625.8000 1145.4000 627.0000 1145.5500 ;
	    RECT 693.0000 1145.4000 694.2000 1145.5500 ;
	    RECT 700.2000 1143.3000 701.4000 1155.9000 ;
	    RECT 707.7000 1155.3000 714.9000 1155.9000 ;
	    RECT 702.6000 1143.3000 703.8000 1155.0000 ;
	    RECT 705.0000 1153.5000 713.1000 1154.4000 ;
	    RECT 705.0000 1153.2001 706.2000 1153.5000 ;
	    RECT 711.9000 1153.2001 713.1000 1153.5000 ;
	    RECT 714.0000 1153.5000 714.9000 1155.3000 ;
	    RECT 717.0000 1155.6000 717.9000 1160.4000 ;
	    RECT 726.6000 1159.5000 727.8000 1162.2001 ;
	    RECT 745.8000 1160.4000 747.0000 1161.6000 ;
	    RECT 748.2000 1159.5000 749.4000 1163.7001 ;
	    RECT 765.0000 1162.5000 766.2000 1169.7001 ;
	    RECT 767.4000 1166.7001 768.6000 1169.7001 ;
	    RECT 796.2000 1168.8000 802.2000 1169.7001 ;
	    RECT 767.4000 1165.5000 768.6000 1165.8000 ;
	    RECT 767.4000 1164.4501 768.6000 1164.6000 ;
	    RECT 777.0000 1164.4501 778.2000 1164.6000 ;
	    RECT 767.4000 1163.5500 778.2000 1164.4501 ;
	    RECT 796.2000 1163.7001 797.4000 1168.8000 ;
	    RECT 798.6000 1163.7001 799.8000 1167.9000 ;
	    RECT 801.0000 1164.0000 802.2000 1168.8000 ;
	    RECT 803.4000 1164.9000 804.6000 1169.7001 ;
	    RECT 805.8000 1164.0000 807.0000 1169.7001 ;
	    RECT 801.0000 1163.7001 807.0000 1164.0000 ;
	    RECT 767.4000 1163.4000 768.6000 1163.5500 ;
	    RECT 777.0000 1163.4000 778.2000 1163.5500 ;
	    RECT 798.6000 1161.6000 799.5000 1163.7001 ;
	    RECT 801.3000 1163.1000 806.7000 1163.7001 ;
	    RECT 817.8000 1162.5000 819.0000 1169.7001 ;
	    RECT 820.2000 1166.7001 821.4000 1169.7001 ;
	    RECT 820.2000 1165.5000 821.4000 1165.8000 ;
	    RECT 820.2000 1163.4000 821.4000 1164.6000 ;
	    RECT 832.2000 1162.5000 833.4000 1169.7001 ;
	    RECT 834.6000 1166.7001 835.8000 1169.7001 ;
	    RECT 849.0000 1166.7001 850.2000 1169.7001 ;
	    RECT 834.6000 1165.5000 835.8000 1165.8000 ;
	    RECT 849.0000 1165.5000 850.2000 1165.8000 ;
	    RECT 834.6000 1164.4501 835.8000 1164.6000 ;
	    RECT 849.0000 1164.4501 850.2000 1164.6000 ;
	    RECT 834.6000 1163.5500 850.2000 1164.4501 ;
	    RECT 834.6000 1163.4000 835.8000 1163.5500 ;
	    RECT 849.0000 1163.4000 850.2000 1163.5500 ;
	    RECT 851.4000 1162.5000 852.6000 1169.7001 ;
	    RECT 870.6000 1166.7001 871.8000 1169.7001 ;
	    RECT 873.0000 1166.7001 874.2000 1169.7001 ;
	    RECT 875.4000 1166.7001 876.6000 1169.7001 ;
	    RECT 911.4000 1168.8000 917.4000 1169.7001 ;
	    RECT 870.6000 1165.5000 871.8000 1165.8000 ;
	    RECT 870.6000 1163.4000 871.8000 1164.6000 ;
	    RECT 873.3000 1162.5000 874.2000 1166.7001 ;
	    RECT 911.4000 1163.7001 912.6000 1168.8000 ;
	    RECT 913.8000 1163.7001 915.0000 1167.9000 ;
	    RECT 916.2000 1164.0000 917.4000 1168.8000 ;
	    RECT 918.6000 1164.9000 919.8000 1169.7001 ;
	    RECT 921.0000 1164.0000 922.2000 1169.7001 ;
	    RECT 964.2000 1167.4501 965.4000 1167.6000 ;
	    RECT 1043.4000 1167.4501 1044.6000 1167.6000 ;
	    RECT 964.2000 1166.5500 1044.6000 1167.4501 ;
	    RECT 1045.8000 1166.7001 1047.0000 1169.7001 ;
	    RECT 964.2000 1166.4000 965.4000 1166.5500 ;
	    RECT 1043.4000 1166.4000 1044.6000 1166.5500 ;
	    RECT 916.2000 1163.7001 922.2000 1164.0000 ;
	    RECT 961.8000 1164.4501 963.0000 1164.6000 ;
	    RECT 1014.6000 1164.4501 1015.8000 1164.6000 ;
	    RECT 765.0000 1161.4501 766.2000 1161.6000 ;
	    RECT 796.2000 1161.4501 797.4000 1161.6000 ;
	    RECT 765.0000 1160.5500 797.4000 1161.4501 ;
	    RECT 798.6000 1160.7001 800.1000 1161.6000 ;
	    RECT 765.0000 1160.4000 766.2000 1160.5500 ;
	    RECT 796.2000 1160.4000 797.4000 1160.5500 ;
	    RECT 801.0000 1160.4000 802.2000 1161.6000 ;
	    RECT 804.6000 1160.7001 804.9000 1162.2001 ;
	    RECT 913.8000 1161.6000 914.7000 1163.7001 ;
	    RECT 916.5000 1163.1000 921.9000 1163.7001 ;
	    RECT 961.8000 1163.5500 1015.8000 1164.4501 ;
	    RECT 1048.2001 1164.0000 1049.4000 1169.7001 ;
	    RECT 961.8000 1163.4000 963.0000 1163.5500 ;
	    RECT 1014.6000 1163.4000 1015.8000 1163.5500 ;
	    RECT 1047.9000 1162.8000 1049.4000 1164.0000 ;
	    RECT 805.8000 1160.4000 807.0000 1161.6000 ;
	    RECT 815.4000 1161.4501 816.6000 1161.6000 ;
	    RECT 817.8000 1161.4501 819.0000 1161.6000 ;
	    RECT 815.4000 1160.5500 819.0000 1161.4501 ;
	    RECT 815.4000 1160.4000 816.6000 1160.5500 ;
	    RECT 817.8000 1160.4000 819.0000 1160.5500 ;
	    RECT 832.2000 1161.4501 833.4000 1161.6000 ;
	    RECT 846.6000 1161.4501 847.8000 1161.6000 ;
	    RECT 832.2000 1160.5500 847.8000 1161.4501 ;
	    RECT 832.2000 1160.4000 833.4000 1160.5500 ;
	    RECT 846.6000 1160.4000 847.8000 1160.5500 ;
	    RECT 849.0000 1161.4501 850.2000 1161.6000 ;
	    RECT 851.4000 1161.4501 852.6000 1161.6000 ;
	    RECT 849.0000 1160.5500 852.6000 1161.4501 ;
	    RECT 849.0000 1160.4000 850.2000 1160.5500 ;
	    RECT 851.4000 1160.4000 852.6000 1160.5500 ;
	    RECT 873.0000 1161.4501 874.2000 1161.6000 ;
	    RECT 875.4000 1161.4501 876.6000 1161.6000 ;
	    RECT 873.0000 1160.5500 876.6000 1161.4501 ;
	    RECT 873.0000 1160.4000 874.2000 1160.5500 ;
	    RECT 875.4000 1160.4000 876.6000 1160.5500 ;
	    RECT 911.4000 1160.4000 912.6000 1161.6000 ;
	    RECT 913.8000 1160.7001 915.3000 1161.6000 ;
	    RECT 916.2000 1160.4000 917.4000 1161.6000 ;
	    RECT 919.8000 1160.7001 920.1000 1162.2001 ;
	    RECT 921.0000 1160.4000 922.2000 1161.6000 ;
	    RECT 798.6000 1159.5000 799.8000 1159.8000 ;
	    RECT 803.4000 1159.5000 804.6000 1159.8000 ;
	    RECT 913.8000 1159.5000 915.0000 1159.8000 ;
	    RECT 918.6000 1159.5000 919.8000 1159.8000 ;
	    RECT 719.4000 1159.2001 720.6000 1159.5000 ;
	    RECT 719.4000 1158.3000 725.1000 1159.2001 ;
	    RECT 723.9000 1158.0000 725.1000 1158.3000 ;
	    RECT 726.6000 1158.4501 727.8000 1158.6000 ;
	    RECT 743.4000 1158.4501 744.6000 1158.6000 ;
	    RECT 726.6000 1157.5500 744.6000 1158.4501 ;
	    RECT 726.6000 1157.4000 727.8000 1157.5500 ;
	    RECT 743.4000 1157.4000 744.6000 1157.5500 ;
	    RECT 748.2000 1158.4501 749.4000 1158.6000 ;
	    RECT 753.0000 1158.4501 754.2000 1158.6000 ;
	    RECT 748.2000 1157.5500 754.2000 1158.4501 ;
	    RECT 748.2000 1157.4000 749.4000 1157.5500 ;
	    RECT 753.0000 1157.4000 754.2000 1157.5500 ;
	    RECT 721.5000 1157.1000 722.7000 1157.4000 ;
	    RECT 721.5000 1156.5000 725.7000 1157.1000 ;
	    RECT 721.5000 1156.2001 727.8000 1156.5000 ;
	    RECT 717.0000 1154.7001 720.6000 1155.6000 ;
	    RECT 716.1000 1153.5000 717.3000 1153.8000 ;
	    RECT 714.0000 1152.6000 717.3000 1153.5000 ;
	    RECT 719.7000 1153.2001 720.6000 1154.7001 ;
	    RECT 719.7000 1152.0000 721.8000 1153.2001 ;
	    RECT 710.1000 1151.1000 711.3000 1151.4000 ;
	    RECT 714.3000 1151.1000 715.5000 1151.4000 ;
	    RECT 705.0000 1149.3000 706.2000 1150.5000 ;
	    RECT 710.1000 1150.2001 715.5000 1151.1000 ;
	    RECT 713.4000 1149.3000 714.3000 1150.2001 ;
	    RECT 719.4000 1149.3000 720.6000 1150.5000 ;
	    RECT 705.0000 1148.4000 708.0000 1149.3000 ;
	    RECT 706.8000 1143.3000 708.0000 1148.4000 ;
	    RECT 711.0000 1143.3000 712.2000 1149.3000 ;
	    RECT 713.4000 1143.3000 714.6000 1149.3000 ;
	    RECT 715.8000 1143.3000 717.0000 1149.3000 ;
	    RECT 719.7000 1143.3000 721.5000 1149.3000 ;
	    RECT 724.2000 1143.3000 725.4000 1155.3000 ;
	    RECT 726.6000 1143.3000 727.8000 1156.2001 ;
	    RECT 745.8000 1143.3000 747.0000 1149.3000 ;
	    RECT 748.2000 1143.3000 749.4000 1156.5000 ;
	    RECT 750.6000 1155.4501 751.8000 1155.6000 ;
	    RECT 755.4000 1155.4501 756.6000 1155.6000 ;
	    RECT 750.6000 1154.5500 756.6000 1155.4501 ;
	    RECT 750.6000 1154.4000 751.8000 1154.5500 ;
	    RECT 755.4000 1154.4000 756.6000 1154.5500 ;
	    RECT 750.6000 1153.2001 751.8000 1153.5000 ;
	    RECT 750.6000 1143.3000 751.8000 1149.3000 ;
	    RECT 765.0000 1143.3000 766.2000 1159.5000 ;
	    RECT 796.2000 1159.2001 797.4000 1159.5000 ;
	    RECT 798.6000 1157.4000 799.8000 1158.6000 ;
	    RECT 801.3000 1155.3000 802.2000 1159.5000 ;
	    RECT 803.4000 1158.4501 804.6000 1158.6000 ;
	    RECT 808.2000 1158.4501 809.4000 1158.6000 ;
	    RECT 803.4000 1157.5500 809.4000 1158.4501 ;
	    RECT 803.4000 1157.4000 804.6000 1157.5500 ;
	    RECT 808.2000 1157.4000 809.4000 1157.5500 ;
	    RECT 767.4000 1143.3000 768.6000 1149.3000 ;
	    RECT 796.2000 1143.3000 797.4000 1155.3000 ;
	    RECT 800.1000 1143.3000 803.1000 1155.3000 ;
	    RECT 805.8000 1143.3000 807.0000 1155.3000 ;
	    RECT 817.8000 1143.3000 819.0000 1159.5000 ;
	    RECT 820.2000 1143.3000 821.4000 1149.3000 ;
	    RECT 832.2000 1143.3000 833.4000 1159.5000 ;
	    RECT 834.6000 1143.3000 835.8000 1149.3000 ;
	    RECT 849.0000 1143.3000 850.2000 1149.3000 ;
	    RECT 851.4000 1143.3000 852.6000 1159.5000 ;
	    RECT 873.3000 1155.3000 874.2000 1159.5000 ;
	    RECT 911.4000 1159.2001 912.6000 1159.5000 ;
	    RECT 875.4000 1158.4501 876.6000 1158.6000 ;
	    RECT 877.8000 1158.4501 879.0000 1158.6000 ;
	    RECT 875.4000 1157.5500 879.0000 1158.4501 ;
	    RECT 875.4000 1157.4000 876.6000 1157.5500 ;
	    RECT 877.8000 1157.4000 879.0000 1157.5500 ;
	    RECT 913.8000 1157.4000 915.0000 1158.6000 ;
	    RECT 875.4000 1156.2001 876.6000 1156.5000 ;
	    RECT 916.5000 1155.3000 917.4000 1159.5000 ;
	    RECT 918.6000 1158.4501 919.8000 1158.6000 ;
	    RECT 954.6000 1158.4501 955.8000 1158.6000 ;
	    RECT 1007.4000 1158.4501 1008.6000 1158.6000 ;
	    RECT 918.6000 1157.5500 1008.6000 1158.4501 ;
	    RECT 918.6000 1157.4000 919.8000 1157.5500 ;
	    RECT 954.6000 1157.4000 955.8000 1157.5500 ;
	    RECT 1007.4000 1157.4000 1008.6000 1157.5500 ;
	    RECT 1047.9000 1156.2001 1049.1000 1162.8000 ;
	    RECT 1050.6000 1161.9000 1051.8000 1169.7001 ;
	    RECT 1055.4000 1163.7001 1056.6000 1169.7001 ;
	    RECT 1060.2001 1164.9000 1061.4000 1169.7001 ;
	    RECT 1062.6000 1165.5000 1063.8000 1169.7001 ;
	    RECT 1065.0000 1165.5000 1066.2001 1169.7001 ;
	    RECT 1067.4000 1165.5000 1068.6000 1169.7001 ;
	    RECT 1069.8000 1165.5000 1071.0000 1169.7001 ;
	    RECT 1072.2001 1166.7001 1073.4000 1169.7001 ;
	    RECT 1074.6000 1165.5000 1075.8000 1169.7001 ;
	    RECT 1077.0000 1166.7001 1078.2001 1169.7001 ;
	    RECT 1079.4000 1165.5000 1080.6000 1169.7001 ;
	    RECT 1081.8000 1165.5000 1083.0000 1169.7001 ;
	    RECT 1084.2001 1165.5000 1085.4000 1169.7001 ;
	    RECT 1057.8000 1163.7001 1061.4000 1164.9000 ;
	    RECT 1086.6000 1164.9000 1087.8000 1169.7001 ;
	    RECT 1057.8000 1162.8000 1059.0000 1163.7001 ;
	    RECT 1050.0000 1161.0000 1051.8000 1161.9000 ;
	    RECT 1056.3000 1161.9000 1059.0000 1162.8000 ;
	    RECT 1065.0000 1163.4000 1066.5000 1164.6000 ;
	    RECT 1071.0000 1163.4000 1071.3000 1164.6000 ;
	    RECT 1072.2001 1163.4000 1073.4000 1164.6000 ;
	    RECT 1074.6000 1163.7001 1081.5000 1164.6000 ;
	    RECT 1086.6000 1163.7001 1090.5000 1164.9000 ;
	    RECT 1091.4000 1163.7001 1092.6000 1169.7001 ;
	    RECT 1074.6000 1163.4000 1075.8000 1163.7001 ;
	    RECT 1050.0000 1158.0000 1050.9000 1161.0000 ;
	    RECT 1056.3000 1160.1000 1057.5000 1161.9000 ;
	    RECT 1051.8000 1158.9000 1057.5000 1160.1000 ;
	    RECT 1065.0000 1159.2001 1066.2001 1163.4000 ;
	    RECT 1077.0000 1162.5000 1078.2001 1162.8000 ;
	    RECT 1074.6000 1162.2001 1075.8000 1162.5000 ;
	    RECT 1069.2001 1161.3000 1075.8000 1162.2001 ;
	    RECT 1069.2001 1161.0000 1070.4000 1161.3000 ;
	    RECT 1077.0000 1160.4000 1078.2001 1161.6000 ;
	    RECT 1080.3000 1160.1000 1081.5000 1163.7001 ;
	    RECT 1089.3000 1162.8000 1090.5000 1163.7001 ;
	    RECT 1089.3000 1161.6000 1093.8000 1162.8000 ;
	    RECT 1096.2001 1160.7001 1097.4000 1169.7001 ;
	    RECT 1115.4000 1163.7001 1116.6000 1169.7001 ;
	    RECT 1119.3000 1164.6000 1120.5000 1169.7001 ;
	    RECT 1117.8000 1163.7001 1120.5000 1164.6000 ;
	    RECT 1115.4000 1162.5000 1116.6000 1162.8000 ;
	    RECT 1069.8000 1158.9000 1074.6000 1160.1000 ;
	    RECT 1080.3000 1158.9000 1083.3000 1160.1000 ;
	    RECT 1084.2001 1159.5000 1097.4000 1160.7001 ;
	    RECT 1110.6000 1161.4501 1111.8000 1161.6000 ;
	    RECT 1115.4000 1161.4501 1116.6000 1161.6000 ;
	    RECT 1110.6000 1160.5500 1116.6000 1161.4501 ;
	    RECT 1110.6000 1160.4000 1111.8000 1160.5500 ;
	    RECT 1115.4000 1160.4000 1116.6000 1160.5500 ;
	    RECT 1117.8000 1159.5000 1119.0000 1163.7001 ;
	    RECT 1141.8000 1162.5000 1143.0000 1169.7001 ;
	    RECT 1144.2001 1166.7001 1145.4000 1169.7001 ;
	    RECT 1156.2001 1166.7001 1157.4000 1169.7001 ;
	    RECT 1144.2001 1165.5000 1145.4000 1165.8000 ;
	    RECT 1156.2001 1165.5000 1157.4000 1165.8000 ;
	    RECT 1144.2001 1163.4000 1145.4000 1164.6000 ;
	    RECT 1156.2001 1163.4000 1157.4000 1164.6000 ;
	    RECT 1158.6000 1162.5000 1159.8000 1169.7001 ;
	    RECT 1185.0000 1163.7001 1186.2001 1169.7001 ;
	    RECT 1187.4000 1164.0000 1188.6000 1169.7001 ;
	    RECT 1189.8000 1164.9000 1191.0000 1169.7001 ;
	    RECT 1192.2001 1164.0000 1193.4000 1169.7001 ;
	    RECT 1317.0000 1166.7001 1318.2001 1169.7001 ;
	    RECT 1319.4000 1164.0000 1320.6000 1169.7001 ;
	    RECT 1187.4000 1163.7001 1193.4000 1164.0000 ;
	    RECT 1185.3000 1162.5000 1186.2001 1163.7001 ;
	    RECT 1187.7001 1163.1000 1193.1000 1163.7001 ;
	    RECT 1319.1000 1162.8000 1320.6000 1164.0000 ;
	    RECT 1122.6000 1161.4501 1123.8000 1161.6000 ;
	    RECT 1141.8000 1161.4501 1143.0000 1161.6000 ;
	    RECT 1122.6000 1160.5500 1143.0000 1161.4501 ;
	    RECT 1122.6000 1160.4000 1123.8000 1160.5500 ;
	    RECT 1141.8000 1160.4000 1143.0000 1160.5500 ;
	    RECT 1158.6000 1161.4501 1159.8000 1161.6000 ;
	    RECT 1182.6000 1161.4501 1183.8000 1161.6000 ;
	    RECT 1158.6000 1160.5500 1183.8000 1161.4501 ;
	    RECT 1158.6000 1160.4000 1159.8000 1160.5500 ;
	    RECT 1182.6000 1160.4000 1183.8000 1160.5500 ;
	    RECT 1185.0000 1160.4000 1186.2001 1161.6000 ;
	    RECT 1187.1000 1160.4000 1188.9000 1161.6000 ;
	    RECT 1191.0000 1160.7001 1191.3000 1162.2001 ;
	    RECT 1192.2001 1161.4501 1193.4000 1161.6000 ;
	    RECT 1223.4000 1161.4501 1224.6000 1161.6000 ;
	    RECT 1192.2001 1160.5500 1224.6000 1161.4501 ;
	    RECT 1192.2001 1160.4000 1193.4000 1160.5500 ;
	    RECT 1223.4000 1160.4000 1224.6000 1160.5500 ;
	    RECT 1060.2001 1158.0000 1061.4000 1158.9000 ;
	    RECT 1050.0000 1157.1000 1051.2001 1158.0000 ;
	    RECT 1060.2001 1157.1000 1085.7001 1158.0000 ;
	    RECT 1086.6000 1157.4000 1087.8000 1158.6000 ;
	    RECT 1094.1000 1158.0000 1095.3000 1158.3000 ;
	    RECT 1088.7001 1157.1000 1095.3000 1158.0000 ;
	    RECT 870.6000 1143.3000 871.8000 1155.3000 ;
	    RECT 873.0000 1154.1000 875.7000 1155.3000 ;
	    RECT 874.5000 1143.3000 875.7000 1154.1000 ;
	    RECT 911.4000 1143.3000 912.6000 1155.3000 ;
	    RECT 915.3000 1143.3000 918.3000 1155.3000 ;
	    RECT 921.0000 1143.3000 922.2000 1155.3000 ;
	    RECT 1047.9000 1155.0000 1049.4000 1156.2001 ;
	    RECT 1048.2001 1153.5000 1049.4000 1155.0000 ;
	    RECT 1050.3000 1154.4000 1051.2001 1157.1000 ;
	    RECT 1052.1000 1156.2001 1053.3000 1156.5000 ;
	    RECT 1052.1000 1155.3000 1090.5000 1156.2001 ;
	    RECT 1086.3000 1155.0000 1087.5000 1155.3000 ;
	    RECT 1091.4000 1154.4000 1092.6000 1155.6000 ;
	    RECT 1050.3000 1153.5000 1063.8000 1154.4000 ;
	    RECT 973.8000 1152.4501 975.0000 1152.6000 ;
	    RECT 1048.2001 1152.4501 1049.4000 1152.6000 ;
	    RECT 973.8000 1151.5500 1049.4000 1152.4501 ;
	    RECT 973.8000 1151.4000 975.0000 1151.5500 ;
	    RECT 1048.2001 1151.4000 1049.4000 1151.5500 ;
	    RECT 1050.3000 1151.1000 1051.2001 1153.5000 ;
	    RECT 1062.6000 1153.2001 1063.8000 1153.5000 ;
	    RECT 1067.4000 1153.5000 1080.3000 1154.4000 ;
	    RECT 1067.4000 1153.2001 1068.6000 1153.5000 ;
	    RECT 1055.1000 1151.4000 1059.0000 1152.6000 ;
	    RECT 1005.0000 1149.4501 1006.2000 1149.6000 ;
	    RECT 1017.0000 1149.4501 1018.2000 1149.6000 ;
	    RECT 1005.0000 1148.5500 1018.2000 1149.4501 ;
	    RECT 1005.0000 1148.4000 1006.2000 1148.5500 ;
	    RECT 1017.0000 1148.4000 1018.2000 1148.5500 ;
	    RECT 923.4000 1146.4501 924.6000 1146.6000 ;
	    RECT 1043.4000 1146.4501 1044.6000 1146.6000 ;
	    RECT 923.4000 1145.5500 1044.6000 1146.4501 ;
	    RECT 923.4000 1145.4000 924.6000 1145.5500 ;
	    RECT 1043.4000 1145.4000 1044.6000 1145.5500 ;
	    RECT 1045.8000 1143.3000 1047.0000 1149.3000 ;
	    RECT 1048.2001 1143.3000 1049.4000 1150.5000 ;
	    RECT 1050.3000 1150.2001 1054.2001 1151.1000 ;
	    RECT 1050.6000 1143.3000 1051.8000 1149.3000 ;
	    RECT 1053.0000 1143.3000 1054.2001 1150.2001 ;
	    RECT 1055.4000 1143.3000 1056.6000 1149.3000 ;
	    RECT 1057.8000 1143.3000 1059.0000 1151.4000 ;
	    RECT 1059.9000 1150.2001 1066.2001 1151.4000 ;
	    RECT 1060.2001 1143.3000 1061.4000 1149.3000 ;
	    RECT 1062.6000 1143.3000 1063.8000 1147.5000 ;
	    RECT 1065.0000 1143.3000 1066.2001 1147.5000 ;
	    RECT 1067.4000 1143.3000 1068.6000 1147.5000 ;
	    RECT 1069.8000 1143.3000 1071.0000 1152.6000 ;
	    RECT 1074.6000 1151.4000 1078.5000 1152.6000 ;
	    RECT 1079.4000 1152.3000 1080.3000 1153.5000 ;
	    RECT 1081.8000 1154.1000 1083.0000 1154.4000 ;
	    RECT 1081.8000 1153.5000 1089.9000 1154.1000 ;
	    RECT 1081.8000 1153.2001 1091.1000 1153.5000 ;
	    RECT 1089.0000 1152.3000 1091.1000 1153.2001 ;
	    RECT 1079.4000 1151.4000 1088.1000 1152.3000 ;
	    RECT 1092.6000 1152.0000 1095.0000 1153.2001 ;
	    RECT 1092.6000 1151.4000 1093.5000 1152.0000 ;
	    RECT 1072.2001 1143.3000 1073.4000 1149.3000 ;
	    RECT 1074.6000 1143.3000 1075.8000 1150.5000 ;
	    RECT 1077.0000 1143.3000 1078.2001 1149.3000 ;
	    RECT 1079.4000 1143.3000 1080.6000 1150.5000 ;
	    RECT 1087.2001 1150.2001 1093.5000 1151.4000 ;
	    RECT 1096.2001 1151.1000 1097.4000 1159.5000 ;
	    RECT 1101.0000 1158.4501 1102.2001 1158.6000 ;
	    RECT 1117.8000 1158.4501 1119.0000 1158.6000 ;
	    RECT 1101.0000 1157.5500 1119.0000 1158.4501 ;
	    RECT 1101.0000 1157.4000 1102.2001 1157.5500 ;
	    RECT 1117.8000 1157.4000 1119.0000 1157.5500 ;
	    RECT 1094.4000 1150.2001 1097.4000 1151.1000 ;
	    RECT 1081.8000 1143.3000 1083.0000 1147.5000 ;
	    RECT 1084.2001 1143.3000 1085.4000 1147.5000 ;
	    RECT 1086.6000 1143.3000 1087.8000 1149.3000 ;
	    RECT 1089.0000 1143.3000 1090.2001 1150.2001 ;
	    RECT 1094.4000 1149.3000 1095.3000 1150.2001 ;
	    RECT 1091.4000 1142.4000 1092.6000 1149.3000 ;
	    RECT 1093.8000 1148.4000 1095.3000 1149.3000 ;
	    RECT 1093.8000 1143.3000 1095.0000 1148.4000 ;
	    RECT 1096.2001 1143.3000 1097.4000 1149.3000 ;
	    RECT 1115.4000 1143.3000 1116.6000 1149.3000 ;
	    RECT 1117.8000 1143.3000 1119.0000 1156.5000 ;
	    RECT 1120.2001 1154.4000 1121.4000 1155.6000 ;
	    RECT 1120.2001 1153.2001 1121.4000 1153.5000 ;
	    RECT 1120.2001 1143.3000 1121.4000 1149.3000 ;
	    RECT 1141.8000 1143.3000 1143.0000 1159.5000 ;
	    RECT 1144.2001 1143.3000 1145.4000 1149.3000 ;
	    RECT 1156.2001 1143.3000 1157.4000 1149.3000 ;
	    RECT 1158.6000 1143.3000 1159.8000 1159.5000 ;
	    RECT 1180.2001 1155.4501 1181.4000 1155.6000 ;
	    RECT 1185.0000 1155.4501 1186.2001 1155.6000 ;
	    RECT 1180.2001 1154.5500 1186.2001 1155.4501 ;
	    RECT 1180.2001 1154.4000 1181.4000 1154.5500 ;
	    RECT 1185.0000 1154.4000 1186.2001 1154.5500 ;
	    RECT 1188.0000 1155.3000 1188.9000 1160.4000 ;
	    RECT 1189.8000 1159.5000 1191.0000 1159.8000 ;
	    RECT 1189.8000 1157.4000 1191.0000 1158.6000 ;
	    RECT 1319.1000 1156.2001 1320.3000 1162.8000 ;
	    RECT 1321.8000 1161.9000 1323.0000 1169.7001 ;
	    RECT 1326.6000 1163.7001 1327.8000 1169.7001 ;
	    RECT 1331.4000 1164.9000 1332.6000 1169.7001 ;
	    RECT 1333.8000 1165.5000 1335.0000 1169.7001 ;
	    RECT 1336.2001 1165.5000 1337.4000 1169.7001 ;
	    RECT 1338.6000 1165.5000 1339.8000 1169.7001 ;
	    RECT 1341.0000 1165.5000 1342.2001 1169.7001 ;
	    RECT 1343.4000 1166.7001 1344.6000 1169.7001 ;
	    RECT 1345.8000 1165.5000 1347.0000 1169.7001 ;
	    RECT 1348.2001 1166.7001 1349.4000 1169.7001 ;
	    RECT 1350.6000 1165.5000 1351.8000 1169.7001 ;
	    RECT 1353.0000 1165.5000 1354.2001 1169.7001 ;
	    RECT 1355.4000 1165.5000 1356.6000 1169.7001 ;
	    RECT 1329.0000 1163.7001 1332.6000 1164.9000 ;
	    RECT 1357.8000 1164.9000 1359.0000 1169.7001 ;
	    RECT 1329.0000 1162.8000 1330.2001 1163.7001 ;
	    RECT 1321.2001 1161.0000 1323.0000 1161.9000 ;
	    RECT 1327.5000 1161.9000 1330.2001 1162.8000 ;
	    RECT 1336.2001 1163.4000 1337.7001 1164.6000 ;
	    RECT 1342.2001 1163.4000 1342.5000 1164.6000 ;
	    RECT 1343.4000 1163.4000 1344.6000 1164.6000 ;
	    RECT 1345.8000 1163.7001 1352.7001 1164.6000 ;
	    RECT 1357.8000 1163.7001 1361.7001 1164.9000 ;
	    RECT 1362.6000 1163.7001 1363.8000 1169.7001 ;
	    RECT 1345.8000 1163.4000 1347.0000 1163.7001 ;
	    RECT 1321.2001 1158.0000 1322.1000 1161.0000 ;
	    RECT 1327.5000 1160.1000 1328.7001 1161.9000 ;
	    RECT 1323.0000 1158.9000 1328.7001 1160.1000 ;
	    RECT 1336.2001 1159.2001 1337.4000 1163.4000 ;
	    RECT 1348.2001 1162.5000 1349.4000 1162.8000 ;
	    RECT 1345.8000 1162.2001 1347.0000 1162.5000 ;
	    RECT 1340.4000 1161.3000 1347.0000 1162.2001 ;
	    RECT 1340.4000 1161.0000 1341.6000 1161.3000 ;
	    RECT 1348.2001 1160.4000 1349.4000 1161.6000 ;
	    RECT 1351.5000 1160.1000 1352.7001 1163.7001 ;
	    RECT 1360.5000 1162.8000 1361.7001 1163.7001 ;
	    RECT 1360.5000 1161.6000 1365.0000 1162.8000 ;
	    RECT 1367.4000 1160.7001 1368.6000 1169.7001 ;
	    RECT 1341.0000 1158.9000 1345.8000 1160.1000 ;
	    RECT 1351.5000 1158.9000 1354.5000 1160.1000 ;
	    RECT 1355.4000 1159.5000 1368.6000 1160.7001 ;
	    RECT 1331.4000 1158.0000 1332.6000 1158.9000 ;
	    RECT 1321.2001 1157.1000 1322.4000 1158.0000 ;
	    RECT 1331.4000 1157.1000 1356.9000 1158.0000 ;
	    RECT 1357.8000 1157.4000 1359.0000 1158.6000 ;
	    RECT 1365.3000 1158.0000 1366.5000 1158.3000 ;
	    RECT 1359.9000 1157.1000 1366.5000 1158.0000 ;
	    RECT 1188.0000 1154.4000 1189.5000 1155.3000 ;
	    RECT 1186.2001 1152.6000 1187.1000 1153.5000 ;
	    RECT 1186.2001 1151.4000 1187.4000 1152.6000 ;
	    RECT 1185.9000 1143.3000 1187.1000 1149.3000 ;
	    RECT 1188.3000 1143.3000 1189.5000 1154.4000 ;
	    RECT 1192.2001 1143.3000 1193.4000 1155.3000 ;
	    RECT 1319.1000 1155.0000 1320.6000 1156.2001 ;
	    RECT 1319.4000 1153.5000 1320.6000 1155.0000 ;
	    RECT 1321.5000 1154.4000 1322.4000 1157.1000 ;
	    RECT 1323.3000 1156.2001 1324.5000 1156.5000 ;
	    RECT 1323.3000 1155.3000 1361.7001 1156.2001 ;
	    RECT 1357.5000 1155.0000 1358.7001 1155.3000 ;
	    RECT 1362.6000 1154.4000 1363.8000 1155.6000 ;
	    RECT 1321.5000 1153.5000 1335.0000 1154.4000 ;
	    RECT 1288.2001 1152.4501 1289.4000 1152.6000 ;
	    RECT 1319.4000 1152.4501 1320.6000 1152.6000 ;
	    RECT 1288.2001 1151.5500 1320.6000 1152.4501 ;
	    RECT 1288.2001 1151.4000 1289.4000 1151.5500 ;
	    RECT 1319.4000 1151.4000 1320.6000 1151.5500 ;
	    RECT 1321.5000 1151.1000 1322.4000 1153.5000 ;
	    RECT 1333.8000 1153.2001 1335.0000 1153.5000 ;
	    RECT 1338.6000 1153.5000 1351.5000 1154.4000 ;
	    RECT 1338.6000 1153.2001 1339.8000 1153.5000 ;
	    RECT 1326.3000 1151.4000 1330.2001 1152.6000 ;
	    RECT 1216.2001 1146.4501 1217.4000 1146.6000 ;
	    RECT 1228.2001 1146.4501 1229.4000 1146.6000 ;
	    RECT 1216.2001 1145.5500 1229.4000 1146.4501 ;
	    RECT 1216.2001 1145.4000 1217.4000 1145.5500 ;
	    RECT 1228.2001 1145.4000 1229.4000 1145.5500 ;
	    RECT 1317.0000 1143.3000 1318.2001 1149.3000 ;
	    RECT 1319.4000 1143.3000 1320.6000 1150.5000 ;
	    RECT 1321.5000 1150.2001 1325.4000 1151.1000 ;
	    RECT 1321.8000 1143.3000 1323.0000 1149.3000 ;
	    RECT 1324.2001 1143.3000 1325.4000 1150.2001 ;
	    RECT 1326.6000 1143.3000 1327.8000 1149.3000 ;
	    RECT 1329.0000 1143.3000 1330.2001 1151.4000 ;
	    RECT 1331.1000 1150.2001 1337.4000 1151.4000 ;
	    RECT 1331.4000 1143.3000 1332.6000 1149.3000 ;
	    RECT 1333.8000 1143.3000 1335.0000 1147.5000 ;
	    RECT 1336.2001 1143.3000 1337.4000 1147.5000 ;
	    RECT 1338.6000 1143.3000 1339.8000 1147.5000 ;
	    RECT 1341.0000 1143.3000 1342.2001 1152.6000 ;
	    RECT 1345.8000 1151.4000 1349.7001 1152.6000 ;
	    RECT 1350.6000 1152.3000 1351.5000 1153.5000 ;
	    RECT 1353.0000 1154.1000 1354.2001 1154.4000 ;
	    RECT 1353.0000 1153.5000 1361.1000 1154.1000 ;
	    RECT 1353.0000 1153.2001 1362.3000 1153.5000 ;
	    RECT 1360.2001 1152.3000 1362.3000 1153.2001 ;
	    RECT 1350.6000 1151.4000 1359.3000 1152.3000 ;
	    RECT 1363.8000 1152.0000 1366.2001 1153.2001 ;
	    RECT 1363.8000 1151.4000 1364.7001 1152.0000 ;
	    RECT 1343.4000 1143.3000 1344.6000 1149.3000 ;
	    RECT 1345.8000 1143.3000 1347.0000 1150.5000 ;
	    RECT 1348.2001 1143.3000 1349.4000 1149.3000 ;
	    RECT 1350.6000 1143.3000 1351.8000 1150.5000 ;
	    RECT 1358.4000 1150.2001 1364.7001 1151.4000 ;
	    RECT 1367.4000 1151.1000 1368.6000 1159.5000 ;
	    RECT 1365.6000 1150.2001 1368.6000 1151.1000 ;
	    RECT 1499.4000 1160.7001 1500.6000 1169.7001 ;
	    RECT 1504.2001 1163.7001 1505.4000 1169.7001 ;
	    RECT 1509.0000 1164.9000 1510.2001 1169.7001 ;
	    RECT 1511.4000 1165.5000 1512.6000 1169.7001 ;
	    RECT 1513.8000 1165.5000 1515.0000 1169.7001 ;
	    RECT 1516.2001 1165.5000 1517.4000 1169.7001 ;
	    RECT 1518.6000 1166.7001 1519.8000 1169.7001 ;
	    RECT 1521.0000 1165.5000 1522.2001 1169.7001 ;
	    RECT 1523.4000 1166.7001 1524.6000 1169.7001 ;
	    RECT 1525.8000 1165.5000 1527.0000 1169.7001 ;
	    RECT 1528.2001 1165.5000 1529.4000 1169.7001 ;
	    RECT 1530.6000 1165.5000 1531.8000 1169.7001 ;
	    RECT 1533.0000 1165.5000 1534.2001 1169.7001 ;
	    RECT 1506.3000 1163.7001 1510.2001 1164.9000 ;
	    RECT 1535.4000 1164.9000 1536.6000 1169.7001 ;
	    RECT 1515.3000 1163.7001 1522.2001 1164.6000 ;
	    RECT 1506.3000 1162.8000 1507.5000 1163.7001 ;
	    RECT 1503.0000 1161.6000 1507.5000 1162.8000 ;
	    RECT 1499.4000 1159.5000 1512.6000 1160.7001 ;
	    RECT 1515.3000 1160.1000 1516.5000 1163.7001 ;
	    RECT 1521.0000 1163.4000 1522.2001 1163.7001 ;
	    RECT 1523.4000 1163.4000 1524.6000 1164.6000 ;
	    RECT 1525.5000 1163.4000 1525.8000 1164.6000 ;
	    RECT 1530.3000 1163.4000 1531.8000 1164.6000 ;
	    RECT 1535.4000 1163.7001 1539.0000 1164.9000 ;
	    RECT 1540.2001 1163.7001 1541.4000 1169.7001 ;
	    RECT 1518.6000 1162.5000 1519.8000 1162.8000 ;
	    RECT 1521.0000 1162.2001 1522.2001 1162.5000 ;
	    RECT 1518.6000 1160.4000 1519.8000 1161.6000 ;
	    RECT 1521.0000 1161.3000 1527.6000 1162.2001 ;
	    RECT 1526.4000 1161.0000 1527.6000 1161.3000 ;
	    RECT 1499.4000 1151.1000 1500.6000 1159.5000 ;
	    RECT 1513.5000 1158.9000 1516.5000 1160.1000 ;
	    RECT 1522.2001 1158.9000 1527.0000 1160.1000 ;
	    RECT 1530.6000 1159.2001 1531.8000 1163.4000 ;
	    RECT 1537.8000 1162.8000 1539.0000 1163.7001 ;
	    RECT 1537.8000 1161.9000 1540.5000 1162.8000 ;
	    RECT 1539.3000 1160.1000 1540.5000 1161.9000 ;
	    RECT 1545.0000 1161.9000 1546.2001 1169.7001 ;
	    RECT 1547.4000 1164.0000 1548.6000 1169.7001 ;
	    RECT 1549.8000 1166.7001 1551.0000 1169.7001 ;
	    RECT 1547.4000 1162.8000 1548.9000 1164.0000 ;
	    RECT 1545.0000 1161.0000 1546.8000 1161.9000 ;
	    RECT 1539.3000 1158.9000 1545.0000 1160.1000 ;
	    RECT 1501.5000 1158.0000 1502.7001 1158.3000 ;
	    RECT 1501.5000 1157.1000 1508.1000 1158.0000 ;
	    RECT 1509.0000 1157.4000 1510.2001 1158.6000 ;
	    RECT 1535.4000 1158.0000 1536.6000 1158.9000 ;
	    RECT 1545.9000 1158.0000 1546.8000 1161.0000 ;
	    RECT 1511.1000 1157.1000 1536.6000 1158.0000 ;
	    RECT 1545.6000 1157.1000 1546.8000 1158.0000 ;
	    RECT 1543.5000 1156.2001 1544.7001 1156.5000 ;
	    RECT 1501.8000 1155.4501 1503.0000 1155.6000 ;
	    RECT 1504.2001 1155.4501 1505.4000 1155.6000 ;
	    RECT 1501.8000 1154.5500 1505.4000 1155.4501 ;
	    RECT 1506.3000 1155.3000 1544.7001 1156.2001 ;
	    RECT 1509.3000 1155.0000 1510.5000 1155.3000 ;
	    RECT 1501.8000 1154.4000 1503.0000 1154.5500 ;
	    RECT 1504.2001 1154.4000 1505.4000 1154.5500 ;
	    RECT 1545.6000 1154.4000 1546.5000 1157.1000 ;
	    RECT 1547.7001 1156.2001 1548.9000 1162.8000 ;
	    RECT 1513.8000 1154.1000 1515.0000 1154.4000 ;
	    RECT 1506.9000 1153.5000 1515.0000 1154.1000 ;
	    RECT 1505.7001 1153.2001 1515.0000 1153.5000 ;
	    RECT 1516.5000 1153.5000 1529.4000 1154.4000 ;
	    RECT 1501.8000 1152.0000 1504.2001 1153.2001 ;
	    RECT 1505.7001 1152.3000 1507.8000 1153.2001 ;
	    RECT 1516.5000 1152.3000 1517.4000 1153.5000 ;
	    RECT 1528.2001 1153.2001 1529.4000 1153.5000 ;
	    RECT 1533.0000 1153.5000 1546.5000 1154.4000 ;
	    RECT 1547.4000 1155.0000 1548.9000 1156.2001 ;
	    RECT 1547.4000 1153.5000 1548.6000 1155.0000 ;
	    RECT 1533.0000 1153.2001 1534.2001 1153.5000 ;
	    RECT 1503.3000 1151.4000 1504.2001 1152.0000 ;
	    RECT 1508.7001 1151.4000 1517.4000 1152.3000 ;
	    RECT 1518.3000 1151.4000 1522.2001 1152.6000 ;
	    RECT 1499.4000 1150.2001 1502.4000 1151.1000 ;
	    RECT 1503.3000 1150.2001 1509.6000 1151.4000 ;
	    RECT 1353.0000 1143.3000 1354.2001 1147.5000 ;
	    RECT 1355.4000 1143.3000 1356.6000 1147.5000 ;
	    RECT 1357.8000 1143.3000 1359.0000 1149.3000 ;
	    RECT 1360.2001 1143.3000 1361.4000 1150.2001 ;
	    RECT 1365.6000 1149.3000 1366.5000 1150.2001 ;
	    RECT 1501.5000 1149.3000 1502.4000 1150.2001 ;
	    RECT 1362.6000 1142.4000 1363.8000 1149.3000 ;
	    RECT 1365.0000 1148.4000 1366.5000 1149.3000 ;
	    RECT 1365.0000 1143.3000 1366.2001 1148.4000 ;
	    RECT 1367.4000 1143.3000 1368.6000 1149.3000 ;
	    RECT 1499.4000 1143.3000 1500.6000 1149.3000 ;
	    RECT 1501.5000 1148.4000 1503.0000 1149.3000 ;
	    RECT 1501.8000 1143.3000 1503.0000 1148.4000 ;
	    RECT 1504.2001 1142.4000 1505.4000 1149.3000 ;
	    RECT 1506.6000 1143.3000 1507.8000 1150.2001 ;
	    RECT 1509.0000 1143.3000 1510.2001 1149.3000 ;
	    RECT 1511.4000 1143.3000 1512.6000 1147.5000 ;
	    RECT 1513.8000 1143.3000 1515.0000 1147.5000 ;
	    RECT 1516.2001 1143.3000 1517.4000 1150.5000 ;
	    RECT 1518.6000 1143.3000 1519.8000 1149.3000 ;
	    RECT 1521.0000 1143.3000 1522.2001 1150.5000 ;
	    RECT 1523.4000 1143.3000 1524.6000 1149.3000 ;
	    RECT 1525.8000 1143.3000 1527.0000 1152.6000 ;
	    RECT 1537.8000 1151.4000 1541.7001 1152.6000 ;
	    RECT 1530.6000 1150.2001 1536.9000 1151.4000 ;
	    RECT 1528.2001 1143.3000 1529.4000 1147.5000 ;
	    RECT 1530.6000 1143.3000 1531.8000 1147.5000 ;
	    RECT 1533.0000 1143.3000 1534.2001 1147.5000 ;
	    RECT 1535.4000 1143.3000 1536.6000 1149.3000 ;
	    RECT 1537.8000 1143.3000 1539.0000 1151.4000 ;
	    RECT 1545.6000 1151.1000 1546.5000 1153.5000 ;
	    RECT 1547.4000 1152.4501 1548.6000 1152.6000 ;
	    RECT 1557.0000 1152.4501 1558.2001 1152.6000 ;
	    RECT 1547.4000 1151.5500 1558.2001 1152.4501 ;
	    RECT 1547.4000 1151.4000 1548.6000 1151.5500 ;
	    RECT 1557.0000 1151.4000 1558.2001 1151.5500 ;
	    RECT 1542.6000 1150.2001 1546.5000 1151.1000 ;
	    RECT 1540.2001 1143.3000 1541.4000 1149.3000 ;
	    RECT 1542.6000 1143.3000 1543.8000 1150.2001 ;
	    RECT 1545.0000 1143.3000 1546.2001 1149.3000 ;
	    RECT 1547.4000 1143.3000 1548.6000 1150.5000 ;
	    RECT 1549.8000 1143.3000 1551.0000 1149.3000 ;
	    RECT 1.2000 1140.6000 1569.0000 1142.4000 ;
	    RECT 124.2000 1133.7001 125.4000 1139.7001 ;
	    RECT 126.6000 1132.5000 127.8000 1139.7001 ;
	    RECT 129.0000 1133.7001 130.2000 1139.7001 ;
	    RECT 131.4000 1132.8000 132.6000 1139.7001 ;
	    RECT 133.8000 1133.7001 135.0000 1139.7001 ;
	    RECT 128.7000 1131.9000 132.6000 1132.8000 ;
	    RECT 126.6000 1130.4000 127.8000 1131.6000 ;
	    RECT 128.7000 1129.5000 129.6000 1131.9000 ;
	    RECT 136.2000 1131.6000 137.4000 1139.7001 ;
	    RECT 138.6000 1133.7001 139.8000 1139.7001 ;
	    RECT 141.0000 1135.5000 142.2000 1139.7001 ;
	    RECT 143.4000 1135.5000 144.6000 1139.7001 ;
	    RECT 145.8000 1135.5000 147.0000 1139.7001 ;
	    RECT 138.3000 1131.6000 144.6000 1132.8000 ;
	    RECT 133.5000 1130.4000 137.4000 1131.6000 ;
	    RECT 148.2000 1130.4000 149.4000 1139.7001 ;
	    RECT 150.6000 1133.7001 151.8000 1139.7001 ;
	    RECT 153.0000 1132.5000 154.2000 1139.7001 ;
	    RECT 155.4000 1133.7001 156.6000 1139.7001 ;
	    RECT 157.8000 1132.5000 159.0000 1139.7001 ;
	    RECT 160.2000 1135.5000 161.4000 1139.7001 ;
	    RECT 162.6000 1135.5000 163.8000 1139.7001 ;
	    RECT 165.0000 1133.7001 166.2000 1139.7001 ;
	    RECT 167.4000 1132.8000 168.6000 1139.7001 ;
	    RECT 169.8000 1133.7001 171.0000 1140.6000 ;
	    RECT 172.2000 1134.6000 173.4000 1139.7001 ;
	    RECT 172.2000 1133.7001 173.7000 1134.6000 ;
	    RECT 174.6000 1133.7001 175.8000 1139.7001 ;
	    RECT 189.0000 1133.7001 190.2000 1139.7001 ;
	    RECT 172.8000 1132.8000 173.7000 1133.7001 ;
	    RECT 165.6000 1131.6000 171.9000 1132.8000 ;
	    RECT 172.8000 1131.9000 175.8000 1132.8000 ;
	    RECT 153.0000 1130.4000 156.9000 1131.6000 ;
	    RECT 157.8000 1130.7001 166.5000 1131.6000 ;
	    RECT 171.0000 1131.0000 171.9000 1131.6000 ;
	    RECT 141.0000 1129.5000 142.2000 1129.8000 ;
	    RECT 126.6000 1128.0000 127.8000 1129.5000 ;
	    RECT 126.3000 1126.8000 127.8000 1128.0000 ;
	    RECT 128.7000 1128.6000 142.2000 1129.5000 ;
	    RECT 145.8000 1129.5000 147.0000 1129.8000 ;
	    RECT 157.8000 1129.5000 158.7000 1130.7001 ;
	    RECT 167.4000 1129.8000 169.5000 1130.7001 ;
	    RECT 171.0000 1129.8000 173.4000 1131.0000 ;
	    RECT 145.8000 1128.6000 158.7000 1129.5000 ;
	    RECT 160.2000 1129.5000 169.5000 1129.8000 ;
	    RECT 160.2000 1128.9000 168.3000 1129.5000 ;
	    RECT 160.2000 1128.6000 161.4000 1128.9000 ;
	    RECT 126.3000 1120.2001 127.5000 1126.8000 ;
	    RECT 128.7000 1125.9000 129.6000 1128.6000 ;
	    RECT 164.7000 1127.7001 165.9000 1128.0000 ;
	    RECT 130.5000 1126.8000 168.9000 1127.7001 ;
	    RECT 169.8000 1127.4000 171.0000 1128.6000 ;
	    RECT 130.5000 1126.5000 131.7000 1126.8000 ;
	    RECT 128.4000 1125.0000 129.6000 1125.9000 ;
	    RECT 138.6000 1125.0000 164.1000 1125.9000 ;
	    RECT 128.4000 1122.0000 129.3000 1125.0000 ;
	    RECT 138.6000 1124.1000 139.8000 1125.0000 ;
	    RECT 165.0000 1124.4000 166.2000 1125.6000 ;
	    RECT 167.1000 1125.0000 173.7000 1125.9000 ;
	    RECT 172.5000 1124.7001 173.7000 1125.0000 ;
	    RECT 130.2000 1122.9000 135.9000 1124.1000 ;
	    RECT 128.4000 1121.1000 130.2000 1122.0000 ;
	    RECT 126.3000 1119.0000 127.8000 1120.2001 ;
	    RECT 124.2000 1113.3000 125.4000 1116.3000 ;
	    RECT 126.6000 1113.3000 127.8000 1119.0000 ;
	    RECT 129.0000 1113.3000 130.2000 1121.1000 ;
	    RECT 134.7000 1121.1000 135.9000 1122.9000 ;
	    RECT 134.7000 1120.2001 137.4000 1121.1000 ;
	    RECT 136.2000 1119.3000 137.4000 1120.2001 ;
	    RECT 143.4000 1119.6000 144.6000 1123.8000 ;
	    RECT 148.2000 1122.9000 153.0000 1124.1000 ;
	    RECT 158.7000 1122.9000 161.7000 1124.1000 ;
	    RECT 174.6000 1123.5000 175.8000 1131.9000 ;
	    RECT 191.4000 1123.5000 192.6000 1139.7001 ;
	    RECT 222.6000 1127.7001 223.8000 1139.7001 ;
	    RECT 226.5000 1128.6000 227.7000 1139.7001 ;
	    RECT 228.9000 1133.7001 230.1000 1139.7001 ;
	    RECT 249.0000 1133.7001 250.2000 1139.7001 ;
	    RECT 228.6000 1130.4000 229.8000 1131.6000 ;
	    RECT 228.9000 1129.5000 229.8000 1130.4000 ;
	    RECT 226.5000 1127.7001 228.0000 1128.6000 ;
	    RECT 225.0000 1125.4501 226.2000 1125.6000 ;
	    RECT 220.3500 1124.5500 226.2000 1125.4501 ;
	    RECT 147.6000 1121.7001 148.8000 1122.0000 ;
	    RECT 147.6000 1120.8000 154.2000 1121.7001 ;
	    RECT 155.4000 1121.4000 156.6000 1122.6000 ;
	    RECT 153.0000 1120.5000 154.2000 1120.8000 ;
	    RECT 155.4000 1120.2001 156.6000 1120.5000 ;
	    RECT 133.8000 1113.3000 135.0000 1119.3000 ;
	    RECT 136.2000 1118.1000 139.8000 1119.3000 ;
	    RECT 143.4000 1118.4000 144.9000 1119.6000 ;
	    RECT 149.4000 1118.4000 149.7000 1119.6000 ;
	    RECT 150.6000 1118.4000 151.8000 1119.6000 ;
	    RECT 153.0000 1119.3000 154.2000 1119.6000 ;
	    RECT 158.7000 1119.3000 159.9000 1122.9000 ;
	    RECT 162.6000 1122.3000 175.8000 1123.5000 ;
	    RECT 167.7000 1120.2001 172.2000 1121.4000 ;
	    RECT 167.7000 1119.3000 168.9000 1120.2001 ;
	    RECT 153.0000 1118.4000 159.9000 1119.3000 ;
	    RECT 138.6000 1113.3000 139.8000 1118.1000 ;
	    RECT 165.0000 1118.1000 168.9000 1119.3000 ;
	    RECT 141.0000 1113.3000 142.2000 1117.5000 ;
	    RECT 143.4000 1113.3000 144.6000 1117.5000 ;
	    RECT 145.8000 1113.3000 147.0000 1117.5000 ;
	    RECT 148.2000 1113.3000 149.4000 1117.5000 ;
	    RECT 150.6000 1113.3000 151.8000 1116.3000 ;
	    RECT 153.0000 1113.3000 154.2000 1117.5000 ;
	    RECT 155.4000 1113.3000 156.6000 1116.3000 ;
	    RECT 157.8000 1113.3000 159.0000 1117.5000 ;
	    RECT 160.2000 1113.3000 161.4000 1117.5000 ;
	    RECT 162.6000 1113.3000 163.8000 1117.5000 ;
	    RECT 165.0000 1113.3000 166.2000 1118.1000 ;
	    RECT 169.8000 1113.3000 171.0000 1119.3000 ;
	    RECT 174.6000 1113.3000 175.8000 1122.3000 ;
	    RECT 191.4000 1122.4501 192.6000 1122.6000 ;
	    RECT 220.3500 1122.4501 221.2500 1124.5500 ;
	    RECT 225.0000 1124.4000 226.2000 1124.5500 ;
	    RECT 225.0000 1123.2001 226.2000 1123.5000 ;
	    RECT 227.1000 1122.6000 228.0000 1127.7001 ;
	    RECT 229.8000 1127.4000 231.0000 1128.6000 ;
	    RECT 251.4000 1126.5000 252.6000 1139.7001 ;
	    RECT 253.8000 1133.7001 255.0000 1139.7001 ;
	    RECT 273.0000 1133.7001 274.2000 1139.7001 ;
	    RECT 253.8000 1129.5000 255.0000 1129.8000 ;
	    RECT 253.8000 1127.4000 255.0000 1128.6000 ;
	    RECT 275.4000 1126.5000 276.6000 1139.7001 ;
	    RECT 277.8000 1133.7001 279.0000 1139.7001 ;
	    RECT 277.8000 1129.5000 279.0000 1129.8000 ;
	    RECT 277.8000 1127.4000 279.0000 1128.6000 ;
	    RECT 297.0000 1127.7001 298.2000 1139.7001 ;
	    RECT 300.9000 1128.9000 302.1000 1139.7001 ;
	    RECT 299.4000 1127.7001 302.1000 1128.9000 ;
	    RECT 325.8000 1127.7001 327.0000 1139.7001 ;
	    RECT 329.7000 1128.6000 330.9000 1139.7001 ;
	    RECT 332.1000 1133.7001 333.3000 1139.7001 ;
	    RECT 331.8000 1130.4000 333.0000 1131.6000 ;
	    RECT 332.1000 1129.5000 333.0000 1130.4000 ;
	    RECT 329.7000 1127.7001 331.2000 1128.6000 ;
	    RECT 234.6000 1125.4501 235.8000 1125.6000 ;
	    RECT 251.4000 1125.4501 252.6000 1125.6000 ;
	    RECT 234.6000 1124.5500 252.6000 1125.4501 ;
	    RECT 234.6000 1124.4000 235.8000 1124.5500 ;
	    RECT 251.4000 1124.4000 252.6000 1124.5500 ;
	    RECT 256.2000 1125.4501 257.4000 1125.6000 ;
	    RECT 275.4000 1125.4501 276.6000 1125.6000 ;
	    RECT 256.2000 1124.5500 276.6000 1125.4501 ;
	    RECT 256.2000 1124.4000 257.4000 1124.5500 ;
	    RECT 275.4000 1124.4000 276.6000 1124.5500 ;
	    RECT 299.7000 1123.5000 300.6000 1127.7001 ;
	    RECT 301.8000 1126.5000 303.0000 1126.8000 ;
	    RECT 301.8000 1125.4501 303.0000 1125.6000 ;
	    RECT 306.6000 1125.4501 307.8000 1125.6000 ;
	    RECT 301.8000 1124.5500 307.8000 1125.4501 ;
	    RECT 301.8000 1124.4000 303.0000 1124.5500 ;
	    RECT 306.6000 1124.4000 307.8000 1124.5500 ;
	    RECT 328.2000 1124.4000 329.4000 1125.6000 ;
	    RECT 191.4000 1121.5500 221.2500 1122.4501 ;
	    RECT 191.4000 1121.4000 192.6000 1121.5500 ;
	    RECT 222.6000 1121.4000 223.8000 1122.6000 ;
	    RECT 224.7000 1120.8000 225.0000 1122.3000 ;
	    RECT 227.1000 1121.4000 228.9000 1122.6000 ;
	    RECT 229.8000 1121.4000 231.0000 1122.6000 ;
	    RECT 232.2000 1122.4501 233.4000 1122.6000 ;
	    RECT 249.0000 1122.4501 250.2000 1122.6000 ;
	    RECT 232.2000 1121.5500 250.2000 1122.4501 ;
	    RECT 232.2000 1121.4000 233.4000 1121.5500 ;
	    RECT 249.0000 1121.4000 250.2000 1121.5500 ;
	    RECT 177.0000 1119.4501 178.2000 1119.6000 ;
	    RECT 179.4000 1119.4501 180.6000 1119.6000 ;
	    RECT 189.0000 1119.4501 190.2000 1119.6000 ;
	    RECT 177.0000 1118.5500 190.2000 1119.4501 ;
	    RECT 177.0000 1118.4000 178.2000 1118.5500 ;
	    RECT 179.4000 1118.4000 180.6000 1118.5500 ;
	    RECT 189.0000 1118.4000 190.2000 1118.5500 ;
	    RECT 189.0000 1117.2001 190.2000 1117.5000 ;
	    RECT 189.0000 1113.3000 190.2000 1116.3000 ;
	    RECT 191.4000 1113.3000 192.6000 1120.5000 ;
	    RECT 222.9000 1119.3000 228.3000 1119.9000 ;
	    RECT 229.8000 1119.3000 230.7000 1120.5000 ;
	    RECT 249.0000 1120.2001 250.2000 1120.5000 ;
	    RECT 251.4000 1119.3000 252.6000 1123.5000 ;
	    RECT 273.0000 1121.4000 274.2000 1122.6000 ;
	    RECT 273.0000 1120.2001 274.2000 1120.5000 ;
	    RECT 275.4000 1119.3000 276.6000 1123.5000 ;
	    RECT 328.2000 1123.2001 329.4000 1123.5000 ;
	    RECT 330.3000 1122.6000 331.2000 1127.7001 ;
	    RECT 333.0000 1127.4000 334.2000 1128.6000 ;
	    RECT 345.0000 1125.4501 346.2000 1125.6000 ;
	    RECT 333.1500 1124.5500 346.2000 1125.4501 ;
	    RECT 333.1500 1122.6000 334.0500 1124.5500 ;
	    RECT 345.0000 1124.4000 346.2000 1124.5500 ;
	    RECT 347.4000 1123.5000 348.6000 1139.7001 ;
	    RECT 349.8000 1133.7001 351.0000 1139.7001 ;
	    RECT 364.2000 1133.7001 365.4000 1139.7001 ;
	    RECT 366.6000 1123.5000 367.8000 1139.7001 ;
	    RECT 390.6000 1127.7001 391.8000 1139.7001 ;
	    RECT 394.5000 1128.6000 395.7000 1139.7001 ;
	    RECT 396.9000 1133.7001 398.1000 1139.7001 ;
	    RECT 417.0000 1133.7001 418.2000 1139.7001 ;
	    RECT 396.6000 1130.4000 397.8000 1131.6000 ;
	    RECT 396.9000 1129.5000 397.8000 1130.4000 ;
	    RECT 417.0000 1129.5000 418.2000 1129.8000 ;
	    RECT 394.5000 1127.7001 396.0000 1128.6000 ;
	    RECT 393.0000 1125.4501 394.2000 1125.6000 ;
	    RECT 388.3500 1124.5500 394.2000 1125.4501 ;
	    RECT 299.4000 1121.4000 300.6000 1122.6000 ;
	    RECT 301.8000 1122.4501 303.0000 1122.6000 ;
	    RECT 325.8000 1122.4501 327.0000 1122.6000 ;
	    RECT 301.8000 1121.5500 327.0000 1122.4501 ;
	    RECT 301.8000 1121.4000 303.0000 1121.5500 ;
	    RECT 325.8000 1121.4000 327.0000 1121.5500 ;
	    RECT 327.9000 1120.8000 328.2000 1122.3000 ;
	    RECT 330.3000 1121.4000 332.1000 1122.6000 ;
	    RECT 333.0000 1121.4000 334.2000 1122.6000 ;
	    RECT 335.4000 1122.4501 336.6000 1122.6000 ;
	    RECT 347.4000 1122.4501 348.6000 1122.6000 ;
	    RECT 335.4000 1121.5500 348.6000 1122.4501 ;
	    RECT 335.4000 1121.4000 336.6000 1121.5500 ;
	    RECT 347.4000 1121.4000 348.6000 1121.5500 ;
	    RECT 366.6000 1122.4501 367.8000 1122.6000 ;
	    RECT 388.3500 1122.4501 389.2500 1124.5500 ;
	    RECT 393.0000 1124.4000 394.2000 1124.5500 ;
	    RECT 393.0000 1123.2001 394.2000 1123.5000 ;
	    RECT 395.1000 1122.6000 396.0000 1127.7001 ;
	    RECT 397.8000 1127.4000 399.0000 1128.6000 ;
	    RECT 417.0000 1127.4000 418.2000 1128.6000 ;
	    RECT 397.9500 1125.4501 398.8500 1127.4000 ;
	    RECT 419.4000 1126.5000 420.6000 1139.7001 ;
	    RECT 421.8000 1133.7001 423.0000 1139.7001 ;
	    RECT 448.2000 1128.6000 449.4000 1139.7001 ;
	    RECT 450.6000 1129.5000 451.8000 1139.7001 ;
	    RECT 448.2000 1127.7001 451.5000 1128.6000 ;
	    RECT 453.0000 1127.7001 454.2000 1139.7001 ;
	    RECT 472.2000 1133.7001 473.4000 1139.7001 ;
	    RECT 450.6000 1126.8000 451.5000 1127.7001 ;
	    RECT 450.6000 1125.6000 452.4000 1126.8000 ;
	    RECT 419.4000 1125.4501 420.6000 1125.6000 ;
	    RECT 397.9500 1124.5500 420.6000 1125.4501 ;
	    RECT 419.4000 1124.4000 420.6000 1124.5500 ;
	    RECT 426.6000 1125.4501 427.8000 1125.6000 ;
	    RECT 448.2000 1125.4501 449.4000 1125.6000 ;
	    RECT 426.6000 1124.5500 449.4000 1125.4501 ;
	    RECT 426.6000 1124.4000 427.8000 1124.5500 ;
	    RECT 448.2000 1124.4000 449.4000 1124.5500 ;
	    RECT 366.6000 1121.5500 389.2500 1122.4501 ;
	    RECT 366.6000 1121.4000 367.8000 1121.5500 ;
	    RECT 390.6000 1121.4000 391.8000 1122.6000 ;
	    RECT 392.7000 1120.8000 393.0000 1122.3000 ;
	    RECT 395.1000 1121.4000 396.9000 1122.6000 ;
	    RECT 397.8000 1122.4501 399.0000 1122.6000 ;
	    RECT 414.6000 1122.4501 415.8000 1122.6000 ;
	    RECT 397.8000 1121.5500 415.8000 1122.4501 ;
	    RECT 397.8000 1121.4000 399.0000 1121.5500 ;
	    RECT 414.6000 1121.4000 415.8000 1121.5500 ;
	    RECT 280.2000 1119.4501 281.4000 1119.6000 ;
	    RECT 297.0000 1119.4501 298.2000 1119.6000 ;
	    RECT 222.6000 1119.0000 228.6000 1119.3000 ;
	    RECT 222.6000 1113.3000 223.8000 1119.0000 ;
	    RECT 225.0000 1113.3000 226.2000 1118.1000 ;
	    RECT 227.4000 1113.3000 228.6000 1119.0000 ;
	    RECT 229.8000 1113.3000 231.0000 1119.3000 ;
	    RECT 249.0000 1113.3000 250.2000 1119.3000 ;
	    RECT 251.4000 1118.4000 254.1000 1119.3000 ;
	    RECT 252.9000 1113.3000 254.1000 1118.4000 ;
	    RECT 273.0000 1113.3000 274.2000 1119.3000 ;
	    RECT 275.4000 1118.4000 278.1000 1119.3000 ;
	    RECT 280.2000 1118.5500 298.2000 1119.4501 ;
	    RECT 280.2000 1118.4000 281.4000 1118.5500 ;
	    RECT 297.0000 1118.4000 298.2000 1118.5500 ;
	    RECT 276.9000 1113.3000 278.1000 1118.4000 ;
	    RECT 297.0000 1117.2001 298.2000 1117.5000 ;
	    RECT 299.7000 1116.3000 300.6000 1120.5000 ;
	    RECT 326.1000 1119.3000 331.5000 1119.9000 ;
	    RECT 333.0000 1119.3000 333.9000 1120.5000 ;
	    RECT 325.8000 1119.0000 331.8000 1119.3000 ;
	    RECT 297.0000 1113.3000 298.2000 1116.3000 ;
	    RECT 299.4000 1113.3000 300.6000 1116.3000 ;
	    RECT 301.8000 1113.3000 303.0000 1116.3000 ;
	    RECT 325.8000 1113.3000 327.0000 1119.0000 ;
	    RECT 328.2000 1113.3000 329.4000 1118.1000 ;
	    RECT 330.6000 1113.3000 331.8000 1119.0000 ;
	    RECT 333.0000 1113.3000 334.2000 1119.3000 ;
	    RECT 347.4000 1113.3000 348.6000 1120.5000 ;
	    RECT 349.8000 1119.4501 351.0000 1119.6000 ;
	    RECT 357.0000 1119.4501 358.2000 1119.6000 ;
	    RECT 349.8000 1118.5500 358.2000 1119.4501 ;
	    RECT 349.8000 1118.4000 351.0000 1118.5500 ;
	    RECT 357.0000 1118.4000 358.2000 1118.5500 ;
	    RECT 364.2000 1118.4000 365.4000 1119.6000 ;
	    RECT 349.8000 1117.2001 351.0000 1117.5000 ;
	    RECT 364.2000 1117.2001 365.4000 1117.5000 ;
	    RECT 349.8000 1113.3000 351.0000 1116.3000 ;
	    RECT 364.2000 1113.3000 365.4000 1116.3000 ;
	    RECT 366.6000 1113.3000 367.8000 1120.5000 ;
	    RECT 390.9000 1119.3000 396.3000 1119.9000 ;
	    RECT 397.8000 1119.3000 398.7000 1120.5000 ;
	    RECT 419.4000 1119.3000 420.6000 1123.5000 ;
	    RECT 448.2000 1123.2001 449.4000 1123.5000 ;
	    RECT 421.8000 1122.4501 423.0000 1122.6000 ;
	    RECT 443.4000 1122.4501 444.6000 1122.6000 ;
	    RECT 421.8000 1121.5500 444.6000 1122.4501 ;
	    RECT 421.8000 1121.4000 423.0000 1121.5500 ;
	    RECT 443.4000 1121.4000 444.6000 1121.5500 ;
	    RECT 450.6000 1121.1000 451.5000 1125.6000 ;
	    RECT 453.3000 1124.4000 454.2000 1127.7001 ;
	    RECT 474.6000 1126.5000 475.8000 1139.7001 ;
	    RECT 477.0000 1133.7001 478.2000 1139.7001 ;
	    RECT 477.0000 1129.5000 478.2000 1129.8000 ;
	    RECT 477.0000 1127.4000 478.2000 1128.6000 ;
	    RECT 501.0000 1127.7001 502.2000 1139.7001 ;
	    RECT 504.9000 1128.6000 506.1000 1139.7001 ;
	    RECT 507.3000 1133.7001 508.5000 1139.7001 ;
	    RECT 633.0000 1133.7001 634.2000 1139.7001 ;
	    RECT 635.4000 1134.6000 636.6000 1139.7001 ;
	    RECT 635.1000 1133.7001 636.6000 1134.6000 ;
	    RECT 637.8000 1133.7001 639.0000 1140.6000 ;
	    RECT 635.1000 1132.8000 636.0000 1133.7001 ;
	    RECT 640.2000 1132.8000 641.4000 1139.7001 ;
	    RECT 642.6000 1133.7001 643.8000 1139.7001 ;
	    RECT 645.0000 1135.5000 646.2000 1139.7001 ;
	    RECT 647.4000 1135.5000 648.6000 1139.7001 ;
	    RECT 633.0000 1131.9000 636.0000 1132.8000 ;
	    RECT 507.0000 1130.4000 508.2000 1131.6000 ;
	    RECT 507.3000 1129.5000 508.2000 1130.4000 ;
	    RECT 504.9000 1127.7001 506.4000 1128.6000 ;
	    RECT 474.6000 1125.4501 475.8000 1125.6000 ;
	    RECT 501.0000 1125.4501 502.2000 1125.6000 ;
	    RECT 474.6000 1124.5500 502.2000 1125.4501 ;
	    RECT 474.6000 1124.4000 475.8000 1124.5500 ;
	    RECT 501.0000 1124.4000 502.2000 1124.5500 ;
	    RECT 503.4000 1124.4000 504.6000 1125.6000 ;
	    RECT 453.0000 1123.5000 454.2000 1124.4000 ;
	    RECT 453.0000 1121.4000 454.2000 1122.6000 ;
	    RECT 460.2000 1122.4501 461.4000 1122.6000 ;
	    RECT 472.2000 1122.4501 473.4000 1122.6000 ;
	    RECT 460.2000 1121.5500 473.4000 1122.4501 ;
	    RECT 460.2000 1121.4000 461.4000 1121.5500 ;
	    RECT 472.2000 1121.4000 473.4000 1121.5500 ;
	    RECT 421.8000 1120.2001 423.0000 1120.5000 ;
	    RECT 448.2000 1120.2001 451.5000 1121.1000 ;
	    RECT 390.6000 1119.0000 396.6000 1119.3000 ;
	    RECT 390.6000 1113.3000 391.8000 1119.0000 ;
	    RECT 393.0000 1113.3000 394.2000 1118.1000 ;
	    RECT 395.4000 1113.3000 396.6000 1119.0000 ;
	    RECT 397.8000 1113.3000 399.0000 1119.3000 ;
	    RECT 417.9000 1118.4000 420.6000 1119.3000 ;
	    RECT 417.9000 1113.3000 419.1000 1118.4000 ;
	    RECT 421.8000 1113.3000 423.0000 1119.3000 ;
	    RECT 448.2000 1113.3000 449.4000 1120.2001 ;
	    RECT 450.6000 1113.3000 451.8000 1119.3000 ;
	    RECT 453.0000 1113.3000 454.2000 1120.5000 ;
	    RECT 472.2000 1120.2001 473.4000 1120.5000 ;
	    RECT 474.6000 1119.3000 475.8000 1123.5000 ;
	    RECT 503.4000 1123.2001 504.6000 1123.5000 ;
	    RECT 505.5000 1122.6000 506.4000 1127.7001 ;
	    RECT 508.2000 1127.4000 509.4000 1128.6000 ;
	    RECT 633.0000 1123.5000 634.2000 1131.9000 ;
	    RECT 636.9000 1131.6000 643.2000 1132.8000 ;
	    RECT 649.8000 1132.5000 651.0000 1139.7001 ;
	    RECT 652.2000 1133.7001 653.4000 1139.7001 ;
	    RECT 654.6000 1132.5000 655.8000 1139.7001 ;
	    RECT 657.0000 1133.7001 658.2000 1139.7001 ;
	    RECT 636.9000 1131.0000 637.8000 1131.6000 ;
	    RECT 635.4000 1129.8000 637.8000 1131.0000 ;
	    RECT 642.3000 1130.7001 651.0000 1131.6000 ;
	    RECT 639.3000 1129.8000 641.4000 1130.7001 ;
	    RECT 639.3000 1129.5000 648.6000 1129.8000 ;
	    RECT 640.5000 1128.9000 648.6000 1129.5000 ;
	    RECT 647.4000 1128.6000 648.6000 1128.9000 ;
	    RECT 650.1000 1129.5000 651.0000 1130.7001 ;
	    RECT 651.9000 1130.4000 655.8000 1131.6000 ;
	    RECT 659.4000 1130.4000 660.6000 1139.7001 ;
	    RECT 661.8000 1135.5000 663.0000 1139.7001 ;
	    RECT 664.2000 1135.5000 665.4000 1139.7001 ;
	    RECT 666.6000 1135.5000 667.8000 1139.7001 ;
	    RECT 669.0000 1133.7001 670.2000 1139.7001 ;
	    RECT 664.2000 1131.6000 670.5000 1132.8000 ;
	    RECT 671.4000 1131.6000 672.6000 1139.7001 ;
	    RECT 673.8000 1133.7001 675.0000 1139.7001 ;
	    RECT 676.2000 1132.8000 677.4000 1139.7001 ;
	    RECT 678.6000 1133.7001 679.8000 1139.7001 ;
	    RECT 676.2000 1131.9000 680.1000 1132.8000 ;
	    RECT 681.0000 1132.5000 682.2000 1139.7001 ;
	    RECT 683.4000 1133.7001 684.6000 1139.7001 ;
	    RECT 712.2000 1139.4000 713.4000 1140.6000 ;
	    RECT 671.4000 1130.4000 675.3000 1131.6000 ;
	    RECT 661.8000 1129.5000 663.0000 1129.8000 ;
	    RECT 650.1000 1128.6000 663.0000 1129.5000 ;
	    RECT 666.6000 1129.5000 667.8000 1129.8000 ;
	    RECT 679.2000 1129.5000 680.1000 1131.9000 ;
	    RECT 681.0000 1131.4501 682.2000 1131.6000 ;
	    RECT 683.4000 1131.4501 684.6000 1131.6000 ;
	    RECT 681.0000 1130.5500 684.6000 1131.4501 ;
	    RECT 681.0000 1130.4000 682.2000 1130.5500 ;
	    RECT 683.4000 1130.4000 684.6000 1130.5500 ;
	    RECT 666.6000 1128.6000 680.1000 1129.5000 ;
	    RECT 637.8000 1127.4000 639.0000 1128.6000 ;
	    RECT 642.9000 1127.7001 644.1000 1128.0000 ;
	    RECT 639.9000 1126.8000 678.3000 1127.7001 ;
	    RECT 677.1000 1126.5000 678.3000 1126.8000 ;
	    RECT 679.2000 1125.9000 680.1000 1128.6000 ;
	    RECT 681.0000 1128.0000 682.2000 1129.5000 ;
	    RECT 681.0000 1126.8000 682.5000 1128.0000 ;
	    RECT 714.6000 1127.7001 715.8000 1139.7001 ;
	    RECT 718.5000 1128.6000 719.7000 1139.7001 ;
	    RECT 720.9000 1133.7001 722.1000 1139.7001 ;
	    RECT 720.6000 1130.4000 721.8000 1131.6000 ;
	    RECT 720.9000 1129.5000 721.8000 1130.4000 ;
	    RECT 718.5000 1127.7001 720.0000 1128.6000 ;
	    RECT 635.1000 1125.0000 641.7000 1125.9000 ;
	    RECT 635.1000 1124.7001 636.3000 1125.0000 ;
	    RECT 642.6000 1124.4000 643.8000 1125.6000 ;
	    RECT 644.7000 1125.0000 670.2000 1125.9000 ;
	    RECT 679.2000 1125.0000 680.4000 1125.9000 ;
	    RECT 669.0000 1124.1000 670.2000 1125.0000 ;
	    RECT 479.4000 1122.4501 480.6000 1122.6000 ;
	    RECT 501.0000 1122.4501 502.2000 1122.6000 ;
	    RECT 479.4000 1121.5500 502.2000 1122.4501 ;
	    RECT 479.4000 1121.4000 480.6000 1121.5500 ;
	    RECT 501.0000 1121.4000 502.2000 1121.5500 ;
	    RECT 503.1000 1120.8000 503.4000 1122.3000 ;
	    RECT 505.5000 1121.4000 507.3000 1122.6000 ;
	    RECT 508.2000 1122.4501 509.4000 1122.6000 ;
	    RECT 587.4000 1122.4501 588.6000 1122.6000 ;
	    RECT 508.2000 1121.5500 588.6000 1122.4501 ;
	    RECT 508.2000 1121.4000 509.4000 1121.5500 ;
	    RECT 587.4000 1121.4000 588.6000 1121.5500 ;
	    RECT 633.0000 1122.3000 646.2000 1123.5000 ;
	    RECT 647.1000 1122.9000 650.1000 1124.1000 ;
	    RECT 655.8000 1122.9000 660.6000 1124.1000 ;
	    RECT 501.3000 1119.3000 506.7000 1119.9000 ;
	    RECT 508.2000 1119.3000 509.1000 1120.5000 ;
	    RECT 472.2000 1113.3000 473.4000 1119.3000 ;
	    RECT 474.6000 1118.4000 477.3000 1119.3000 ;
	    RECT 476.1000 1113.3000 477.3000 1118.4000 ;
	    RECT 501.0000 1119.0000 507.0000 1119.3000 ;
	    RECT 501.0000 1113.3000 502.2000 1119.0000 ;
	    RECT 503.4000 1113.3000 504.6000 1118.1000 ;
	    RECT 505.8000 1113.3000 507.0000 1119.0000 ;
	    RECT 508.2000 1113.3000 509.4000 1119.3000 ;
	    RECT 633.0000 1113.3000 634.2000 1122.3000 ;
	    RECT 636.6000 1120.2001 641.1000 1121.4000 ;
	    RECT 639.9000 1119.3000 641.1000 1120.2001 ;
	    RECT 648.9000 1119.3000 650.1000 1122.9000 ;
	    RECT 652.2000 1121.4000 653.4000 1122.6000 ;
	    RECT 660.0000 1121.7001 661.2000 1122.0000 ;
	    RECT 654.6000 1120.8000 661.2000 1121.7001 ;
	    RECT 654.6000 1120.5000 655.8000 1120.8000 ;
	    RECT 652.2000 1120.2001 653.4000 1120.5000 ;
	    RECT 664.2000 1119.6000 665.4000 1123.8000 ;
	    RECT 672.9000 1122.9000 678.6000 1124.1000 ;
	    RECT 672.9000 1121.1000 674.1000 1122.9000 ;
	    RECT 679.5000 1122.0000 680.4000 1125.0000 ;
	    RECT 654.6000 1119.3000 655.8000 1119.6000 ;
	    RECT 637.8000 1113.3000 639.0000 1119.3000 ;
	    RECT 639.9000 1118.1000 643.8000 1119.3000 ;
	    RECT 648.9000 1118.4000 655.8000 1119.3000 ;
	    RECT 657.0000 1118.4000 658.2000 1119.6000 ;
	    RECT 659.1000 1118.4000 659.4000 1119.6000 ;
	    RECT 663.9000 1118.4000 665.4000 1119.6000 ;
	    RECT 671.4000 1120.2001 674.1000 1121.1000 ;
	    RECT 678.6000 1121.1000 680.4000 1122.0000 ;
	    RECT 671.4000 1119.3000 672.6000 1120.2001 ;
	    RECT 642.6000 1113.3000 643.8000 1118.1000 ;
	    RECT 669.0000 1118.1000 672.6000 1119.3000 ;
	    RECT 645.0000 1113.3000 646.2000 1117.5000 ;
	    RECT 647.4000 1113.3000 648.6000 1117.5000 ;
	    RECT 649.8000 1113.3000 651.0000 1117.5000 ;
	    RECT 652.2000 1113.3000 653.4000 1116.3000 ;
	    RECT 654.6000 1113.3000 655.8000 1117.5000 ;
	    RECT 657.0000 1113.3000 658.2000 1116.3000 ;
	    RECT 659.4000 1113.3000 660.6000 1117.5000 ;
	    RECT 661.8000 1113.3000 663.0000 1117.5000 ;
	    RECT 664.2000 1113.3000 665.4000 1117.5000 ;
	    RECT 666.6000 1113.3000 667.8000 1117.5000 ;
	    RECT 669.0000 1113.3000 670.2000 1118.1000 ;
	    RECT 673.8000 1113.3000 675.0000 1119.3000 ;
	    RECT 678.6000 1113.3000 679.8000 1121.1000 ;
	    RECT 681.3000 1120.2001 682.5000 1126.8000 ;
	    RECT 717.0000 1124.4000 718.2000 1125.6000 ;
	    RECT 717.0000 1123.2001 718.2000 1123.5000 ;
	    RECT 719.1000 1122.6000 720.0000 1127.7001 ;
	    RECT 721.8000 1128.4501 723.0000 1128.6000 ;
	    RECT 726.6000 1128.4501 727.8000 1128.6000 ;
	    RECT 721.8000 1127.5500 727.8000 1128.4501 ;
	    RECT 721.8000 1127.4000 723.0000 1127.5500 ;
	    RECT 726.6000 1127.4000 727.8000 1127.5500 ;
	    RECT 736.2000 1123.5000 737.4000 1139.7001 ;
	    RECT 738.6000 1133.7001 739.8000 1139.7001 ;
	    RECT 757.8000 1133.7001 759.0000 1139.7001 ;
	    RECT 757.8000 1129.5000 759.0000 1129.8000 ;
	    RECT 757.8000 1127.4000 759.0000 1128.6000 ;
	    RECT 760.2000 1126.5000 761.4000 1139.7001 ;
	    RECT 762.6000 1133.7001 763.8000 1139.7001 ;
	    RECT 765.1500 1137.4501 766.0500 1140.6000 ;
	    RECT 767.4000 1137.4501 768.6000 1137.6000 ;
	    RECT 765.1500 1136.5500 768.6000 1137.4501 ;
	    RECT 767.4000 1136.4000 768.6000 1136.5500 ;
	    RECT 781.8000 1127.7001 783.0000 1139.7001 ;
	    RECT 785.7000 1128.9000 786.9000 1139.7001 ;
	    RECT 832.2000 1139.4000 833.4000 1140.6000 ;
	    RECT 808.2000 1137.4501 809.4000 1137.6000 ;
	    RECT 918.6000 1137.4501 919.8000 1137.6000 ;
	    RECT 808.2000 1136.5500 919.8000 1137.4501 ;
	    RECT 808.2000 1136.4000 809.4000 1136.5500 ;
	    RECT 918.6000 1136.4000 919.8000 1136.5500 ;
	    RECT 921.0000 1133.7001 922.2000 1139.7001 ;
	    RECT 923.4000 1134.6000 924.6000 1139.7001 ;
	    RECT 923.1000 1133.7001 924.6000 1134.6000 ;
	    RECT 925.8000 1133.7001 927.0000 1140.6000 ;
	    RECT 923.1000 1132.8000 924.0000 1133.7001 ;
	    RECT 928.2000 1132.8000 929.4000 1139.7001 ;
	    RECT 930.6000 1133.7001 931.8000 1139.7001 ;
	    RECT 933.0000 1135.5000 934.2000 1139.7001 ;
	    RECT 935.4000 1135.5000 936.6000 1139.7001 ;
	    RECT 784.2000 1127.7001 786.9000 1128.9000 ;
	    RECT 921.0000 1131.9000 924.0000 1132.8000 ;
	    RECT 760.2000 1124.4000 761.4000 1125.6000 ;
	    RECT 784.5000 1123.5000 785.4000 1127.7001 ;
	    RECT 786.6000 1126.5000 787.8000 1126.8000 ;
	    RECT 786.6000 1125.4501 787.8000 1125.6000 ;
	    RECT 827.4000 1125.4501 828.6000 1125.6000 ;
	    RECT 786.6000 1124.5500 828.6000 1125.4501 ;
	    RECT 786.6000 1124.4000 787.8000 1124.5500 ;
	    RECT 827.4000 1124.4000 828.6000 1124.5500 ;
	    RECT 921.0000 1123.5000 922.2000 1131.9000 ;
	    RECT 924.9000 1131.6000 931.2000 1132.8000 ;
	    RECT 937.8000 1132.5000 939.0000 1139.7001 ;
	    RECT 940.2000 1133.7001 941.4000 1139.7001 ;
	    RECT 942.6000 1132.5000 943.8000 1139.7001 ;
	    RECT 945.0000 1133.7001 946.2000 1139.7001 ;
	    RECT 924.9000 1131.0000 925.8000 1131.6000 ;
	    RECT 923.4000 1129.8000 925.8000 1131.0000 ;
	    RECT 930.3000 1130.7001 939.0000 1131.6000 ;
	    RECT 927.3000 1129.8000 929.4000 1130.7001 ;
	    RECT 927.3000 1129.5000 936.6000 1129.8000 ;
	    RECT 928.5000 1128.9000 936.6000 1129.5000 ;
	    RECT 935.4000 1128.6000 936.6000 1128.9000 ;
	    RECT 938.1000 1129.5000 939.0000 1130.7001 ;
	    RECT 939.9000 1130.4000 943.8000 1131.6000 ;
	    RECT 947.4000 1130.4000 948.6000 1139.7001 ;
	    RECT 949.8000 1135.5000 951.0000 1139.7001 ;
	    RECT 952.2000 1135.5000 953.4000 1139.7001 ;
	    RECT 954.6000 1135.5000 955.8000 1139.7001 ;
	    RECT 957.0000 1133.7001 958.2000 1139.7001 ;
	    RECT 952.2000 1131.6000 958.5000 1132.8000 ;
	    RECT 959.4000 1131.6000 960.6000 1139.7001 ;
	    RECT 961.8000 1133.7001 963.0000 1139.7001 ;
	    RECT 964.2000 1132.8000 965.4000 1139.7001 ;
	    RECT 966.6000 1133.7001 967.8000 1139.7001 ;
	    RECT 964.2000 1131.9000 968.1000 1132.8000 ;
	    RECT 969.0000 1132.5000 970.2000 1139.7001 ;
	    RECT 971.4000 1133.7001 972.6000 1139.7001 ;
	    RECT 959.4000 1130.4000 963.3000 1131.6000 ;
	    RECT 949.8000 1129.5000 951.0000 1129.8000 ;
	    RECT 938.1000 1128.6000 951.0000 1129.5000 ;
	    RECT 954.6000 1129.5000 955.8000 1129.8000 ;
	    RECT 967.2000 1129.5000 968.1000 1131.9000 ;
	    RECT 969.0000 1130.4000 970.2000 1131.6000 ;
	    RECT 954.6000 1128.6000 968.1000 1129.5000 ;
	    RECT 925.8000 1127.4000 927.0000 1128.6000 ;
	    RECT 930.9000 1127.7001 932.1000 1128.0000 ;
	    RECT 927.9000 1126.8000 966.3000 1127.7001 ;
	    RECT 965.1000 1126.5000 966.3000 1126.8000 ;
	    RECT 967.2000 1125.9000 968.1000 1128.6000 ;
	    RECT 969.0000 1128.0000 970.2000 1129.5000 ;
	    RECT 969.0000 1126.8000 970.5000 1128.0000 ;
	    RECT 1000.2000 1127.7001 1001.4000 1139.7001 ;
	    RECT 1004.1000 1127.7001 1007.1000 1139.7001 ;
	    RECT 1009.8000 1127.7001 1011.0000 1139.7001 ;
	    RECT 1038.6000 1127.7001 1039.8000 1139.7001 ;
	    RECT 1042.5000 1127.7001 1045.5000 1139.7001 ;
	    RECT 1048.2001 1127.7001 1049.4000 1139.7001 ;
	    RECT 1053.0000 1131.4501 1054.2001 1131.6000 ;
	    RECT 1053.0000 1130.5500 1056.4501 1131.4501 ;
	    RECT 1053.0000 1130.4000 1054.2001 1130.5500 ;
	    RECT 923.1000 1125.0000 929.7000 1125.9000 ;
	    RECT 923.1000 1124.7001 924.3000 1125.0000 ;
	    RECT 930.6000 1124.4000 931.8000 1125.6000 ;
	    RECT 932.7000 1125.0000 958.2000 1125.9000 ;
	    RECT 967.2000 1125.0000 968.4000 1125.9000 ;
	    RECT 957.0000 1124.1000 958.2000 1125.0000 ;
	    RECT 712.2000 1122.4501 713.4000 1122.6000 ;
	    RECT 714.6000 1122.4501 715.8000 1122.6000 ;
	    RECT 712.2000 1121.5500 715.8000 1122.4501 ;
	    RECT 712.2000 1121.4000 713.4000 1121.5500 ;
	    RECT 714.6000 1121.4000 715.8000 1121.5500 ;
	    RECT 716.7000 1120.8000 717.0000 1122.3000 ;
	    RECT 719.1000 1121.4000 720.9000 1122.6000 ;
	    RECT 721.8000 1121.4000 723.0000 1122.6000 ;
	    RECT 724.2000 1122.4501 725.4000 1122.6000 ;
	    RECT 736.2000 1122.4501 737.4000 1122.6000 ;
	    RECT 724.2000 1121.5500 737.4000 1122.4501 ;
	    RECT 724.2000 1121.4000 725.4000 1121.5500 ;
	    RECT 736.2000 1121.4000 737.4000 1121.5500 ;
	    RECT 681.0000 1119.0000 682.5000 1120.2001 ;
	    RECT 714.9000 1119.3000 720.3000 1119.9000 ;
	    RECT 721.8000 1119.3000 722.7000 1120.5000 ;
	    RECT 714.6000 1119.0000 720.6000 1119.3000 ;
	    RECT 681.0000 1113.3000 682.2000 1119.0000 ;
	    RECT 683.4000 1113.3000 684.6000 1116.3000 ;
	    RECT 714.6000 1113.3000 715.8000 1119.0000 ;
	    RECT 717.0000 1113.3000 718.2000 1118.1000 ;
	    RECT 719.4000 1113.3000 720.6000 1119.0000 ;
	    RECT 721.8000 1113.3000 723.0000 1119.3000 ;
	    RECT 736.2000 1113.3000 737.4000 1120.5000 ;
	    RECT 738.6000 1119.4501 739.8000 1119.6000 ;
	    RECT 748.2000 1119.4501 749.4000 1119.6000 ;
	    RECT 738.6000 1118.5500 749.4000 1119.4501 ;
	    RECT 760.2000 1119.3000 761.4000 1123.5000 ;
	    RECT 762.6000 1122.4501 763.8000 1122.6000 ;
	    RECT 767.4000 1122.4501 768.6000 1122.6000 ;
	    RECT 762.6000 1121.5500 768.6000 1122.4501 ;
	    RECT 762.6000 1121.4000 763.8000 1121.5500 ;
	    RECT 767.4000 1121.4000 768.6000 1121.5500 ;
	    RECT 784.2000 1122.4501 785.4000 1122.6000 ;
	    RECT 789.0000 1122.4501 790.2000 1122.6000 ;
	    RECT 784.2000 1121.5500 790.2000 1122.4501 ;
	    RECT 784.2000 1121.4000 785.4000 1121.5500 ;
	    RECT 789.0000 1121.4000 790.2000 1121.5500 ;
	    RECT 921.0000 1122.3000 934.2000 1123.5000 ;
	    RECT 935.1000 1122.9000 938.1000 1124.1000 ;
	    RECT 943.8000 1122.9000 948.6000 1124.1000 ;
	    RECT 762.6000 1120.2001 763.8000 1120.5000 ;
	    RECT 738.6000 1118.4000 739.8000 1118.5500 ;
	    RECT 748.2000 1118.4000 749.4000 1118.5500 ;
	    RECT 758.7000 1118.4000 761.4000 1119.3000 ;
	    RECT 738.6000 1117.2001 739.8000 1117.5000 ;
	    RECT 738.6000 1113.3000 739.8000 1116.3000 ;
	    RECT 758.7000 1113.3000 759.9000 1118.4000 ;
	    RECT 762.6000 1113.3000 763.8000 1119.3000 ;
	    RECT 781.8000 1118.4000 783.0000 1119.6000 ;
	    RECT 781.8000 1117.2001 783.0000 1117.5000 ;
	    RECT 784.5000 1116.3000 785.4000 1120.5000 ;
	    RECT 781.8000 1113.3000 783.0000 1116.3000 ;
	    RECT 784.2000 1113.3000 785.4000 1116.3000 ;
	    RECT 786.6000 1113.3000 787.8000 1116.3000 ;
	    RECT 921.0000 1113.3000 922.2000 1122.3000 ;
	    RECT 924.6000 1120.2001 929.1000 1121.4000 ;
	    RECT 927.9000 1119.3000 929.1000 1120.2001 ;
	    RECT 936.9000 1119.3000 938.1000 1122.9000 ;
	    RECT 940.2000 1121.4000 941.4000 1122.6000 ;
	    RECT 948.0000 1121.7001 949.2000 1122.0000 ;
	    RECT 942.6000 1120.8000 949.2000 1121.7001 ;
	    RECT 942.6000 1120.5000 943.8000 1120.8000 ;
	    RECT 940.2000 1120.2001 941.4000 1120.5000 ;
	    RECT 952.2000 1119.6000 953.4000 1123.8000 ;
	    RECT 960.9000 1122.9000 966.6000 1124.1000 ;
	    RECT 960.9000 1121.1000 962.1000 1122.9000 ;
	    RECT 967.5000 1122.0000 968.4000 1125.0000 ;
	    RECT 942.6000 1119.3000 943.8000 1119.6000 ;
	    RECT 925.8000 1113.3000 927.0000 1119.3000 ;
	    RECT 927.9000 1118.1000 931.8000 1119.3000 ;
	    RECT 936.9000 1118.4000 943.8000 1119.3000 ;
	    RECT 945.0000 1118.4000 946.2000 1119.6000 ;
	    RECT 947.1000 1118.4000 947.4000 1119.6000 ;
	    RECT 951.9000 1118.4000 953.4000 1119.6000 ;
	    RECT 959.4000 1120.2001 962.1000 1121.1000 ;
	    RECT 966.6000 1121.1000 968.4000 1122.0000 ;
	    RECT 959.4000 1119.3000 960.6000 1120.2001 ;
	    RECT 930.6000 1113.3000 931.8000 1118.1000 ;
	    RECT 957.0000 1118.1000 960.6000 1119.3000 ;
	    RECT 933.0000 1113.3000 934.2000 1117.5000 ;
	    RECT 935.4000 1113.3000 936.6000 1117.5000 ;
	    RECT 937.8000 1113.3000 939.0000 1117.5000 ;
	    RECT 940.2000 1113.3000 941.4000 1116.3000 ;
	    RECT 942.6000 1113.3000 943.8000 1117.5000 ;
	    RECT 945.0000 1113.3000 946.2000 1116.3000 ;
	    RECT 947.4000 1113.3000 948.6000 1117.5000 ;
	    RECT 949.8000 1113.3000 951.0000 1117.5000 ;
	    RECT 952.2000 1113.3000 953.4000 1117.5000 ;
	    RECT 954.6000 1113.3000 955.8000 1117.5000 ;
	    RECT 957.0000 1113.3000 958.2000 1118.1000 ;
	    RECT 961.8000 1113.3000 963.0000 1119.3000 ;
	    RECT 966.6000 1113.3000 967.8000 1121.1000 ;
	    RECT 969.3000 1120.2001 970.5000 1126.8000 ;
	    RECT 1002.6000 1124.4000 1003.8000 1125.6000 ;
	    RECT 1000.2000 1123.5000 1001.4000 1123.8000 ;
	    RECT 1005.3000 1123.5000 1006.2000 1127.7001 ;
	    RECT 1007.4000 1124.4000 1008.6000 1125.6000 ;
	    RECT 1041.0000 1124.4000 1042.2001 1125.6000 ;
	    RECT 1038.6000 1123.5000 1039.8000 1123.8000 ;
	    RECT 1043.7001 1123.5000 1044.6000 1127.7001 ;
	    RECT 1045.8000 1124.4000 1047.0000 1125.6000 ;
	    RECT 1048.2001 1125.4501 1049.4000 1125.6000 ;
	    RECT 1053.0000 1125.4501 1054.2001 1125.6000 ;
	    RECT 1048.2001 1124.5500 1054.2001 1125.4501 ;
	    RECT 1048.2001 1124.4000 1049.4000 1124.5500 ;
	    RECT 1053.0000 1124.4000 1054.2001 1124.5500 ;
	    RECT 1002.6000 1123.2001 1003.8000 1123.5000 ;
	    RECT 1007.4000 1123.2001 1008.6000 1123.5000 ;
	    RECT 1041.0000 1123.2001 1042.2001 1123.5000 ;
	    RECT 1045.8000 1123.2001 1047.0000 1123.5000 ;
	    RECT 1000.2000 1121.4000 1001.4000 1122.6000 ;
	    RECT 1002.6000 1121.4000 1004.1000 1122.3000 ;
	    RECT 1005.0000 1121.4000 1006.2000 1122.6000 ;
	    RECT 1009.8000 1122.4501 1011.0000 1122.6000 ;
	    RECT 1019.4000 1122.4501 1020.6000 1122.6000 ;
	    RECT 969.0000 1119.0000 970.5000 1120.2001 ;
	    RECT 1002.6000 1119.3000 1003.5000 1121.4000 ;
	    RECT 1008.6000 1120.8000 1008.9000 1122.3000 ;
	    RECT 1009.8000 1121.5500 1020.6000 1122.4501 ;
	    RECT 1009.8000 1121.4000 1011.0000 1121.5500 ;
	    RECT 1019.4000 1121.4000 1020.6000 1121.5500 ;
	    RECT 1038.6000 1121.4000 1039.8000 1122.6000 ;
	    RECT 1041.0000 1121.4000 1042.5000 1122.3000 ;
	    RECT 1043.4000 1121.4000 1044.6000 1122.6000 ;
	    RECT 1048.2001 1122.4501 1049.4000 1122.6000 ;
	    RECT 1055.5500 1122.4501 1056.4501 1130.5500 ;
	    RECT 1060.2001 1123.5000 1061.4000 1139.7001 ;
	    RECT 1062.6000 1133.7001 1063.8000 1139.7001 ;
	    RECT 1081.8000 1133.7001 1083.0000 1139.7001 ;
	    RECT 1084.2001 1126.5000 1085.4000 1139.7001 ;
	    RECT 1086.6000 1133.7001 1087.8000 1139.7001 ;
	    RECT 1218.6000 1133.7001 1219.8000 1139.7001 ;
	    RECT 1221.0000 1134.6000 1222.2001 1139.7001 ;
	    RECT 1220.7001 1133.7001 1222.2001 1134.6000 ;
	    RECT 1223.4000 1133.7001 1224.6000 1140.6000 ;
	    RECT 1220.7001 1132.8000 1221.6000 1133.7001 ;
	    RECT 1225.8000 1132.8000 1227.0000 1139.7001 ;
	    RECT 1228.2001 1133.7001 1229.4000 1139.7001 ;
	    RECT 1230.6000 1135.5000 1231.8000 1139.7001 ;
	    RECT 1233.0000 1135.5000 1234.2001 1139.7001 ;
	    RECT 1218.6000 1131.9000 1221.6000 1132.8000 ;
	    RECT 1086.6000 1129.5000 1087.8000 1129.8000 ;
	    RECT 1086.6000 1128.4501 1087.8000 1128.6000 ;
	    RECT 1091.4000 1128.4501 1092.6000 1128.6000 ;
	    RECT 1086.6000 1127.5500 1092.6000 1128.4501 ;
	    RECT 1086.6000 1127.4000 1087.8000 1127.5500 ;
	    RECT 1091.4000 1127.4000 1092.6000 1127.5500 ;
	    RECT 1084.2001 1125.4501 1085.4000 1125.6000 ;
	    RECT 1216.2001 1125.4501 1217.4000 1125.6000 ;
	    RECT 1084.2001 1124.5500 1217.4000 1125.4501 ;
	    RECT 1084.2001 1124.4000 1085.4000 1124.5500 ;
	    RECT 1216.2001 1124.4000 1217.4000 1124.5500 ;
	    RECT 1218.6000 1123.5000 1219.8000 1131.9000 ;
	    RECT 1222.5000 1131.6000 1228.8000 1132.8000 ;
	    RECT 1235.4000 1132.5000 1236.6000 1139.7001 ;
	    RECT 1237.8000 1133.7001 1239.0000 1139.7001 ;
	    RECT 1240.2001 1132.5000 1241.4000 1139.7001 ;
	    RECT 1242.6000 1133.7001 1243.8000 1139.7001 ;
	    RECT 1222.5000 1131.0000 1223.4000 1131.6000 ;
	    RECT 1221.0000 1129.8000 1223.4000 1131.0000 ;
	    RECT 1227.9000 1130.7001 1236.6000 1131.6000 ;
	    RECT 1224.9000 1129.8000 1227.0000 1130.7001 ;
	    RECT 1224.9000 1129.5000 1234.2001 1129.8000 ;
	    RECT 1226.1000 1128.9000 1234.2001 1129.5000 ;
	    RECT 1233.0000 1128.6000 1234.2001 1128.9000 ;
	    RECT 1235.7001 1129.5000 1236.6000 1130.7001 ;
	    RECT 1237.5000 1130.4000 1241.4000 1131.6000 ;
	    RECT 1245.0000 1130.4000 1246.2001 1139.7001 ;
	    RECT 1247.4000 1135.5000 1248.6000 1139.7001 ;
	    RECT 1249.8000 1135.5000 1251.0000 1139.7001 ;
	    RECT 1252.2001 1135.5000 1253.4000 1139.7001 ;
	    RECT 1254.6000 1133.7001 1255.8000 1139.7001 ;
	    RECT 1249.8000 1131.6000 1256.1000 1132.8000 ;
	    RECT 1257.0000 1131.6000 1258.2001 1139.7001 ;
	    RECT 1259.4000 1133.7001 1260.6000 1139.7001 ;
	    RECT 1261.8000 1132.8000 1263.0000 1139.7001 ;
	    RECT 1264.2001 1133.7001 1265.4000 1139.7001 ;
	    RECT 1261.8000 1131.9000 1265.7001 1132.8000 ;
	    RECT 1266.6000 1132.5000 1267.8000 1139.7001 ;
	    RECT 1269.0000 1133.7001 1270.2001 1139.7001 ;
	    RECT 1281.0000 1133.7001 1282.2001 1139.7001 ;
	    RECT 1257.0000 1130.4000 1260.9000 1131.6000 ;
	    RECT 1247.4000 1129.5000 1248.6000 1129.8000 ;
	    RECT 1235.7001 1128.6000 1248.6000 1129.5000 ;
	    RECT 1252.2001 1129.5000 1253.4000 1129.8000 ;
	    RECT 1264.8000 1129.5000 1265.7001 1131.9000 ;
	    RECT 1266.6000 1131.4501 1267.8000 1131.6000 ;
	    RECT 1269.0000 1131.4501 1270.2001 1131.6000 ;
	    RECT 1266.6000 1130.5500 1270.2001 1131.4501 ;
	    RECT 1266.6000 1130.4000 1267.8000 1130.5500 ;
	    RECT 1269.0000 1130.4000 1270.2001 1130.5500 ;
	    RECT 1252.2001 1128.6000 1265.7001 1129.5000 ;
	    RECT 1223.4000 1127.4000 1224.6000 1128.6000 ;
	    RECT 1228.5000 1127.7001 1229.7001 1128.0000 ;
	    RECT 1225.5000 1126.8000 1263.9000 1127.7001 ;
	    RECT 1262.7001 1126.5000 1263.9000 1126.8000 ;
	    RECT 1264.8000 1125.9000 1265.7001 1128.6000 ;
	    RECT 1266.6000 1128.0000 1267.8000 1129.5000 ;
	    RECT 1266.6000 1126.8000 1268.1000 1128.0000 ;
	    RECT 1220.7001 1125.0000 1227.3000 1125.9000 ;
	    RECT 1220.7001 1124.7001 1221.9000 1125.0000 ;
	    RECT 1228.2001 1124.4000 1229.4000 1125.6000 ;
	    RECT 1230.3000 1125.0000 1255.8000 1125.9000 ;
	    RECT 1264.8000 1125.0000 1266.0000 1125.9000 ;
	    RECT 1254.6000 1124.1000 1255.8000 1125.0000 ;
	    RECT 1005.3000 1119.3000 1010.7000 1119.9000 ;
	    RECT 1041.0000 1119.3000 1041.9000 1121.4000 ;
	    RECT 1047.0000 1120.8000 1047.3000 1122.3000 ;
	    RECT 1048.2001 1121.5500 1056.4501 1122.4501 ;
	    RECT 1048.2001 1121.4000 1049.4000 1121.5500 ;
	    RECT 1060.2001 1121.4000 1061.4000 1122.6000 ;
	    RECT 1081.8000 1122.4501 1083.0000 1122.6000 ;
	    RECT 1062.7500 1121.5500 1083.0000 1122.4501 ;
	    RECT 1043.7001 1119.3000 1049.1000 1119.9000 ;
	    RECT 969.0000 1113.3000 970.2000 1119.0000 ;
	    RECT 971.4000 1113.3000 972.6000 1116.3000 ;
	    RECT 1000.2000 1114.2001 1001.4000 1119.3000 ;
	    RECT 1002.6000 1115.1000 1003.8000 1119.3000 ;
	    RECT 1005.0000 1119.0000 1011.0000 1119.3000 ;
	    RECT 1005.0000 1114.2001 1006.2000 1119.0000 ;
	    RECT 1000.2000 1113.3000 1006.2000 1114.2001 ;
	    RECT 1007.4000 1113.3000 1008.6000 1118.1000 ;
	    RECT 1009.8000 1113.3000 1011.0000 1119.0000 ;
	    RECT 1038.6000 1114.2001 1039.8000 1119.3000 ;
	    RECT 1041.0000 1115.1000 1042.2001 1119.3000 ;
	    RECT 1043.4000 1119.0000 1049.4000 1119.3000 ;
	    RECT 1043.4000 1114.2001 1044.6000 1119.0000 ;
	    RECT 1038.6000 1113.3000 1044.6000 1114.2001 ;
	    RECT 1045.8000 1113.3000 1047.0000 1118.1000 ;
	    RECT 1048.2001 1113.3000 1049.4000 1119.0000 ;
	    RECT 1060.2001 1113.3000 1061.4000 1120.5000 ;
	    RECT 1062.7500 1119.6000 1063.6500 1121.5500 ;
	    RECT 1081.8000 1121.4000 1083.0000 1121.5500 ;
	    RECT 1081.8000 1120.2001 1083.0000 1120.5000 ;
	    RECT 1062.6000 1118.4000 1063.8000 1119.6000 ;
	    RECT 1084.2001 1119.3000 1085.4000 1123.5000 ;
	    RECT 1218.6000 1122.3000 1231.8000 1123.5000 ;
	    RECT 1232.7001 1122.9000 1235.7001 1124.1000 ;
	    RECT 1241.4000 1122.9000 1246.2001 1124.1000 ;
	    RECT 1062.6000 1117.2001 1063.8000 1117.5000 ;
	    RECT 1062.6000 1113.3000 1063.8000 1116.3000 ;
	    RECT 1081.8000 1113.3000 1083.0000 1119.3000 ;
	    RECT 1084.2001 1118.4000 1086.9000 1119.3000 ;
	    RECT 1085.7001 1113.3000 1086.9000 1118.4000 ;
	    RECT 1218.6000 1113.3000 1219.8000 1122.3000 ;
	    RECT 1222.2001 1120.2001 1226.7001 1121.4000 ;
	    RECT 1225.5000 1119.3000 1226.7001 1120.2001 ;
	    RECT 1234.5000 1119.3000 1235.7001 1122.9000 ;
	    RECT 1237.8000 1121.4000 1239.0000 1122.6000 ;
	    RECT 1245.6000 1121.7001 1246.8000 1122.0000 ;
	    RECT 1240.2001 1120.8000 1246.8000 1121.7001 ;
	    RECT 1240.2001 1120.5000 1241.4000 1120.8000 ;
	    RECT 1237.8000 1120.2001 1239.0000 1120.5000 ;
	    RECT 1249.8000 1119.6000 1251.0000 1123.8000 ;
	    RECT 1258.5000 1122.9000 1264.2001 1124.1000 ;
	    RECT 1258.5000 1121.1000 1259.7001 1122.9000 ;
	    RECT 1265.1000 1122.0000 1266.0000 1125.0000 ;
	    RECT 1240.2001 1119.3000 1241.4000 1119.6000 ;
	    RECT 1223.4000 1113.3000 1224.6000 1119.3000 ;
	    RECT 1225.5000 1118.1000 1229.4000 1119.3000 ;
	    RECT 1234.5000 1118.4000 1241.4000 1119.3000 ;
	    RECT 1242.6000 1118.4000 1243.8000 1119.6000 ;
	    RECT 1244.7001 1118.4000 1245.0000 1119.6000 ;
	    RECT 1249.5000 1118.4000 1251.0000 1119.6000 ;
	    RECT 1257.0000 1120.2001 1259.7001 1121.1000 ;
	    RECT 1264.2001 1121.1000 1266.0000 1122.0000 ;
	    RECT 1257.0000 1119.3000 1258.2001 1120.2001 ;
	    RECT 1228.2001 1113.3000 1229.4000 1118.1000 ;
	    RECT 1254.6000 1118.1000 1258.2001 1119.3000 ;
	    RECT 1230.6000 1113.3000 1231.8000 1117.5000 ;
	    RECT 1233.0000 1113.3000 1234.2001 1117.5000 ;
	    RECT 1235.4000 1113.3000 1236.6000 1117.5000 ;
	    RECT 1237.8000 1113.3000 1239.0000 1116.3000 ;
	    RECT 1240.2001 1113.3000 1241.4000 1117.5000 ;
	    RECT 1242.6000 1113.3000 1243.8000 1116.3000 ;
	    RECT 1245.0000 1113.3000 1246.2001 1117.5000 ;
	    RECT 1247.4000 1113.3000 1248.6000 1117.5000 ;
	    RECT 1249.8000 1113.3000 1251.0000 1117.5000 ;
	    RECT 1252.2001 1113.3000 1253.4000 1117.5000 ;
	    RECT 1254.6000 1113.3000 1255.8000 1118.1000 ;
	    RECT 1259.4000 1113.3000 1260.6000 1119.3000 ;
	    RECT 1264.2001 1113.3000 1265.4000 1121.1000 ;
	    RECT 1266.9000 1120.2001 1268.1000 1126.8000 ;
	    RECT 1283.4000 1123.5000 1284.6000 1139.7001 ;
	    RECT 1310.7001 1133.7001 1311.9000 1139.7001 ;
	    RECT 1311.0000 1130.4000 1312.2001 1131.6000 ;
	    RECT 1311.0000 1129.5000 1311.9000 1130.4000 ;
	    RECT 1313.1000 1128.6000 1314.3000 1139.7001 ;
	    RECT 1309.8000 1127.4000 1311.0000 1128.6000 ;
	    RECT 1312.8000 1127.7001 1314.3000 1128.6000 ;
	    RECT 1317.0000 1127.7001 1318.2001 1139.7001 ;
	    RECT 1344.3000 1133.7001 1345.5000 1139.7001 ;
	    RECT 1344.6000 1130.4000 1345.8000 1131.6000 ;
	    RECT 1344.6000 1129.5000 1345.5000 1130.4000 ;
	    RECT 1346.7001 1128.6000 1347.9000 1139.7001 ;
	    RECT 1285.8000 1125.4501 1287.0000 1125.6000 ;
	    RECT 1285.8000 1124.5500 1310.8500 1125.4501 ;
	    RECT 1285.8000 1124.4000 1287.0000 1124.5500 ;
	    RECT 1309.9501 1122.6000 1310.8500 1124.5500 ;
	    RECT 1312.8000 1122.6000 1313.7001 1127.7001 ;
	    RECT 1343.4000 1127.4000 1344.6000 1128.6000 ;
	    RECT 1346.4000 1127.7001 1347.9000 1128.6000 ;
	    RECT 1350.6000 1127.7001 1351.8000 1139.7001 ;
	    RECT 1314.6000 1124.4000 1315.8000 1125.6000 ;
	    RECT 1314.6000 1123.2001 1315.8000 1123.5000 ;
	    RECT 1346.4000 1122.6000 1347.3000 1127.7001 ;
	    RECT 1348.2001 1125.4501 1349.4000 1125.6000 ;
	    RECT 1348.2001 1124.5500 1366.0500 1125.4501 ;
	    RECT 1348.2001 1124.4000 1349.4000 1124.5500 ;
	    RECT 1348.2001 1123.2001 1349.4000 1123.5000 ;
	    RECT 1283.4000 1122.4501 1284.6000 1122.6000 ;
	    RECT 1307.4000 1122.4501 1308.6000 1122.6000 ;
	    RECT 1283.4000 1121.5500 1308.6000 1122.4501 ;
	    RECT 1283.4000 1121.4000 1284.6000 1121.5500 ;
	    RECT 1307.4000 1121.4000 1308.6000 1121.5500 ;
	    RECT 1309.8000 1121.4000 1311.0000 1122.6000 ;
	    RECT 1311.9000 1121.4000 1313.7001 1122.6000 ;
	    RECT 1315.8000 1120.8000 1316.1000 1122.3000 ;
	    RECT 1317.0000 1121.4000 1318.2001 1122.6000 ;
	    RECT 1319.4000 1122.4501 1320.6000 1122.6000 ;
	    RECT 1343.4000 1122.4501 1344.6000 1122.6000 ;
	    RECT 1319.4000 1121.5500 1344.6000 1122.4501 ;
	    RECT 1319.4000 1121.4000 1320.6000 1121.5500 ;
	    RECT 1343.4000 1121.4000 1344.6000 1121.5500 ;
	    RECT 1345.5000 1121.4000 1347.3000 1122.6000 ;
	    RECT 1350.6000 1122.4501 1351.8000 1122.6000 ;
	    RECT 1362.6000 1122.4501 1363.8000 1122.6000 ;
	    RECT 1349.4000 1120.8000 1349.7001 1122.3000 ;
	    RECT 1350.6000 1121.5500 1363.8000 1122.4501 ;
	    RECT 1365.1500 1122.4501 1366.0500 1124.5500 ;
	    RECT 1369.8000 1123.5000 1371.0000 1139.7001 ;
	    RECT 1372.2001 1133.7001 1373.4000 1139.7001 ;
	    RECT 1386.6000 1133.7001 1387.8000 1139.7001 ;
	    RECT 1389.0000 1123.5000 1390.2001 1139.7001 ;
	    RECT 1408.2001 1133.7001 1409.4000 1139.7001 ;
	    RECT 1408.2001 1129.5000 1409.4000 1129.8000 ;
	    RECT 1391.4000 1128.4501 1392.6000 1128.6000 ;
	    RECT 1408.2001 1128.4501 1409.4000 1128.6000 ;
	    RECT 1391.4000 1127.5500 1409.4000 1128.4501 ;
	    RECT 1391.4000 1127.4000 1392.6000 1127.5500 ;
	    RECT 1408.2001 1127.4000 1409.4000 1127.5500 ;
	    RECT 1410.6000 1126.5000 1411.8000 1139.7001 ;
	    RECT 1413.0000 1133.7001 1414.2001 1139.7001 ;
	    RECT 1393.8000 1125.4501 1395.0000 1125.6000 ;
	    RECT 1410.6000 1125.4501 1411.8000 1125.6000 ;
	    RECT 1393.8000 1124.5500 1411.8000 1125.4501 ;
	    RECT 1393.8000 1124.4000 1395.0000 1124.5500 ;
	    RECT 1410.6000 1124.4000 1411.8000 1124.5500 ;
	    RECT 1425.0000 1123.5000 1426.2001 1139.7001 ;
	    RECT 1427.4000 1133.7001 1428.6000 1139.7001 ;
	    RECT 1497.0000 1126.8000 1498.2001 1139.7001 ;
	    RECT 1499.4000 1127.7001 1500.6000 1139.7001 ;
	    RECT 1503.3000 1133.7001 1505.1000 1139.7001 ;
	    RECT 1507.8000 1133.7001 1509.0000 1139.7001 ;
	    RECT 1510.2001 1133.7001 1511.4000 1139.7001 ;
	    RECT 1512.6000 1133.7001 1513.8000 1139.7001 ;
	    RECT 1516.8000 1134.6000 1518.0000 1139.7001 ;
	    RECT 1516.8000 1133.7001 1519.8000 1134.6000 ;
	    RECT 1504.2001 1132.5000 1505.4000 1133.7001 ;
	    RECT 1510.5000 1132.8000 1511.4000 1133.7001 ;
	    RECT 1509.3000 1131.9000 1514.7001 1132.8000 ;
	    RECT 1518.6000 1132.5000 1519.8000 1133.7001 ;
	    RECT 1509.3000 1131.6000 1510.5000 1131.9000 ;
	    RECT 1513.5000 1131.6000 1514.7001 1131.9000 ;
	    RECT 1503.0000 1129.8000 1505.1000 1131.0000 ;
	    RECT 1504.2001 1128.3000 1505.1000 1129.8000 ;
	    RECT 1507.5000 1129.5000 1510.8000 1130.4000 ;
	    RECT 1507.5000 1129.2001 1508.7001 1129.5000 ;
	    RECT 1504.2001 1127.4000 1507.8000 1128.3000 ;
	    RECT 1497.0000 1126.5000 1503.3000 1126.8000 ;
	    RECT 1499.1000 1125.9000 1503.3000 1126.5000 ;
	    RECT 1502.1000 1125.6000 1503.3000 1125.9000 ;
	    RECT 1449.0000 1125.4501 1450.2001 1125.6000 ;
	    RECT 1497.0000 1125.4501 1498.2001 1125.6000 ;
	    RECT 1449.0000 1124.5500 1498.2001 1125.4501 ;
	    RECT 1449.0000 1124.4000 1450.2001 1124.5500 ;
	    RECT 1497.0000 1124.4000 1498.2001 1124.5500 ;
	    RECT 1499.7001 1124.7001 1500.9000 1125.0000 ;
	    RECT 1499.7001 1123.8000 1505.4000 1124.7001 ;
	    RECT 1504.2001 1123.5000 1505.4000 1123.8000 ;
	    RECT 1369.8000 1122.4501 1371.0000 1122.6000 ;
	    RECT 1365.1500 1121.5500 1371.0000 1122.4501 ;
	    RECT 1350.6000 1121.4000 1351.8000 1121.5500 ;
	    RECT 1362.6000 1121.4000 1363.8000 1121.5500 ;
	    RECT 1369.8000 1121.4000 1371.0000 1121.5500 ;
	    RECT 1374.6000 1122.4501 1375.8000 1122.6000 ;
	    RECT 1389.0000 1122.4501 1390.2001 1122.6000 ;
	    RECT 1374.6000 1121.5500 1390.2001 1122.4501 ;
	    RECT 1374.6000 1121.4000 1375.8000 1121.5500 ;
	    RECT 1389.0000 1121.4000 1390.2001 1121.5500 ;
	    RECT 1266.6000 1119.0000 1268.1000 1120.2001 ;
	    RECT 1269.0000 1119.4501 1270.2001 1119.6000 ;
	    RECT 1281.0000 1119.4501 1282.2001 1119.6000 ;
	    RECT 1266.6000 1113.3000 1267.8000 1119.0000 ;
	    RECT 1269.0000 1118.5500 1282.2001 1119.4501 ;
	    RECT 1269.0000 1118.4000 1270.2001 1118.5500 ;
	    RECT 1281.0000 1118.4000 1282.2001 1118.5500 ;
	    RECT 1281.0000 1117.2001 1282.2001 1117.5000 ;
	    RECT 1269.0000 1113.3000 1270.2001 1116.3000 ;
	    RECT 1281.0000 1113.3000 1282.2001 1116.3000 ;
	    RECT 1283.4000 1113.3000 1284.6000 1120.5000 ;
	    RECT 1310.1000 1119.3000 1311.0000 1120.5000 ;
	    RECT 1312.5000 1119.3000 1317.9000 1119.9000 ;
	    RECT 1343.7001 1119.3000 1344.6000 1120.5000 ;
	    RECT 1346.1000 1119.3000 1351.5000 1119.9000 ;
	    RECT 1309.8000 1113.3000 1311.0000 1119.3000 ;
	    RECT 1312.2001 1119.0000 1318.2001 1119.3000 ;
	    RECT 1312.2001 1113.3000 1313.4000 1119.0000 ;
	    RECT 1314.6000 1113.3000 1315.8000 1118.1000 ;
	    RECT 1317.0000 1113.3000 1318.2001 1119.0000 ;
	    RECT 1343.4000 1113.3000 1344.6000 1119.3000 ;
	    RECT 1345.8000 1119.0000 1351.8000 1119.3000 ;
	    RECT 1345.8000 1113.3000 1347.0000 1119.0000 ;
	    RECT 1348.2001 1113.3000 1349.4000 1118.1000 ;
	    RECT 1350.6000 1113.3000 1351.8000 1119.0000 ;
	    RECT 1369.8000 1113.3000 1371.0000 1120.5000 ;
	    RECT 1372.2001 1118.4000 1373.4000 1119.6000 ;
	    RECT 1384.2001 1119.4501 1385.4000 1119.6000 ;
	    RECT 1386.6000 1119.4501 1387.8000 1119.6000 ;
	    RECT 1384.2001 1118.5500 1387.8000 1119.4501 ;
	    RECT 1384.2001 1118.4000 1385.4000 1118.5500 ;
	    RECT 1386.6000 1118.4000 1387.8000 1118.5500 ;
	    RECT 1372.2001 1117.2001 1373.4000 1117.5000 ;
	    RECT 1386.6000 1117.2001 1387.8000 1117.5000 ;
	    RECT 1372.2001 1113.3000 1373.4000 1116.3000 ;
	    RECT 1386.6000 1113.3000 1387.8000 1116.3000 ;
	    RECT 1389.0000 1113.3000 1390.2001 1120.5000 ;
	    RECT 1410.6000 1119.3000 1411.8000 1123.5000 ;
	    RECT 1413.0000 1121.4000 1414.2001 1122.6000 ;
	    RECT 1425.0000 1122.4501 1426.2001 1122.6000 ;
	    RECT 1470.6000 1122.4501 1471.8000 1122.6000 ;
	    RECT 1425.0000 1121.5500 1471.8000 1122.4501 ;
	    RECT 1425.0000 1121.4000 1426.2001 1121.5500 ;
	    RECT 1470.6000 1121.4000 1471.8000 1121.5500 ;
	    RECT 1497.0000 1120.8000 1498.2001 1123.5000 ;
	    RECT 1506.9000 1122.6000 1507.8000 1127.4000 ;
	    RECT 1509.9000 1127.7001 1510.8000 1129.5000 ;
	    RECT 1511.7001 1129.5000 1512.9000 1129.8000 ;
	    RECT 1518.6000 1129.5000 1519.8000 1129.8000 ;
	    RECT 1511.7001 1128.6000 1519.8000 1129.5000 ;
	    RECT 1521.0000 1128.0000 1522.2001 1139.7001 ;
	    RECT 1509.9000 1127.1000 1517.1000 1127.7001 ;
	    RECT 1523.4000 1127.1000 1524.6000 1139.7001 ;
	    RECT 1533.0000 1139.4000 1534.2001 1140.6000 ;
	    RECT 1542.6000 1133.7001 1543.8000 1139.7001 ;
	    RECT 1509.9000 1126.8000 1524.6000 1127.1000 ;
	    RECT 1515.9000 1126.5000 1524.6000 1126.8000 ;
	    RECT 1545.0000 1126.5000 1546.2001 1139.7001 ;
	    RECT 1547.4000 1133.7001 1548.6000 1139.7001 ;
	    RECT 1547.4000 1129.5000 1548.6000 1129.8000 ;
	    RECT 1516.2001 1126.2001 1524.6000 1126.5000 ;
	    RECT 1513.8000 1124.4000 1515.0000 1125.6000 ;
	    RECT 1525.8000 1125.4501 1527.0000 1125.6000 ;
	    RECT 1545.0000 1125.4501 1546.2001 1125.6000 ;
	    RECT 1515.9000 1124.4000 1521.3000 1125.3000 ;
	    RECT 1525.8000 1124.5500 1546.2001 1125.4501 ;
	    RECT 1525.8000 1124.4000 1527.0000 1124.5500 ;
	    RECT 1545.0000 1124.4000 1546.2001 1124.5500 ;
	    RECT 1520.1000 1124.1000 1521.3000 1124.4000 ;
	    RECT 1517.7001 1122.6000 1518.9000 1122.9000 ;
	    RECT 1506.9000 1121.7001 1520.1000 1122.6000 ;
	    RECT 1507.5000 1121.4000 1508.7001 1121.7001 ;
	    RECT 1413.0000 1120.2001 1414.2001 1120.5000 ;
	    RECT 1409.1000 1118.4000 1411.8000 1119.3000 ;
	    RECT 1409.1000 1113.3000 1410.3000 1118.4000 ;
	    RECT 1413.0000 1113.3000 1414.2001 1119.3000 ;
	    RECT 1425.0000 1113.3000 1426.2001 1120.5000 ;
	    RECT 1497.0000 1119.9000 1502.7001 1120.8000 ;
	    RECT 1427.4000 1118.4000 1428.6000 1119.6000 ;
	    RECT 1427.4000 1117.2001 1428.6000 1117.5000 ;
	    RECT 1427.4000 1113.3000 1428.6000 1116.3000 ;
	    RECT 1497.0000 1113.3000 1498.2001 1119.9000 ;
	    RECT 1501.5000 1119.6000 1502.7001 1119.9000 ;
	    RECT 1499.4000 1113.3000 1500.6000 1119.0000 ;
	    RECT 1516.2001 1118.4000 1517.1000 1121.7001 ;
	    RECT 1521.0000 1121.4000 1522.2001 1122.6000 ;
	    RECT 1523.1000 1121.4000 1523.4000 1122.6000 ;
	    RECT 1533.0000 1122.4501 1534.2001 1122.6000 ;
	    RECT 1542.6000 1122.4501 1543.8000 1122.6000 ;
	    RECT 1533.0000 1121.5500 1543.8000 1122.4501 ;
	    RECT 1533.0000 1121.4000 1534.2001 1121.5500 ;
	    RECT 1542.6000 1121.4000 1543.8000 1121.5500 ;
	    RECT 1513.5000 1118.1000 1514.7001 1118.4000 ;
	    RECT 1504.2001 1116.3000 1505.4000 1117.5000 ;
	    RECT 1510.5000 1117.2001 1514.7001 1118.1000 ;
	    RECT 1516.2001 1117.2001 1517.4000 1118.4000 ;
	    RECT 1510.5000 1116.3000 1511.4000 1117.2001 ;
	    RECT 1518.6000 1116.3000 1519.8000 1117.5000 ;
	    RECT 1503.3000 1115.4000 1505.4000 1116.3000 ;
	    RECT 1503.3000 1113.3000 1505.1000 1115.4000 ;
	    RECT 1507.8000 1113.3000 1509.0000 1116.3000 ;
	    RECT 1510.2001 1113.3000 1511.4000 1116.3000 ;
	    RECT 1512.6000 1113.3000 1514.1000 1116.3000 ;
	    RECT 1516.8000 1115.4000 1519.8000 1116.3000 ;
	    RECT 1516.8000 1113.3000 1518.0000 1115.4000 ;
	    RECT 1521.0000 1113.3000 1522.2001 1119.3000 ;
	    RECT 1523.4000 1113.3000 1524.6000 1120.5000 ;
	    RECT 1542.6000 1120.2001 1543.8000 1120.5000 ;
	    RECT 1545.0000 1119.3000 1546.2001 1123.5000 ;
	    RECT 1542.6000 1113.3000 1543.8000 1119.3000 ;
	    RECT 1545.0000 1118.4000 1547.7001 1119.3000 ;
	    RECT 1546.5000 1113.3000 1547.7001 1118.4000 ;
	    RECT 1.2000 1110.6000 1569.0000 1112.4000 ;
	    RECT 124.2000 1100.7001 125.4000 1109.7001 ;
	    RECT 129.0000 1103.7001 130.2000 1109.7001 ;
	    RECT 133.8000 1104.9000 135.0000 1109.7001 ;
	    RECT 136.2000 1105.5000 137.4000 1109.7001 ;
	    RECT 138.6000 1105.5000 139.8000 1109.7001 ;
	    RECT 141.0000 1105.5000 142.2000 1109.7001 ;
	    RECT 143.4000 1106.7001 144.6000 1109.7001 ;
	    RECT 145.8000 1105.5000 147.0000 1109.7001 ;
	    RECT 148.2000 1106.7001 149.4000 1109.7001 ;
	    RECT 150.6000 1105.5000 151.8000 1109.7001 ;
	    RECT 153.0000 1105.5000 154.2000 1109.7001 ;
	    RECT 155.4000 1105.5000 156.6000 1109.7001 ;
	    RECT 157.8000 1105.5000 159.0000 1109.7001 ;
	    RECT 131.1000 1103.7001 135.0000 1104.9000 ;
	    RECT 160.2000 1104.9000 161.4000 1109.7001 ;
	    RECT 140.1000 1103.7001 147.0000 1104.6000 ;
	    RECT 131.1000 1102.8000 132.3000 1103.7001 ;
	    RECT 127.8000 1101.6000 132.3000 1102.8000 ;
	    RECT 124.2000 1099.5000 137.4000 1100.7001 ;
	    RECT 140.1000 1100.1000 141.3000 1103.7001 ;
	    RECT 145.8000 1103.4000 147.0000 1103.7001 ;
	    RECT 148.2000 1103.4000 149.4000 1104.6000 ;
	    RECT 150.3000 1103.4000 150.6000 1104.6000 ;
	    RECT 155.1000 1103.4000 156.6000 1104.6000 ;
	    RECT 160.2000 1103.7001 163.8000 1104.9000 ;
	    RECT 165.0000 1103.7001 166.2000 1109.7001 ;
	    RECT 143.4000 1102.5000 144.6000 1102.8000 ;
	    RECT 145.8000 1102.2001 147.0000 1102.5000 ;
	    RECT 143.4000 1100.4000 144.6000 1101.6000 ;
	    RECT 145.8000 1101.3000 152.4000 1102.2001 ;
	    RECT 151.2000 1101.0000 152.4000 1101.3000 ;
	    RECT 124.2000 1091.1000 125.4000 1099.5000 ;
	    RECT 138.3000 1098.9000 141.3000 1100.1000 ;
	    RECT 147.0000 1098.9000 151.8000 1100.1000 ;
	    RECT 155.4000 1099.2001 156.6000 1103.4000 ;
	    RECT 162.6000 1102.8000 163.8000 1103.7001 ;
	    RECT 162.6000 1101.9000 165.3000 1102.8000 ;
	    RECT 164.1000 1100.1000 165.3000 1101.9000 ;
	    RECT 169.8000 1101.9000 171.0000 1109.7001 ;
	    RECT 172.2000 1104.0000 173.4000 1109.7001 ;
	    RECT 174.6000 1106.7001 175.8000 1109.7001 ;
	    RECT 172.2000 1102.8000 173.7000 1104.0000 ;
	    RECT 169.8000 1101.0000 171.6000 1101.9000 ;
	    RECT 164.1000 1098.9000 169.8000 1100.1000 ;
	    RECT 126.3000 1098.0000 127.5000 1098.3000 ;
	    RECT 126.3000 1097.1000 132.9000 1098.0000 ;
	    RECT 133.8000 1097.4000 135.0000 1098.6000 ;
	    RECT 160.2000 1098.0000 161.4000 1098.9000 ;
	    RECT 170.7000 1098.0000 171.6000 1101.0000 ;
	    RECT 135.9000 1097.1000 161.4000 1098.0000 ;
	    RECT 170.4000 1097.1000 171.6000 1098.0000 ;
	    RECT 168.3000 1096.2001 169.5000 1096.5000 ;
	    RECT 129.0000 1094.4000 130.2000 1095.6000 ;
	    RECT 131.1000 1095.3000 169.5000 1096.2001 ;
	    RECT 134.1000 1095.0000 135.3000 1095.3000 ;
	    RECT 170.4000 1094.4000 171.3000 1097.1000 ;
	    RECT 172.5000 1096.2001 173.7000 1102.8000 ;
	    RECT 189.0000 1102.5000 190.2000 1109.7001 ;
	    RECT 191.4000 1106.7001 192.6000 1109.7001 ;
	    RECT 210.6000 1106.7001 211.8000 1109.7001 ;
	    RECT 191.4000 1105.5000 192.6000 1105.8000 ;
	    RECT 210.6000 1105.5000 211.8000 1105.8000 ;
	    RECT 191.4000 1104.4501 192.6000 1104.6000 ;
	    RECT 196.2000 1104.4501 197.4000 1104.6000 ;
	    RECT 191.4000 1103.5500 197.4000 1104.4501 ;
	    RECT 191.4000 1103.4000 192.6000 1103.5500 ;
	    RECT 196.2000 1103.4000 197.4000 1103.5500 ;
	    RECT 210.6000 1103.4000 211.8000 1104.6000 ;
	    RECT 213.0000 1102.5000 214.2000 1109.7001 ;
	    RECT 244.2000 1104.0000 245.4000 1109.7001 ;
	    RECT 246.6000 1104.9000 247.8000 1109.7001 ;
	    RECT 249.0000 1108.8000 255.0000 1109.7001 ;
	    RECT 249.0000 1104.0000 250.2000 1108.8000 ;
	    RECT 244.2000 1103.7001 250.2000 1104.0000 ;
	    RECT 251.4000 1103.7001 252.6000 1107.9000 ;
	    RECT 253.8000 1103.7001 255.0000 1108.8000 ;
	    RECT 273.0000 1106.7001 274.2000 1109.7001 ;
	    RECT 275.4000 1106.7001 276.6000 1109.7001 ;
	    RECT 277.8000 1106.7001 279.0000 1109.7001 ;
	    RECT 244.5000 1103.1000 249.9000 1103.7001 ;
	    RECT 189.0000 1101.4501 190.2000 1101.6000 ;
	    RECT 196.2000 1101.4501 197.4000 1101.6000 ;
	    RECT 189.0000 1100.5500 197.4000 1101.4501 ;
	    RECT 189.0000 1100.4000 190.2000 1100.5500 ;
	    RECT 196.2000 1100.4000 197.4000 1100.5500 ;
	    RECT 213.0000 1101.4501 214.2000 1101.6000 ;
	    RECT 225.0000 1101.4501 226.2000 1101.6000 ;
	    RECT 213.0000 1100.5500 226.2000 1101.4501 ;
	    RECT 213.0000 1100.4000 214.2000 1100.5500 ;
	    RECT 225.0000 1100.4000 226.2000 1100.5500 ;
	    RECT 239.4000 1101.4501 240.6000 1101.6000 ;
	    RECT 244.2000 1101.4501 245.4000 1101.6000 ;
	    RECT 239.4000 1100.5500 245.4000 1101.4501 ;
	    RECT 246.3000 1100.7001 246.6000 1102.2001 ;
	    RECT 251.7000 1101.6000 252.6000 1103.7001 ;
	    RECT 275.4000 1102.5000 276.3000 1106.7001 ;
	    RECT 277.8000 1105.5000 279.0000 1105.8000 ;
	    RECT 297.9000 1104.6000 299.1000 1109.7001 ;
	    RECT 277.8000 1103.4000 279.0000 1104.6000 ;
	    RECT 297.9000 1103.7001 300.6000 1104.6000 ;
	    RECT 301.8000 1103.7001 303.0000 1109.7001 ;
	    RECT 333.0000 1104.0000 334.2000 1109.7001 ;
	    RECT 335.4000 1104.9000 336.6000 1109.7001 ;
	    RECT 337.8000 1108.8000 343.8000 1109.7001 ;
	    RECT 337.8000 1104.0000 339.0000 1108.8000 ;
	    RECT 333.0000 1103.7001 339.0000 1104.0000 ;
	    RECT 340.2000 1103.7001 341.4000 1107.9000 ;
	    RECT 342.6000 1103.7001 343.8000 1108.8000 ;
	    RECT 239.4000 1100.4000 240.6000 1100.5500 ;
	    RECT 244.2000 1100.4000 245.4000 1100.5500 ;
	    RECT 249.0000 1100.4000 250.2000 1101.6000 ;
	    RECT 251.1000 1100.7001 252.6000 1101.6000 ;
	    RECT 253.8000 1101.4501 255.0000 1101.6000 ;
	    RECT 263.4000 1101.4501 264.6000 1101.6000 ;
	    RECT 253.8000 1100.5500 264.6000 1101.4501 ;
	    RECT 253.8000 1100.4000 255.0000 1100.5500 ;
	    RECT 263.4000 1100.4000 264.6000 1100.5500 ;
	    RECT 275.4000 1101.4501 276.6000 1101.6000 ;
	    RECT 294.6000 1101.4501 295.8000 1101.6000 ;
	    RECT 275.4000 1100.5500 295.8000 1101.4501 ;
	    RECT 275.4000 1100.4000 276.6000 1100.5500 ;
	    RECT 294.6000 1100.4000 295.8000 1100.5500 ;
	    RECT 246.6000 1099.5000 247.8000 1099.8000 ;
	    RECT 251.4000 1099.5000 252.6000 1099.8000 ;
	    RECT 299.4000 1099.5000 300.6000 1103.7001 ;
	    RECT 333.3000 1103.1000 338.7000 1103.7001 ;
	    RECT 301.8000 1102.5000 303.0000 1102.8000 ;
	    RECT 301.8000 1100.4000 303.0000 1101.6000 ;
	    RECT 330.6000 1101.4501 331.8000 1101.6000 ;
	    RECT 333.0000 1101.4501 334.2000 1101.6000 ;
	    RECT 330.6000 1100.5500 334.2000 1101.4501 ;
	    RECT 335.1000 1100.7001 335.4000 1102.2001 ;
	    RECT 340.5000 1101.6000 341.4000 1103.7001 ;
	    RECT 354.6000 1102.5000 355.8000 1109.7001 ;
	    RECT 357.0000 1106.7001 358.2000 1109.7001 ;
	    RECT 357.0000 1105.5000 358.2000 1105.8000 ;
	    RECT 357.0000 1103.4000 358.2000 1104.6000 ;
	    RECT 369.0000 1102.5000 370.2000 1109.7001 ;
	    RECT 371.4000 1106.7001 372.6000 1109.7001 ;
	    RECT 385.8000 1106.7001 387.0000 1109.7001 ;
	    RECT 371.4000 1105.5000 372.6000 1105.8000 ;
	    RECT 385.8000 1105.5000 387.0000 1105.8000 ;
	    RECT 371.4000 1104.4501 372.6000 1104.6000 ;
	    RECT 376.2000 1104.4501 377.4000 1104.6000 ;
	    RECT 371.4000 1103.5500 377.4000 1104.4501 ;
	    RECT 371.4000 1103.4000 372.6000 1103.5500 ;
	    RECT 376.2000 1103.4000 377.4000 1103.5500 ;
	    RECT 385.8000 1103.4000 387.0000 1104.6000 ;
	    RECT 388.2000 1102.5000 389.4000 1109.7001 ;
	    RECT 412.2000 1104.0000 413.4000 1109.7001 ;
	    RECT 414.6000 1104.9000 415.8000 1109.7001 ;
	    RECT 417.0000 1104.0000 418.2000 1109.7001 ;
	    RECT 412.2000 1103.7001 418.2000 1104.0000 ;
	    RECT 419.4000 1103.7001 420.6000 1109.7001 ;
	    RECT 412.5000 1103.1000 417.9000 1103.7001 ;
	    RECT 419.4000 1102.5000 420.3000 1103.7001 ;
	    RECT 441.0000 1102.5000 442.2000 1109.7001 ;
	    RECT 443.4000 1106.7001 444.6000 1109.7001 ;
	    RECT 443.4000 1105.5000 444.6000 1105.8000 ;
	    RECT 443.4000 1104.4501 444.6000 1104.6000 ;
	    RECT 445.8000 1104.4501 447.0000 1104.6000 ;
	    RECT 443.4000 1103.5500 447.0000 1104.4501 ;
	    RECT 443.4000 1103.4000 444.6000 1103.5500 ;
	    RECT 445.8000 1103.4000 447.0000 1103.5500 ;
	    RECT 330.6000 1100.4000 331.8000 1100.5500 ;
	    RECT 333.0000 1100.4000 334.2000 1100.5500 ;
	    RECT 337.8000 1100.4000 339.0000 1101.6000 ;
	    RECT 339.9000 1100.7001 341.4000 1101.6000 ;
	    RECT 342.6000 1101.4501 343.8000 1101.6000 ;
	    RECT 354.6000 1101.4501 355.8000 1101.6000 ;
	    RECT 342.6000 1100.5500 355.8000 1101.4501 ;
	    RECT 342.6000 1100.4000 343.8000 1100.5500 ;
	    RECT 354.6000 1100.4000 355.8000 1100.5500 ;
	    RECT 357.0000 1101.4501 358.2000 1101.6000 ;
	    RECT 369.0000 1101.4501 370.2000 1101.6000 ;
	    RECT 357.0000 1100.5500 370.2000 1101.4501 ;
	    RECT 357.0000 1100.4000 358.2000 1100.5500 ;
	    RECT 369.0000 1100.4000 370.2000 1100.5500 ;
	    RECT 388.2000 1100.4000 389.4000 1101.6000 ;
	    RECT 390.6000 1101.4501 391.8000 1101.6000 ;
	    RECT 412.2000 1101.4501 413.4000 1101.6000 ;
	    RECT 390.6000 1100.5500 413.4000 1101.4501 ;
	    RECT 414.3000 1100.7001 414.6000 1102.2001 ;
	    RECT 390.6000 1100.4000 391.8000 1100.5500 ;
	    RECT 412.2000 1100.4000 413.4000 1100.5500 ;
	    RECT 416.7000 1100.4000 418.5000 1101.6000 ;
	    RECT 419.4000 1101.4501 420.6000 1101.6000 ;
	    RECT 438.6000 1101.4501 439.8000 1101.6000 ;
	    RECT 419.4000 1100.5500 439.8000 1101.4501 ;
	    RECT 419.4000 1100.4000 420.6000 1100.5500 ;
	    RECT 438.6000 1100.4000 439.8000 1100.5500 ;
	    RECT 441.0000 1101.4501 442.2000 1101.6000 ;
	    RECT 503.4000 1101.4501 504.6000 1101.6000 ;
	    RECT 441.0000 1100.5500 504.6000 1101.4501 ;
	    RECT 441.0000 1100.4000 442.2000 1100.5500 ;
	    RECT 503.4000 1100.4000 504.6000 1100.5500 ;
	    RECT 568.2000 1100.7001 569.4000 1109.7001 ;
	    RECT 573.0000 1103.7001 574.2000 1109.7001 ;
	    RECT 577.8000 1104.9000 579.0000 1109.7001 ;
	    RECT 580.2000 1105.5000 581.4000 1109.7001 ;
	    RECT 582.6000 1105.5000 583.8000 1109.7001 ;
	    RECT 585.0000 1105.5000 586.2000 1109.7001 ;
	    RECT 587.4000 1106.7001 588.6000 1109.7001 ;
	    RECT 589.8000 1105.5000 591.0000 1109.7001 ;
	    RECT 592.2000 1106.7001 593.4000 1109.7001 ;
	    RECT 594.6000 1105.5000 595.8000 1109.7001 ;
	    RECT 597.0000 1105.5000 598.2000 1109.7001 ;
	    RECT 599.4000 1105.5000 600.6000 1109.7001 ;
	    RECT 601.8000 1105.5000 603.0000 1109.7001 ;
	    RECT 575.1000 1103.7001 579.0000 1104.9000 ;
	    RECT 604.2000 1104.9000 605.4000 1109.7001 ;
	    RECT 584.1000 1103.7001 591.0000 1104.6000 ;
	    RECT 575.1000 1102.8000 576.3000 1103.7001 ;
	    RECT 571.8000 1101.6000 576.3000 1102.8000 ;
	    RECT 335.4000 1099.5000 336.6000 1099.8000 ;
	    RECT 340.2000 1099.5000 341.4000 1099.8000 ;
	    RECT 414.6000 1099.5000 415.8000 1099.8000 ;
	    RECT 138.6000 1094.1000 139.8000 1094.4000 ;
	    RECT 131.7000 1093.5000 139.8000 1094.1000 ;
	    RECT 130.5000 1093.2001 139.8000 1093.5000 ;
	    RECT 141.3000 1093.5000 154.2000 1094.4000 ;
	    RECT 126.6000 1092.0000 129.0000 1093.2001 ;
	    RECT 130.5000 1092.3000 132.6000 1093.2001 ;
	    RECT 141.3000 1092.3000 142.2000 1093.5000 ;
	    RECT 153.0000 1093.2001 154.2000 1093.5000 ;
	    RECT 157.8000 1093.5000 171.3000 1094.4000 ;
	    RECT 172.2000 1095.0000 173.7000 1096.2001 ;
	    RECT 172.2000 1093.5000 173.4000 1095.0000 ;
	    RECT 157.8000 1093.2001 159.0000 1093.5000 ;
	    RECT 128.1000 1091.4000 129.0000 1092.0000 ;
	    RECT 133.5000 1091.4000 142.2000 1092.3000 ;
	    RECT 143.1000 1091.4000 147.0000 1092.6000 ;
	    RECT 124.2000 1090.2001 127.2000 1091.1000 ;
	    RECT 128.1000 1090.2001 134.4000 1091.4000 ;
	    RECT 126.3000 1089.3000 127.2000 1090.2001 ;
	    RECT 124.2000 1083.3000 125.4000 1089.3000 ;
	    RECT 126.3000 1088.4000 127.8000 1089.3000 ;
	    RECT 126.6000 1083.3000 127.8000 1088.4000 ;
	    RECT 129.0000 1082.4000 130.2000 1089.3000 ;
	    RECT 131.4000 1083.3000 132.6000 1090.2001 ;
	    RECT 133.8000 1083.3000 135.0000 1089.3000 ;
	    RECT 136.2000 1083.3000 137.4000 1087.5000 ;
	    RECT 138.6000 1083.3000 139.8000 1087.5000 ;
	    RECT 141.0000 1083.3000 142.2000 1090.5000 ;
	    RECT 143.4000 1083.3000 144.6000 1089.3000 ;
	    RECT 145.8000 1083.3000 147.0000 1090.5000 ;
	    RECT 148.2000 1083.3000 149.4000 1089.3000 ;
	    RECT 150.6000 1083.3000 151.8000 1092.6000 ;
	    RECT 162.6000 1091.4000 166.5000 1092.6000 ;
	    RECT 155.4000 1090.2001 161.7000 1091.4000 ;
	    RECT 153.0000 1083.3000 154.2000 1087.5000 ;
	    RECT 155.4000 1083.3000 156.6000 1087.5000 ;
	    RECT 157.8000 1083.3000 159.0000 1087.5000 ;
	    RECT 160.2000 1083.3000 161.4000 1089.3000 ;
	    RECT 162.6000 1083.3000 163.8000 1091.4000 ;
	    RECT 170.4000 1091.1000 171.3000 1093.5000 ;
	    RECT 172.2000 1091.4000 173.4000 1092.6000 ;
	    RECT 167.4000 1090.2001 171.3000 1091.1000 ;
	    RECT 165.0000 1083.3000 166.2000 1089.3000 ;
	    RECT 167.4000 1083.3000 168.6000 1090.2001 ;
	    RECT 169.8000 1083.3000 171.0000 1089.3000 ;
	    RECT 172.2000 1083.3000 173.4000 1090.5000 ;
	    RECT 174.6000 1083.3000 175.8000 1089.3000 ;
	    RECT 189.0000 1083.3000 190.2000 1099.5000 ;
	    RECT 191.4000 1083.3000 192.6000 1089.3000 ;
	    RECT 210.6000 1083.3000 211.8000 1089.3000 ;
	    RECT 213.0000 1083.3000 214.2000 1099.5000 ;
	    RECT 220.2000 1098.4501 221.4000 1098.6000 ;
	    RECT 246.6000 1098.4501 247.8000 1098.6000 ;
	    RECT 220.2000 1097.5500 247.8000 1098.4501 ;
	    RECT 220.2000 1097.4000 221.4000 1097.5500 ;
	    RECT 246.6000 1097.4000 247.8000 1097.5500 ;
	    RECT 249.0000 1095.3000 249.9000 1099.5000 ;
	    RECT 253.8000 1099.2001 255.0000 1099.5000 ;
	    RECT 251.4000 1097.4000 252.6000 1098.6000 ;
	    RECT 273.0000 1097.4000 274.2000 1098.6000 ;
	    RECT 273.0000 1096.2001 274.2000 1096.5000 ;
	    RECT 275.4000 1095.3000 276.3000 1099.5000 ;
	    RECT 299.4000 1097.4000 300.6000 1098.6000 ;
	    RECT 301.8000 1098.4501 303.0000 1098.6000 ;
	    RECT 335.4000 1098.4501 336.6000 1098.6000 ;
	    RECT 301.8000 1097.5500 336.6000 1098.4501 ;
	    RECT 301.8000 1097.4000 303.0000 1097.5500 ;
	    RECT 335.4000 1097.4000 336.6000 1097.5500 ;
	    RECT 294.6000 1095.4501 295.8000 1095.6000 ;
	    RECT 297.0000 1095.4501 298.2000 1095.6000 ;
	    RECT 244.2000 1083.3000 245.4000 1095.3000 ;
	    RECT 248.1000 1083.3000 251.1000 1095.3000 ;
	    RECT 253.8000 1083.3000 255.0000 1095.3000 ;
	    RECT 273.9000 1094.1000 276.6000 1095.3000 ;
	    RECT 256.2000 1092.4501 257.4000 1092.6000 ;
	    RECT 270.6000 1092.4501 271.8000 1092.6000 ;
	    RECT 256.2000 1091.5500 271.8000 1092.4501 ;
	    RECT 256.2000 1091.4000 257.4000 1091.5500 ;
	    RECT 270.6000 1091.4000 271.8000 1091.5500 ;
	    RECT 273.9000 1083.3000 275.1000 1094.1000 ;
	    RECT 277.8000 1083.3000 279.0000 1095.3000 ;
	    RECT 294.6000 1094.5500 298.2000 1095.4501 ;
	    RECT 294.6000 1094.4000 295.8000 1094.5500 ;
	    RECT 297.0000 1094.4000 298.2000 1094.5500 ;
	    RECT 297.0000 1093.2001 298.2000 1093.5000 ;
	    RECT 297.0000 1083.3000 298.2000 1089.3000 ;
	    RECT 299.4000 1083.3000 300.6000 1096.5000 ;
	    RECT 337.8000 1095.3000 338.7000 1099.5000 ;
	    RECT 342.6000 1099.2001 343.8000 1099.5000 ;
	    RECT 340.2000 1097.4000 341.4000 1098.6000 ;
	    RECT 301.8000 1083.3000 303.0000 1089.3000 ;
	    RECT 306.6000 1086.4501 307.8000 1086.6000 ;
	    RECT 313.8000 1086.4501 315.0000 1086.6000 ;
	    RECT 306.6000 1085.5500 315.0000 1086.4501 ;
	    RECT 306.6000 1085.4000 307.8000 1085.5500 ;
	    RECT 313.8000 1085.4000 315.0000 1085.5500 ;
	    RECT 333.0000 1083.3000 334.2000 1095.3000 ;
	    RECT 336.9000 1083.3000 339.9000 1095.3000 ;
	    RECT 342.6000 1083.3000 343.8000 1095.3000 ;
	    RECT 354.6000 1083.3000 355.8000 1099.5000 ;
	    RECT 357.0000 1083.3000 358.2000 1089.3000 ;
	    RECT 369.0000 1083.3000 370.2000 1099.5000 ;
	    RECT 371.4000 1083.3000 372.6000 1089.3000 ;
	    RECT 385.8000 1083.3000 387.0000 1089.3000 ;
	    RECT 388.2000 1083.3000 389.4000 1099.5000 ;
	    RECT 400.2000 1098.4501 401.4000 1098.6000 ;
	    RECT 414.6000 1098.4501 415.8000 1098.6000 ;
	    RECT 400.2000 1097.5500 415.8000 1098.4501 ;
	    RECT 400.2000 1097.4000 401.4000 1097.5500 ;
	    RECT 414.6000 1097.4000 415.8000 1097.5500 ;
	    RECT 416.7000 1095.3000 417.6000 1100.4000 ;
	    RECT 568.2000 1099.5000 581.4000 1100.7001 ;
	    RECT 584.1000 1100.1000 585.3000 1103.7001 ;
	    RECT 589.8000 1103.4000 591.0000 1103.7001 ;
	    RECT 592.2000 1103.4000 593.4000 1104.6000 ;
	    RECT 594.3000 1103.4000 594.6000 1104.6000 ;
	    RECT 599.1000 1103.4000 600.6000 1104.6000 ;
	    RECT 604.2000 1103.7001 607.8000 1104.9000 ;
	    RECT 609.0000 1103.7001 610.2000 1109.7001 ;
	    RECT 587.4000 1102.5000 588.6000 1102.8000 ;
	    RECT 589.8000 1102.2001 591.0000 1102.5000 ;
	    RECT 587.4000 1100.4000 588.6000 1101.6000 ;
	    RECT 589.8000 1101.3000 596.4000 1102.2001 ;
	    RECT 595.2000 1101.0000 596.4000 1101.3000 ;
	    RECT 412.2000 1083.3000 413.4000 1095.3000 ;
	    RECT 416.1000 1094.4000 417.6000 1095.3000 ;
	    RECT 419.4000 1094.4000 420.6000 1095.6000 ;
	    RECT 416.1000 1083.3000 417.3000 1094.4000 ;
	    RECT 418.5000 1092.6000 419.4000 1093.5000 ;
	    RECT 418.2000 1091.4000 419.4000 1092.6000 ;
	    RECT 418.5000 1083.3000 419.7000 1089.3000 ;
	    RECT 441.0000 1083.3000 442.2000 1099.5000 ;
	    RECT 568.2000 1091.1000 569.4000 1099.5000 ;
	    RECT 582.3000 1098.9000 585.3000 1100.1000 ;
	    RECT 591.0000 1098.9000 595.8000 1100.1000 ;
	    RECT 599.4000 1099.2001 600.6000 1103.4000 ;
	    RECT 606.6000 1102.8000 607.8000 1103.7001 ;
	    RECT 606.6000 1101.9000 609.3000 1102.8000 ;
	    RECT 608.1000 1100.1000 609.3000 1101.9000 ;
	    RECT 613.8000 1101.9000 615.0000 1109.7001 ;
	    RECT 616.2000 1104.0000 617.4000 1109.7001 ;
	    RECT 618.6000 1106.7001 619.8000 1109.7001 ;
	    RECT 638.7000 1104.6000 639.9000 1109.7001 ;
	    RECT 616.2000 1102.8000 617.7000 1104.0000 ;
	    RECT 638.7000 1103.7001 641.4000 1104.6000 ;
	    RECT 642.6000 1103.7001 643.8000 1109.7001 ;
	    RECT 673.8000 1103.7001 675.0000 1109.7001 ;
	    RECT 676.2000 1104.0000 677.4000 1109.7001 ;
	    RECT 678.6000 1104.9000 679.8000 1109.7001 ;
	    RECT 681.0000 1104.0000 682.2000 1109.7001 ;
	    RECT 695.4000 1106.7001 696.6000 1109.7001 ;
	    RECT 695.4000 1105.5000 696.6000 1105.8000 ;
	    RECT 676.2000 1103.7001 682.2000 1104.0000 ;
	    RECT 683.4000 1104.4501 684.6000 1104.6000 ;
	    RECT 695.4000 1104.4501 696.6000 1104.6000 ;
	    RECT 613.8000 1101.0000 615.6000 1101.9000 ;
	    RECT 608.1000 1098.9000 613.8000 1100.1000 ;
	    RECT 570.3000 1098.0000 571.5000 1098.3000 ;
	    RECT 570.3000 1097.1000 576.9000 1098.0000 ;
	    RECT 577.8000 1097.4000 579.0000 1098.6000 ;
	    RECT 604.2000 1098.0000 605.4000 1098.9000 ;
	    RECT 614.7000 1098.0000 615.6000 1101.0000 ;
	    RECT 579.9000 1097.1000 605.4000 1098.0000 ;
	    RECT 614.4000 1097.1000 615.6000 1098.0000 ;
	    RECT 612.3000 1096.2001 613.5000 1096.5000 ;
	    RECT 573.0000 1094.4000 574.2000 1095.6000 ;
	    RECT 575.1000 1095.3000 613.5000 1096.2001 ;
	    RECT 578.1000 1095.0000 579.3000 1095.3000 ;
	    RECT 614.4000 1094.4000 615.3000 1097.1000 ;
	    RECT 616.5000 1096.2001 617.7000 1102.8000 ;
	    RECT 640.2000 1099.5000 641.4000 1103.7001 ;
	    RECT 642.6000 1102.5000 643.8000 1102.8000 ;
	    RECT 674.1000 1102.5000 675.0000 1103.7001 ;
	    RECT 676.5000 1103.1000 681.9000 1103.7001 ;
	    RECT 683.4000 1103.5500 696.6000 1104.4501 ;
	    RECT 683.4000 1103.4000 684.6000 1103.5500 ;
	    RECT 695.4000 1103.4000 696.6000 1103.5500 ;
	    RECT 697.8000 1102.5000 699.0000 1109.7001 ;
	    RECT 738.6000 1103.7001 739.8000 1109.7001 ;
	    RECT 741.0000 1104.6000 742.5000 1109.7001 ;
	    RECT 745.2000 1104.3000 747.6000 1109.7001 ;
	    RECT 750.3000 1104.6000 751.8000 1109.7001 ;
	    RECT 738.6000 1102.8000 742.2000 1103.7001 ;
	    RECT 741.0000 1102.5000 742.2000 1102.8000 ;
	    RECT 743.1000 1102.2001 744.3000 1103.4000 ;
	    RECT 642.6000 1100.4000 643.8000 1101.6000 ;
	    RECT 652.2000 1101.4501 653.4000 1101.6000 ;
	    RECT 673.8000 1101.4501 675.0000 1101.6000 ;
	    RECT 652.2000 1100.5500 675.0000 1101.4501 ;
	    RECT 652.2000 1100.4000 653.4000 1100.5500 ;
	    RECT 673.8000 1100.4000 675.0000 1100.5500 ;
	    RECT 675.9000 1100.4000 677.7000 1101.6000 ;
	    RECT 679.8000 1100.7001 680.1000 1102.2001 ;
	    RECT 743.1000 1101.6000 744.0000 1102.2001 ;
	    RECT 681.0000 1100.4000 682.2000 1101.6000 ;
	    RECT 697.8000 1101.4501 699.0000 1101.6000 ;
	    RECT 683.5500 1100.5500 699.0000 1101.4501 ;
	    RECT 640.2000 1098.4501 641.4000 1098.6000 ;
	    RECT 640.2000 1097.5500 674.8500 1098.4501 ;
	    RECT 640.2000 1097.4000 641.4000 1097.5500 ;
	    RECT 582.6000 1094.1000 583.8000 1094.4000 ;
	    RECT 575.7000 1093.5000 583.8000 1094.1000 ;
	    RECT 574.5000 1093.2001 583.8000 1093.5000 ;
	    RECT 585.3000 1093.5000 598.2000 1094.4000 ;
	    RECT 570.6000 1092.0000 573.0000 1093.2001 ;
	    RECT 574.5000 1092.3000 576.6000 1093.2001 ;
	    RECT 585.3000 1092.3000 586.2000 1093.5000 ;
	    RECT 597.0000 1093.2001 598.2000 1093.5000 ;
	    RECT 601.8000 1093.5000 615.3000 1094.4000 ;
	    RECT 616.2000 1095.0000 617.7000 1096.2001 ;
	    RECT 618.6000 1095.4501 619.8000 1095.6000 ;
	    RECT 637.8000 1095.4501 639.0000 1095.6000 ;
	    RECT 616.2000 1093.5000 617.4000 1095.0000 ;
	    RECT 618.6000 1094.5500 639.0000 1095.4501 ;
	    RECT 618.6000 1094.4000 619.8000 1094.5500 ;
	    RECT 637.8000 1094.4000 639.0000 1094.5500 ;
	    RECT 601.8000 1093.2001 603.0000 1093.5000 ;
	    RECT 572.1000 1091.4000 573.0000 1092.0000 ;
	    RECT 577.5000 1091.4000 586.2000 1092.3000 ;
	    RECT 587.1000 1091.4000 591.0000 1092.6000 ;
	    RECT 568.2000 1090.2001 571.2000 1091.1000 ;
	    RECT 572.1000 1090.2001 578.4000 1091.4000 ;
	    RECT 570.3000 1089.3000 571.2000 1090.2001 ;
	    RECT 443.4000 1083.3000 444.6000 1089.3000 ;
	    RECT 568.2000 1083.3000 569.4000 1089.3000 ;
	    RECT 570.3000 1088.4000 571.8000 1089.3000 ;
	    RECT 570.6000 1083.3000 571.8000 1088.4000 ;
	    RECT 573.0000 1082.4000 574.2000 1089.3000 ;
	    RECT 575.4000 1083.3000 576.6000 1090.2001 ;
	    RECT 577.8000 1083.3000 579.0000 1089.3000 ;
	    RECT 580.2000 1083.3000 581.4000 1087.5000 ;
	    RECT 582.6000 1083.3000 583.8000 1087.5000 ;
	    RECT 585.0000 1083.3000 586.2000 1090.5000 ;
	    RECT 587.4000 1083.3000 588.6000 1089.3000 ;
	    RECT 589.8000 1083.3000 591.0000 1090.5000 ;
	    RECT 592.2000 1083.3000 593.4000 1089.3000 ;
	    RECT 594.6000 1083.3000 595.8000 1092.6000 ;
	    RECT 606.6000 1091.4000 610.5000 1092.6000 ;
	    RECT 599.4000 1090.2001 605.7000 1091.4000 ;
	    RECT 597.0000 1083.3000 598.2000 1087.5000 ;
	    RECT 599.4000 1083.3000 600.6000 1087.5000 ;
	    RECT 601.8000 1083.3000 603.0000 1087.5000 ;
	    RECT 604.2000 1083.3000 605.4000 1089.3000 ;
	    RECT 606.6000 1083.3000 607.8000 1091.4000 ;
	    RECT 614.4000 1091.1000 615.3000 1093.5000 ;
	    RECT 637.8000 1093.2001 639.0000 1093.5000 ;
	    RECT 616.2000 1091.4000 617.4000 1092.6000 ;
	    RECT 611.4000 1090.2001 615.3000 1091.1000 ;
	    RECT 609.0000 1083.3000 610.2000 1089.3000 ;
	    RECT 611.4000 1083.3000 612.6000 1090.2001 ;
	    RECT 613.8000 1083.3000 615.0000 1089.3000 ;
	    RECT 616.2000 1083.3000 617.4000 1090.5000 ;
	    RECT 618.6000 1083.3000 619.8000 1089.3000 ;
	    RECT 637.8000 1083.3000 639.0000 1089.3000 ;
	    RECT 640.2000 1083.3000 641.4000 1096.5000 ;
	    RECT 673.9500 1095.6000 674.8500 1097.5500 ;
	    RECT 673.8000 1094.4000 675.0000 1095.6000 ;
	    RECT 676.8000 1095.3000 677.7000 1100.4000 ;
	    RECT 678.6000 1099.5000 679.8000 1099.8000 ;
	    RECT 678.6000 1098.4501 679.8000 1098.6000 ;
	    RECT 683.5500 1098.4501 684.4500 1100.5500 ;
	    RECT 697.8000 1100.4000 699.0000 1100.5500 ;
	    RECT 707.4000 1101.4501 708.6000 1101.6000 ;
	    RECT 738.6000 1101.4501 739.8000 1101.6000 ;
	    RECT 707.4000 1100.5500 739.8000 1101.4501 ;
	    RECT 707.4000 1100.4000 708.6000 1100.5500 ;
	    RECT 738.6000 1100.4000 739.8000 1100.5500 ;
	    RECT 740.7000 1100.4000 741.0000 1101.6000 ;
	    RECT 742.8000 1100.4000 744.0000 1101.6000 ;
	    RECT 745.2000 1101.3000 746.1000 1104.3000 ;
	    RECT 753.0000 1103.7001 754.2000 1109.7001 ;
	    RECT 773.1000 1104.6000 774.3000 1109.7001 ;
	    RECT 773.1000 1103.7001 775.8000 1104.6000 ;
	    RECT 777.0000 1103.7001 778.2000 1109.7001 ;
	    RECT 791.4000 1106.7001 792.6000 1109.7001 ;
	    RECT 791.4000 1105.5000 792.6000 1105.8000 ;
	    RECT 747.0000 1102.2001 749.4000 1103.4000 ;
	    RECT 750.3000 1102.8000 754.2000 1103.7001 ;
	    RECT 750.3000 1102.5000 751.5000 1102.8000 ;
	    RECT 751.8000 1101.3000 752.1000 1101.6000 ;
	    RECT 745.2000 1100.4000 746.7000 1101.3000 ;
	    RECT 750.9000 1101.0000 752.1000 1101.3000 ;
	    RECT 745.8000 1099.5000 746.7000 1100.4000 ;
	    RECT 747.6000 1100.4000 752.1000 1101.0000 ;
	    RECT 753.0000 1100.4000 754.2000 1101.6000 ;
	    RECT 747.6000 1100.1000 751.8000 1100.4000 ;
	    RECT 747.6000 1099.8000 748.8000 1100.1000 ;
	    RECT 774.6000 1099.5000 775.8000 1103.7001 ;
	    RECT 791.4000 1103.4000 792.6000 1104.6000 ;
	    RECT 777.0000 1102.5000 778.2000 1102.8000 ;
	    RECT 793.8000 1102.5000 795.0000 1109.7001 ;
	    RECT 822.6000 1108.8000 828.6000 1109.7001 ;
	    RECT 822.6000 1103.7001 823.8000 1108.8000 ;
	    RECT 825.0000 1103.7001 826.2000 1107.9000 ;
	    RECT 827.4000 1104.0000 828.6000 1108.8000 ;
	    RECT 829.8000 1104.9000 831.0000 1109.7001 ;
	    RECT 832.2000 1104.0000 833.4000 1109.7001 ;
	    RECT 904.2000 1107.4501 905.4000 1107.6000 ;
	    RECT 928.2000 1107.4501 929.4000 1107.6000 ;
	    RECT 904.2000 1106.5500 929.4000 1107.4501 ;
	    RECT 964.2000 1106.7001 965.4000 1109.7001 ;
	    RECT 904.2000 1106.4000 905.4000 1106.5500 ;
	    RECT 928.2000 1106.4000 929.4000 1106.5500 ;
	    RECT 827.4000 1103.7001 833.4000 1104.0000 ;
	    RECT 901.8000 1104.4501 903.0000 1104.6000 ;
	    RECT 909.0000 1104.4501 910.2000 1104.6000 ;
	    RECT 825.0000 1101.6000 825.9000 1103.7001 ;
	    RECT 827.7000 1103.1000 833.1000 1103.7001 ;
	    RECT 901.8000 1103.5500 910.2000 1104.4501 ;
	    RECT 901.8000 1103.4000 903.0000 1103.5500 ;
	    RECT 909.0000 1103.4000 910.2000 1103.5500 ;
	    RECT 930.6000 1104.4501 931.8000 1104.6000 ;
	    RECT 964.2000 1104.4501 965.4000 1104.6000 ;
	    RECT 930.6000 1103.5500 965.4000 1104.4501 ;
	    RECT 966.6000 1104.0000 967.8000 1109.7001 ;
	    RECT 930.6000 1103.4000 931.8000 1103.5500 ;
	    RECT 964.2000 1103.4000 965.4000 1103.5500 ;
	    RECT 966.3000 1102.8000 967.8000 1104.0000 ;
	    RECT 777.0000 1100.4000 778.2000 1101.6000 ;
	    RECT 793.8000 1101.4501 795.0000 1101.6000 ;
	    RECT 820.2000 1101.4501 821.4000 1101.6000 ;
	    RECT 793.8000 1100.5500 821.4000 1101.4501 ;
	    RECT 793.8000 1100.4000 795.0000 1100.5500 ;
	    RECT 820.2000 1100.4000 821.4000 1100.5500 ;
	    RECT 822.6000 1100.4000 823.8000 1101.6000 ;
	    RECT 825.0000 1100.7001 826.5000 1101.6000 ;
	    RECT 827.4000 1100.4000 828.6000 1101.6000 ;
	    RECT 831.0000 1100.7001 831.3000 1102.2001 ;
	    RECT 832.2000 1100.4000 833.4000 1101.6000 ;
	    RECT 825.0000 1099.5000 826.2000 1099.8000 ;
	    RECT 829.8000 1099.5000 831.0000 1099.8000 ;
	    RECT 678.6000 1097.5500 684.4500 1098.4501 ;
	    RECT 678.6000 1097.4000 679.8000 1097.5500 ;
	    RECT 676.8000 1094.4000 678.3000 1095.3000 ;
	    RECT 675.0000 1092.6000 675.9000 1093.5000 ;
	    RECT 675.0000 1091.4000 676.2000 1092.6000 ;
	    RECT 642.6000 1083.3000 643.8000 1089.3000 ;
	    RECT 674.7000 1083.3000 675.9000 1089.3000 ;
	    RECT 677.1000 1083.3000 678.3000 1094.4000 ;
	    RECT 681.0000 1083.3000 682.2000 1095.3000 ;
	    RECT 695.4000 1083.3000 696.6000 1089.3000 ;
	    RECT 697.8000 1083.3000 699.0000 1099.5000 ;
	    RECT 733.8000 1098.4501 735.0000 1098.6000 ;
	    RECT 745.8000 1098.4501 747.0000 1098.6000 ;
	    RECT 733.8000 1097.5500 747.0000 1098.4501 ;
	    RECT 749.7000 1098.3000 750.9000 1098.6000 ;
	    RECT 733.8000 1097.4000 735.0000 1097.5500 ;
	    RECT 745.8000 1097.4000 747.0000 1097.5500 ;
	    RECT 748.5000 1097.4000 750.9000 1098.3000 ;
	    RECT 753.0000 1098.4501 754.2000 1098.6000 ;
	    RECT 774.6000 1098.4501 775.8000 1098.6000 ;
	    RECT 753.0000 1097.5500 775.8000 1098.4501 ;
	    RECT 753.0000 1097.4000 754.2000 1097.5500 ;
	    RECT 774.6000 1097.4000 775.8000 1097.5500 ;
	    RECT 748.5000 1097.1000 749.7000 1097.4000 ;
	    RECT 745.8000 1095.3000 746.7000 1096.5000 ;
	    RECT 767.4000 1095.4501 768.6000 1095.6000 ;
	    RECT 772.2000 1095.4501 773.4000 1095.6000 ;
	    RECT 738.6000 1094.4000 742.2000 1095.3000 ;
	    RECT 738.6000 1083.3000 739.8000 1094.4000 ;
	    RECT 741.0000 1094.1000 742.2000 1094.4000 ;
	    RECT 741.0000 1083.3000 742.5000 1093.2001 ;
	    RECT 745.2000 1083.3000 747.6000 1095.3000 ;
	    RECT 750.3000 1094.4000 754.2000 1095.3000 ;
	    RECT 767.4000 1094.5500 773.4000 1095.4501 ;
	    RECT 767.4000 1094.4000 768.6000 1094.5500 ;
	    RECT 772.2000 1094.4000 773.4000 1094.5500 ;
	    RECT 750.3000 1094.1000 751.5000 1094.4000 ;
	    RECT 750.3000 1083.3000 751.8000 1093.2001 ;
	    RECT 753.0000 1083.3000 754.2000 1094.4000 ;
	    RECT 772.2000 1093.2001 773.4000 1093.5000 ;
	    RECT 772.2000 1083.3000 773.4000 1089.3000 ;
	    RECT 774.6000 1083.3000 775.8000 1096.5000 ;
	    RECT 777.0000 1083.3000 778.2000 1089.3000 ;
	    RECT 791.4000 1083.3000 792.6000 1089.3000 ;
	    RECT 793.8000 1083.3000 795.0000 1099.5000 ;
	    RECT 822.6000 1099.2001 823.8000 1099.5000 ;
	    RECT 825.0000 1097.4000 826.2000 1098.6000 ;
	    RECT 827.7000 1095.3000 828.6000 1099.5000 ;
	    RECT 829.8000 1098.4501 831.0000 1098.6000 ;
	    RECT 832.2000 1098.4501 833.4000 1098.6000 ;
	    RECT 829.8000 1097.5500 833.4000 1098.4501 ;
	    RECT 829.8000 1097.4000 831.0000 1097.5500 ;
	    RECT 832.2000 1097.4000 833.4000 1097.5500 ;
	    RECT 873.0000 1098.4501 874.2000 1098.6000 ;
	    RECT 940.2000 1098.4501 941.4000 1098.6000 ;
	    RECT 873.0000 1097.5500 941.4000 1098.4501 ;
	    RECT 873.0000 1097.4000 874.2000 1097.5500 ;
	    RECT 940.2000 1097.4000 941.4000 1097.5500 ;
	    RECT 966.3000 1096.2001 967.5000 1102.8000 ;
	    RECT 969.0000 1101.9000 970.2000 1109.7001 ;
	    RECT 973.8000 1103.7001 975.0000 1109.7001 ;
	    RECT 978.6000 1104.9000 979.8000 1109.7001 ;
	    RECT 981.0000 1105.5000 982.2000 1109.7001 ;
	    RECT 983.4000 1105.5000 984.6000 1109.7001 ;
	    RECT 985.8000 1105.5000 987.0000 1109.7001 ;
	    RECT 988.2000 1105.5000 989.4000 1109.7001 ;
	    RECT 990.6000 1106.7001 991.8000 1109.7001 ;
	    RECT 993.0000 1105.5000 994.2000 1109.7001 ;
	    RECT 995.4000 1106.7001 996.6000 1109.7001 ;
	    RECT 997.8000 1105.5000 999.0000 1109.7001 ;
	    RECT 1000.2000 1105.5000 1001.4000 1109.7001 ;
	    RECT 1002.6000 1105.5000 1003.8000 1109.7001 ;
	    RECT 976.2000 1103.7001 979.8000 1104.9000 ;
	    RECT 1005.0000 1104.9000 1006.2000 1109.7001 ;
	    RECT 976.2000 1102.8000 977.4000 1103.7001 ;
	    RECT 968.4000 1101.0000 970.2000 1101.9000 ;
	    RECT 974.7000 1101.9000 977.4000 1102.8000 ;
	    RECT 983.4000 1103.4000 984.9000 1104.6000 ;
	    RECT 989.4000 1103.4000 989.7000 1104.6000 ;
	    RECT 990.6000 1103.4000 991.8000 1104.6000 ;
	    RECT 993.0000 1103.7001 999.9000 1104.6000 ;
	    RECT 1005.0000 1103.7001 1008.9000 1104.9000 ;
	    RECT 1009.8000 1103.7001 1011.0000 1109.7001 ;
	    RECT 993.0000 1103.4000 994.2000 1103.7001 ;
	    RECT 968.4000 1098.0000 969.3000 1101.0000 ;
	    RECT 974.7000 1100.1000 975.9000 1101.9000 ;
	    RECT 970.2000 1098.9000 975.9000 1100.1000 ;
	    RECT 983.4000 1099.2001 984.6000 1103.4000 ;
	    RECT 995.4000 1102.5000 996.6000 1102.8000 ;
	    RECT 993.0000 1102.2001 994.2000 1102.5000 ;
	    RECT 987.6000 1101.3000 994.2000 1102.2001 ;
	    RECT 987.6000 1101.0000 988.8000 1101.3000 ;
	    RECT 995.4000 1100.4000 996.6000 1101.6000 ;
	    RECT 998.7000 1100.1000 999.9000 1103.7001 ;
	    RECT 1007.7000 1102.8000 1008.9000 1103.7001 ;
	    RECT 1007.7000 1101.6000 1012.2000 1102.8000 ;
	    RECT 1014.6000 1100.7001 1015.8000 1109.7001 ;
	    RECT 1045.8000 1104.0000 1047.0000 1109.7001 ;
	    RECT 1048.2001 1104.9000 1049.4000 1109.7001 ;
	    RECT 1050.6000 1108.8000 1056.6000 1109.7001 ;
	    RECT 1050.6000 1104.0000 1051.8000 1108.8000 ;
	    RECT 1045.8000 1103.7001 1051.8000 1104.0000 ;
	    RECT 1053.0000 1103.7001 1054.2001 1107.9000 ;
	    RECT 1055.4000 1103.7001 1056.6000 1108.8000 ;
	    RECT 1108.2001 1103.7001 1109.4000 1109.7001 ;
	    RECT 1046.1000 1103.1000 1051.5000 1103.7001 ;
	    RECT 988.2000 1098.9000 993.0000 1100.1000 ;
	    RECT 998.7000 1098.9000 1001.7000 1100.1000 ;
	    RECT 1002.6000 1099.5000 1015.8000 1100.7001 ;
	    RECT 1045.8000 1100.4000 1047.0000 1101.6000 ;
	    RECT 1047.9000 1100.7001 1048.2001 1102.2001 ;
	    RECT 1053.3000 1101.6000 1054.2001 1103.7001 ;
	    RECT 1110.6000 1102.8000 1111.8000 1109.7001 ;
	    RECT 1113.0000 1103.7001 1114.2001 1109.7001 ;
	    RECT 1115.4000 1102.8000 1116.6000 1109.7001 ;
	    RECT 1117.8000 1103.7001 1119.0000 1109.7001 ;
	    RECT 1120.2001 1102.8000 1121.4000 1109.7001 ;
	    RECT 1122.6000 1103.7001 1123.8000 1109.7001 ;
	    RECT 1125.0000 1102.8000 1126.2001 1109.7001 ;
	    RECT 1127.4000 1103.7001 1128.6000 1109.7001 ;
	    RECT 1110.6000 1101.6000 1113.3000 1102.8000 ;
	    RECT 1115.4000 1101.6000 1118.7001 1102.8000 ;
	    RECT 1120.2001 1101.6000 1123.5000 1102.8000 ;
	    RECT 1125.0000 1101.6000 1128.6000 1102.8000 ;
	    RECT 1149.0000 1102.5000 1150.2001 1109.7001 ;
	    RECT 1151.4000 1106.7001 1152.6000 1109.7001 ;
	    RECT 1151.4000 1105.5000 1152.6000 1105.8000 ;
	    RECT 1151.4000 1104.4501 1152.6000 1104.6000 ;
	    RECT 1223.4000 1104.4501 1224.6000 1104.6000 ;
	    RECT 1151.4000 1103.5500 1224.6000 1104.4501 ;
	    RECT 1151.4000 1103.4000 1152.6000 1103.5500 ;
	    RECT 1223.4000 1103.4000 1224.6000 1103.5500 ;
	    RECT 1050.6000 1100.4000 1051.8000 1101.6000 ;
	    RECT 1052.7001 1100.7001 1054.2001 1101.6000 ;
	    RECT 1055.4000 1101.4501 1056.6000 1101.6000 ;
	    RECT 1060.2001 1101.4501 1061.4000 1101.6000 ;
	    RECT 1055.4000 1100.5500 1061.4000 1101.4501 ;
	    RECT 1112.1000 1100.7001 1113.3000 1101.6000 ;
	    RECT 1117.5000 1100.7001 1118.7001 1101.6000 ;
	    RECT 1122.3000 1100.7001 1123.5000 1101.6000 ;
	    RECT 1055.4000 1100.4000 1056.6000 1100.5500 ;
	    RECT 1060.2001 1100.4000 1061.4000 1100.5500 ;
	    RECT 1048.2001 1099.5000 1049.4000 1099.8000 ;
	    RECT 1053.0000 1099.5000 1054.2001 1099.8000 ;
	    RECT 1110.3000 1099.5000 1110.9000 1100.7001 ;
	    RECT 1112.1000 1099.5000 1116.0000 1100.7001 ;
	    RECT 1117.5000 1099.5000 1121.1000 1100.7001 ;
	    RECT 1122.3000 1099.5000 1126.2001 1100.7001 ;
	    RECT 1127.4000 1099.5000 1128.6000 1101.6000 ;
	    RECT 1129.8000 1101.4501 1131.0000 1101.6000 ;
	    RECT 1149.0000 1101.4501 1150.2001 1101.6000 ;
	    RECT 1129.8000 1100.5500 1150.2001 1101.4501 ;
	    RECT 1129.8000 1100.4000 1131.0000 1100.5500 ;
	    RECT 1149.0000 1100.4000 1150.2001 1100.5500 ;
	    RECT 1278.6000 1100.7001 1279.8000 1109.7001 ;
	    RECT 1283.4000 1103.7001 1284.6000 1109.7001 ;
	    RECT 1288.2001 1104.9000 1289.4000 1109.7001 ;
	    RECT 1290.6000 1105.5000 1291.8000 1109.7001 ;
	    RECT 1293.0000 1105.5000 1294.2001 1109.7001 ;
	    RECT 1295.4000 1105.5000 1296.6000 1109.7001 ;
	    RECT 1297.8000 1106.7001 1299.0000 1109.7001 ;
	    RECT 1300.2001 1105.5000 1301.4000 1109.7001 ;
	    RECT 1302.6000 1106.7001 1303.8000 1109.7001 ;
	    RECT 1305.0000 1105.5000 1306.2001 1109.7001 ;
	    RECT 1307.4000 1105.5000 1308.6000 1109.7001 ;
	    RECT 1309.8000 1105.5000 1311.0000 1109.7001 ;
	    RECT 1312.2001 1105.5000 1313.4000 1109.7001 ;
	    RECT 1285.5000 1103.7001 1289.4000 1104.9000 ;
	    RECT 1314.6000 1104.9000 1315.8000 1109.7001 ;
	    RECT 1294.5000 1103.7001 1301.4000 1104.6000 ;
	    RECT 1285.5000 1102.8000 1286.7001 1103.7001 ;
	    RECT 1282.2001 1101.6000 1286.7001 1102.8000 ;
	    RECT 1278.6000 1099.5000 1291.8000 1100.7001 ;
	    RECT 1294.5000 1100.1000 1295.7001 1103.7001 ;
	    RECT 1300.2001 1103.4000 1301.4000 1103.7001 ;
	    RECT 1302.6000 1103.4000 1303.8000 1104.6000 ;
	    RECT 1304.7001 1103.4000 1305.0000 1104.6000 ;
	    RECT 1309.5000 1103.4000 1311.0000 1104.6000 ;
	    RECT 1314.6000 1103.7001 1318.2001 1104.9000 ;
	    RECT 1319.4000 1103.7001 1320.6000 1109.7001 ;
	    RECT 1297.8000 1102.5000 1299.0000 1102.8000 ;
	    RECT 1300.2001 1102.2001 1301.4000 1102.5000 ;
	    RECT 1297.8000 1100.4000 1299.0000 1101.6000 ;
	    RECT 1300.2001 1101.3000 1306.8000 1102.2001 ;
	    RECT 1305.6000 1101.0000 1306.8000 1101.3000 ;
	    RECT 978.6000 1098.0000 979.8000 1098.9000 ;
	    RECT 968.4000 1097.1000 969.6000 1098.0000 ;
	    RECT 978.6000 1097.1000 1004.1000 1098.0000 ;
	    RECT 1005.0000 1097.4000 1006.2000 1098.6000 ;
	    RECT 1012.5000 1098.0000 1013.7000 1098.3000 ;
	    RECT 1007.1000 1097.1000 1013.7000 1098.0000 ;
	    RECT 880.2000 1095.4501 881.4000 1095.6000 ;
	    RECT 940.2000 1095.4501 941.4000 1095.6000 ;
	    RECT 822.6000 1083.3000 823.8000 1095.3000 ;
	    RECT 826.5000 1083.3000 829.5000 1095.3000 ;
	    RECT 832.2000 1083.3000 833.4000 1095.3000 ;
	    RECT 880.2000 1094.5500 941.4000 1095.4501 ;
	    RECT 966.3000 1095.0000 967.8000 1096.2001 ;
	    RECT 880.2000 1094.4000 881.4000 1094.5500 ;
	    RECT 940.2000 1094.4000 941.4000 1094.5500 ;
	    RECT 966.6000 1093.5000 967.8000 1095.0000 ;
	    RECT 968.7000 1094.4000 969.6000 1097.1000 ;
	    RECT 970.5000 1096.2001 971.7000 1096.5000 ;
	    RECT 970.5000 1095.3000 1008.9000 1096.2001 ;
	    RECT 1004.7000 1095.0000 1005.9000 1095.3000 ;
	    RECT 1009.8000 1094.4000 1011.0000 1095.6000 ;
	    RECT 968.7000 1093.5000 982.2000 1094.4000 ;
	    RECT 851.4000 1092.4501 852.6000 1092.6000 ;
	    RECT 885.0000 1092.4501 886.2000 1092.6000 ;
	    RECT 851.4000 1091.5500 886.2000 1092.4501 ;
	    RECT 851.4000 1091.4000 852.6000 1091.5500 ;
	    RECT 885.0000 1091.4000 886.2000 1091.5500 ;
	    RECT 887.4000 1092.4501 888.6000 1092.6000 ;
	    RECT 966.6000 1092.4501 967.8000 1092.6000 ;
	    RECT 887.4000 1091.5500 967.8000 1092.4501 ;
	    RECT 887.4000 1091.4000 888.6000 1091.5500 ;
	    RECT 966.6000 1091.4000 967.8000 1091.5500 ;
	    RECT 968.7000 1091.1000 969.6000 1093.5000 ;
	    RECT 981.0000 1093.2001 982.2000 1093.5000 ;
	    RECT 985.8000 1093.5000 998.7000 1094.4000 ;
	    RECT 985.8000 1093.2001 987.0000 1093.5000 ;
	    RECT 973.5000 1091.4000 977.4000 1092.6000 ;
	    RECT 863.4000 1086.4501 864.6000 1086.6000 ;
	    RECT 930.6000 1086.4501 931.8000 1086.6000 ;
	    RECT 863.4000 1085.5500 931.8000 1086.4501 ;
	    RECT 863.4000 1085.4000 864.6000 1085.5500 ;
	    RECT 930.6000 1085.4000 931.8000 1085.5500 ;
	    RECT 964.2000 1083.3000 965.4000 1089.3000 ;
	    RECT 966.6000 1083.3000 967.8000 1090.5000 ;
	    RECT 968.7000 1090.2001 972.6000 1091.1000 ;
	    RECT 969.0000 1083.3000 970.2000 1089.3000 ;
	    RECT 971.4000 1083.3000 972.6000 1090.2001 ;
	    RECT 973.8000 1083.3000 975.0000 1089.3000 ;
	    RECT 976.2000 1083.3000 977.4000 1091.4000 ;
	    RECT 978.3000 1090.2001 984.6000 1091.4000 ;
	    RECT 978.6000 1083.3000 979.8000 1089.3000 ;
	    RECT 981.0000 1083.3000 982.2000 1087.5000 ;
	    RECT 983.4000 1083.3000 984.6000 1087.5000 ;
	    RECT 985.8000 1083.3000 987.0000 1087.5000 ;
	    RECT 988.2000 1083.3000 989.4000 1092.6000 ;
	    RECT 993.0000 1091.4000 996.9000 1092.6000 ;
	    RECT 997.8000 1092.3000 998.7000 1093.5000 ;
	    RECT 1000.2000 1094.1000 1001.4000 1094.4000 ;
	    RECT 1000.2000 1093.5000 1008.3000 1094.1000 ;
	    RECT 1000.2000 1093.2001 1009.5000 1093.5000 ;
	    RECT 1007.4000 1092.3000 1009.5000 1093.2001 ;
	    RECT 997.8000 1091.4000 1006.5000 1092.3000 ;
	    RECT 1011.0000 1092.0000 1013.4000 1093.2001 ;
	    RECT 1011.0000 1091.4000 1011.9000 1092.0000 ;
	    RECT 990.6000 1083.3000 991.8000 1089.3000 ;
	    RECT 993.0000 1083.3000 994.2000 1090.5000 ;
	    RECT 995.4000 1083.3000 996.6000 1089.3000 ;
	    RECT 997.8000 1083.3000 999.0000 1090.5000 ;
	    RECT 1005.6000 1090.2001 1011.9000 1091.4000 ;
	    RECT 1014.6000 1091.1000 1015.8000 1099.5000 ;
	    RECT 1021.8000 1098.4501 1023.0000 1098.6000 ;
	    RECT 1048.2001 1098.4501 1049.4000 1098.6000 ;
	    RECT 1021.8000 1097.5500 1049.4000 1098.4501 ;
	    RECT 1021.8000 1097.4000 1023.0000 1097.5500 ;
	    RECT 1048.2001 1097.4000 1049.4000 1097.5500 ;
	    RECT 1050.6000 1095.3000 1051.5000 1099.5000 ;
	    RECT 1055.4000 1099.2001 1056.6000 1099.5000 ;
	    RECT 1053.0000 1097.4000 1054.2001 1098.6000 ;
	    RECT 1112.1000 1097.4000 1113.3000 1099.5000 ;
	    RECT 1117.5000 1097.4000 1118.7001 1099.5000 ;
	    RECT 1122.3000 1097.4000 1123.5000 1099.5000 ;
	    RECT 1127.4000 1098.4501 1128.6000 1098.6000 ;
	    RECT 1134.6000 1098.4501 1135.8000 1098.6000 ;
	    RECT 1146.6000 1098.4501 1147.8000 1098.6000 ;
	    RECT 1127.4000 1097.5500 1147.8000 1098.4501 ;
	    RECT 1127.4000 1097.4000 1128.6000 1097.5500 ;
	    RECT 1134.6000 1097.4000 1135.8000 1097.5500 ;
	    RECT 1146.6000 1097.4000 1147.8000 1097.5500 ;
	    RECT 1110.6000 1096.2001 1113.3000 1097.4000 ;
	    RECT 1115.4000 1096.2001 1118.7001 1097.4000 ;
	    RECT 1120.2001 1096.2001 1123.5000 1097.4000 ;
	    RECT 1125.0000 1096.5000 1126.5000 1097.4000 ;
	    RECT 1125.0000 1096.2001 1128.6000 1096.5000 ;
	    RECT 1012.8000 1090.2001 1015.8000 1091.1000 ;
	    RECT 1000.2000 1083.3000 1001.4000 1087.5000 ;
	    RECT 1002.6000 1083.3000 1003.8000 1087.5000 ;
	    RECT 1005.0000 1083.3000 1006.2000 1089.3000 ;
	    RECT 1007.4000 1083.3000 1008.6000 1090.2001 ;
	    RECT 1012.8000 1089.3000 1013.7000 1090.2001 ;
	    RECT 1009.8000 1082.4000 1011.0000 1089.3000 ;
	    RECT 1012.2000 1088.4000 1013.7000 1089.3000 ;
	    RECT 1012.2000 1083.3000 1013.4000 1088.4000 ;
	    RECT 1014.6000 1083.3000 1015.8000 1089.3000 ;
	    RECT 1045.8000 1083.3000 1047.0000 1095.3000 ;
	    RECT 1049.7001 1083.3000 1052.7001 1095.3000 ;
	    RECT 1055.4000 1083.3000 1056.6000 1095.3000 ;
	    RECT 1108.2001 1083.3000 1109.4000 1095.3000 ;
	    RECT 1110.6000 1083.3000 1111.8000 1096.2001 ;
	    RECT 1113.0000 1083.3000 1114.2001 1095.3000 ;
	    RECT 1115.4000 1083.3000 1116.6000 1096.2001 ;
	    RECT 1117.8000 1083.3000 1119.0000 1095.3000 ;
	    RECT 1120.2001 1083.3000 1121.4000 1096.2001 ;
	    RECT 1122.6000 1083.3000 1123.8000 1095.3000 ;
	    RECT 1125.0000 1083.3000 1126.2001 1096.2001 ;
	    RECT 1127.4000 1083.3000 1128.6000 1095.3000 ;
	    RECT 1149.0000 1083.3000 1150.2001 1099.5000 ;
	    RECT 1278.6000 1091.1000 1279.8000 1099.5000 ;
	    RECT 1292.7001 1098.9000 1295.7001 1100.1000 ;
	    RECT 1301.4000 1098.9000 1306.2001 1100.1000 ;
	    RECT 1309.8000 1099.2001 1311.0000 1103.4000 ;
	    RECT 1317.0000 1102.8000 1318.2001 1103.7001 ;
	    RECT 1317.0000 1101.9000 1319.7001 1102.8000 ;
	    RECT 1318.5000 1100.1000 1319.7001 1101.9000 ;
	    RECT 1324.2001 1101.9000 1325.4000 1109.7001 ;
	    RECT 1326.6000 1104.0000 1327.8000 1109.7001 ;
	    RECT 1329.0000 1106.7001 1330.2001 1109.7001 ;
	    RECT 1326.6000 1102.8000 1328.1000 1104.0000 ;
	    RECT 1348.2001 1103.7001 1349.4000 1109.7001 ;
	    RECT 1352.1000 1104.6000 1353.3000 1109.7001 ;
	    RECT 1350.6000 1103.7001 1353.3000 1104.6000 ;
	    RECT 1386.6000 1104.0000 1387.8000 1109.7001 ;
	    RECT 1389.0000 1104.9000 1390.2001 1109.7001 ;
	    RECT 1391.4000 1104.0000 1392.6000 1109.7001 ;
	    RECT 1386.6000 1103.7001 1392.6000 1104.0000 ;
	    RECT 1393.8000 1103.7001 1395.0000 1109.7001 ;
	    RECT 1408.2001 1106.7001 1409.4000 1109.7001 ;
	    RECT 1408.2001 1105.5000 1409.4000 1105.8000 ;
	    RECT 1324.2001 1101.0000 1326.0000 1101.9000 ;
	    RECT 1318.5000 1098.9000 1324.2001 1100.1000 ;
	    RECT 1280.7001 1098.0000 1281.9000 1098.3000 ;
	    RECT 1280.7001 1097.1000 1287.3000 1098.0000 ;
	    RECT 1288.2001 1097.4000 1289.4000 1098.6000 ;
	    RECT 1314.6000 1098.0000 1315.8000 1098.9000 ;
	    RECT 1325.1000 1098.0000 1326.0000 1101.0000 ;
	    RECT 1290.3000 1097.1000 1315.8000 1098.0000 ;
	    RECT 1324.8000 1097.1000 1326.0000 1098.0000 ;
	    RECT 1322.7001 1096.2001 1323.9000 1096.5000 ;
	    RECT 1283.4000 1094.4000 1284.6000 1095.6000 ;
	    RECT 1285.5000 1095.3000 1323.9000 1096.2001 ;
	    RECT 1288.5000 1095.0000 1289.7001 1095.3000 ;
	    RECT 1324.8000 1094.4000 1325.7001 1097.1000 ;
	    RECT 1326.9000 1096.2001 1328.1000 1102.8000 ;
	    RECT 1348.2001 1102.5000 1349.4000 1102.8000 ;
	    RECT 1348.2001 1100.4000 1349.4000 1101.6000 ;
	    RECT 1350.6000 1099.5000 1351.8000 1103.7001 ;
	    RECT 1386.9000 1103.1000 1392.3000 1103.7001 ;
	    RECT 1393.8000 1102.5000 1394.7001 1103.7001 ;
	    RECT 1408.2001 1103.4000 1409.4000 1104.6000 ;
	    RECT 1410.6000 1102.5000 1411.8000 1109.7001 ;
	    RECT 1434.6000 1103.7001 1435.8000 1109.7001 ;
	    RECT 1437.0000 1104.0000 1438.2001 1109.7001 ;
	    RECT 1439.4000 1104.9000 1440.6000 1109.7001 ;
	    RECT 1441.8000 1104.0000 1443.0000 1109.7001 ;
	    RECT 1437.0000 1103.7001 1443.0000 1104.0000 ;
	    RECT 1468.2001 1104.0000 1469.4000 1109.7001 ;
	    RECT 1470.6000 1104.9000 1471.8000 1109.7001 ;
	    RECT 1473.0000 1104.0000 1474.2001 1109.7001 ;
	    RECT 1468.2001 1103.7001 1474.2001 1104.0000 ;
	    RECT 1475.4000 1103.7001 1476.6000 1109.7001 ;
	    RECT 1501.8000 1104.0000 1503.0000 1109.7001 ;
	    RECT 1504.2001 1104.9000 1505.4000 1109.7001 ;
	    RECT 1506.6000 1104.0000 1507.8000 1109.7001 ;
	    RECT 1501.8000 1103.7001 1507.8000 1104.0000 ;
	    RECT 1509.0000 1103.7001 1510.2001 1109.7001 ;
	    RECT 1528.2001 1103.7001 1529.4000 1109.7001 ;
	    RECT 1532.1000 1104.6000 1533.3000 1109.7001 ;
	    RECT 1530.6000 1103.7001 1533.3000 1104.6000 ;
	    RECT 1434.9000 1102.5000 1435.8000 1103.7001 ;
	    RECT 1437.3000 1103.1000 1442.7001 1103.7001 ;
	    RECT 1468.5000 1103.1000 1473.9000 1103.7001 ;
	    RECT 1475.4000 1102.5000 1476.3000 1103.7001 ;
	    RECT 1502.1000 1103.1000 1507.5000 1103.7001 ;
	    RECT 1509.0000 1102.5000 1509.9000 1103.7001 ;
	    RECT 1528.2001 1102.5000 1529.4000 1102.8000 ;
	    RECT 1374.6000 1101.4501 1375.8000 1101.6000 ;
	    RECT 1386.6000 1101.4501 1387.8000 1101.6000 ;
	    RECT 1374.6000 1100.5500 1387.8000 1101.4501 ;
	    RECT 1388.7001 1100.7001 1389.0000 1102.2001 ;
	    RECT 1374.6000 1100.4000 1375.8000 1100.5500 ;
	    RECT 1386.6000 1100.4000 1387.8000 1100.5500 ;
	    RECT 1391.1000 1100.4000 1392.9000 1101.6000 ;
	    RECT 1393.8000 1101.4501 1395.0000 1101.6000 ;
	    RECT 1405.8000 1101.4501 1407.0000 1101.6000 ;
	    RECT 1393.8000 1100.5500 1407.0000 1101.4501 ;
	    RECT 1393.8000 1100.4000 1395.0000 1100.5500 ;
	    RECT 1405.8000 1100.4000 1407.0000 1100.5500 ;
	    RECT 1410.6000 1101.4501 1411.8000 1101.6000 ;
	    RECT 1429.8000 1101.4501 1431.0000 1101.6000 ;
	    RECT 1410.6000 1100.5500 1431.0000 1101.4501 ;
	    RECT 1410.6000 1100.4000 1411.8000 1100.5500 ;
	    RECT 1429.8000 1100.4000 1431.0000 1100.5500 ;
	    RECT 1432.2001 1101.4501 1433.4000 1101.6000 ;
	    RECT 1434.6000 1101.4501 1435.8000 1101.6000 ;
	    RECT 1432.2001 1100.5500 1435.8000 1101.4501 ;
	    RECT 1432.2001 1100.4000 1433.4000 1100.5500 ;
	    RECT 1434.6000 1100.4000 1435.8000 1100.5500 ;
	    RECT 1436.7001 1100.4000 1438.5000 1101.6000 ;
	    RECT 1440.6000 1100.7001 1440.9000 1102.2001 ;
	    RECT 1441.8000 1100.4000 1443.0000 1101.6000 ;
	    RECT 1444.2001 1101.4501 1445.4000 1101.6000 ;
	    RECT 1468.2001 1101.4501 1469.4000 1101.6000 ;
	    RECT 1444.2001 1100.5500 1469.4000 1101.4501 ;
	    RECT 1470.3000 1100.7001 1470.6000 1102.2001 ;
	    RECT 1444.2001 1100.4000 1445.4000 1100.5500 ;
	    RECT 1468.2001 1100.4000 1469.4000 1100.5500 ;
	    RECT 1472.7001 1100.4000 1474.5000 1101.6000 ;
	    RECT 1475.4000 1101.4501 1476.6000 1101.6000 ;
	    RECT 1482.6000 1101.4501 1483.8000 1101.6000 ;
	    RECT 1475.4000 1100.5500 1483.8000 1101.4501 ;
	    RECT 1475.4000 1100.4000 1476.6000 1100.5500 ;
	    RECT 1482.6000 1100.4000 1483.8000 1100.5500 ;
	    RECT 1492.2001 1101.4501 1493.4000 1101.6000 ;
	    RECT 1501.8000 1101.4501 1503.0000 1101.6000 ;
	    RECT 1492.2001 1100.5500 1503.0000 1101.4501 ;
	    RECT 1503.9000 1100.7001 1504.2001 1102.2001 ;
	    RECT 1492.2001 1100.4000 1493.4000 1100.5500 ;
	    RECT 1501.8000 1100.4000 1503.0000 1100.5500 ;
	    RECT 1506.3000 1100.4000 1508.1000 1101.6000 ;
	    RECT 1509.0000 1100.4000 1510.2001 1101.6000 ;
	    RECT 1513.8000 1101.4501 1515.0000 1101.6000 ;
	    RECT 1528.2001 1101.4501 1529.4000 1101.6000 ;
	    RECT 1513.8000 1100.5500 1529.4000 1101.4501 ;
	    RECT 1513.8000 1100.4000 1515.0000 1100.5500 ;
	    RECT 1528.2001 1100.4000 1529.4000 1100.5500 ;
	    RECT 1389.0000 1099.5000 1390.2001 1099.8000 ;
	    RECT 1350.6000 1098.4501 1351.8000 1098.6000 ;
	    RECT 1367.4000 1098.4501 1368.6000 1098.6000 ;
	    RECT 1350.6000 1097.5500 1368.6000 1098.4501 ;
	    RECT 1350.6000 1097.4000 1351.8000 1097.5500 ;
	    RECT 1367.4000 1097.4000 1368.6000 1097.5500 ;
	    RECT 1386.6000 1098.4501 1387.8000 1098.6000 ;
	    RECT 1389.0000 1098.4501 1390.2001 1098.6000 ;
	    RECT 1386.6000 1097.5500 1390.2001 1098.4501 ;
	    RECT 1386.6000 1097.4000 1387.8000 1097.5500 ;
	    RECT 1389.0000 1097.4000 1390.2001 1097.5500 ;
	    RECT 1293.0000 1094.1000 1294.2001 1094.4000 ;
	    RECT 1286.1000 1093.5000 1294.2001 1094.1000 ;
	    RECT 1284.9000 1093.2001 1294.2001 1093.5000 ;
	    RECT 1295.7001 1093.5000 1308.6000 1094.4000 ;
	    RECT 1281.0000 1092.0000 1283.4000 1093.2001 ;
	    RECT 1284.9000 1092.3000 1287.0000 1093.2001 ;
	    RECT 1295.7001 1092.3000 1296.6000 1093.5000 ;
	    RECT 1307.4000 1093.2001 1308.6000 1093.5000 ;
	    RECT 1312.2001 1093.5000 1325.7001 1094.4000 ;
	    RECT 1326.6000 1095.0000 1328.1000 1096.2001 ;
	    RECT 1326.6000 1093.5000 1327.8000 1095.0000 ;
	    RECT 1312.2001 1093.2001 1313.4000 1093.5000 ;
	    RECT 1282.5000 1091.4000 1283.4000 1092.0000 ;
	    RECT 1287.9000 1091.4000 1296.6000 1092.3000 ;
	    RECT 1297.5000 1091.4000 1301.4000 1092.6000 ;
	    RECT 1278.6000 1090.2001 1281.6000 1091.1000 ;
	    RECT 1282.5000 1090.2001 1288.8000 1091.4000 ;
	    RECT 1280.7001 1089.3000 1281.6000 1090.2001 ;
	    RECT 1151.4000 1083.3000 1152.6000 1089.3000 ;
	    RECT 1278.6000 1083.3000 1279.8000 1089.3000 ;
	    RECT 1280.7001 1088.4000 1282.2001 1089.3000 ;
	    RECT 1281.0000 1083.3000 1282.2001 1088.4000 ;
	    RECT 1283.4000 1082.4000 1284.6000 1089.3000 ;
	    RECT 1285.8000 1083.3000 1287.0000 1090.2001 ;
	    RECT 1288.2001 1083.3000 1289.4000 1089.3000 ;
	    RECT 1290.6000 1083.3000 1291.8000 1087.5000 ;
	    RECT 1293.0000 1083.3000 1294.2001 1087.5000 ;
	    RECT 1295.4000 1083.3000 1296.6000 1090.5000 ;
	    RECT 1297.8000 1083.3000 1299.0000 1089.3000 ;
	    RECT 1300.2001 1083.3000 1301.4000 1090.5000 ;
	    RECT 1302.6000 1083.3000 1303.8000 1089.3000 ;
	    RECT 1305.0000 1083.3000 1306.2001 1092.6000 ;
	    RECT 1317.0000 1091.4000 1320.9000 1092.6000 ;
	    RECT 1309.8000 1090.2001 1316.1000 1091.4000 ;
	    RECT 1307.4000 1083.3000 1308.6000 1087.5000 ;
	    RECT 1309.8000 1083.3000 1311.0000 1087.5000 ;
	    RECT 1312.2001 1083.3000 1313.4000 1087.5000 ;
	    RECT 1314.6000 1083.3000 1315.8000 1089.3000 ;
	    RECT 1317.0000 1083.3000 1318.2001 1091.4000 ;
	    RECT 1324.8000 1091.1000 1325.7001 1093.5000 ;
	    RECT 1326.6000 1091.4000 1327.8000 1092.6000 ;
	    RECT 1321.8000 1090.2001 1325.7001 1091.1000 ;
	    RECT 1319.4000 1083.3000 1320.6000 1089.3000 ;
	    RECT 1321.8000 1083.3000 1323.0000 1090.2001 ;
	    RECT 1324.2001 1083.3000 1325.4000 1089.3000 ;
	    RECT 1326.6000 1083.3000 1327.8000 1090.5000 ;
	    RECT 1329.0000 1083.3000 1330.2001 1089.3000 ;
	    RECT 1348.2001 1083.3000 1349.4000 1089.3000 ;
	    RECT 1350.6000 1083.3000 1351.8000 1096.5000 ;
	    RECT 1353.0000 1095.4501 1354.2001 1095.6000 ;
	    RECT 1379.4000 1095.4501 1380.6000 1095.6000 ;
	    RECT 1353.0000 1094.5500 1380.6000 1095.4501 ;
	    RECT 1391.1000 1095.3000 1392.0000 1100.4000 ;
	    RECT 1353.0000 1094.4000 1354.2001 1094.5500 ;
	    RECT 1379.4000 1094.4000 1380.6000 1094.5500 ;
	    RECT 1353.0000 1093.2001 1354.2001 1093.5000 ;
	    RECT 1353.0000 1083.3000 1354.2001 1089.3000 ;
	    RECT 1386.6000 1083.3000 1387.8000 1095.3000 ;
	    RECT 1390.5000 1094.4000 1392.0000 1095.3000 ;
	    RECT 1393.8000 1094.4000 1395.0000 1095.6000 ;
	    RECT 1390.5000 1083.3000 1391.7001 1094.4000 ;
	    RECT 1392.9000 1092.6000 1393.8000 1093.5000 ;
	    RECT 1392.6000 1091.4000 1393.8000 1092.6000 ;
	    RECT 1392.9000 1083.3000 1394.1000 1089.3000 ;
	    RECT 1408.2001 1083.3000 1409.4000 1089.3000 ;
	    RECT 1410.6000 1083.3000 1411.8000 1099.5000 ;
	    RECT 1434.6000 1094.4000 1435.8000 1095.6000 ;
	    RECT 1437.6000 1095.3000 1438.5000 1100.4000 ;
	    RECT 1439.4000 1099.5000 1440.6000 1099.8000 ;
	    RECT 1470.6000 1099.5000 1471.8000 1099.8000 ;
	    RECT 1439.4000 1097.4000 1440.6000 1098.6000 ;
	    RECT 1470.6000 1097.4000 1471.8000 1098.6000 ;
	    RECT 1472.7001 1095.3000 1473.6000 1100.4000 ;
	    RECT 1504.2001 1099.5000 1505.4000 1099.8000 ;
	    RECT 1504.2001 1097.4000 1505.4000 1098.6000 ;
	    RECT 1437.6000 1094.4000 1439.1000 1095.3000 ;
	    RECT 1435.8000 1092.6000 1436.7001 1093.5000 ;
	    RECT 1435.8000 1091.4000 1437.0000 1092.6000 ;
	    RECT 1435.5000 1083.3000 1436.7001 1089.3000 ;
	    RECT 1437.9000 1083.3000 1439.1000 1094.4000 ;
	    RECT 1441.8000 1083.3000 1443.0000 1095.3000 ;
	    RECT 1468.2001 1083.3000 1469.4000 1095.3000 ;
	    RECT 1472.1000 1094.4000 1473.6000 1095.3000 ;
	    RECT 1475.4000 1095.4501 1476.6000 1095.6000 ;
	    RECT 1499.4000 1095.4501 1500.6000 1095.6000 ;
	    RECT 1475.4000 1094.5500 1500.6000 1095.4501 ;
	    RECT 1506.3000 1095.3000 1507.2001 1100.4000 ;
	    RECT 1530.6000 1099.5000 1531.8000 1103.7001 ;
	    RECT 1559.4000 1100.7001 1560.6000 1109.7001 ;
	    RECT 1564.8000 1101.3000 1566.0000 1109.7001 ;
	    RECT 1564.8000 1100.7001 1567.5000 1101.3000 ;
	    RECT 1565.1000 1100.4000 1567.5000 1100.7001 ;
	    RECT 1509.0000 1098.4501 1510.2001 1098.6000 ;
	    RECT 1525.8000 1098.4501 1527.0000 1098.6000 ;
	    RECT 1509.0000 1097.5500 1527.0000 1098.4501 ;
	    RECT 1509.0000 1097.4000 1510.2001 1097.5500 ;
	    RECT 1525.8000 1097.4000 1527.0000 1097.5500 ;
	    RECT 1530.6000 1098.4501 1531.8000 1098.6000 ;
	    RECT 1549.8000 1098.4501 1551.0000 1098.6000 ;
	    RECT 1530.6000 1097.5500 1551.0000 1098.4501 ;
	    RECT 1530.6000 1097.4000 1531.8000 1097.5500 ;
	    RECT 1549.8000 1097.4000 1551.0000 1097.5500 ;
	    RECT 1561.8000 1097.4000 1563.0000 1098.6000 ;
	    RECT 1563.9000 1097.4000 1564.2001 1098.6000 ;
	    RECT 1559.4000 1096.5000 1560.6000 1096.8000 ;
	    RECT 1566.6000 1096.5000 1567.5000 1100.4000 ;
	    RECT 1475.4000 1094.4000 1476.6000 1094.5500 ;
	    RECT 1499.4000 1094.4000 1500.6000 1094.5500 ;
	    RECT 1472.1000 1083.3000 1473.3000 1094.4000 ;
	    RECT 1474.5000 1092.6000 1475.4000 1093.5000 ;
	    RECT 1474.2001 1091.4000 1475.4000 1092.6000 ;
	    RECT 1474.5000 1083.3000 1475.7001 1089.3000 ;
	    RECT 1501.8000 1083.3000 1503.0000 1095.3000 ;
	    RECT 1505.7001 1094.4000 1507.2001 1095.3000 ;
	    RECT 1509.0000 1095.4501 1510.2001 1095.6000 ;
	    RECT 1528.2001 1095.4501 1529.4000 1095.6000 ;
	    RECT 1509.0000 1094.5500 1529.4000 1095.4501 ;
	    RECT 1509.0000 1094.4000 1510.2001 1094.5500 ;
	    RECT 1528.2001 1094.4000 1529.4000 1094.5500 ;
	    RECT 1505.7001 1083.3000 1506.9000 1094.4000 ;
	    RECT 1508.1000 1092.6000 1509.0000 1093.5000 ;
	    RECT 1507.8000 1091.4000 1509.0000 1092.6000 ;
	    RECT 1508.1000 1083.3000 1509.3000 1089.3000 ;
	    RECT 1528.2001 1083.3000 1529.4000 1089.3000 ;
	    RECT 1530.6000 1083.3000 1531.8000 1096.5000 ;
	    RECT 1533.0000 1094.4000 1534.2001 1095.6000 ;
	    RECT 1535.4000 1095.4501 1536.6000 1095.6000 ;
	    RECT 1559.4000 1095.4501 1560.6000 1095.6000 ;
	    RECT 1535.4000 1094.5500 1560.6000 1095.4501 ;
	    RECT 1535.4000 1094.4000 1536.6000 1094.5500 ;
	    RECT 1559.4000 1094.4000 1560.6000 1094.5500 ;
	    RECT 1566.6000 1094.4000 1567.8000 1095.6000 ;
	    RECT 1564.2001 1093.5000 1565.4000 1093.8000 ;
	    RECT 1533.0000 1093.2001 1534.2001 1093.5000 ;
	    RECT 1564.2001 1091.4000 1565.4000 1092.6000 ;
	    RECT 1566.6000 1090.5000 1567.5000 1093.5000 ;
	    RECT 1562.1000 1089.6000 1567.5000 1090.5000 ;
	    RECT 1562.1000 1089.3000 1563.0000 1089.6000 ;
	    RECT 1533.0000 1083.3000 1534.2001 1089.3000 ;
	    RECT 1559.4000 1083.3000 1560.6000 1089.3000 ;
	    RECT 1561.8000 1083.3000 1563.0000 1089.3000 ;
	    RECT 1566.6000 1089.3000 1567.5000 1089.6000 ;
	    RECT 1564.2001 1083.3000 1565.4000 1088.7001 ;
	    RECT 1566.6000 1083.3000 1567.8000 1089.3000 ;
	    RECT 1.2000 1080.6000 1569.0000 1082.4000 ;
	    RECT 124.2000 1073.7001 125.4000 1079.7001 ;
	    RECT 126.6000 1074.6000 127.8000 1079.7001 ;
	    RECT 126.3000 1073.7001 127.8000 1074.6000 ;
	    RECT 129.0000 1073.7001 130.2000 1080.6000 ;
	    RECT 126.3000 1072.8000 127.2000 1073.7001 ;
	    RECT 131.4000 1072.8000 132.6000 1079.7001 ;
	    RECT 133.8000 1073.7001 135.0000 1079.7001 ;
	    RECT 136.2000 1075.5000 137.4000 1079.7001 ;
	    RECT 138.6000 1075.5000 139.8000 1079.7001 ;
	    RECT 124.2000 1071.9000 127.2000 1072.8000 ;
	    RECT 124.2000 1063.5000 125.4000 1071.9000 ;
	    RECT 128.1000 1071.6000 134.4000 1072.8000 ;
	    RECT 141.0000 1072.5000 142.2000 1079.7001 ;
	    RECT 143.4000 1073.7001 144.6000 1079.7001 ;
	    RECT 145.8000 1072.5000 147.0000 1079.7001 ;
	    RECT 148.2000 1073.7001 149.4000 1079.7001 ;
	    RECT 128.1000 1071.0000 129.0000 1071.6000 ;
	    RECT 126.6000 1069.8000 129.0000 1071.0000 ;
	    RECT 133.5000 1070.7001 142.2000 1071.6000 ;
	    RECT 130.5000 1069.8000 132.6000 1070.7001 ;
	    RECT 130.5000 1069.5000 139.8000 1069.8000 ;
	    RECT 131.7000 1068.9000 139.8000 1069.5000 ;
	    RECT 138.6000 1068.6000 139.8000 1068.9000 ;
	    RECT 141.3000 1069.5000 142.2000 1070.7001 ;
	    RECT 143.1000 1070.4000 147.0000 1071.6000 ;
	    RECT 150.6000 1070.4000 151.8000 1079.7001 ;
	    RECT 153.0000 1075.5000 154.2000 1079.7001 ;
	    RECT 155.4000 1075.5000 156.6000 1079.7001 ;
	    RECT 157.8000 1075.5000 159.0000 1079.7001 ;
	    RECT 160.2000 1073.7001 161.4000 1079.7001 ;
	    RECT 155.4000 1071.6000 161.7000 1072.8000 ;
	    RECT 162.6000 1071.6000 163.8000 1079.7001 ;
	    RECT 165.0000 1073.7001 166.2000 1079.7001 ;
	    RECT 167.4000 1072.8000 168.6000 1079.7001 ;
	    RECT 169.8000 1073.7001 171.0000 1079.7001 ;
	    RECT 167.4000 1071.9000 171.3000 1072.8000 ;
	    RECT 172.2000 1072.5000 173.4000 1079.7001 ;
	    RECT 174.6000 1073.7001 175.8000 1079.7001 ;
	    RECT 162.6000 1070.4000 166.5000 1071.6000 ;
	    RECT 153.0000 1069.5000 154.2000 1069.8000 ;
	    RECT 141.3000 1068.6000 154.2000 1069.5000 ;
	    RECT 157.8000 1069.5000 159.0000 1069.8000 ;
	    RECT 170.4000 1069.5000 171.3000 1071.9000 ;
	    RECT 172.2000 1070.4000 173.4000 1071.6000 ;
	    RECT 157.8000 1068.6000 171.3000 1069.5000 ;
	    RECT 129.0000 1067.4000 130.2000 1068.6000 ;
	    RECT 134.1000 1067.7001 135.3000 1068.0000 ;
	    RECT 131.1000 1066.8000 169.5000 1067.7001 ;
	    RECT 168.3000 1066.5000 169.5000 1066.8000 ;
	    RECT 170.4000 1065.9000 171.3000 1068.6000 ;
	    RECT 172.2000 1068.0000 173.4000 1069.5000 ;
	    RECT 172.2000 1066.8000 173.7000 1068.0000 ;
	    RECT 213.0000 1067.7001 214.2000 1079.7001 ;
	    RECT 216.9000 1067.7001 219.9000 1079.7001 ;
	    RECT 222.6000 1067.7001 223.8000 1079.7001 ;
	    RECT 126.3000 1065.0000 132.9000 1065.9000 ;
	    RECT 126.3000 1064.7001 127.5000 1065.0000 ;
	    RECT 133.8000 1064.4000 135.0000 1065.6000 ;
	    RECT 135.9000 1065.0000 161.4000 1065.9000 ;
	    RECT 170.4000 1065.0000 171.6000 1065.9000 ;
	    RECT 160.2000 1064.1000 161.4000 1065.0000 ;
	    RECT 124.2000 1062.3000 137.4000 1063.5000 ;
	    RECT 138.3000 1062.9000 141.3000 1064.1000 ;
	    RECT 147.0000 1062.9000 151.8000 1064.1000 ;
	    RECT 124.2000 1053.3000 125.4000 1062.3000 ;
	    RECT 127.8000 1060.2001 132.3000 1061.4000 ;
	    RECT 131.1000 1059.3000 132.3000 1060.2001 ;
	    RECT 140.1000 1059.3000 141.3000 1062.9000 ;
	    RECT 143.4000 1061.4000 144.6000 1062.6000 ;
	    RECT 151.2000 1061.7001 152.4000 1062.0000 ;
	    RECT 145.8000 1060.8000 152.4000 1061.7001 ;
	    RECT 145.8000 1060.5000 147.0000 1060.8000 ;
	    RECT 143.4000 1060.2001 144.6000 1060.5000 ;
	    RECT 155.4000 1059.6000 156.6000 1063.8000 ;
	    RECT 164.1000 1062.9000 169.8000 1064.1000 ;
	    RECT 164.1000 1061.1000 165.3000 1062.9000 ;
	    RECT 170.7000 1062.0000 171.6000 1065.0000 ;
	    RECT 145.8000 1059.3000 147.0000 1059.6000 ;
	    RECT 129.0000 1053.3000 130.2000 1059.3000 ;
	    RECT 131.1000 1058.1000 135.0000 1059.3000 ;
	    RECT 140.1000 1058.4000 147.0000 1059.3000 ;
	    RECT 148.2000 1058.4000 149.4000 1059.6000 ;
	    RECT 150.3000 1058.4000 150.6000 1059.6000 ;
	    RECT 155.1000 1058.4000 156.6000 1059.6000 ;
	    RECT 162.6000 1060.2001 165.3000 1061.1000 ;
	    RECT 169.8000 1061.1000 171.6000 1062.0000 ;
	    RECT 162.6000 1059.3000 163.8000 1060.2001 ;
	    RECT 133.8000 1053.3000 135.0000 1058.1000 ;
	    RECT 160.2000 1058.1000 163.8000 1059.3000 ;
	    RECT 136.2000 1053.3000 137.4000 1057.5000 ;
	    RECT 138.6000 1053.3000 139.8000 1057.5000 ;
	    RECT 141.0000 1053.3000 142.2000 1057.5000 ;
	    RECT 143.4000 1053.3000 144.6000 1056.3000 ;
	    RECT 145.8000 1053.3000 147.0000 1057.5000 ;
	    RECT 148.2000 1053.3000 149.4000 1056.3000 ;
	    RECT 150.6000 1053.3000 151.8000 1057.5000 ;
	    RECT 153.0000 1053.3000 154.2000 1057.5000 ;
	    RECT 155.4000 1053.3000 156.6000 1057.5000 ;
	    RECT 157.8000 1053.3000 159.0000 1057.5000 ;
	    RECT 160.2000 1053.3000 161.4000 1058.1000 ;
	    RECT 165.0000 1053.3000 166.2000 1059.3000 ;
	    RECT 169.8000 1053.3000 171.0000 1061.1000 ;
	    RECT 172.5000 1060.2001 173.7000 1066.8000 ;
	    RECT 215.4000 1064.4000 216.6000 1065.6000 ;
	    RECT 217.8000 1063.5000 218.7000 1067.7001 ;
	    RECT 220.2000 1064.4000 221.4000 1065.6000 ;
	    RECT 222.6000 1063.5000 223.8000 1063.8000 ;
	    RECT 234.6000 1063.5000 235.8000 1079.7001 ;
	    RECT 237.0000 1073.7001 238.2000 1079.7001 ;
	    RECT 256.2000 1067.7001 257.4000 1079.7001 ;
	    RECT 258.6000 1069.5000 259.8000 1079.7001 ;
	    RECT 261.0000 1068.6000 262.2000 1079.7001 ;
	    RECT 258.9000 1067.7001 262.2000 1068.6000 ;
	    RECT 280.2000 1067.7001 281.4000 1079.7001 ;
	    RECT 284.1000 1068.9000 285.3000 1079.7001 ;
	    RECT 304.2000 1073.7001 305.4000 1079.7001 ;
	    RECT 304.2000 1069.5000 305.4000 1069.8000 ;
	    RECT 282.6000 1067.7001 285.3000 1068.9000 ;
	    RECT 256.2000 1064.4000 257.1000 1067.7001 ;
	    RECT 258.9000 1066.8000 259.8000 1067.7001 ;
	    RECT 258.0000 1065.6000 259.8000 1066.8000 ;
	    RECT 256.2000 1063.5000 257.4000 1064.4000 ;
	    RECT 215.4000 1063.2001 216.6000 1063.5000 ;
	    RECT 220.2000 1063.2001 221.4000 1063.5000 ;
	    RECT 196.2000 1062.4501 197.4000 1062.6000 ;
	    RECT 213.0000 1062.4501 214.2000 1062.6000 ;
	    RECT 196.2000 1061.5500 214.2000 1062.4501 ;
	    RECT 196.2000 1061.4000 197.4000 1061.5500 ;
	    RECT 213.0000 1061.4000 214.2000 1061.5500 ;
	    RECT 215.1000 1060.8000 215.4000 1062.3000 ;
	    RECT 217.8000 1061.4000 219.0000 1062.6000 ;
	    RECT 219.9000 1061.4000 221.4000 1062.3000 ;
	    RECT 222.6000 1061.4000 223.8000 1062.6000 ;
	    RECT 227.4000 1062.4501 228.6000 1062.6000 ;
	    RECT 234.6000 1062.4501 235.8000 1062.6000 ;
	    RECT 227.4000 1061.5500 235.8000 1062.4501 ;
	    RECT 227.4000 1061.4000 228.6000 1061.5500 ;
	    RECT 234.6000 1061.4000 235.8000 1061.5500 ;
	    RECT 256.2000 1061.4000 257.4000 1062.6000 ;
	    RECT 172.2000 1059.0000 173.7000 1060.2001 ;
	    RECT 213.3000 1059.3000 218.7000 1059.9000 ;
	    RECT 220.5000 1059.3000 221.4000 1061.4000 ;
	    RECT 258.9000 1061.1000 259.8000 1065.6000 ;
	    RECT 261.0000 1064.4000 262.2000 1065.6000 ;
	    RECT 282.9000 1063.5000 283.8000 1067.7001 ;
	    RECT 304.2000 1067.4000 305.4000 1068.6000 ;
	    RECT 285.0000 1066.5000 286.2000 1066.8000 ;
	    RECT 306.6000 1066.5000 307.8000 1079.7001 ;
	    RECT 309.0000 1073.7001 310.2000 1079.7001 ;
	    RECT 328.2000 1073.7001 329.4000 1079.7001 ;
	    RECT 330.6000 1066.5000 331.8000 1079.7001 ;
	    RECT 333.0000 1073.7001 334.2000 1079.7001 ;
	    RECT 345.0000 1073.7001 346.2000 1079.7001 ;
	    RECT 333.0000 1069.5000 334.2000 1069.8000 ;
	    RECT 333.0000 1068.4501 334.2000 1068.6000 ;
	    RECT 335.4000 1068.4501 336.6000 1068.6000 ;
	    RECT 333.0000 1067.5500 336.6000 1068.4501 ;
	    RECT 333.0000 1067.4000 334.2000 1067.5500 ;
	    RECT 335.4000 1067.4000 336.6000 1067.5500 ;
	    RECT 285.0000 1065.4501 286.2000 1065.6000 ;
	    RECT 304.2000 1065.4501 305.4000 1065.6000 ;
	    RECT 285.0000 1064.5500 305.4000 1065.4501 ;
	    RECT 285.0000 1064.4000 286.2000 1064.5500 ;
	    RECT 304.2000 1064.4000 305.4000 1064.5500 ;
	    RECT 306.6000 1065.4501 307.8000 1065.6000 ;
	    RECT 328.2000 1065.4501 329.4000 1065.6000 ;
	    RECT 306.6000 1064.5500 329.4000 1065.4501 ;
	    RECT 306.6000 1064.4000 307.8000 1064.5500 ;
	    RECT 328.2000 1064.4000 329.4000 1064.5500 ;
	    RECT 330.6000 1065.4501 331.8000 1065.6000 ;
	    RECT 333.0000 1065.4501 334.2000 1065.6000 ;
	    RECT 330.6000 1064.5500 334.2000 1065.4501 ;
	    RECT 330.6000 1064.4000 331.8000 1064.5500 ;
	    RECT 333.0000 1064.4000 334.2000 1064.5500 ;
	    RECT 347.4000 1063.5000 348.6000 1079.7001 ;
	    RECT 373.8000 1067.7001 375.0000 1079.7001 ;
	    RECT 377.7000 1068.6000 378.9000 1079.7001 ;
	    RECT 380.1000 1073.7001 381.3000 1079.7001 ;
	    RECT 515.4000 1073.7001 516.6000 1079.7001 ;
	    RECT 517.8000 1072.5000 519.0000 1079.7001 ;
	    RECT 520.2000 1073.7001 521.4000 1079.7001 ;
	    RECT 522.6000 1072.8000 523.8000 1079.7001 ;
	    RECT 525.0000 1073.7001 526.2000 1079.7001 ;
	    RECT 519.9000 1071.9000 523.8000 1072.8000 ;
	    RECT 379.8000 1070.4000 381.0000 1071.6000 ;
	    RECT 385.8000 1071.4501 387.0000 1071.6000 ;
	    RECT 517.8000 1071.4501 519.0000 1071.6000 ;
	    RECT 385.8000 1070.5500 519.0000 1071.4501 ;
	    RECT 385.8000 1070.4000 387.0000 1070.5500 ;
	    RECT 517.8000 1070.4000 519.0000 1070.5500 ;
	    RECT 380.1000 1069.5000 381.0000 1070.4000 ;
	    RECT 519.9000 1069.5000 520.8000 1071.9000 ;
	    RECT 527.4000 1071.6000 528.6000 1079.7001 ;
	    RECT 529.8000 1073.7001 531.0000 1079.7001 ;
	    RECT 532.2000 1075.5000 533.4000 1079.7001 ;
	    RECT 534.6000 1075.5000 535.8000 1079.7001 ;
	    RECT 537.0000 1075.5000 538.2000 1079.7001 ;
	    RECT 529.5000 1071.6000 535.8000 1072.8000 ;
	    RECT 524.7000 1070.4000 528.6000 1071.6000 ;
	    RECT 539.4000 1070.4000 540.6000 1079.7001 ;
	    RECT 541.8000 1073.7001 543.0000 1079.7001 ;
	    RECT 544.2000 1072.5000 545.4000 1079.7001 ;
	    RECT 546.6000 1073.7001 547.8000 1079.7001 ;
	    RECT 549.0000 1072.5000 550.2000 1079.7001 ;
	    RECT 551.4000 1075.5000 552.6000 1079.7001 ;
	    RECT 553.8000 1075.5000 555.0000 1079.7001 ;
	    RECT 556.2000 1073.7001 557.4000 1079.7001 ;
	    RECT 558.6000 1072.8000 559.8000 1079.7001 ;
	    RECT 561.0000 1073.7001 562.2000 1080.6000 ;
	    RECT 563.4000 1074.6000 564.6000 1079.7001 ;
	    RECT 563.4000 1073.7001 564.9000 1074.6000 ;
	    RECT 565.8000 1073.7001 567.0000 1079.7001 ;
	    RECT 585.0000 1073.7001 586.2000 1079.7001 ;
	    RECT 564.0000 1072.8000 564.9000 1073.7001 ;
	    RECT 556.8000 1071.6000 563.1000 1072.8000 ;
	    RECT 564.0000 1071.9000 567.0000 1072.8000 ;
	    RECT 544.2000 1070.4000 548.1000 1071.6000 ;
	    RECT 549.0000 1070.7001 557.7000 1071.6000 ;
	    RECT 562.2000 1071.0000 563.1000 1071.6000 ;
	    RECT 532.2000 1069.5000 533.4000 1069.8000 ;
	    RECT 377.7000 1067.7001 379.2000 1068.6000 ;
	    RECT 376.2000 1065.4501 377.4000 1065.6000 ;
	    RECT 371.5500 1064.5500 377.4000 1065.4501 ;
	    RECT 261.0000 1063.2001 262.2000 1063.5000 ;
	    RECT 282.6000 1062.4501 283.8000 1062.6000 ;
	    RECT 294.6000 1062.4501 295.8000 1062.6000 ;
	    RECT 282.6000 1061.5500 295.8000 1062.4501 ;
	    RECT 282.6000 1061.4000 283.8000 1061.5500 ;
	    RECT 294.6000 1061.4000 295.8000 1061.5500 ;
	    RECT 213.0000 1059.0000 219.0000 1059.3000 ;
	    RECT 172.2000 1053.3000 173.4000 1059.0000 ;
	    RECT 174.6000 1053.3000 175.8000 1056.3000 ;
	    RECT 213.0000 1053.3000 214.2000 1059.0000 ;
	    RECT 215.4000 1053.3000 216.6000 1058.1000 ;
	    RECT 217.8000 1054.2001 219.0000 1059.0000 ;
	    RECT 220.2000 1055.1000 221.4000 1059.3000 ;
	    RECT 222.6000 1054.2001 223.8000 1059.3000 ;
	    RECT 217.8000 1053.3000 223.8000 1054.2001 ;
	    RECT 234.6000 1053.3000 235.8000 1060.5000 ;
	    RECT 237.0000 1059.4501 238.2000 1059.6000 ;
	    RECT 239.4000 1059.4501 240.6000 1059.6000 ;
	    RECT 237.0000 1058.5500 240.6000 1059.4501 ;
	    RECT 237.0000 1058.4000 238.2000 1058.5500 ;
	    RECT 239.4000 1058.4000 240.6000 1058.5500 ;
	    RECT 237.0000 1057.2001 238.2000 1057.5000 ;
	    RECT 237.0000 1053.3000 238.2000 1056.3000 ;
	    RECT 256.2000 1053.3000 257.4000 1060.5000 ;
	    RECT 258.9000 1060.2001 262.2000 1061.1000 ;
	    RECT 258.6000 1053.3000 259.8000 1059.3000 ;
	    RECT 261.0000 1053.3000 262.2000 1060.2001 ;
	    RECT 268.2000 1059.4501 269.4000 1059.6000 ;
	    RECT 280.2000 1059.4501 281.4000 1059.6000 ;
	    RECT 268.2000 1058.5500 281.4000 1059.4501 ;
	    RECT 268.2000 1058.4000 269.4000 1058.5500 ;
	    RECT 280.2000 1058.4000 281.4000 1058.5500 ;
	    RECT 280.2000 1057.2001 281.4000 1057.5000 ;
	    RECT 282.9000 1056.3000 283.8000 1060.5000 ;
	    RECT 306.6000 1059.3000 307.8000 1063.5000 ;
	    RECT 309.0000 1062.4501 310.2000 1062.6000 ;
	    RECT 311.4000 1062.4501 312.6000 1062.6000 ;
	    RECT 328.2000 1062.4501 329.4000 1062.6000 ;
	    RECT 309.0000 1061.5500 329.4000 1062.4501 ;
	    RECT 309.0000 1061.4000 310.2000 1061.5500 ;
	    RECT 311.4000 1061.4000 312.6000 1061.5500 ;
	    RECT 328.2000 1061.4000 329.4000 1061.5500 ;
	    RECT 309.0000 1060.2001 310.2000 1060.5000 ;
	    RECT 328.2000 1060.2001 329.4000 1060.5000 ;
	    RECT 330.6000 1059.3000 331.8000 1063.5000 ;
	    RECT 347.4000 1062.4501 348.6000 1062.6000 ;
	    RECT 371.5500 1062.4501 372.4500 1064.5500 ;
	    RECT 376.2000 1064.4000 377.4000 1064.5500 ;
	    RECT 376.2000 1063.2001 377.4000 1063.5000 ;
	    RECT 378.3000 1062.6000 379.2000 1067.7001 ;
	    RECT 381.0000 1067.4000 382.2000 1068.6000 ;
	    RECT 517.8000 1068.0000 519.0000 1069.5000 ;
	    RECT 517.5000 1066.8000 519.0000 1068.0000 ;
	    RECT 519.9000 1068.6000 533.4000 1069.5000 ;
	    RECT 537.0000 1069.5000 538.2000 1069.8000 ;
	    RECT 549.0000 1069.5000 549.9000 1070.7001 ;
	    RECT 558.6000 1069.8000 560.7000 1070.7001 ;
	    RECT 562.2000 1069.8000 564.6000 1071.0000 ;
	    RECT 537.0000 1068.6000 549.9000 1069.5000 ;
	    RECT 551.4000 1069.5000 560.7000 1069.8000 ;
	    RECT 551.4000 1068.9000 559.5000 1069.5000 ;
	    RECT 551.4000 1068.6000 552.6000 1068.9000 ;
	    RECT 347.4000 1061.5500 372.4500 1062.4501 ;
	    RECT 347.4000 1061.4000 348.6000 1061.5500 ;
	    RECT 373.8000 1061.4000 375.0000 1062.6000 ;
	    RECT 375.9000 1060.8000 376.2000 1062.3000 ;
	    RECT 378.3000 1061.4000 380.1000 1062.6000 ;
	    RECT 381.0000 1062.4501 382.2000 1062.6000 ;
	    RECT 467.4000 1062.4501 468.6000 1062.6000 ;
	    RECT 381.0000 1061.5500 468.6000 1062.4501 ;
	    RECT 381.0000 1061.4000 382.2000 1061.5500 ;
	    RECT 467.4000 1061.4000 468.6000 1061.5500 ;
	    RECT 337.8000 1059.4501 339.0000 1059.6000 ;
	    RECT 345.0000 1059.4501 346.2000 1059.6000 ;
	    RECT 305.1000 1058.4000 307.8000 1059.3000 ;
	    RECT 280.2000 1053.3000 281.4000 1056.3000 ;
	    RECT 282.6000 1053.3000 283.8000 1056.3000 ;
	    RECT 285.0000 1053.3000 286.2000 1056.3000 ;
	    RECT 305.1000 1053.3000 306.3000 1058.4000 ;
	    RECT 309.0000 1053.3000 310.2000 1059.3000 ;
	    RECT 328.2000 1053.3000 329.4000 1059.3000 ;
	    RECT 330.6000 1058.4000 333.3000 1059.3000 ;
	    RECT 337.8000 1058.5500 346.2000 1059.4501 ;
	    RECT 337.8000 1058.4000 339.0000 1058.5500 ;
	    RECT 345.0000 1058.4000 346.2000 1058.5500 ;
	    RECT 332.1000 1053.3000 333.3000 1058.4000 ;
	    RECT 345.0000 1057.2001 346.2000 1057.5000 ;
	    RECT 345.0000 1053.3000 346.2000 1056.3000 ;
	    RECT 347.4000 1053.3000 348.6000 1060.5000 ;
	    RECT 374.1000 1059.3000 379.5000 1059.9000 ;
	    RECT 381.0000 1059.3000 381.9000 1060.5000 ;
	    RECT 517.5000 1060.2001 518.7000 1066.8000 ;
	    RECT 519.9000 1065.9000 520.8000 1068.6000 ;
	    RECT 555.9000 1067.7001 557.1000 1068.0000 ;
	    RECT 521.7000 1066.8000 560.1000 1067.7001 ;
	    RECT 561.0000 1067.4000 562.2000 1068.6000 ;
	    RECT 521.7000 1066.5000 522.9000 1066.8000 ;
	    RECT 519.6000 1065.0000 520.8000 1065.9000 ;
	    RECT 529.8000 1065.0000 555.3000 1065.9000 ;
	    RECT 519.6000 1062.0000 520.5000 1065.0000 ;
	    RECT 529.8000 1064.1000 531.0000 1065.0000 ;
	    RECT 556.2000 1064.4000 557.4000 1065.6000 ;
	    RECT 558.3000 1065.0000 564.9000 1065.9000 ;
	    RECT 563.7000 1064.7001 564.9000 1065.0000 ;
	    RECT 521.4000 1062.9000 527.1000 1064.1000 ;
	    RECT 519.6000 1061.1000 521.4000 1062.0000 ;
	    RECT 373.8000 1059.0000 379.8000 1059.3000 ;
	    RECT 373.8000 1053.3000 375.0000 1059.0000 ;
	    RECT 376.2000 1053.3000 377.4000 1058.1000 ;
	    RECT 378.6000 1053.3000 379.8000 1059.0000 ;
	    RECT 381.0000 1053.3000 382.2000 1059.3000 ;
	    RECT 517.5000 1059.0000 519.0000 1060.2001 ;
	    RECT 515.4000 1053.3000 516.6000 1056.3000 ;
	    RECT 517.8000 1053.3000 519.0000 1059.0000 ;
	    RECT 520.2000 1053.3000 521.4000 1061.1000 ;
	    RECT 525.9000 1061.1000 527.1000 1062.9000 ;
	    RECT 525.9000 1060.2001 528.6000 1061.1000 ;
	    RECT 527.4000 1059.3000 528.6000 1060.2001 ;
	    RECT 534.6000 1059.6000 535.8000 1063.8000 ;
	    RECT 539.4000 1062.9000 544.2000 1064.1000 ;
	    RECT 549.9000 1062.9000 552.9000 1064.1000 ;
	    RECT 565.8000 1063.5000 567.0000 1071.9000 ;
	    RECT 585.0000 1069.5000 586.2000 1069.8000 ;
	    RECT 573.0000 1068.4501 574.2000 1068.6000 ;
	    RECT 585.0000 1068.4501 586.2000 1068.6000 ;
	    RECT 573.0000 1067.5500 586.2000 1068.4501 ;
	    RECT 573.0000 1067.4000 574.2000 1067.5500 ;
	    RECT 585.0000 1067.4000 586.2000 1067.5500 ;
	    RECT 587.4000 1066.5000 588.6000 1079.7001 ;
	    RECT 589.8000 1073.7001 591.0000 1079.7001 ;
	    RECT 594.6000 1079.4000 595.8000 1080.6000 ;
	    RECT 601.8000 1073.7001 603.0000 1079.7001 ;
	    RECT 587.4000 1065.4501 588.6000 1065.6000 ;
	    RECT 592.2000 1065.4501 593.4000 1065.6000 ;
	    RECT 587.4000 1064.5500 593.4000 1065.4501 ;
	    RECT 587.4000 1064.4000 588.6000 1064.5500 ;
	    RECT 592.2000 1064.4000 593.4000 1064.5500 ;
	    RECT 604.2000 1063.5000 605.4000 1079.7001 ;
	    RECT 624.3000 1068.9000 625.5000 1079.7001 ;
	    RECT 624.3000 1067.7001 627.0000 1068.9000 ;
	    RECT 628.2000 1067.7001 629.4000 1079.7001 ;
	    RECT 647.4000 1073.7001 648.6000 1079.7001 ;
	    RECT 647.4000 1069.5000 648.6000 1069.8000 ;
	    RECT 635.4000 1068.4501 636.6000 1068.6000 ;
	    RECT 647.4000 1068.4501 648.6000 1068.6000 ;
	    RECT 623.4000 1066.5000 624.6000 1066.8000 ;
	    RECT 623.4000 1064.4000 624.6000 1065.6000 ;
	    RECT 538.8000 1061.7001 540.0000 1062.0000 ;
	    RECT 538.8000 1060.8000 545.4000 1061.7001 ;
	    RECT 546.6000 1061.4000 547.8000 1062.6000 ;
	    RECT 544.2000 1060.5000 545.4000 1060.8000 ;
	    RECT 546.6000 1060.2001 547.8000 1060.5000 ;
	    RECT 525.0000 1053.3000 526.2000 1059.3000 ;
	    RECT 527.4000 1058.1000 531.0000 1059.3000 ;
	    RECT 534.6000 1058.4000 536.1000 1059.6000 ;
	    RECT 540.6000 1058.4000 540.9000 1059.6000 ;
	    RECT 541.8000 1058.4000 543.0000 1059.6000 ;
	    RECT 544.2000 1059.3000 545.4000 1059.6000 ;
	    RECT 549.9000 1059.3000 551.1000 1062.9000 ;
	    RECT 553.8000 1062.3000 567.0000 1063.5000 ;
	    RECT 558.9000 1060.2001 563.4000 1061.4000 ;
	    RECT 558.9000 1059.3000 560.1000 1060.2001 ;
	    RECT 544.2000 1058.4000 551.1000 1059.3000 ;
	    RECT 529.8000 1053.3000 531.0000 1058.1000 ;
	    RECT 556.2000 1058.1000 560.1000 1059.3000 ;
	    RECT 532.2000 1053.3000 533.4000 1057.5000 ;
	    RECT 534.6000 1053.3000 535.8000 1057.5000 ;
	    RECT 537.0000 1053.3000 538.2000 1057.5000 ;
	    RECT 539.4000 1053.3000 540.6000 1057.5000 ;
	    RECT 541.8000 1053.3000 543.0000 1056.3000 ;
	    RECT 544.2000 1053.3000 545.4000 1057.5000 ;
	    RECT 546.6000 1053.3000 547.8000 1056.3000 ;
	    RECT 549.0000 1053.3000 550.2000 1057.5000 ;
	    RECT 551.4000 1053.3000 552.6000 1057.5000 ;
	    RECT 553.8000 1053.3000 555.0000 1057.5000 ;
	    RECT 556.2000 1053.3000 557.4000 1058.1000 ;
	    RECT 561.0000 1053.3000 562.2000 1059.3000 ;
	    RECT 565.8000 1053.3000 567.0000 1062.3000 ;
	    RECT 587.4000 1059.3000 588.6000 1063.5000 ;
	    RECT 589.8000 1062.4501 591.0000 1062.6000 ;
	    RECT 594.6000 1062.4501 595.8000 1062.6000 ;
	    RECT 589.8000 1061.5500 595.8000 1062.4501 ;
	    RECT 589.8000 1061.4000 591.0000 1061.5500 ;
	    RECT 594.6000 1061.4000 595.8000 1061.5500 ;
	    RECT 604.2000 1062.4501 605.4000 1062.6000 ;
	    RECT 623.5500 1062.4501 624.4500 1064.4000 ;
	    RECT 625.8000 1063.5000 626.7000 1067.7001 ;
	    RECT 635.4000 1067.5500 648.6000 1068.4501 ;
	    RECT 635.4000 1067.4000 636.6000 1067.5500 ;
	    RECT 647.4000 1067.4000 648.6000 1067.5500 ;
	    RECT 649.8000 1066.5000 651.0000 1079.7001 ;
	    RECT 652.2000 1073.7001 653.4000 1079.7001 ;
	    RECT 637.8000 1065.4501 639.0000 1065.6000 ;
	    RECT 649.8000 1065.4501 651.0000 1065.6000 ;
	    RECT 637.8000 1064.5500 651.0000 1065.4501 ;
	    RECT 637.8000 1064.4000 639.0000 1064.5500 ;
	    RECT 649.8000 1064.4000 651.0000 1064.5500 ;
	    RECT 673.8000 1063.5000 675.0000 1079.7001 ;
	    RECT 676.2000 1073.7001 677.4000 1079.7001 ;
	    RECT 745.8000 1067.1000 747.0000 1079.7001 ;
	    RECT 748.2000 1068.0000 749.4000 1079.7001 ;
	    RECT 752.4000 1074.6000 753.6000 1079.7001 ;
	    RECT 750.6000 1073.7001 753.6000 1074.6000 ;
	    RECT 756.6000 1073.7001 757.8000 1079.7001 ;
	    RECT 759.0000 1073.7001 760.2000 1079.7001 ;
	    RECT 761.4000 1073.7001 762.6000 1079.7001 ;
	    RECT 765.3000 1073.7001 767.1000 1079.7001 ;
	    RECT 750.6000 1072.5000 751.8000 1073.7001 ;
	    RECT 759.0000 1072.8000 759.9000 1073.7001 ;
	    RECT 755.7000 1071.9000 761.1000 1072.8000 ;
	    RECT 765.0000 1072.5000 766.2000 1073.7001 ;
	    RECT 755.7000 1071.6000 756.9000 1071.9000 ;
	    RECT 759.9000 1071.6000 761.1000 1071.9000 ;
	    RECT 750.6000 1069.5000 751.8000 1069.8000 ;
	    RECT 757.5000 1069.5000 758.7000 1069.8000 ;
	    RECT 750.6000 1068.6000 758.7000 1069.5000 ;
	    RECT 759.6000 1069.5000 762.9000 1070.4000 ;
	    RECT 759.6000 1067.7001 760.5000 1069.5000 ;
	    RECT 761.7000 1069.2001 762.9000 1069.5000 ;
	    RECT 765.3000 1069.8000 767.4000 1071.0000 ;
	    RECT 765.3000 1068.3000 766.2000 1069.8000 ;
	    RECT 753.3000 1067.1000 760.5000 1067.7001 ;
	    RECT 745.8000 1066.8000 760.5000 1067.1000 ;
	    RECT 762.6000 1067.4000 766.2000 1068.3000 ;
	    RECT 769.8000 1067.7001 771.0000 1079.7001 ;
	    RECT 745.8000 1066.5000 754.5000 1066.8000 ;
	    RECT 745.8000 1066.2001 754.2000 1066.5000 ;
	    RECT 749.1000 1064.4000 754.5000 1065.3000 ;
	    RECT 755.4000 1064.4000 756.6000 1065.6000 ;
	    RECT 749.1000 1064.1000 750.3000 1064.4000 ;
	    RECT 604.2000 1061.5500 624.4500 1062.4501 ;
	    RECT 604.2000 1061.4000 605.4000 1061.5500 ;
	    RECT 625.8000 1061.4000 627.0000 1062.6000 ;
	    RECT 589.8000 1060.2001 591.0000 1060.5000 ;
	    RECT 585.9000 1058.4000 588.6000 1059.3000 ;
	    RECT 585.9000 1053.3000 587.1000 1058.4000 ;
	    RECT 589.8000 1053.3000 591.0000 1059.3000 ;
	    RECT 601.8000 1058.4000 603.0000 1059.6000 ;
	    RECT 601.8000 1057.2001 603.0000 1057.5000 ;
	    RECT 601.8000 1053.3000 603.0000 1056.3000 ;
	    RECT 604.2000 1053.3000 605.4000 1060.5000 ;
	    RECT 625.8000 1056.3000 626.7000 1060.5000 ;
	    RECT 628.2000 1058.4000 629.4000 1059.6000 ;
	    RECT 649.8000 1059.3000 651.0000 1063.5000 ;
	    RECT 751.5000 1062.6000 752.7000 1062.9000 ;
	    RECT 762.6000 1062.6000 763.5000 1067.4000 ;
	    RECT 772.2000 1066.8000 773.4000 1079.7001 ;
	    RECT 774.6000 1079.4000 775.8000 1080.6000 ;
	    RECT 791.4000 1073.7001 792.6000 1079.7001 ;
	    RECT 767.1000 1066.5000 773.4000 1066.8000 ;
	    RECT 793.8000 1066.5000 795.0000 1079.7001 ;
	    RECT 796.2000 1073.7001 797.4000 1079.7001 ;
	    RECT 796.2000 1069.5000 797.4000 1069.8000 ;
	    RECT 796.2000 1067.4000 797.4000 1068.6000 ;
	    RECT 815.4000 1067.7001 816.6000 1079.7001 ;
	    RECT 819.3000 1068.9000 820.5000 1079.7001 ;
	    RECT 817.8000 1067.7001 820.5000 1068.9000 ;
	    RECT 849.0000 1067.7001 850.2000 1079.7001 ;
	    RECT 852.9000 1067.7001 855.9000 1079.7001 ;
	    RECT 858.6000 1067.7001 859.8000 1079.7001 ;
	    RECT 767.1000 1065.9000 771.3000 1066.5000 ;
	    RECT 767.1000 1065.6000 768.3000 1065.9000 ;
	    RECT 769.5000 1064.7001 770.7000 1065.0000 ;
	    RECT 765.0000 1063.8000 770.7000 1064.7001 ;
	    RECT 772.2000 1064.4000 773.4000 1065.6000 ;
	    RECT 793.8000 1064.4000 795.0000 1065.6000 ;
	    RECT 765.0000 1063.5000 766.2000 1063.8000 ;
	    RECT 818.1000 1063.5000 819.0000 1067.7001 ;
	    RECT 820.2000 1066.5000 821.4000 1066.8000 ;
	    RECT 820.2000 1065.4501 821.4000 1065.6000 ;
	    RECT 846.6000 1065.4501 847.8000 1065.6000 ;
	    RECT 820.2000 1064.5500 847.8000 1065.4501 ;
	    RECT 820.2000 1064.4000 821.4000 1064.5500 ;
	    RECT 846.6000 1064.4000 847.8000 1064.5500 ;
	    RECT 851.4000 1064.4000 852.6000 1065.6000 ;
	    RECT 853.8000 1063.5000 854.7000 1067.7001 ;
	    RECT 856.2000 1064.4000 857.4000 1065.6000 ;
	    RECT 858.6000 1063.5000 859.8000 1063.8000 ;
	    RECT 870.6000 1063.5000 871.8000 1079.7001 ;
	    RECT 873.0000 1073.7001 874.2000 1079.7001 ;
	    RECT 907.5000 1073.7001 908.7000 1079.7001 ;
	    RECT 907.8000 1070.4000 909.0000 1071.6000 ;
	    RECT 907.8000 1069.5000 908.7000 1070.4000 ;
	    RECT 909.9000 1068.6000 911.1000 1079.7001 ;
	    RECT 906.6000 1067.4000 907.8000 1068.6000 ;
	    RECT 909.6000 1067.7001 911.1000 1068.6000 ;
	    RECT 913.8000 1067.7001 915.0000 1079.7001 ;
	    RECT 933.9000 1068.9000 935.1000 1079.7001 ;
	    RECT 933.9000 1067.7001 936.6000 1068.9000 ;
	    RECT 937.8000 1067.7001 939.0000 1079.7001 ;
	    RECT 940.2000 1077.4501 941.4000 1077.6000 ;
	    RECT 1005.0000 1077.4501 1006.2000 1077.6000 ;
	    RECT 940.2000 1076.5500 1006.2000 1077.4501 ;
	    RECT 940.2000 1076.4000 941.4000 1076.5500 ;
	    RECT 1005.0000 1076.4000 1006.2000 1076.5500 ;
	    RECT 1062.6000 1073.7001 1063.8000 1079.7001 ;
	    RECT 1065.0000 1074.6000 1066.2001 1079.7001 ;
	    RECT 1064.7001 1073.7001 1066.2001 1074.6000 ;
	    RECT 1067.4000 1073.7001 1068.6000 1080.6000 ;
	    RECT 1064.7001 1072.8000 1065.6000 1073.7001 ;
	    RECT 1069.8000 1072.8000 1071.0000 1079.7001 ;
	    RECT 1072.2001 1073.7001 1073.4000 1079.7001 ;
	    RECT 1074.6000 1075.5000 1075.8000 1079.7001 ;
	    RECT 1077.0000 1075.5000 1078.2001 1079.7001 ;
	    RECT 1062.6000 1071.9000 1065.6000 1072.8000 ;
	    RECT 652.2000 1062.4501 653.4000 1062.6000 ;
	    RECT 673.8000 1062.4501 675.0000 1062.6000 ;
	    RECT 652.2000 1061.5500 675.0000 1062.4501 ;
	    RECT 652.2000 1061.4000 653.4000 1061.5500 ;
	    RECT 673.8000 1061.4000 675.0000 1061.5500 ;
	    RECT 747.0000 1061.4000 747.3000 1062.6000 ;
	    RECT 748.2000 1061.4000 749.4000 1062.6000 ;
	    RECT 750.3000 1061.7001 763.5000 1062.6000 ;
	    RECT 652.2000 1060.2001 653.4000 1060.5000 ;
	    RECT 648.3000 1058.4000 651.0000 1059.3000 ;
	    RECT 628.2000 1057.2001 629.4000 1057.5000 ;
	    RECT 623.4000 1053.3000 624.6000 1056.3000 ;
	    RECT 625.8000 1053.3000 627.0000 1056.3000 ;
	    RECT 628.2000 1053.3000 629.4000 1056.3000 ;
	    RECT 648.3000 1053.3000 649.5000 1058.4000 ;
	    RECT 652.2000 1053.3000 653.4000 1059.3000 ;
	    RECT 673.8000 1053.3000 675.0000 1060.5000 ;
	    RECT 676.2000 1058.4000 677.4000 1059.6000 ;
	    RECT 676.2000 1057.2001 677.4000 1057.5000 ;
	    RECT 676.2000 1053.3000 677.4000 1056.3000 ;
	    RECT 745.8000 1053.3000 747.0000 1060.5000 ;
	    RECT 748.2000 1053.3000 749.4000 1059.3000 ;
	    RECT 753.3000 1058.4000 754.2000 1061.7001 ;
	    RECT 761.7000 1061.4000 762.9000 1061.7001 ;
	    RECT 772.2000 1060.8000 773.4000 1063.5000 ;
	    RECT 789.0000 1062.4501 790.2000 1062.6000 ;
	    RECT 791.4000 1062.4501 792.6000 1062.6000 ;
	    RECT 789.0000 1061.5500 792.6000 1062.4501 ;
	    RECT 789.0000 1061.4000 790.2000 1061.5500 ;
	    RECT 791.4000 1061.4000 792.6000 1061.5500 ;
	    RECT 767.7000 1059.9000 773.4000 1060.8000 ;
	    RECT 791.4000 1060.2001 792.6000 1060.5000 ;
	    RECT 767.7000 1059.6000 768.9000 1059.9000 ;
	    RECT 750.6000 1056.3000 751.8000 1057.5000 ;
	    RECT 753.0000 1057.2001 754.2000 1058.4000 ;
	    RECT 755.7000 1058.1000 756.9000 1058.4000 ;
	    RECT 755.7000 1057.2001 759.9000 1058.1000 ;
	    RECT 759.0000 1056.3000 759.9000 1057.2001 ;
	    RECT 765.0000 1056.3000 766.2000 1057.5000 ;
	    RECT 750.6000 1055.4000 753.6000 1056.3000 ;
	    RECT 752.4000 1053.3000 753.6000 1055.4000 ;
	    RECT 756.3000 1053.3000 757.8000 1056.3000 ;
	    RECT 759.0000 1053.3000 760.2000 1056.3000 ;
	    RECT 761.4000 1053.3000 762.6000 1056.3000 ;
	    RECT 765.0000 1055.4000 767.1000 1056.3000 ;
	    RECT 765.3000 1053.3000 767.1000 1055.4000 ;
	    RECT 769.8000 1053.3000 771.0000 1059.0000 ;
	    RECT 772.2000 1053.3000 773.4000 1059.9000 ;
	    RECT 793.8000 1059.3000 795.0000 1063.5000 ;
	    RECT 851.4000 1063.2001 852.6000 1063.5000 ;
	    RECT 856.2000 1063.2001 857.4000 1063.5000 ;
	    RECT 909.6000 1062.6000 910.5000 1067.7001 ;
	    RECT 933.0000 1066.5000 934.2000 1066.8000 ;
	    RECT 911.4000 1064.4000 912.6000 1065.6000 ;
	    RECT 923.4000 1065.4501 924.6000 1065.6000 ;
	    RECT 933.0000 1065.4501 934.2000 1065.6000 ;
	    RECT 923.4000 1064.5500 934.2000 1065.4501 ;
	    RECT 923.4000 1064.4000 924.6000 1064.5500 ;
	    RECT 933.0000 1064.4000 934.2000 1064.5500 ;
	    RECT 935.4000 1063.5000 936.3000 1067.7001 ;
	    RECT 1062.6000 1063.5000 1063.8000 1071.9000 ;
	    RECT 1066.5000 1071.6000 1072.8000 1072.8000 ;
	    RECT 1079.4000 1072.5000 1080.6000 1079.7001 ;
	    RECT 1081.8000 1073.7001 1083.0000 1079.7001 ;
	    RECT 1084.2001 1072.5000 1085.4000 1079.7001 ;
	    RECT 1086.6000 1073.7001 1087.8000 1079.7001 ;
	    RECT 1066.5000 1071.0000 1067.4000 1071.6000 ;
	    RECT 1065.0000 1069.8000 1067.4000 1071.0000 ;
	    RECT 1071.9000 1070.7001 1080.6000 1071.6000 ;
	    RECT 1068.9000 1069.8000 1071.0000 1070.7001 ;
	    RECT 1068.9000 1069.5000 1078.2001 1069.8000 ;
	    RECT 1070.1000 1068.9000 1078.2001 1069.5000 ;
	    RECT 1077.0000 1068.6000 1078.2001 1068.9000 ;
	    RECT 1079.7001 1069.5000 1080.6000 1070.7001 ;
	    RECT 1081.5000 1070.4000 1085.4000 1071.6000 ;
	    RECT 1089.0000 1070.4000 1090.2001 1079.7001 ;
	    RECT 1091.4000 1075.5000 1092.6000 1079.7001 ;
	    RECT 1093.8000 1075.5000 1095.0000 1079.7001 ;
	    RECT 1096.2001 1075.5000 1097.4000 1079.7001 ;
	    RECT 1098.6000 1073.7001 1099.8000 1079.7001 ;
	    RECT 1093.8000 1071.6000 1100.1000 1072.8000 ;
	    RECT 1101.0000 1071.6000 1102.2001 1079.7001 ;
	    RECT 1103.4000 1073.7001 1104.6000 1079.7001 ;
	    RECT 1105.8000 1072.8000 1107.0000 1079.7001 ;
	    RECT 1108.2001 1073.7001 1109.4000 1079.7001 ;
	    RECT 1105.8000 1071.9000 1109.7001 1072.8000 ;
	    RECT 1110.6000 1072.5000 1111.8000 1079.7001 ;
	    RECT 1113.0000 1073.7001 1114.2001 1079.7001 ;
	    RECT 1101.0000 1070.4000 1104.9000 1071.6000 ;
	    RECT 1091.4000 1069.5000 1092.6000 1069.8000 ;
	    RECT 1079.7001 1068.6000 1092.6000 1069.5000 ;
	    RECT 1096.2001 1069.5000 1097.4000 1069.8000 ;
	    RECT 1108.8000 1069.5000 1109.7001 1071.9000 ;
	    RECT 1110.6000 1070.4000 1111.8000 1071.6000 ;
	    RECT 1096.2001 1068.6000 1109.7001 1069.5000 ;
	    RECT 1067.4000 1067.4000 1068.6000 1068.6000 ;
	    RECT 1072.5000 1067.7001 1073.7001 1068.0000 ;
	    RECT 1069.5000 1066.8000 1107.9000 1067.7001 ;
	    RECT 1106.7001 1066.5000 1107.9000 1066.8000 ;
	    RECT 1108.8000 1065.9000 1109.7001 1068.6000 ;
	    RECT 1110.6000 1068.0000 1111.8000 1069.5000 ;
	    RECT 1110.6000 1066.8000 1112.1000 1068.0000 ;
	    RECT 1064.7001 1065.0000 1071.3000 1065.9000 ;
	    RECT 1064.7001 1064.7001 1065.9000 1065.0000 ;
	    RECT 1072.2001 1064.4000 1073.4000 1065.6000 ;
	    RECT 1074.3000 1065.0000 1099.8000 1065.9000 ;
	    RECT 1108.8000 1065.0000 1110.0000 1065.9000 ;
	    RECT 1098.6000 1064.1000 1099.8000 1065.0000 ;
	    RECT 911.4000 1063.2001 912.6000 1063.5000 ;
	    RECT 796.2000 1062.4501 797.4000 1062.6000 ;
	    RECT 817.8000 1062.4501 819.0000 1062.6000 ;
	    RECT 796.2000 1061.5500 819.0000 1062.4501 ;
	    RECT 796.2000 1061.4000 797.4000 1061.5500 ;
	    RECT 817.8000 1061.4000 819.0000 1061.5500 ;
	    RECT 849.0000 1061.4000 850.2000 1062.6000 ;
	    RECT 851.1000 1060.8000 851.4000 1062.3000 ;
	    RECT 853.8000 1061.4000 855.0000 1062.6000 ;
	    RECT 855.9000 1061.4000 857.4000 1062.3000 ;
	    RECT 858.6000 1061.4000 859.8000 1062.6000 ;
	    RECT 870.6000 1062.4501 871.8000 1062.6000 ;
	    RECT 877.8000 1062.4501 879.0000 1062.6000 ;
	    RECT 870.6000 1061.5500 879.0000 1062.4501 ;
	    RECT 870.6000 1061.4000 871.8000 1061.5500 ;
	    RECT 877.8000 1061.4000 879.0000 1061.5500 ;
	    RECT 904.2000 1062.4501 905.4000 1062.6000 ;
	    RECT 906.6000 1062.4501 907.8000 1062.6000 ;
	    RECT 904.2000 1061.5500 907.8000 1062.4501 ;
	    RECT 904.2000 1061.4000 905.4000 1061.5500 ;
	    RECT 906.6000 1061.4000 907.8000 1061.5500 ;
	    RECT 908.7000 1061.4000 910.5000 1062.6000 ;
	    RECT 913.8000 1062.4501 915.0000 1062.6000 ;
	    RECT 925.8000 1062.4501 927.0000 1062.6000 ;
	    RECT 805.8000 1059.4501 807.0000 1059.6000 ;
	    RECT 815.4000 1059.4501 816.6000 1059.6000 ;
	    RECT 791.4000 1053.3000 792.6000 1059.3000 ;
	    RECT 793.8000 1058.4000 796.5000 1059.3000 ;
	    RECT 805.8000 1058.5500 816.6000 1059.4501 ;
	    RECT 805.8000 1058.4000 807.0000 1058.5500 ;
	    RECT 815.4000 1058.4000 816.6000 1058.5500 ;
	    RECT 795.3000 1053.3000 796.5000 1058.4000 ;
	    RECT 815.4000 1057.2001 816.6000 1057.5000 ;
	    RECT 818.1000 1056.3000 819.0000 1060.5000 ;
	    RECT 849.3000 1059.3000 854.7000 1059.9000 ;
	    RECT 856.5000 1059.3000 857.4000 1061.4000 ;
	    RECT 912.6000 1060.8000 912.9000 1062.3000 ;
	    RECT 913.8000 1061.5500 927.0000 1062.4501 ;
	    RECT 913.8000 1061.4000 915.0000 1061.5500 ;
	    RECT 925.8000 1061.4000 927.0000 1061.5500 ;
	    RECT 928.2000 1062.4501 929.4000 1062.6000 ;
	    RECT 935.4000 1062.4501 936.6000 1062.6000 ;
	    RECT 928.2000 1061.5500 936.6000 1062.4501 ;
	    RECT 928.2000 1061.4000 929.4000 1061.5500 ;
	    RECT 935.4000 1061.4000 936.6000 1061.5500 ;
	    RECT 1062.6000 1062.3000 1075.8000 1063.5000 ;
	    RECT 1076.7001 1062.9000 1079.7001 1064.1000 ;
	    RECT 1085.4000 1062.9000 1090.2001 1064.1000 ;
	    RECT 849.0000 1059.0000 855.0000 1059.3000 ;
	    RECT 815.4000 1053.3000 816.6000 1056.3000 ;
	    RECT 817.8000 1053.3000 819.0000 1056.3000 ;
	    RECT 820.2000 1053.3000 821.4000 1056.3000 ;
	    RECT 849.0000 1053.3000 850.2000 1059.0000 ;
	    RECT 851.4000 1053.3000 852.6000 1058.1000 ;
	    RECT 853.8000 1054.2001 855.0000 1059.0000 ;
	    RECT 856.2000 1055.1000 857.4000 1059.3000 ;
	    RECT 858.6000 1054.2001 859.8000 1059.3000 ;
	    RECT 853.8000 1053.3000 859.8000 1054.2001 ;
	    RECT 870.6000 1053.3000 871.8000 1060.5000 ;
	    RECT 873.0000 1059.4501 874.2000 1059.6000 ;
	    RECT 901.8000 1059.4501 903.0000 1059.6000 ;
	    RECT 873.0000 1058.5500 903.0000 1059.4501 ;
	    RECT 906.9000 1059.3000 907.8000 1060.5000 ;
	    RECT 909.3000 1059.3000 914.7000 1059.9000 ;
	    RECT 921.0000 1059.4501 922.2000 1059.6000 ;
	    RECT 928.2000 1059.4501 929.4000 1059.6000 ;
	    RECT 873.0000 1058.4000 874.2000 1058.5500 ;
	    RECT 901.8000 1058.4000 903.0000 1058.5500 ;
	    RECT 873.0000 1057.2001 874.2000 1057.5000 ;
	    RECT 873.0000 1053.3000 874.2000 1056.3000 ;
	    RECT 906.6000 1053.3000 907.8000 1059.3000 ;
	    RECT 909.0000 1059.0000 915.0000 1059.3000 ;
	    RECT 909.0000 1053.3000 910.2000 1059.0000 ;
	    RECT 911.4000 1053.3000 912.6000 1058.1000 ;
	    RECT 913.8000 1053.3000 915.0000 1059.0000 ;
	    RECT 921.0000 1058.5500 929.4000 1059.4501 ;
	    RECT 921.0000 1058.4000 922.2000 1058.5500 ;
	    RECT 928.2000 1058.4000 929.4000 1058.5500 ;
	    RECT 935.4000 1056.3000 936.3000 1060.5000 ;
	    RECT 937.8000 1059.4501 939.0000 1059.6000 ;
	    RECT 1050.6000 1059.4501 1051.8000 1059.6000 ;
	    RECT 937.8000 1058.5500 1051.8000 1059.4501 ;
	    RECT 937.8000 1058.4000 939.0000 1058.5500 ;
	    RECT 1050.6000 1058.4000 1051.8000 1058.5500 ;
	    RECT 937.8000 1057.2001 939.0000 1057.5000 ;
	    RECT 933.0000 1053.3000 934.2000 1056.3000 ;
	    RECT 935.4000 1053.3000 936.6000 1056.3000 ;
	    RECT 937.8000 1053.3000 939.0000 1056.3000 ;
	    RECT 1062.6000 1053.3000 1063.8000 1062.3000 ;
	    RECT 1066.2001 1060.2001 1070.7001 1061.4000 ;
	    RECT 1069.5000 1059.3000 1070.7001 1060.2001 ;
	    RECT 1078.5000 1059.3000 1079.7001 1062.9000 ;
	    RECT 1081.8000 1061.4000 1083.0000 1062.6000 ;
	    RECT 1089.6000 1061.7001 1090.8000 1062.0000 ;
	    RECT 1084.2001 1060.8000 1090.8000 1061.7001 ;
	    RECT 1084.2001 1060.5000 1085.4000 1060.8000 ;
	    RECT 1081.8000 1060.2001 1083.0000 1060.5000 ;
	    RECT 1093.8000 1059.6000 1095.0000 1063.8000 ;
	    RECT 1102.5000 1062.9000 1108.2001 1064.1000 ;
	    RECT 1102.5000 1061.1000 1103.7001 1062.9000 ;
	    RECT 1109.1000 1062.0000 1110.0000 1065.0000 ;
	    RECT 1084.2001 1059.3000 1085.4000 1059.6000 ;
	    RECT 1067.4000 1053.3000 1068.6000 1059.3000 ;
	    RECT 1069.5000 1058.1000 1073.4000 1059.3000 ;
	    RECT 1078.5000 1058.4000 1085.4000 1059.3000 ;
	    RECT 1086.6000 1058.4000 1087.8000 1059.6000 ;
	    RECT 1088.7001 1058.4000 1089.0000 1059.6000 ;
	    RECT 1093.5000 1058.4000 1095.0000 1059.6000 ;
	    RECT 1101.0000 1060.2001 1103.7001 1061.1000 ;
	    RECT 1108.2001 1061.1000 1110.0000 1062.0000 ;
	    RECT 1101.0000 1059.3000 1102.2001 1060.2001 ;
	    RECT 1072.2001 1053.3000 1073.4000 1058.1000 ;
	    RECT 1098.6000 1058.1000 1102.2001 1059.3000 ;
	    RECT 1074.6000 1053.3000 1075.8000 1057.5000 ;
	    RECT 1077.0000 1053.3000 1078.2001 1057.5000 ;
	    RECT 1079.4000 1053.3000 1080.6000 1057.5000 ;
	    RECT 1081.8000 1053.3000 1083.0000 1056.3000 ;
	    RECT 1084.2001 1053.3000 1085.4000 1057.5000 ;
	    RECT 1086.6000 1053.3000 1087.8000 1056.3000 ;
	    RECT 1089.0000 1053.3000 1090.2001 1057.5000 ;
	    RECT 1091.4000 1053.3000 1092.6000 1057.5000 ;
	    RECT 1093.8000 1053.3000 1095.0000 1057.5000 ;
	    RECT 1096.2001 1053.3000 1097.4000 1057.5000 ;
	    RECT 1098.6000 1053.3000 1099.8000 1058.1000 ;
	    RECT 1103.4000 1053.3000 1104.6000 1059.3000 ;
	    RECT 1108.2001 1053.3000 1109.4000 1061.1000 ;
	    RECT 1110.9000 1060.2001 1112.1000 1066.8000 ;
	    RECT 1132.2001 1063.5000 1133.4000 1079.7001 ;
	    RECT 1134.6000 1073.7001 1135.8000 1079.7001 ;
	    RECT 1153.8000 1073.7001 1155.0000 1079.7001 ;
	    RECT 1156.2001 1066.5000 1157.4000 1079.7001 ;
	    RECT 1158.6000 1073.7001 1159.8000 1079.7001 ;
	    RECT 1158.6000 1069.5000 1159.8000 1069.8000 ;
	    RECT 1158.6000 1067.4000 1159.8000 1068.6000 ;
	    RECT 1182.6000 1067.7001 1183.8000 1079.7001 ;
	    RECT 1185.0000 1068.3000 1186.2001 1079.7001 ;
	    RECT 1187.4000 1073.7001 1188.6000 1079.7001 ;
	    RECT 1189.8000 1073.7001 1191.0000 1079.7001 ;
	    RECT 1182.6000 1066.5000 1183.5000 1067.7001 ;
	    RECT 1187.4000 1067.4000 1188.3000 1073.7001 ;
	    RECT 1209.0000 1067.7001 1210.2001 1079.7001 ;
	    RECT 1212.9000 1068.9000 1214.1000 1079.7001 ;
	    RECT 1211.4000 1067.7001 1214.1000 1068.9000 ;
	    RECT 1240.2001 1067.7001 1241.4000 1079.7001 ;
	    RECT 1244.1000 1068.6000 1245.3000 1079.7001 ;
	    RECT 1246.5000 1073.7001 1247.7001 1079.7001 ;
	    RECT 1246.2001 1070.4000 1247.4000 1071.6000 ;
	    RECT 1246.5000 1069.5000 1247.4000 1070.4000 ;
	    RECT 1267.5000 1068.9000 1268.7001 1079.7001 ;
	    RECT 1244.1000 1067.7001 1245.6000 1068.6000 ;
	    RECT 1184.7001 1066.5000 1188.3000 1067.4000 ;
	    RECT 1156.2001 1065.4501 1157.4000 1065.6000 ;
	    RECT 1180.2001 1065.4501 1181.4000 1065.6000 ;
	    RECT 1156.2001 1064.5500 1181.4000 1065.4501 ;
	    RECT 1156.2001 1064.4000 1157.4000 1064.5500 ;
	    RECT 1180.2001 1064.4000 1181.4000 1064.5500 ;
	    RECT 1182.6000 1064.4000 1183.8000 1065.6000 ;
	    RECT 1113.0000 1062.4501 1114.2001 1062.6000 ;
	    RECT 1132.2001 1062.4501 1133.4000 1062.6000 ;
	    RECT 1153.8000 1062.4501 1155.0000 1062.6000 ;
	    RECT 1113.0000 1061.5500 1133.4000 1062.4501 ;
	    RECT 1113.0000 1061.4000 1114.2001 1061.5500 ;
	    RECT 1132.2001 1061.4000 1133.4000 1061.5500 ;
	    RECT 1134.7500 1061.5500 1155.0000 1062.4501 ;
	    RECT 1110.6000 1059.0000 1112.1000 1060.2001 ;
	    RECT 1110.6000 1053.3000 1111.8000 1059.0000 ;
	    RECT 1113.0000 1053.3000 1114.2001 1056.3000 ;
	    RECT 1132.2001 1053.3000 1133.4000 1060.5000 ;
	    RECT 1134.7500 1059.6000 1135.6500 1061.5500 ;
	    RECT 1153.8000 1061.4000 1155.0000 1061.5500 ;
	    RECT 1153.8000 1060.2001 1155.0000 1060.5000 ;
	    RECT 1134.6000 1058.4000 1135.8000 1059.6000 ;
	    RECT 1156.2001 1059.3000 1157.4000 1063.5000 ;
	    RECT 1182.6000 1059.3000 1183.5000 1063.5000 ;
	    RECT 1184.7001 1061.4000 1185.6000 1066.5000 ;
	    RECT 1187.4000 1064.4000 1188.6000 1065.6000 ;
	    RECT 1189.8000 1063.5000 1191.0000 1063.8000 ;
	    RECT 1211.7001 1063.5000 1212.6000 1067.7001 ;
	    RECT 1213.8000 1066.5000 1215.0000 1066.8000 ;
	    RECT 1213.8000 1064.4000 1215.0000 1065.6000 ;
	    RECT 1242.6000 1064.4000 1243.8000 1065.6000 ;
	    RECT 1187.4000 1063.2001 1188.3000 1063.5000 ;
	    RECT 1242.6000 1063.2001 1243.8000 1063.5000 ;
	    RECT 1186.8000 1062.3000 1188.3000 1063.2001 ;
	    RECT 1244.7001 1062.6000 1245.6000 1067.7001 ;
	    RECT 1247.4000 1067.4000 1248.6000 1068.6000 ;
	    RECT 1267.5000 1067.7001 1270.2001 1068.9000 ;
	    RECT 1271.4000 1067.7001 1272.6000 1079.7001 ;
	    RECT 1283.4000 1073.7001 1284.6000 1079.7001 ;
	    RECT 1266.6000 1066.5000 1267.8000 1066.8000 ;
	    RECT 1266.6000 1064.4000 1267.8000 1065.6000 ;
	    RECT 1269.0000 1063.5000 1269.9000 1067.7001 ;
	    RECT 1285.8000 1063.5000 1287.0000 1079.7001 ;
	    RECT 1312.2001 1068.6000 1313.4000 1079.7001 ;
	    RECT 1314.6000 1069.5000 1315.8000 1079.7001 ;
	    RECT 1317.0000 1068.6000 1318.2001 1079.7001 ;
	    RECT 1312.2001 1067.7001 1318.2001 1068.6000 ;
	    RECT 1319.4000 1067.7001 1320.6000 1079.7001 ;
	    RECT 1345.8000 1077.4501 1347.0000 1077.6000 ;
	    RECT 1384.2001 1077.4501 1385.4000 1077.6000 ;
	    RECT 1345.8000 1076.5500 1385.4000 1077.4501 ;
	    RECT 1345.8000 1076.4000 1347.0000 1076.5500 ;
	    RECT 1384.2001 1076.4000 1385.4000 1076.5500 ;
	    RECT 1451.4000 1073.7001 1452.6000 1079.7001 ;
	    RECT 1453.8000 1072.5000 1455.0000 1079.7001 ;
	    RECT 1456.2001 1073.7001 1457.4000 1079.7001 ;
	    RECT 1458.6000 1072.8000 1459.8000 1079.7001 ;
	    RECT 1461.0000 1073.7001 1462.2001 1079.7001 ;
	    RECT 1455.9000 1071.9000 1459.8000 1072.8000 ;
	    RECT 1408.2001 1071.4501 1409.4000 1071.6000 ;
	    RECT 1453.8000 1071.4501 1455.0000 1071.6000 ;
	    RECT 1408.2001 1070.5500 1455.0000 1071.4501 ;
	    RECT 1408.2001 1070.4000 1409.4000 1070.5500 ;
	    RECT 1453.8000 1070.4000 1455.0000 1070.5500 ;
	    RECT 1455.9000 1069.5000 1456.8000 1071.9000 ;
	    RECT 1463.4000 1071.6000 1464.6000 1079.7001 ;
	    RECT 1465.8000 1073.7001 1467.0000 1079.7001 ;
	    RECT 1468.2001 1075.5000 1469.4000 1079.7001 ;
	    RECT 1470.6000 1075.5000 1471.8000 1079.7001 ;
	    RECT 1473.0000 1075.5000 1474.2001 1079.7001 ;
	    RECT 1465.5000 1071.6000 1471.8000 1072.8000 ;
	    RECT 1460.7001 1070.4000 1464.6000 1071.6000 ;
	    RECT 1475.4000 1070.4000 1476.6000 1079.7001 ;
	    RECT 1477.8000 1073.7001 1479.0000 1079.7001 ;
	    RECT 1480.2001 1072.5000 1481.4000 1079.7001 ;
	    RECT 1482.6000 1073.7001 1483.8000 1079.7001 ;
	    RECT 1485.0000 1072.5000 1486.2001 1079.7001 ;
	    RECT 1487.4000 1075.5000 1488.6000 1079.7001 ;
	    RECT 1489.8000 1075.5000 1491.0000 1079.7001 ;
	    RECT 1492.2001 1073.7001 1493.4000 1079.7001 ;
	    RECT 1494.6000 1072.8000 1495.8000 1079.7001 ;
	    RECT 1497.0000 1073.7001 1498.2001 1080.6000 ;
	    RECT 1499.4000 1074.6000 1500.6000 1079.7001 ;
	    RECT 1499.4000 1073.7001 1500.9000 1074.6000 ;
	    RECT 1501.8000 1073.7001 1503.0000 1079.7001 ;
	    RECT 1521.0000 1073.7001 1522.2001 1079.7001 ;
	    RECT 1500.0000 1072.8000 1500.9000 1073.7001 ;
	    RECT 1492.8000 1071.6000 1499.1000 1072.8000 ;
	    RECT 1500.0000 1071.9000 1503.0000 1072.8000 ;
	    RECT 1480.2001 1070.4000 1484.1000 1071.6000 ;
	    RECT 1485.0000 1070.7001 1493.7001 1071.6000 ;
	    RECT 1498.2001 1071.0000 1499.1000 1071.6000 ;
	    RECT 1468.2001 1069.5000 1469.4000 1069.8000 ;
	    RECT 1453.8000 1068.0000 1455.0000 1069.5000 ;
	    RECT 1319.4000 1066.5000 1320.3000 1067.7001 ;
	    RECT 1453.5000 1066.8000 1455.0000 1068.0000 ;
	    RECT 1455.9000 1068.6000 1469.4000 1069.5000 ;
	    RECT 1473.0000 1069.5000 1474.2001 1069.8000 ;
	    RECT 1485.0000 1069.5000 1485.9000 1070.7001 ;
	    RECT 1494.6000 1069.8000 1496.7001 1070.7001 ;
	    RECT 1498.2001 1069.8000 1500.6000 1071.0000 ;
	    RECT 1473.0000 1068.6000 1485.9000 1069.5000 ;
	    RECT 1487.4000 1069.5000 1496.7001 1069.8000 ;
	    RECT 1487.4000 1068.9000 1495.5000 1069.5000 ;
	    RECT 1487.4000 1068.6000 1488.6000 1068.9000 ;
	    RECT 1312.2001 1064.4000 1313.4000 1065.6000 ;
	    RECT 1314.3000 1064.7001 1314.6000 1066.2001 ;
	    RECT 1317.0000 1064.7001 1318.5000 1065.6000 ;
	    RECT 1319.4000 1065.4501 1320.6000 1065.6000 ;
	    RECT 1350.6000 1065.4501 1351.8000 1065.6000 ;
	    RECT 1189.8000 1062.4501 1191.0000 1062.6000 ;
	    RECT 1192.2001 1062.4501 1193.4000 1062.6000 ;
	    RECT 1186.8000 1062.0000 1188.0000 1062.3000 ;
	    RECT 1189.8000 1061.5500 1193.4000 1062.4501 ;
	    RECT 1189.8000 1061.4000 1191.0000 1061.5500 ;
	    RECT 1192.2001 1061.4000 1193.4000 1061.5500 ;
	    RECT 1211.4000 1062.4501 1212.6000 1062.6000 ;
	    RECT 1240.2001 1062.4501 1241.4000 1062.6000 ;
	    RECT 1211.4000 1061.5500 1241.4000 1062.4501 ;
	    RECT 1211.4000 1061.4000 1212.6000 1061.5500 ;
	    RECT 1240.2001 1061.4000 1241.4000 1061.5500 ;
	    RECT 1184.4000 1061.1000 1185.6000 1061.4000 ;
	    RECT 1184.4000 1060.5000 1188.9000 1061.1000 ;
	    RECT 1242.3000 1060.8000 1242.6000 1062.3000 ;
	    RECT 1244.7001 1061.4000 1246.5000 1062.6000 ;
	    RECT 1247.4000 1061.4000 1248.6000 1062.6000 ;
	    RECT 1249.8000 1062.4501 1251.0000 1062.6000 ;
	    RECT 1269.0000 1062.4501 1270.2001 1062.6000 ;
	    RECT 1249.8000 1061.5500 1270.2001 1062.4501 ;
	    RECT 1249.8000 1061.4000 1251.0000 1061.5500 ;
	    RECT 1269.0000 1061.4000 1270.2001 1061.5500 ;
	    RECT 1285.8000 1062.4501 1287.0000 1062.6000 ;
	    RECT 1312.3500 1062.4501 1313.2500 1064.4000 ;
	    RECT 1314.6000 1063.5000 1315.8000 1063.8000 ;
	    RECT 1285.8000 1061.5500 1313.2500 1062.4501 ;
	    RECT 1285.8000 1061.4000 1287.0000 1061.5500 ;
	    RECT 1314.6000 1061.4000 1315.8000 1062.6000 ;
	    RECT 1184.4000 1060.2001 1190.7001 1060.5000 ;
	    RECT 1188.0000 1059.6000 1190.7001 1060.2001 ;
	    RECT 1189.8000 1059.3000 1190.7001 1059.6000 ;
	    RECT 1134.6000 1057.2001 1135.8000 1057.5000 ;
	    RECT 1134.6000 1053.3000 1135.8000 1056.3000 ;
	    RECT 1153.8000 1053.3000 1155.0000 1059.3000 ;
	    RECT 1156.2001 1058.4000 1158.9000 1059.3000 ;
	    RECT 1157.7001 1053.3000 1158.9000 1058.4000 ;
	    RECT 1182.6000 1057.8000 1184.7001 1059.3000 ;
	    RECT 1183.5000 1053.3000 1184.7001 1057.8000 ;
	    RECT 1185.9000 1053.3000 1187.1000 1059.0000 ;
	    RECT 1189.8000 1053.3000 1191.0000 1059.3000 ;
	    RECT 1209.0000 1058.4000 1210.2001 1059.6000 ;
	    RECT 1209.0000 1057.2001 1210.2001 1057.5000 ;
	    RECT 1211.7001 1056.3000 1212.6000 1060.5000 ;
	    RECT 1240.5000 1059.3000 1245.9000 1059.9000 ;
	    RECT 1247.4000 1059.3000 1248.3000 1060.5000 ;
	    RECT 1240.2001 1059.0000 1246.2001 1059.3000 ;
	    RECT 1209.0000 1053.3000 1210.2001 1056.3000 ;
	    RECT 1211.4000 1053.3000 1212.6000 1056.3000 ;
	    RECT 1213.8000 1053.3000 1215.0000 1056.3000 ;
	    RECT 1240.2001 1053.3000 1241.4000 1059.0000 ;
	    RECT 1242.6000 1053.3000 1243.8000 1058.1000 ;
	    RECT 1245.0000 1053.3000 1246.2001 1059.0000 ;
	    RECT 1247.4000 1053.3000 1248.6000 1059.3000 ;
	    RECT 1269.0000 1056.3000 1269.9000 1060.5000 ;
	    RECT 1271.4000 1059.4501 1272.6000 1059.6000 ;
	    RECT 1283.4000 1059.4501 1284.6000 1059.6000 ;
	    RECT 1271.4000 1058.5500 1284.6000 1059.4501 ;
	    RECT 1271.4000 1058.4000 1272.6000 1058.5500 ;
	    RECT 1283.4000 1058.4000 1284.6000 1058.5500 ;
	    RECT 1271.4000 1057.2001 1272.6000 1057.5000 ;
	    RECT 1283.4000 1057.2001 1284.6000 1057.5000 ;
	    RECT 1266.6000 1053.3000 1267.8000 1056.3000 ;
	    RECT 1269.0000 1053.3000 1270.2001 1056.3000 ;
	    RECT 1271.4000 1053.3000 1272.6000 1056.3000 ;
	    RECT 1283.4000 1053.3000 1284.6000 1056.3000 ;
	    RECT 1285.8000 1053.3000 1287.0000 1060.5000 ;
	    RECT 1317.0000 1059.3000 1317.9000 1064.7001 ;
	    RECT 1319.4000 1064.5500 1351.8000 1065.4501 ;
	    RECT 1319.4000 1064.4000 1320.6000 1064.5500 ;
	    RECT 1350.6000 1064.4000 1351.8000 1064.5500 ;
	    RECT 1453.5000 1060.2001 1454.7001 1066.8000 ;
	    RECT 1455.9000 1065.9000 1456.8000 1068.6000 ;
	    RECT 1491.9000 1067.7001 1493.1000 1068.0000 ;
	    RECT 1457.7001 1066.8000 1496.1000 1067.7001 ;
	    RECT 1497.0000 1067.4000 1498.2001 1068.6000 ;
	    RECT 1457.7001 1066.5000 1458.9000 1066.8000 ;
	    RECT 1455.6000 1065.0000 1456.8000 1065.9000 ;
	    RECT 1465.8000 1065.0000 1491.3000 1065.9000 ;
	    RECT 1455.6000 1062.0000 1456.5000 1065.0000 ;
	    RECT 1465.8000 1064.1000 1467.0000 1065.0000 ;
	    RECT 1492.2001 1064.4000 1493.4000 1065.6000 ;
	    RECT 1494.3000 1065.0000 1500.9000 1065.9000 ;
	    RECT 1499.7001 1064.7001 1500.9000 1065.0000 ;
	    RECT 1457.4000 1062.9000 1463.1000 1064.1000 ;
	    RECT 1455.6000 1061.1000 1457.4000 1062.0000 ;
	    RECT 1313.1000 1053.3000 1314.3000 1059.3000 ;
	    RECT 1317.0000 1053.3000 1318.2001 1059.3000 ;
	    RECT 1319.4000 1058.4000 1320.6000 1059.6000 ;
	    RECT 1453.5000 1059.0000 1455.0000 1060.2001 ;
	    RECT 1319.1000 1057.2001 1320.3000 1057.5000 ;
	    RECT 1319.4000 1053.3000 1320.6000 1056.3000 ;
	    RECT 1451.4000 1053.3000 1452.6000 1056.3000 ;
	    RECT 1453.8000 1053.3000 1455.0000 1059.0000 ;
	    RECT 1456.2001 1053.3000 1457.4000 1061.1000 ;
	    RECT 1461.9000 1061.1000 1463.1000 1062.9000 ;
	    RECT 1461.9000 1060.2001 1464.6000 1061.1000 ;
	    RECT 1463.4000 1059.3000 1464.6000 1060.2001 ;
	    RECT 1470.6000 1059.6000 1471.8000 1063.8000 ;
	    RECT 1475.4000 1062.9000 1480.2001 1064.1000 ;
	    RECT 1485.9000 1062.9000 1488.9000 1064.1000 ;
	    RECT 1501.8000 1063.5000 1503.0000 1071.9000 ;
	    RECT 1521.0000 1069.5000 1522.2001 1069.8000 ;
	    RECT 1521.0000 1067.4000 1522.2001 1068.6000 ;
	    RECT 1523.4000 1066.5000 1524.6000 1079.7001 ;
	    RECT 1525.8000 1073.7001 1527.0000 1079.7001 ;
	    RECT 1553.1000 1073.7001 1554.3000 1079.7001 ;
	    RECT 1553.4000 1070.4000 1554.6000 1071.6000 ;
	    RECT 1553.4000 1069.5000 1554.3000 1070.4000 ;
	    RECT 1555.5000 1068.6000 1556.7001 1079.7001 ;
	    RECT 1540.2001 1068.4501 1541.4000 1068.6000 ;
	    RECT 1552.2001 1068.4501 1553.4000 1068.6000 ;
	    RECT 1540.2001 1067.5500 1553.4000 1068.4501 ;
	    RECT 1540.2001 1067.4000 1541.4000 1067.5500 ;
	    RECT 1552.2001 1067.4000 1553.4000 1067.5500 ;
	    RECT 1555.2001 1067.7001 1556.7001 1068.6000 ;
	    RECT 1559.4000 1067.7001 1560.6000 1079.7001 ;
	    RECT 1521.0000 1065.4501 1522.2001 1065.6000 ;
	    RECT 1523.4000 1065.4501 1524.6000 1065.6000 ;
	    RECT 1521.0000 1064.5500 1524.6000 1065.4501 ;
	    RECT 1521.0000 1064.4000 1522.2001 1064.5500 ;
	    RECT 1523.4000 1064.4000 1524.6000 1064.5500 ;
	    RECT 1474.8000 1061.7001 1476.0000 1062.0000 ;
	    RECT 1474.8000 1060.8000 1481.4000 1061.7001 ;
	    RECT 1482.6000 1061.4000 1483.8000 1062.6000 ;
	    RECT 1480.2001 1060.5000 1481.4000 1060.8000 ;
	    RECT 1482.6000 1060.2001 1483.8000 1060.5000 ;
	    RECT 1461.0000 1053.3000 1462.2001 1059.3000 ;
	    RECT 1463.4000 1058.1000 1467.0000 1059.3000 ;
	    RECT 1470.6000 1058.4000 1472.1000 1059.6000 ;
	    RECT 1476.6000 1058.4000 1476.9000 1059.6000 ;
	    RECT 1477.8000 1058.4000 1479.0000 1059.6000 ;
	    RECT 1480.2001 1059.3000 1481.4000 1059.6000 ;
	    RECT 1485.9000 1059.3000 1487.1000 1062.9000 ;
	    RECT 1489.8000 1062.3000 1503.0000 1063.5000 ;
	    RECT 1494.9000 1060.2001 1499.4000 1061.4000 ;
	    RECT 1494.9000 1059.3000 1496.1000 1060.2001 ;
	    RECT 1480.2001 1058.4000 1487.1000 1059.3000 ;
	    RECT 1465.8000 1053.3000 1467.0000 1058.1000 ;
	    RECT 1492.2001 1058.1000 1496.1000 1059.3000 ;
	    RECT 1468.2001 1053.3000 1469.4000 1057.5000 ;
	    RECT 1470.6000 1053.3000 1471.8000 1057.5000 ;
	    RECT 1473.0000 1053.3000 1474.2001 1057.5000 ;
	    RECT 1475.4000 1053.3000 1476.6000 1057.5000 ;
	    RECT 1477.8000 1053.3000 1479.0000 1056.3000 ;
	    RECT 1480.2001 1053.3000 1481.4000 1057.5000 ;
	    RECT 1482.6000 1053.3000 1483.8000 1056.3000 ;
	    RECT 1485.0000 1053.3000 1486.2001 1057.5000 ;
	    RECT 1487.4000 1053.3000 1488.6000 1057.5000 ;
	    RECT 1489.8000 1053.3000 1491.0000 1057.5000 ;
	    RECT 1492.2001 1053.3000 1493.4000 1058.1000 ;
	    RECT 1497.0000 1053.3000 1498.2001 1059.3000 ;
	    RECT 1501.8000 1053.3000 1503.0000 1062.3000 ;
	    RECT 1523.4000 1059.3000 1524.6000 1063.5000 ;
	    RECT 1555.2001 1062.6000 1556.1000 1067.7001 ;
	    RECT 1557.0000 1064.4000 1558.2001 1065.6000 ;
	    RECT 1557.0000 1063.2001 1558.2001 1063.5000 ;
	    RECT 1525.8000 1062.4501 1527.0000 1062.6000 ;
	    RECT 1542.6000 1062.4501 1543.8000 1062.6000 ;
	    RECT 1525.8000 1061.5500 1543.8000 1062.4501 ;
	    RECT 1525.8000 1061.4000 1527.0000 1061.5500 ;
	    RECT 1542.6000 1061.4000 1543.8000 1061.5500 ;
	    RECT 1552.2001 1061.4000 1553.4000 1062.6000 ;
	    RECT 1554.3000 1061.4000 1556.1000 1062.6000 ;
	    RECT 1558.2001 1060.8000 1558.5000 1062.3000 ;
	    RECT 1559.4000 1061.4000 1560.6000 1062.6000 ;
	    RECT 1525.8000 1060.2001 1527.0000 1060.5000 ;
	    RECT 1552.5000 1059.3000 1553.4000 1060.5000 ;
	    RECT 1554.9000 1059.3000 1560.3000 1059.9000 ;
	    RECT 1521.9000 1058.4000 1524.6000 1059.3000 ;
	    RECT 1521.9000 1053.3000 1523.1000 1058.4000 ;
	    RECT 1525.8000 1053.3000 1527.0000 1059.3000 ;
	    RECT 1552.2001 1053.3000 1553.4000 1059.3000 ;
	    RECT 1554.6000 1059.0000 1560.6000 1059.3000 ;
	    RECT 1554.6000 1053.3000 1555.8000 1059.0000 ;
	    RECT 1557.0000 1053.3000 1558.2001 1058.1000 ;
	    RECT 1559.4000 1053.3000 1560.6000 1059.0000 ;
	    RECT 1.2000 1050.6000 1569.0000 1052.4000 ;
	    RECT 18.6000 1043.7001 19.8000 1049.7001 ;
	    RECT 22.5000 1044.6000 23.7000 1049.7001 ;
	    RECT 21.0000 1043.7001 23.7000 1044.6000 ;
	    RECT 49.8000 1043.7001 51.0000 1049.7001 ;
	    RECT 52.2000 1044.0000 53.4000 1049.7001 ;
	    RECT 54.6000 1044.9000 55.8000 1049.7001 ;
	    RECT 57.0000 1044.0000 58.2000 1049.7001 ;
	    RECT 52.2000 1043.7001 58.2000 1044.0000 ;
	    RECT 18.6000 1042.5000 19.8000 1042.8000 ;
	    RECT 18.6000 1040.4000 19.8000 1041.6000 ;
	    RECT 21.0000 1039.5000 22.2000 1043.7001 ;
	    RECT 50.1000 1042.5000 51.0000 1043.7001 ;
	    RECT 52.5000 1043.1000 57.9000 1043.7001 ;
	    RECT 69.0000 1042.5000 70.2000 1049.7001 ;
	    RECT 71.4000 1046.7001 72.6000 1049.7001 ;
	    RECT 85.8000 1046.7001 87.0000 1049.7001 ;
	    RECT 71.4000 1045.5000 72.6000 1045.8000 ;
	    RECT 85.8000 1045.5000 87.0000 1045.8000 ;
	    RECT 71.4000 1044.4501 72.6000 1044.6000 ;
	    RECT 83.4000 1044.4501 84.6000 1044.6000 ;
	    RECT 71.4000 1043.5500 84.6000 1044.4501 ;
	    RECT 71.4000 1043.4000 72.6000 1043.5500 ;
	    RECT 83.4000 1043.4000 84.6000 1043.5500 ;
	    RECT 85.8000 1043.4000 87.0000 1044.6000 ;
	    RECT 88.2000 1042.5000 89.4000 1049.7001 ;
	    RECT 100.2000 1046.7001 101.4000 1049.7001 ;
	    RECT 100.2000 1045.5000 101.4000 1045.8000 ;
	    RECT 100.2000 1043.4000 101.4000 1044.6000 ;
	    RECT 102.6000 1042.5000 103.8000 1049.7001 ;
	    RECT 133.8000 1048.8000 139.8000 1049.7001 ;
	    RECT 133.8000 1043.7001 135.0000 1048.8000 ;
	    RECT 136.2000 1043.7001 137.4000 1047.9000 ;
	    RECT 138.6000 1044.0000 139.8000 1048.8000 ;
	    RECT 141.0000 1044.9000 142.2000 1049.7001 ;
	    RECT 143.4000 1044.0000 144.6000 1049.7001 ;
	    RECT 138.6000 1043.7001 144.6000 1044.0000 ;
	    RECT 49.8000 1040.4000 51.0000 1041.6000 ;
	    RECT 51.9000 1040.4000 53.7000 1041.6000 ;
	    RECT 55.8000 1040.7001 56.1000 1042.2001 ;
	    RECT 136.2000 1041.6000 137.1000 1043.7001 ;
	    RECT 138.9000 1043.1000 144.3000 1043.7001 ;
	    RECT 157.8000 1042.5000 159.0000 1049.7001 ;
	    RECT 160.2000 1046.7001 161.4000 1049.7001 ;
	    RECT 160.2000 1045.5000 161.4000 1045.8000 ;
	    RECT 160.2000 1044.4501 161.4000 1044.6000 ;
	    RECT 172.2000 1044.4501 173.4000 1044.6000 ;
	    RECT 160.2000 1043.5500 173.4000 1044.4501 ;
	    RECT 184.2000 1043.7001 185.4000 1049.7001 ;
	    RECT 186.6000 1044.0000 187.8000 1049.7001 ;
	    RECT 189.0000 1044.9000 190.2000 1049.7001 ;
	    RECT 191.4000 1044.0000 192.6000 1049.7001 ;
	    RECT 186.6000 1043.7001 192.6000 1044.0000 ;
	    RECT 217.8000 1043.7001 219.0000 1049.7001 ;
	    RECT 221.7000 1044.6000 222.9000 1049.7001 ;
	    RECT 241.8000 1046.7001 243.0000 1049.7001 ;
	    RECT 244.2000 1046.7001 245.4000 1049.7001 ;
	    RECT 246.6000 1046.7001 247.8000 1049.7001 ;
	    RECT 265.8000 1046.7001 267.0000 1049.7001 ;
	    RECT 268.2000 1046.7001 269.4000 1049.7001 ;
	    RECT 270.6000 1046.7001 271.8000 1049.7001 ;
	    RECT 220.2000 1043.7001 222.9000 1044.6000 ;
	    RECT 160.2000 1043.4000 161.4000 1043.5500 ;
	    RECT 172.2000 1043.4000 173.4000 1043.5500 ;
	    RECT 184.5000 1042.5000 185.4000 1043.7001 ;
	    RECT 186.9000 1043.1000 192.3000 1043.7001 ;
	    RECT 217.8000 1042.5000 219.0000 1042.8000 ;
	    RECT 57.0000 1040.4000 58.2000 1041.6000 ;
	    RECT 69.0000 1041.4501 70.2000 1041.6000 ;
	    RECT 59.5500 1040.5500 70.2000 1041.4501 ;
	    RECT 21.0000 1038.4501 22.2000 1038.6000 ;
	    RECT 21.0000 1037.5500 50.8500 1038.4501 ;
	    RECT 21.0000 1037.4000 22.2000 1037.5500 ;
	    RECT 18.6000 1023.3000 19.8000 1029.3000 ;
	    RECT 21.0000 1023.3000 22.2000 1036.5000 ;
	    RECT 49.9500 1035.6000 50.8500 1037.5500 ;
	    RECT 23.4000 1034.4000 24.6000 1035.6000 ;
	    RECT 49.8000 1034.4000 51.0000 1035.6000 ;
	    RECT 52.8000 1035.3000 53.7000 1040.4000 ;
	    RECT 54.6000 1039.5000 55.8000 1039.8000 ;
	    RECT 54.6000 1038.4501 55.8000 1038.6000 ;
	    RECT 59.5500 1038.4501 60.4500 1040.5500 ;
	    RECT 69.0000 1040.4000 70.2000 1040.5500 ;
	    RECT 88.2000 1041.4501 89.4000 1041.6000 ;
	    RECT 100.2000 1041.4501 101.4000 1041.6000 ;
	    RECT 88.2000 1040.5500 101.4000 1041.4501 ;
	    RECT 88.2000 1040.4000 89.4000 1040.5500 ;
	    RECT 100.2000 1040.4000 101.4000 1040.5500 ;
	    RECT 102.6000 1041.4501 103.8000 1041.6000 ;
	    RECT 133.8000 1041.4501 135.0000 1041.6000 ;
	    RECT 102.6000 1040.5500 135.0000 1041.4501 ;
	    RECT 136.2000 1040.7001 137.7000 1041.6000 ;
	    RECT 102.6000 1040.4000 103.8000 1040.5500 ;
	    RECT 133.8000 1040.4000 135.0000 1040.5500 ;
	    RECT 138.6000 1040.4000 139.8000 1041.6000 ;
	    RECT 142.2000 1040.7001 142.5000 1042.2001 ;
	    RECT 143.4000 1041.4501 144.6000 1041.6000 ;
	    RECT 145.8000 1041.4501 147.0000 1041.6000 ;
	    RECT 143.4000 1040.5500 147.0000 1041.4501 ;
	    RECT 143.4000 1040.4000 144.6000 1040.5500 ;
	    RECT 145.8000 1040.4000 147.0000 1040.5500 ;
	    RECT 157.8000 1041.4501 159.0000 1041.6000 ;
	    RECT 181.8000 1041.4501 183.0000 1041.6000 ;
	    RECT 157.8000 1040.5500 183.0000 1041.4501 ;
	    RECT 157.8000 1040.4000 159.0000 1040.5500 ;
	    RECT 181.8000 1040.4000 183.0000 1040.5500 ;
	    RECT 184.2000 1040.4000 185.4000 1041.6000 ;
	    RECT 186.3000 1040.4000 188.1000 1041.6000 ;
	    RECT 190.2000 1040.7001 190.5000 1042.2001 ;
	    RECT 191.4000 1041.4501 192.6000 1041.6000 ;
	    RECT 217.8000 1041.4501 219.0000 1041.6000 ;
	    RECT 191.4000 1040.5500 219.0000 1041.4501 ;
	    RECT 191.4000 1040.4000 192.6000 1040.5500 ;
	    RECT 217.8000 1040.4000 219.0000 1040.5500 ;
	    RECT 136.2000 1039.5000 137.4000 1039.8000 ;
	    RECT 141.0000 1039.5000 142.2000 1039.8000 ;
	    RECT 54.6000 1037.5500 60.4500 1038.4501 ;
	    RECT 54.6000 1037.4000 55.8000 1037.5500 ;
	    RECT 52.8000 1034.4000 54.3000 1035.3000 ;
	    RECT 23.4000 1033.2001 24.6000 1033.5000 ;
	    RECT 51.0000 1032.6000 51.9000 1033.5000 ;
	    RECT 51.0000 1031.4000 52.2000 1032.6000 ;
	    RECT 23.4000 1023.3000 24.6000 1029.3000 ;
	    RECT 50.7000 1023.3000 51.9000 1029.3000 ;
	    RECT 53.1000 1023.3000 54.3000 1034.4000 ;
	    RECT 57.0000 1023.3000 58.2000 1035.3000 ;
	    RECT 69.0000 1023.3000 70.2000 1039.5000 ;
	    RECT 71.4000 1023.3000 72.6000 1029.3000 ;
	    RECT 85.8000 1023.3000 87.0000 1029.3000 ;
	    RECT 88.2000 1023.3000 89.4000 1039.5000 ;
	    RECT 100.2000 1023.3000 101.4000 1029.3000 ;
	    RECT 102.6000 1023.3000 103.8000 1039.5000 ;
	    RECT 133.8000 1039.2001 135.0000 1039.5000 ;
	    RECT 136.2000 1037.4000 137.4000 1038.6000 ;
	    RECT 138.9000 1035.3000 139.8000 1039.5000 ;
	    RECT 141.0000 1038.4501 142.2000 1038.6000 ;
	    RECT 143.4000 1038.4501 144.6000 1038.6000 ;
	    RECT 141.0000 1037.5500 144.6000 1038.4501 ;
	    RECT 141.0000 1037.4000 142.2000 1037.5500 ;
	    RECT 143.4000 1037.4000 144.6000 1037.5500 ;
	    RECT 133.8000 1023.3000 135.0000 1035.3000 ;
	    RECT 137.7000 1023.3000 140.7000 1035.3000 ;
	    RECT 143.4000 1023.3000 144.6000 1035.3000 ;
	    RECT 157.8000 1023.3000 159.0000 1039.5000 ;
	    RECT 184.2000 1034.4000 185.4000 1035.6000 ;
	    RECT 187.2000 1035.3000 188.1000 1040.4000 ;
	    RECT 189.0000 1039.5000 190.2000 1039.8000 ;
	    RECT 220.2000 1039.5000 221.4000 1043.7001 ;
	    RECT 244.2000 1042.5000 245.1000 1046.7001 ;
	    RECT 246.6000 1045.5000 247.8000 1045.8000 ;
	    RECT 246.6000 1043.4000 247.8000 1044.6000 ;
	    RECT 268.2000 1042.5000 269.1000 1046.7001 ;
	    RECT 270.6000 1045.5000 271.8000 1045.8000 ;
	    RECT 290.7000 1044.6000 291.9000 1049.7001 ;
	    RECT 270.6000 1044.4501 271.8000 1044.6000 ;
	    RECT 273.0000 1044.4501 274.2000 1044.6000 ;
	    RECT 270.6000 1043.5500 274.2000 1044.4501 ;
	    RECT 290.7000 1043.7001 293.4000 1044.6000 ;
	    RECT 294.6000 1043.7001 295.8000 1049.7001 ;
	    RECT 309.0000 1046.7001 310.2000 1049.7001 ;
	    RECT 309.0000 1045.5000 310.2000 1045.8000 ;
	    RECT 270.6000 1043.4000 271.8000 1043.5500 ;
	    RECT 273.0000 1043.4000 274.2000 1043.5500 ;
	    RECT 244.2000 1041.4501 245.4000 1041.6000 ;
	    RECT 263.4000 1041.4501 264.6000 1041.6000 ;
	    RECT 244.2000 1040.5500 264.6000 1041.4501 ;
	    RECT 244.2000 1040.4000 245.4000 1040.5500 ;
	    RECT 263.4000 1040.4000 264.6000 1040.5500 ;
	    RECT 268.2000 1040.4000 269.4000 1041.6000 ;
	    RECT 292.2000 1039.5000 293.4000 1043.7001 ;
	    RECT 309.0000 1043.4000 310.2000 1044.6000 ;
	    RECT 294.6000 1042.5000 295.8000 1042.8000 ;
	    RECT 311.4000 1042.5000 312.6000 1049.7001 ;
	    RECT 313.8000 1044.4501 315.0000 1044.6000 ;
	    RECT 340.2000 1044.4501 341.4000 1044.6000 ;
	    RECT 313.8000 1043.5500 341.4000 1044.4501 ;
	    RECT 342.6000 1044.0000 343.8000 1049.7001 ;
	    RECT 345.0000 1044.9000 346.2000 1049.7001 ;
	    RECT 347.4000 1048.8000 353.4000 1049.7001 ;
	    RECT 347.4000 1044.0000 348.6000 1048.8000 ;
	    RECT 342.6000 1043.7001 348.6000 1044.0000 ;
	    RECT 349.8000 1043.7001 351.0000 1047.9000 ;
	    RECT 352.2000 1043.7001 353.4000 1048.8000 ;
	    RECT 484.2000 1046.7001 485.4000 1049.7001 ;
	    RECT 486.6000 1044.0000 487.8000 1049.7001 ;
	    RECT 313.8000 1043.4000 315.0000 1043.5500 ;
	    RECT 340.2000 1043.4000 341.4000 1043.5500 ;
	    RECT 342.9000 1043.1000 348.3000 1043.7001 ;
	    RECT 294.6000 1040.4000 295.8000 1041.6000 ;
	    RECT 311.4000 1041.4501 312.6000 1041.6000 ;
	    RECT 342.6000 1041.4501 343.8000 1041.6000 ;
	    RECT 311.4000 1040.5500 343.8000 1041.4501 ;
	    RECT 344.7000 1040.7001 345.0000 1042.2001 ;
	    RECT 350.1000 1041.6000 351.0000 1043.7001 ;
	    RECT 486.3000 1042.8000 487.8000 1044.0000 ;
	    RECT 311.4000 1040.4000 312.6000 1040.5500 ;
	    RECT 342.6000 1040.4000 343.8000 1040.5500 ;
	    RECT 347.4000 1040.4000 348.6000 1041.6000 ;
	    RECT 349.5000 1040.7001 351.0000 1041.6000 ;
	    RECT 352.2000 1041.4501 353.4000 1041.6000 ;
	    RECT 357.0000 1041.4501 358.2000 1041.6000 ;
	    RECT 352.2000 1040.5500 358.2000 1041.4501 ;
	    RECT 352.2000 1040.4000 353.4000 1040.5500 ;
	    RECT 357.0000 1040.4000 358.2000 1040.5500 ;
	    RECT 345.0000 1039.5000 346.2000 1039.8000 ;
	    RECT 349.8000 1039.5000 351.0000 1039.8000 ;
	    RECT 189.0000 1037.4000 190.2000 1038.6000 ;
	    RECT 191.4000 1038.4501 192.6000 1038.6000 ;
	    RECT 220.2000 1038.4501 221.4000 1038.6000 ;
	    RECT 191.4000 1037.5500 221.4000 1038.4501 ;
	    RECT 191.4000 1037.4000 192.6000 1037.5500 ;
	    RECT 220.2000 1037.4000 221.4000 1037.5500 ;
	    RECT 229.8000 1038.4501 231.0000 1038.6000 ;
	    RECT 241.8000 1038.4501 243.0000 1038.6000 ;
	    RECT 229.8000 1037.5500 243.0000 1038.4501 ;
	    RECT 229.8000 1037.4000 231.0000 1037.5500 ;
	    RECT 241.8000 1037.4000 243.0000 1037.5500 ;
	    RECT 187.2000 1034.4000 188.7000 1035.3000 ;
	    RECT 185.4000 1032.6000 186.3000 1033.5000 ;
	    RECT 185.4000 1031.4000 186.6000 1032.6000 ;
	    RECT 160.2000 1023.3000 161.4000 1029.3000 ;
	    RECT 185.1000 1023.3000 186.3000 1029.3000 ;
	    RECT 187.5000 1023.3000 188.7000 1034.4000 ;
	    RECT 191.4000 1023.3000 192.6000 1035.3000 ;
	    RECT 217.8000 1023.3000 219.0000 1029.3000 ;
	    RECT 220.2000 1023.3000 221.4000 1036.5000 ;
	    RECT 241.8000 1036.2001 243.0000 1036.5000 ;
	    RECT 222.6000 1034.4000 223.8000 1035.6000 ;
	    RECT 244.2000 1035.3000 245.1000 1039.5000 ;
	    RECT 265.8000 1037.4000 267.0000 1038.6000 ;
	    RECT 265.8000 1036.2001 267.0000 1036.5000 ;
	    RECT 268.2000 1035.3000 269.1000 1039.5000 ;
	    RECT 292.2000 1037.4000 293.4000 1038.6000 ;
	    RECT 273.0000 1035.4501 274.2000 1035.6000 ;
	    RECT 289.8000 1035.4501 291.0000 1035.6000 ;
	    RECT 242.7000 1034.1000 245.4000 1035.3000 ;
	    RECT 222.6000 1033.2001 223.8000 1033.5000 ;
	    RECT 222.6000 1023.3000 223.8000 1029.3000 ;
	    RECT 242.7000 1023.3000 243.9000 1034.1000 ;
	    RECT 246.6000 1023.3000 247.8000 1035.3000 ;
	    RECT 266.7000 1034.1000 269.4000 1035.3000 ;
	    RECT 266.7000 1023.3000 267.9000 1034.1000 ;
	    RECT 270.6000 1023.3000 271.8000 1035.3000 ;
	    RECT 273.0000 1034.5500 291.0000 1035.4501 ;
	    RECT 273.0000 1034.4000 274.2000 1034.5500 ;
	    RECT 289.8000 1034.4000 291.0000 1034.5500 ;
	    RECT 289.8000 1033.2001 291.0000 1033.5000 ;
	    RECT 289.8000 1023.3000 291.0000 1029.3000 ;
	    RECT 292.2000 1023.3000 293.4000 1036.5000 ;
	    RECT 294.6000 1023.3000 295.8000 1029.3000 ;
	    RECT 309.0000 1023.3000 310.2000 1029.3000 ;
	    RECT 311.4000 1023.3000 312.6000 1039.5000 ;
	    RECT 337.8000 1038.4501 339.0000 1038.6000 ;
	    RECT 345.0000 1038.4501 346.2000 1038.6000 ;
	    RECT 337.8000 1037.5500 346.2000 1038.4501 ;
	    RECT 337.8000 1037.4000 339.0000 1037.5500 ;
	    RECT 345.0000 1037.4000 346.2000 1037.5500 ;
	    RECT 347.4000 1035.3000 348.3000 1039.5000 ;
	    RECT 352.2000 1039.2001 353.4000 1039.5000 ;
	    RECT 349.8000 1037.4000 351.0000 1038.6000 ;
	    RECT 486.3000 1036.2001 487.5000 1042.8000 ;
	    RECT 489.0000 1041.9000 490.2000 1049.7001 ;
	    RECT 493.8000 1043.7001 495.0000 1049.7001 ;
	    RECT 498.6000 1044.9000 499.8000 1049.7001 ;
	    RECT 501.0000 1045.5000 502.2000 1049.7001 ;
	    RECT 503.4000 1045.5000 504.6000 1049.7001 ;
	    RECT 505.8000 1045.5000 507.0000 1049.7001 ;
	    RECT 508.2000 1045.5000 509.4000 1049.7001 ;
	    RECT 510.6000 1046.7001 511.8000 1049.7001 ;
	    RECT 513.0000 1045.5000 514.2000 1049.7001 ;
	    RECT 515.4000 1046.7001 516.6000 1049.7001 ;
	    RECT 517.8000 1045.5000 519.0000 1049.7001 ;
	    RECT 520.2000 1045.5000 521.4000 1049.7001 ;
	    RECT 522.6000 1045.5000 523.8000 1049.7001 ;
	    RECT 496.2000 1043.7001 499.8000 1044.9000 ;
	    RECT 525.0000 1044.9000 526.2000 1049.7001 ;
	    RECT 496.2000 1042.8000 497.4000 1043.7001 ;
	    RECT 488.4000 1041.0000 490.2000 1041.9000 ;
	    RECT 494.7000 1041.9000 497.4000 1042.8000 ;
	    RECT 503.4000 1043.4000 504.9000 1044.6000 ;
	    RECT 509.4000 1043.4000 509.7000 1044.6000 ;
	    RECT 510.6000 1043.4000 511.8000 1044.6000 ;
	    RECT 513.0000 1043.7001 519.9000 1044.6000 ;
	    RECT 525.0000 1043.7001 528.9000 1044.9000 ;
	    RECT 529.8000 1043.7001 531.0000 1049.7001 ;
	    RECT 513.0000 1043.4000 514.2000 1043.7001 ;
	    RECT 488.4000 1038.0000 489.3000 1041.0000 ;
	    RECT 494.7000 1040.1000 495.9000 1041.9000 ;
	    RECT 490.2000 1038.9000 495.9000 1040.1000 ;
	    RECT 503.4000 1039.2001 504.6000 1043.4000 ;
	    RECT 515.4000 1042.5000 516.6000 1042.8000 ;
	    RECT 513.0000 1042.2001 514.2000 1042.5000 ;
	    RECT 507.6000 1041.3000 514.2000 1042.2001 ;
	    RECT 507.6000 1041.0000 508.8000 1041.3000 ;
	    RECT 515.4000 1040.4000 516.6000 1041.6000 ;
	    RECT 518.7000 1040.1000 519.9000 1043.7001 ;
	    RECT 527.7000 1042.8000 528.9000 1043.7001 ;
	    RECT 527.7000 1041.6000 532.2000 1042.8000 ;
	    RECT 534.6000 1040.7001 535.8000 1049.7001 ;
	    RECT 587.4000 1043.7001 588.6000 1049.7001 ;
	    RECT 589.8000 1042.8000 591.0000 1049.7001 ;
	    RECT 592.2000 1043.7001 593.4000 1049.7001 ;
	    RECT 594.6000 1042.8000 595.8000 1049.7001 ;
	    RECT 597.0000 1043.7001 598.2000 1049.7001 ;
	    RECT 599.4000 1042.8000 600.6000 1049.7001 ;
	    RECT 601.8000 1043.7001 603.0000 1049.7001 ;
	    RECT 604.2000 1042.8000 605.4000 1049.7001 ;
	    RECT 606.6000 1043.7001 607.8000 1049.7001 ;
	    RECT 633.0000 1046.7001 634.2000 1049.7001 ;
	    RECT 633.3000 1045.5000 634.5000 1045.8000 ;
	    RECT 625.8000 1044.4501 627.0000 1044.6000 ;
	    RECT 633.0000 1044.4501 634.2000 1044.6000 ;
	    RECT 625.8000 1043.5500 634.2000 1044.4501 ;
	    RECT 635.4000 1043.7001 636.6000 1049.7001 ;
	    RECT 639.3000 1043.7001 640.5000 1049.7001 ;
	    RECT 672.3000 1043.7001 673.5000 1049.7001 ;
	    RECT 676.2000 1043.7001 677.4000 1049.7001 ;
	    RECT 678.6000 1046.7001 679.8000 1049.7001 ;
	    RECT 678.3000 1045.5000 679.5000 1045.8000 ;
	    RECT 625.8000 1043.4000 627.0000 1043.5500 ;
	    RECT 633.0000 1043.4000 634.2000 1043.5500 ;
	    RECT 508.2000 1038.9000 513.0000 1040.1000 ;
	    RECT 518.7000 1038.9000 521.7000 1040.1000 ;
	    RECT 522.6000 1039.5000 535.8000 1040.7001 ;
	    RECT 587.4000 1041.6000 591.0000 1042.8000 ;
	    RECT 592.5000 1041.6000 595.8000 1042.8000 ;
	    RECT 597.3000 1041.6000 600.6000 1042.8000 ;
	    RECT 602.7000 1041.6000 605.4000 1042.8000 ;
	    RECT 587.4000 1039.5000 588.6000 1041.6000 ;
	    RECT 592.5000 1040.7001 593.7000 1041.6000 ;
	    RECT 597.3000 1040.7001 598.5000 1041.6000 ;
	    RECT 602.7000 1040.7001 603.9000 1041.6000 ;
	    RECT 589.8000 1039.5000 593.7000 1040.7001 ;
	    RECT 594.9000 1039.5000 598.5000 1040.7001 ;
	    RECT 600.0000 1039.5000 603.9000 1040.7001 ;
	    RECT 605.1000 1039.5000 605.7000 1040.7001 ;
	    RECT 498.6000 1038.0000 499.8000 1038.9000 ;
	    RECT 488.4000 1037.1000 489.6000 1038.0000 ;
	    RECT 498.6000 1037.1000 524.1000 1038.0000 ;
	    RECT 525.0000 1037.4000 526.2000 1038.6000 ;
	    RECT 532.5000 1038.0000 533.7000 1038.3000 ;
	    RECT 527.1000 1037.1000 533.7000 1038.0000 ;
	    RECT 342.6000 1023.3000 343.8000 1035.3000 ;
	    RECT 346.5000 1023.3000 349.5000 1035.3000 ;
	    RECT 352.2000 1023.3000 353.4000 1035.3000 ;
	    RECT 486.3000 1035.0000 487.8000 1036.2001 ;
	    RECT 486.6000 1033.5000 487.8000 1035.0000 ;
	    RECT 488.7000 1034.4000 489.6000 1037.1000 ;
	    RECT 490.5000 1036.2001 491.7000 1036.5000 ;
	    RECT 490.5000 1035.3000 528.9000 1036.2001 ;
	    RECT 524.7000 1035.0000 525.9000 1035.3000 ;
	    RECT 529.8000 1034.4000 531.0000 1035.6000 ;
	    RECT 488.7000 1033.5000 502.2000 1034.4000 ;
	    RECT 409.8000 1032.4501 411.0000 1032.6000 ;
	    RECT 486.6000 1032.4501 487.8000 1032.6000 ;
	    RECT 409.8000 1031.5500 487.8000 1032.4501 ;
	    RECT 409.8000 1031.4000 411.0000 1031.5500 ;
	    RECT 486.6000 1031.4000 487.8000 1031.5500 ;
	    RECT 488.7000 1031.1000 489.6000 1033.5000 ;
	    RECT 501.0000 1033.2001 502.2000 1033.5000 ;
	    RECT 505.8000 1033.5000 518.7000 1034.4000 ;
	    RECT 505.8000 1033.2001 507.0000 1033.5000 ;
	    RECT 493.5000 1031.4000 497.4000 1032.6000 ;
	    RECT 484.2000 1023.3000 485.4000 1029.3000 ;
	    RECT 486.6000 1023.3000 487.8000 1030.5000 ;
	    RECT 488.7000 1030.2001 492.6000 1031.1000 ;
	    RECT 489.0000 1023.3000 490.2000 1029.3000 ;
	    RECT 491.4000 1023.3000 492.6000 1030.2001 ;
	    RECT 493.8000 1023.3000 495.0000 1029.3000 ;
	    RECT 496.2000 1023.3000 497.4000 1031.4000 ;
	    RECT 498.3000 1030.2001 504.6000 1031.4000 ;
	    RECT 498.6000 1023.3000 499.8000 1029.3000 ;
	    RECT 501.0000 1023.3000 502.2000 1027.5000 ;
	    RECT 503.4000 1023.3000 504.6000 1027.5000 ;
	    RECT 505.8000 1023.3000 507.0000 1027.5000 ;
	    RECT 508.2000 1023.3000 509.4000 1032.6000 ;
	    RECT 513.0000 1031.4000 516.9000 1032.6000 ;
	    RECT 517.8000 1032.3000 518.7000 1033.5000 ;
	    RECT 520.2000 1034.1000 521.4000 1034.4000 ;
	    RECT 520.2000 1033.5000 528.3000 1034.1000 ;
	    RECT 520.2000 1033.2001 529.5000 1033.5000 ;
	    RECT 527.4000 1032.3000 529.5000 1033.2001 ;
	    RECT 517.8000 1031.4000 526.5000 1032.3000 ;
	    RECT 531.0000 1032.0000 533.4000 1033.2001 ;
	    RECT 531.0000 1031.4000 531.9000 1032.0000 ;
	    RECT 510.6000 1023.3000 511.8000 1029.3000 ;
	    RECT 513.0000 1023.3000 514.2000 1030.5000 ;
	    RECT 515.4000 1023.3000 516.6000 1029.3000 ;
	    RECT 517.8000 1023.3000 519.0000 1030.5000 ;
	    RECT 525.6000 1030.2001 531.9000 1031.4000 ;
	    RECT 534.6000 1031.1000 535.8000 1039.5000 ;
	    RECT 539.4000 1038.4501 540.6000 1038.6000 ;
	    RECT 587.4000 1038.4501 588.6000 1038.6000 ;
	    RECT 539.4000 1037.5500 588.6000 1038.4501 ;
	    RECT 539.4000 1037.4000 540.6000 1037.5500 ;
	    RECT 587.4000 1037.4000 588.6000 1037.5500 ;
	    RECT 592.5000 1037.4000 593.7000 1039.5000 ;
	    RECT 597.3000 1037.4000 598.5000 1039.5000 ;
	    RECT 602.7000 1037.4000 603.9000 1039.5000 ;
	    RECT 633.0000 1037.4000 634.2000 1038.6000 ;
	    RECT 635.7000 1038.3000 636.6000 1043.7001 ;
	    RECT 637.8000 1040.4000 639.0000 1041.6000 ;
	    RECT 673.8000 1040.4000 675.0000 1041.6000 ;
	    RECT 637.8000 1039.2001 639.0000 1039.5000 ;
	    RECT 673.8000 1039.2001 675.0000 1039.5000 ;
	    RECT 635.1000 1037.4000 636.6000 1038.3000 ;
	    RECT 589.5000 1036.5000 591.0000 1037.4000 ;
	    RECT 587.4000 1036.2001 591.0000 1036.5000 ;
	    RECT 592.5000 1036.2001 595.8000 1037.4000 ;
	    RECT 597.3000 1036.2001 600.6000 1037.4000 ;
	    RECT 602.7000 1036.2001 605.4000 1037.4000 ;
	    RECT 639.0000 1036.8000 639.3000 1038.3000 ;
	    RECT 640.2000 1037.4000 641.4000 1038.6000 ;
	    RECT 642.6000 1038.4501 643.8000 1038.6000 ;
	    RECT 657.0000 1038.4501 658.2000 1038.6000 ;
	    RECT 671.4000 1038.4501 672.6000 1038.6000 ;
	    RECT 642.6000 1037.5500 672.6000 1038.4501 ;
	    RECT 676.2000 1038.3000 677.1000 1043.7001 ;
	    RECT 678.6000 1043.4000 679.8000 1044.6000 ;
	    RECT 719.4000 1043.7001 720.6000 1049.7001 ;
	    RECT 721.8000 1044.6000 723.3000 1049.7001 ;
	    RECT 726.0000 1044.3000 728.4000 1049.7001 ;
	    RECT 731.1000 1044.6000 732.6000 1049.7001 ;
	    RECT 719.4000 1042.8000 723.3000 1043.7001 ;
	    RECT 722.1000 1042.5000 723.3000 1042.8000 ;
	    RECT 724.2000 1042.2001 726.6000 1043.4000 ;
	    RECT 700.2000 1041.4501 701.4000 1041.6000 ;
	    RECT 719.4000 1041.4501 720.6000 1041.6000 ;
	    RECT 700.2000 1040.5500 720.6000 1041.4501 ;
	    RECT 700.2000 1040.4000 701.4000 1040.5500 ;
	    RECT 719.4000 1040.4000 720.6000 1040.5500 ;
	    RECT 721.5000 1041.3000 721.8000 1041.6000 ;
	    RECT 727.5000 1041.3000 728.4000 1044.3000 ;
	    RECT 733.8000 1043.7001 735.0000 1049.7001 ;
	    RECT 748.2000 1046.7001 749.4000 1049.7001 ;
	    RECT 748.2000 1045.5000 749.4000 1045.8000 ;
	    RECT 729.3000 1042.2001 730.5000 1043.4000 ;
	    RECT 731.4000 1042.8000 735.0000 1043.7001 ;
	    RECT 745.8000 1044.4501 747.0000 1044.6000 ;
	    RECT 748.2000 1044.4501 749.4000 1044.6000 ;
	    RECT 745.8000 1043.5500 749.4000 1044.4501 ;
	    RECT 745.8000 1043.4000 747.0000 1043.5500 ;
	    RECT 748.2000 1043.4000 749.4000 1043.5500 ;
	    RECT 731.4000 1042.5000 732.6000 1042.8000 ;
	    RECT 750.6000 1042.5000 751.8000 1049.7001 ;
	    RECT 765.0000 1042.5000 766.2000 1049.7001 ;
	    RECT 767.4000 1046.7001 768.6000 1049.7001 ;
	    RECT 781.8000 1046.7001 783.0000 1049.7001 ;
	    RECT 767.4000 1045.5000 768.6000 1045.8000 ;
	    RECT 781.8000 1045.5000 783.0000 1045.8000 ;
	    RECT 767.4000 1043.4000 768.6000 1044.6000 ;
	    RECT 781.8000 1043.4000 783.0000 1044.6000 ;
	    RECT 784.2000 1042.5000 785.4000 1049.7001 ;
	    RECT 813.0000 1044.0000 814.2000 1049.7001 ;
	    RECT 815.4000 1044.9000 816.6000 1049.7001 ;
	    RECT 817.8000 1048.8000 823.8000 1049.7001 ;
	    RECT 817.8000 1044.0000 819.0000 1048.8000 ;
	    RECT 813.0000 1043.7001 819.0000 1044.0000 ;
	    RECT 820.2000 1043.7001 821.4000 1047.9000 ;
	    RECT 822.6000 1043.7001 823.8000 1048.8000 ;
	    RECT 842.7000 1044.6000 843.9000 1049.7001 ;
	    RECT 842.7000 1043.7001 845.4000 1044.6000 ;
	    RECT 846.6000 1043.7001 847.8000 1049.7001 ;
	    RECT 873.0000 1043.7001 874.2000 1049.7001 ;
	    RECT 875.4000 1044.0000 876.6000 1049.7001 ;
	    RECT 877.8000 1044.9000 879.0000 1049.7001 ;
	    RECT 880.2000 1044.0000 881.4000 1049.7001 ;
	    RECT 892.2000 1046.7001 893.4000 1049.7001 ;
	    RECT 892.2000 1045.5000 893.4000 1045.8000 ;
	    RECT 875.4000 1043.7001 881.4000 1044.0000 ;
	    RECT 813.3000 1043.1000 818.7000 1043.7001 ;
	    RECT 721.5000 1041.0000 722.7000 1041.3000 ;
	    RECT 721.5000 1040.4000 726.0000 1041.0000 ;
	    RECT 721.8000 1040.1000 726.0000 1040.4000 ;
	    RECT 724.8000 1039.8000 726.0000 1040.1000 ;
	    RECT 726.9000 1040.4000 728.4000 1041.3000 ;
	    RECT 729.6000 1041.6000 730.5000 1042.2001 ;
	    RECT 729.6000 1040.4000 730.8000 1041.6000 ;
	    RECT 732.6000 1040.4000 732.9000 1041.6000 ;
	    RECT 733.8000 1040.4000 735.0000 1041.6000 ;
	    RECT 750.6000 1041.4501 751.8000 1041.6000 ;
	    RECT 762.6000 1041.4501 763.8000 1041.6000 ;
	    RECT 750.6000 1040.5500 763.8000 1041.4501 ;
	    RECT 750.6000 1040.4000 751.8000 1040.5500 ;
	    RECT 762.6000 1040.4000 763.8000 1040.5500 ;
	    RECT 765.0000 1041.4501 766.2000 1041.6000 ;
	    RECT 779.4000 1041.4501 780.6000 1041.6000 ;
	    RECT 765.0000 1040.5500 780.6000 1041.4501 ;
	    RECT 765.0000 1040.4000 766.2000 1040.5500 ;
	    RECT 779.4000 1040.4000 780.6000 1040.5500 ;
	    RECT 784.2000 1041.4501 785.4000 1041.6000 ;
	    RECT 813.0000 1041.4501 814.2000 1041.6000 ;
	    RECT 784.2000 1040.5500 814.2000 1041.4501 ;
	    RECT 815.1000 1040.7001 815.4000 1042.2001 ;
	    RECT 820.5000 1041.6000 821.4000 1043.7001 ;
	    RECT 784.2000 1040.4000 785.4000 1040.5500 ;
	    RECT 813.0000 1040.4000 814.2000 1040.5500 ;
	    RECT 817.8000 1040.4000 819.0000 1041.6000 ;
	    RECT 819.9000 1040.7001 821.4000 1041.6000 ;
	    RECT 822.6000 1040.4000 823.8000 1041.6000 ;
	    RECT 726.9000 1039.5000 727.8000 1040.4000 ;
	    RECT 815.4000 1039.5000 816.6000 1039.8000 ;
	    RECT 820.2000 1039.5000 821.4000 1039.8000 ;
	    RECT 844.2000 1039.5000 845.4000 1043.7001 ;
	    RECT 846.6000 1042.5000 847.8000 1042.8000 ;
	    RECT 873.3000 1042.5000 874.2000 1043.7001 ;
	    RECT 875.7000 1043.1000 881.1000 1043.7001 ;
	    RECT 892.2000 1043.4000 893.4000 1044.6000 ;
	    RECT 894.6000 1042.5000 895.8000 1049.7001 ;
	    RECT 901.8000 1047.4501 903.0000 1047.6000 ;
	    RECT 916.2000 1047.4501 917.4000 1047.6000 ;
	    RECT 901.8000 1046.5500 917.4000 1047.4501 ;
	    RECT 901.8000 1046.4000 903.0000 1046.5500 ;
	    RECT 916.2000 1046.4000 917.4000 1046.5500 ;
	    RECT 921.0000 1043.7001 922.2000 1049.7001 ;
	    RECT 924.9000 1044.6000 926.1000 1049.7001 ;
	    RECT 923.4000 1043.7001 926.1000 1044.6000 ;
	    RECT 978.6000 1043.7001 979.8000 1049.7001 ;
	    RECT 921.0000 1042.5000 922.2000 1042.8000 ;
	    RECT 846.6000 1041.4501 847.8000 1041.6000 ;
	    RECT 856.2000 1041.4501 857.4000 1041.6000 ;
	    RECT 846.6000 1040.5500 857.4000 1041.4501 ;
	    RECT 846.6000 1040.4000 847.8000 1040.5500 ;
	    RECT 856.2000 1040.4000 857.4000 1040.5500 ;
	    RECT 873.0000 1040.4000 874.2000 1041.6000 ;
	    RECT 875.1000 1040.4000 876.9000 1041.6000 ;
	    RECT 879.0000 1040.7001 879.3000 1042.2001 ;
	    RECT 880.2000 1041.4501 881.4000 1041.6000 ;
	    RECT 889.8000 1041.4501 891.0000 1041.6000 ;
	    RECT 880.2000 1040.5500 891.0000 1041.4501 ;
	    RECT 880.2000 1040.4000 881.4000 1040.5500 ;
	    RECT 889.8000 1040.4000 891.0000 1040.5500 ;
	    RECT 894.6000 1041.4501 895.8000 1041.6000 ;
	    RECT 911.4000 1041.4501 912.6000 1041.6000 ;
	    RECT 894.6000 1040.5500 912.6000 1041.4501 ;
	    RECT 894.6000 1040.4000 895.8000 1040.5500 ;
	    RECT 911.4000 1040.4000 912.6000 1040.5500 ;
	    RECT 921.0000 1040.4000 922.2000 1041.6000 ;
	    RECT 678.6000 1038.4501 679.8000 1038.6000 ;
	    RECT 719.4000 1038.4501 720.6000 1038.6000 ;
	    RECT 642.6000 1037.4000 643.8000 1037.5500 ;
	    RECT 657.0000 1037.4000 658.2000 1037.5500 ;
	    RECT 671.4000 1037.4000 672.6000 1037.5500 ;
	    RECT 673.5000 1036.8000 673.8000 1038.3000 ;
	    RECT 676.2000 1037.4000 677.7000 1038.3000 ;
	    RECT 678.6000 1037.5500 720.6000 1038.4501 ;
	    RECT 678.6000 1037.4000 679.8000 1037.5500 ;
	    RECT 719.4000 1037.4000 720.6000 1037.5500 ;
	    RECT 722.7000 1038.3000 723.9000 1038.6000 ;
	    RECT 726.6000 1038.4501 727.8000 1038.6000 ;
	    RECT 748.2000 1038.4501 749.4000 1038.6000 ;
	    RECT 722.7000 1037.4000 725.1000 1038.3000 ;
	    RECT 726.6000 1037.5500 749.4000 1038.4501 ;
	    RECT 726.6000 1037.4000 727.8000 1037.5500 ;
	    RECT 748.2000 1037.4000 749.4000 1037.5500 ;
	    RECT 723.9000 1037.1000 725.1000 1037.4000 ;
	    RECT 532.8000 1030.2001 535.8000 1031.1000 ;
	    RECT 520.2000 1023.3000 521.4000 1027.5000 ;
	    RECT 522.6000 1023.3000 523.8000 1027.5000 ;
	    RECT 525.0000 1023.3000 526.2000 1029.3000 ;
	    RECT 527.4000 1023.3000 528.6000 1030.2001 ;
	    RECT 532.8000 1029.3000 533.7000 1030.2001 ;
	    RECT 529.8000 1022.4000 531.0000 1029.3000 ;
	    RECT 532.2000 1028.4000 533.7000 1029.3000 ;
	    RECT 532.2000 1023.3000 533.4000 1028.4000 ;
	    RECT 534.6000 1023.3000 535.8000 1029.3000 ;
	    RECT 587.4000 1023.3000 588.6000 1035.3000 ;
	    RECT 589.8000 1023.3000 591.0000 1036.2001 ;
	    RECT 592.2000 1023.3000 593.4000 1035.3000 ;
	    RECT 594.6000 1023.3000 595.8000 1036.2001 ;
	    RECT 597.0000 1023.3000 598.2000 1035.3000 ;
	    RECT 599.4000 1023.3000 600.6000 1036.2001 ;
	    RECT 601.8000 1023.3000 603.0000 1035.3000 ;
	    RECT 604.2000 1023.3000 605.4000 1036.2001 ;
	    RECT 633.3000 1035.3000 634.2000 1036.5000 ;
	    RECT 678.6000 1035.3000 679.5000 1036.5000 ;
	    RECT 726.9000 1035.3000 727.8000 1036.5000 ;
	    RECT 606.6000 1023.3000 607.8000 1035.3000 ;
	    RECT 633.0000 1023.3000 634.2000 1035.3000 ;
	    RECT 635.4000 1034.4000 641.4000 1035.3000 ;
	    RECT 635.4000 1023.3000 636.6000 1034.4000 ;
	    RECT 637.8000 1023.3000 639.0000 1033.5000 ;
	    RECT 640.2000 1023.3000 641.4000 1034.4000 ;
	    RECT 671.4000 1034.4000 677.4000 1035.3000 ;
	    RECT 671.4000 1023.3000 672.6000 1034.4000 ;
	    RECT 673.8000 1023.3000 675.0000 1033.5000 ;
	    RECT 676.2000 1023.3000 677.4000 1034.4000 ;
	    RECT 678.6000 1023.3000 679.8000 1035.3000 ;
	    RECT 719.4000 1034.4000 723.3000 1035.3000 ;
	    RECT 719.4000 1023.3000 720.6000 1034.4000 ;
	    RECT 722.1000 1034.1000 723.3000 1034.4000 ;
	    RECT 721.8000 1023.3000 723.3000 1033.2001 ;
	    RECT 726.0000 1023.3000 728.4000 1035.3000 ;
	    RECT 731.4000 1034.4000 735.0000 1035.3000 ;
	    RECT 731.4000 1034.1000 732.6000 1034.4000 ;
	    RECT 731.1000 1023.3000 732.6000 1033.2001 ;
	    RECT 733.8000 1023.3000 735.0000 1034.4000 ;
	    RECT 748.2000 1023.3000 749.4000 1029.3000 ;
	    RECT 750.6000 1023.3000 751.8000 1039.5000 ;
	    RECT 765.0000 1023.3000 766.2000 1039.5000 ;
	    RECT 767.4000 1023.3000 768.6000 1029.3000 ;
	    RECT 781.8000 1023.3000 783.0000 1029.3000 ;
	    RECT 784.2000 1023.3000 785.4000 1039.5000 ;
	    RECT 808.2000 1038.4501 809.4000 1038.6000 ;
	    RECT 813.0000 1038.4501 814.2000 1038.6000 ;
	    RECT 808.2000 1037.5500 814.2000 1038.4501 ;
	    RECT 808.2000 1037.4000 809.4000 1037.5500 ;
	    RECT 813.0000 1037.4000 814.2000 1037.5500 ;
	    RECT 815.4000 1037.4000 816.6000 1038.6000 ;
	    RECT 817.8000 1035.3000 818.7000 1039.5000 ;
	    RECT 822.6000 1039.2001 823.8000 1039.5000 ;
	    RECT 820.2000 1037.4000 821.4000 1038.6000 ;
	    RECT 844.2000 1038.4501 845.4000 1038.6000 ;
	    RECT 844.2000 1037.5500 874.0500 1038.4501 ;
	    RECT 844.2000 1037.4000 845.4000 1037.5500 ;
	    RECT 839.4000 1035.4501 840.6000 1035.6000 ;
	    RECT 841.8000 1035.4501 843.0000 1035.6000 ;
	    RECT 813.0000 1023.3000 814.2000 1035.3000 ;
	    RECT 816.9000 1023.3000 819.9000 1035.3000 ;
	    RECT 822.6000 1023.3000 823.8000 1035.3000 ;
	    RECT 839.4000 1034.5500 843.0000 1035.4501 ;
	    RECT 839.4000 1034.4000 840.6000 1034.5500 ;
	    RECT 841.8000 1034.4000 843.0000 1034.5500 ;
	    RECT 841.8000 1033.2001 843.0000 1033.5000 ;
	    RECT 841.8000 1023.3000 843.0000 1029.3000 ;
	    RECT 844.2000 1023.3000 845.4000 1036.5000 ;
	    RECT 873.1500 1035.6000 874.0500 1037.5500 ;
	    RECT 873.0000 1034.4000 874.2000 1035.6000 ;
	    RECT 876.0000 1035.3000 876.9000 1040.4000 ;
	    RECT 877.8000 1039.5000 879.0000 1039.8000 ;
	    RECT 923.4000 1039.5000 924.6000 1043.7001 ;
	    RECT 981.0000 1042.8000 982.2000 1049.7001 ;
	    RECT 983.4000 1043.7001 984.6000 1049.7001 ;
	    RECT 985.8000 1042.8000 987.0000 1049.7001 ;
	    RECT 988.2000 1043.7001 989.4000 1049.7001 ;
	    RECT 990.6000 1042.8000 991.8000 1049.7001 ;
	    RECT 993.0000 1043.7001 994.2000 1049.7001 ;
	    RECT 995.4000 1042.8000 996.6000 1049.7001 ;
	    RECT 997.8000 1043.7001 999.0000 1049.7001 ;
	    RECT 1017.9000 1044.6000 1019.1000 1049.7001 ;
	    RECT 1017.9000 1043.7001 1020.6000 1044.6000 ;
	    RECT 1021.8000 1043.7001 1023.0000 1049.7001 ;
	    RECT 1036.2001 1046.7001 1037.4000 1049.7001 ;
	    RECT 1036.2001 1045.5000 1037.4000 1045.8000 ;
	    RECT 981.0000 1041.6000 983.7000 1042.8000 ;
	    RECT 985.8000 1041.6000 989.1000 1042.8000 ;
	    RECT 990.6000 1041.6000 993.9000 1042.8000 ;
	    RECT 995.4000 1041.6000 999.0000 1042.8000 ;
	    RECT 957.0000 1041.4501 958.2000 1041.6000 ;
	    RECT 978.6000 1041.4501 979.8000 1041.6000 ;
	    RECT 957.0000 1040.5500 979.8000 1041.4501 ;
	    RECT 982.5000 1040.7001 983.7000 1041.6000 ;
	    RECT 987.9000 1040.7001 989.1000 1041.6000 ;
	    RECT 992.7000 1040.7001 993.9000 1041.6000 ;
	    RECT 957.0000 1040.4000 958.2000 1040.5500 ;
	    RECT 978.6000 1040.4000 979.8000 1040.5500 ;
	    RECT 980.7000 1039.5000 981.3000 1040.7001 ;
	    RECT 982.5000 1039.5000 986.4000 1040.7001 ;
	    RECT 987.9000 1039.5000 991.5000 1040.7001 ;
	    RECT 992.7000 1039.5000 996.6000 1040.7001 ;
	    RECT 997.8000 1039.5000 999.0000 1041.6000 ;
	    RECT 1019.4000 1039.5000 1020.6000 1043.7001 ;
	    RECT 1036.2001 1043.4000 1037.4000 1044.6000 ;
	    RECT 1021.8000 1042.5000 1023.0000 1042.8000 ;
	    RECT 1038.6000 1042.5000 1039.8000 1049.7001 ;
	    RECT 1091.4000 1043.7001 1092.6000 1049.7001 ;
	    RECT 1093.8000 1042.8000 1095.0000 1049.7001 ;
	    RECT 1096.2001 1043.7001 1097.4000 1049.7001 ;
	    RECT 1098.6000 1042.8000 1099.8000 1049.7001 ;
	    RECT 1101.0000 1043.7001 1102.2001 1049.7001 ;
	    RECT 1103.4000 1042.8000 1104.6000 1049.7001 ;
	    RECT 1105.8000 1043.7001 1107.0000 1049.7001 ;
	    RECT 1108.2001 1042.8000 1109.4000 1049.7001 ;
	    RECT 1110.6000 1043.7001 1111.8000 1049.7001 ;
	    RECT 1093.8000 1041.6000 1096.5000 1042.8000 ;
	    RECT 1098.6000 1041.6000 1101.9000 1042.8000 ;
	    RECT 1103.4000 1041.6000 1106.7001 1042.8000 ;
	    RECT 1108.2001 1041.6000 1111.8000 1042.8000 ;
	    RECT 1187.4000 1042.5000 1188.6000 1049.7001 ;
	    RECT 1189.8000 1043.7001 1191.0000 1049.7001 ;
	    RECT 1194.0000 1047.6000 1195.2001 1049.7001 ;
	    RECT 1192.2001 1046.7001 1195.2001 1047.6000 ;
	    RECT 1197.9000 1046.7001 1199.4000 1049.7001 ;
	    RECT 1200.6000 1046.7001 1201.8000 1049.7001 ;
	    RECT 1203.0000 1046.7001 1204.2001 1049.7001 ;
	    RECT 1206.9000 1047.6000 1208.7001 1049.7001 ;
	    RECT 1206.6000 1046.7001 1208.7001 1047.6000 ;
	    RECT 1192.2001 1045.5000 1193.4000 1046.7001 ;
	    RECT 1200.6000 1045.8000 1201.5000 1046.7001 ;
	    RECT 1194.6000 1044.6000 1195.8000 1045.8000 ;
	    RECT 1197.3000 1044.9000 1201.5000 1045.8000 ;
	    RECT 1206.6000 1045.5000 1207.8000 1046.7001 ;
	    RECT 1197.3000 1044.6000 1198.5000 1044.9000 ;
	    RECT 1021.8000 1040.4000 1023.0000 1041.6000 ;
	    RECT 1026.6000 1041.4501 1027.8000 1041.6000 ;
	    RECT 1038.6000 1041.4501 1039.8000 1041.6000 ;
	    RECT 1026.6000 1040.5500 1039.8000 1041.4501 ;
	    RECT 1095.3000 1040.7001 1096.5000 1041.6000 ;
	    RECT 1100.7001 1040.7001 1101.9000 1041.6000 ;
	    RECT 1105.5000 1040.7001 1106.7001 1041.6000 ;
	    RECT 1026.6000 1040.4000 1027.8000 1040.5500 ;
	    RECT 1038.6000 1040.4000 1039.8000 1040.5500 ;
	    RECT 1093.5000 1039.5000 1094.1000 1040.7001 ;
	    RECT 1095.3000 1039.5000 1099.2001 1040.7001 ;
	    RECT 1100.7001 1039.5000 1104.3000 1040.7001 ;
	    RECT 1105.5000 1039.5000 1109.4000 1040.7001 ;
	    RECT 1110.6000 1039.5000 1111.8000 1041.6000 ;
	    RECT 1188.6000 1040.4000 1188.9000 1041.6000 ;
	    RECT 1189.8000 1040.4000 1191.0000 1041.6000 ;
	    RECT 1194.9000 1041.3000 1195.8000 1044.6000 ;
	    RECT 1211.4000 1044.0000 1212.6000 1049.7001 ;
	    RECT 1209.3000 1043.1000 1210.5000 1043.4000 ;
	    RECT 1213.8000 1043.1000 1215.0000 1049.7001 ;
	    RECT 1237.8000 1043.7001 1239.0000 1049.7001 ;
	    RECT 1240.2001 1044.0000 1241.4000 1049.7001 ;
	    RECT 1242.6000 1044.9000 1243.8000 1049.7001 ;
	    RECT 1245.0000 1044.0000 1246.2001 1049.7001 ;
	    RECT 1259.4000 1046.7001 1260.6000 1049.7001 ;
	    RECT 1259.4000 1045.5000 1260.6000 1045.8000 ;
	    RECT 1240.2001 1043.7001 1246.2001 1044.0000 ;
	    RECT 1209.3000 1042.2001 1215.0000 1043.1000 ;
	    RECT 1238.1000 1042.5000 1239.0000 1043.7001 ;
	    RECT 1240.5000 1043.1000 1245.9000 1043.7001 ;
	    RECT 1259.4000 1043.4000 1260.6000 1044.6000 ;
	    RECT 1261.8000 1042.5000 1263.0000 1049.7001 ;
	    RECT 1285.8000 1044.0000 1287.0000 1049.7001 ;
	    RECT 1288.2001 1044.9000 1289.4000 1049.7001 ;
	    RECT 1290.6000 1044.0000 1291.8000 1049.7001 ;
	    RECT 1285.8000 1043.7001 1291.8000 1044.0000 ;
	    RECT 1293.0000 1043.7001 1294.2001 1049.7001 ;
	    RECT 1307.4000 1046.7001 1308.6000 1049.7001 ;
	    RECT 1307.4000 1045.5000 1308.6000 1045.8000 ;
	    RECT 1286.1000 1043.1000 1291.5000 1043.7001 ;
	    RECT 1293.0000 1042.5000 1293.9000 1043.7001 ;
	    RECT 1307.4000 1043.4000 1308.6000 1044.6000 ;
	    RECT 1309.8000 1042.5000 1311.0000 1049.7001 ;
	    RECT 1357.8000 1043.7001 1359.0000 1049.7001 ;
	    RECT 1360.2001 1044.6000 1361.7001 1049.7001 ;
	    RECT 1364.4000 1044.3000 1366.8000 1049.7001 ;
	    RECT 1369.5000 1044.6000 1371.0000 1049.7001 ;
	    RECT 1357.8000 1042.8000 1361.7001 1043.7001 ;
	    RECT 1360.5000 1042.5000 1361.7001 1042.8000 ;
	    RECT 1362.6000 1042.2001 1365.0000 1043.4000 ;
	    RECT 1203.3000 1041.3000 1204.5000 1041.6000 ;
	    RECT 1191.9000 1040.4000 1205.1000 1041.3000 ;
	    RECT 1193.1000 1040.1000 1194.3000 1040.4000 ;
	    RECT 877.8000 1037.4000 879.0000 1038.6000 ;
	    RECT 876.0000 1034.4000 877.5000 1035.3000 ;
	    RECT 874.2000 1032.6000 875.1000 1033.5000 ;
	    RECT 874.2000 1031.4000 875.4000 1032.6000 ;
	    RECT 846.6000 1023.3000 847.8000 1029.3000 ;
	    RECT 873.9000 1023.3000 875.1000 1029.3000 ;
	    RECT 876.3000 1023.3000 877.5000 1034.4000 ;
	    RECT 880.2000 1023.3000 881.4000 1035.3000 ;
	    RECT 892.2000 1023.3000 893.4000 1029.3000 ;
	    RECT 894.6000 1023.3000 895.8000 1039.5000 ;
	    RECT 906.6000 1038.4501 907.8000 1038.6000 ;
	    RECT 923.4000 1038.4501 924.6000 1038.6000 ;
	    RECT 906.6000 1037.5500 924.6000 1038.4501 ;
	    RECT 906.6000 1037.4000 907.8000 1037.5500 ;
	    RECT 923.4000 1037.4000 924.6000 1037.5500 ;
	    RECT 982.5000 1037.4000 983.7000 1039.5000 ;
	    RECT 987.9000 1037.4000 989.1000 1039.5000 ;
	    RECT 992.7000 1037.4000 993.9000 1039.5000 ;
	    RECT 997.8000 1037.4000 999.0000 1038.6000 ;
	    RECT 1019.4000 1038.4501 1020.6000 1038.6000 ;
	    RECT 1036.2001 1038.4501 1037.4000 1038.6000 ;
	    RECT 1019.4000 1037.5500 1037.4000 1038.4501 ;
	    RECT 1019.4000 1037.4000 1020.6000 1037.5500 ;
	    RECT 1036.2001 1037.4000 1037.4000 1037.5500 ;
	    RECT 916.2000 1032.4501 917.4000 1032.6000 ;
	    RECT 921.0000 1032.4501 922.2000 1032.6000 ;
	    RECT 916.2000 1031.5500 922.2000 1032.4501 ;
	    RECT 916.2000 1031.4000 917.4000 1031.5500 ;
	    RECT 921.0000 1031.4000 922.2000 1031.5500 ;
	    RECT 921.0000 1023.3000 922.2000 1029.3000 ;
	    RECT 923.4000 1023.3000 924.6000 1036.5000 ;
	    RECT 981.0000 1036.2001 983.7000 1037.4000 ;
	    RECT 985.8000 1036.2001 989.1000 1037.4000 ;
	    RECT 990.6000 1036.2001 993.9000 1037.4000 ;
	    RECT 995.4000 1036.5000 996.9000 1037.4000 ;
	    RECT 995.4000 1036.2001 999.0000 1036.5000 ;
	    RECT 925.8000 1035.4501 927.0000 1035.6000 ;
	    RECT 973.8000 1035.4501 975.0000 1035.6000 ;
	    RECT 925.8000 1034.5500 975.0000 1035.4501 ;
	    RECT 925.8000 1034.4000 927.0000 1034.5500 ;
	    RECT 973.8000 1034.4000 975.0000 1034.5500 ;
	    RECT 925.8000 1033.2001 927.0000 1033.5000 ;
	    RECT 925.8000 1023.3000 927.0000 1029.3000 ;
	    RECT 978.6000 1023.3000 979.8000 1035.3000 ;
	    RECT 981.0000 1023.3000 982.2000 1036.2001 ;
	    RECT 983.4000 1023.3000 984.6000 1035.3000 ;
	    RECT 985.8000 1023.3000 987.0000 1036.2001 ;
	    RECT 988.2000 1023.3000 989.4000 1035.3000 ;
	    RECT 990.6000 1023.3000 991.8000 1036.2001 ;
	    RECT 993.0000 1023.3000 994.2000 1035.3000 ;
	    RECT 995.4000 1023.3000 996.6000 1036.2001 ;
	    RECT 997.8000 1023.3000 999.0000 1035.3000 ;
	    RECT 1017.0000 1034.4000 1018.2000 1035.6000 ;
	    RECT 1017.0000 1033.2001 1018.2000 1033.5000 ;
	    RECT 1017.0000 1023.3000 1018.2000 1029.3000 ;
	    RECT 1019.4000 1023.3000 1020.6000 1036.5000 ;
	    RECT 1021.8000 1023.3000 1023.0000 1029.3000 ;
	    RECT 1036.2001 1023.3000 1037.4000 1029.3000 ;
	    RECT 1038.6000 1023.3000 1039.8000 1039.5000 ;
	    RECT 1095.3000 1037.4000 1096.5000 1039.5000 ;
	    RECT 1100.7001 1037.4000 1101.9000 1039.5000 ;
	    RECT 1105.5000 1037.4000 1106.7001 1039.5000 ;
	    RECT 1190.7001 1038.6000 1191.9000 1038.9000 ;
	    RECT 1110.6000 1037.4000 1111.8000 1038.6000 ;
	    RECT 1190.7001 1037.7001 1196.1000 1038.6000 ;
	    RECT 1197.0000 1037.4000 1198.2001 1038.6000 ;
	    RECT 1093.8000 1036.2001 1096.5000 1037.4000 ;
	    RECT 1098.6000 1036.2001 1101.9000 1037.4000 ;
	    RECT 1103.4000 1036.2001 1106.7001 1037.4000 ;
	    RECT 1108.2001 1036.5000 1109.7001 1037.4000 ;
	    RECT 1187.4000 1036.5000 1195.8000 1036.8000 ;
	    RECT 1108.2001 1036.2001 1111.8000 1036.5000 ;
	    RECT 1187.4000 1036.2001 1196.1000 1036.5000 ;
	    RECT 1091.4000 1023.3000 1092.6000 1035.3000 ;
	    RECT 1093.8000 1023.3000 1095.0000 1036.2001 ;
	    RECT 1096.2001 1023.3000 1097.4000 1035.3000 ;
	    RECT 1098.6000 1023.3000 1099.8000 1036.2001 ;
	    RECT 1101.0000 1023.3000 1102.2001 1035.3000 ;
	    RECT 1103.4000 1023.3000 1104.6000 1036.2001 ;
	    RECT 1105.8000 1023.3000 1107.0000 1035.3000 ;
	    RECT 1108.2001 1023.3000 1109.4000 1036.2001 ;
	    RECT 1187.4000 1035.9000 1202.1000 1036.2001 ;
	    RECT 1110.6000 1023.3000 1111.8000 1035.3000 ;
	    RECT 1187.4000 1023.3000 1188.6000 1035.9000 ;
	    RECT 1194.9000 1035.3000 1202.1000 1035.9000 ;
	    RECT 1189.8000 1023.3000 1191.0000 1035.0000 ;
	    RECT 1192.2001 1033.5000 1200.3000 1034.4000 ;
	    RECT 1192.2001 1033.2001 1193.4000 1033.5000 ;
	    RECT 1199.1000 1033.2001 1200.3000 1033.5000 ;
	    RECT 1201.2001 1033.5000 1202.1000 1035.3000 ;
	    RECT 1204.2001 1035.6000 1205.1000 1040.4000 ;
	    RECT 1213.8000 1039.5000 1215.0000 1042.2001 ;
	    RECT 1216.2001 1041.4501 1217.4000 1041.6000 ;
	    RECT 1237.8000 1041.4501 1239.0000 1041.6000 ;
	    RECT 1216.2001 1040.5500 1239.0000 1041.4501 ;
	    RECT 1216.2001 1040.4000 1217.4000 1040.5500 ;
	    RECT 1237.8000 1040.4000 1239.0000 1040.5500 ;
	    RECT 1239.9000 1040.4000 1241.7001 1041.6000 ;
	    RECT 1243.8000 1040.7001 1244.1000 1042.2001 ;
	    RECT 1245.0000 1040.4000 1246.2001 1041.6000 ;
	    RECT 1261.8000 1041.4501 1263.0000 1041.6000 ;
	    RECT 1266.6000 1041.4501 1267.8000 1041.6000 ;
	    RECT 1261.8000 1040.5500 1267.8000 1041.4501 ;
	    RECT 1261.8000 1040.4000 1263.0000 1040.5500 ;
	    RECT 1266.6000 1040.4000 1267.8000 1040.5500 ;
	    RECT 1285.8000 1040.4000 1287.0000 1041.6000 ;
	    RECT 1287.9000 1040.7001 1288.2001 1042.2001 ;
	    RECT 1290.3000 1040.4000 1292.1000 1041.6000 ;
	    RECT 1293.0000 1041.4501 1294.2001 1041.6000 ;
	    RECT 1295.4000 1041.4501 1296.6000 1041.6000 ;
	    RECT 1293.0000 1040.5500 1296.6000 1041.4501 ;
	    RECT 1293.0000 1040.4000 1294.2001 1040.5500 ;
	    RECT 1295.4000 1040.4000 1296.6000 1040.5500 ;
	    RECT 1297.8000 1041.4501 1299.0000 1041.6000 ;
	    RECT 1309.8000 1041.4501 1311.0000 1041.6000 ;
	    RECT 1297.8000 1040.5500 1311.0000 1041.4501 ;
	    RECT 1297.8000 1040.4000 1299.0000 1040.5500 ;
	    RECT 1309.8000 1040.4000 1311.0000 1040.5500 ;
	    RECT 1357.8000 1040.4000 1359.0000 1041.6000 ;
	    RECT 1359.9000 1041.3000 1360.2001 1041.6000 ;
	    RECT 1365.9000 1041.3000 1366.8000 1044.3000 ;
	    RECT 1372.2001 1043.7001 1373.4000 1049.7001 ;
	    RECT 1377.0000 1047.4501 1378.2001 1047.6000 ;
	    RECT 1475.4000 1047.4501 1476.6000 1047.6000 ;
	    RECT 1492.2001 1047.4501 1493.4000 1047.6000 ;
	    RECT 1377.0000 1046.5500 1493.4000 1047.4501 ;
	    RECT 1497.0000 1046.7001 1498.2001 1049.7001 ;
	    RECT 1377.0000 1046.4000 1378.2001 1046.5500 ;
	    RECT 1475.4000 1046.4000 1476.6000 1046.5500 ;
	    RECT 1492.2001 1046.4000 1493.4000 1046.5500 ;
	    RECT 1367.7001 1042.2001 1368.9000 1043.4000 ;
	    RECT 1369.8000 1042.8000 1373.4000 1043.7001 ;
	    RECT 1379.4000 1044.4501 1380.6000 1044.6000 ;
	    RECT 1389.0000 1044.4501 1390.2001 1044.6000 ;
	    RECT 1379.4000 1043.5500 1390.2001 1044.4501 ;
	    RECT 1499.4000 1044.0000 1500.6000 1049.7001 ;
	    RECT 1379.4000 1043.4000 1380.6000 1043.5500 ;
	    RECT 1389.0000 1043.4000 1390.2001 1043.5500 ;
	    RECT 1499.1000 1042.8000 1500.6000 1044.0000 ;
	    RECT 1369.8000 1042.5000 1371.0000 1042.8000 ;
	    RECT 1359.9000 1041.0000 1361.1000 1041.3000 ;
	    RECT 1359.9000 1040.4000 1364.4000 1041.0000 ;
	    RECT 1206.6000 1039.2001 1207.8000 1039.5000 ;
	    RECT 1206.6000 1038.3000 1212.3000 1039.2001 ;
	    RECT 1211.1000 1038.0000 1212.3000 1038.3000 ;
	    RECT 1213.8000 1038.4501 1215.0000 1038.6000 ;
	    RECT 1223.4000 1038.4501 1224.6000 1038.6000 ;
	    RECT 1213.8000 1037.5500 1224.6000 1038.4501 ;
	    RECT 1213.8000 1037.4000 1215.0000 1037.5500 ;
	    RECT 1223.4000 1037.4000 1224.6000 1037.5500 ;
	    RECT 1208.7001 1037.1000 1209.9000 1037.4000 ;
	    RECT 1208.7001 1036.5000 1212.9000 1037.1000 ;
	    RECT 1208.7001 1036.2001 1215.0000 1036.5000 ;
	    RECT 1204.2001 1034.7001 1207.8000 1035.6000 ;
	    RECT 1203.3000 1033.5000 1204.5000 1033.8000 ;
	    RECT 1201.2001 1032.6000 1204.5000 1033.5000 ;
	    RECT 1206.9000 1033.2001 1207.8000 1034.7001 ;
	    RECT 1206.9000 1032.0000 1209.0000 1033.2001 ;
	    RECT 1197.3000 1031.1000 1198.5000 1031.4000 ;
	    RECT 1201.5000 1031.1000 1202.7001 1031.4000 ;
	    RECT 1192.2001 1029.3000 1193.4000 1030.5000 ;
	    RECT 1197.3000 1030.2001 1202.7001 1031.1000 ;
	    RECT 1200.6000 1029.3000 1201.5000 1030.2001 ;
	    RECT 1206.6000 1029.3000 1207.8000 1030.5000 ;
	    RECT 1192.2001 1028.4000 1195.2001 1029.3000 ;
	    RECT 1194.0000 1023.3000 1195.2001 1028.4000 ;
	    RECT 1198.2001 1023.3000 1199.4000 1029.3000 ;
	    RECT 1200.6000 1023.3000 1201.8000 1029.3000 ;
	    RECT 1203.0000 1023.3000 1204.2001 1029.3000 ;
	    RECT 1206.9000 1023.3000 1208.7001 1029.3000 ;
	    RECT 1211.4000 1023.3000 1212.6000 1035.3000 ;
	    RECT 1213.8000 1023.3000 1215.0000 1036.2001 ;
	    RECT 1237.8000 1034.4000 1239.0000 1035.6000 ;
	    RECT 1240.8000 1035.3000 1241.7001 1040.4000 ;
	    RECT 1242.6000 1039.5000 1243.8000 1039.8000 ;
	    RECT 1288.2001 1039.5000 1289.4000 1039.8000 ;
	    RECT 1242.6000 1038.4501 1243.8000 1038.6000 ;
	    RECT 1245.0000 1038.4501 1246.2001 1038.6000 ;
	    RECT 1242.6000 1037.5500 1246.2001 1038.4501 ;
	    RECT 1242.6000 1037.4000 1243.8000 1037.5500 ;
	    RECT 1245.0000 1037.4000 1246.2001 1037.5500 ;
	    RECT 1240.8000 1034.4000 1242.3000 1035.3000 ;
	    RECT 1239.0000 1032.6000 1239.9000 1033.5000 ;
	    RECT 1239.0000 1031.4000 1240.2001 1032.6000 ;
	    RECT 1238.7001 1023.3000 1239.9000 1029.3000 ;
	    RECT 1241.1000 1023.3000 1242.3000 1034.4000 ;
	    RECT 1245.0000 1023.3000 1246.2001 1035.3000 ;
	    RECT 1259.4000 1023.3000 1260.6000 1029.3000 ;
	    RECT 1261.8000 1023.3000 1263.0000 1039.5000 ;
	    RECT 1288.2001 1037.4000 1289.4000 1038.6000 ;
	    RECT 1290.3000 1035.3000 1291.2001 1040.4000 ;
	    RECT 1360.2001 1040.1000 1364.4000 1040.4000 ;
	    RECT 1363.2001 1039.8000 1364.4000 1040.1000 ;
	    RECT 1365.3000 1040.4000 1366.8000 1041.3000 ;
	    RECT 1368.0000 1041.6000 1368.9000 1042.2001 ;
	    RECT 1368.0000 1040.4000 1369.2001 1041.6000 ;
	    RECT 1371.0000 1040.4000 1371.3000 1041.6000 ;
	    RECT 1372.2001 1041.4501 1373.4000 1041.6000 ;
	    RECT 1429.8000 1041.4501 1431.0000 1041.6000 ;
	    RECT 1372.2001 1040.5500 1431.0000 1041.4501 ;
	    RECT 1372.2001 1040.4000 1373.4000 1040.5500 ;
	    RECT 1429.8000 1040.4000 1431.0000 1040.5500 ;
	    RECT 1365.3000 1039.5000 1366.2001 1040.4000 ;
	    RECT 1285.8000 1023.3000 1287.0000 1035.3000 ;
	    RECT 1289.7001 1034.4000 1291.2001 1035.3000 ;
	    RECT 1293.0000 1035.4501 1294.2001 1035.6000 ;
	    RECT 1297.8000 1035.4501 1299.0000 1035.6000 ;
	    RECT 1293.0000 1034.5500 1299.0000 1035.4501 ;
	    RECT 1293.0000 1034.4000 1294.2001 1034.5500 ;
	    RECT 1297.8000 1034.4000 1299.0000 1034.5500 ;
	    RECT 1289.7001 1023.3000 1290.9000 1034.4000 ;
	    RECT 1292.1000 1032.6000 1293.0000 1033.5000 ;
	    RECT 1291.8000 1031.4000 1293.0000 1032.6000 ;
	    RECT 1292.1000 1023.3000 1293.3000 1029.3000 ;
	    RECT 1307.4000 1023.3000 1308.6000 1029.3000 ;
	    RECT 1309.8000 1023.3000 1311.0000 1039.5000 ;
	    RECT 1361.1000 1038.3000 1362.3000 1038.6000 ;
	    RECT 1365.0000 1038.4501 1366.2001 1038.6000 ;
	    RECT 1386.6000 1038.4501 1387.8000 1038.6000 ;
	    RECT 1361.1000 1037.4000 1363.5000 1038.3000 ;
	    RECT 1365.0000 1037.5500 1387.8000 1038.4501 ;
	    RECT 1365.0000 1037.4000 1366.2001 1037.5500 ;
	    RECT 1386.6000 1037.4000 1387.8000 1037.5500 ;
	    RECT 1362.3000 1037.1000 1363.5000 1037.4000 ;
	    RECT 1365.3000 1035.3000 1366.2001 1036.5000 ;
	    RECT 1499.1000 1036.2001 1500.3000 1042.8000 ;
	    RECT 1501.8000 1041.9000 1503.0000 1049.7001 ;
	    RECT 1506.6000 1043.7001 1507.8000 1049.7001 ;
	    RECT 1511.4000 1044.9000 1512.6000 1049.7001 ;
	    RECT 1513.8000 1045.5000 1515.0000 1049.7001 ;
	    RECT 1516.2001 1045.5000 1517.4000 1049.7001 ;
	    RECT 1518.6000 1045.5000 1519.8000 1049.7001 ;
	    RECT 1521.0000 1045.5000 1522.2001 1049.7001 ;
	    RECT 1523.4000 1046.7001 1524.6000 1049.7001 ;
	    RECT 1525.8000 1045.5000 1527.0000 1049.7001 ;
	    RECT 1528.2001 1046.7001 1529.4000 1049.7001 ;
	    RECT 1530.6000 1045.5000 1531.8000 1049.7001 ;
	    RECT 1533.0000 1045.5000 1534.2001 1049.7001 ;
	    RECT 1535.4000 1045.5000 1536.6000 1049.7001 ;
	    RECT 1509.0000 1043.7001 1512.6000 1044.9000 ;
	    RECT 1537.8000 1044.9000 1539.0000 1049.7001 ;
	    RECT 1509.0000 1042.8000 1510.2001 1043.7001 ;
	    RECT 1501.2001 1041.0000 1503.0000 1041.9000 ;
	    RECT 1507.5000 1041.9000 1510.2001 1042.8000 ;
	    RECT 1516.2001 1043.4000 1517.7001 1044.6000 ;
	    RECT 1522.2001 1043.4000 1522.5000 1044.6000 ;
	    RECT 1523.4000 1043.4000 1524.6000 1044.6000 ;
	    RECT 1525.8000 1043.7001 1532.7001 1044.6000 ;
	    RECT 1537.8000 1043.7001 1541.7001 1044.9000 ;
	    RECT 1542.6000 1043.7001 1543.8000 1049.7001 ;
	    RECT 1525.8000 1043.4000 1527.0000 1043.7001 ;
	    RECT 1501.2001 1038.0000 1502.1000 1041.0000 ;
	    RECT 1507.5000 1040.1000 1508.7001 1041.9000 ;
	    RECT 1503.0000 1038.9000 1508.7001 1040.1000 ;
	    RECT 1516.2001 1039.2001 1517.4000 1043.4000 ;
	    RECT 1528.2001 1042.5000 1529.4000 1042.8000 ;
	    RECT 1525.8000 1042.2001 1527.0000 1042.5000 ;
	    RECT 1520.4000 1041.3000 1527.0000 1042.2001 ;
	    RECT 1520.4000 1041.0000 1521.6000 1041.3000 ;
	    RECT 1528.2001 1040.4000 1529.4000 1041.6000 ;
	    RECT 1531.5000 1040.1000 1532.7001 1043.7001 ;
	    RECT 1540.5000 1042.8000 1541.7001 1043.7001 ;
	    RECT 1540.5000 1041.6000 1545.0000 1042.8000 ;
	    RECT 1547.4000 1040.7001 1548.6000 1049.7001 ;
	    RECT 1521.0000 1038.9000 1525.8000 1040.1000 ;
	    RECT 1531.5000 1038.9000 1534.5000 1040.1000 ;
	    RECT 1535.4000 1039.5000 1548.6000 1040.7001 ;
	    RECT 1511.4000 1038.0000 1512.6000 1038.9000 ;
	    RECT 1501.2001 1037.1000 1502.4000 1038.0000 ;
	    RECT 1511.4000 1037.1000 1536.9000 1038.0000 ;
	    RECT 1537.8000 1037.4000 1539.0000 1038.6000 ;
	    RECT 1545.3000 1038.0000 1546.5000 1038.3000 ;
	    RECT 1539.9000 1037.1000 1546.5000 1038.0000 ;
	    RECT 1357.8000 1034.4000 1361.7001 1035.3000 ;
	    RECT 1357.8000 1023.3000 1359.0000 1034.4000 ;
	    RECT 1360.5000 1034.1000 1361.7001 1034.4000 ;
	    RECT 1360.2001 1023.3000 1361.7001 1033.2001 ;
	    RECT 1364.4000 1023.3000 1366.8000 1035.3000 ;
	    RECT 1369.8000 1034.4000 1373.4000 1035.3000 ;
	    RECT 1499.1000 1035.0000 1500.6000 1036.2001 ;
	    RECT 1369.8000 1034.1000 1371.0000 1034.4000 ;
	    RECT 1369.5000 1023.3000 1371.0000 1033.2001 ;
	    RECT 1372.2001 1023.3000 1373.4000 1034.4000 ;
	    RECT 1499.4000 1033.5000 1500.6000 1035.0000 ;
	    RECT 1501.5000 1034.4000 1502.4000 1037.1000 ;
	    RECT 1503.3000 1036.2001 1504.5000 1036.5000 ;
	    RECT 1503.3000 1035.3000 1541.7001 1036.2001 ;
	    RECT 1542.6000 1035.4501 1543.8000 1035.6000 ;
	    RECT 1545.0000 1035.4501 1546.2001 1035.6000 ;
	    RECT 1537.5000 1035.0000 1538.7001 1035.3000 ;
	    RECT 1542.6000 1034.5500 1546.2001 1035.4501 ;
	    RECT 1542.6000 1034.4000 1543.8000 1034.5500 ;
	    RECT 1545.0000 1034.4000 1546.2001 1034.5500 ;
	    RECT 1501.5000 1033.5000 1515.0000 1034.4000 ;
	    RECT 1427.4000 1032.4501 1428.6000 1032.6000 ;
	    RECT 1499.4000 1032.4501 1500.6000 1032.6000 ;
	    RECT 1427.4000 1031.5500 1500.6000 1032.4501 ;
	    RECT 1427.4000 1031.4000 1428.6000 1031.5500 ;
	    RECT 1499.4000 1031.4000 1500.6000 1031.5500 ;
	    RECT 1501.5000 1031.1000 1502.4000 1033.5000 ;
	    RECT 1513.8000 1033.2001 1515.0000 1033.5000 ;
	    RECT 1518.6000 1033.5000 1531.5000 1034.4000 ;
	    RECT 1518.6000 1033.2001 1519.8000 1033.5000 ;
	    RECT 1506.3000 1031.4000 1510.2001 1032.6000 ;
	    RECT 1497.0000 1023.3000 1498.2001 1029.3000 ;
	    RECT 1499.4000 1023.3000 1500.6000 1030.5000 ;
	    RECT 1501.5000 1030.2001 1505.4000 1031.1000 ;
	    RECT 1501.8000 1023.3000 1503.0000 1029.3000 ;
	    RECT 1504.2001 1023.3000 1505.4000 1030.2001 ;
	    RECT 1506.6000 1023.3000 1507.8000 1029.3000 ;
	    RECT 1509.0000 1023.3000 1510.2001 1031.4000 ;
	    RECT 1511.1000 1030.2001 1517.4000 1031.4000 ;
	    RECT 1511.4000 1023.3000 1512.6000 1029.3000 ;
	    RECT 1513.8000 1023.3000 1515.0000 1027.5000 ;
	    RECT 1516.2001 1023.3000 1517.4000 1027.5000 ;
	    RECT 1518.6000 1023.3000 1519.8000 1027.5000 ;
	    RECT 1521.0000 1023.3000 1522.2001 1032.6000 ;
	    RECT 1525.8000 1031.4000 1529.7001 1032.6000 ;
	    RECT 1530.6000 1032.3000 1531.5000 1033.5000 ;
	    RECT 1533.0000 1034.1000 1534.2001 1034.4000 ;
	    RECT 1533.0000 1033.5000 1541.1000 1034.1000 ;
	    RECT 1533.0000 1033.2001 1542.3000 1033.5000 ;
	    RECT 1540.2001 1032.3000 1542.3000 1033.2001 ;
	    RECT 1530.6000 1031.4000 1539.3000 1032.3000 ;
	    RECT 1543.8000 1032.0000 1546.2001 1033.2001 ;
	    RECT 1543.8000 1031.4000 1544.7001 1032.0000 ;
	    RECT 1523.4000 1023.3000 1524.6000 1029.3000 ;
	    RECT 1525.8000 1023.3000 1527.0000 1030.5000 ;
	    RECT 1528.2001 1023.3000 1529.4000 1029.3000 ;
	    RECT 1530.6000 1023.3000 1531.8000 1030.5000 ;
	    RECT 1538.4000 1030.2001 1544.7001 1031.4000 ;
	    RECT 1547.4000 1031.1000 1548.6000 1039.5000 ;
	    RECT 1545.6000 1030.2001 1548.6000 1031.1000 ;
	    RECT 1533.0000 1023.3000 1534.2001 1027.5000 ;
	    RECT 1535.4000 1023.3000 1536.6000 1027.5000 ;
	    RECT 1537.8000 1023.3000 1539.0000 1029.3000 ;
	    RECT 1540.2001 1023.3000 1541.4000 1030.2001 ;
	    RECT 1545.6000 1029.3000 1546.5000 1030.2001 ;
	    RECT 1542.6000 1022.4000 1543.8000 1029.3000 ;
	    RECT 1545.0000 1028.4000 1546.5000 1029.3000 ;
	    RECT 1545.0000 1023.3000 1546.2001 1028.4000 ;
	    RECT 1547.4000 1023.3000 1548.6000 1029.3000 ;
	    RECT 1566.6000 1025.4000 1567.8000 1026.6000 ;
	    RECT 1566.7500 1022.4000 1567.6500 1025.4000 ;
	    RECT 1.2000 1020.6000 1569.0000 1022.4000 ;
	    RECT 126.6000 1013.7000 127.8000 1019.7000 ;
	    RECT 129.0000 1014.6000 130.2000 1019.7000 ;
	    RECT 128.7000 1013.7000 130.2000 1014.6000 ;
	    RECT 131.4000 1013.7000 132.6000 1020.6000 ;
	    RECT 128.7000 1012.8000 129.6000 1013.7000 ;
	    RECT 133.8000 1012.8000 135.0000 1019.7000 ;
	    RECT 136.2000 1013.7000 137.4000 1019.7000 ;
	    RECT 138.6000 1015.5000 139.8000 1019.7000 ;
	    RECT 141.0000 1015.5000 142.2000 1019.7000 ;
	    RECT 126.6000 1011.9000 129.6000 1012.8000 ;
	    RECT 126.6000 1003.5000 127.8000 1011.9000 ;
	    RECT 130.5000 1011.6000 136.8000 1012.8000 ;
	    RECT 143.4000 1012.5000 144.6000 1019.7000 ;
	    RECT 145.8000 1013.7000 147.0000 1019.7000 ;
	    RECT 148.2000 1012.5000 149.4000 1019.7000 ;
	    RECT 150.6000 1013.7000 151.8000 1019.7000 ;
	    RECT 130.5000 1011.0000 131.4000 1011.6000 ;
	    RECT 129.0000 1009.8000 131.4000 1011.0000 ;
	    RECT 135.9000 1010.7000 144.6000 1011.6000 ;
	    RECT 132.9000 1009.8000 135.0000 1010.7000 ;
	    RECT 132.9000 1009.5000 142.2000 1009.8000 ;
	    RECT 134.1000 1008.9000 142.2000 1009.5000 ;
	    RECT 141.0000 1008.6000 142.2000 1008.9000 ;
	    RECT 143.7000 1009.5000 144.6000 1010.7000 ;
	    RECT 145.5000 1010.4000 149.4000 1011.6000 ;
	    RECT 153.0000 1010.4000 154.2000 1019.7000 ;
	    RECT 155.4000 1015.5000 156.6000 1019.7000 ;
	    RECT 157.8000 1015.5000 159.0000 1019.7000 ;
	    RECT 160.2000 1015.5000 161.4000 1019.7000 ;
	    RECT 162.6000 1013.7000 163.8000 1019.7000 ;
	    RECT 157.8000 1011.6000 164.1000 1012.8000 ;
	    RECT 165.0000 1011.6000 166.2000 1019.7000 ;
	    RECT 167.4000 1013.7000 168.6000 1019.7000 ;
	    RECT 169.8000 1012.8000 171.0000 1019.7000 ;
	    RECT 172.2000 1013.7000 173.4000 1019.7000 ;
	    RECT 169.8000 1011.9000 173.7000 1012.8000 ;
	    RECT 174.6000 1012.5000 175.8000 1019.7000 ;
	    RECT 177.0000 1013.7000 178.2000 1019.7000 ;
	    RECT 191.4000 1013.7000 192.6000 1019.7000 ;
	    RECT 165.0000 1010.4000 168.9000 1011.6000 ;
	    RECT 155.4000 1009.5000 156.6000 1009.8000 ;
	    RECT 143.7000 1008.6000 156.6000 1009.5000 ;
	    RECT 160.2000 1009.5000 161.4000 1009.8000 ;
	    RECT 172.8000 1009.5000 173.7000 1011.9000 ;
	    RECT 174.6000 1011.4500 175.8000 1011.6000 ;
	    RECT 177.0000 1011.4500 178.2000 1011.6000 ;
	    RECT 174.6000 1010.5500 178.2000 1011.4500 ;
	    RECT 174.6000 1010.4000 175.8000 1010.5500 ;
	    RECT 177.0000 1010.4000 178.2000 1010.5500 ;
	    RECT 160.2000 1008.6000 173.7000 1009.5000 ;
	    RECT 131.4000 1007.4000 132.6000 1008.6000 ;
	    RECT 136.5000 1007.7000 137.7000 1008.0000 ;
	    RECT 133.5000 1006.8000 171.9000 1007.7000 ;
	    RECT 170.7000 1006.5000 171.9000 1006.8000 ;
	    RECT 172.8000 1005.9000 173.7000 1008.6000 ;
	    RECT 174.6000 1008.0000 175.8000 1009.5000 ;
	    RECT 174.6000 1006.8000 176.1000 1008.0000 ;
	    RECT 128.7000 1005.0000 135.3000 1005.9000 ;
	    RECT 128.7000 1004.7000 129.9000 1005.0000 ;
	    RECT 136.2000 1004.4000 137.4000 1005.6000 ;
	    RECT 138.3000 1005.0000 163.8000 1005.9000 ;
	    RECT 172.8000 1005.0000 174.0000 1005.9000 ;
	    RECT 162.6000 1004.1000 163.8000 1005.0000 ;
	    RECT 126.6000 1002.3000 139.8000 1003.5000 ;
	    RECT 140.7000 1002.9000 143.7000 1004.1000 ;
	    RECT 149.4000 1002.9000 154.2000 1004.1000 ;
	    RECT 126.6000 993.3000 127.8000 1002.3000 ;
	    RECT 130.2000 1000.2000 134.7000 1001.4000 ;
	    RECT 133.5000 999.3000 134.7000 1000.2000 ;
	    RECT 142.5000 999.3000 143.7000 1002.9000 ;
	    RECT 145.8000 1001.4000 147.0000 1002.6000 ;
	    RECT 153.6000 1001.7000 154.8000 1002.0000 ;
	    RECT 148.2000 1000.8000 154.8000 1001.7000 ;
	    RECT 148.2000 1000.5000 149.4000 1000.8000 ;
	    RECT 145.8000 1000.2000 147.0000 1000.5000 ;
	    RECT 157.8000 999.6000 159.0000 1003.8000 ;
	    RECT 166.5000 1002.9000 172.2000 1004.1000 ;
	    RECT 166.5000 1001.1000 167.7000 1002.9000 ;
	    RECT 173.1000 1002.0000 174.0000 1005.0000 ;
	    RECT 148.2000 999.3000 149.4000 999.6000 ;
	    RECT 131.4000 993.3000 132.6000 999.3000 ;
	    RECT 133.5000 998.1000 137.4000 999.3000 ;
	    RECT 142.5000 998.4000 149.4000 999.3000 ;
	    RECT 150.6000 998.4000 151.8000 999.6000 ;
	    RECT 152.7000 998.4000 153.0000 999.6000 ;
	    RECT 157.5000 998.4000 159.0000 999.6000 ;
	    RECT 165.0000 1000.2000 167.7000 1001.1000 ;
	    RECT 172.2000 1001.1000 174.0000 1002.0000 ;
	    RECT 165.0000 999.3000 166.2000 1000.2000 ;
	    RECT 136.2000 993.3000 137.4000 998.1000 ;
	    RECT 162.6000 998.1000 166.2000 999.3000 ;
	    RECT 138.6000 993.3000 139.8000 997.5000 ;
	    RECT 141.0000 993.3000 142.2000 997.5000 ;
	    RECT 143.4000 993.3000 144.6000 997.5000 ;
	    RECT 145.8000 993.3000 147.0000 996.3000 ;
	    RECT 148.2000 993.3000 149.4000 997.5000 ;
	    RECT 150.6000 993.3000 151.8000 996.3000 ;
	    RECT 153.0000 993.3000 154.2000 997.5000 ;
	    RECT 155.4000 993.3000 156.6000 997.5000 ;
	    RECT 157.8000 993.3000 159.0000 997.5000 ;
	    RECT 160.2000 993.3000 161.4000 997.5000 ;
	    RECT 162.6000 993.3000 163.8000 998.1000 ;
	    RECT 167.4000 993.3000 168.6000 999.3000 ;
	    RECT 172.2000 993.3000 173.4000 1001.1000 ;
	    RECT 174.9000 1000.2000 176.1000 1006.8000 ;
	    RECT 193.8000 1003.5000 195.0000 1019.7000 ;
	    RECT 232.2000 1007.7000 233.4000 1019.7000 ;
	    RECT 236.1000 1007.7000 239.1000 1019.7000 ;
	    RECT 241.8000 1007.7000 243.0000 1019.7000 ;
	    RECT 232.2000 1005.4500 233.4000 1005.6000 ;
	    RECT 234.6000 1005.4500 235.8000 1005.6000 ;
	    RECT 232.2000 1004.5500 235.8000 1005.4500 ;
	    RECT 232.2000 1004.4000 233.4000 1004.5500 ;
	    RECT 234.6000 1004.4000 235.8000 1004.5500 ;
	    RECT 237.0000 1003.5000 237.9000 1007.7000 ;
	    RECT 239.4000 1004.4000 240.6000 1005.6000 ;
	    RECT 241.8000 1003.5000 243.0000 1003.8000 ;
	    RECT 256.2000 1003.5000 257.4000 1019.7000 ;
	    RECT 258.6000 1013.7000 259.8000 1019.7000 ;
	    RECT 289.8000 1007.7000 291.0000 1019.7000 ;
	    RECT 293.7000 1007.7000 296.7000 1019.7000 ;
	    RECT 299.4000 1007.7000 300.6000 1019.7000 ;
	    RECT 292.2000 1004.4000 293.4000 1005.6000 ;
	    RECT 289.8000 1003.5000 291.0000 1003.8000 ;
	    RECT 294.9000 1003.5000 295.8000 1007.7000 ;
	    RECT 297.0000 1005.4500 298.2000 1005.6000 ;
	    RECT 306.6000 1005.4500 307.8000 1005.6000 ;
	    RECT 311.4000 1005.4500 312.6000 1005.6000 ;
	    RECT 297.0000 1004.5500 312.6000 1005.4500 ;
	    RECT 297.0000 1004.4000 298.2000 1004.5500 ;
	    RECT 306.6000 1004.4000 307.8000 1004.5500 ;
	    RECT 311.4000 1004.4000 312.6000 1004.5500 ;
	    RECT 313.8000 1003.5000 315.0000 1019.7000 ;
	    RECT 316.2000 1013.7000 317.4000 1019.7000 ;
	    RECT 448.2000 1013.7000 449.4000 1019.7000 ;
	    RECT 450.6000 1014.6000 451.8000 1019.7000 ;
	    RECT 450.3000 1013.7000 451.8000 1014.6000 ;
	    RECT 453.0000 1013.7000 454.2000 1020.6000 ;
	    RECT 450.3000 1012.8000 451.2000 1013.7000 ;
	    RECT 455.4000 1012.8000 456.6000 1019.7000 ;
	    RECT 457.8000 1013.7000 459.0000 1019.7000 ;
	    RECT 460.2000 1015.5000 461.4000 1019.7000 ;
	    RECT 462.6000 1015.5000 463.8000 1019.7000 ;
	    RECT 448.2000 1011.9000 451.2000 1012.8000 ;
	    RECT 448.2000 1003.5000 449.4000 1011.9000 ;
	    RECT 452.1000 1011.6000 458.4000 1012.8000 ;
	    RECT 465.0000 1012.5000 466.2000 1019.7000 ;
	    RECT 467.4000 1013.7000 468.6000 1019.7000 ;
	    RECT 469.8000 1012.5000 471.0000 1019.7000 ;
	    RECT 472.2000 1013.7000 473.4000 1019.7000 ;
	    RECT 452.1000 1011.0000 453.0000 1011.6000 ;
	    RECT 450.6000 1009.8000 453.0000 1011.0000 ;
	    RECT 457.5000 1010.7000 466.2000 1011.6000 ;
	    RECT 454.5000 1009.8000 456.6000 1010.7000 ;
	    RECT 454.5000 1009.5000 463.8000 1009.8000 ;
	    RECT 455.7000 1008.9000 463.8000 1009.5000 ;
	    RECT 462.6000 1008.6000 463.8000 1008.9000 ;
	    RECT 465.3000 1009.5000 466.2000 1010.7000 ;
	    RECT 467.1000 1010.4000 471.0000 1011.6000 ;
	    RECT 474.6000 1010.4000 475.8000 1019.7000 ;
	    RECT 477.0000 1015.5000 478.2000 1019.7000 ;
	    RECT 479.4000 1015.5000 480.6000 1019.7000 ;
	    RECT 481.8000 1015.5000 483.0000 1019.7000 ;
	    RECT 484.2000 1013.7000 485.4000 1019.7000 ;
	    RECT 479.4000 1011.6000 485.7000 1012.8000 ;
	    RECT 486.6000 1011.6000 487.8000 1019.7000 ;
	    RECT 489.0000 1013.7000 490.2000 1019.7000 ;
	    RECT 491.4000 1012.8000 492.6000 1019.7000 ;
	    RECT 493.8000 1013.7000 495.0000 1019.7000 ;
	    RECT 491.4000 1011.9000 495.3000 1012.8000 ;
	    RECT 496.2000 1012.5000 497.4000 1019.7000 ;
	    RECT 498.6000 1013.7000 499.8000 1019.7000 ;
	    RECT 510.6000 1013.7000 511.8000 1019.7000 ;
	    RECT 486.6000 1010.4000 490.5000 1011.6000 ;
	    RECT 477.0000 1009.5000 478.2000 1009.8000 ;
	    RECT 465.3000 1008.6000 478.2000 1009.5000 ;
	    RECT 481.8000 1009.5000 483.0000 1009.8000 ;
	    RECT 494.4000 1009.5000 495.3000 1011.9000 ;
	    RECT 496.2000 1010.4000 497.4000 1011.6000 ;
	    RECT 481.8000 1008.6000 495.3000 1009.5000 ;
	    RECT 453.0000 1007.4000 454.2000 1008.6000 ;
	    RECT 458.1000 1007.7000 459.3000 1008.0000 ;
	    RECT 455.1000 1006.8000 493.5000 1007.7000 ;
	    RECT 492.3000 1006.5000 493.5000 1006.8000 ;
	    RECT 494.4000 1005.9000 495.3000 1008.6000 ;
	    RECT 496.2000 1008.0000 497.4000 1009.5000 ;
	    RECT 496.2000 1006.8000 497.7000 1008.0000 ;
	    RECT 450.3000 1005.0000 456.9000 1005.9000 ;
	    RECT 450.3000 1004.7000 451.5000 1005.0000 ;
	    RECT 457.8000 1004.4000 459.0000 1005.6000 ;
	    RECT 459.9000 1005.0000 485.4000 1005.9000 ;
	    RECT 494.4000 1005.0000 495.6000 1005.9000 ;
	    RECT 484.2000 1004.1000 485.4000 1005.0000 ;
	    RECT 234.6000 1003.2000 235.8000 1003.5000 ;
	    RECT 239.4000 1003.2000 240.6000 1003.5000 ;
	    RECT 292.2000 1003.2000 293.4000 1003.5000 ;
	    RECT 297.0000 1003.2000 298.2000 1003.5000 ;
	    RECT 193.8000 1002.4500 195.0000 1002.6000 ;
	    RECT 210.6000 1002.4500 211.8000 1002.6000 ;
	    RECT 193.8000 1001.5500 211.8000 1002.4500 ;
	    RECT 193.8000 1001.4000 195.0000 1001.5500 ;
	    RECT 210.6000 1001.4000 211.8000 1001.5500 ;
	    RECT 225.0000 1002.4500 226.2000 1002.6000 ;
	    RECT 232.2000 1002.4500 233.4000 1002.6000 ;
	    RECT 225.0000 1001.5500 233.4000 1002.4500 ;
	    RECT 225.0000 1001.4000 226.2000 1001.5500 ;
	    RECT 232.2000 1001.4000 233.4000 1001.5500 ;
	    RECT 234.3000 1000.8000 234.6000 1002.3000 ;
	    RECT 237.0000 1001.4000 238.2000 1002.6000 ;
	    RECT 241.8000 1002.4500 243.0000 1002.6000 ;
	    RECT 256.2000 1002.4500 257.4000 1002.6000 ;
	    RECT 239.1000 1001.4000 240.6000 1002.3000 ;
	    RECT 241.8000 1001.5500 257.4000 1002.4500 ;
	    RECT 241.8000 1001.4000 243.0000 1001.5500 ;
	    RECT 256.2000 1001.4000 257.4000 1001.5500 ;
	    RECT 285.0000 1002.4500 286.2000 1002.6000 ;
	    RECT 289.8000 1002.4500 291.0000 1002.6000 ;
	    RECT 285.0000 1001.5500 291.0000 1002.4500 ;
	    RECT 285.0000 1001.4000 286.2000 1001.5500 ;
	    RECT 289.8000 1001.4000 291.0000 1001.5500 ;
	    RECT 292.2000 1001.4000 293.7000 1002.3000 ;
	    RECT 294.6000 1001.4000 295.8000 1002.6000 ;
	    RECT 299.4000 1002.4500 300.6000 1002.6000 ;
	    RECT 313.8000 1002.4500 315.0000 1002.6000 ;
	    RECT 174.6000 999.0000 176.1000 1000.2000 ;
	    RECT 174.6000 993.3000 175.8000 999.0000 ;
	    RECT 191.4000 998.4000 192.6000 999.6000 ;
	    RECT 191.4000 997.2000 192.6000 997.5000 ;
	    RECT 177.0000 993.3000 178.2000 996.3000 ;
	    RECT 191.4000 993.3000 192.6000 996.3000 ;
	    RECT 193.8000 993.3000 195.0000 1000.5000 ;
	    RECT 232.5000 999.3000 237.9000 999.9000 ;
	    RECT 239.7000 999.3000 240.6000 1001.4000 ;
	    RECT 232.2000 999.0000 238.2000 999.3000 ;
	    RECT 232.2000 993.3000 233.4000 999.0000 ;
	    RECT 234.6000 993.3000 235.8000 998.1000 ;
	    RECT 237.0000 994.2000 238.2000 999.0000 ;
	    RECT 239.4000 995.1000 240.6000 999.3000 ;
	    RECT 241.8000 994.2000 243.0000 999.3000 ;
	    RECT 237.0000 993.3000 243.0000 994.2000 ;
	    RECT 256.2000 993.3000 257.4000 1000.5000 ;
	    RECT 258.6000 999.4500 259.8000 999.6000 ;
	    RECT 270.6000 999.4500 271.8000 999.6000 ;
	    RECT 258.6000 998.5500 271.8000 999.4500 ;
	    RECT 292.2000 999.3000 293.1000 1001.4000 ;
	    RECT 298.2000 1000.8000 298.5000 1002.3000 ;
	    RECT 299.4000 1001.5500 315.0000 1002.4500 ;
	    RECT 299.4000 1001.4000 300.6000 1001.5500 ;
	    RECT 313.8000 1001.4000 315.0000 1001.5500 ;
	    RECT 448.2000 1002.3000 461.4000 1003.5000 ;
	    RECT 462.3000 1002.9000 465.3000 1004.1000 ;
	    RECT 471.0000 1002.9000 475.8000 1004.1000 ;
	    RECT 294.9000 999.3000 300.3000 999.9000 ;
	    RECT 258.6000 998.4000 259.8000 998.5500 ;
	    RECT 270.6000 998.4000 271.8000 998.5500 ;
	    RECT 258.6000 997.2000 259.8000 997.5000 ;
	    RECT 258.6000 993.3000 259.8000 996.3000 ;
	    RECT 289.8000 994.2000 291.0000 999.3000 ;
	    RECT 292.2000 995.1000 293.4000 999.3000 ;
	    RECT 294.6000 999.0000 300.6000 999.3000 ;
	    RECT 294.6000 994.2000 295.8000 999.0000 ;
	    RECT 289.8000 993.3000 295.8000 994.2000 ;
	    RECT 297.0000 993.3000 298.2000 998.1000 ;
	    RECT 299.4000 993.3000 300.6000 999.0000 ;
	    RECT 313.8000 993.3000 315.0000 1000.5000 ;
	    RECT 316.2000 998.4000 317.4000 999.6000 ;
	    RECT 316.2000 997.2000 317.4000 997.5000 ;
	    RECT 316.2000 993.3000 317.4000 996.3000 ;
	    RECT 448.2000 993.3000 449.4000 1002.3000 ;
	    RECT 451.8000 1000.2000 456.3000 1001.4000 ;
	    RECT 455.1000 999.3000 456.3000 1000.2000 ;
	    RECT 464.1000 999.3000 465.3000 1002.9000 ;
	    RECT 467.4000 1001.4000 468.6000 1002.6000 ;
	    RECT 475.2000 1001.7000 476.4000 1002.0000 ;
	    RECT 469.8000 1000.8000 476.4000 1001.7000 ;
	    RECT 469.8000 1000.5000 471.0000 1000.8000 ;
	    RECT 467.4000 1000.2000 468.6000 1000.5000 ;
	    RECT 479.4000 999.6000 480.6000 1003.8000 ;
	    RECT 488.1000 1002.9000 493.8000 1004.1000 ;
	    RECT 488.1000 1001.1000 489.3000 1002.9000 ;
	    RECT 494.7000 1002.0000 495.6000 1005.0000 ;
	    RECT 469.8000 999.3000 471.0000 999.6000 ;
	    RECT 453.0000 993.3000 454.2000 999.3000 ;
	    RECT 455.1000 998.1000 459.0000 999.3000 ;
	    RECT 464.1000 998.4000 471.0000 999.3000 ;
	    RECT 472.2000 998.4000 473.4000 999.6000 ;
	    RECT 474.3000 998.4000 474.6000 999.6000 ;
	    RECT 479.1000 998.4000 480.6000 999.6000 ;
	    RECT 486.6000 1000.2000 489.3000 1001.1000 ;
	    RECT 493.8000 1001.1000 495.6000 1002.0000 ;
	    RECT 486.6000 999.3000 487.8000 1000.2000 ;
	    RECT 457.8000 993.3000 459.0000 998.1000 ;
	    RECT 484.2000 998.1000 487.8000 999.3000 ;
	    RECT 460.2000 993.3000 461.4000 997.5000 ;
	    RECT 462.6000 993.3000 463.8000 997.5000 ;
	    RECT 465.0000 993.3000 466.2000 997.5000 ;
	    RECT 467.4000 993.3000 468.6000 996.3000 ;
	    RECT 469.8000 993.3000 471.0000 997.5000 ;
	    RECT 472.2000 993.3000 473.4000 996.3000 ;
	    RECT 474.6000 993.3000 475.8000 997.5000 ;
	    RECT 477.0000 993.3000 478.2000 997.5000 ;
	    RECT 479.4000 993.3000 480.6000 997.5000 ;
	    RECT 481.8000 993.3000 483.0000 997.5000 ;
	    RECT 484.2000 993.3000 485.4000 998.1000 ;
	    RECT 489.0000 993.3000 490.2000 999.3000 ;
	    RECT 493.8000 993.3000 495.0000 1001.1000 ;
	    RECT 496.5000 1000.2000 497.7000 1006.8000 ;
	    RECT 513.0000 1003.5000 514.2000 1019.7000 ;
	    RECT 532.2000 1013.7000 533.4000 1019.7000 ;
	    RECT 532.2000 1009.5000 533.4000 1009.8000 ;
	    RECT 515.4000 1008.4500 516.6000 1008.6000 ;
	    RECT 532.2000 1008.4500 533.4000 1008.6000 ;
	    RECT 515.4000 1007.5500 533.4000 1008.4500 ;
	    RECT 515.4000 1007.4000 516.6000 1007.5500 ;
	    RECT 532.2000 1007.4000 533.4000 1007.5500 ;
	    RECT 534.6000 1006.5000 535.8000 1019.7000 ;
	    RECT 537.0000 1013.7000 538.2000 1019.7000 ;
	    RECT 561.9000 1013.7000 563.1000 1019.7000 ;
	    RECT 562.2000 1010.4000 563.4000 1011.6000 ;
	    RECT 562.2000 1009.5000 563.1000 1010.4000 ;
	    RECT 564.3000 1008.6000 565.5000 1019.7000 ;
	    RECT 561.0000 1007.4000 562.2000 1008.6000 ;
	    RECT 564.0000 1007.7000 565.5000 1008.6000 ;
	    RECT 568.2000 1007.7000 569.4000 1019.7000 ;
	    RECT 534.6000 1005.4500 535.8000 1005.6000 ;
	    RECT 561.1500 1005.4500 562.0500 1007.4000 ;
	    RECT 534.6000 1004.5500 562.0500 1005.4500 ;
	    RECT 534.6000 1004.4000 535.8000 1004.5500 ;
	    RECT 513.0000 1002.4500 514.2000 1002.6000 ;
	    RECT 532.2000 1002.4500 533.4000 1002.6000 ;
	    RECT 513.0000 1001.5500 533.4000 1002.4500 ;
	    RECT 513.0000 1001.4000 514.2000 1001.5500 ;
	    RECT 532.2000 1001.4000 533.4000 1001.5500 ;
	    RECT 496.2000 999.0000 497.7000 1000.2000 ;
	    RECT 496.2000 993.3000 497.4000 999.0000 ;
	    RECT 510.6000 998.4000 511.8000 999.6000 ;
	    RECT 510.6000 997.2000 511.8000 997.5000 ;
	    RECT 498.6000 993.3000 499.8000 996.3000 ;
	    RECT 510.6000 993.3000 511.8000 996.3000 ;
	    RECT 513.0000 993.3000 514.2000 1000.5000 ;
	    RECT 534.6000 999.3000 535.8000 1003.5000 ;
	    RECT 564.0000 1002.6000 564.9000 1007.7000 ;
	    RECT 565.8000 1005.4500 567.0000 1005.6000 ;
	    RECT 565.8000 1004.5500 571.6500 1005.4500 ;
	    RECT 565.8000 1004.4000 567.0000 1004.5500 ;
	    RECT 565.8000 1003.2000 567.0000 1003.5000 ;
	    RECT 537.0000 1001.4000 538.2000 1002.6000 ;
	    RECT 561.0000 1001.4000 562.2000 1002.6000 ;
	    RECT 563.1000 1001.4000 564.9000 1002.6000 ;
	    RECT 567.0000 1000.8000 567.3000 1002.3000 ;
	    RECT 568.2000 1001.4000 569.4000 1002.6000 ;
	    RECT 570.7500 1002.4500 571.6500 1004.5500 ;
	    RECT 582.6000 1003.5000 583.8000 1019.7000 ;
	    RECT 585.0000 1013.7000 586.2000 1019.7000 ;
	    RECT 625.8000 1008.6000 627.0000 1019.7000 ;
	    RECT 628.2000 1009.8000 629.7000 1019.7000 ;
	    RECT 628.2000 1008.6000 629.4000 1008.9000 ;
	    RECT 625.8000 1007.7000 629.4000 1008.6000 ;
	    RECT 632.4000 1007.7000 634.8000 1019.7000 ;
	    RECT 637.5000 1009.8000 639.0000 1019.7000 ;
	    RECT 637.5000 1008.6000 638.7000 1008.9000 ;
	    RECT 640.2000 1008.6000 641.4000 1019.7000 ;
	    RECT 671.4000 1013.7000 672.6000 1019.7000 ;
	    RECT 673.8000 1013.7000 675.0000 1019.7000 ;
	    RECT 676.2000 1014.3000 677.4000 1019.7000 ;
	    RECT 674.1000 1013.4000 675.0000 1013.7000 ;
	    RECT 678.6000 1013.7000 679.8000 1019.7000 ;
	    RECT 678.6000 1013.4000 679.5000 1013.7000 ;
	    RECT 674.1000 1012.5000 679.5000 1013.4000 ;
	    RECT 657.0000 1011.4500 658.2000 1011.6000 ;
	    RECT 676.2000 1011.4500 677.4000 1011.6000 ;
	    RECT 657.0000 1010.5500 677.4000 1011.4500 ;
	    RECT 657.0000 1010.4000 658.2000 1010.5500 ;
	    RECT 676.2000 1010.4000 677.4000 1010.5500 ;
	    RECT 678.6000 1009.5000 679.5000 1012.5000 ;
	    RECT 676.2000 1009.2000 677.4000 1009.5000 ;
	    RECT 721.8000 1008.6000 723.0000 1019.7000 ;
	    RECT 724.2000 1009.8000 725.7000 1019.7000 ;
	    RECT 723.9000 1008.6000 725.1000 1008.9000 ;
	    RECT 637.5000 1007.7000 641.4000 1008.6000 ;
	    RECT 671.4000 1008.4500 672.6000 1008.6000 ;
	    RECT 673.8000 1008.4500 675.0000 1008.6000 ;
	    RECT 633.0000 1006.5000 633.9000 1007.7000 ;
	    RECT 671.4000 1007.5500 675.0000 1008.4500 ;
	    RECT 671.4000 1007.4000 672.6000 1007.5500 ;
	    RECT 673.8000 1007.4000 675.0000 1007.5500 ;
	    RECT 678.6000 1008.4500 679.8000 1008.6000 ;
	    RECT 709.8000 1008.4500 711.0000 1008.6000 ;
	    RECT 678.6000 1007.5500 711.0000 1008.4500 ;
	    RECT 721.8000 1007.7000 725.1000 1008.6000 ;
	    RECT 728.4000 1008.6000 730.8000 1019.7000 ;
	    RECT 733.5000 1009.8000 735.0000 1019.7000 ;
	    RECT 733.8000 1008.6000 735.0000 1008.9000 ;
	    RECT 736.2000 1008.6000 737.4000 1019.7000 ;
	    RECT 763.5000 1013.7000 764.7000 1019.7000 ;
	    RECT 763.8000 1010.4000 765.0000 1011.6000 ;
	    RECT 763.8000 1009.5000 764.7000 1010.4000 ;
	    RECT 765.9000 1008.6000 767.1000 1019.7000 ;
	    RECT 728.4000 1007.7000 731.4000 1008.6000 ;
	    RECT 733.8000 1007.7000 737.4000 1008.6000 ;
	    RECT 760.2000 1008.4500 761.4000 1008.6000 ;
	    RECT 762.6000 1008.4500 763.8000 1008.6000 ;
	    RECT 678.6000 1007.4000 679.8000 1007.5500 ;
	    RECT 709.8000 1007.4000 711.0000 1007.5500 ;
	    RECT 724.2000 1006.8000 725.1000 1007.7000 ;
	    RECT 671.4000 1006.2000 672.6000 1006.5000 ;
	    RECT 635.7000 1005.6000 636.9000 1005.9000 ;
	    RECT 630.6000 1005.4500 631.8000 1005.6000 ;
	    RECT 633.0000 1005.4500 634.2000 1005.6000 ;
	    RECT 630.6000 1004.5500 634.2000 1005.4500 ;
	    RECT 635.7000 1004.7000 638.1000 1005.6000 ;
	    RECT 630.6000 1004.4000 631.8000 1004.5500 ;
	    RECT 633.0000 1004.4000 634.2000 1004.5500 ;
	    RECT 636.9000 1004.4000 638.1000 1004.7000 ;
	    RECT 673.8000 1004.4000 675.0000 1005.6000 ;
	    RECT 675.9000 1004.4000 676.2000 1005.6000 ;
	    RECT 633.0000 1002.6000 633.9000 1003.5000 ;
	    RECT 582.6000 1002.4500 583.8000 1002.6000 ;
	    RECT 570.7500 1001.5500 583.8000 1002.4500 ;
	    RECT 582.6000 1001.4000 583.8000 1001.5500 ;
	    RECT 601.8000 1002.4500 603.0000 1002.6000 ;
	    RECT 618.6000 1002.4500 619.8000 1002.6000 ;
	    RECT 625.8000 1002.4500 627.0000 1002.6000 ;
	    RECT 601.8000 1001.5500 627.0000 1002.4500 ;
	    RECT 601.8000 1001.4000 603.0000 1001.5500 ;
	    RECT 618.6000 1001.4000 619.8000 1001.5500 ;
	    RECT 625.8000 1001.4000 627.0000 1001.5500 ;
	    RECT 627.9000 1001.4000 628.2000 1002.6000 ;
	    RECT 630.0000 1001.4000 631.2000 1002.6000 ;
	    RECT 630.3000 1000.8000 631.2000 1001.4000 ;
	    RECT 632.4000 1001.7000 633.9000 1002.6000 ;
	    RECT 634.8000 1002.9000 636.0000 1003.2000 ;
	    RECT 634.8000 1002.6000 639.0000 1002.9000 ;
	    RECT 678.6000 1002.6000 679.5000 1006.5000 ;
	    RECT 724.2000 1005.9000 729.3000 1006.8000 ;
	    RECT 730.5000 1006.5000 731.4000 1007.7000 ;
	    RECT 760.2000 1007.5500 763.8000 1008.4500 ;
	    RECT 760.2000 1007.4000 761.4000 1007.5500 ;
	    RECT 762.6000 1007.4000 763.8000 1007.5500 ;
	    RECT 765.6000 1007.7000 767.1000 1008.6000 ;
	    RECT 769.8000 1007.7000 771.0000 1019.7000 ;
	    RECT 781.8000 1019.4000 783.0000 1020.6000 ;
	    RECT 728.1000 1005.6000 729.3000 1005.9000 ;
	    RECT 731.4000 1005.4500 732.6000 1005.6000 ;
	    RECT 748.2000 1005.4500 749.4000 1005.6000 ;
	    RECT 724.8000 1004.7000 726.0000 1005.0000 ;
	    RECT 724.8000 1003.8000 728.7000 1004.7000 ;
	    RECT 727.8000 1002.9000 728.7000 1003.8000 ;
	    RECT 729.9000 1003.5000 730.5000 1004.7000 ;
	    RECT 731.4000 1004.5500 749.4000 1005.4500 ;
	    RECT 731.4000 1004.4000 732.6000 1004.5500 ;
	    RECT 748.2000 1004.4000 749.4000 1004.5500 ;
	    RECT 634.8000 1002.0000 639.3000 1002.6000 ;
	    RECT 638.1000 1001.7000 639.3000 1002.0000 ;
	    RECT 537.0000 1000.2000 538.2000 1000.5000 ;
	    RECT 561.3000 999.3000 562.2000 1000.5000 ;
	    RECT 563.7000 999.3000 569.1000 999.9000 ;
	    RECT 533.1000 998.4000 535.8000 999.3000 ;
	    RECT 533.1000 993.3000 534.3000 998.4000 ;
	    RECT 537.0000 993.3000 538.2000 999.3000 ;
	    RECT 561.0000 993.3000 562.2000 999.3000 ;
	    RECT 563.4000 999.0000 569.4000 999.3000 ;
	    RECT 563.4000 993.3000 564.6000 999.0000 ;
	    RECT 565.8000 993.3000 567.0000 998.1000 ;
	    RECT 568.2000 993.3000 569.4000 999.0000 ;
	    RECT 582.6000 993.3000 583.8000 1000.5000 ;
	    RECT 628.2000 1000.2000 629.4000 1000.5000 ;
	    RECT 585.0000 999.4500 586.2000 999.6000 ;
	    RECT 623.4000 999.4500 624.6000 999.6000 ;
	    RECT 585.0000 998.5500 624.6000 999.4500 ;
	    RECT 585.0000 998.4000 586.2000 998.5500 ;
	    RECT 623.4000 998.4000 624.6000 998.5500 ;
	    RECT 625.8000 999.3000 629.4000 1000.2000 ;
	    RECT 630.3000 999.6000 631.5000 1000.8000 ;
	    RECT 585.0000 997.2000 586.2000 997.5000 ;
	    RECT 585.0000 993.3000 586.2000 996.3000 ;
	    RECT 625.8000 993.3000 627.0000 999.3000 ;
	    RECT 632.4000 998.7000 633.3000 1001.7000 ;
	    RECT 639.0000 1001.4000 639.3000 1001.7000 ;
	    RECT 640.2000 1002.4500 641.4000 1002.6000 ;
	    RECT 642.6000 1002.4500 643.8000 1002.6000 ;
	    RECT 640.2000 1001.5500 643.8000 1002.4500 ;
	    RECT 677.1000 1002.3000 679.5000 1002.6000 ;
	    RECT 640.2000 1001.4000 641.4000 1001.5500 ;
	    RECT 642.6000 1001.4000 643.8000 1001.5500 ;
	    RECT 634.2000 999.6000 636.6000 1000.8000 ;
	    RECT 637.5000 1000.2000 638.7000 1000.5000 ;
	    RECT 637.5000 999.3000 641.4000 1000.2000 ;
	    RECT 628.2000 993.3000 629.7000 998.4000 ;
	    RECT 632.4000 993.3000 634.8000 998.7000 ;
	    RECT 637.5000 993.3000 639.0000 998.4000 ;
	    RECT 640.2000 993.3000 641.4000 999.3000 ;
	    RECT 671.4000 993.3000 672.6000 1002.3000 ;
	    RECT 676.8000 1001.7000 679.5000 1002.3000 ;
	    RECT 719.4000 1002.4500 720.6000 1002.6000 ;
	    RECT 721.8000 1002.4500 723.0000 1002.6000 ;
	    RECT 676.8000 993.3000 678.0000 1001.7000 ;
	    RECT 719.4000 1001.5500 723.0000 1002.4500 ;
	    RECT 719.4000 1001.4000 720.6000 1001.5500 ;
	    RECT 721.8000 1001.4000 723.0000 1001.5500 ;
	    RECT 723.9000 1002.3000 724.2000 1002.6000 ;
	    RECT 723.9000 1001.4000 726.9000 1002.3000 ;
	    RECT 727.8000 1001.7000 729.0000 1002.9000 ;
	    RECT 726.0000 1000.8000 726.9000 1001.4000 ;
	    RECT 723.9000 1000.2000 725.1000 1000.5000 ;
	    RECT 721.8000 999.3000 725.1000 1000.2000 ;
	    RECT 726.0000 999.9000 729.0000 1000.8000 ;
	    RECT 726.6000 999.6000 729.0000 999.9000 ;
	    RECT 721.8000 993.3000 723.0000 999.3000 ;
	    RECT 729.9000 998.7000 730.8000 1003.5000 ;
	    RECT 765.6000 1002.6000 766.5000 1007.7000 ;
	    RECT 767.4000 1004.4000 768.6000 1005.6000 ;
	    RECT 784.2000 1003.5000 785.4000 1019.7000 ;
	    RECT 786.6000 1013.7000 787.8000 1019.7000 ;
	    RECT 837.0000 1017.4500 838.2000 1017.6000 ;
	    RECT 906.6000 1017.4500 907.8000 1017.6000 ;
	    RECT 837.0000 1016.5500 907.8000 1017.4500 ;
	    RECT 837.0000 1016.4000 838.2000 1016.5500 ;
	    RECT 906.6000 1016.4000 907.8000 1016.5500 ;
	    RECT 827.4000 1014.4500 828.6000 1014.6000 ;
	    RECT 901.8000 1014.4500 903.0000 1014.6000 ;
	    RECT 827.4000 1013.5500 903.0000 1014.4500 ;
	    RECT 921.0000 1013.7000 922.2000 1019.7000 ;
	    RECT 923.4000 1014.6000 924.6000 1019.7000 ;
	    RECT 923.1000 1013.7000 924.6000 1014.6000 ;
	    RECT 925.8000 1013.7000 927.0000 1020.6000 ;
	    RECT 827.4000 1013.4000 828.6000 1013.5500 ;
	    RECT 901.8000 1013.4000 903.0000 1013.5500 ;
	    RECT 923.1000 1012.8000 924.0000 1013.7000 ;
	    RECT 928.2000 1012.8000 929.4000 1019.7000 ;
	    RECT 930.6000 1013.7000 931.8000 1019.7000 ;
	    RECT 933.0000 1015.5000 934.2000 1019.7000 ;
	    RECT 935.4000 1015.5000 936.6000 1019.7000 ;
	    RECT 921.0000 1011.9000 924.0000 1012.8000 ;
	    RECT 921.0000 1003.5000 922.2000 1011.9000 ;
	    RECT 924.9000 1011.6000 931.2000 1012.8000 ;
	    RECT 937.8000 1012.5000 939.0000 1019.7000 ;
	    RECT 940.2000 1013.7000 941.4000 1019.7000 ;
	    RECT 942.6000 1012.5000 943.8000 1019.7000 ;
	    RECT 945.0000 1013.7000 946.2000 1019.7000 ;
	    RECT 924.9000 1011.0000 925.8000 1011.6000 ;
	    RECT 923.4000 1009.8000 925.8000 1011.0000 ;
	    RECT 930.3000 1010.7000 939.0000 1011.6000 ;
	    RECT 927.3000 1009.8000 929.4000 1010.7000 ;
	    RECT 927.3000 1009.5000 936.6000 1009.8000 ;
	    RECT 928.5000 1008.9000 936.6000 1009.5000 ;
	    RECT 935.4000 1008.6000 936.6000 1008.9000 ;
	    RECT 938.1000 1009.5000 939.0000 1010.7000 ;
	    RECT 939.9000 1010.4000 943.8000 1011.6000 ;
	    RECT 947.4000 1010.4000 948.6000 1019.7000 ;
	    RECT 949.8000 1015.5000 951.0000 1019.7000 ;
	    RECT 952.2000 1015.5000 953.4000 1019.7000 ;
	    RECT 954.6000 1015.5000 955.8000 1019.7000 ;
	    RECT 957.0000 1013.7000 958.2000 1019.7000 ;
	    RECT 952.2000 1011.6000 958.5000 1012.8000 ;
	    RECT 959.4000 1011.6000 960.6000 1019.7000 ;
	    RECT 961.8000 1013.7000 963.0000 1019.7000 ;
	    RECT 964.2000 1012.8000 965.4000 1019.7000 ;
	    RECT 966.6000 1013.7000 967.8000 1019.7000 ;
	    RECT 964.2000 1011.9000 968.1000 1012.8000 ;
	    RECT 969.0000 1012.5000 970.2000 1019.7000 ;
	    RECT 971.4000 1013.7000 972.6000 1019.7000 ;
	    RECT 959.4000 1010.4000 963.3000 1011.6000 ;
	    RECT 949.8000 1009.5000 951.0000 1009.8000 ;
	    RECT 938.1000 1008.6000 951.0000 1009.5000 ;
	    RECT 954.6000 1009.5000 955.8000 1009.8000 ;
	    RECT 967.2000 1009.5000 968.1000 1011.9000 ;
	    RECT 969.0000 1010.4000 970.2000 1011.6000 ;
	    RECT 954.6000 1008.6000 968.1000 1009.5000 ;
	    RECT 925.8000 1007.4000 927.0000 1008.6000 ;
	    RECT 930.9000 1007.7000 932.1000 1008.0000 ;
	    RECT 927.9000 1006.8000 966.3000 1007.7000 ;
	    RECT 965.1000 1006.5000 966.3000 1006.8000 ;
	    RECT 967.2000 1005.9000 968.1000 1008.6000 ;
	    RECT 969.0000 1008.0000 970.2000 1009.5000 ;
	    RECT 969.0000 1006.8000 970.5000 1008.0000 ;
	    RECT 923.1000 1005.0000 929.7000 1005.9000 ;
	    RECT 923.1000 1004.7000 924.3000 1005.0000 ;
	    RECT 930.6000 1004.4000 931.8000 1005.6000 ;
	    RECT 932.7000 1005.0000 958.2000 1005.9000 ;
	    RECT 967.2000 1005.0000 968.4000 1005.9000 ;
	    RECT 957.0000 1004.1000 958.2000 1005.0000 ;
	    RECT 767.4000 1003.2000 768.6000 1003.5000 ;
	    RECT 732.0000 1001.4000 733.2000 1002.6000 ;
	    RECT 735.0000 1001.4000 735.3000 1002.6000 ;
	    RECT 736.2000 1001.4000 737.4000 1002.6000 ;
	    RECT 762.6000 1001.4000 763.8000 1002.6000 ;
	    RECT 764.7000 1001.4000 766.5000 1002.6000 ;
	    RECT 769.8000 1002.4500 771.0000 1002.6000 ;
	    RECT 781.8000 1002.4500 783.0000 1002.6000 ;
	    RECT 732.0000 1000.8000 732.9000 1001.4000 ;
	    RECT 768.6000 1000.8000 768.9000 1002.3000 ;
	    RECT 769.8000 1001.5500 783.0000 1002.4500 ;
	    RECT 769.8000 1001.4000 771.0000 1001.5500 ;
	    RECT 781.8000 1001.4000 783.0000 1001.5500 ;
	    RECT 784.2000 1002.4500 785.4000 1002.6000 ;
	    RECT 858.6000 1002.4500 859.8000 1002.6000 ;
	    RECT 784.2000 1001.5500 859.8000 1002.4500 ;
	    RECT 784.2000 1001.4000 785.4000 1001.5500 ;
	    RECT 858.6000 1001.4000 859.8000 1001.5500 ;
	    RECT 921.0000 1002.3000 934.2000 1003.5000 ;
	    RECT 935.1000 1002.9000 938.1000 1004.1000 ;
	    RECT 943.8000 1002.9000 948.6000 1004.1000 ;
	    RECT 731.7000 999.6000 732.9000 1000.8000 ;
	    RECT 733.8000 1000.2000 735.0000 1000.5000 ;
	    RECT 733.8000 999.3000 737.4000 1000.2000 ;
	    RECT 762.9000 999.3000 763.8000 1000.5000 ;
	    RECT 765.3000 999.3000 770.7000 999.9000 ;
	    RECT 724.2000 993.3000 725.7000 998.4000 ;
	    RECT 728.4000 993.3000 730.8000 998.7000 ;
	    RECT 733.5000 993.3000 735.0000 998.4000 ;
	    RECT 736.2000 993.3000 737.4000 999.3000 ;
	    RECT 762.6000 993.3000 763.8000 999.3000 ;
	    RECT 765.0000 999.0000 771.0000 999.3000 ;
	    RECT 765.0000 993.3000 766.2000 999.0000 ;
	    RECT 767.4000 993.3000 768.6000 998.1000 ;
	    RECT 769.8000 993.3000 771.0000 999.0000 ;
	    RECT 784.2000 993.3000 785.4000 1000.5000 ;
	    RECT 786.6000 998.4000 787.8000 999.6000 ;
	    RECT 786.6000 997.2000 787.8000 997.5000 ;
	    RECT 892.2000 996.4500 893.4000 996.6000 ;
	    RECT 904.2000 996.4500 905.4000 996.6000 ;
	    RECT 916.2000 996.4500 917.4000 996.6000 ;
	    RECT 786.6000 993.3000 787.8000 996.3000 ;
	    RECT 892.2000 995.5500 917.4000 996.4500 ;
	    RECT 892.2000 995.4000 893.4000 995.5500 ;
	    RECT 904.2000 995.4000 905.4000 995.5500 ;
	    RECT 916.2000 995.4000 917.4000 995.5500 ;
	    RECT 921.0000 993.3000 922.2000 1002.3000 ;
	    RECT 924.6000 1000.2000 929.1000 1001.4000 ;
	    RECT 927.9000 999.3000 929.1000 1000.2000 ;
	    RECT 936.9000 999.3000 938.1000 1002.9000 ;
	    RECT 940.2000 1001.4000 941.4000 1002.6000 ;
	    RECT 948.0000 1001.7000 949.2000 1002.0000 ;
	    RECT 942.6000 1000.8000 949.2000 1001.7000 ;
	    RECT 942.6000 1000.5000 943.8000 1000.8000 ;
	    RECT 940.2000 1000.2000 941.4000 1000.5000 ;
	    RECT 952.2000 999.6000 953.4000 1003.8000 ;
	    RECT 960.9000 1002.9000 966.6000 1004.1000 ;
	    RECT 960.9000 1001.1000 962.1000 1002.9000 ;
	    RECT 967.5000 1002.0000 968.4000 1005.0000 ;
	    RECT 942.6000 999.3000 943.8000 999.6000 ;
	    RECT 925.8000 993.3000 927.0000 999.3000 ;
	    RECT 927.9000 998.1000 931.8000 999.3000 ;
	    RECT 936.9000 998.4000 943.8000 999.3000 ;
	    RECT 945.0000 998.4000 946.2000 999.6000 ;
	    RECT 947.1000 998.4000 947.4000 999.6000 ;
	    RECT 951.9000 998.4000 953.4000 999.6000 ;
	    RECT 959.4000 1000.2000 962.1000 1001.1000 ;
	    RECT 966.6000 1001.1000 968.4000 1002.0000 ;
	    RECT 959.4000 999.3000 960.6000 1000.2000 ;
	    RECT 930.6000 993.3000 931.8000 998.1000 ;
	    RECT 957.0000 998.1000 960.6000 999.3000 ;
	    RECT 933.0000 993.3000 934.2000 997.5000 ;
	    RECT 935.4000 993.3000 936.6000 997.5000 ;
	    RECT 937.8000 993.3000 939.0000 997.5000 ;
	    RECT 940.2000 993.3000 941.4000 996.3000 ;
	    RECT 942.6000 993.3000 943.8000 997.5000 ;
	    RECT 945.0000 993.3000 946.2000 996.3000 ;
	    RECT 947.4000 993.3000 948.6000 997.5000 ;
	    RECT 949.8000 993.3000 951.0000 997.5000 ;
	    RECT 952.2000 993.3000 953.4000 997.5000 ;
	    RECT 954.6000 993.3000 955.8000 997.5000 ;
	    RECT 957.0000 993.3000 958.2000 998.1000 ;
	    RECT 961.8000 993.3000 963.0000 999.3000 ;
	    RECT 966.6000 993.3000 967.8000 1001.1000 ;
	    RECT 969.3000 1000.2000 970.5000 1006.8000 ;
	    RECT 985.8000 1003.5000 987.0000 1019.7000 ;
	    RECT 988.2000 1013.7000 989.4000 1019.7000 ;
	    RECT 1013.1000 1013.7000 1014.3000 1019.7000 ;
	    RECT 1013.4000 1010.4000 1014.6000 1011.6000 ;
	    RECT 1013.4000 1009.5000 1014.3000 1010.4000 ;
	    RECT 1015.5000 1008.6000 1016.7000 1019.7000 ;
	    RECT 1000.2000 1008.4500 1001.4000 1008.6000 ;
	    RECT 1012.2000 1008.4500 1013.4000 1008.6000 ;
	    RECT 1000.2000 1007.5500 1013.4000 1008.4500 ;
	    RECT 1000.2000 1007.4000 1001.4000 1007.5500 ;
	    RECT 1012.2000 1007.4000 1013.4000 1007.5500 ;
	    RECT 1015.2000 1007.7000 1016.7000 1008.6000 ;
	    RECT 1019.4000 1007.7000 1020.6000 1019.7000 ;
	    RECT 1015.2000 1002.6000 1016.1000 1007.7000 ;
	    RECT 1017.0000 1005.4500 1018.2000 1005.6000 ;
	    RECT 1026.6000 1005.4500 1027.8000 1005.6000 ;
	    RECT 1017.0000 1004.5500 1027.8000 1005.4500 ;
	    RECT 1017.0000 1004.4000 1018.2000 1004.5500 ;
	    RECT 1026.6000 1004.4000 1027.8000 1004.5500 ;
	    RECT 1033.8000 1003.5000 1035.0000 1019.7000 ;
	    RECT 1036.2001 1013.7000 1037.4000 1019.7000 ;
	    RECT 1055.4000 1013.7000 1056.6000 1019.7000 ;
	    RECT 1055.4000 1009.5000 1056.6000 1009.8000 ;
	    RECT 1055.4000 1007.4000 1056.6000 1008.6000 ;
	    RECT 1057.8000 1006.5000 1059.0000 1019.7000 ;
	    RECT 1060.2001 1013.7000 1061.4000 1019.7000 ;
	    RECT 1192.2001 1013.7000 1193.4000 1019.7000 ;
	    RECT 1194.6000 1012.5000 1195.8000 1019.7000 ;
	    RECT 1197.0000 1013.7000 1198.2001 1019.7000 ;
	    RECT 1199.4000 1012.8000 1200.6000 1019.7000 ;
	    RECT 1201.8000 1013.7000 1203.0000 1019.7000 ;
	    RECT 1196.7001 1011.9000 1200.6000 1012.8000 ;
	    RECT 1163.4000 1011.4500 1164.6000 1011.6000 ;
	    RECT 1194.6000 1011.4500 1195.8000 1011.6000 ;
	    RECT 1163.4000 1010.5500 1195.8000 1011.4500 ;
	    RECT 1163.4000 1010.4000 1164.6000 1010.5500 ;
	    RECT 1194.6000 1010.4000 1195.8000 1010.5500 ;
	    RECT 1196.7001 1009.5000 1197.6000 1011.9000 ;
	    RECT 1204.2001 1011.6000 1205.4000 1019.7000 ;
	    RECT 1206.6000 1013.7000 1207.8000 1019.7000 ;
	    RECT 1209.0000 1015.5000 1210.2001 1019.7000 ;
	    RECT 1211.4000 1015.5000 1212.6000 1019.7000 ;
	    RECT 1213.8000 1015.5000 1215.0000 1019.7000 ;
	    RECT 1206.3000 1011.6000 1212.6000 1012.8000 ;
	    RECT 1201.5000 1010.4000 1205.4000 1011.6000 ;
	    RECT 1216.2001 1010.4000 1217.4000 1019.7000 ;
	    RECT 1218.6000 1013.7000 1219.8000 1019.7000 ;
	    RECT 1221.0000 1012.5000 1222.2001 1019.7000 ;
	    RECT 1223.4000 1013.7000 1224.6000 1019.7000 ;
	    RECT 1225.8000 1012.5000 1227.0000 1019.7000 ;
	    RECT 1228.2001 1015.5000 1229.4000 1019.7000 ;
	    RECT 1230.6000 1015.5000 1231.8000 1019.7000 ;
	    RECT 1233.0000 1013.7000 1234.2001 1019.7000 ;
	    RECT 1235.4000 1012.8000 1236.6000 1019.7000 ;
	    RECT 1237.8000 1013.7000 1239.0000 1020.6000 ;
	    RECT 1240.2001 1014.6000 1241.4000 1019.7000 ;
	    RECT 1240.2001 1013.7000 1241.7001 1014.6000 ;
	    RECT 1242.6000 1013.7000 1243.8000 1019.7000 ;
	    RECT 1261.8000 1013.7000 1263.0000 1019.7000 ;
	    RECT 1240.8000 1012.8000 1241.7001 1013.7000 ;
	    RECT 1233.6000 1011.6000 1239.9000 1012.8000 ;
	    RECT 1240.8000 1011.9000 1243.8000 1012.8000 ;
	    RECT 1221.0000 1010.4000 1224.9000 1011.6000 ;
	    RECT 1225.8000 1010.7000 1234.5000 1011.6000 ;
	    RECT 1239.0000 1011.0000 1239.9000 1011.6000 ;
	    RECT 1209.0000 1009.5000 1210.2001 1009.8000 ;
	    RECT 1194.6000 1008.0000 1195.8000 1009.5000 ;
	    RECT 1194.3000 1006.8000 1195.8000 1008.0000 ;
	    RECT 1196.7001 1008.6000 1210.2001 1009.5000 ;
	    RECT 1213.8000 1009.5000 1215.0000 1009.8000 ;
	    RECT 1225.8000 1009.5000 1226.7001 1010.7000 ;
	    RECT 1235.4000 1009.8000 1237.5000 1010.7000 ;
	    RECT 1239.0000 1009.8000 1241.4000 1011.0000 ;
	    RECT 1213.8000 1008.6000 1226.7001 1009.5000 ;
	    RECT 1228.2001 1009.5000 1237.5000 1009.8000 ;
	    RECT 1228.2001 1008.9000 1236.3000 1009.5000 ;
	    RECT 1228.2001 1008.6000 1229.4000 1008.9000 ;
	    RECT 1057.8000 1005.4500 1059.0000 1005.6000 ;
	    RECT 1093.8000 1005.4500 1095.0000 1005.6000 ;
	    RECT 1057.8000 1004.5500 1095.0000 1005.4500 ;
	    RECT 1057.8000 1004.4000 1059.0000 1004.5500 ;
	    RECT 1093.8000 1004.4000 1095.0000 1004.5500 ;
	    RECT 1017.0000 1003.2000 1018.2000 1003.5000 ;
	    RECT 985.8000 1002.4500 987.0000 1002.6000 ;
	    RECT 1009.8000 1002.4500 1011.0000 1002.6000 ;
	    RECT 985.8000 1001.5500 1011.0000 1002.4500 ;
	    RECT 985.8000 1001.4000 987.0000 1001.5500 ;
	    RECT 1009.8000 1001.4000 1011.0000 1001.5500 ;
	    RECT 1012.2000 1001.4000 1013.4000 1002.6000 ;
	    RECT 1014.3000 1001.4000 1016.1000 1002.6000 ;
	    RECT 1018.2000 1000.8000 1018.5000 1002.3000 ;
	    RECT 1019.4000 1001.4000 1020.6000 1002.6000 ;
	    RECT 1033.8000 1002.4500 1035.0000 1002.6000 ;
	    RECT 1036.2001 1002.4500 1037.4000 1002.6000 ;
	    RECT 1033.8000 1001.5500 1037.4000 1002.4500 ;
	    RECT 1033.8000 1001.4000 1035.0000 1001.5500 ;
	    RECT 1036.2001 1001.4000 1037.4000 1001.5500 ;
	    RECT 969.0000 999.0000 970.5000 1000.2000 ;
	    RECT 969.0000 993.3000 970.2000 999.0000 ;
	    RECT 971.4000 993.3000 972.6000 996.3000 ;
	    RECT 985.8000 993.3000 987.0000 1000.5000 ;
	    RECT 988.2000 999.4500 989.4000 999.6000 ;
	    RECT 990.6000 999.4500 991.8000 999.6000 ;
	    RECT 988.2000 998.5500 991.8000 999.4500 ;
	    RECT 1012.5000 999.3000 1013.4000 1000.5000 ;
	    RECT 1014.9000 999.3000 1020.3000 999.9000 ;
	    RECT 988.2000 998.4000 989.4000 998.5500 ;
	    RECT 990.6000 998.4000 991.8000 998.5500 ;
	    RECT 988.2000 997.2000 989.4000 997.5000 ;
	    RECT 988.2000 993.3000 989.4000 996.3000 ;
	    RECT 1012.2000 993.3000 1013.4000 999.3000 ;
	    RECT 1014.6000 999.0000 1020.6000 999.3000 ;
	    RECT 1014.6000 993.3000 1015.8000 999.0000 ;
	    RECT 1017.0000 993.3000 1018.2000 998.1000 ;
	    RECT 1019.4000 993.3000 1020.6000 999.0000 ;
	    RECT 1033.8000 993.3000 1035.0000 1000.5000 ;
	    RECT 1036.2001 999.4500 1037.4000 999.6000 ;
	    RECT 1038.6000 999.4500 1039.8000 999.6000 ;
	    RECT 1036.2001 998.5500 1039.8000 999.4500 ;
	    RECT 1057.8000 999.3000 1059.0000 1003.5000 ;
	    RECT 1060.2001 1001.4000 1061.4000 1002.6000 ;
	    RECT 1060.2001 1000.2000 1061.4000 1000.5000 ;
	    RECT 1194.3000 1000.2000 1195.5000 1006.8000 ;
	    RECT 1196.7001 1005.9000 1197.6000 1008.6000 ;
	    RECT 1232.7001 1007.7000 1233.9000 1008.0000 ;
	    RECT 1198.5000 1006.8000 1236.9000 1007.7000 ;
	    RECT 1237.8000 1007.4000 1239.0000 1008.6000 ;
	    RECT 1198.5000 1006.5000 1199.7001 1006.8000 ;
	    RECT 1196.4000 1005.0000 1197.6000 1005.9000 ;
	    RECT 1206.6000 1005.0000 1232.1000 1005.9000 ;
	    RECT 1196.4000 1002.0000 1197.3000 1005.0000 ;
	    RECT 1206.6000 1004.1000 1207.8000 1005.0000 ;
	    RECT 1233.0000 1004.4000 1234.2001 1005.6000 ;
	    RECT 1235.1000 1005.0000 1241.7001 1005.9000 ;
	    RECT 1240.5000 1004.7000 1241.7001 1005.0000 ;
	    RECT 1198.2001 1002.9000 1203.9000 1004.1000 ;
	    RECT 1196.4000 1001.1000 1198.2001 1002.0000 ;
	    RECT 1036.2001 998.4000 1037.4000 998.5500 ;
	    RECT 1038.6000 998.4000 1039.8000 998.5500 ;
	    RECT 1056.3000 998.4000 1059.0000 999.3000 ;
	    RECT 1036.2001 997.2000 1037.4000 997.5000 ;
	    RECT 1036.2001 993.3000 1037.4000 996.3000 ;
	    RECT 1056.3000 993.3000 1057.5000 998.4000 ;
	    RECT 1060.2001 993.3000 1061.4000 999.3000 ;
	    RECT 1194.3000 999.0000 1195.8000 1000.2000 ;
	    RECT 1062.6000 996.4500 1063.8000 996.6000 ;
	    RECT 1137.0000 996.4500 1138.2001 996.6000 ;
	    RECT 1062.6000 995.5500 1138.2001 996.4500 ;
	    RECT 1062.6000 995.4000 1063.8000 995.5500 ;
	    RECT 1137.0000 995.4000 1138.2001 995.5500 ;
	    RECT 1192.2001 993.3000 1193.4000 996.3000 ;
	    RECT 1194.6000 993.3000 1195.8000 999.0000 ;
	    RECT 1197.0000 993.3000 1198.2001 1001.1000 ;
	    RECT 1202.7001 1001.1000 1203.9000 1002.9000 ;
	    RECT 1202.7001 1000.2000 1205.4000 1001.1000 ;
	    RECT 1204.2001 999.3000 1205.4000 1000.2000 ;
	    RECT 1211.4000 999.6000 1212.6000 1003.8000 ;
	    RECT 1216.2001 1002.9000 1221.0000 1004.1000 ;
	    RECT 1226.7001 1002.9000 1229.7001 1004.1000 ;
	    RECT 1242.6000 1003.5000 1243.8000 1011.9000 ;
	    RECT 1264.2001 1006.5000 1265.4000 1019.7000 ;
	    RECT 1266.6000 1013.7000 1267.8000 1019.7000 ;
	    RECT 1290.6000 1013.7000 1291.8000 1019.7000 ;
	    RECT 1293.0000 1013.7000 1294.2001 1019.7000 ;
	    RECT 1295.4000 1014.3000 1296.6000 1019.7000 ;
	    RECT 1293.3000 1013.4000 1294.2001 1013.7000 ;
	    RECT 1297.8000 1013.7000 1299.0000 1019.7000 ;
	    RECT 1317.0000 1013.7000 1318.2001 1019.7000 ;
	    RECT 1297.8000 1013.4000 1298.7001 1013.7000 ;
	    RECT 1293.3000 1012.5000 1298.7001 1013.4000 ;
	    RECT 1288.2001 1011.4500 1289.4000 1011.6000 ;
	    RECT 1295.4000 1011.4500 1296.6000 1011.6000 ;
	    RECT 1288.2001 1010.5500 1296.6000 1011.4500 ;
	    RECT 1288.2001 1010.4000 1289.4000 1010.5500 ;
	    RECT 1295.4000 1010.4000 1296.6000 1010.5500 ;
	    RECT 1266.6000 1009.5000 1267.8000 1009.8000 ;
	    RECT 1297.8000 1009.5000 1298.7001 1012.5000 ;
	    RECT 1317.0000 1009.5000 1318.2001 1009.8000 ;
	    RECT 1295.4000 1009.2000 1296.6000 1009.5000 ;
	    RECT 1266.6000 1008.4500 1267.8000 1008.6000 ;
	    RECT 1288.2001 1008.4500 1289.4000 1008.6000 ;
	    RECT 1266.6000 1007.5500 1289.4000 1008.4500 ;
	    RECT 1266.6000 1007.4000 1267.8000 1007.5500 ;
	    RECT 1288.2001 1007.4000 1289.4000 1007.5500 ;
	    RECT 1290.6000 1007.4000 1291.8000 1008.6000 ;
	    RECT 1297.8000 1007.4000 1299.0000 1008.6000 ;
	    RECT 1317.0000 1007.4000 1318.2001 1008.6000 ;
	    RECT 1319.4000 1006.5000 1320.6000 1019.7000 ;
	    RECT 1321.8000 1013.7000 1323.0000 1019.7000 ;
	    RECT 1341.0000 1013.7000 1342.2001 1019.7000 ;
	    RECT 1341.0000 1009.5000 1342.2001 1009.8000 ;
	    RECT 1341.0000 1007.4000 1342.2001 1008.6000 ;
	    RECT 1343.4000 1006.5000 1344.6000 1019.7000 ;
	    RECT 1345.8000 1013.7000 1347.0000 1019.7000 ;
	    RECT 1377.0000 1007.7000 1378.2001 1019.7000 ;
	    RECT 1380.9000 1008.6000 1382.1000 1019.7000 ;
	    RECT 1383.3000 1013.7000 1384.5000 1019.7000 ;
	    RECT 1396.2001 1013.7000 1397.4000 1019.7000 ;
	    RECT 1383.0000 1010.4000 1384.2001 1011.6000 ;
	    RECT 1383.3000 1009.5000 1384.2001 1010.4000 ;
	    RECT 1380.9000 1007.7000 1382.4000 1008.6000 ;
	    RECT 1290.6000 1006.2000 1291.8000 1006.5000 ;
	    RECT 1245.0000 1005.4500 1246.2001 1005.6000 ;
	    RECT 1264.2001 1005.4500 1265.4000 1005.6000 ;
	    RECT 1245.0000 1004.5500 1265.4000 1005.4500 ;
	    RECT 1245.0000 1004.4000 1246.2001 1004.5500 ;
	    RECT 1264.2001 1004.4000 1265.4000 1004.5500 ;
	    RECT 1293.0000 1004.4000 1294.2001 1005.6000 ;
	    RECT 1295.1000 1004.4000 1295.4000 1005.6000 ;
	    RECT 1215.6000 1001.7000 1216.8000 1002.0000 ;
	    RECT 1215.6000 1000.8000 1222.2001 1001.7000 ;
	    RECT 1223.4000 1001.4000 1224.6000 1002.6000 ;
	    RECT 1221.0000 1000.5000 1222.2001 1000.8000 ;
	    RECT 1223.4000 1000.2000 1224.6000 1000.5000 ;
	    RECT 1201.8000 993.3000 1203.0000 999.3000 ;
	    RECT 1204.2001 998.1000 1207.8000 999.3000 ;
	    RECT 1211.4000 998.4000 1212.9000 999.6000 ;
	    RECT 1217.4000 998.4000 1217.7001 999.6000 ;
	    RECT 1218.6000 998.4000 1219.8000 999.6000 ;
	    RECT 1221.0000 999.3000 1222.2001 999.6000 ;
	    RECT 1226.7001 999.3000 1227.9000 1002.9000 ;
	    RECT 1230.6000 1002.3000 1243.8000 1003.5000 ;
	    RECT 1235.7001 1000.2000 1240.2001 1001.4000 ;
	    RECT 1235.7001 999.3000 1236.9000 1000.2000 ;
	    RECT 1221.0000 998.4000 1227.9000 999.3000 ;
	    RECT 1206.6000 993.3000 1207.8000 998.1000 ;
	    RECT 1233.0000 998.1000 1236.9000 999.3000 ;
	    RECT 1209.0000 993.3000 1210.2001 997.5000 ;
	    RECT 1211.4000 993.3000 1212.6000 997.5000 ;
	    RECT 1213.8000 993.3000 1215.0000 997.5000 ;
	    RECT 1216.2001 993.3000 1217.4000 997.5000 ;
	    RECT 1218.6000 993.3000 1219.8000 996.3000 ;
	    RECT 1221.0000 993.3000 1222.2001 997.5000 ;
	    RECT 1223.4000 993.3000 1224.6000 996.3000 ;
	    RECT 1225.8000 993.3000 1227.0000 997.5000 ;
	    RECT 1228.2001 993.3000 1229.4000 997.5000 ;
	    RECT 1230.6000 993.3000 1231.8000 997.5000 ;
	    RECT 1233.0000 993.3000 1234.2001 998.1000 ;
	    RECT 1237.8000 993.3000 1239.0000 999.3000 ;
	    RECT 1242.6000 993.3000 1243.8000 1002.3000 ;
	    RECT 1261.8000 1001.4000 1263.0000 1002.6000 ;
	    RECT 1261.8000 1000.2000 1263.0000 1000.5000 ;
	    RECT 1264.2001 999.3000 1265.4000 1003.5000 ;
	    RECT 1297.8000 1002.6000 1298.7001 1006.5000 ;
	    RECT 1319.4000 1005.4500 1320.6000 1005.6000 ;
	    RECT 1326.6000 1005.4500 1327.8000 1005.6000 ;
	    RECT 1319.4000 1004.5500 1327.8000 1005.4500 ;
	    RECT 1319.4000 1004.4000 1320.6000 1004.5500 ;
	    RECT 1326.6000 1004.4000 1327.8000 1004.5500 ;
	    RECT 1343.4000 1005.4500 1344.6000 1005.6000 ;
	    RECT 1357.8000 1005.4500 1359.0000 1005.6000 ;
	    RECT 1343.4000 1004.5500 1359.0000 1005.4500 ;
	    RECT 1343.4000 1004.4000 1344.6000 1004.5500 ;
	    RECT 1357.8000 1004.4000 1359.0000 1004.5500 ;
	    RECT 1379.4000 1004.4000 1380.6000 1005.6000 ;
	    RECT 1296.3000 1002.3000 1298.7001 1002.6000 ;
	    RECT 1261.8000 993.3000 1263.0000 999.3000 ;
	    RECT 1264.2001 998.4000 1266.9000 999.3000 ;
	    RECT 1265.7001 993.3000 1266.9000 998.4000 ;
	    RECT 1290.6000 993.3000 1291.8000 1002.3000 ;
	    RECT 1296.0000 1001.7000 1298.7001 1002.3000 ;
	    RECT 1296.0000 993.3000 1297.2001 1001.7000 ;
	    RECT 1319.4000 999.3000 1320.6000 1003.5000 ;
	    RECT 1321.8000 1001.4000 1323.0000 1002.6000 ;
	    RECT 1321.8000 1000.2000 1323.0000 1000.5000 ;
	    RECT 1343.4000 999.3000 1344.6000 1003.5000 ;
	    RECT 1379.4000 1003.2000 1380.6000 1003.5000 ;
	    RECT 1381.5000 1002.6000 1382.4000 1007.7000 ;
	    RECT 1384.2001 1007.4000 1385.4000 1008.6000 ;
	    RECT 1398.6000 1003.5000 1399.8000 1019.7000 ;
	    RECT 1425.0000 1007.7000 1426.2001 1019.7000 ;
	    RECT 1427.4000 1008.6000 1428.6000 1019.7000 ;
	    RECT 1429.8000 1009.5000 1431.0000 1019.7000 ;
	    RECT 1432.2001 1008.6000 1433.4000 1019.7000 ;
	    RECT 1427.4000 1007.7000 1433.4000 1008.6000 ;
	    RECT 1458.6000 1008.6000 1459.8000 1019.7000 ;
	    RECT 1461.0000 1009.5000 1462.2001 1019.7000 ;
	    RECT 1463.4000 1008.6000 1464.6000 1019.7000 ;
	    RECT 1458.6000 1007.7000 1464.6000 1008.6000 ;
	    RECT 1465.8000 1007.7000 1467.0000 1019.7000 ;
	    RECT 1489.8000 1007.7000 1491.0000 1019.7000 ;
	    RECT 1493.7001 1008.6000 1494.9000 1019.7000 ;
	    RECT 1496.1000 1013.7000 1497.3000 1019.7000 ;
	    RECT 1495.8000 1010.4000 1497.0000 1011.6000 ;
	    RECT 1496.1000 1009.5000 1497.0000 1010.4000 ;
	    RECT 1493.7001 1007.7000 1495.2001 1008.6000 ;
	    RECT 1425.3000 1006.5000 1426.2001 1007.7000 ;
	    RECT 1465.8000 1006.5000 1466.7001 1007.7000 ;
	    RECT 1425.0000 1004.4000 1426.2001 1005.6000 ;
	    RECT 1427.1000 1004.7000 1428.6000 1005.6000 ;
	    RECT 1431.0000 1004.7000 1431.3000 1006.2000 ;
	    RECT 1345.8000 1002.4500 1347.0000 1002.6000 ;
	    RECT 1350.6000 1002.4500 1351.8000 1002.6000 ;
	    RECT 1345.8000 1001.5500 1351.8000 1002.4500 ;
	    RECT 1345.8000 1001.4000 1347.0000 1001.5500 ;
	    RECT 1350.6000 1001.4000 1351.8000 1001.5500 ;
	    RECT 1353.0000 1002.4500 1354.2001 1002.6000 ;
	    RECT 1377.0000 1002.4500 1378.2001 1002.6000 ;
	    RECT 1353.0000 1001.5500 1378.2001 1002.4500 ;
	    RECT 1353.0000 1001.4000 1354.2001 1001.5500 ;
	    RECT 1377.0000 1001.4000 1378.2001 1001.5500 ;
	    RECT 1379.1000 1000.8000 1379.4000 1002.3000 ;
	    RECT 1381.5000 1001.4000 1383.3000 1002.6000 ;
	    RECT 1384.2001 1002.4500 1385.4000 1002.6000 ;
	    RECT 1396.2001 1002.4500 1397.4000 1002.6000 ;
	    RECT 1384.2001 1001.5500 1397.4000 1002.4500 ;
	    RECT 1384.2001 1001.4000 1385.4000 1001.5500 ;
	    RECT 1396.2001 1001.4000 1397.4000 1001.5500 ;
	    RECT 1398.6000 1002.4500 1399.8000 1002.6000 ;
	    RECT 1398.6000 1001.5500 1426.0500 1002.4500 ;
	    RECT 1398.6000 1001.4000 1399.8000 1001.5500 ;
	    RECT 1345.8000 1000.2000 1347.0000 1000.5000 ;
	    RECT 1377.3000 999.3000 1382.7001 999.9000 ;
	    RECT 1384.2001 999.3000 1385.1000 1000.5000 ;
	    RECT 1386.6000 999.4500 1387.8000 999.6000 ;
	    RECT 1396.2001 999.4500 1397.4000 999.6000 ;
	    RECT 1317.9000 998.4000 1320.6000 999.3000 ;
	    RECT 1317.9000 993.3000 1319.1000 998.4000 ;
	    RECT 1321.8000 993.3000 1323.0000 999.3000 ;
	    RECT 1341.9000 998.4000 1344.6000 999.3000 ;
	    RECT 1341.9000 993.3000 1343.1000 998.4000 ;
	    RECT 1345.8000 993.3000 1347.0000 999.3000 ;
	    RECT 1377.0000 999.0000 1383.0000 999.3000 ;
	    RECT 1377.0000 993.3000 1378.2001 999.0000 ;
	    RECT 1379.4000 993.3000 1380.6000 998.1000 ;
	    RECT 1381.8000 993.3000 1383.0000 999.0000 ;
	    RECT 1384.2001 993.3000 1385.4000 999.3000 ;
	    RECT 1386.6000 998.5500 1397.4000 999.4500 ;
	    RECT 1386.6000 998.4000 1387.8000 998.5500 ;
	    RECT 1396.2001 998.4000 1397.4000 998.5500 ;
	    RECT 1396.2001 997.2000 1397.4000 997.5000 ;
	    RECT 1396.2001 993.3000 1397.4000 996.3000 ;
	    RECT 1398.6000 993.3000 1399.8000 1000.5000 ;
	    RECT 1425.1500 999.6000 1426.0500 1001.5500 ;
	    RECT 1425.0000 998.4000 1426.2001 999.6000 ;
	    RECT 1427.7001 999.3000 1428.6000 1004.7000 ;
	    RECT 1432.2001 1004.4000 1433.4000 1005.6000 ;
	    RECT 1453.8000 1005.4500 1455.0000 1005.6000 ;
	    RECT 1458.6000 1005.4500 1459.8000 1005.6000 ;
	    RECT 1453.8000 1004.5500 1459.8000 1005.4500 ;
	    RECT 1460.7001 1004.7000 1461.0000 1006.2000 ;
	    RECT 1463.4000 1004.7000 1464.9000 1005.6000 ;
	    RECT 1465.8000 1005.4500 1467.0000 1005.6000 ;
	    RECT 1489.8000 1005.4500 1491.0000 1005.6000 ;
	    RECT 1453.8000 1004.4000 1455.0000 1004.5500 ;
	    RECT 1458.6000 1004.4000 1459.8000 1004.5500 ;
	    RECT 1429.8000 1003.5000 1431.0000 1003.8000 ;
	    RECT 1461.0000 1003.5000 1462.2001 1003.8000 ;
	    RECT 1429.8000 1001.4000 1431.0000 1002.6000 ;
	    RECT 1444.2001 1002.4500 1445.4000 1002.6000 ;
	    RECT 1461.0000 1002.4500 1462.2001 1002.6000 ;
	    RECT 1444.2001 1001.5500 1462.2001 1002.4500 ;
	    RECT 1444.2001 1001.4000 1445.4000 1001.5500 ;
	    RECT 1461.0000 1001.4000 1462.2001 1001.5500 ;
	    RECT 1463.4000 999.3000 1464.3000 1004.7000 ;
	    RECT 1465.8000 1004.5500 1491.0000 1005.4500 ;
	    RECT 1465.8000 1004.4000 1467.0000 1004.5500 ;
	    RECT 1489.8000 1004.4000 1491.0000 1004.5500 ;
	    RECT 1492.2001 1004.4000 1493.4000 1005.6000 ;
	    RECT 1489.9501 1002.6000 1490.8500 1004.4000 ;
	    RECT 1492.2001 1003.2000 1493.4000 1003.5000 ;
	    RECT 1494.3000 1002.6000 1495.2001 1007.7000 ;
	    RECT 1497.0000 1007.4000 1498.2001 1008.6000 ;
	    RECT 1509.0000 1003.5000 1510.2001 1019.7000 ;
	    RECT 1511.4000 1013.7000 1512.6000 1019.7000 ;
	    RECT 1513.8000 1019.4000 1515.0000 1020.6000 ;
	    RECT 1516.2001 1014.4500 1517.4000 1014.6000 ;
	    RECT 1535.4000 1014.4500 1536.6000 1014.6000 ;
	    RECT 1516.2001 1013.5500 1536.6000 1014.4500 ;
	    RECT 1537.8000 1013.7000 1539.0000 1019.7000 ;
	    RECT 1540.2001 1013.7000 1541.4000 1019.7000 ;
	    RECT 1542.6000 1014.3000 1543.8000 1019.7000 ;
	    RECT 1516.2001 1013.4000 1517.4000 1013.5500 ;
	    RECT 1535.4000 1013.4000 1536.6000 1013.5500 ;
	    RECT 1540.5000 1013.4000 1541.4000 1013.7000 ;
	    RECT 1545.0000 1013.7000 1546.2001 1019.7000 ;
	    RECT 1545.0000 1013.4000 1545.9000 1013.7000 ;
	    RECT 1540.5000 1012.5000 1545.9000 1013.4000 ;
	    RECT 1521.0000 1011.4500 1522.2001 1011.6000 ;
	    RECT 1542.6000 1011.4500 1543.8000 1011.6000 ;
	    RECT 1521.0000 1010.5500 1543.8000 1011.4500 ;
	    RECT 1521.0000 1010.4000 1522.2001 1010.5500 ;
	    RECT 1542.6000 1010.4000 1543.8000 1010.5500 ;
	    RECT 1545.0000 1009.5000 1545.9000 1012.5000 ;
	    RECT 1542.6000 1009.2000 1543.8000 1009.5000 ;
	    RECT 1533.0000 1008.4500 1534.2001 1008.6000 ;
	    RECT 1537.8000 1008.4500 1539.0000 1008.6000 ;
	    RECT 1540.2001 1008.4500 1541.4000 1008.6000 ;
	    RECT 1533.0000 1007.5500 1541.4000 1008.4500 ;
	    RECT 1533.0000 1007.4000 1534.2001 1007.5500 ;
	    RECT 1537.8000 1007.4000 1539.0000 1007.5500 ;
	    RECT 1540.2001 1007.4000 1541.4000 1007.5500 ;
	    RECT 1545.0000 1008.4500 1546.2001 1008.6000 ;
	    RECT 1547.4000 1008.4500 1548.6000 1008.6000 ;
	    RECT 1545.0000 1007.5500 1548.6000 1008.4500 ;
	    RECT 1545.0000 1007.4000 1546.2001 1007.5500 ;
	    RECT 1547.4000 1007.4000 1548.6000 1007.5500 ;
	    RECT 1537.8000 1006.2000 1539.0000 1006.5000 ;
	    RECT 1540.2001 1004.4000 1541.4000 1005.6000 ;
	    RECT 1542.3000 1004.4000 1542.6000 1005.6000 ;
	    RECT 1545.0000 1002.6000 1545.9000 1006.5000 ;
	    RECT 1489.8000 1001.4000 1491.0000 1002.6000 ;
	    RECT 1491.9000 1000.8000 1492.2001 1002.3000 ;
	    RECT 1494.3000 1001.4000 1496.1000 1002.6000 ;
	    RECT 1497.0000 1001.4000 1498.2001 1002.6000 ;
	    RECT 1499.4000 1002.4500 1500.6000 1002.6000 ;
	    RECT 1509.0000 1002.4500 1510.2001 1002.6000 ;
	    RECT 1523.4000 1002.4500 1524.6000 1002.6000 ;
	    RECT 1499.4000 1001.5500 1524.6000 1002.4500 ;
	    RECT 1543.5000 1002.3000 1545.9000 1002.6000 ;
	    RECT 1499.4000 1001.4000 1500.6000 1001.5500 ;
	    RECT 1509.0000 1001.4000 1510.2001 1001.5500 ;
	    RECT 1523.4000 1001.4000 1524.6000 1001.5500 ;
	    RECT 1425.3000 997.2000 1426.5000 997.5000 ;
	    RECT 1425.0000 993.3000 1426.2001 996.3000 ;
	    RECT 1427.4000 993.3000 1428.6000 999.3000 ;
	    RECT 1431.3000 993.3000 1432.5000 999.3000 ;
	    RECT 1459.5000 993.3000 1460.7001 999.3000 ;
	    RECT 1463.4000 993.3000 1464.6000 999.3000 ;
	    RECT 1465.8000 998.4000 1467.0000 999.6000 ;
	    RECT 1490.1000 999.3000 1495.5000 999.9000 ;
	    RECT 1497.0000 999.3000 1497.9000 1000.5000 ;
	    RECT 1489.8000 999.0000 1495.8000 999.3000 ;
	    RECT 1465.5000 997.2000 1466.7001 997.5000 ;
	    RECT 1465.8000 993.3000 1467.0000 996.3000 ;
	    RECT 1489.8000 993.3000 1491.0000 999.0000 ;
	    RECT 1492.2001 993.3000 1493.4000 998.1000 ;
	    RECT 1494.6000 993.3000 1495.8000 999.0000 ;
	    RECT 1497.0000 993.3000 1498.2001 999.3000 ;
	    RECT 1509.0000 993.3000 1510.2001 1000.5000 ;
	    RECT 1511.4000 999.4500 1512.6000 999.6000 ;
	    RECT 1533.0000 999.4500 1534.2001 999.6000 ;
	    RECT 1511.4000 998.5500 1534.2001 999.4500 ;
	    RECT 1511.4000 998.4000 1512.6000 998.5500 ;
	    RECT 1533.0000 998.4000 1534.2001 998.5500 ;
	    RECT 1511.4000 997.2000 1512.6000 997.5000 ;
	    RECT 1511.4000 993.3000 1512.6000 996.3000 ;
	    RECT 1537.8000 993.3000 1539.0000 1002.3000 ;
	    RECT 1543.2001 1001.7000 1545.9000 1002.3000 ;
	    RECT 1543.2001 993.3000 1544.4000 1001.7000 ;
	    RECT 1.2000 990.6000 1569.0000 992.4000 ;
	    RECT 126.6000 980.7000 127.8000 989.7000 ;
	    RECT 131.4000 983.7000 132.6000 989.7000 ;
	    RECT 136.2000 984.9000 137.4000 989.7000 ;
	    RECT 138.6000 985.5000 139.8000 989.7000 ;
	    RECT 141.0000 985.5000 142.2000 989.7000 ;
	    RECT 143.4000 985.5000 144.6000 989.7000 ;
	    RECT 145.8000 986.7000 147.0000 989.7000 ;
	    RECT 148.2000 985.5000 149.4000 989.7000 ;
	    RECT 150.6000 986.7000 151.8000 989.7000 ;
	    RECT 153.0000 985.5000 154.2000 989.7000 ;
	    RECT 155.4000 985.5000 156.6000 989.7000 ;
	    RECT 157.8000 985.5000 159.0000 989.7000 ;
	    RECT 160.2000 985.5000 161.4000 989.7000 ;
	    RECT 133.5000 983.7000 137.4000 984.9000 ;
	    RECT 162.6000 984.9000 163.8000 989.7000 ;
	    RECT 142.5000 983.7000 149.4000 984.6000 ;
	    RECT 133.5000 982.8000 134.7000 983.7000 ;
	    RECT 130.2000 981.6000 134.7000 982.8000 ;
	    RECT 126.6000 979.5000 139.8000 980.7000 ;
	    RECT 142.5000 980.1000 143.7000 983.7000 ;
	    RECT 148.2000 983.4000 149.4000 983.7000 ;
	    RECT 150.6000 983.4000 151.8000 984.6000 ;
	    RECT 152.7000 983.4000 153.0000 984.6000 ;
	    RECT 157.5000 983.4000 159.0000 984.6000 ;
	    RECT 162.6000 983.7000 166.2000 984.9000 ;
	    RECT 167.4000 983.7000 168.6000 989.7000 ;
	    RECT 145.8000 982.5000 147.0000 982.8000 ;
	    RECT 148.2000 982.2000 149.4000 982.5000 ;
	    RECT 145.8000 980.4000 147.0000 981.6000 ;
	    RECT 148.2000 981.3000 154.8000 982.2000 ;
	    RECT 153.6000 981.0000 154.8000 981.3000 ;
	    RECT 126.6000 971.1000 127.8000 979.5000 ;
	    RECT 140.7000 978.9000 143.7000 980.1000 ;
	    RECT 149.4000 978.9000 154.2000 980.1000 ;
	    RECT 157.8000 979.2000 159.0000 983.4000 ;
	    RECT 165.0000 982.8000 166.2000 983.7000 ;
	    RECT 165.0000 981.9000 167.7000 982.8000 ;
	    RECT 166.5000 980.1000 167.7000 981.9000 ;
	    RECT 172.2000 981.9000 173.4000 989.7000 ;
	    RECT 174.6000 984.0000 175.8000 989.7000 ;
	    RECT 177.0000 986.7000 178.2000 989.7000 ;
	    RECT 215.4000 984.0000 216.6000 989.7000 ;
	    RECT 217.8000 984.9000 219.0000 989.7000 ;
	    RECT 220.2000 988.8000 226.2000 989.7000 ;
	    RECT 220.2000 984.0000 221.4000 988.8000 ;
	    RECT 174.6000 982.8000 176.1000 984.0000 ;
	    RECT 215.4000 983.7000 221.4000 984.0000 ;
	    RECT 222.6000 983.7000 223.8000 987.9000 ;
	    RECT 225.0000 983.7000 226.2000 988.8000 ;
	    RECT 244.2000 986.7000 245.4000 989.7000 ;
	    RECT 246.6000 986.7000 247.8000 989.7000 ;
	    RECT 249.0000 986.7000 250.2000 989.7000 ;
	    RECT 244.2000 985.5000 245.4000 985.8000 ;
	    RECT 237.0000 984.4500 238.2000 984.6000 ;
	    RECT 244.2000 984.4500 245.4000 984.6000 ;
	    RECT 215.7000 983.1000 221.1000 983.7000 ;
	    RECT 172.2000 981.0000 174.0000 981.9000 ;
	    RECT 166.5000 978.9000 172.2000 980.1000 ;
	    RECT 128.7000 978.0000 129.9000 978.3000 ;
	    RECT 128.7000 977.1000 135.3000 978.0000 ;
	    RECT 136.2000 977.4000 137.4000 978.6000 ;
	    RECT 162.6000 978.0000 163.8000 978.9000 ;
	    RECT 173.1000 978.0000 174.0000 981.0000 ;
	    RECT 138.3000 977.1000 163.8000 978.0000 ;
	    RECT 172.8000 977.1000 174.0000 978.0000 ;
	    RECT 170.7000 976.2000 171.9000 976.5000 ;
	    RECT 131.4000 974.4000 132.6000 975.6000 ;
	    RECT 133.5000 975.3000 171.9000 976.2000 ;
	    RECT 136.5000 975.0000 137.7000 975.3000 ;
	    RECT 172.8000 974.4000 173.7000 977.1000 ;
	    RECT 174.9000 976.2000 176.1000 982.8000 ;
	    RECT 210.6000 981.4500 211.8000 981.6000 ;
	    RECT 215.4000 981.4500 216.6000 981.6000 ;
	    RECT 210.6000 980.5500 216.6000 981.4500 ;
	    RECT 217.5000 980.7000 217.8000 982.2000 ;
	    RECT 222.9000 981.6000 223.8000 983.7000 ;
	    RECT 237.0000 983.5500 245.4000 984.4500 ;
	    RECT 237.0000 983.4000 238.2000 983.5500 ;
	    RECT 244.2000 983.4000 245.4000 983.5500 ;
	    RECT 246.9000 982.5000 247.8000 986.7000 ;
	    RECT 268.2000 983.7000 269.4000 989.7000 ;
	    RECT 272.1000 984.6000 273.3000 989.7000 ;
	    RECT 270.6000 983.7000 273.3000 984.6000 ;
	    RECT 268.2000 982.5000 269.4000 982.8000 ;
	    RECT 210.6000 980.4000 211.8000 980.5500 ;
	    RECT 215.4000 980.4000 216.6000 980.5500 ;
	    RECT 220.2000 980.4000 221.4000 981.6000 ;
	    RECT 222.3000 980.7000 223.8000 981.6000 ;
	    RECT 225.0000 981.4500 226.2000 981.6000 ;
	    RECT 227.4000 981.4500 228.6000 981.6000 ;
	    RECT 225.0000 980.5500 228.6000 981.4500 ;
	    RECT 225.0000 980.4000 226.2000 980.5500 ;
	    RECT 227.4000 980.4000 228.6000 980.5500 ;
	    RECT 246.6000 981.4500 247.8000 981.6000 ;
	    RECT 265.8000 981.4500 267.0000 981.6000 ;
	    RECT 246.6000 980.5500 267.0000 981.4500 ;
	    RECT 246.6000 980.4000 247.8000 980.5500 ;
	    RECT 265.8000 980.4000 267.0000 980.5500 ;
	    RECT 268.2000 980.4000 269.4000 981.6000 ;
	    RECT 217.8000 979.5000 219.0000 979.8000 ;
	    RECT 222.6000 979.5000 223.8000 979.8000 ;
	    RECT 270.6000 979.5000 271.8000 983.7000 ;
	    RECT 298.8000 981.3000 300.0000 989.7000 ;
	    RECT 297.3000 980.7000 300.0000 981.3000 ;
	    RECT 304.2000 980.7000 305.4000 989.7000 ;
	    RECT 373.8000 983.1000 375.0000 989.7000 ;
	    RECT 376.2000 984.0000 377.4000 989.7000 ;
	    RECT 380.1000 987.6000 381.9000 989.7000 ;
	    RECT 380.1000 986.7000 382.2000 987.6000 ;
	    RECT 384.6000 986.7000 385.8000 989.7000 ;
	    RECT 387.0000 986.7000 388.2000 989.7000 ;
	    RECT 389.4000 986.7000 390.9000 989.7000 ;
	    RECT 393.6000 987.6000 394.8000 989.7000 ;
	    RECT 393.6000 986.7000 396.6000 987.6000 ;
	    RECT 381.0000 985.5000 382.2000 986.7000 ;
	    RECT 387.3000 985.8000 388.2000 986.7000 ;
	    RECT 387.3000 984.9000 391.5000 985.8000 ;
	    RECT 390.3000 984.6000 391.5000 984.9000 ;
	    RECT 393.0000 984.6000 394.2000 985.8000 ;
	    RECT 395.4000 985.5000 396.6000 986.7000 ;
	    RECT 378.3000 983.1000 379.5000 983.4000 ;
	    RECT 373.8000 982.2000 379.5000 983.1000 ;
	    RECT 297.3000 980.4000 299.7000 980.7000 ;
	    RECT 191.4000 978.4500 192.6000 978.6000 ;
	    RECT 217.8000 978.4500 219.0000 978.6000 ;
	    RECT 191.4000 977.5500 219.0000 978.4500 ;
	    RECT 191.4000 977.4000 192.6000 977.5500 ;
	    RECT 217.8000 977.4000 219.0000 977.5500 ;
	    RECT 141.0000 974.1000 142.2000 974.4000 ;
	    RECT 134.1000 973.5000 142.2000 974.1000 ;
	    RECT 132.9000 973.2000 142.2000 973.5000 ;
	    RECT 143.7000 973.5000 156.6000 974.4000 ;
	    RECT 129.0000 972.0000 131.4000 973.2000 ;
	    RECT 132.9000 972.3000 135.0000 973.2000 ;
	    RECT 143.7000 972.3000 144.6000 973.5000 ;
	    RECT 155.4000 973.2000 156.6000 973.5000 ;
	    RECT 160.2000 973.5000 173.7000 974.4000 ;
	    RECT 174.6000 975.0000 176.1000 976.2000 ;
	    RECT 220.2000 975.3000 221.1000 979.5000 ;
	    RECT 225.0000 979.2000 226.2000 979.5000 ;
	    RECT 222.6000 977.4000 223.8000 978.6000 ;
	    RECT 246.9000 975.3000 247.8000 979.5000 ;
	    RECT 249.0000 977.4000 250.2000 978.6000 ;
	    RECT 270.6000 977.4000 271.8000 978.6000 ;
	    RECT 297.3000 976.5000 298.2000 980.4000 ;
	    RECT 373.8000 979.5000 375.0000 982.2000 ;
	    RECT 384.3000 981.3000 385.5000 981.6000 ;
	    RECT 393.0000 981.3000 393.9000 984.6000 ;
	    RECT 397.8000 983.7000 399.0000 989.7000 ;
	    RECT 400.2000 982.5000 401.4000 989.7000 ;
	    RECT 419.4000 983.7000 420.6000 989.7000 ;
	    RECT 423.3000 984.6000 424.5000 989.7000 ;
	    RECT 465.0000 987.4500 466.2000 987.6000 ;
	    RECT 486.6000 987.4500 487.8000 987.6000 ;
	    RECT 465.0000 986.5500 487.8000 987.4500 ;
	    RECT 465.0000 986.4000 466.2000 986.5500 ;
	    RECT 486.6000 986.4000 487.8000 986.5500 ;
	    RECT 421.8000 983.7000 424.5000 984.6000 ;
	    RECT 419.4000 982.5000 420.6000 982.8000 ;
	    RECT 383.7000 980.4000 396.9000 981.3000 ;
	    RECT 397.8000 980.4000 399.0000 981.6000 ;
	    RECT 399.9000 980.4000 400.2000 981.6000 ;
	    RECT 419.4000 980.4000 420.6000 981.6000 ;
	    RECT 381.0000 979.2000 382.2000 979.5000 ;
	    RECT 300.6000 977.4000 300.9000 978.6000 ;
	    RECT 301.8000 977.4000 303.0000 978.6000 ;
	    RECT 313.8000 978.4500 315.0000 978.6000 ;
	    RECT 373.8000 978.4500 375.0000 978.6000 ;
	    RECT 313.8000 977.5500 375.0000 978.4500 ;
	    RECT 376.5000 978.3000 382.2000 979.2000 ;
	    RECT 376.5000 978.0000 377.7000 978.3000 ;
	    RECT 313.8000 977.4000 315.0000 977.5500 ;
	    RECT 373.8000 977.4000 375.0000 977.5500 ;
	    RECT 378.9000 977.1000 380.1000 977.4000 ;
	    RECT 304.2000 976.5000 305.4000 976.8000 ;
	    RECT 375.9000 976.5000 380.1000 977.1000 ;
	    RECT 249.0000 976.2000 250.2000 976.5000 ;
	    RECT 174.6000 973.5000 175.8000 975.0000 ;
	    RECT 160.2000 973.2000 161.4000 973.5000 ;
	    RECT 130.5000 971.4000 131.4000 972.0000 ;
	    RECT 135.9000 971.4000 144.6000 972.3000 ;
	    RECT 145.5000 971.4000 149.4000 972.6000 ;
	    RECT 126.6000 970.2000 129.6000 971.1000 ;
	    RECT 130.5000 970.2000 136.8000 971.4000 ;
	    RECT 128.7000 969.3000 129.6000 970.2000 ;
	    RECT 126.6000 963.3000 127.8000 969.3000 ;
	    RECT 128.7000 968.4000 130.2000 969.3000 ;
	    RECT 129.0000 963.3000 130.2000 968.4000 ;
	    RECT 131.4000 962.4000 132.6000 969.3000 ;
	    RECT 133.8000 963.3000 135.0000 970.2000 ;
	    RECT 136.2000 963.3000 137.4000 969.3000 ;
	    RECT 138.6000 963.3000 139.8000 967.5000 ;
	    RECT 141.0000 963.3000 142.2000 967.5000 ;
	    RECT 143.4000 963.3000 144.6000 970.5000 ;
	    RECT 145.8000 963.3000 147.0000 969.3000 ;
	    RECT 148.2000 963.3000 149.4000 970.5000 ;
	    RECT 150.6000 963.3000 151.8000 969.3000 ;
	    RECT 153.0000 963.3000 154.2000 972.6000 ;
	    RECT 165.0000 971.4000 168.9000 972.6000 ;
	    RECT 157.8000 970.2000 164.1000 971.4000 ;
	    RECT 155.4000 963.3000 156.6000 967.5000 ;
	    RECT 157.8000 963.3000 159.0000 967.5000 ;
	    RECT 160.2000 963.3000 161.4000 967.5000 ;
	    RECT 162.6000 963.3000 163.8000 969.3000 ;
	    RECT 165.0000 963.3000 166.2000 971.4000 ;
	    RECT 172.8000 971.1000 173.7000 973.5000 ;
	    RECT 174.6000 971.4000 175.8000 972.6000 ;
	    RECT 169.8000 970.2000 173.7000 971.1000 ;
	    RECT 167.4000 963.3000 168.6000 969.3000 ;
	    RECT 169.8000 963.3000 171.0000 970.2000 ;
	    RECT 172.2000 963.3000 173.4000 969.3000 ;
	    RECT 174.6000 963.3000 175.8000 970.5000 ;
	    RECT 177.0000 963.3000 178.2000 969.3000 ;
	    RECT 215.4000 963.3000 216.6000 975.3000 ;
	    RECT 219.3000 963.3000 222.3000 975.3000 ;
	    RECT 225.0000 963.3000 226.2000 975.3000 ;
	    RECT 244.2000 963.3000 245.4000 975.3000 ;
	    RECT 246.6000 974.1000 249.3000 975.3000 ;
	    RECT 248.1000 963.3000 249.3000 974.1000 ;
	    RECT 268.2000 963.3000 269.4000 969.3000 ;
	    RECT 270.6000 963.3000 271.8000 976.5000 ;
	    RECT 373.8000 976.2000 380.1000 976.5000 ;
	    RECT 273.0000 974.4000 274.2000 975.6000 ;
	    RECT 275.4000 975.4500 276.6000 975.6000 ;
	    RECT 297.0000 975.4500 298.2000 975.6000 ;
	    RECT 275.4000 974.5500 298.2000 975.4500 ;
	    RECT 275.4000 974.4000 276.6000 974.5500 ;
	    RECT 297.0000 974.4000 298.2000 974.5500 ;
	    RECT 304.2000 974.4000 305.4000 975.6000 ;
	    RECT 299.4000 973.5000 300.6000 973.8000 ;
	    RECT 273.0000 973.2000 274.2000 973.5000 ;
	    RECT 297.3000 970.5000 298.2000 973.5000 ;
	    RECT 299.4000 972.4500 300.6000 972.6000 ;
	    RECT 313.8000 972.4500 315.0000 972.6000 ;
	    RECT 299.4000 971.5500 315.0000 972.4500 ;
	    RECT 299.4000 971.4000 300.6000 971.5500 ;
	    RECT 313.8000 971.4000 315.0000 971.5500 ;
	    RECT 297.3000 969.6000 302.7000 970.5000 ;
	    RECT 297.3000 969.3000 298.2000 969.6000 ;
	    RECT 273.0000 963.3000 274.2000 969.3000 ;
	    RECT 297.0000 963.3000 298.2000 969.3000 ;
	    RECT 301.8000 969.3000 302.7000 969.6000 ;
	    RECT 299.4000 963.3000 300.6000 968.7000 ;
	    RECT 301.8000 963.3000 303.0000 969.3000 ;
	    RECT 304.2000 963.3000 305.4000 969.3000 ;
	    RECT 309.0000 966.4500 310.2000 966.6000 ;
	    RECT 337.8000 966.4500 339.0000 966.6000 ;
	    RECT 309.0000 965.5500 339.0000 966.4500 ;
	    RECT 309.0000 965.4000 310.2000 965.5500 ;
	    RECT 337.8000 965.4000 339.0000 965.5500 ;
	    RECT 373.8000 963.3000 375.0000 976.2000 ;
	    RECT 383.7000 975.6000 384.6000 980.4000 ;
	    RECT 394.5000 980.1000 395.7000 980.4000 ;
	    RECT 421.8000 979.5000 423.0000 983.7000 ;
	    RECT 501.0000 983.1000 502.2000 989.7000 ;
	    RECT 503.4000 984.0000 504.6000 989.7000 ;
	    RECT 507.3000 987.6000 509.1000 989.7000 ;
	    RECT 507.3000 986.7000 509.4000 987.6000 ;
	    RECT 511.8000 986.7000 513.0000 989.7000 ;
	    RECT 514.2000 986.7000 515.4000 989.7000 ;
	    RECT 516.6000 986.7000 518.1000 989.7000 ;
	    RECT 520.8000 987.6000 522.0000 989.7000 ;
	    RECT 520.8000 986.7000 523.8000 987.6000 ;
	    RECT 508.2000 985.5000 509.4000 986.7000 ;
	    RECT 514.5000 985.8000 515.4000 986.7000 ;
	    RECT 514.5000 984.9000 518.7000 985.8000 ;
	    RECT 517.5000 984.6000 518.7000 984.9000 ;
	    RECT 520.2000 984.6000 521.4000 985.8000 ;
	    RECT 522.6000 985.5000 523.8000 986.7000 ;
	    RECT 505.5000 983.1000 506.7000 983.4000 ;
	    RECT 501.0000 982.2000 506.7000 983.1000 ;
	    RECT 501.0000 979.5000 502.2000 982.2000 ;
	    RECT 511.5000 981.3000 512.7000 981.6000 ;
	    RECT 520.2000 981.3000 521.1000 984.6000 ;
	    RECT 525.0000 983.7000 526.2000 989.7000 ;
	    RECT 527.4000 982.5000 528.6000 989.7000 ;
	    RECT 613.8000 987.4500 615.0000 987.6000 ;
	    RECT 633.0000 987.4500 634.2000 987.6000 ;
	    RECT 613.8000 986.5500 634.2000 987.4500 ;
	    RECT 613.8000 986.4000 615.0000 986.5500 ;
	    RECT 633.0000 986.4000 634.2000 986.5500 ;
	    RECT 623.4000 984.4500 624.6000 984.6000 ;
	    RECT 637.8000 984.4500 639.0000 984.6000 ;
	    RECT 623.4000 983.5500 639.0000 984.4500 ;
	    RECT 623.4000 983.4000 624.6000 983.5500 ;
	    RECT 637.8000 983.4000 639.0000 983.5500 ;
	    RECT 510.9000 980.4000 524.1000 981.3000 ;
	    RECT 525.0000 980.4000 526.2000 981.6000 ;
	    RECT 527.1000 980.4000 527.4000 981.6000 ;
	    RECT 659.4000 980.7000 660.6000 989.7000 ;
	    RECT 664.2000 983.7000 665.4000 989.7000 ;
	    RECT 669.0000 984.9000 670.2000 989.7000 ;
	    RECT 671.4000 985.5000 672.6000 989.7000 ;
	    RECT 673.8000 985.5000 675.0000 989.7000 ;
	    RECT 676.2000 985.5000 677.4000 989.7000 ;
	    RECT 678.6000 986.7000 679.8000 989.7000 ;
	    RECT 681.0000 985.5000 682.2000 989.7000 ;
	    RECT 683.4000 986.7000 684.6000 989.7000 ;
	    RECT 685.8000 985.5000 687.0000 989.7000 ;
	    RECT 688.2000 985.5000 689.4000 989.7000 ;
	    RECT 690.6000 985.5000 691.8000 989.7000 ;
	    RECT 693.0000 985.5000 694.2000 989.7000 ;
	    RECT 666.3000 983.7000 670.2000 984.9000 ;
	    RECT 695.4000 984.9000 696.6000 989.7000 ;
	    RECT 675.3000 983.7000 682.2000 984.6000 ;
	    RECT 666.3000 982.8000 667.5000 983.7000 ;
	    RECT 663.0000 981.6000 667.5000 982.8000 ;
	    RECT 508.2000 979.2000 509.4000 979.5000 ;
	    RECT 396.9000 978.6000 398.1000 978.9000 ;
	    RECT 390.6000 977.4000 391.8000 978.6000 ;
	    RECT 392.7000 977.7000 398.1000 978.6000 ;
	    RECT 421.8000 978.4500 423.0000 978.6000 ;
	    RECT 453.0000 978.4500 454.2000 978.6000 ;
	    RECT 421.8000 977.5500 454.2000 978.4500 ;
	    RECT 421.8000 977.4000 423.0000 977.5500 ;
	    RECT 453.0000 977.4000 454.2000 977.5500 ;
	    RECT 455.4000 978.4500 456.6000 978.6000 ;
	    RECT 501.0000 978.4500 502.2000 978.6000 ;
	    RECT 455.4000 977.5500 502.2000 978.4500 ;
	    RECT 503.7000 978.3000 509.4000 979.2000 ;
	    RECT 503.7000 978.0000 504.9000 978.3000 ;
	    RECT 455.4000 977.4000 456.6000 977.5500 ;
	    RECT 501.0000 977.4000 502.2000 977.5500 ;
	    RECT 506.1000 977.1000 507.3000 977.4000 ;
	    RECT 393.0000 976.5000 401.4000 976.8000 ;
	    RECT 503.1000 976.5000 507.3000 977.1000 ;
	    RECT 392.7000 976.2000 401.4000 976.5000 ;
	    RECT 376.2000 963.3000 377.4000 975.3000 ;
	    RECT 381.0000 974.7000 384.6000 975.6000 ;
	    RECT 386.7000 975.9000 401.4000 976.2000 ;
	    RECT 386.7000 975.3000 393.9000 975.9000 ;
	    RECT 381.0000 973.2000 381.9000 974.7000 ;
	    RECT 379.8000 972.0000 381.9000 973.2000 ;
	    RECT 384.3000 973.5000 385.5000 973.8000 ;
	    RECT 386.7000 973.5000 387.6000 975.3000 ;
	    RECT 384.3000 972.6000 387.6000 973.5000 ;
	    RECT 388.5000 973.5000 396.6000 974.4000 ;
	    RECT 388.5000 973.2000 389.7000 973.5000 ;
	    RECT 395.4000 973.2000 396.6000 973.5000 ;
	    RECT 386.1000 971.1000 387.3000 971.4000 ;
	    RECT 390.3000 971.1000 391.5000 971.4000 ;
	    RECT 381.0000 969.3000 382.2000 970.5000 ;
	    RECT 386.1000 970.2000 391.5000 971.1000 ;
	    RECT 387.3000 969.3000 388.2000 970.2000 ;
	    RECT 395.4000 969.3000 396.6000 970.5000 ;
	    RECT 380.1000 963.3000 381.9000 969.3000 ;
	    RECT 384.6000 963.3000 385.8000 969.3000 ;
	    RECT 387.0000 963.3000 388.2000 969.3000 ;
	    RECT 389.4000 963.3000 390.6000 969.3000 ;
	    RECT 393.6000 968.4000 396.6000 969.3000 ;
	    RECT 393.6000 963.3000 394.8000 968.4000 ;
	    RECT 397.8000 963.3000 399.0000 975.0000 ;
	    RECT 400.2000 963.3000 401.4000 975.9000 ;
	    RECT 419.4000 963.3000 420.6000 969.3000 ;
	    RECT 421.8000 963.3000 423.0000 976.5000 ;
	    RECT 501.0000 976.2000 507.3000 976.5000 ;
	    RECT 424.2000 975.4500 425.4000 975.6000 ;
	    RECT 460.2000 975.4500 461.4000 975.6000 ;
	    RECT 424.2000 974.5500 461.4000 975.4500 ;
	    RECT 424.2000 974.4000 425.4000 974.5500 ;
	    RECT 460.2000 974.4000 461.4000 974.5500 ;
	    RECT 424.2000 973.2000 425.4000 973.5000 ;
	    RECT 424.2000 963.3000 425.4000 969.3000 ;
	    RECT 501.0000 963.3000 502.2000 976.2000 ;
	    RECT 510.9000 975.6000 511.8000 980.4000 ;
	    RECT 521.7000 980.1000 522.9000 980.4000 ;
	    RECT 659.4000 979.5000 672.6000 980.7000 ;
	    RECT 675.3000 980.1000 676.5000 983.7000 ;
	    RECT 681.0000 983.4000 682.2000 983.7000 ;
	    RECT 683.4000 983.4000 684.6000 984.6000 ;
	    RECT 685.5000 983.4000 685.8000 984.6000 ;
	    RECT 690.3000 983.4000 691.8000 984.6000 ;
	    RECT 695.4000 983.7000 699.0000 984.9000 ;
	    RECT 700.2000 983.7000 701.4000 989.7000 ;
	    RECT 678.6000 982.5000 679.8000 982.8000 ;
	    RECT 681.0000 982.2000 682.2000 982.5000 ;
	    RECT 678.6000 980.4000 679.8000 981.6000 ;
	    RECT 681.0000 981.3000 687.6000 982.2000 ;
	    RECT 686.4000 981.0000 687.6000 981.3000 ;
	    RECT 524.1000 978.6000 525.3000 978.9000 ;
	    RECT 517.8000 977.4000 519.0000 978.6000 ;
	    RECT 519.9000 977.7000 525.3000 978.6000 ;
	    RECT 520.2000 976.5000 528.6000 976.8000 ;
	    RECT 519.9000 976.2000 528.6000 976.5000 ;
	    RECT 503.4000 963.3000 504.6000 975.3000 ;
	    RECT 508.2000 974.7000 511.8000 975.6000 ;
	    RECT 513.9000 975.9000 528.6000 976.2000 ;
	    RECT 513.9000 975.3000 521.1000 975.9000 ;
	    RECT 508.2000 973.2000 509.1000 974.7000 ;
	    RECT 507.0000 972.0000 509.1000 973.2000 ;
	    RECT 511.5000 973.5000 512.7000 973.8000 ;
	    RECT 513.9000 973.5000 514.8000 975.3000 ;
	    RECT 511.5000 972.6000 514.8000 973.5000 ;
	    RECT 515.7000 973.5000 523.8000 974.4000 ;
	    RECT 515.7000 973.2000 516.9000 973.5000 ;
	    RECT 522.6000 973.2000 523.8000 973.5000 ;
	    RECT 513.3000 971.1000 514.5000 971.4000 ;
	    RECT 517.5000 971.1000 518.7000 971.4000 ;
	    RECT 508.2000 969.3000 509.4000 970.5000 ;
	    RECT 513.3000 970.2000 518.7000 971.1000 ;
	    RECT 514.5000 969.3000 515.4000 970.2000 ;
	    RECT 522.6000 969.3000 523.8000 970.5000 ;
	    RECT 507.3000 963.3000 509.1000 969.3000 ;
	    RECT 511.8000 963.3000 513.0000 969.3000 ;
	    RECT 514.2000 963.3000 515.4000 969.3000 ;
	    RECT 516.6000 963.3000 517.8000 969.3000 ;
	    RECT 520.8000 968.4000 523.8000 969.3000 ;
	    RECT 520.8000 963.3000 522.0000 968.4000 ;
	    RECT 525.0000 963.3000 526.2000 975.0000 ;
	    RECT 527.4000 963.3000 528.6000 975.9000 ;
	    RECT 659.4000 971.1000 660.6000 979.5000 ;
	    RECT 673.5000 978.9000 676.5000 980.1000 ;
	    RECT 682.2000 978.9000 687.0000 980.1000 ;
	    RECT 690.6000 979.2000 691.8000 983.4000 ;
	    RECT 697.8000 982.8000 699.0000 983.7000 ;
	    RECT 697.8000 981.9000 700.5000 982.8000 ;
	    RECT 699.3000 980.1000 700.5000 981.9000 ;
	    RECT 705.0000 981.9000 706.2000 989.7000 ;
	    RECT 707.4000 984.0000 708.6000 989.7000 ;
	    RECT 709.8000 986.7000 711.0000 989.7000 ;
	    RECT 729.9000 984.6000 731.1000 989.7000 ;
	    RECT 707.4000 982.8000 708.9000 984.0000 ;
	    RECT 729.9000 983.7000 732.6000 984.6000 ;
	    RECT 733.8000 983.7000 735.0000 989.7000 ;
	    RECT 745.8000 986.7000 747.0000 989.7000 ;
	    RECT 745.8000 985.5000 747.0000 985.8000 ;
	    RECT 705.0000 981.0000 706.8000 981.9000 ;
	    RECT 699.3000 978.9000 705.0000 980.1000 ;
	    RECT 661.5000 978.0000 662.7000 978.3000 ;
	    RECT 661.5000 977.1000 668.1000 978.0000 ;
	    RECT 669.0000 977.4000 670.2000 978.6000 ;
	    RECT 695.4000 978.0000 696.6000 978.9000 ;
	    RECT 705.9000 978.0000 706.8000 981.0000 ;
	    RECT 671.1000 977.1000 696.6000 978.0000 ;
	    RECT 705.6000 977.1000 706.8000 978.0000 ;
	    RECT 703.5000 976.2000 704.7000 976.5000 ;
	    RECT 664.2000 974.4000 665.4000 975.6000 ;
	    RECT 666.3000 975.3000 704.7000 976.2000 ;
	    RECT 669.3000 975.0000 670.5000 975.3000 ;
	    RECT 705.6000 974.4000 706.5000 977.1000 ;
	    RECT 707.7000 976.2000 708.9000 982.8000 ;
	    RECT 731.4000 979.5000 732.6000 983.7000 ;
	    RECT 745.8000 983.4000 747.0000 984.6000 ;
	    RECT 733.8000 982.5000 735.0000 982.8000 ;
	    RECT 748.2000 982.5000 749.4000 989.7000 ;
	    RECT 789.0000 983.7000 790.2000 989.7000 ;
	    RECT 791.4000 984.6000 792.9000 989.7000 ;
	    RECT 795.6000 984.3000 798.0000 989.7000 ;
	    RECT 800.7000 984.6000 802.2000 989.7000 ;
	    RECT 789.0000 982.8000 792.9000 983.7000 ;
	    RECT 791.7000 982.5000 792.9000 982.8000 ;
	    RECT 793.8000 982.2000 796.2000 983.4000 ;
	    RECT 733.8000 981.4500 735.0000 981.6000 ;
	    RECT 743.4000 981.4500 744.6000 981.6000 ;
	    RECT 733.8000 980.5500 744.6000 981.4500 ;
	    RECT 733.8000 980.4000 735.0000 980.5500 ;
	    RECT 743.4000 980.4000 744.6000 980.5500 ;
	    RECT 748.2000 981.4500 749.4000 981.6000 ;
	    RECT 767.4000 981.4500 768.6000 981.6000 ;
	    RECT 748.2000 980.5500 768.6000 981.4500 ;
	    RECT 748.2000 980.4000 749.4000 980.5500 ;
	    RECT 767.4000 980.4000 768.6000 980.5500 ;
	    RECT 789.0000 980.4000 790.2000 981.6000 ;
	    RECT 791.1000 981.3000 791.4000 981.6000 ;
	    RECT 797.1000 981.3000 798.0000 984.3000 ;
	    RECT 803.4000 983.7000 804.6000 989.7000 ;
	    RECT 817.8000 986.7000 819.0000 989.7000 ;
	    RECT 817.8000 985.5000 819.0000 985.8000 ;
	    RECT 798.9000 982.2000 800.1000 983.4000 ;
	    RECT 801.0000 982.8000 804.6000 983.7000 ;
	    RECT 815.4000 984.4500 816.6000 984.6000 ;
	    RECT 817.8000 984.4500 819.0000 984.6000 ;
	    RECT 815.4000 983.5500 819.0000 984.4500 ;
	    RECT 815.4000 983.4000 816.6000 983.5500 ;
	    RECT 817.8000 983.4000 819.0000 983.5500 ;
	    RECT 801.0000 982.5000 802.2000 982.8000 ;
	    RECT 820.2000 982.5000 821.4000 989.7000 ;
	    RECT 834.6000 982.5000 835.8000 989.7000 ;
	    RECT 837.0000 986.7000 838.2000 989.7000 ;
	    RECT 837.0000 985.5000 838.2000 985.8000 ;
	    RECT 837.0000 983.4000 838.2000 984.6000 ;
	    RECT 791.1000 981.0000 792.3000 981.3000 ;
	    RECT 791.1000 980.4000 795.6000 981.0000 ;
	    RECT 791.4000 980.1000 795.6000 980.4000 ;
	    RECT 794.4000 979.8000 795.6000 980.1000 ;
	    RECT 796.5000 980.4000 798.0000 981.3000 ;
	    RECT 799.2000 981.6000 800.1000 982.2000 ;
	    RECT 799.2000 980.4000 800.4000 981.6000 ;
	    RECT 802.2000 980.4000 802.5000 981.6000 ;
	    RECT 803.4000 980.4000 804.6000 981.6000 ;
	    RECT 820.2000 980.4000 821.4000 981.6000 ;
	    RECT 822.6000 981.4500 823.8000 981.6000 ;
	    RECT 834.6000 981.4500 835.8000 981.6000 ;
	    RECT 822.6000 980.5500 835.8000 981.4500 ;
	    RECT 863.4000 980.7000 864.6000 989.7000 ;
	    RECT 868.8000 981.3000 870.0000 989.7000 ;
	    RECT 889.8000 983.7000 891.0000 989.7000 ;
	    RECT 893.7000 984.6000 894.9000 989.7000 ;
	    RECT 916.2000 986.7000 917.4000 989.7000 ;
	    RECT 916.2000 985.5000 917.4000 985.8000 ;
	    RECT 892.2000 983.7000 894.9000 984.6000 ;
	    RECT 889.8000 982.5000 891.0000 982.8000 ;
	    RECT 868.8000 980.7000 871.5000 981.3000 ;
	    RECT 822.6000 980.4000 823.8000 980.5500 ;
	    RECT 834.6000 980.4000 835.8000 980.5500 ;
	    RECT 869.1000 980.4000 871.5000 980.7000 ;
	    RECT 889.8000 980.4000 891.0000 981.6000 ;
	    RECT 796.5000 979.5000 797.4000 980.4000 ;
	    RECT 731.4000 978.4500 732.6000 978.6000 ;
	    RECT 738.6000 978.4500 739.8000 978.6000 ;
	    RECT 731.4000 977.5500 739.8000 978.4500 ;
	    RECT 731.4000 977.4000 732.6000 977.5500 ;
	    RECT 738.6000 977.4000 739.8000 977.5500 ;
	    RECT 673.8000 974.1000 675.0000 974.4000 ;
	    RECT 666.9000 973.5000 675.0000 974.1000 ;
	    RECT 665.7000 973.2000 675.0000 973.5000 ;
	    RECT 676.5000 973.5000 689.4000 974.4000 ;
	    RECT 661.8000 972.0000 664.2000 973.2000 ;
	    RECT 665.7000 972.3000 667.8000 973.2000 ;
	    RECT 676.5000 972.3000 677.4000 973.5000 ;
	    RECT 688.2000 973.2000 689.4000 973.5000 ;
	    RECT 693.0000 973.5000 706.5000 974.4000 ;
	    RECT 707.4000 975.0000 708.9000 976.2000 ;
	    RECT 707.4000 973.5000 708.6000 975.0000 ;
	    RECT 729.0000 974.4000 730.2000 975.6000 ;
	    RECT 693.0000 973.2000 694.2000 973.5000 ;
	    RECT 663.3000 971.4000 664.2000 972.0000 ;
	    RECT 668.7000 971.4000 677.4000 972.3000 ;
	    RECT 678.3000 971.4000 682.2000 972.6000 ;
	    RECT 659.4000 970.2000 662.4000 971.1000 ;
	    RECT 663.3000 970.2000 669.6000 971.4000 ;
	    RECT 661.5000 969.3000 662.4000 970.2000 ;
	    RECT 659.4000 963.3000 660.6000 969.3000 ;
	    RECT 661.5000 968.4000 663.0000 969.3000 ;
	    RECT 661.8000 963.3000 663.0000 968.4000 ;
	    RECT 664.2000 962.4000 665.4000 969.3000 ;
	    RECT 666.6000 963.3000 667.8000 970.2000 ;
	    RECT 669.0000 963.3000 670.2000 969.3000 ;
	    RECT 671.4000 963.3000 672.6000 967.5000 ;
	    RECT 673.8000 963.3000 675.0000 967.5000 ;
	    RECT 676.2000 963.3000 677.4000 970.5000 ;
	    RECT 678.6000 963.3000 679.8000 969.3000 ;
	    RECT 681.0000 963.3000 682.2000 970.5000 ;
	    RECT 683.4000 963.3000 684.6000 969.3000 ;
	    RECT 685.8000 963.3000 687.0000 972.6000 ;
	    RECT 697.8000 971.4000 701.7000 972.6000 ;
	    RECT 690.6000 970.2000 696.9000 971.4000 ;
	    RECT 688.2000 963.3000 689.4000 967.5000 ;
	    RECT 690.6000 963.3000 691.8000 967.5000 ;
	    RECT 693.0000 963.3000 694.2000 967.5000 ;
	    RECT 695.4000 963.3000 696.6000 969.3000 ;
	    RECT 697.8000 963.3000 699.0000 971.4000 ;
	    RECT 705.6000 971.1000 706.5000 973.5000 ;
	    RECT 729.0000 973.2000 730.2000 973.5000 ;
	    RECT 707.4000 971.4000 708.6000 972.6000 ;
	    RECT 702.6000 970.2000 706.5000 971.1000 ;
	    RECT 700.2000 963.3000 701.4000 969.3000 ;
	    RECT 702.6000 963.3000 703.8000 970.2000 ;
	    RECT 705.0000 963.3000 706.2000 969.3000 ;
	    RECT 707.4000 963.3000 708.6000 970.5000 ;
	    RECT 709.8000 963.3000 711.0000 969.3000 ;
	    RECT 729.0000 963.3000 730.2000 969.3000 ;
	    RECT 731.4000 963.3000 732.6000 976.5000 ;
	    RECT 733.8000 963.3000 735.0000 969.3000 ;
	    RECT 745.8000 963.3000 747.0000 969.3000 ;
	    RECT 748.2000 963.3000 749.4000 979.5000 ;
	    RECT 792.3000 978.3000 793.5000 978.6000 ;
	    RECT 796.2000 978.4500 797.4000 978.6000 ;
	    RECT 817.8000 978.4500 819.0000 978.6000 ;
	    RECT 792.3000 977.4000 794.7000 978.3000 ;
	    RECT 796.2000 977.5500 819.0000 978.4500 ;
	    RECT 796.2000 977.4000 797.4000 977.5500 ;
	    RECT 817.8000 977.4000 819.0000 977.5500 ;
	    RECT 793.5000 977.1000 794.7000 977.4000 ;
	    RECT 796.5000 975.3000 797.4000 976.5000 ;
	    RECT 789.0000 974.4000 792.9000 975.3000 ;
	    RECT 765.0000 969.4500 766.2000 969.6000 ;
	    RECT 786.6000 969.4500 787.8000 969.6000 ;
	    RECT 765.0000 968.5500 787.8000 969.4500 ;
	    RECT 765.0000 968.4000 766.2000 968.5500 ;
	    RECT 786.6000 968.4000 787.8000 968.5500 ;
	    RECT 762.6000 966.4500 763.8000 966.6000 ;
	    RECT 769.8000 966.4500 771.0000 966.6000 ;
	    RECT 762.6000 965.5500 771.0000 966.4500 ;
	    RECT 762.6000 965.4000 763.8000 965.5500 ;
	    RECT 769.8000 965.4000 771.0000 965.5500 ;
	    RECT 789.0000 963.3000 790.2000 974.4000 ;
	    RECT 791.7000 974.1000 792.9000 974.4000 ;
	    RECT 791.4000 963.3000 792.9000 973.2000 ;
	    RECT 795.6000 963.3000 798.0000 975.3000 ;
	    RECT 801.0000 974.4000 804.6000 975.3000 ;
	    RECT 801.0000 974.1000 802.2000 974.4000 ;
	    RECT 800.7000 963.3000 802.2000 973.2000 ;
	    RECT 803.4000 963.3000 804.6000 974.4000 ;
	    RECT 817.8000 963.3000 819.0000 969.3000 ;
	    RECT 820.2000 963.3000 821.4000 979.5000 ;
	    RECT 834.6000 963.3000 835.8000 979.5000 ;
	    RECT 865.8000 977.4000 867.0000 978.6000 ;
	    RECT 867.9000 977.4000 868.2000 978.6000 ;
	    RECT 863.4000 976.5000 864.6000 976.8000 ;
	    RECT 870.6000 976.5000 871.5000 980.4000 ;
	    RECT 892.2000 979.5000 893.4000 983.7000 ;
	    RECT 916.2000 983.4000 917.4000 984.6000 ;
	    RECT 918.6000 982.5000 919.8000 989.7000 ;
	    RECT 923.4000 987.4500 924.6000 987.6000 ;
	    RECT 935.4000 987.4500 936.6000 987.6000 ;
	    RECT 923.4000 986.5500 936.6000 987.4500 ;
	    RECT 923.4000 986.4000 924.6000 986.5500 ;
	    RECT 935.4000 986.4000 936.6000 986.5500 ;
	    RECT 947.4000 984.0000 948.6000 989.7000 ;
	    RECT 949.8000 984.9000 951.0000 989.7000 ;
	    RECT 952.2000 988.8000 958.2000 989.7000 ;
	    RECT 952.2000 984.0000 953.4000 988.8000 ;
	    RECT 947.4000 983.7000 953.4000 984.0000 ;
	    RECT 954.6000 983.7000 955.8000 987.9000 ;
	    RECT 957.0000 983.7000 958.2000 988.8000 ;
	    RECT 947.7000 983.1000 953.1000 983.7000 ;
	    RECT 918.6000 981.4500 919.8000 981.6000 ;
	    RECT 947.4000 981.4500 948.6000 981.6000 ;
	    RECT 918.6000 980.5500 948.6000 981.4500 ;
	    RECT 949.5000 980.7000 949.8000 982.2000 ;
	    RECT 954.9000 981.6000 955.8000 983.7000 ;
	    RECT 971.4000 982.5000 972.6000 989.7000 ;
	    RECT 973.8000 986.7000 975.0000 989.7000 ;
	    RECT 988.2000 986.7000 989.4000 989.7000 ;
	    RECT 973.8000 985.5000 975.0000 985.8000 ;
	    RECT 988.2000 985.5000 989.4000 985.8000 ;
	    RECT 973.8000 983.4000 975.0000 984.6000 ;
	    RECT 988.2000 983.4000 989.4000 984.6000 ;
	    RECT 990.6000 982.5000 991.8000 989.7000 ;
	    RECT 1021.8000 984.0000 1023.0000 989.7000 ;
	    RECT 1024.2001 984.9000 1025.4000 989.7000 ;
	    RECT 1026.6000 988.8000 1032.6000 989.7000 ;
	    RECT 1026.6000 984.0000 1027.8000 988.8000 ;
	    RECT 1021.8000 983.7000 1027.8000 984.0000 ;
	    RECT 1029.0000 983.7000 1030.2001 987.9000 ;
	    RECT 1031.4000 983.7000 1032.6000 988.8000 ;
	    RECT 1043.4000 986.7000 1044.6000 989.7000 ;
	    RECT 1043.4000 985.5000 1044.6000 985.8000 ;
	    RECT 1022.1000 983.1000 1027.5000 983.7000 ;
	    RECT 918.6000 980.4000 919.8000 980.5500 ;
	    RECT 947.4000 980.4000 948.6000 980.5500 ;
	    RECT 952.2000 980.4000 953.4000 981.6000 ;
	    RECT 954.3000 980.7000 955.8000 981.6000 ;
	    RECT 957.0000 981.4500 958.2000 981.6000 ;
	    RECT 971.4000 981.4500 972.6000 981.6000 ;
	    RECT 957.0000 980.5500 972.6000 981.4500 ;
	    RECT 957.0000 980.4000 958.2000 980.5500 ;
	    RECT 971.4000 980.4000 972.6000 980.5500 ;
	    RECT 990.6000 981.4500 991.8000 981.6000 ;
	    RECT 1021.8000 981.4500 1023.0000 981.6000 ;
	    RECT 990.6000 980.5500 1023.0000 981.4500 ;
	    RECT 1023.9000 980.7000 1024.2001 982.2000 ;
	    RECT 1029.3000 981.6000 1030.2001 983.7000 ;
	    RECT 1043.4000 983.4000 1044.6000 984.6000 ;
	    RECT 1045.8000 982.5000 1047.0000 989.7000 ;
	    RECT 1072.2001 984.0000 1073.4000 989.7000 ;
	    RECT 1074.6000 984.9000 1075.8000 989.7000 ;
	    RECT 1077.0000 984.0000 1078.2001 989.7000 ;
	    RECT 1072.2001 983.7000 1078.2001 984.0000 ;
	    RECT 1079.4000 983.7000 1080.6000 989.7000 ;
	    RECT 1103.4000 983.7000 1104.6000 989.7000 ;
	    RECT 1105.8000 984.0000 1107.0000 989.7000 ;
	    RECT 1108.2001 984.9000 1109.4000 989.7000 ;
	    RECT 1110.6000 984.0000 1111.8000 989.7000 ;
	    RECT 1105.8000 983.7000 1111.8000 984.0000 ;
	    RECT 1072.5000 983.1000 1077.9000 983.7000 ;
	    RECT 1079.4000 982.5000 1080.3000 983.7000 ;
	    RECT 1103.7001 982.5000 1104.6000 983.7000 ;
	    RECT 1106.1000 983.1000 1111.5000 983.7000 ;
	    RECT 1132.2001 982.5000 1133.4000 989.7000 ;
	    RECT 1134.6000 986.7000 1135.8000 989.7000 ;
	    RECT 1134.6000 985.5000 1135.8000 985.8000 ;
	    RECT 1134.6000 983.4000 1135.8000 984.6000 ;
	    RECT 1146.6000 982.5000 1147.8000 989.7000 ;
	    RECT 1149.0000 986.7000 1150.2001 989.7000 ;
	    RECT 1163.4000 986.7000 1164.6000 989.7000 ;
	    RECT 1149.0000 985.5000 1150.2001 985.8000 ;
	    RECT 1163.4000 985.5000 1164.6000 985.8000 ;
	    RECT 1149.0000 983.4000 1150.2001 984.6000 ;
	    RECT 1163.4000 983.4000 1164.6000 984.6000 ;
	    RECT 1165.8000 982.5000 1167.0000 989.7000 ;
	    RECT 1192.2001 984.0000 1193.4000 989.7000 ;
	    RECT 1194.6000 984.9000 1195.8000 989.7000 ;
	    RECT 1197.0000 984.0000 1198.2001 989.7000 ;
	    RECT 1192.2001 983.7000 1198.2001 984.0000 ;
	    RECT 1199.4000 983.7000 1200.6000 989.7000 ;
	    RECT 1219.5000 984.6000 1220.7001 989.7000 ;
	    RECT 1219.5000 983.7000 1222.2001 984.6000 ;
	    RECT 1223.4000 983.7000 1224.6000 989.7000 ;
	    RECT 1192.5000 983.1000 1197.9000 983.7000 ;
	    RECT 1199.4000 982.5000 1200.3000 983.7000 ;
	    RECT 990.6000 980.4000 991.8000 980.5500 ;
	    RECT 1021.8000 980.4000 1023.0000 980.5500 ;
	    RECT 1026.6000 980.4000 1027.8000 981.6000 ;
	    RECT 1028.7001 980.7000 1030.2001 981.6000 ;
	    RECT 1031.4000 980.4000 1032.6000 981.6000 ;
	    RECT 1045.8000 981.4500 1047.0000 981.6000 ;
	    RECT 1045.8000 980.5500 1066.0500 981.4500 ;
	    RECT 1045.8000 980.4000 1047.0000 980.5500 ;
	    RECT 949.8000 979.5000 951.0000 979.8000 ;
	    RECT 954.6000 979.5000 955.8000 979.8000 ;
	    RECT 1024.2001 979.5000 1025.4000 979.8000 ;
	    RECT 1029.0000 979.5000 1030.2001 979.8000 ;
	    RECT 892.2000 978.4500 893.4000 978.6000 ;
	    RECT 913.8000 978.4500 915.0000 978.6000 ;
	    RECT 892.2000 977.5500 915.0000 978.4500 ;
	    RECT 892.2000 977.4000 893.4000 977.5500 ;
	    RECT 913.8000 977.4000 915.0000 977.5500 ;
	    RECT 839.4000 975.4500 840.6000 975.6000 ;
	    RECT 863.4000 975.4500 864.6000 975.6000 ;
	    RECT 839.4000 974.5500 864.6000 975.4500 ;
	    RECT 839.4000 974.4000 840.6000 974.5500 ;
	    RECT 863.4000 974.4000 864.6000 974.5500 ;
	    RECT 870.6000 975.4500 871.8000 975.6000 ;
	    RECT 889.8000 975.4500 891.0000 975.6000 ;
	    RECT 870.6000 974.5500 891.0000 975.4500 ;
	    RECT 870.6000 974.4000 871.8000 974.5500 ;
	    RECT 889.8000 974.4000 891.0000 974.5500 ;
	    RECT 868.2000 973.5000 869.4000 973.8000 ;
	    RECT 868.2000 971.4000 869.4000 972.6000 ;
	    RECT 870.6000 970.5000 871.5000 973.5000 ;
	    RECT 866.1000 969.6000 871.5000 970.5000 ;
	    RECT 866.1000 969.3000 867.0000 969.6000 ;
	    RECT 837.0000 963.3000 838.2000 969.3000 ;
	    RECT 863.4000 963.3000 864.6000 969.3000 ;
	    RECT 865.8000 963.3000 867.0000 969.3000 ;
	    RECT 870.6000 969.3000 871.5000 969.6000 ;
	    RECT 868.2000 963.3000 869.4000 968.7000 ;
	    RECT 870.6000 963.3000 871.8000 969.3000 ;
	    RECT 889.8000 963.3000 891.0000 969.3000 ;
	    RECT 892.2000 963.3000 893.4000 976.5000 ;
	    RECT 894.6000 974.4000 895.8000 975.6000 ;
	    RECT 894.6000 973.2000 895.8000 973.5000 ;
	    RECT 894.6000 963.3000 895.8000 969.3000 ;
	    RECT 916.2000 963.3000 917.4000 969.3000 ;
	    RECT 918.6000 963.3000 919.8000 979.5000 ;
	    RECT 921.0000 978.4500 922.2000 978.6000 ;
	    RECT 949.8000 978.4500 951.0000 978.6000 ;
	    RECT 921.0000 977.5500 951.0000 978.4500 ;
	    RECT 921.0000 977.4000 922.2000 977.5500 ;
	    RECT 949.8000 977.4000 951.0000 977.5500 ;
	    RECT 952.2000 975.3000 953.1000 979.5000 ;
	    RECT 957.0000 979.2000 958.2000 979.5000 ;
	    RECT 954.6000 977.4000 955.8000 978.6000 ;
	    RECT 947.4000 963.3000 948.6000 975.3000 ;
	    RECT 951.3000 963.3000 954.3000 975.3000 ;
	    RECT 957.0000 963.3000 958.2000 975.3000 ;
	    RECT 971.4000 963.3000 972.6000 979.5000 ;
	    RECT 973.8000 963.3000 975.0000 969.3000 ;
	    RECT 988.2000 963.3000 989.4000 969.3000 ;
	    RECT 990.6000 963.3000 991.8000 979.5000 ;
	    RECT 993.0000 978.4500 994.2000 978.6000 ;
	    RECT 1002.6000 978.4500 1003.8000 978.6000 ;
	    RECT 1024.2001 978.4500 1025.4000 978.6000 ;
	    RECT 993.0000 977.5500 1025.4000 978.4500 ;
	    RECT 993.0000 977.4000 994.2000 977.5500 ;
	    RECT 1002.6000 977.4000 1003.8000 977.5500 ;
	    RECT 1024.2001 977.4000 1025.4000 977.5500 ;
	    RECT 1026.6000 975.3000 1027.5000 979.5000 ;
	    RECT 1031.4000 979.2000 1032.6000 979.5000 ;
	    RECT 1029.0000 977.4000 1030.2001 978.6000 ;
	    RECT 1021.8000 963.3000 1023.0000 975.3000 ;
	    RECT 1025.7001 963.3000 1028.7001 975.3000 ;
	    RECT 1031.4000 963.3000 1032.6000 975.3000 ;
	    RECT 1043.4000 963.3000 1044.6000 969.3000 ;
	    RECT 1045.8000 963.3000 1047.0000 979.5000 ;
	    RECT 1065.1500 978.4500 1066.0500 980.5500 ;
	    RECT 1072.2001 980.4000 1073.4000 981.6000 ;
	    RECT 1074.3000 980.7000 1074.6000 982.2000 ;
	    RECT 1076.7001 980.4000 1078.5000 981.6000 ;
	    RECT 1079.4000 981.4500 1080.6000 981.6000 ;
	    RECT 1084.2001 981.4500 1085.4000 981.6000 ;
	    RECT 1079.4000 980.5500 1085.4000 981.4500 ;
	    RECT 1079.4000 980.4000 1080.6000 980.5500 ;
	    RECT 1084.2001 980.4000 1085.4000 980.5500 ;
	    RECT 1103.4000 980.4000 1104.6000 981.6000 ;
	    RECT 1105.5000 980.4000 1107.3000 981.6000 ;
	    RECT 1109.4000 980.7000 1109.7001 982.2000 ;
	    RECT 1110.6000 981.4500 1111.8000 981.6000 ;
	    RECT 1129.8000 981.4500 1131.0000 981.6000 ;
	    RECT 1110.6000 980.5500 1131.0000 981.4500 ;
	    RECT 1110.6000 980.4000 1111.8000 980.5500 ;
	    RECT 1129.8000 980.4000 1131.0000 980.5500 ;
	    RECT 1132.2001 980.4000 1133.4000 981.6000 ;
	    RECT 1137.0000 981.4500 1138.2001 981.6000 ;
	    RECT 1146.6000 981.4500 1147.8000 981.6000 ;
	    RECT 1137.0000 980.5500 1147.8000 981.4500 ;
	    RECT 1137.0000 980.4000 1138.2001 980.5500 ;
	    RECT 1146.6000 980.4000 1147.8000 980.5500 ;
	    RECT 1165.8000 981.4500 1167.0000 981.6000 ;
	    RECT 1189.8000 981.4500 1191.0000 981.6000 ;
	    RECT 1192.2001 981.4500 1193.4000 981.6000 ;
	    RECT 1165.8000 980.5500 1188.4501 981.4500 ;
	    RECT 1165.8000 980.4000 1167.0000 980.5500 ;
	    RECT 1074.6000 979.5000 1075.8000 979.8000 ;
	    RECT 1074.6000 978.4500 1075.8000 978.6000 ;
	    RECT 1065.1500 977.5500 1075.8000 978.4500 ;
	    RECT 1074.6000 977.4000 1075.8000 977.5500 ;
	    RECT 1076.7001 975.3000 1077.6000 980.4000 ;
	    RECT 1072.2001 963.3000 1073.4000 975.3000 ;
	    RECT 1076.1000 974.4000 1077.6000 975.3000 ;
	    RECT 1079.4000 974.4000 1080.6000 975.6000 ;
	    RECT 1093.8000 975.4500 1095.0000 975.6000 ;
	    RECT 1103.4000 975.4500 1104.6000 975.6000 ;
	    RECT 1093.8000 974.5500 1104.6000 975.4500 ;
	    RECT 1093.8000 974.4000 1095.0000 974.5500 ;
	    RECT 1103.4000 974.4000 1104.6000 974.5500 ;
	    RECT 1106.4000 975.3000 1107.3000 980.4000 ;
	    RECT 1108.2001 979.5000 1109.4000 979.8000 ;
	    RECT 1108.2001 978.4500 1109.4000 978.6000 ;
	    RECT 1122.6000 978.4500 1123.8000 978.6000 ;
	    RECT 1108.2001 977.5500 1123.8000 978.4500 ;
	    RECT 1108.2001 977.4000 1109.4000 977.5500 ;
	    RECT 1122.6000 977.4000 1123.8000 977.5500 ;
	    RECT 1106.4000 974.4000 1107.9000 975.3000 ;
	    RECT 1076.1000 963.3000 1077.3000 974.4000 ;
	    RECT 1078.5000 972.6000 1079.4000 973.5000 ;
	    RECT 1078.2001 971.4000 1079.4000 972.6000 ;
	    RECT 1104.6000 972.6000 1105.5000 973.5000 ;
	    RECT 1104.6000 971.4000 1105.8000 972.6000 ;
	    RECT 1078.5000 963.3000 1079.7001 969.3000 ;
	    RECT 1104.3000 963.3000 1105.5000 969.3000 ;
	    RECT 1106.7001 963.3000 1107.9000 974.4000 ;
	    RECT 1110.6000 963.3000 1111.8000 975.3000 ;
	    RECT 1132.2001 963.3000 1133.4000 979.5000 ;
	    RECT 1134.6000 963.3000 1135.8000 969.3000 ;
	    RECT 1146.6000 963.3000 1147.8000 979.5000 ;
	    RECT 1149.0000 963.3000 1150.2001 969.3000 ;
	    RECT 1163.4000 963.3000 1164.6000 969.3000 ;
	    RECT 1165.8000 963.3000 1167.0000 979.5000 ;
	    RECT 1187.5500 978.4500 1188.4501 980.5500 ;
	    RECT 1189.8000 980.5500 1193.4000 981.4500 ;
	    RECT 1194.3000 980.7000 1194.6000 982.2000 ;
	    RECT 1189.8000 980.4000 1191.0000 980.5500 ;
	    RECT 1192.2001 980.4000 1193.4000 980.5500 ;
	    RECT 1196.7001 980.4000 1198.5000 981.6000 ;
	    RECT 1199.4000 981.4500 1200.6000 981.6000 ;
	    RECT 1201.8000 981.4500 1203.0000 981.6000 ;
	    RECT 1199.4000 980.5500 1203.0000 981.4500 ;
	    RECT 1199.4000 980.4000 1200.6000 980.5500 ;
	    RECT 1201.8000 980.4000 1203.0000 980.5500 ;
	    RECT 1194.6000 979.5000 1195.8000 979.8000 ;
	    RECT 1194.6000 978.4500 1195.8000 978.6000 ;
	    RECT 1187.5500 977.5500 1195.8000 978.4500 ;
	    RECT 1194.6000 977.4000 1195.8000 977.5500 ;
	    RECT 1196.7001 975.3000 1197.6000 980.4000 ;
	    RECT 1221.0000 979.5000 1222.2001 983.7000 ;
	    RECT 1223.4000 982.5000 1224.6000 982.8000 ;
	    RECT 1237.8000 982.5000 1239.0000 989.7000 ;
	    RECT 1240.2001 986.7000 1241.4000 989.7000 ;
	    RECT 1240.2001 985.5000 1241.4000 985.8000 ;
	    RECT 1240.2001 984.4500 1241.4000 984.6000 ;
	    RECT 1261.8000 984.4500 1263.0000 984.6000 ;
	    RECT 1240.2001 983.5500 1263.0000 984.4500 ;
	    RECT 1264.2001 984.0000 1265.4000 989.7000 ;
	    RECT 1266.6000 984.9000 1267.8000 989.7000 ;
	    RECT 1269.0000 984.0000 1270.2001 989.7000 ;
	    RECT 1264.2001 983.7000 1270.2001 984.0000 ;
	    RECT 1271.4000 983.7000 1272.6000 989.7000 ;
	    RECT 1295.4000 986.7000 1296.6000 989.7000 ;
	    RECT 1295.7001 985.5000 1296.9000 985.8000 ;
	    RECT 1293.0000 984.4500 1294.2001 984.6000 ;
	    RECT 1295.4000 984.4500 1296.6000 984.6000 ;
	    RECT 1240.2001 983.4000 1241.4000 983.5500 ;
	    RECT 1261.8000 983.4000 1263.0000 983.5500 ;
	    RECT 1264.5000 983.1000 1269.9000 983.7000 ;
	    RECT 1271.4000 982.5000 1272.3000 983.7000 ;
	    RECT 1293.0000 983.5500 1296.6000 984.4500 ;
	    RECT 1297.8000 983.7000 1299.0000 989.7000 ;
	    RECT 1301.7001 983.7000 1302.9000 989.7000 ;
	    RECT 1326.6000 983.7000 1327.8000 989.7000 ;
	    RECT 1329.0000 984.0000 1330.2001 989.7000 ;
	    RECT 1331.4000 984.9000 1332.6000 989.7000 ;
	    RECT 1333.8000 984.0000 1335.0000 989.7000 ;
	    RECT 1348.2001 986.7000 1349.4000 989.7000 ;
	    RECT 1348.2001 985.5000 1349.4000 985.8000 ;
	    RECT 1329.0000 983.7000 1335.0000 984.0000 ;
	    RECT 1345.8000 984.4500 1347.0000 984.6000 ;
	    RECT 1348.2001 984.4500 1349.4000 984.6000 ;
	    RECT 1293.0000 983.4000 1294.2001 983.5500 ;
	    RECT 1295.4000 983.4000 1296.6000 983.5500 ;
	    RECT 1223.4000 981.4500 1224.6000 981.6000 ;
	    RECT 1235.4000 981.4500 1236.6000 981.6000 ;
	    RECT 1223.4000 980.5500 1236.6000 981.4500 ;
	    RECT 1223.4000 980.4000 1224.6000 980.5500 ;
	    RECT 1235.4000 980.4000 1236.6000 980.5500 ;
	    RECT 1237.8000 981.4500 1239.0000 981.6000 ;
	    RECT 1237.8000 980.5500 1262.8500 981.4500 ;
	    RECT 1237.8000 980.4000 1239.0000 980.5500 ;
	    RECT 1221.0000 978.4500 1222.2001 978.6000 ;
	    RECT 1235.4000 978.4500 1236.6000 978.6000 ;
	    RECT 1221.0000 977.5500 1236.6000 978.4500 ;
	    RECT 1221.0000 977.4000 1222.2001 977.5500 ;
	    RECT 1235.4000 977.4000 1236.6000 977.5500 ;
	    RECT 1192.2001 963.3000 1193.4000 975.3000 ;
	    RECT 1196.1000 974.4000 1197.6000 975.3000 ;
	    RECT 1199.4000 974.4000 1200.6000 975.6000 ;
	    RECT 1204.2001 975.4500 1205.4000 975.6000 ;
	    RECT 1218.6000 975.4500 1219.8000 975.6000 ;
	    RECT 1204.2001 974.5500 1219.8000 975.4500 ;
	    RECT 1204.2001 974.4000 1205.4000 974.5500 ;
	    RECT 1218.6000 974.4000 1219.8000 974.5500 ;
	    RECT 1196.1000 963.3000 1197.3000 974.4000 ;
	    RECT 1198.5000 972.6000 1199.4000 973.5000 ;
	    RECT 1218.6000 973.2000 1219.8000 973.5000 ;
	    RECT 1198.2001 971.4000 1199.4000 972.6000 ;
	    RECT 1198.5000 963.3000 1199.7001 969.3000 ;
	    RECT 1218.6000 963.3000 1219.8000 969.3000 ;
	    RECT 1221.0000 963.3000 1222.2001 976.5000 ;
	    RECT 1223.4000 963.3000 1224.6000 969.3000 ;
	    RECT 1237.8000 963.3000 1239.0000 979.5000 ;
	    RECT 1261.9501 978.4500 1262.8500 980.5500 ;
	    RECT 1264.2001 980.4000 1265.4000 981.6000 ;
	    RECT 1266.3000 980.7000 1266.6000 982.2000 ;
	    RECT 1268.7001 980.4000 1270.5000 981.6000 ;
	    RECT 1271.4000 981.4500 1272.6000 981.6000 ;
	    RECT 1295.4000 981.4500 1296.6000 981.6000 ;
	    RECT 1271.4000 980.5500 1296.6000 981.4500 ;
	    RECT 1271.4000 980.4000 1272.6000 980.5500 ;
	    RECT 1295.4000 980.4000 1296.6000 980.5500 ;
	    RECT 1266.6000 979.5000 1267.8000 979.8000 ;
	    RECT 1266.6000 978.4500 1267.8000 978.6000 ;
	    RECT 1261.9501 977.5500 1267.8000 978.4500 ;
	    RECT 1266.6000 977.4000 1267.8000 977.5500 ;
	    RECT 1268.7001 975.3000 1269.6000 980.4000 ;
	    RECT 1285.8000 978.4500 1287.0000 978.6000 ;
	    RECT 1295.4000 978.4500 1296.6000 978.6000 ;
	    RECT 1285.8000 977.5500 1296.6000 978.4500 ;
	    RECT 1298.1000 978.3000 1299.0000 983.7000 ;
	    RECT 1326.9000 982.5000 1327.8000 983.7000 ;
	    RECT 1329.3000 983.1000 1334.7001 983.7000 ;
	    RECT 1345.8000 983.5500 1349.4000 984.4500 ;
	    RECT 1345.8000 983.4000 1347.0000 983.5500 ;
	    RECT 1348.2001 983.4000 1349.4000 983.5500 ;
	    RECT 1350.6000 982.5000 1351.8000 989.7000 ;
	    RECT 1377.0000 983.7000 1378.2001 989.7000 ;
	    RECT 1380.9000 984.6000 1382.1000 989.7000 ;
	    RECT 1379.4000 983.7000 1382.1000 984.6000 ;
	    RECT 1377.0000 982.5000 1378.2001 982.8000 ;
	    RECT 1300.2001 980.4000 1301.4000 981.6000 ;
	    RECT 1317.0000 981.4500 1318.2001 981.6000 ;
	    RECT 1326.6000 981.4500 1327.8000 981.6000 ;
	    RECT 1317.0000 980.5500 1327.8000 981.4500 ;
	    RECT 1317.0000 980.4000 1318.2001 980.5500 ;
	    RECT 1326.6000 980.4000 1327.8000 980.5500 ;
	    RECT 1328.7001 980.4000 1330.5000 981.6000 ;
	    RECT 1332.6000 980.7000 1332.9000 982.2000 ;
	    RECT 1333.8000 980.4000 1335.0000 981.6000 ;
	    RECT 1350.6000 981.4500 1351.8000 981.6000 ;
	    RECT 1336.3500 980.5500 1351.8000 981.4500 ;
	    RECT 1300.2001 979.2000 1301.4000 979.5000 ;
	    RECT 1285.8000 977.4000 1287.0000 977.5500 ;
	    RECT 1295.4000 977.4000 1296.6000 977.5500 ;
	    RECT 1297.5000 977.4000 1299.0000 978.3000 ;
	    RECT 1301.4000 976.8000 1301.7001 978.3000 ;
	    RECT 1302.6000 977.4000 1303.8000 978.6000 ;
	    RECT 1240.2001 963.3000 1241.4000 969.3000 ;
	    RECT 1264.2001 963.3000 1265.4000 975.3000 ;
	    RECT 1268.1000 974.4000 1269.6000 975.3000 ;
	    RECT 1271.4000 974.4000 1272.6000 975.6000 ;
	    RECT 1295.7001 975.3000 1296.6000 976.5000 ;
	    RECT 1268.1000 963.3000 1269.3000 974.4000 ;
	    RECT 1270.5000 972.6000 1271.4000 973.5000 ;
	    RECT 1270.2001 971.4000 1271.4000 972.6000 ;
	    RECT 1270.5000 963.3000 1271.7001 969.3000 ;
	    RECT 1295.4000 963.3000 1296.6000 975.3000 ;
	    RECT 1297.8000 974.4000 1303.8000 975.3000 ;
	    RECT 1326.6000 974.4000 1327.8000 975.6000 ;
	    RECT 1329.6000 975.3000 1330.5000 980.4000 ;
	    RECT 1331.4000 979.5000 1332.6000 979.8000 ;
	    RECT 1331.4000 978.4500 1332.6000 978.6000 ;
	    RECT 1336.3500 978.4500 1337.2500 980.5500 ;
	    RECT 1350.6000 980.4000 1351.8000 980.5500 ;
	    RECT 1377.0000 980.4000 1378.2001 981.6000 ;
	    RECT 1379.4000 979.5000 1380.6000 983.7000 ;
	    RECT 1407.6000 981.3000 1408.8000 989.7000 ;
	    RECT 1406.1000 980.7000 1408.8000 981.3000 ;
	    RECT 1413.0000 980.7000 1414.2001 989.7000 ;
	    RECT 1433.1000 984.6000 1434.3000 989.7000 ;
	    RECT 1433.1000 983.7000 1435.8000 984.6000 ;
	    RECT 1437.0000 983.7000 1438.2001 989.7000 ;
	    RECT 1461.0000 986.7000 1462.2001 989.7000 ;
	    RECT 1461.3000 985.5000 1462.5000 985.8000 ;
	    RECT 1451.4000 984.4500 1452.6000 984.6000 ;
	    RECT 1461.0000 984.4500 1462.2001 984.6000 ;
	    RECT 1406.1000 980.4000 1408.5000 980.7000 ;
	    RECT 1331.4000 977.5500 1337.2500 978.4500 ;
	    RECT 1331.4000 977.4000 1332.6000 977.5500 ;
	    RECT 1329.6000 974.4000 1331.1000 975.3000 ;
	    RECT 1297.8000 963.3000 1299.0000 974.4000 ;
	    RECT 1300.2001 963.3000 1301.4000 973.5000 ;
	    RECT 1302.6000 963.3000 1303.8000 974.4000 ;
	    RECT 1327.8000 972.6000 1328.7001 973.5000 ;
	    RECT 1327.8000 971.4000 1329.0000 972.6000 ;
	    RECT 1327.5000 963.3000 1328.7001 969.3000 ;
	    RECT 1329.9000 963.3000 1331.1000 974.4000 ;
	    RECT 1333.8000 963.3000 1335.0000 975.3000 ;
	    RECT 1348.2001 963.3000 1349.4000 969.3000 ;
	    RECT 1350.6000 963.3000 1351.8000 979.5000 ;
	    RECT 1353.0000 978.4500 1354.2001 978.6000 ;
	    RECT 1379.4000 978.4500 1380.6000 978.6000 ;
	    RECT 1353.0000 977.5500 1380.6000 978.4500 ;
	    RECT 1353.0000 977.4000 1354.2001 977.5500 ;
	    RECT 1379.4000 977.4000 1380.6000 977.5500 ;
	    RECT 1406.1000 976.5000 1407.0000 980.4000 ;
	    RECT 1434.6000 979.5000 1435.8000 983.7000 ;
	    RECT 1451.4000 983.5500 1462.2001 984.4500 ;
	    RECT 1463.4000 983.7000 1464.6000 989.7000 ;
	    RECT 1467.3000 983.7000 1468.5000 989.7000 ;
	    RECT 1487.4000 983.7000 1488.6000 989.7000 ;
	    RECT 1491.3000 984.6000 1492.5000 989.7000 ;
	    RECT 1489.8000 983.7000 1492.5000 984.6000 ;
	    RECT 1517.1000 983.7000 1518.3000 989.7000 ;
	    RECT 1521.0000 983.7000 1522.2001 989.7000 ;
	    RECT 1523.4000 986.7000 1524.6000 989.7000 ;
	    RECT 1523.1000 985.5000 1524.3000 985.8000 ;
	    RECT 1451.4000 983.4000 1452.6000 983.5500 ;
	    RECT 1461.0000 983.4000 1462.2001 983.5500 ;
	    RECT 1437.0000 982.5000 1438.2001 982.8000 ;
	    RECT 1437.0000 980.4000 1438.2001 981.6000 ;
	    RECT 1409.4000 977.4000 1409.7001 978.6000 ;
	    RECT 1410.6000 977.4000 1411.8000 978.6000 ;
	    RECT 1434.6000 977.4000 1435.8000 978.6000 ;
	    RECT 1439.4000 978.4500 1440.6000 978.6000 ;
	    RECT 1461.0000 978.4500 1462.2001 978.6000 ;
	    RECT 1439.4000 977.5500 1462.2001 978.4500 ;
	    RECT 1463.7001 978.3000 1464.6000 983.7000 ;
	    RECT 1487.4000 982.5000 1488.6000 982.8000 ;
	    RECT 1465.8000 980.4000 1467.0000 981.6000 ;
	    RECT 1482.6000 981.4500 1483.8000 981.6000 ;
	    RECT 1487.4000 981.4500 1488.6000 981.6000 ;
	    RECT 1482.6000 980.5500 1488.6000 981.4500 ;
	    RECT 1482.6000 980.4000 1483.8000 980.5500 ;
	    RECT 1487.4000 980.4000 1488.6000 980.5500 ;
	    RECT 1489.8000 979.5000 1491.0000 983.7000 ;
	    RECT 1518.6000 980.4000 1519.8000 981.6000 ;
	    RECT 1465.8000 979.2000 1467.0000 979.5000 ;
	    RECT 1518.6000 979.2000 1519.8000 979.5000 ;
	    RECT 1439.4000 977.4000 1440.6000 977.5500 ;
	    RECT 1461.0000 977.4000 1462.2001 977.5500 ;
	    RECT 1463.1000 977.4000 1464.6000 978.3000 ;
	    RECT 1467.0000 976.8000 1467.3000 978.3000 ;
	    RECT 1468.2001 977.4000 1469.4000 978.6000 ;
	    RECT 1489.8000 977.4000 1491.0000 978.6000 ;
	    RECT 1516.2001 977.4000 1517.4000 978.6000 ;
	    RECT 1521.0000 978.3000 1521.9000 983.7000 ;
	    RECT 1523.4000 983.4000 1524.6000 984.6000 ;
	    RECT 1542.6000 983.7000 1543.8000 989.7000 ;
	    RECT 1546.5000 984.6000 1547.7001 989.7000 ;
	    RECT 1545.0000 983.7000 1547.7001 984.6000 ;
	    RECT 1542.6000 982.5000 1543.8000 982.8000 ;
	    RECT 1542.6000 980.4000 1543.8000 981.6000 ;
	    RECT 1545.0000 979.5000 1546.2001 983.7000 ;
	    RECT 1518.3000 976.8000 1518.6000 978.3000 ;
	    RECT 1521.0000 977.4000 1522.5000 978.3000 ;
	    RECT 1523.4000 977.4000 1524.6000 978.6000 ;
	    RECT 1545.0000 978.4500 1546.2001 978.6000 ;
	    RECT 1561.8000 978.4500 1563.0000 978.6000 ;
	    RECT 1545.0000 977.5500 1563.0000 978.4500 ;
	    RECT 1545.0000 977.4000 1546.2001 977.5500 ;
	    RECT 1561.8000 977.4000 1563.0000 977.5500 ;
	    RECT 1413.0000 976.5000 1414.2001 976.8000 ;
	    RECT 1377.0000 963.3000 1378.2001 969.3000 ;
	    RECT 1379.4000 963.3000 1380.6000 976.5000 ;
	    RECT 1381.8000 975.4500 1383.0000 975.6000 ;
	    RECT 1386.6000 975.4500 1387.8000 975.6000 ;
	    RECT 1381.8000 974.5500 1387.8000 975.4500 ;
	    RECT 1381.8000 974.4000 1383.0000 974.5500 ;
	    RECT 1386.6000 974.4000 1387.8000 974.5500 ;
	    RECT 1393.8000 975.4500 1395.0000 975.6000 ;
	    RECT 1405.8000 975.4500 1407.0000 975.6000 ;
	    RECT 1393.8000 974.5500 1407.0000 975.4500 ;
	    RECT 1393.8000 974.4000 1395.0000 974.5500 ;
	    RECT 1405.8000 974.4000 1407.0000 974.5500 ;
	    RECT 1413.0000 975.4500 1414.2001 975.6000 ;
	    RECT 1432.2001 975.4500 1433.4000 975.6000 ;
	    RECT 1413.0000 974.5500 1433.4000 975.4500 ;
	    RECT 1413.0000 974.4000 1414.2001 974.5500 ;
	    RECT 1432.2001 974.4000 1433.4000 974.5500 ;
	    RECT 1408.2001 973.5000 1409.4000 973.8000 ;
	    RECT 1381.8000 973.2000 1383.0000 973.5000 ;
	    RECT 1406.1000 970.5000 1407.0000 973.5000 ;
	    RECT 1432.2001 973.2000 1433.4000 973.5000 ;
	    RECT 1408.2001 971.4000 1409.4000 972.6000 ;
	    RECT 1406.1000 969.6000 1411.5000 970.5000 ;
	    RECT 1406.1000 969.3000 1407.0000 969.6000 ;
	    RECT 1381.8000 963.3000 1383.0000 969.3000 ;
	    RECT 1405.8000 963.3000 1407.0000 969.3000 ;
	    RECT 1410.6000 969.3000 1411.5000 969.6000 ;
	    RECT 1408.2001 963.3000 1409.4000 968.7000 ;
	    RECT 1410.6000 963.3000 1411.8000 969.3000 ;
	    RECT 1413.0000 963.3000 1414.2001 969.3000 ;
	    RECT 1432.2001 963.3000 1433.4000 969.3000 ;
	    RECT 1434.6000 963.3000 1435.8000 976.5000 ;
	    RECT 1461.3000 975.3000 1462.2001 976.5000 ;
	    RECT 1437.0000 963.3000 1438.2001 969.3000 ;
	    RECT 1461.0000 963.3000 1462.2001 975.3000 ;
	    RECT 1463.4000 974.4000 1469.4000 975.3000 ;
	    RECT 1463.4000 963.3000 1464.6000 974.4000 ;
	    RECT 1465.8000 963.3000 1467.0000 973.5000 ;
	    RECT 1468.2001 963.3000 1469.4000 974.4000 ;
	    RECT 1487.4000 963.3000 1488.6000 969.3000 ;
	    RECT 1489.8000 963.3000 1491.0000 976.5000 ;
	    RECT 1492.2001 974.4000 1493.4000 975.6000 ;
	    RECT 1523.4000 975.3000 1524.3000 976.5000 ;
	    RECT 1516.2001 974.4000 1522.2001 975.3000 ;
	    RECT 1492.2001 973.2000 1493.4000 973.5000 ;
	    RECT 1492.2001 963.3000 1493.4000 969.3000 ;
	    RECT 1516.2001 963.3000 1517.4000 974.4000 ;
	    RECT 1518.6000 963.3000 1519.8000 973.5000 ;
	    RECT 1521.0000 963.3000 1522.2001 974.4000 ;
	    RECT 1523.4000 963.3000 1524.6000 975.3000 ;
	    RECT 1535.4000 972.4500 1536.6000 972.6000 ;
	    RECT 1542.6000 972.4500 1543.8000 972.6000 ;
	    RECT 1535.4000 971.5500 1543.8000 972.4500 ;
	    RECT 1535.4000 971.4000 1536.6000 971.5500 ;
	    RECT 1542.6000 971.4000 1543.8000 971.5500 ;
	    RECT 1542.6000 963.3000 1543.8000 969.3000 ;
	    RECT 1545.0000 963.3000 1546.2001 976.5000 ;
	    RECT 1547.4000 974.4000 1548.6000 975.6000 ;
	    RECT 1547.4000 973.2000 1548.6000 973.5000 ;
	    RECT 1547.4000 963.3000 1548.6000 969.3000 ;
	    RECT 1.2000 960.6000 1569.0000 962.4000 ;
	    RECT 25.8000 947.7000 27.0000 959.7000 ;
	    RECT 29.7000 948.6000 30.9000 959.7000 ;
	    RECT 32.1000 953.7000 33.3000 959.7000 ;
	    RECT 31.8000 950.4000 33.0000 951.6000 ;
	    RECT 32.1000 949.5000 33.0000 950.4000 ;
	    RECT 29.7000 947.7000 31.2000 948.6000 ;
	    RECT 18.6000 945.4500 19.8000 945.6000 ;
	    RECT 25.8000 945.4500 27.0000 945.6000 ;
	    RECT 18.6000 944.5500 27.0000 945.4500 ;
	    RECT 18.6000 944.4000 19.8000 944.5500 ;
	    RECT 25.8000 944.4000 27.0000 944.5500 ;
	    RECT 28.2000 944.4000 29.4000 945.6000 ;
	    RECT 28.2000 943.2000 29.4000 943.5000 ;
	    RECT 30.3000 942.6000 31.2000 947.7000 ;
	    RECT 33.0000 947.4000 34.2000 948.6000 ;
	    RECT 45.0000 943.5000 46.2000 959.7000 ;
	    RECT 47.4000 953.7000 48.6000 959.7000 ;
	    RECT 66.6000 953.7000 67.8000 959.7000 ;
	    RECT 66.6000 949.5000 67.8000 949.8000 ;
	    RECT 66.6000 947.4000 67.8000 948.6000 ;
	    RECT 69.0000 946.5000 70.2000 959.7000 ;
	    RECT 71.4000 953.7000 72.6000 959.7000 ;
	    RECT 96.3000 953.7000 97.5000 959.7000 ;
	    RECT 96.6000 950.4000 97.8000 951.6000 ;
	    RECT 96.6000 949.5000 97.5000 950.4000 ;
	    RECT 98.7000 948.6000 99.9000 959.7000 ;
	    RECT 95.4000 947.4000 96.6000 948.6000 ;
	    RECT 98.4000 947.7000 99.9000 948.6000 ;
	    RECT 102.6000 947.7000 103.8000 959.7000 ;
	    RECT 69.0000 945.4500 70.2000 945.6000 ;
	    RECT 95.5500 945.4500 96.4500 947.4000 ;
	    RECT 69.0000 944.5500 96.4500 945.4500 ;
	    RECT 69.0000 944.4000 70.2000 944.5500 ;
	    RECT 25.8000 941.4000 27.0000 942.6000 ;
	    RECT 27.9000 940.8000 28.2000 942.3000 ;
	    RECT 30.3000 941.4000 32.1000 942.6000 ;
	    RECT 33.0000 942.4500 34.2000 942.6000 ;
	    RECT 35.4000 942.4500 36.6000 942.6000 ;
	    RECT 33.0000 941.5500 36.6000 942.4500 ;
	    RECT 33.0000 941.4000 34.2000 941.5500 ;
	    RECT 35.4000 941.4000 36.6000 941.5500 ;
	    RECT 37.8000 942.4500 39.0000 942.6000 ;
	    RECT 45.0000 942.4500 46.2000 942.6000 ;
	    RECT 37.8000 941.5500 46.2000 942.4500 ;
	    RECT 37.8000 941.4000 39.0000 941.5500 ;
	    RECT 45.0000 941.4000 46.2000 941.5500 ;
	    RECT 26.1000 939.3000 31.5000 939.9000 ;
	    RECT 33.0000 939.3000 33.9000 940.5000 ;
	    RECT 25.8000 939.0000 31.8000 939.3000 ;
	    RECT 25.8000 933.3000 27.0000 939.0000 ;
	    RECT 28.2000 933.3000 29.4000 938.1000 ;
	    RECT 30.6000 933.3000 31.8000 939.0000 ;
	    RECT 33.0000 933.3000 34.2000 939.3000 ;
	    RECT 45.0000 933.3000 46.2000 940.5000 ;
	    RECT 47.4000 939.4500 48.6000 939.6000 ;
	    RECT 64.2000 939.4500 65.4000 939.6000 ;
	    RECT 47.4000 938.5500 65.4000 939.4500 ;
	    RECT 69.0000 939.3000 70.2000 943.5000 ;
	    RECT 98.4000 942.6000 99.3000 947.7000 ;
	    RECT 100.2000 945.4500 101.4000 945.6000 ;
	    RECT 100.2000 944.5500 106.0500 945.4500 ;
	    RECT 100.2000 944.4000 101.4000 944.5500 ;
	    RECT 100.2000 943.2000 101.4000 943.5000 ;
	    RECT 71.4000 941.4000 72.6000 942.6000 ;
	    RECT 95.4000 941.4000 96.6000 942.6000 ;
	    RECT 97.5000 941.4000 99.3000 942.6000 ;
	    RECT 101.4000 940.8000 101.7000 942.3000 ;
	    RECT 102.6000 941.4000 103.8000 942.6000 ;
	    RECT 105.1500 942.4500 106.0500 944.5500 ;
	    RECT 117.0000 943.5000 118.2000 959.7000 ;
	    RECT 119.4000 953.7000 120.6000 959.7000 ;
	    RECT 133.8000 953.7000 135.0000 959.7000 ;
	    RECT 136.2000 943.5000 137.4000 959.7000 ;
	    RECT 155.4000 953.7000 156.6000 959.7000 ;
	    RECT 155.4000 949.5000 156.6000 949.8000 ;
	    RECT 153.0000 948.4500 154.2000 948.6000 ;
	    RECT 155.4000 948.4500 156.6000 948.6000 ;
	    RECT 153.0000 947.5500 156.6000 948.4500 ;
	    RECT 153.0000 947.4000 154.2000 947.5500 ;
	    RECT 155.4000 947.4000 156.6000 947.5500 ;
	    RECT 157.8000 946.5000 159.0000 959.7000 ;
	    RECT 160.2000 953.7000 161.4000 959.7000 ;
	    RECT 179.4000 954.4500 180.6000 954.6000 ;
	    RECT 184.2000 954.4500 185.4000 954.6000 ;
	    RECT 179.4000 953.5500 185.4000 954.4500 ;
	    RECT 179.4000 953.4000 180.6000 953.5500 ;
	    RECT 184.2000 953.4000 185.4000 953.5500 ;
	    RECT 191.4000 947.7000 192.6000 959.7000 ;
	    RECT 195.3000 947.7000 198.3000 959.7000 ;
	    RECT 201.0000 947.7000 202.2000 959.7000 ;
	    RECT 157.8000 944.4000 159.0000 945.6000 ;
	    RECT 179.4000 945.4500 180.6000 945.6000 ;
	    RECT 191.4000 945.4500 192.6000 945.6000 ;
	    RECT 193.8000 945.4500 195.0000 945.6000 ;
	    RECT 179.4000 944.5500 195.0000 945.4500 ;
	    RECT 179.4000 944.4000 180.6000 944.5500 ;
	    RECT 191.4000 944.4000 192.6000 944.5500 ;
	    RECT 193.8000 944.4000 195.0000 944.5500 ;
	    RECT 196.2000 943.5000 197.1000 947.7000 ;
	    RECT 198.6000 944.4000 199.8000 945.6000 ;
	    RECT 201.0000 943.5000 202.2000 943.8000 ;
	    RECT 220.2000 943.5000 221.4000 959.7000 ;
	    RECT 222.6000 953.7000 223.8000 959.7000 ;
	    RECT 249.0000 953.7000 250.2000 959.7000 ;
	    RECT 251.4000 954.3000 252.6000 959.7000 ;
	    RECT 249.3000 953.4000 250.2000 953.7000 ;
	    RECT 253.8000 953.7000 255.0000 959.7000 ;
	    RECT 256.2000 953.7000 257.4000 959.7000 ;
	    RECT 280.2000 953.7000 281.4000 959.7000 ;
	    RECT 282.6000 953.7000 283.8000 959.7000 ;
	    RECT 285.0000 954.3000 286.2000 959.7000 ;
	    RECT 253.8000 953.4000 254.7000 953.7000 ;
	    RECT 249.3000 952.5000 254.7000 953.4000 ;
	    RECT 282.9000 953.4000 283.8000 953.7000 ;
	    RECT 287.4000 953.7000 288.6000 959.7000 ;
	    RECT 313.8000 953.7000 315.0000 959.7000 ;
	    RECT 316.2000 954.3000 317.4000 959.7000 ;
	    RECT 287.4000 953.4000 288.3000 953.7000 ;
	    RECT 282.9000 952.5000 288.3000 953.4000 ;
	    RECT 249.3000 949.5000 250.2000 952.5000 ;
	    RECT 251.4000 951.4500 252.6000 951.6000 ;
	    RECT 275.4000 951.4500 276.6000 951.6000 ;
	    RECT 251.4000 950.5500 276.6000 951.4500 ;
	    RECT 251.4000 950.4000 252.6000 950.5500 ;
	    RECT 275.4000 950.4000 276.6000 950.5500 ;
	    RECT 285.0000 950.4000 286.2000 951.6000 ;
	    RECT 287.4000 949.5000 288.3000 952.5000 ;
	    RECT 314.1000 953.4000 315.0000 953.7000 ;
	    RECT 318.6000 953.7000 319.8000 959.7000 ;
	    RECT 321.0000 953.7000 322.2000 959.7000 ;
	    RECT 345.0000 953.7000 346.2000 959.7000 ;
	    RECT 347.4000 953.7000 348.6000 959.7000 ;
	    RECT 349.8000 954.3000 351.0000 959.7000 ;
	    RECT 318.6000 953.4000 319.5000 953.7000 ;
	    RECT 314.1000 952.5000 319.5000 953.4000 ;
	    RECT 347.7000 953.4000 348.6000 953.7000 ;
	    RECT 352.2000 953.7000 353.4000 959.7000 ;
	    RECT 376.2000 953.7000 377.4000 959.7000 ;
	    RECT 378.6000 954.3000 379.8000 959.7000 ;
	    RECT 352.2000 953.4000 353.1000 953.7000 ;
	    RECT 347.7000 952.5000 353.1000 953.4000 ;
	    RECT 314.1000 949.5000 315.0000 952.5000 ;
	    RECT 316.2000 950.4000 317.4000 951.6000 ;
	    RECT 318.6000 951.4500 319.8000 951.6000 ;
	    RECT 328.2000 951.4500 329.4000 951.6000 ;
	    RECT 349.8000 951.4500 351.0000 951.6000 ;
	    RECT 318.6000 950.5500 324.4500 951.4500 ;
	    RECT 318.6000 950.4000 319.8000 950.5500 ;
	    RECT 251.4000 949.2000 252.6000 949.5000 ;
	    RECT 285.0000 949.2000 286.2000 949.5000 ;
	    RECT 316.2000 949.2000 317.4000 949.5000 ;
	    RECT 249.0000 947.4000 250.2000 948.6000 ;
	    RECT 256.2000 948.4500 257.4000 948.6000 ;
	    RECT 280.2000 948.4500 281.4000 948.6000 ;
	    RECT 256.2000 947.5500 281.4000 948.4500 ;
	    RECT 256.2000 947.4000 257.4000 947.5500 ;
	    RECT 280.2000 947.4000 281.4000 947.5500 ;
	    RECT 287.4000 948.4500 288.6000 948.6000 ;
	    RECT 309.0000 948.4500 310.2000 948.6000 ;
	    RECT 287.4000 947.5500 310.2000 948.4500 ;
	    RECT 287.4000 947.4000 288.6000 947.5500 ;
	    RECT 309.0000 947.4000 310.2000 947.5500 ;
	    RECT 311.4000 948.4500 312.6000 948.6000 ;
	    RECT 313.8000 948.4500 315.0000 948.6000 ;
	    RECT 311.4000 947.5500 315.0000 948.4500 ;
	    RECT 311.4000 947.4000 312.6000 947.5500 ;
	    RECT 313.8000 947.4000 315.0000 947.5500 ;
	    RECT 321.0000 947.4000 322.2000 948.6000 ;
	    RECT 323.5500 948.4500 324.4500 950.5500 ;
	    RECT 328.2000 950.5500 351.0000 951.4500 ;
	    RECT 328.2000 950.4000 329.4000 950.5500 ;
	    RECT 349.8000 950.4000 351.0000 950.5500 ;
	    RECT 352.2000 949.5000 353.1000 952.5000 ;
	    RECT 376.5000 953.4000 377.4000 953.7000 ;
	    RECT 381.0000 953.7000 382.2000 959.7000 ;
	    RECT 383.4000 953.7000 384.6000 959.7000 ;
	    RECT 407.4000 953.7000 408.6000 959.7000 ;
	    RECT 409.8000 954.3000 411.0000 959.7000 ;
	    RECT 381.0000 953.4000 381.9000 953.7000 ;
	    RECT 376.5000 952.5000 381.9000 953.4000 ;
	    RECT 407.7000 953.4000 408.6000 953.7000 ;
	    RECT 412.2000 953.7000 413.4000 959.7000 ;
	    RECT 414.6000 953.7000 415.8000 959.7000 ;
	    RECT 449.1000 953.7000 450.3000 959.7000 ;
	    RECT 412.2000 953.4000 413.1000 953.7000 ;
	    RECT 407.7000 952.5000 413.1000 953.4000 ;
	    RECT 376.5000 949.5000 377.4000 952.5000 ;
	    RECT 378.6000 950.4000 379.8000 951.6000 ;
	    RECT 407.7000 949.5000 408.6000 952.5000 ;
	    RECT 409.8000 950.4000 411.0000 951.6000 ;
	    RECT 417.0000 951.4500 418.2000 951.6000 ;
	    RECT 412.3500 950.5500 418.2000 951.4500 ;
	    RECT 349.8000 949.2000 351.0000 949.5000 ;
	    RECT 378.6000 949.2000 379.8000 949.5000 ;
	    RECT 409.8000 949.2000 411.0000 949.5000 ;
	    RECT 342.6000 948.4500 343.8000 948.6000 ;
	    RECT 345.0000 948.4500 346.2000 948.6000 ;
	    RECT 323.5500 947.5500 346.2000 948.4500 ;
	    RECT 342.6000 947.4000 343.8000 947.5500 ;
	    RECT 345.0000 947.4000 346.2000 947.5500 ;
	    RECT 352.2000 948.4500 353.4000 948.6000 ;
	    RECT 357.0000 948.4500 358.2000 948.6000 ;
	    RECT 376.2000 948.4500 377.4000 948.6000 ;
	    RECT 352.2000 947.5500 355.6500 948.4500 ;
	    RECT 352.2000 947.4000 353.4000 947.5500 ;
	    RECT 117.0000 942.4500 118.2000 942.6000 ;
	    RECT 105.1500 941.5500 118.2000 942.4500 ;
	    RECT 117.0000 941.4000 118.2000 941.5500 ;
	    RECT 136.2000 942.4500 137.4000 942.6000 ;
	    RECT 138.6000 942.4500 139.8000 942.6000 ;
	    RECT 136.2000 941.5500 139.8000 942.4500 ;
	    RECT 136.2000 941.4000 137.4000 941.5500 ;
	    RECT 138.6000 941.4000 139.8000 941.5500 ;
	    RECT 71.4000 940.2000 72.6000 940.5000 ;
	    RECT 95.7000 939.3000 96.6000 940.5000 ;
	    RECT 98.1000 939.3000 103.5000 939.9000 ;
	    RECT 47.4000 938.4000 48.6000 938.5500 ;
	    RECT 64.2000 938.4000 65.4000 938.5500 ;
	    RECT 67.5000 938.4000 70.2000 939.3000 ;
	    RECT 47.4000 937.2000 48.6000 937.5000 ;
	    RECT 47.4000 933.3000 48.6000 936.3000 ;
	    RECT 67.5000 933.3000 68.7000 938.4000 ;
	    RECT 71.4000 933.3000 72.6000 939.3000 ;
	    RECT 95.4000 933.3000 96.6000 939.3000 ;
	    RECT 97.8000 939.0000 103.8000 939.3000 ;
	    RECT 97.8000 933.3000 99.0000 939.0000 ;
	    RECT 100.2000 933.3000 101.4000 938.1000 ;
	    RECT 102.6000 933.3000 103.8000 939.0000 ;
	    RECT 117.0000 933.3000 118.2000 940.5000 ;
	    RECT 119.4000 939.4500 120.6000 939.6000 ;
	    RECT 131.4000 939.4500 132.6000 939.6000 ;
	    RECT 119.4000 938.5500 132.6000 939.4500 ;
	    RECT 119.4000 938.4000 120.6000 938.5500 ;
	    RECT 131.4000 938.4000 132.6000 938.5500 ;
	    RECT 133.8000 938.4000 135.0000 939.6000 ;
	    RECT 119.4000 937.2000 120.6000 937.5000 ;
	    RECT 133.8000 937.2000 135.0000 937.5000 ;
	    RECT 119.4000 933.3000 120.6000 936.3000 ;
	    RECT 133.8000 933.3000 135.0000 936.3000 ;
	    RECT 136.2000 933.3000 137.4000 940.5000 ;
	    RECT 157.8000 939.3000 159.0000 943.5000 ;
	    RECT 193.8000 943.2000 195.0000 943.5000 ;
	    RECT 198.6000 943.2000 199.8000 943.5000 ;
	    RECT 249.3000 942.6000 250.2000 946.5000 ;
	    RECT 256.2000 946.2000 257.4000 946.5000 ;
	    RECT 280.2000 946.2000 281.4000 946.5000 ;
	    RECT 252.6000 944.4000 252.9000 945.6000 ;
	    RECT 253.8000 944.4000 255.0000 945.6000 ;
	    RECT 282.6000 944.4000 283.8000 945.6000 ;
	    RECT 284.7000 944.4000 285.0000 945.6000 ;
	    RECT 287.4000 942.6000 288.3000 946.5000 ;
	    RECT 160.2000 942.4500 161.4000 942.6000 ;
	    RECT 162.6000 942.4500 163.8000 942.6000 ;
	    RECT 174.6000 942.4500 175.8000 942.6000 ;
	    RECT 160.2000 941.5500 175.8000 942.4500 ;
	    RECT 160.2000 941.4000 161.4000 941.5500 ;
	    RECT 162.6000 941.4000 163.8000 941.5500 ;
	    RECT 174.6000 941.4000 175.8000 941.5500 ;
	    RECT 191.4000 941.4000 192.6000 942.6000 ;
	    RECT 193.5000 940.8000 193.8000 942.3000 ;
	    RECT 196.2000 941.4000 197.4000 942.6000 ;
	    RECT 201.0000 942.4500 202.2000 942.6000 ;
	    RECT 220.2000 942.4500 221.4000 942.6000 ;
	    RECT 198.3000 941.4000 199.8000 942.3000 ;
	    RECT 201.0000 941.5500 221.4000 942.4500 ;
	    RECT 249.3000 942.3000 251.7000 942.6000 ;
	    RECT 285.9000 942.3000 288.3000 942.6000 ;
	    RECT 249.3000 941.7000 252.0000 942.3000 ;
	    RECT 201.0000 941.4000 202.2000 941.5500 ;
	    RECT 220.2000 941.4000 221.4000 941.5500 ;
	    RECT 160.2000 940.2000 161.4000 940.5000 ;
	    RECT 162.6000 939.4500 163.8000 939.6000 ;
	    RECT 169.8000 939.4500 171.0000 939.6000 ;
	    RECT 156.3000 938.4000 159.0000 939.3000 ;
	    RECT 156.3000 933.3000 157.5000 938.4000 ;
	    RECT 160.2000 933.3000 161.4000 939.3000 ;
	    RECT 162.6000 938.5500 171.0000 939.4500 ;
	    RECT 191.7000 939.3000 197.1000 939.9000 ;
	    RECT 198.9000 939.3000 199.8000 941.4000 ;
	    RECT 162.6000 938.4000 163.8000 938.5500 ;
	    RECT 169.8000 938.4000 171.0000 938.5500 ;
	    RECT 191.4000 939.0000 197.4000 939.3000 ;
	    RECT 191.4000 933.3000 192.6000 939.0000 ;
	    RECT 193.8000 933.3000 195.0000 938.1000 ;
	    RECT 196.2000 934.2000 197.4000 939.0000 ;
	    RECT 198.6000 935.1000 199.8000 939.3000 ;
	    RECT 201.0000 934.2000 202.2000 939.3000 ;
	    RECT 196.2000 933.3000 202.2000 934.2000 ;
	    RECT 220.2000 933.3000 221.4000 940.5000 ;
	    RECT 222.6000 939.4500 223.8000 939.6000 ;
	    RECT 244.2000 939.4500 245.4000 939.6000 ;
	    RECT 222.6000 938.5500 245.4000 939.4500 ;
	    RECT 222.6000 938.4000 223.8000 938.5500 ;
	    RECT 244.2000 938.4000 245.4000 938.5500 ;
	    RECT 222.6000 937.2000 223.8000 937.5000 ;
	    RECT 222.6000 933.3000 223.8000 936.3000 ;
	    RECT 250.8000 933.3000 252.0000 941.7000 ;
	    RECT 256.2000 933.3000 257.4000 942.3000 ;
	    RECT 280.2000 933.3000 281.4000 942.3000 ;
	    RECT 285.6000 941.7000 288.3000 942.3000 ;
	    RECT 314.1000 942.6000 315.0000 946.5000 ;
	    RECT 321.0000 946.2000 322.2000 946.5000 ;
	    RECT 345.0000 946.2000 346.2000 946.5000 ;
	    RECT 317.4000 944.4000 317.7000 945.6000 ;
	    RECT 318.6000 944.4000 319.8000 945.6000 ;
	    RECT 347.4000 944.4000 348.6000 945.6000 ;
	    RECT 349.5000 944.4000 349.8000 945.6000 ;
	    RECT 352.2000 942.6000 353.1000 946.5000 ;
	    RECT 354.7500 945.4500 355.6500 947.5500 ;
	    RECT 357.0000 947.5500 377.4000 948.4500 ;
	    RECT 357.0000 947.4000 358.2000 947.5500 ;
	    RECT 376.2000 947.4000 377.4000 947.5500 ;
	    RECT 383.4000 948.4500 384.6000 948.6000 ;
	    RECT 385.8000 948.4500 387.0000 948.6000 ;
	    RECT 383.4000 947.5500 387.0000 948.4500 ;
	    RECT 383.4000 947.4000 384.6000 947.5500 ;
	    RECT 385.8000 947.4000 387.0000 947.5500 ;
	    RECT 390.6000 948.4500 391.8000 948.6000 ;
	    RECT 407.4000 948.4500 408.6000 948.6000 ;
	    RECT 390.6000 947.5500 408.6000 948.4500 ;
	    RECT 390.6000 947.4000 391.8000 947.5500 ;
	    RECT 407.4000 947.4000 408.6000 947.5500 ;
	    RECT 373.8000 945.4500 375.0000 945.6000 ;
	    RECT 354.7500 944.5500 375.0000 945.4500 ;
	    RECT 373.8000 944.4000 375.0000 944.5500 ;
	    RECT 314.1000 942.3000 316.5000 942.6000 ;
	    RECT 350.7000 942.3000 353.1000 942.6000 ;
	    RECT 314.1000 941.7000 316.8000 942.3000 ;
	    RECT 285.6000 933.3000 286.8000 941.7000 ;
	    RECT 315.6000 933.3000 316.8000 941.7000 ;
	    RECT 321.0000 933.3000 322.2000 942.3000 ;
	    RECT 345.0000 933.3000 346.2000 942.3000 ;
	    RECT 350.4000 941.7000 353.1000 942.3000 ;
	    RECT 376.5000 942.6000 377.4000 946.5000 ;
	    RECT 383.4000 946.2000 384.6000 946.5000 ;
	    RECT 379.8000 944.4000 380.1000 945.6000 ;
	    RECT 381.0000 944.4000 382.2000 945.6000 ;
	    RECT 407.7000 942.6000 408.6000 946.5000 ;
	    RECT 412.3500 945.6000 413.2500 950.5500 ;
	    RECT 417.0000 950.4000 418.2000 950.5500 ;
	    RECT 449.4000 950.4000 450.6000 951.6000 ;
	    RECT 449.4000 949.5000 450.3000 950.4000 ;
	    RECT 451.5000 948.6000 452.7000 959.7000 ;
	    RECT 414.6000 948.4500 415.8000 948.6000 ;
	    RECT 424.2000 948.4500 425.4000 948.6000 ;
	    RECT 414.6000 947.5500 425.4000 948.4500 ;
	    RECT 414.6000 947.4000 415.8000 947.5500 ;
	    RECT 424.2000 947.4000 425.4000 947.5500 ;
	    RECT 433.8000 948.4500 435.0000 948.6000 ;
	    RECT 448.2000 948.4500 449.4000 948.6000 ;
	    RECT 433.8000 947.5500 449.4000 948.4500 ;
	    RECT 433.8000 947.4000 435.0000 947.5500 ;
	    RECT 448.2000 947.4000 449.4000 947.5500 ;
	    RECT 451.2000 947.7000 452.7000 948.6000 ;
	    RECT 455.4000 947.7000 456.6000 959.7000 ;
	    RECT 414.6000 946.2000 415.8000 946.5000 ;
	    RECT 411.0000 944.4000 411.3000 945.6000 ;
	    RECT 412.2000 944.4000 413.4000 945.6000 ;
	    RECT 451.2000 942.6000 452.1000 947.7000 ;
	    RECT 453.0000 944.4000 454.2000 945.6000 ;
	    RECT 469.8000 943.5000 471.0000 959.7000 ;
	    RECT 472.2000 953.7000 473.4000 959.7000 ;
	    RECT 525.0000 959.4000 526.2000 960.6000 ;
	    RECT 597.0000 953.7000 598.2000 959.7000 ;
	    RECT 599.4000 954.6000 600.6000 959.7000 ;
	    RECT 599.1000 953.7000 600.6000 954.6000 ;
	    RECT 601.8000 953.7000 603.0000 960.6000 ;
	    RECT 599.1000 952.8000 600.0000 953.7000 ;
	    RECT 604.2000 952.8000 605.4000 959.7000 ;
	    RECT 606.6000 953.7000 607.8000 959.7000 ;
	    RECT 609.0000 955.5000 610.2000 959.7000 ;
	    RECT 611.4000 955.5000 612.6000 959.7000 ;
	    RECT 597.0000 951.9000 600.0000 952.8000 ;
	    RECT 597.0000 943.5000 598.2000 951.9000 ;
	    RECT 600.9000 951.6000 607.2000 952.8000 ;
	    RECT 613.8000 952.5000 615.0000 959.7000 ;
	    RECT 616.2000 953.7000 617.4000 959.7000 ;
	    RECT 618.6000 952.5000 619.8000 959.7000 ;
	    RECT 621.0000 953.7000 622.2000 959.7000 ;
	    RECT 600.9000 951.0000 601.8000 951.6000 ;
	    RECT 599.4000 949.8000 601.8000 951.0000 ;
	    RECT 606.3000 950.7000 615.0000 951.6000 ;
	    RECT 603.3000 949.8000 605.4000 950.7000 ;
	    RECT 603.3000 949.5000 612.6000 949.8000 ;
	    RECT 604.5000 948.9000 612.6000 949.5000 ;
	    RECT 611.4000 948.6000 612.6000 948.9000 ;
	    RECT 614.1000 949.5000 615.0000 950.7000 ;
	    RECT 615.9000 950.4000 619.8000 951.6000 ;
	    RECT 623.4000 950.4000 624.6000 959.7000 ;
	    RECT 625.8000 955.5000 627.0000 959.7000 ;
	    RECT 628.2000 955.5000 629.4000 959.7000 ;
	    RECT 630.6000 955.5000 631.8000 959.7000 ;
	    RECT 633.0000 953.7000 634.2000 959.7000 ;
	    RECT 628.2000 951.6000 634.5000 952.8000 ;
	    RECT 635.4000 951.6000 636.6000 959.7000 ;
	    RECT 637.8000 953.7000 639.0000 959.7000 ;
	    RECT 640.2000 952.8000 641.4000 959.7000 ;
	    RECT 642.6000 953.7000 643.8000 959.7000 ;
	    RECT 640.2000 951.9000 644.1000 952.8000 ;
	    RECT 645.0000 952.5000 646.2000 959.7000 ;
	    RECT 647.4000 953.7000 648.6000 959.7000 ;
	    RECT 678.6000 953.7000 679.8000 959.7000 ;
	    RECT 681.0000 953.7000 682.2000 959.7000 ;
	    RECT 635.4000 950.4000 639.3000 951.6000 ;
	    RECT 625.8000 949.5000 627.0000 949.8000 ;
	    RECT 614.1000 948.6000 627.0000 949.5000 ;
	    RECT 630.6000 949.5000 631.8000 949.8000 ;
	    RECT 643.2000 949.5000 644.1000 951.9000 ;
	    RECT 645.0000 950.4000 646.2000 951.6000 ;
	    RECT 630.6000 948.6000 644.1000 949.5000 ;
	    RECT 601.8000 947.4000 603.0000 948.6000 ;
	    RECT 606.9000 947.7000 608.1000 948.0000 ;
	    RECT 603.9000 946.8000 642.3000 947.7000 ;
	    RECT 641.1000 946.5000 642.3000 946.8000 ;
	    RECT 643.2000 945.9000 644.1000 948.6000 ;
	    RECT 645.0000 948.0000 646.2000 949.5000 ;
	    RECT 645.0000 946.8000 646.5000 948.0000 ;
	    RECT 599.1000 945.0000 605.7000 945.9000 ;
	    RECT 599.1000 944.7000 600.3000 945.0000 ;
	    RECT 606.6000 944.4000 607.8000 945.6000 ;
	    RECT 608.7000 945.0000 634.2000 945.9000 ;
	    RECT 643.2000 945.0000 644.4000 945.9000 ;
	    RECT 633.0000 944.1000 634.2000 945.0000 ;
	    RECT 453.0000 943.2000 454.2000 943.5000 ;
	    RECT 376.5000 942.3000 378.9000 942.6000 ;
	    RECT 407.7000 942.3000 410.1000 942.6000 ;
	    RECT 417.0000 942.4500 418.2000 942.6000 ;
	    RECT 448.2000 942.4500 449.4000 942.6000 ;
	    RECT 376.5000 941.7000 379.2000 942.3000 ;
	    RECT 350.4000 933.3000 351.6000 941.7000 ;
	    RECT 354.6000 939.4500 355.8000 939.6000 ;
	    RECT 361.8000 939.4500 363.0000 939.6000 ;
	    RECT 354.6000 938.5500 363.0000 939.4500 ;
	    RECT 354.6000 938.4000 355.8000 938.5500 ;
	    RECT 361.8000 938.4000 363.0000 938.5500 ;
	    RECT 378.0000 933.3000 379.2000 941.7000 ;
	    RECT 383.4000 933.3000 384.6000 942.3000 ;
	    RECT 407.7000 941.7000 410.4000 942.3000 ;
	    RECT 409.2000 933.3000 410.4000 941.7000 ;
	    RECT 414.6000 933.3000 415.8000 942.3000 ;
	    RECT 417.0000 941.5500 449.4000 942.4500 ;
	    RECT 417.0000 941.4000 418.2000 941.5500 ;
	    RECT 448.2000 941.4000 449.4000 941.5500 ;
	    RECT 450.3000 941.4000 452.1000 942.6000 ;
	    RECT 454.2000 940.8000 454.5000 942.3000 ;
	    RECT 455.4000 941.4000 456.6000 942.6000 ;
	    RECT 460.2000 942.4500 461.4000 942.6000 ;
	    RECT 469.8000 942.4500 471.0000 942.6000 ;
	    RECT 460.2000 941.5500 471.0000 942.4500 ;
	    RECT 460.2000 941.4000 461.4000 941.5500 ;
	    RECT 469.8000 941.4000 471.0000 941.5500 ;
	    RECT 597.0000 942.3000 610.2000 943.5000 ;
	    RECT 611.1000 942.9000 614.1000 944.1000 ;
	    RECT 619.8000 942.9000 624.6000 944.1000 ;
	    RECT 448.5000 939.3000 449.4000 940.5000 ;
	    RECT 450.9000 939.3000 456.3000 939.9000 ;
	    RECT 448.2000 933.3000 449.4000 939.3000 ;
	    RECT 450.6000 939.0000 456.6000 939.3000 ;
	    RECT 450.6000 933.3000 451.8000 939.0000 ;
	    RECT 453.0000 933.3000 454.2000 938.1000 ;
	    RECT 455.4000 933.3000 456.6000 939.0000 ;
	    RECT 469.8000 933.3000 471.0000 940.5000 ;
	    RECT 472.2000 939.4500 473.4000 939.6000 ;
	    RECT 479.4000 939.4500 480.6000 939.6000 ;
	    RECT 510.6000 939.4500 511.8000 939.6000 ;
	    RECT 472.2000 938.5500 511.8000 939.4500 ;
	    RECT 472.2000 938.4000 473.4000 938.5500 ;
	    RECT 479.4000 938.4000 480.6000 938.5500 ;
	    RECT 510.6000 938.4000 511.8000 938.5500 ;
	    RECT 472.2000 937.2000 473.4000 937.5000 ;
	    RECT 472.2000 933.3000 473.4000 936.3000 ;
	    RECT 597.0000 933.3000 598.2000 942.3000 ;
	    RECT 600.6000 940.2000 605.1000 941.4000 ;
	    RECT 603.9000 939.3000 605.1000 940.2000 ;
	    RECT 612.9000 939.3000 614.1000 942.9000 ;
	    RECT 616.2000 941.4000 617.4000 942.6000 ;
	    RECT 624.0000 941.7000 625.2000 942.0000 ;
	    RECT 618.6000 940.8000 625.2000 941.7000 ;
	    RECT 618.6000 940.5000 619.8000 940.8000 ;
	    RECT 616.2000 940.2000 617.4000 940.5000 ;
	    RECT 628.2000 939.6000 629.4000 943.8000 ;
	    RECT 636.9000 942.9000 642.6000 944.1000 ;
	    RECT 636.9000 941.1000 638.1000 942.9000 ;
	    RECT 643.5000 942.0000 644.4000 945.0000 ;
	    RECT 618.6000 939.3000 619.8000 939.6000 ;
	    RECT 601.8000 933.3000 603.0000 939.3000 ;
	    RECT 603.9000 938.1000 607.8000 939.3000 ;
	    RECT 612.9000 938.4000 619.8000 939.3000 ;
	    RECT 621.0000 938.4000 622.2000 939.6000 ;
	    RECT 623.1000 938.4000 623.4000 939.6000 ;
	    RECT 627.9000 938.4000 629.4000 939.6000 ;
	    RECT 635.4000 940.2000 638.1000 941.1000 ;
	    RECT 642.6000 941.1000 644.4000 942.0000 ;
	    RECT 635.4000 939.3000 636.6000 940.2000 ;
	    RECT 606.6000 933.3000 607.8000 938.1000 ;
	    RECT 633.0000 938.1000 636.6000 939.3000 ;
	    RECT 609.0000 933.3000 610.2000 937.5000 ;
	    RECT 611.4000 933.3000 612.6000 937.5000 ;
	    RECT 613.8000 933.3000 615.0000 937.5000 ;
	    RECT 616.2000 933.3000 617.4000 936.3000 ;
	    RECT 618.6000 933.3000 619.8000 937.5000 ;
	    RECT 621.0000 933.3000 622.2000 936.3000 ;
	    RECT 623.4000 933.3000 624.6000 937.5000 ;
	    RECT 625.8000 933.3000 627.0000 937.5000 ;
	    RECT 628.2000 933.3000 629.4000 937.5000 ;
	    RECT 630.6000 933.3000 631.8000 937.5000 ;
	    RECT 633.0000 933.3000 634.2000 938.1000 ;
	    RECT 637.8000 933.3000 639.0000 939.3000 ;
	    RECT 642.6000 933.3000 643.8000 941.1000 ;
	    RECT 645.3000 940.2000 646.5000 946.8000 ;
	    RECT 681.3000 947.4000 682.2000 953.7000 ;
	    RECT 683.4000 948.3000 684.6000 959.7000 ;
	    RECT 685.8000 947.7000 687.0000 959.7000 ;
	    RECT 709.8000 948.6000 711.0000 959.7000 ;
	    RECT 712.2000 949.5000 713.4000 959.7000 ;
	    RECT 714.6000 948.6000 715.8000 959.7000 ;
	    RECT 709.8000 947.7000 715.8000 948.6000 ;
	    RECT 717.0000 947.7000 718.2000 959.7000 ;
	    RECT 741.0000 947.7000 742.2000 959.7000 ;
	    RECT 744.9000 948.6000 746.1000 959.7000 ;
	    RECT 747.3000 953.7000 748.5000 959.7000 ;
	    RECT 767.4000 953.7000 768.6000 959.7000 ;
	    RECT 747.0000 950.4000 748.2000 951.6000 ;
	    RECT 747.3000 949.5000 748.2000 950.4000 ;
	    RECT 767.4000 949.5000 768.6000 949.8000 ;
	    RECT 744.9000 947.7000 746.4000 948.6000 ;
	    RECT 681.3000 946.5000 684.9000 947.4000 ;
	    RECT 686.1000 946.5000 687.0000 947.7000 ;
	    RECT 717.0000 946.5000 717.9000 947.7000 ;
	    RECT 681.0000 944.4000 682.2000 945.6000 ;
	    RECT 678.6000 943.5000 679.8000 943.8000 ;
	    RECT 681.3000 943.2000 682.2000 943.5000 ;
	    RECT 678.6000 941.4000 679.8000 942.6000 ;
	    RECT 681.3000 942.3000 682.8000 943.2000 ;
	    RECT 681.6000 942.0000 682.8000 942.3000 ;
	    RECT 684.0000 941.4000 684.9000 946.5000 ;
	    RECT 685.8000 945.4500 687.0000 945.6000 ;
	    RECT 688.2000 945.4500 689.4000 945.6000 ;
	    RECT 685.8000 944.5500 689.4000 945.4500 ;
	    RECT 685.8000 944.4000 687.0000 944.5500 ;
	    RECT 688.2000 944.4000 689.4000 944.5500 ;
	    RECT 709.8000 944.4000 711.0000 945.6000 ;
	    RECT 711.9000 944.7000 712.2000 946.2000 ;
	    RECT 714.6000 944.7000 716.1000 945.6000 ;
	    RECT 717.0000 945.4500 718.2000 945.6000 ;
	    RECT 743.4000 945.4500 744.6000 945.6000 ;
	    RECT 712.2000 943.5000 713.4000 943.8000 ;
	    RECT 684.0000 941.1000 685.2000 941.4000 ;
	    RECT 680.7000 940.5000 685.2000 941.1000 ;
	    RECT 645.0000 939.0000 646.5000 940.2000 ;
	    RECT 678.9000 940.2000 685.2000 940.5000 ;
	    RECT 678.9000 939.6000 681.6000 940.2000 ;
	    RECT 678.9000 939.3000 679.8000 939.6000 ;
	    RECT 686.1000 939.3000 687.0000 943.5000 ;
	    RECT 712.2000 941.4000 713.4000 942.6000 ;
	    RECT 714.6000 939.3000 715.5000 944.7000 ;
	    RECT 717.0000 944.5500 744.6000 945.4500 ;
	    RECT 717.0000 944.4000 718.2000 944.5500 ;
	    RECT 743.4000 944.4000 744.6000 944.5500 ;
	    RECT 743.4000 943.2000 744.6000 943.5000 ;
	    RECT 745.5000 942.6000 746.4000 947.7000 ;
	    RECT 748.2000 948.4500 749.4000 948.6000 ;
	    RECT 753.0000 948.4500 754.2000 948.6000 ;
	    RECT 748.2000 947.5500 754.2000 948.4500 ;
	    RECT 748.2000 947.4000 749.4000 947.5500 ;
	    RECT 753.0000 947.4000 754.2000 947.5500 ;
	    RECT 767.4000 947.4000 768.6000 948.6000 ;
	    RECT 769.8000 946.5000 771.0000 959.7000 ;
	    RECT 772.2000 953.7000 773.4000 959.7000 ;
	    RECT 796.2000 947.7000 797.4000 959.7000 ;
	    RECT 800.1000 948.6000 801.3000 959.7000 ;
	    RECT 802.5000 953.7000 803.7000 959.7000 ;
	    RECT 817.8000 959.4000 819.0000 960.6000 ;
	    RECT 830.7000 953.7000 831.9000 959.7000 ;
	    RECT 802.2000 950.4000 803.4000 951.6000 ;
	    RECT 802.5000 949.5000 803.4000 950.4000 ;
	    RECT 831.0000 950.4000 832.2000 951.6000 ;
	    RECT 831.0000 949.5000 831.9000 950.4000 ;
	    RECT 833.1000 948.6000 834.3000 959.7000 ;
	    RECT 800.1000 947.7000 801.6000 948.6000 ;
	    RECT 769.8000 945.4500 771.0000 945.6000 ;
	    RECT 786.6000 945.4500 787.8000 945.6000 ;
	    RECT 769.8000 944.5500 787.8000 945.4500 ;
	    RECT 769.8000 944.4000 771.0000 944.5500 ;
	    RECT 786.6000 944.4000 787.8000 944.5500 ;
	    RECT 791.4000 945.4500 792.6000 945.6000 ;
	    RECT 798.6000 945.4500 799.8000 945.6000 ;
	    RECT 791.4000 944.5500 799.8000 945.4500 ;
	    RECT 791.4000 944.4000 792.6000 944.5500 ;
	    RECT 798.6000 944.4000 799.8000 944.5500 ;
	    RECT 724.2000 942.4500 725.4000 942.6000 ;
	    RECT 741.0000 942.4500 742.2000 942.6000 ;
	    RECT 724.2000 941.5500 742.2000 942.4500 ;
	    RECT 724.2000 941.4000 725.4000 941.5500 ;
	    RECT 741.0000 941.4000 742.2000 941.5500 ;
	    RECT 743.1000 940.8000 743.4000 942.3000 ;
	    RECT 745.5000 941.4000 747.3000 942.6000 ;
	    RECT 748.2000 942.4500 749.4000 942.6000 ;
	    RECT 765.0000 942.4500 766.2000 942.6000 ;
	    RECT 748.2000 941.5500 766.2000 942.4500 ;
	    RECT 748.2000 941.4000 749.4000 941.5500 ;
	    RECT 765.0000 941.4000 766.2000 941.5500 ;
	    RECT 645.0000 933.3000 646.2000 939.0000 ;
	    RECT 647.4000 933.3000 648.6000 936.3000 ;
	    RECT 678.6000 933.3000 679.8000 939.3000 ;
	    RECT 682.5000 933.3000 683.7000 939.0000 ;
	    RECT 684.9000 937.8000 687.0000 939.3000 ;
	    RECT 684.9000 933.3000 686.1000 937.8000 ;
	    RECT 710.7000 933.3000 711.9000 939.3000 ;
	    RECT 714.6000 933.3000 715.8000 939.3000 ;
	    RECT 717.0000 938.4000 718.2000 939.6000 ;
	    RECT 741.3000 939.3000 746.7000 939.9000 ;
	    RECT 748.2000 939.3000 749.1000 940.5000 ;
	    RECT 769.8000 939.3000 771.0000 943.5000 ;
	    RECT 798.6000 943.2000 799.8000 943.5000 ;
	    RECT 800.7000 942.6000 801.6000 947.7000 ;
	    RECT 803.4000 948.4500 804.6000 948.6000 ;
	    RECT 822.6000 948.4500 823.8000 948.6000 ;
	    RECT 803.4000 947.5500 823.8000 948.4500 ;
	    RECT 803.4000 947.4000 804.6000 947.5500 ;
	    RECT 822.6000 947.4000 823.8000 947.5500 ;
	    RECT 829.8000 947.4000 831.0000 948.6000 ;
	    RECT 832.8000 947.7000 834.3000 948.6000 ;
	    RECT 837.0000 947.7000 838.2000 959.7000 ;
	    RECT 856.2000 953.7000 857.4000 959.7000 ;
	    RECT 832.8000 942.6000 833.7000 947.7000 ;
	    RECT 858.6000 946.5000 859.8000 959.7000 ;
	    RECT 861.0000 953.7000 862.2000 959.7000 ;
	    RECT 863.4000 959.4000 864.6000 960.6000 ;
	    RECT 873.0000 953.7000 874.2000 959.7000 ;
	    RECT 861.0000 949.5000 862.2000 949.8000 ;
	    RECT 861.0000 947.4000 862.2000 948.6000 ;
	    RECT 834.6000 944.4000 835.8000 945.6000 ;
	    RECT 839.4000 945.4500 840.6000 945.6000 ;
	    RECT 858.6000 945.4500 859.8000 945.6000 ;
	    RECT 839.4000 944.5500 859.8000 945.4500 ;
	    RECT 839.4000 944.4000 840.6000 944.5500 ;
	    RECT 858.6000 944.4000 859.8000 944.5500 ;
	    RECT 875.4000 943.5000 876.6000 959.7000 ;
	    RECT 889.8000 953.7000 891.0000 959.7000 ;
	    RECT 892.2000 943.5000 893.4000 959.7000 ;
	    RECT 930.6000 947.7000 931.8000 959.7000 ;
	    RECT 934.5000 947.7000 937.5000 959.7000 ;
	    RECT 940.2000 947.7000 941.4000 959.7000 ;
	    RECT 959.4000 953.7000 960.6000 959.7000 ;
	    RECT 933.0000 944.4000 934.2000 945.6000 ;
	    RECT 930.6000 943.5000 931.8000 943.8000 ;
	    RECT 935.7000 943.5000 936.6000 947.7000 ;
	    RECT 961.8000 946.5000 963.0000 959.7000 ;
	    RECT 964.2000 953.7000 965.4000 959.7000 ;
	    RECT 1072.2001 959.4000 1073.4000 960.6000 ;
	    RECT 1019.4000 957.4500 1020.6000 957.6000 ;
	    RECT 1033.8000 957.4500 1035.0000 957.6000 ;
	    RECT 1019.4000 956.5500 1035.0000 957.4500 ;
	    RECT 1019.4000 956.4000 1020.6000 956.5500 ;
	    RECT 1033.8000 956.4000 1035.0000 956.5500 ;
	    RECT 1089.0000 953.7000 1090.2001 959.7000 ;
	    RECT 1091.4000 952.5000 1092.6000 959.7000 ;
	    RECT 1093.8000 953.7000 1095.0000 959.7000 ;
	    RECT 1096.2001 952.8000 1097.4000 959.7000 ;
	    RECT 1098.6000 953.7000 1099.8000 959.7000 ;
	    RECT 1093.5000 951.9000 1097.4000 952.8000 ;
	    RECT 990.6000 951.4500 991.8000 951.6000 ;
	    RECT 1089.0000 951.4500 1090.2001 951.6000 ;
	    RECT 1091.4000 951.4500 1092.6000 951.6000 ;
	    RECT 990.6000 950.5500 1092.6000 951.4500 ;
	    RECT 990.6000 950.4000 991.8000 950.5500 ;
	    RECT 1089.0000 950.4000 1090.2001 950.5500 ;
	    RECT 1091.4000 950.4000 1092.6000 950.5500 ;
	    RECT 964.2000 949.5000 965.4000 949.8000 ;
	    RECT 1093.5000 949.5000 1094.4000 951.9000 ;
	    RECT 1101.0000 951.6000 1102.2001 959.7000 ;
	    RECT 1103.4000 953.7000 1104.6000 959.7000 ;
	    RECT 1105.8000 955.5000 1107.0000 959.7000 ;
	    RECT 1108.2001 955.5000 1109.4000 959.7000 ;
	    RECT 1110.6000 955.5000 1111.8000 959.7000 ;
	    RECT 1103.1000 951.6000 1109.4000 952.8000 ;
	    RECT 1098.3000 950.4000 1102.2001 951.6000 ;
	    RECT 1113.0000 950.4000 1114.2001 959.7000 ;
	    RECT 1115.4000 953.7000 1116.6000 959.7000 ;
	    RECT 1117.8000 952.5000 1119.0000 959.7000 ;
	    RECT 1120.2001 953.7000 1121.4000 959.7000 ;
	    RECT 1122.6000 952.5000 1123.8000 959.7000 ;
	    RECT 1125.0000 955.5000 1126.2001 959.7000 ;
	    RECT 1127.4000 955.5000 1128.6000 959.7000 ;
	    RECT 1129.8000 953.7000 1131.0000 959.7000 ;
	    RECT 1132.2001 952.8000 1133.4000 959.7000 ;
	    RECT 1134.6000 953.7000 1135.8000 960.6000 ;
	    RECT 1137.0000 954.6000 1138.2001 959.7000 ;
	    RECT 1137.0000 953.7000 1138.5000 954.6000 ;
	    RECT 1139.4000 953.7000 1140.6000 959.7000 ;
	    RECT 1165.8000 953.7000 1167.0000 959.7000 ;
	    RECT 1137.6000 952.8000 1138.5000 953.7000 ;
	    RECT 1130.4000 951.6000 1136.7001 952.8000 ;
	    RECT 1137.6000 951.9000 1140.6000 952.8000 ;
	    RECT 1117.8000 950.4000 1121.7001 951.6000 ;
	    RECT 1122.6000 950.7000 1131.3000 951.6000 ;
	    RECT 1135.8000 951.0000 1136.7001 951.6000 ;
	    RECT 1105.8000 949.5000 1107.0000 949.8000 ;
	    RECT 964.2000 948.4500 965.4000 948.6000 ;
	    RECT 976.2000 948.4500 977.4000 948.6000 ;
	    RECT 964.2000 947.5500 977.4000 948.4500 ;
	    RECT 1091.4000 948.0000 1092.6000 949.5000 ;
	    RECT 964.2000 947.4000 965.4000 947.5500 ;
	    RECT 976.2000 947.4000 977.4000 947.5500 ;
	    RECT 1091.1000 946.8000 1092.6000 948.0000 ;
	    RECT 1093.5000 948.6000 1107.0000 949.5000 ;
	    RECT 1110.6000 949.5000 1111.8000 949.8000 ;
	    RECT 1122.6000 949.5000 1123.5000 950.7000 ;
	    RECT 1132.2001 949.8000 1134.3000 950.7000 ;
	    RECT 1135.8000 949.8000 1138.2001 951.0000 ;
	    RECT 1110.6000 948.6000 1123.5000 949.5000 ;
	    RECT 1125.0000 949.5000 1134.3000 949.8000 ;
	    RECT 1125.0000 948.9000 1133.1000 949.5000 ;
	    RECT 1125.0000 948.6000 1126.2001 948.9000 ;
	    RECT 937.8000 944.4000 939.0000 945.6000 ;
	    RECT 961.8000 945.4500 963.0000 945.6000 ;
	    RECT 1000.2000 945.4500 1001.4000 945.6000 ;
	    RECT 961.8000 944.5500 1001.4000 945.4500 ;
	    RECT 961.8000 944.4000 963.0000 944.5500 ;
	    RECT 1000.2000 944.4000 1001.4000 944.5500 ;
	    RECT 834.6000 943.2000 835.8000 943.5000 ;
	    RECT 772.2000 941.4000 773.4000 942.6000 ;
	    RECT 796.2000 941.4000 797.4000 942.6000 ;
	    RECT 798.3000 940.8000 798.6000 942.3000 ;
	    RECT 800.7000 941.4000 802.5000 942.6000 ;
	    RECT 803.4000 942.4500 804.6000 942.6000 ;
	    RECT 825.0000 942.4500 826.2000 942.6000 ;
	    RECT 803.4000 941.5500 826.2000 942.4500 ;
	    RECT 803.4000 941.4000 804.6000 941.5500 ;
	    RECT 825.0000 941.4000 826.2000 941.5500 ;
	    RECT 827.4000 942.4500 828.6000 942.6000 ;
	    RECT 829.8000 942.4500 831.0000 942.6000 ;
	    RECT 827.4000 941.5500 831.0000 942.4500 ;
	    RECT 827.4000 941.4000 828.6000 941.5500 ;
	    RECT 829.8000 941.4000 831.0000 941.5500 ;
	    RECT 831.9000 941.4000 833.7000 942.6000 ;
	    RECT 835.8000 940.8000 836.1000 942.3000 ;
	    RECT 837.0000 941.4000 838.2000 942.6000 ;
	    RECT 856.2000 941.4000 857.4000 942.6000 ;
	    RECT 772.2000 940.2000 773.4000 940.5000 ;
	    RECT 796.5000 939.3000 801.9000 939.9000 ;
	    RECT 803.4000 939.3000 804.3000 940.5000 ;
	    RECT 830.1000 939.3000 831.0000 940.5000 ;
	    RECT 856.2000 940.2000 857.4000 940.5000 ;
	    RECT 832.5000 939.3000 837.9000 939.9000 ;
	    RECT 858.6000 939.3000 859.8000 943.5000 ;
	    RECT 933.0000 943.2000 934.2000 943.5000 ;
	    RECT 937.8000 943.2000 939.0000 943.5000 ;
	    RECT 863.4000 942.4500 864.6000 942.6000 ;
	    RECT 875.4000 942.4500 876.6000 942.6000 ;
	    RECT 863.4000 941.5500 876.6000 942.4500 ;
	    RECT 863.4000 941.4000 864.6000 941.5500 ;
	    RECT 875.4000 941.4000 876.6000 941.5500 ;
	    RECT 892.2000 942.4500 893.4000 942.6000 ;
	    RECT 930.6000 942.4500 931.8000 942.6000 ;
	    RECT 892.2000 941.5500 931.8000 942.4500 ;
	    RECT 892.2000 941.4000 893.4000 941.5500 ;
	    RECT 930.6000 941.4000 931.8000 941.5500 ;
	    RECT 933.0000 941.4000 934.5000 942.3000 ;
	    RECT 935.4000 941.4000 936.6000 942.6000 ;
	    RECT 940.2000 942.4500 941.4000 942.6000 ;
	    RECT 942.6000 942.4500 943.8000 942.6000 ;
	    RECT 865.8000 939.4500 867.0000 939.6000 ;
	    RECT 873.0000 939.4500 874.2000 939.6000 ;
	    RECT 741.0000 939.0000 747.0000 939.3000 ;
	    RECT 716.7000 937.2000 717.9000 937.5000 ;
	    RECT 717.0000 933.3000 718.2000 936.3000 ;
	    RECT 741.0000 933.3000 742.2000 939.0000 ;
	    RECT 743.4000 933.3000 744.6000 938.1000 ;
	    RECT 745.8000 933.3000 747.0000 939.0000 ;
	    RECT 748.2000 933.3000 749.4000 939.3000 ;
	    RECT 768.3000 938.4000 771.0000 939.3000 ;
	    RECT 768.3000 933.3000 769.5000 938.4000 ;
	    RECT 772.2000 933.3000 773.4000 939.3000 ;
	    RECT 796.2000 939.0000 802.2000 939.3000 ;
	    RECT 796.2000 933.3000 797.4000 939.0000 ;
	    RECT 798.6000 933.3000 799.8000 938.1000 ;
	    RECT 801.0000 933.3000 802.2000 939.0000 ;
	    RECT 803.4000 933.3000 804.6000 939.3000 ;
	    RECT 829.8000 933.3000 831.0000 939.3000 ;
	    RECT 832.2000 939.0000 838.2000 939.3000 ;
	    RECT 832.2000 933.3000 833.4000 939.0000 ;
	    RECT 834.6000 933.3000 835.8000 938.1000 ;
	    RECT 837.0000 933.3000 838.2000 939.0000 ;
	    RECT 856.2000 933.3000 857.4000 939.3000 ;
	    RECT 858.6000 938.4000 861.3000 939.3000 ;
	    RECT 865.8000 938.5500 874.2000 939.4500 ;
	    RECT 865.8000 938.4000 867.0000 938.5500 ;
	    RECT 873.0000 938.4000 874.2000 938.5500 ;
	    RECT 860.1000 933.3000 861.3000 938.4000 ;
	    RECT 873.0000 937.2000 874.2000 937.5000 ;
	    RECT 873.0000 933.3000 874.2000 936.3000 ;
	    RECT 875.4000 933.3000 876.6000 940.5000 ;
	    RECT 889.8000 938.4000 891.0000 939.6000 ;
	    RECT 889.8000 937.2000 891.0000 937.5000 ;
	    RECT 889.8000 933.3000 891.0000 936.3000 ;
	    RECT 892.2000 933.3000 893.4000 940.5000 ;
	    RECT 933.0000 939.3000 933.9000 941.4000 ;
	    RECT 939.0000 940.8000 939.3000 942.3000 ;
	    RECT 940.2000 941.5500 943.8000 942.4500 ;
	    RECT 940.2000 941.4000 941.4000 941.5500 ;
	    RECT 942.6000 941.4000 943.8000 941.5500 ;
	    RECT 959.4000 941.4000 960.6000 942.6000 ;
	    RECT 959.4000 940.2000 960.6000 940.5000 ;
	    RECT 935.7000 939.3000 941.1000 939.9000 ;
	    RECT 961.8000 939.3000 963.0000 943.5000 ;
	    RECT 973.8000 942.4500 975.0000 942.6000 ;
	    RECT 1069.8000 942.4500 1071.0000 942.6000 ;
	    RECT 973.8000 941.5500 1071.0000 942.4500 ;
	    RECT 973.8000 941.4000 975.0000 941.5500 ;
	    RECT 1069.8000 941.4000 1071.0000 941.5500 ;
	    RECT 1091.1000 940.2000 1092.3000 946.8000 ;
	    RECT 1093.5000 945.9000 1094.4000 948.6000 ;
	    RECT 1129.5000 947.7000 1130.7001 948.0000 ;
	    RECT 1095.3000 946.8000 1133.7001 947.7000 ;
	    RECT 1134.6000 947.4000 1135.8000 948.6000 ;
	    RECT 1095.3000 946.5000 1096.5000 946.8000 ;
	    RECT 1093.2001 945.0000 1094.4000 945.9000 ;
	    RECT 1103.4000 945.0000 1128.9000 945.9000 ;
	    RECT 1093.2001 942.0000 1094.1000 945.0000 ;
	    RECT 1103.4000 944.1000 1104.6000 945.0000 ;
	    RECT 1129.8000 944.4000 1131.0000 945.6000 ;
	    RECT 1131.9000 945.0000 1138.5000 945.9000 ;
	    RECT 1137.3000 944.7000 1138.5000 945.0000 ;
	    RECT 1095.0000 942.9000 1100.7001 944.1000 ;
	    RECT 1093.2001 941.1000 1095.0000 942.0000 ;
	    RECT 930.6000 934.2000 931.8000 939.3000 ;
	    RECT 933.0000 935.1000 934.2000 939.3000 ;
	    RECT 935.4000 939.0000 941.4000 939.3000 ;
	    RECT 935.4000 934.2000 936.6000 939.0000 ;
	    RECT 930.6000 933.3000 936.6000 934.2000 ;
	    RECT 937.8000 933.3000 939.0000 938.1000 ;
	    RECT 940.2000 933.3000 941.4000 939.0000 ;
	    RECT 959.4000 933.3000 960.6000 939.3000 ;
	    RECT 961.8000 938.4000 964.5000 939.3000 ;
	    RECT 1091.1000 939.0000 1092.6000 940.2000 ;
	    RECT 963.3000 933.3000 964.5000 938.4000 ;
	    RECT 1089.0000 933.3000 1090.2001 936.3000 ;
	    RECT 1091.4000 933.3000 1092.6000 939.0000 ;
	    RECT 1093.8000 933.3000 1095.0000 941.1000 ;
	    RECT 1099.5000 941.1000 1100.7001 942.9000 ;
	    RECT 1099.5000 940.2000 1102.2001 941.1000 ;
	    RECT 1101.0000 939.3000 1102.2001 940.2000 ;
	    RECT 1108.2001 939.6000 1109.4000 943.8000 ;
	    RECT 1113.0000 942.9000 1117.8000 944.1000 ;
	    RECT 1123.5000 942.9000 1126.5000 944.1000 ;
	    RECT 1139.4000 943.5000 1140.6000 951.9000 ;
	    RECT 1165.8000 949.5000 1167.0000 949.8000 ;
	    RECT 1149.0000 948.4500 1150.2001 948.6000 ;
	    RECT 1165.8000 948.4500 1167.0000 948.6000 ;
	    RECT 1149.0000 947.5500 1167.0000 948.4500 ;
	    RECT 1149.0000 947.4000 1150.2001 947.5500 ;
	    RECT 1165.8000 947.4000 1167.0000 947.5500 ;
	    RECT 1168.2001 946.5000 1169.4000 959.7000 ;
	    RECT 1170.6000 953.7000 1171.8000 959.7000 ;
	    RECT 1297.8000 953.7000 1299.0000 959.7000 ;
	    RECT 1300.2001 954.6000 1301.4000 959.7000 ;
	    RECT 1299.9000 953.7000 1301.4000 954.6000 ;
	    RECT 1302.6000 953.7000 1303.8000 960.6000 ;
	    RECT 1299.9000 952.8000 1300.8000 953.7000 ;
	    RECT 1305.0000 952.8000 1306.2001 959.7000 ;
	    RECT 1307.4000 953.7000 1308.6000 959.7000 ;
	    RECT 1309.8000 955.5000 1311.0000 959.7000 ;
	    RECT 1312.2001 955.5000 1313.4000 959.7000 ;
	    RECT 1297.8000 951.9000 1300.8000 952.8000 ;
	    RECT 1168.2001 945.4500 1169.4000 945.6000 ;
	    RECT 1240.2001 945.4500 1241.4000 945.6000 ;
	    RECT 1168.2001 944.5500 1241.4000 945.4500 ;
	    RECT 1168.2001 944.4000 1169.4000 944.5500 ;
	    RECT 1240.2001 944.4000 1241.4000 944.5500 ;
	    RECT 1297.8000 943.5000 1299.0000 951.9000 ;
	    RECT 1301.7001 951.6000 1308.0000 952.8000 ;
	    RECT 1314.6000 952.5000 1315.8000 959.7000 ;
	    RECT 1317.0000 953.7000 1318.2001 959.7000 ;
	    RECT 1319.4000 952.5000 1320.6000 959.7000 ;
	    RECT 1321.8000 953.7000 1323.0000 959.7000 ;
	    RECT 1301.7001 951.0000 1302.6000 951.6000 ;
	    RECT 1300.2001 949.8000 1302.6000 951.0000 ;
	    RECT 1307.1000 950.7000 1315.8000 951.6000 ;
	    RECT 1304.1000 949.8000 1306.2001 950.7000 ;
	    RECT 1304.1000 949.5000 1313.4000 949.8000 ;
	    RECT 1305.3000 948.9000 1313.4000 949.5000 ;
	    RECT 1312.2001 948.6000 1313.4000 948.9000 ;
	    RECT 1314.9000 949.5000 1315.8000 950.7000 ;
	    RECT 1316.7001 950.4000 1320.6000 951.6000 ;
	    RECT 1324.2001 950.4000 1325.4000 959.7000 ;
	    RECT 1326.6000 955.5000 1327.8000 959.7000 ;
	    RECT 1329.0000 955.5000 1330.2001 959.7000 ;
	    RECT 1331.4000 955.5000 1332.6000 959.7000 ;
	    RECT 1333.8000 953.7000 1335.0000 959.7000 ;
	    RECT 1329.0000 951.6000 1335.3000 952.8000 ;
	    RECT 1336.2001 951.6000 1337.4000 959.7000 ;
	    RECT 1338.6000 953.7000 1339.8000 959.7000 ;
	    RECT 1341.0000 952.8000 1342.2001 959.7000 ;
	    RECT 1343.4000 953.7000 1344.6000 959.7000 ;
	    RECT 1341.0000 951.9000 1344.9000 952.8000 ;
	    RECT 1345.8000 952.5000 1347.0000 959.7000 ;
	    RECT 1348.2001 953.7000 1349.4000 959.7000 ;
	    RECT 1377.0000 959.4000 1378.2001 960.6000 ;
	    RECT 1379.4000 953.7000 1380.6000 959.7000 ;
	    RECT 1381.8000 954.3000 1383.0000 959.7000 ;
	    RECT 1379.7001 953.4000 1380.6000 953.7000 ;
	    RECT 1384.2001 953.7000 1385.4000 959.7000 ;
	    RECT 1386.6000 953.7000 1387.8000 959.7000 ;
	    RECT 1444.2001 957.4500 1445.4000 957.6000 ;
	    RECT 1509.0000 957.4500 1510.2001 957.6000 ;
	    RECT 1444.2001 956.5500 1510.2001 957.4500 ;
	    RECT 1444.2001 956.4000 1445.4000 956.5500 ;
	    RECT 1509.0000 956.4000 1510.2001 956.5500 ;
	    RECT 1511.4000 953.7000 1512.6000 959.7000 ;
	    RECT 1384.2001 953.4000 1385.1000 953.7000 ;
	    RECT 1379.7001 952.5000 1385.1000 953.4000 ;
	    RECT 1513.8000 952.5000 1515.0000 959.7000 ;
	    RECT 1516.2001 953.7000 1517.4000 959.7000 ;
	    RECT 1518.6000 952.8000 1519.8000 959.7000 ;
	    RECT 1521.0000 953.7000 1522.2001 959.7000 ;
	    RECT 1336.2001 950.4000 1340.1000 951.6000 ;
	    RECT 1326.6000 949.5000 1327.8000 949.8000 ;
	    RECT 1314.9000 948.6000 1327.8000 949.5000 ;
	    RECT 1331.4000 949.5000 1332.6000 949.8000 ;
	    RECT 1344.0000 949.5000 1344.9000 951.9000 ;
	    RECT 1345.8000 950.4000 1347.0000 951.6000 ;
	    RECT 1379.7001 949.5000 1380.6000 952.5000 ;
	    RECT 1515.9000 951.9000 1519.8000 952.8000 ;
	    RECT 1381.8000 951.4500 1383.0000 951.6000 ;
	    RECT 1408.2001 951.4500 1409.4000 951.6000 ;
	    RECT 1432.2001 951.4500 1433.4000 951.6000 ;
	    RECT 1468.2001 951.4500 1469.4000 951.6000 ;
	    RECT 1381.8000 950.5500 1469.4000 951.4500 ;
	    RECT 1381.8000 950.4000 1383.0000 950.5500 ;
	    RECT 1408.2001 950.4000 1409.4000 950.5500 ;
	    RECT 1432.2001 950.4000 1433.4000 950.5500 ;
	    RECT 1468.2001 950.4000 1469.4000 950.5500 ;
	    RECT 1473.0000 951.4500 1474.2001 951.6000 ;
	    RECT 1513.8000 951.4500 1515.0000 951.6000 ;
	    RECT 1473.0000 950.5500 1515.0000 951.4500 ;
	    RECT 1473.0000 950.4000 1474.2001 950.5500 ;
	    RECT 1513.8000 950.4000 1515.0000 950.5500 ;
	    RECT 1515.9000 949.5000 1516.8000 951.9000 ;
	    RECT 1523.4000 951.6000 1524.6000 959.7000 ;
	    RECT 1525.8000 953.7000 1527.0000 959.7000 ;
	    RECT 1528.2001 955.5000 1529.4000 959.7000 ;
	    RECT 1530.6000 955.5000 1531.8000 959.7000 ;
	    RECT 1533.0000 955.5000 1534.2001 959.7000 ;
	    RECT 1525.5000 951.6000 1531.8000 952.8000 ;
	    RECT 1520.7001 950.4000 1524.6000 951.6000 ;
	    RECT 1535.4000 950.4000 1536.6000 959.7000 ;
	    RECT 1537.8000 953.7000 1539.0000 959.7000 ;
	    RECT 1540.2001 952.5000 1541.4000 959.7000 ;
	    RECT 1542.6000 953.7000 1543.8000 959.7000 ;
	    RECT 1545.0000 952.5000 1546.2001 959.7000 ;
	    RECT 1547.4000 955.5000 1548.6000 959.7000 ;
	    RECT 1549.8000 955.5000 1551.0000 959.7000 ;
	    RECT 1552.2001 953.7000 1553.4000 959.7000 ;
	    RECT 1554.6000 952.8000 1555.8000 959.7000 ;
	    RECT 1557.0000 953.7000 1558.2001 960.6000 ;
	    RECT 1559.4000 954.6000 1560.6000 959.7000 ;
	    RECT 1559.4000 953.7000 1560.9000 954.6000 ;
	    RECT 1561.8000 953.7000 1563.0000 959.7000 ;
	    RECT 1560.0000 952.8000 1560.9000 953.7000 ;
	    RECT 1552.8000 951.6000 1559.1000 952.8000 ;
	    RECT 1560.0000 951.9000 1563.0000 952.8000 ;
	    RECT 1540.2001 950.4000 1544.1000 951.6000 ;
	    RECT 1545.0000 950.7000 1553.7001 951.6000 ;
	    RECT 1558.2001 951.0000 1559.1000 951.6000 ;
	    RECT 1528.2001 949.5000 1529.4000 949.8000 ;
	    RECT 1331.4000 948.6000 1344.9000 949.5000 ;
	    RECT 1302.6000 947.4000 1303.8000 948.6000 ;
	    RECT 1307.7001 947.7000 1308.9000 948.0000 ;
	    RECT 1304.7001 946.8000 1343.1000 947.7000 ;
	    RECT 1341.9000 946.5000 1343.1000 946.8000 ;
	    RECT 1344.0000 945.9000 1344.9000 948.6000 ;
	    RECT 1345.8000 948.0000 1347.0000 949.5000 ;
	    RECT 1381.8000 949.2000 1383.0000 949.5000 ;
	    RECT 1345.8000 946.8000 1347.3000 948.0000 ;
	    RECT 1379.4000 947.4000 1380.6000 948.6000 ;
	    RECT 1386.6000 948.4500 1387.8000 948.6000 ;
	    RECT 1389.0000 948.4500 1390.2001 948.6000 ;
	    RECT 1386.6000 947.5500 1390.2001 948.4500 ;
	    RECT 1513.8000 948.0000 1515.0000 949.5000 ;
	    RECT 1386.6000 947.4000 1387.8000 947.5500 ;
	    RECT 1389.0000 947.4000 1390.2001 947.5500 ;
	    RECT 1299.9000 945.0000 1306.5000 945.9000 ;
	    RECT 1299.9000 944.7000 1301.1000 945.0000 ;
	    RECT 1307.4000 944.4000 1308.6000 945.6000 ;
	    RECT 1309.5000 945.0000 1335.0000 945.9000 ;
	    RECT 1344.0000 945.0000 1345.2001 945.9000 ;
	    RECT 1333.8000 944.1000 1335.0000 945.0000 ;
	    RECT 1112.4000 941.7000 1113.6000 942.0000 ;
	    RECT 1112.4000 940.8000 1119.0000 941.7000 ;
	    RECT 1120.2001 941.4000 1121.4000 942.6000 ;
	    RECT 1117.8000 940.5000 1119.0000 940.8000 ;
	    RECT 1120.2001 940.2000 1121.4000 940.5000 ;
	    RECT 1098.6000 933.3000 1099.8000 939.3000 ;
	    RECT 1101.0000 938.1000 1104.6000 939.3000 ;
	    RECT 1108.2001 938.4000 1109.7001 939.6000 ;
	    RECT 1114.2001 938.4000 1114.5000 939.6000 ;
	    RECT 1115.4000 938.4000 1116.6000 939.6000 ;
	    RECT 1117.8000 939.3000 1119.0000 939.6000 ;
	    RECT 1123.5000 939.3000 1124.7001 942.9000 ;
	    RECT 1127.4000 942.3000 1140.6000 943.5000 ;
	    RECT 1132.5000 940.2000 1137.0000 941.4000 ;
	    RECT 1132.5000 939.3000 1133.7001 940.2000 ;
	    RECT 1117.8000 938.4000 1124.7001 939.3000 ;
	    RECT 1103.4000 933.3000 1104.6000 938.1000 ;
	    RECT 1129.8000 938.1000 1133.7001 939.3000 ;
	    RECT 1105.8000 933.3000 1107.0000 937.5000 ;
	    RECT 1108.2001 933.3000 1109.4000 937.5000 ;
	    RECT 1110.6000 933.3000 1111.8000 937.5000 ;
	    RECT 1113.0000 933.3000 1114.2001 937.5000 ;
	    RECT 1115.4000 933.3000 1116.6000 936.3000 ;
	    RECT 1117.8000 933.3000 1119.0000 937.5000 ;
	    RECT 1120.2001 933.3000 1121.4000 936.3000 ;
	    RECT 1122.6000 933.3000 1123.8000 937.5000 ;
	    RECT 1125.0000 933.3000 1126.2001 937.5000 ;
	    RECT 1127.4000 933.3000 1128.6000 937.5000 ;
	    RECT 1129.8000 933.3000 1131.0000 938.1000 ;
	    RECT 1134.6000 933.3000 1135.8000 939.3000 ;
	    RECT 1139.4000 933.3000 1140.6000 942.3000 ;
	    RECT 1168.2001 939.3000 1169.4000 943.5000 ;
	    RECT 1170.6000 942.4500 1171.8000 942.6000 ;
	    RECT 1189.8000 942.4500 1191.0000 942.6000 ;
	    RECT 1170.6000 941.5500 1191.0000 942.4500 ;
	    RECT 1170.6000 941.4000 1171.8000 941.5500 ;
	    RECT 1189.8000 941.4000 1191.0000 941.5500 ;
	    RECT 1297.8000 942.3000 1311.0000 943.5000 ;
	    RECT 1311.9000 942.9000 1314.9000 944.1000 ;
	    RECT 1320.6000 942.9000 1325.4000 944.1000 ;
	    RECT 1170.6000 940.2000 1171.8000 940.5000 ;
	    RECT 1166.7001 938.4000 1169.4000 939.3000 ;
	    RECT 1166.7001 933.3000 1167.9000 938.4000 ;
	    RECT 1170.6000 933.3000 1171.8000 939.3000 ;
	    RECT 1297.8000 933.3000 1299.0000 942.3000 ;
	    RECT 1301.4000 940.2000 1305.9000 941.4000 ;
	    RECT 1304.7001 939.3000 1305.9000 940.2000 ;
	    RECT 1313.7001 939.3000 1314.9000 942.9000 ;
	    RECT 1317.0000 941.4000 1318.2001 942.6000 ;
	    RECT 1324.8000 941.7000 1326.0000 942.0000 ;
	    RECT 1319.4000 940.8000 1326.0000 941.7000 ;
	    RECT 1319.4000 940.5000 1320.6000 940.8000 ;
	    RECT 1317.0000 940.2000 1318.2001 940.5000 ;
	    RECT 1329.0000 939.6000 1330.2001 943.8000 ;
	    RECT 1337.7001 942.9000 1343.4000 944.1000 ;
	    RECT 1337.7001 941.1000 1338.9000 942.9000 ;
	    RECT 1344.3000 942.0000 1345.2001 945.0000 ;
	    RECT 1319.4000 939.3000 1320.6000 939.6000 ;
	    RECT 1302.6000 933.3000 1303.8000 939.3000 ;
	    RECT 1304.7001 938.1000 1308.6000 939.3000 ;
	    RECT 1313.7001 938.4000 1320.6000 939.3000 ;
	    RECT 1321.8000 938.4000 1323.0000 939.6000 ;
	    RECT 1323.9000 938.4000 1324.2001 939.6000 ;
	    RECT 1328.7001 938.4000 1330.2001 939.6000 ;
	    RECT 1336.2001 940.2000 1338.9000 941.1000 ;
	    RECT 1343.4000 941.1000 1345.2001 942.0000 ;
	    RECT 1336.2001 939.3000 1337.4000 940.2000 ;
	    RECT 1307.4000 933.3000 1308.6000 938.1000 ;
	    RECT 1333.8000 938.1000 1337.4000 939.3000 ;
	    RECT 1309.8000 933.3000 1311.0000 937.5000 ;
	    RECT 1312.2001 933.3000 1313.4000 937.5000 ;
	    RECT 1314.6000 933.3000 1315.8000 937.5000 ;
	    RECT 1317.0000 933.3000 1318.2001 936.3000 ;
	    RECT 1319.4000 933.3000 1320.6000 937.5000 ;
	    RECT 1321.8000 933.3000 1323.0000 936.3000 ;
	    RECT 1324.2001 933.3000 1325.4000 937.5000 ;
	    RECT 1326.6000 933.3000 1327.8000 937.5000 ;
	    RECT 1329.0000 933.3000 1330.2001 937.5000 ;
	    RECT 1331.4000 933.3000 1332.6000 937.5000 ;
	    RECT 1333.8000 933.3000 1335.0000 938.1000 ;
	    RECT 1338.6000 933.3000 1339.8000 939.3000 ;
	    RECT 1343.4000 933.3000 1344.6000 941.1000 ;
	    RECT 1346.1000 940.2000 1347.3000 946.8000 ;
	    RECT 1513.5000 946.8000 1515.0000 948.0000 ;
	    RECT 1515.9000 948.6000 1529.4000 949.5000 ;
	    RECT 1533.0000 949.5000 1534.2001 949.8000 ;
	    RECT 1545.0000 949.5000 1545.9000 950.7000 ;
	    RECT 1554.6000 949.8000 1556.7001 950.7000 ;
	    RECT 1558.2001 949.8000 1560.6000 951.0000 ;
	    RECT 1533.0000 948.6000 1545.9000 949.5000 ;
	    RECT 1547.4000 949.5000 1556.7001 949.8000 ;
	    RECT 1547.4000 948.9000 1555.5000 949.5000 ;
	    RECT 1547.4000 948.6000 1548.6000 948.9000 ;
	    RECT 1379.7001 942.6000 1380.6000 946.5000 ;
	    RECT 1386.6000 946.2000 1387.8000 946.5000 ;
	    RECT 1383.0000 944.4000 1383.3000 945.6000 ;
	    RECT 1384.2001 944.4000 1385.4000 945.6000 ;
	    RECT 1379.7001 942.3000 1382.1000 942.6000 ;
	    RECT 1379.7001 941.7000 1382.4000 942.3000 ;
	    RECT 1345.8000 939.0000 1347.3000 940.2000 ;
	    RECT 1345.8000 933.3000 1347.0000 939.0000 ;
	    RECT 1348.2001 933.3000 1349.4000 936.3000 ;
	    RECT 1381.2001 933.3000 1382.4000 941.7000 ;
	    RECT 1386.6000 933.3000 1387.8000 942.3000 ;
	    RECT 1513.5000 940.2000 1514.7001 946.8000 ;
	    RECT 1515.9000 945.9000 1516.8000 948.6000 ;
	    RECT 1557.0000 948.4500 1558.2001 948.6000 ;
	    RECT 1559.4000 948.4500 1560.6000 948.6000 ;
	    RECT 1551.9000 947.7000 1553.1000 948.0000 ;
	    RECT 1517.7001 946.8000 1556.1000 947.7000 ;
	    RECT 1557.0000 947.5500 1560.6000 948.4500 ;
	    RECT 1557.0000 947.4000 1558.2001 947.5500 ;
	    RECT 1559.4000 947.4000 1560.6000 947.5500 ;
	    RECT 1517.7001 946.5000 1518.9000 946.8000 ;
	    RECT 1515.6000 945.0000 1516.8000 945.9000 ;
	    RECT 1525.8000 945.0000 1551.3000 945.9000 ;
	    RECT 1515.6000 942.0000 1516.5000 945.0000 ;
	    RECT 1525.8000 944.1000 1527.0000 945.0000 ;
	    RECT 1552.2001 944.4000 1553.4000 945.6000 ;
	    RECT 1554.3000 945.0000 1560.9000 945.9000 ;
	    RECT 1559.7001 944.7000 1560.9000 945.0000 ;
	    RECT 1517.4000 942.9000 1523.1000 944.1000 ;
	    RECT 1515.6000 941.1000 1517.4000 942.0000 ;
	    RECT 1513.5000 939.0000 1515.0000 940.2000 ;
	    RECT 1511.4000 933.3000 1512.6000 936.3000 ;
	    RECT 1513.8000 933.3000 1515.0000 939.0000 ;
	    RECT 1516.2001 933.3000 1517.4000 941.1000 ;
	    RECT 1521.9000 941.1000 1523.1000 942.9000 ;
	    RECT 1521.9000 940.2000 1524.6000 941.1000 ;
	    RECT 1523.4000 939.3000 1524.6000 940.2000 ;
	    RECT 1530.6000 939.6000 1531.8000 943.8000 ;
	    RECT 1535.4000 942.9000 1540.2001 944.1000 ;
	    RECT 1545.9000 942.9000 1548.9000 944.1000 ;
	    RECT 1561.8000 943.5000 1563.0000 951.9000 ;
	    RECT 1534.8000 941.7000 1536.0000 942.0000 ;
	    RECT 1534.8000 940.8000 1541.4000 941.7000 ;
	    RECT 1542.6000 941.4000 1543.8000 942.6000 ;
	    RECT 1540.2001 940.5000 1541.4000 940.8000 ;
	    RECT 1542.6000 940.2000 1543.8000 940.5000 ;
	    RECT 1521.0000 933.3000 1522.2001 939.3000 ;
	    RECT 1523.4000 938.1000 1527.0000 939.3000 ;
	    RECT 1530.6000 938.4000 1532.1000 939.6000 ;
	    RECT 1536.6000 938.4000 1536.9000 939.6000 ;
	    RECT 1537.8000 938.4000 1539.0000 939.6000 ;
	    RECT 1540.2001 939.3000 1541.4000 939.6000 ;
	    RECT 1545.9000 939.3000 1547.1000 942.9000 ;
	    RECT 1549.8000 942.3000 1563.0000 943.5000 ;
	    RECT 1554.9000 940.2000 1559.4000 941.4000 ;
	    RECT 1554.9000 939.3000 1556.1000 940.2000 ;
	    RECT 1540.2001 938.4000 1547.1000 939.3000 ;
	    RECT 1525.8000 933.3000 1527.0000 938.1000 ;
	    RECT 1552.2001 938.1000 1556.1000 939.3000 ;
	    RECT 1528.2001 933.3000 1529.4000 937.5000 ;
	    RECT 1530.6000 933.3000 1531.8000 937.5000 ;
	    RECT 1533.0000 933.3000 1534.2001 937.5000 ;
	    RECT 1535.4000 933.3000 1536.6000 937.5000 ;
	    RECT 1537.8000 933.3000 1539.0000 936.3000 ;
	    RECT 1540.2001 933.3000 1541.4000 937.5000 ;
	    RECT 1542.6000 933.3000 1543.8000 936.3000 ;
	    RECT 1545.0000 933.3000 1546.2001 937.5000 ;
	    RECT 1547.4000 933.3000 1548.6000 937.5000 ;
	    RECT 1549.8000 933.3000 1551.0000 937.5000 ;
	    RECT 1552.2001 933.3000 1553.4000 938.1000 ;
	    RECT 1557.0000 933.3000 1558.2001 939.3000 ;
	    RECT 1561.8000 933.3000 1563.0000 942.3000 ;
	    RECT 1.2000 930.6000 1569.0000 932.4000 ;
	    RECT 18.6000 922.8000 19.8000 929.7000 ;
	    RECT 21.0000 923.7000 22.2000 929.7000 ;
	    RECT 18.6000 921.9000 21.9000 922.8000 ;
	    RECT 23.4000 922.5000 24.6000 929.7000 ;
	    RECT 42.6000 923.7000 43.8000 929.7000 ;
	    RECT 46.5000 924.6000 47.7000 929.7000 ;
	    RECT 45.0000 923.7000 47.7000 924.6000 ;
	    RECT 66.6000 923.7000 67.8000 929.7000 ;
	    RECT 70.5000 924.6000 71.7000 929.7000 ;
	    RECT 133.8000 927.4500 135.0000 927.6000 ;
	    RECT 191.4000 927.4500 192.6000 927.6000 ;
	    RECT 133.8000 926.5500 192.6000 927.4500 ;
	    RECT 133.8000 926.4000 135.0000 926.5500 ;
	    RECT 191.4000 926.4000 192.6000 926.5500 ;
	    RECT 69.0000 923.7000 71.7000 924.6000 ;
	    RECT 42.6000 922.5000 43.8000 922.8000 ;
	    RECT 18.6000 919.5000 19.8000 919.8000 ;
	    RECT 18.6000 917.4000 19.8000 918.6000 ;
	    RECT 21.0000 917.4000 21.9000 921.9000 ;
	    RECT 23.4000 921.4500 24.6000 921.6000 ;
	    RECT 25.8000 921.4500 27.0000 921.6000 ;
	    RECT 42.6000 921.4500 43.8000 921.6000 ;
	    RECT 23.4000 920.5500 43.8000 921.4500 ;
	    RECT 23.4000 920.4000 24.6000 920.5500 ;
	    RECT 25.8000 920.4000 27.0000 920.5500 ;
	    RECT 42.6000 920.4000 43.8000 920.5500 ;
	    RECT 45.0000 919.5000 46.2000 923.7000 ;
	    RECT 66.6000 922.5000 67.8000 922.8000 ;
	    RECT 54.6000 921.4500 55.8000 921.6000 ;
	    RECT 66.6000 921.4500 67.8000 921.6000 ;
	    RECT 54.6000 920.5500 67.8000 921.4500 ;
	    RECT 54.6000 920.4000 55.8000 920.5500 ;
	    RECT 66.6000 920.4000 67.8000 920.5500 ;
	    RECT 69.0000 919.5000 70.2000 923.7000 ;
	    RECT 203.4000 920.7000 204.6000 929.7000 ;
	    RECT 208.2000 923.7000 209.4000 929.7000 ;
	    RECT 213.0000 924.9000 214.2000 929.7000 ;
	    RECT 215.4000 925.5000 216.6000 929.7000 ;
	    RECT 217.8000 925.5000 219.0000 929.7000 ;
	    RECT 220.2000 925.5000 221.4000 929.7000 ;
	    RECT 222.6000 926.7000 223.8000 929.7000 ;
	    RECT 225.0000 925.5000 226.2000 929.7000 ;
	    RECT 227.4000 926.7000 228.6000 929.7000 ;
	    RECT 229.8000 925.5000 231.0000 929.7000 ;
	    RECT 232.2000 925.5000 233.4000 929.7000 ;
	    RECT 234.6000 925.5000 235.8000 929.7000 ;
	    RECT 237.0000 925.5000 238.2000 929.7000 ;
	    RECT 210.3000 923.7000 214.2000 924.9000 ;
	    RECT 239.4000 924.9000 240.6000 929.7000 ;
	    RECT 219.3000 923.7000 226.2000 924.6000 ;
	    RECT 210.3000 922.8000 211.5000 923.7000 ;
	    RECT 207.0000 921.6000 211.5000 922.8000 ;
	    RECT 203.4000 919.5000 216.6000 920.7000 ;
	    RECT 219.3000 920.1000 220.5000 923.7000 ;
	    RECT 225.0000 923.4000 226.2000 923.7000 ;
	    RECT 227.4000 923.4000 228.6000 924.6000 ;
	    RECT 229.5000 923.4000 229.8000 924.6000 ;
	    RECT 234.3000 923.4000 235.8000 924.6000 ;
	    RECT 239.4000 923.7000 243.0000 924.9000 ;
	    RECT 244.2000 923.7000 245.4000 929.7000 ;
	    RECT 222.6000 922.5000 223.8000 922.8000 ;
	    RECT 225.0000 922.2000 226.2000 922.5000 ;
	    RECT 222.6000 920.4000 223.8000 921.6000 ;
	    RECT 225.0000 921.3000 231.6000 922.2000 ;
	    RECT 230.4000 921.0000 231.6000 921.3000 ;
	    RECT 23.4000 918.6000 24.6000 919.5000 ;
	    RECT 21.0000 916.2000 22.8000 917.4000 ;
	    RECT 21.0000 915.3000 21.9000 916.2000 ;
	    RECT 23.7000 915.3000 24.6000 918.6000 ;
	    RECT 33.0000 918.4500 34.2000 918.6000 ;
	    RECT 45.0000 918.4500 46.2000 918.6000 ;
	    RECT 33.0000 917.5500 46.2000 918.4500 ;
	    RECT 33.0000 917.4000 34.2000 917.5500 ;
	    RECT 45.0000 917.4000 46.2000 917.5500 ;
	    RECT 47.4000 918.4500 48.6000 918.6000 ;
	    RECT 69.0000 918.4500 70.2000 918.6000 ;
	    RECT 47.4000 917.5500 70.2000 918.4500 ;
	    RECT 47.4000 917.4000 48.6000 917.5500 ;
	    RECT 69.0000 917.4000 70.2000 917.5500 ;
	    RECT 18.6000 914.4000 21.9000 915.3000 ;
	    RECT 18.6000 903.3000 19.8000 914.4000 ;
	    RECT 21.0000 903.3000 22.2000 913.5000 ;
	    RECT 23.4000 903.3000 24.6000 915.3000 ;
	    RECT 42.6000 903.3000 43.8000 909.3000 ;
	    RECT 45.0000 903.3000 46.2000 916.5000 ;
	    RECT 47.4000 914.4000 48.6000 915.6000 ;
	    RECT 47.4000 913.2000 48.6000 913.5000 ;
	    RECT 47.4000 903.3000 48.6000 909.3000 ;
	    RECT 66.6000 903.3000 67.8000 909.3000 ;
	    RECT 69.0000 903.3000 70.2000 916.5000 ;
	    RECT 71.4000 915.4500 72.6000 915.6000 ;
	    RECT 109.8000 915.4500 111.0000 915.6000 ;
	    RECT 71.4000 914.5500 111.0000 915.4500 ;
	    RECT 71.4000 914.4000 72.6000 914.5500 ;
	    RECT 109.8000 914.4000 111.0000 914.5500 ;
	    RECT 71.4000 913.2000 72.6000 913.5000 ;
	    RECT 203.4000 911.1000 204.6000 919.5000 ;
	    RECT 217.5000 918.9000 220.5000 920.1000 ;
	    RECT 226.2000 918.9000 231.0000 920.1000 ;
	    RECT 234.6000 919.2000 235.8000 923.4000 ;
	    RECT 241.8000 922.8000 243.0000 923.7000 ;
	    RECT 241.8000 921.9000 244.5000 922.8000 ;
	    RECT 243.3000 920.1000 244.5000 921.9000 ;
	    RECT 249.0000 921.9000 250.2000 929.7000 ;
	    RECT 251.4000 924.0000 252.6000 929.7000 ;
	    RECT 253.8000 926.7000 255.0000 929.7000 ;
	    RECT 265.8000 926.7000 267.0000 929.7000 ;
	    RECT 265.8000 925.5000 267.0000 925.8000 ;
	    RECT 251.4000 922.8000 252.9000 924.0000 ;
	    RECT 265.8000 923.4000 267.0000 924.6000 ;
	    RECT 249.0000 921.0000 250.8000 921.9000 ;
	    RECT 243.3000 918.9000 249.0000 920.1000 ;
	    RECT 205.5000 918.0000 206.7000 918.3000 ;
	    RECT 205.5000 917.1000 212.1000 918.0000 ;
	    RECT 213.0000 917.4000 214.2000 918.6000 ;
	    RECT 239.4000 918.0000 240.6000 918.9000 ;
	    RECT 249.9000 918.0000 250.8000 921.0000 ;
	    RECT 215.1000 917.1000 240.6000 918.0000 ;
	    RECT 249.6000 917.1000 250.8000 918.0000 ;
	    RECT 247.5000 916.2000 248.7000 916.5000 ;
	    RECT 208.2000 914.4000 209.4000 915.6000 ;
	    RECT 210.3000 915.3000 248.7000 916.2000 ;
	    RECT 213.3000 915.0000 214.5000 915.3000 ;
	    RECT 249.6000 914.4000 250.5000 917.1000 ;
	    RECT 251.7000 916.2000 252.9000 922.8000 ;
	    RECT 268.2000 922.5000 269.4000 929.7000 ;
	    RECT 268.2000 921.4500 269.4000 921.6000 ;
	    RECT 285.0000 921.4500 286.2000 921.6000 ;
	    RECT 268.2000 920.5500 286.2000 921.4500 ;
	    RECT 294.0000 921.3000 295.2000 929.7000 ;
	    RECT 268.2000 920.4000 269.4000 920.5500 ;
	    RECT 285.0000 920.4000 286.2000 920.5500 ;
	    RECT 292.5000 920.7000 295.2000 921.3000 ;
	    RECT 299.4000 920.7000 300.6000 929.7000 ;
	    RECT 313.8000 926.7000 315.0000 929.7000 ;
	    RECT 313.8000 925.5000 315.0000 925.8000 ;
	    RECT 313.8000 923.4000 315.0000 924.6000 ;
	    RECT 316.2000 922.5000 317.4000 929.7000 ;
	    RECT 330.6000 922.5000 331.8000 929.7000 ;
	    RECT 333.0000 926.7000 334.2000 929.7000 ;
	    RECT 333.0000 925.5000 334.2000 925.8000 ;
	    RECT 333.0000 923.4000 334.2000 924.6000 ;
	    RECT 301.8000 921.4500 303.0000 921.6000 ;
	    RECT 316.2000 921.4500 317.4000 921.6000 ;
	    RECT 328.2000 921.4500 329.4000 921.6000 ;
	    RECT 292.5000 920.4000 294.9000 920.7000 ;
	    RECT 301.8000 920.5500 329.4000 921.4500 ;
	    RECT 301.8000 920.4000 303.0000 920.5500 ;
	    RECT 316.2000 920.4000 317.4000 920.5500 ;
	    RECT 328.2000 920.4000 329.4000 920.5500 ;
	    RECT 330.6000 921.4500 331.8000 921.6000 ;
	    RECT 342.6000 921.4500 343.8000 921.6000 ;
	    RECT 330.6000 920.5500 343.8000 921.4500 ;
	    RECT 358.8000 921.3000 360.0000 929.7000 ;
	    RECT 330.6000 920.4000 331.8000 920.5500 ;
	    RECT 342.6000 920.4000 343.8000 920.5500 ;
	    RECT 357.3000 920.7000 360.0000 921.3000 ;
	    RECT 364.2000 920.7000 365.4000 929.7000 ;
	    RECT 376.2000 922.5000 377.4000 929.7000 ;
	    RECT 378.6000 926.7000 379.8000 929.7000 ;
	    RECT 393.0000 926.7000 394.2000 929.7000 ;
	    RECT 378.6000 925.5000 379.8000 925.8000 ;
	    RECT 393.0000 925.5000 394.2000 925.8000 ;
	    RECT 378.6000 924.4500 379.8000 924.6000 ;
	    RECT 388.2000 924.4500 389.4000 924.6000 ;
	    RECT 378.6000 923.5500 389.4000 924.4500 ;
	    RECT 378.6000 923.4000 379.8000 923.5500 ;
	    RECT 388.2000 923.4000 389.4000 923.5500 ;
	    RECT 393.0000 923.4000 394.2000 924.6000 ;
	    RECT 395.4000 922.5000 396.6000 929.7000 ;
	    RECT 376.2000 921.4500 377.4000 921.6000 ;
	    RECT 378.6000 921.4500 379.8000 921.6000 ;
	    RECT 357.3000 920.4000 359.7000 920.7000 ;
	    RECT 376.2000 920.5500 379.8000 921.4500 ;
	    RECT 376.2000 920.4000 377.4000 920.5500 ;
	    RECT 378.6000 920.4000 379.8000 920.5500 ;
	    RECT 395.4000 921.4500 396.6000 921.6000 ;
	    RECT 417.0000 921.4500 418.2000 921.6000 ;
	    RECT 395.4000 920.5500 418.2000 921.4500 ;
	    RECT 421.2000 921.3000 422.4000 929.7000 ;
	    RECT 395.4000 920.4000 396.6000 920.5500 ;
	    RECT 417.0000 920.4000 418.2000 920.5500 ;
	    RECT 419.7000 920.7000 422.4000 921.3000 ;
	    RECT 426.6000 920.7000 427.8000 929.7000 ;
	    RECT 448.2000 922.5000 449.4000 929.7000 ;
	    RECT 450.6000 926.7000 451.8000 929.7000 ;
	    RECT 465.0000 926.7000 466.2000 929.7000 ;
	    RECT 450.6000 925.5000 451.8000 925.8000 ;
	    RECT 465.0000 925.5000 466.2000 925.8000 ;
	    RECT 450.6000 924.4500 451.8000 924.6000 ;
	    RECT 453.0000 924.4500 454.2000 924.6000 ;
	    RECT 450.6000 923.5500 454.2000 924.4500 ;
	    RECT 450.6000 923.4000 451.8000 923.5500 ;
	    RECT 453.0000 923.4000 454.2000 923.5500 ;
	    RECT 465.0000 923.4000 466.2000 924.6000 ;
	    RECT 467.4000 922.5000 468.6000 929.7000 ;
	    RECT 491.4000 924.0000 492.6000 929.7000 ;
	    RECT 493.8000 924.9000 495.0000 929.7000 ;
	    RECT 496.2000 924.0000 497.4000 929.7000 ;
	    RECT 491.4000 923.7000 497.4000 924.0000 ;
	    RECT 498.6000 923.7000 499.8000 929.7000 ;
	    RECT 517.8000 923.7000 519.0000 929.7000 ;
	    RECT 521.7000 924.6000 522.9000 929.7000 ;
	    RECT 520.2000 923.7000 522.9000 924.6000 ;
	    RECT 541.8000 923.7000 543.0000 929.7000 ;
	    RECT 545.7000 924.6000 546.9000 929.7000 ;
	    RECT 544.2000 923.7000 546.9000 924.6000 ;
	    RECT 566.7000 924.6000 567.9000 929.7000 ;
	    RECT 566.7000 923.7000 569.4000 924.6000 ;
	    RECT 570.6000 923.7000 571.8000 929.7000 ;
	    RECT 597.0000 923.7000 598.2000 929.7000 ;
	    RECT 599.4000 924.0000 600.6000 929.7000 ;
	    RECT 601.8000 924.9000 603.0000 929.7000 ;
	    RECT 604.2000 924.0000 605.4000 929.7000 ;
	    RECT 599.4000 923.7000 605.4000 924.0000 ;
	    RECT 491.7000 923.1000 497.1000 923.7000 ;
	    RECT 498.6000 922.5000 499.5000 923.7000 ;
	    RECT 517.8000 922.5000 519.0000 922.8000 ;
	    RECT 429.0000 921.4500 430.2000 921.6000 ;
	    RECT 448.2000 921.4500 449.4000 921.6000 ;
	    RECT 419.7000 920.4000 422.1000 920.7000 ;
	    RECT 429.0000 920.5500 449.4000 921.4500 ;
	    RECT 429.0000 920.4000 430.2000 920.5500 ;
	    RECT 448.2000 920.4000 449.4000 920.5500 ;
	    RECT 467.4000 921.4500 468.6000 921.6000 ;
	    RECT 477.0000 921.4500 478.2000 921.6000 ;
	    RECT 491.4000 921.4500 492.6000 921.6000 ;
	    RECT 467.4000 920.5500 475.6500 921.4500 ;
	    RECT 467.4000 920.4000 468.6000 920.5500 ;
	    RECT 217.8000 914.1000 219.0000 914.4000 ;
	    RECT 210.9000 913.5000 219.0000 914.1000 ;
	    RECT 209.7000 913.2000 219.0000 913.5000 ;
	    RECT 220.5000 913.5000 233.4000 914.4000 ;
	    RECT 205.8000 912.0000 208.2000 913.2000 ;
	    RECT 209.7000 912.3000 211.8000 913.2000 ;
	    RECT 220.5000 912.3000 221.4000 913.5000 ;
	    RECT 232.2000 913.2000 233.4000 913.5000 ;
	    RECT 237.0000 913.5000 250.5000 914.4000 ;
	    RECT 251.4000 915.0000 252.9000 916.2000 ;
	    RECT 251.4000 913.5000 252.6000 915.0000 ;
	    RECT 237.0000 913.2000 238.2000 913.5000 ;
	    RECT 207.3000 911.4000 208.2000 912.0000 ;
	    RECT 212.7000 911.4000 221.4000 912.3000 ;
	    RECT 222.3000 911.4000 226.2000 912.6000 ;
	    RECT 203.4000 910.2000 206.4000 911.1000 ;
	    RECT 207.3000 910.2000 213.6000 911.4000 ;
	    RECT 205.5000 909.3000 206.4000 910.2000 ;
	    RECT 71.4000 903.3000 72.6000 909.3000 ;
	    RECT 203.4000 903.3000 204.6000 909.3000 ;
	    RECT 205.5000 908.4000 207.0000 909.3000 ;
	    RECT 205.8000 903.3000 207.0000 908.4000 ;
	    RECT 208.2000 902.4000 209.4000 909.3000 ;
	    RECT 210.6000 903.3000 211.8000 910.2000 ;
	    RECT 213.0000 903.3000 214.2000 909.3000 ;
	    RECT 215.4000 903.3000 216.6000 907.5000 ;
	    RECT 217.8000 903.3000 219.0000 907.5000 ;
	    RECT 220.2000 903.3000 221.4000 910.5000 ;
	    RECT 222.6000 903.3000 223.8000 909.3000 ;
	    RECT 225.0000 903.3000 226.2000 910.5000 ;
	    RECT 227.4000 903.3000 228.6000 909.3000 ;
	    RECT 229.8000 903.3000 231.0000 912.6000 ;
	    RECT 241.8000 911.4000 245.7000 912.6000 ;
	    RECT 234.6000 910.2000 240.9000 911.4000 ;
	    RECT 232.2000 903.3000 233.4000 907.5000 ;
	    RECT 234.6000 903.3000 235.8000 907.5000 ;
	    RECT 237.0000 903.3000 238.2000 907.5000 ;
	    RECT 239.4000 903.3000 240.6000 909.3000 ;
	    RECT 241.8000 903.3000 243.0000 911.4000 ;
	    RECT 249.6000 911.1000 250.5000 913.5000 ;
	    RECT 251.4000 911.4000 252.6000 912.6000 ;
	    RECT 246.6000 910.2000 250.5000 911.1000 ;
	    RECT 244.2000 903.3000 245.4000 909.3000 ;
	    RECT 246.6000 903.3000 247.8000 910.2000 ;
	    RECT 249.0000 903.3000 250.2000 909.3000 ;
	    RECT 251.4000 903.3000 252.6000 910.5000 ;
	    RECT 253.8000 903.3000 255.0000 909.3000 ;
	    RECT 265.8000 903.3000 267.0000 909.3000 ;
	    RECT 268.2000 903.3000 269.4000 919.5000 ;
	    RECT 292.5000 916.5000 293.4000 920.4000 ;
	    RECT 295.8000 917.4000 296.1000 918.6000 ;
	    RECT 297.0000 917.4000 298.2000 918.6000 ;
	    RECT 299.4000 916.5000 300.6000 916.8000 ;
	    RECT 292.2000 914.4000 293.4000 915.6000 ;
	    RECT 299.4000 914.4000 300.6000 915.6000 ;
	    RECT 294.6000 913.5000 295.8000 913.8000 ;
	    RECT 292.5000 910.5000 293.4000 913.5000 ;
	    RECT 294.6000 912.4500 295.8000 912.6000 ;
	    RECT 301.8000 912.4500 303.0000 912.6000 ;
	    RECT 294.6000 911.5500 303.0000 912.4500 ;
	    RECT 294.6000 911.4000 295.8000 911.5500 ;
	    RECT 301.8000 911.4000 303.0000 911.5500 ;
	    RECT 292.5000 909.6000 297.9000 910.5000 ;
	    RECT 292.5000 909.3000 293.4000 909.6000 ;
	    RECT 292.2000 903.3000 293.4000 909.3000 ;
	    RECT 297.0000 909.3000 297.9000 909.6000 ;
	    RECT 294.6000 903.3000 295.8000 908.7000 ;
	    RECT 297.0000 903.3000 298.2000 909.3000 ;
	    RECT 299.4000 903.3000 300.6000 909.3000 ;
	    RECT 313.8000 903.3000 315.0000 909.3000 ;
	    RECT 316.2000 903.3000 317.4000 919.5000 ;
	    RECT 330.6000 903.3000 331.8000 919.5000 ;
	    RECT 357.3000 916.5000 358.2000 920.4000 ;
	    RECT 360.6000 917.4000 360.9000 918.6000 ;
	    RECT 361.8000 917.4000 363.0000 918.6000 ;
	    RECT 364.2000 916.5000 365.4000 916.8000 ;
	    RECT 352.2000 915.4500 353.4000 915.6000 ;
	    RECT 357.0000 915.4500 358.2000 915.6000 ;
	    RECT 352.2000 914.5500 358.2000 915.4500 ;
	    RECT 352.2000 914.4000 353.4000 914.5500 ;
	    RECT 357.0000 914.4000 358.2000 914.5500 ;
	    RECT 364.2000 914.4000 365.4000 915.6000 ;
	    RECT 359.4000 913.5000 360.6000 913.8000 ;
	    RECT 357.3000 910.5000 358.2000 913.5000 ;
	    RECT 359.4000 912.4500 360.6000 912.6000 ;
	    RECT 371.4000 912.4500 372.6000 912.6000 ;
	    RECT 359.4000 911.5500 372.6000 912.4500 ;
	    RECT 359.4000 911.4000 360.6000 911.5500 ;
	    RECT 371.4000 911.4000 372.6000 911.5500 ;
	    RECT 357.3000 909.6000 362.7000 910.5000 ;
	    RECT 357.3000 909.3000 358.2000 909.6000 ;
	    RECT 333.0000 903.3000 334.2000 909.3000 ;
	    RECT 357.0000 903.3000 358.2000 909.3000 ;
	    RECT 361.8000 909.3000 362.7000 909.6000 ;
	    RECT 359.4000 903.3000 360.6000 908.7000 ;
	    RECT 361.8000 903.3000 363.0000 909.3000 ;
	    RECT 364.2000 903.3000 365.4000 909.3000 ;
	    RECT 376.2000 903.3000 377.4000 919.5000 ;
	    RECT 378.6000 903.3000 379.8000 909.3000 ;
	    RECT 393.0000 903.3000 394.2000 909.3000 ;
	    RECT 395.4000 903.3000 396.6000 919.5000 ;
	    RECT 419.7000 916.5000 420.6000 920.4000 ;
	    RECT 423.0000 917.4000 423.3000 918.6000 ;
	    RECT 424.2000 917.4000 425.4000 918.6000 ;
	    RECT 426.6000 916.5000 427.8000 916.8000 ;
	    RECT 409.8000 915.4500 411.0000 915.6000 ;
	    RECT 419.4000 915.4500 420.6000 915.6000 ;
	    RECT 409.8000 914.5500 420.6000 915.4500 ;
	    RECT 409.8000 914.4000 411.0000 914.5500 ;
	    RECT 419.4000 914.4000 420.6000 914.5500 ;
	    RECT 426.6000 914.4000 427.8000 915.6000 ;
	    RECT 421.8000 913.5000 423.0000 913.8000 ;
	    RECT 419.7000 910.5000 420.6000 913.5000 ;
	    RECT 421.8000 911.4000 423.0000 912.6000 ;
	    RECT 419.7000 909.6000 425.1000 910.5000 ;
	    RECT 419.7000 909.3000 420.6000 909.6000 ;
	    RECT 419.4000 903.3000 420.6000 909.3000 ;
	    RECT 424.2000 909.3000 425.1000 909.6000 ;
	    RECT 421.8000 903.3000 423.0000 908.7000 ;
	    RECT 424.2000 903.3000 425.4000 909.3000 ;
	    RECT 426.6000 903.3000 427.8000 909.3000 ;
	    RECT 448.2000 903.3000 449.4000 919.5000 ;
	    RECT 450.6000 903.3000 451.8000 909.3000 ;
	    RECT 465.0000 903.3000 466.2000 909.3000 ;
	    RECT 467.4000 903.3000 468.6000 919.5000 ;
	    RECT 474.7500 918.4500 475.6500 920.5500 ;
	    RECT 477.0000 920.5500 492.6000 921.4500 ;
	    RECT 493.5000 920.7000 493.8000 922.2000 ;
	    RECT 477.0000 920.4000 478.2000 920.5500 ;
	    RECT 491.4000 920.4000 492.6000 920.5500 ;
	    RECT 495.9000 920.4000 497.7000 921.6000 ;
	    RECT 498.6000 921.4500 499.8000 921.6000 ;
	    RECT 513.0000 921.4500 514.2000 921.6000 ;
	    RECT 498.6000 920.5500 514.2000 921.4500 ;
	    RECT 498.6000 920.4000 499.8000 920.5500 ;
	    RECT 513.0000 920.4000 514.2000 920.5500 ;
	    RECT 517.8000 920.4000 519.0000 921.6000 ;
	    RECT 493.8000 919.5000 495.0000 919.8000 ;
	    RECT 493.8000 918.4500 495.0000 918.6000 ;
	    RECT 474.7500 917.5500 495.0000 918.4500 ;
	    RECT 493.8000 917.4000 495.0000 917.5500 ;
	    RECT 495.9000 915.3000 496.8000 920.4000 ;
	    RECT 520.2000 919.5000 521.4000 923.7000 ;
	    RECT 541.8000 922.5000 543.0000 922.8000 ;
	    RECT 534.6000 921.4500 535.8000 921.6000 ;
	    RECT 541.8000 921.4500 543.0000 921.6000 ;
	    RECT 534.6000 920.5500 543.0000 921.4500 ;
	    RECT 534.6000 920.4000 535.8000 920.5500 ;
	    RECT 541.8000 920.4000 543.0000 920.5500 ;
	    RECT 544.2000 919.5000 545.4000 923.7000 ;
	    RECT 568.2000 919.5000 569.4000 923.7000 ;
	    RECT 570.6000 922.5000 571.8000 922.8000 ;
	    RECT 597.3000 922.5000 598.2000 923.7000 ;
	    RECT 599.7000 923.1000 605.1000 923.7000 ;
	    RECT 616.2000 922.5000 617.4000 929.7000 ;
	    RECT 618.6000 926.7000 619.8000 929.7000 ;
	    RECT 621.0000 927.4500 622.2000 927.6000 ;
	    RECT 729.0000 927.4500 730.2000 927.6000 ;
	    RECT 741.0000 927.4500 742.2000 927.6000 ;
	    RECT 621.0000 926.5500 742.2000 927.4500 ;
	    RECT 621.0000 926.4000 622.2000 926.5500 ;
	    RECT 729.0000 926.4000 730.2000 926.5500 ;
	    RECT 741.0000 926.4000 742.2000 926.5500 ;
	    RECT 618.6000 925.5000 619.8000 925.8000 ;
	    RECT 618.6000 924.4500 619.8000 924.6000 ;
	    RECT 645.0000 924.4500 646.2000 924.6000 ;
	    RECT 618.6000 923.5500 646.2000 924.4500 ;
	    RECT 618.6000 923.4000 619.8000 923.5500 ;
	    RECT 645.0000 923.4000 646.2000 923.5500 ;
	    RECT 570.6000 921.4500 571.8000 921.6000 ;
	    RECT 592.2000 921.4500 593.4000 921.6000 ;
	    RECT 570.6000 920.5500 593.4000 921.4500 ;
	    RECT 570.6000 920.4000 571.8000 920.5500 ;
	    RECT 592.2000 920.4000 593.4000 920.5500 ;
	    RECT 597.0000 920.4000 598.2000 921.6000 ;
	    RECT 599.1000 920.4000 600.9000 921.6000 ;
	    RECT 603.0000 920.7000 603.3000 922.2000 ;
	    RECT 604.2000 920.4000 605.4000 921.6000 ;
	    RECT 616.2000 921.4500 617.4000 921.6000 ;
	    RECT 606.7500 920.5500 617.4000 921.4500 ;
	    RECT 498.6000 918.4500 499.8000 918.6000 ;
	    RECT 520.2000 918.4500 521.4000 918.6000 ;
	    RECT 498.6000 917.5500 521.4000 918.4500 ;
	    RECT 498.6000 917.4000 499.8000 917.5500 ;
	    RECT 520.2000 917.4000 521.4000 917.5500 ;
	    RECT 522.6000 918.4500 523.8000 918.6000 ;
	    RECT 544.2000 918.4500 545.4000 918.6000 ;
	    RECT 522.6000 917.5500 545.4000 918.4500 ;
	    RECT 522.6000 917.4000 523.8000 917.5500 ;
	    RECT 544.2000 917.4000 545.4000 917.5500 ;
	    RECT 568.2000 918.4500 569.4000 918.6000 ;
	    RECT 568.2000 917.5500 598.0500 918.4500 ;
	    RECT 568.2000 917.4000 569.4000 917.5500 ;
	    RECT 491.4000 903.3000 492.6000 915.3000 ;
	    RECT 495.3000 914.4000 496.8000 915.3000 ;
	    RECT 498.6000 915.4500 499.8000 915.6000 ;
	    RECT 517.8000 915.4500 519.0000 915.6000 ;
	    RECT 498.6000 914.5500 519.0000 915.4500 ;
	    RECT 498.6000 914.4000 499.8000 914.5500 ;
	    RECT 517.8000 914.4000 519.0000 914.5500 ;
	    RECT 495.3000 903.3000 496.5000 914.4000 ;
	    RECT 497.7000 912.6000 498.6000 913.5000 ;
	    RECT 497.4000 911.4000 498.6000 912.6000 ;
	    RECT 497.7000 903.3000 498.9000 909.3000 ;
	    RECT 517.8000 903.3000 519.0000 909.3000 ;
	    RECT 520.2000 903.3000 521.4000 916.5000 ;
	    RECT 522.6000 915.4500 523.8000 915.6000 ;
	    RECT 541.8000 915.4500 543.0000 915.6000 ;
	    RECT 522.6000 914.5500 543.0000 915.4500 ;
	    RECT 522.6000 914.4000 523.8000 914.5500 ;
	    RECT 541.8000 914.4000 543.0000 914.5500 ;
	    RECT 522.6000 913.2000 523.8000 913.5000 ;
	    RECT 522.6000 903.3000 523.8000 909.3000 ;
	    RECT 541.8000 903.3000 543.0000 909.3000 ;
	    RECT 544.2000 903.3000 545.4000 916.5000 ;
	    RECT 546.6000 915.4500 547.8000 915.6000 ;
	    RECT 565.8000 915.4500 567.0000 915.6000 ;
	    RECT 546.6000 914.5500 567.0000 915.4500 ;
	    RECT 546.6000 914.4000 547.8000 914.5500 ;
	    RECT 565.8000 914.4000 567.0000 914.5500 ;
	    RECT 546.6000 913.2000 547.8000 913.5000 ;
	    RECT 565.8000 913.2000 567.0000 913.5000 ;
	    RECT 546.6000 903.3000 547.8000 909.3000 ;
	    RECT 565.8000 903.3000 567.0000 909.3000 ;
	    RECT 568.2000 903.3000 569.4000 916.5000 ;
	    RECT 597.1500 915.6000 598.0500 917.5500 ;
	    RECT 597.0000 914.4000 598.2000 915.6000 ;
	    RECT 600.0000 915.3000 600.9000 920.4000 ;
	    RECT 601.8000 919.5000 603.0000 919.8000 ;
	    RECT 601.8000 918.4500 603.0000 918.6000 ;
	    RECT 606.7500 918.4500 607.6500 920.5500 ;
	    RECT 616.2000 920.4000 617.4000 920.5500 ;
	    RECT 750.6000 920.7000 751.8000 929.7000 ;
	    RECT 755.4000 923.7000 756.6000 929.7000 ;
	    RECT 760.2000 924.9000 761.4000 929.7000 ;
	    RECT 762.6000 925.5000 763.8000 929.7000 ;
	    RECT 765.0000 925.5000 766.2000 929.7000 ;
	    RECT 767.4000 925.5000 768.6000 929.7000 ;
	    RECT 769.8000 926.7000 771.0000 929.7000 ;
	    RECT 772.2000 925.5000 773.4000 929.7000 ;
	    RECT 774.6000 926.7000 775.8000 929.7000 ;
	    RECT 777.0000 925.5000 778.2000 929.7000 ;
	    RECT 779.4000 925.5000 780.6000 929.7000 ;
	    RECT 781.8000 925.5000 783.0000 929.7000 ;
	    RECT 784.2000 925.5000 785.4000 929.7000 ;
	    RECT 757.5000 923.7000 761.4000 924.9000 ;
	    RECT 786.6000 924.9000 787.8000 929.7000 ;
	    RECT 766.5000 923.7000 773.4000 924.6000 ;
	    RECT 757.5000 922.8000 758.7000 923.7000 ;
	    RECT 754.2000 921.6000 758.7000 922.8000 ;
	    RECT 750.6000 919.5000 763.8000 920.7000 ;
	    RECT 766.5000 920.1000 767.7000 923.7000 ;
	    RECT 772.2000 923.4000 773.4000 923.7000 ;
	    RECT 774.6000 923.4000 775.8000 924.6000 ;
	    RECT 776.7000 923.4000 777.0000 924.6000 ;
	    RECT 781.5000 923.4000 783.0000 924.6000 ;
	    RECT 786.6000 923.7000 790.2000 924.9000 ;
	    RECT 791.4000 923.7000 792.6000 929.7000 ;
	    RECT 769.8000 922.5000 771.0000 922.8000 ;
	    RECT 772.2000 922.2000 773.4000 922.5000 ;
	    RECT 769.8000 920.4000 771.0000 921.6000 ;
	    RECT 772.2000 921.3000 778.8000 922.2000 ;
	    RECT 777.6000 921.0000 778.8000 921.3000 ;
	    RECT 601.8000 917.5500 607.6500 918.4500 ;
	    RECT 601.8000 917.4000 603.0000 917.5500 ;
	    RECT 600.0000 914.4000 601.5000 915.3000 ;
	    RECT 598.2000 912.6000 599.1000 913.5000 ;
	    RECT 598.2000 911.4000 599.4000 912.6000 ;
	    RECT 570.6000 903.3000 571.8000 909.3000 ;
	    RECT 597.9000 903.3000 599.1000 909.3000 ;
	    RECT 600.3000 903.3000 601.5000 914.4000 ;
	    RECT 604.2000 903.3000 605.4000 915.3000 ;
	    RECT 616.2000 903.3000 617.4000 919.5000 ;
	    RECT 750.6000 911.1000 751.8000 919.5000 ;
	    RECT 764.7000 918.9000 767.7000 920.1000 ;
	    RECT 773.4000 918.9000 778.2000 920.1000 ;
	    RECT 781.8000 919.2000 783.0000 923.4000 ;
	    RECT 789.0000 922.8000 790.2000 923.7000 ;
	    RECT 789.0000 921.9000 791.7000 922.8000 ;
	    RECT 790.5000 920.1000 791.7000 921.9000 ;
	    RECT 796.2000 921.9000 797.4000 929.7000 ;
	    RECT 798.6000 924.0000 799.8000 929.7000 ;
	    RECT 801.0000 926.7000 802.2000 929.7000 ;
	    RECT 861.0000 927.4500 862.2000 927.6000 ;
	    RECT 863.4000 927.4500 864.6000 927.6000 ;
	    RECT 897.0000 927.4500 898.2000 927.6000 ;
	    RECT 861.0000 926.5500 898.2000 927.4500 ;
	    RECT 933.0000 926.7000 934.2000 929.7000 ;
	    RECT 861.0000 926.4000 862.2000 926.5500 ;
	    RECT 863.4000 926.4000 864.6000 926.5500 ;
	    RECT 897.0000 926.4000 898.2000 926.5500 ;
	    RECT 808.2000 924.4500 809.4000 924.6000 ;
	    RECT 933.0000 924.4500 934.2000 924.6000 ;
	    RECT 798.6000 922.8000 800.1000 924.0000 ;
	    RECT 808.2000 923.5500 934.2000 924.4500 ;
	    RECT 935.4000 924.0000 936.6000 929.7000 ;
	    RECT 808.2000 923.4000 809.4000 923.5500 ;
	    RECT 933.0000 923.4000 934.2000 923.5500 ;
	    RECT 796.2000 921.0000 798.0000 921.9000 ;
	    RECT 790.5000 918.9000 796.2000 920.1000 ;
	    RECT 752.7000 918.0000 753.9000 918.3000 ;
	    RECT 752.7000 917.1000 759.3000 918.0000 ;
	    RECT 760.2000 917.4000 761.4000 918.6000 ;
	    RECT 786.6000 918.0000 787.8000 918.9000 ;
	    RECT 797.1000 918.0000 798.0000 921.0000 ;
	    RECT 762.3000 917.1000 787.8000 918.0000 ;
	    RECT 796.8000 917.1000 798.0000 918.0000 ;
	    RECT 794.7000 916.2000 795.9000 916.5000 ;
	    RECT 755.4000 914.4000 756.6000 915.6000 ;
	    RECT 757.5000 915.3000 795.9000 916.2000 ;
	    RECT 760.5000 915.0000 761.7000 915.3000 ;
	    RECT 796.8000 914.4000 797.7000 917.1000 ;
	    RECT 798.9000 916.2000 800.1000 922.8000 ;
	    RECT 765.0000 914.1000 766.2000 914.4000 ;
	    RECT 758.1000 913.5000 766.2000 914.1000 ;
	    RECT 756.9000 913.2000 766.2000 913.5000 ;
	    RECT 767.7000 913.5000 780.6000 914.4000 ;
	    RECT 753.0000 912.0000 755.4000 913.2000 ;
	    RECT 756.9000 912.3000 759.0000 913.2000 ;
	    RECT 767.7000 912.3000 768.6000 913.5000 ;
	    RECT 779.4000 913.2000 780.6000 913.5000 ;
	    RECT 784.2000 913.5000 797.7000 914.4000 ;
	    RECT 798.6000 915.0000 800.1000 916.2000 ;
	    RECT 935.1000 922.8000 936.6000 924.0000 ;
	    RECT 935.1000 916.2000 936.3000 922.8000 ;
	    RECT 937.8000 921.9000 939.0000 929.7000 ;
	    RECT 942.6000 923.7000 943.8000 929.7000 ;
	    RECT 947.4000 924.9000 948.6000 929.7000 ;
	    RECT 949.8000 925.5000 951.0000 929.7000 ;
	    RECT 952.2000 925.5000 953.4000 929.7000 ;
	    RECT 954.6000 925.5000 955.8000 929.7000 ;
	    RECT 957.0000 925.5000 958.2000 929.7000 ;
	    RECT 959.4000 926.7000 960.6000 929.7000 ;
	    RECT 961.8000 925.5000 963.0000 929.7000 ;
	    RECT 964.2000 926.7000 965.4000 929.7000 ;
	    RECT 966.6000 925.5000 967.8000 929.7000 ;
	    RECT 969.0000 925.5000 970.2000 929.7000 ;
	    RECT 971.4000 925.5000 972.6000 929.7000 ;
	    RECT 945.0000 923.7000 948.6000 924.9000 ;
	    RECT 973.8000 924.9000 975.0000 929.7000 ;
	    RECT 945.0000 922.8000 946.2000 923.7000 ;
	    RECT 937.2000 921.0000 939.0000 921.9000 ;
	    RECT 943.5000 921.9000 946.2000 922.8000 ;
	    RECT 952.2000 923.4000 953.7000 924.6000 ;
	    RECT 958.2000 923.4000 958.5000 924.6000 ;
	    RECT 959.4000 923.4000 960.6000 924.6000 ;
	    RECT 961.8000 923.7000 968.7000 924.6000 ;
	    RECT 973.8000 923.7000 977.7000 924.9000 ;
	    RECT 978.6000 923.7000 979.8000 929.7000 ;
	    RECT 961.8000 923.4000 963.0000 923.7000 ;
	    RECT 937.2000 918.0000 938.1000 921.0000 ;
	    RECT 943.5000 920.1000 944.7000 921.9000 ;
	    RECT 939.0000 918.9000 944.7000 920.1000 ;
	    RECT 952.2000 919.2000 953.4000 923.4000 ;
	    RECT 964.2000 922.5000 965.4000 922.8000 ;
	    RECT 961.8000 922.2000 963.0000 922.5000 ;
	    RECT 956.4000 921.3000 963.0000 922.2000 ;
	    RECT 956.4000 921.0000 957.6000 921.3000 ;
	    RECT 964.2000 920.4000 965.4000 921.6000 ;
	    RECT 967.5000 920.1000 968.7000 923.7000 ;
	    RECT 976.5000 922.8000 977.7000 923.7000 ;
	    RECT 976.5000 921.6000 981.0000 922.8000 ;
	    RECT 983.4000 920.7000 984.6000 929.7000 ;
	    RECT 1115.4000 926.7000 1116.6000 929.7000 ;
	    RECT 1117.8000 924.0000 1119.0000 929.7000 ;
	    RECT 957.0000 918.9000 961.8000 920.1000 ;
	    RECT 967.5000 918.9000 970.5000 920.1000 ;
	    RECT 971.4000 919.5000 984.6000 920.7000 ;
	    RECT 947.4000 918.0000 948.6000 918.9000 ;
	    RECT 937.2000 917.1000 938.4000 918.0000 ;
	    RECT 947.4000 917.1000 972.9000 918.0000 ;
	    RECT 973.8000 917.4000 975.0000 918.6000 ;
	    RECT 981.3000 918.0000 982.5000 918.3000 ;
	    RECT 975.9000 917.1000 982.5000 918.0000 ;
	    RECT 858.6000 915.4500 859.8000 915.6000 ;
	    RECT 899.4000 915.4500 900.6000 915.6000 ;
	    RECT 798.6000 913.5000 799.8000 915.0000 ;
	    RECT 858.6000 914.5500 900.6000 915.4500 ;
	    RECT 935.1000 915.0000 936.6000 916.2000 ;
	    RECT 858.6000 914.4000 859.8000 914.5500 ;
	    RECT 899.4000 914.4000 900.6000 914.5500 ;
	    RECT 935.4000 913.5000 936.6000 915.0000 ;
	    RECT 937.5000 914.4000 938.4000 917.1000 ;
	    RECT 939.3000 916.2000 940.5000 916.5000 ;
	    RECT 939.3000 915.3000 977.7000 916.2000 ;
	    RECT 973.5000 915.0000 974.7000 915.3000 ;
	    RECT 978.6000 914.4000 979.8000 915.6000 ;
	    RECT 937.5000 913.5000 951.0000 914.4000 ;
	    RECT 784.2000 913.2000 785.4000 913.5000 ;
	    RECT 754.5000 911.4000 755.4000 912.0000 ;
	    RECT 759.9000 911.4000 768.6000 912.3000 ;
	    RECT 769.5000 911.4000 773.4000 912.6000 ;
	    RECT 750.6000 910.2000 753.6000 911.1000 ;
	    RECT 754.5000 910.2000 760.8000 911.4000 ;
	    RECT 752.7000 909.3000 753.6000 910.2000 ;
	    RECT 618.6000 903.3000 619.8000 909.3000 ;
	    RECT 750.6000 903.3000 751.8000 909.3000 ;
	    RECT 752.7000 908.4000 754.2000 909.3000 ;
	    RECT 753.0000 903.3000 754.2000 908.4000 ;
	    RECT 755.4000 902.4000 756.6000 909.3000 ;
	    RECT 757.8000 903.3000 759.0000 910.2000 ;
	    RECT 760.2000 903.3000 761.4000 909.3000 ;
	    RECT 762.6000 903.3000 763.8000 907.5000 ;
	    RECT 765.0000 903.3000 766.2000 907.5000 ;
	    RECT 767.4000 903.3000 768.6000 910.5000 ;
	    RECT 769.8000 903.3000 771.0000 909.3000 ;
	    RECT 772.2000 903.3000 773.4000 910.5000 ;
	    RECT 774.6000 903.3000 775.8000 909.3000 ;
	    RECT 777.0000 903.3000 778.2000 912.6000 ;
	    RECT 789.0000 911.4000 792.9000 912.6000 ;
	    RECT 781.8000 910.2000 788.1000 911.4000 ;
	    RECT 779.4000 903.3000 780.6000 907.5000 ;
	    RECT 781.8000 903.3000 783.0000 907.5000 ;
	    RECT 784.2000 903.3000 785.4000 907.5000 ;
	    RECT 786.6000 903.3000 787.8000 909.3000 ;
	    RECT 789.0000 903.3000 790.2000 911.4000 ;
	    RECT 796.8000 911.1000 797.7000 913.5000 ;
	    RECT 798.6000 911.4000 799.8000 912.6000 ;
	    RECT 846.6000 912.4500 847.8000 912.6000 ;
	    RECT 921.0000 912.4500 922.2000 912.6000 ;
	    RECT 935.4000 912.4500 936.6000 912.6000 ;
	    RECT 846.6000 911.5500 936.6000 912.4500 ;
	    RECT 846.6000 911.4000 847.8000 911.5500 ;
	    RECT 921.0000 911.4000 922.2000 911.5500 ;
	    RECT 935.4000 911.4000 936.6000 911.5500 ;
	    RECT 793.8000 910.2000 797.7000 911.1000 ;
	    RECT 937.5000 911.1000 938.4000 913.5000 ;
	    RECT 949.8000 913.2000 951.0000 913.5000 ;
	    RECT 954.6000 913.5000 967.5000 914.4000 ;
	    RECT 954.6000 913.2000 955.8000 913.5000 ;
	    RECT 942.3000 911.4000 946.2000 912.6000 ;
	    RECT 791.4000 903.3000 792.6000 909.3000 ;
	    RECT 793.8000 903.3000 795.0000 910.2000 ;
	    RECT 796.2000 903.3000 797.4000 909.3000 ;
	    RECT 798.6000 903.3000 799.8000 910.5000 ;
	    RECT 801.0000 903.3000 802.2000 909.3000 ;
	    RECT 933.0000 903.3000 934.2000 909.3000 ;
	    RECT 935.4000 903.3000 936.6000 910.5000 ;
	    RECT 937.5000 910.2000 941.4000 911.1000 ;
	    RECT 937.8000 903.3000 939.0000 909.3000 ;
	    RECT 940.2000 903.3000 941.4000 910.2000 ;
	    RECT 942.6000 903.3000 943.8000 909.3000 ;
	    RECT 945.0000 903.3000 946.2000 911.4000 ;
	    RECT 947.1000 910.2000 953.4000 911.4000 ;
	    RECT 947.4000 903.3000 948.6000 909.3000 ;
	    RECT 949.8000 903.3000 951.0000 907.5000 ;
	    RECT 952.2000 903.3000 953.4000 907.5000 ;
	    RECT 954.6000 903.3000 955.8000 907.5000 ;
	    RECT 957.0000 903.3000 958.2000 912.6000 ;
	    RECT 961.8000 911.4000 965.7000 912.6000 ;
	    RECT 966.6000 912.3000 967.5000 913.5000 ;
	    RECT 969.0000 914.1000 970.2000 914.4000 ;
	    RECT 969.0000 913.5000 977.1000 914.1000 ;
	    RECT 969.0000 913.2000 978.3000 913.5000 ;
	    RECT 976.2000 912.3000 978.3000 913.2000 ;
	    RECT 966.6000 911.4000 975.3000 912.3000 ;
	    RECT 979.8000 912.0000 982.2000 913.2000 ;
	    RECT 979.8000 911.4000 980.7000 912.0000 ;
	    RECT 959.4000 903.3000 960.6000 909.3000 ;
	    RECT 961.8000 903.3000 963.0000 910.5000 ;
	    RECT 964.2000 903.3000 965.4000 909.3000 ;
	    RECT 966.6000 903.3000 967.8000 910.5000 ;
	    RECT 974.4000 910.2000 980.7000 911.4000 ;
	    RECT 983.4000 911.1000 984.6000 919.5000 ;
	    RECT 1117.5000 922.8000 1119.0000 924.0000 ;
	    RECT 1117.5000 916.2000 1118.7001 922.8000 ;
	    RECT 1120.2001 921.9000 1121.4000 929.7000 ;
	    RECT 1125.0000 923.7000 1126.2001 929.7000 ;
	    RECT 1129.8000 924.9000 1131.0000 929.7000 ;
	    RECT 1132.2001 925.5000 1133.4000 929.7000 ;
	    RECT 1134.6000 925.5000 1135.8000 929.7000 ;
	    RECT 1137.0000 925.5000 1138.2001 929.7000 ;
	    RECT 1139.4000 925.5000 1140.6000 929.7000 ;
	    RECT 1141.8000 926.7000 1143.0000 929.7000 ;
	    RECT 1144.2001 925.5000 1145.4000 929.7000 ;
	    RECT 1146.6000 926.7000 1147.8000 929.7000 ;
	    RECT 1149.0000 925.5000 1150.2001 929.7000 ;
	    RECT 1151.4000 925.5000 1152.6000 929.7000 ;
	    RECT 1153.8000 925.5000 1155.0000 929.7000 ;
	    RECT 1127.4000 923.7000 1131.0000 924.9000 ;
	    RECT 1156.2001 924.9000 1157.4000 929.7000 ;
	    RECT 1127.4000 922.8000 1128.6000 923.7000 ;
	    RECT 1119.6000 921.0000 1121.4000 921.9000 ;
	    RECT 1125.9000 921.9000 1128.6000 922.8000 ;
	    RECT 1134.6000 923.4000 1136.1000 924.6000 ;
	    RECT 1140.6000 923.4000 1140.9000 924.6000 ;
	    RECT 1141.8000 923.4000 1143.0000 924.6000 ;
	    RECT 1144.2001 923.7000 1151.1000 924.6000 ;
	    RECT 1156.2001 923.7000 1160.1000 924.9000 ;
	    RECT 1161.0000 923.7000 1162.2001 929.7000 ;
	    RECT 1144.2001 923.4000 1145.4000 923.7000 ;
	    RECT 1119.6000 918.0000 1120.5000 921.0000 ;
	    RECT 1125.9000 920.1000 1127.1000 921.9000 ;
	    RECT 1121.4000 918.9000 1127.1000 920.1000 ;
	    RECT 1134.6000 919.2000 1135.8000 923.4000 ;
	    RECT 1146.6000 922.5000 1147.8000 922.8000 ;
	    RECT 1144.2001 922.2000 1145.4000 922.5000 ;
	    RECT 1138.8000 921.3000 1145.4000 922.2000 ;
	    RECT 1138.8000 921.0000 1140.0000 921.3000 ;
	    RECT 1146.6000 920.4000 1147.8000 921.6000 ;
	    RECT 1149.9000 920.1000 1151.1000 923.7000 ;
	    RECT 1158.9000 922.8000 1160.1000 923.7000 ;
	    RECT 1158.9000 921.6000 1163.4000 922.8000 ;
	    RECT 1165.8000 920.7000 1167.0000 929.7000 ;
	    RECT 1290.6000 926.7000 1291.8000 929.7000 ;
	    RECT 1293.0000 924.0000 1294.2001 929.7000 ;
	    RECT 1139.4000 918.9000 1144.2001 920.1000 ;
	    RECT 1149.9000 918.9000 1152.9000 920.1000 ;
	    RECT 1153.8000 919.5000 1167.0000 920.7000 ;
	    RECT 1129.8000 918.0000 1131.0000 918.9000 ;
	    RECT 1119.6000 917.1000 1120.8000 918.0000 ;
	    RECT 1129.8000 917.1000 1155.3000 918.0000 ;
	    RECT 1156.2001 917.4000 1157.4000 918.6000 ;
	    RECT 1163.7001 918.0000 1164.9000 918.3000 ;
	    RECT 1158.3000 917.1000 1164.9000 918.0000 ;
	    RECT 1117.5000 915.0000 1119.0000 916.2000 ;
	    RECT 1117.8000 913.5000 1119.0000 915.0000 ;
	    RECT 1119.9000 914.4000 1120.8000 917.1000 ;
	    RECT 1121.7001 916.2000 1122.9000 916.5000 ;
	    RECT 1121.7001 915.3000 1160.1000 916.2000 ;
	    RECT 1155.9000 915.0000 1157.1000 915.3000 ;
	    RECT 1161.0000 914.4000 1162.2001 915.6000 ;
	    RECT 1119.9000 913.5000 1133.4000 914.4000 ;
	    RECT 997.8000 912.4500 999.0000 912.6000 ;
	    RECT 1043.4000 912.4500 1044.6000 912.6000 ;
	    RECT 1117.8000 912.4500 1119.0000 912.6000 ;
	    RECT 997.8000 911.5500 1119.0000 912.4500 ;
	    RECT 997.8000 911.4000 999.0000 911.5500 ;
	    RECT 1043.4000 911.4000 1044.6000 911.5500 ;
	    RECT 1117.8000 911.4000 1119.0000 911.5500 ;
	    RECT 981.6000 910.2000 984.6000 911.1000 ;
	    RECT 1119.9000 911.1000 1120.8000 913.5000 ;
	    RECT 1132.2001 913.2000 1133.4000 913.5000 ;
	    RECT 1137.0000 913.5000 1149.9000 914.4000 ;
	    RECT 1137.0000 913.2000 1138.2001 913.5000 ;
	    RECT 1124.7001 911.4000 1128.6000 912.6000 ;
	    RECT 969.0000 903.3000 970.2000 907.5000 ;
	    RECT 971.4000 903.3000 972.6000 907.5000 ;
	    RECT 973.8000 903.3000 975.0000 909.3000 ;
	    RECT 976.2000 903.3000 977.4000 910.2000 ;
	    RECT 981.6000 909.3000 982.5000 910.2000 ;
	    RECT 978.6000 902.4000 979.8000 909.3000 ;
	    RECT 981.0000 908.4000 982.5000 909.3000 ;
	    RECT 981.0000 903.3000 982.2000 908.4000 ;
	    RECT 983.4000 903.3000 984.6000 909.3000 ;
	    RECT 1115.4000 903.3000 1116.6000 909.3000 ;
	    RECT 1117.8000 903.3000 1119.0000 910.5000 ;
	    RECT 1119.9000 910.2000 1123.8000 911.1000 ;
	    RECT 1120.2001 903.3000 1121.4000 909.3000 ;
	    RECT 1122.6000 903.3000 1123.8000 910.2000 ;
	    RECT 1125.0000 903.3000 1126.2001 909.3000 ;
	    RECT 1127.4000 903.3000 1128.6000 911.4000 ;
	    RECT 1129.5000 910.2000 1135.8000 911.4000 ;
	    RECT 1129.8000 903.3000 1131.0000 909.3000 ;
	    RECT 1132.2001 903.3000 1133.4000 907.5000 ;
	    RECT 1134.6000 903.3000 1135.8000 907.5000 ;
	    RECT 1137.0000 903.3000 1138.2001 907.5000 ;
	    RECT 1139.4000 903.3000 1140.6000 912.6000 ;
	    RECT 1144.2001 911.4000 1148.1000 912.6000 ;
	    RECT 1149.0000 912.3000 1149.9000 913.5000 ;
	    RECT 1151.4000 914.1000 1152.6000 914.4000 ;
	    RECT 1151.4000 913.5000 1159.5000 914.1000 ;
	    RECT 1151.4000 913.2000 1160.7001 913.5000 ;
	    RECT 1158.6000 912.3000 1160.7001 913.2000 ;
	    RECT 1149.0000 911.4000 1157.7001 912.3000 ;
	    RECT 1162.2001 912.0000 1164.6000 913.2000 ;
	    RECT 1162.2001 911.4000 1163.1000 912.0000 ;
	    RECT 1141.8000 903.3000 1143.0000 909.3000 ;
	    RECT 1144.2001 903.3000 1145.4000 910.5000 ;
	    RECT 1146.6000 903.3000 1147.8000 909.3000 ;
	    RECT 1149.0000 903.3000 1150.2001 910.5000 ;
	    RECT 1156.8000 910.2000 1163.1000 911.4000 ;
	    RECT 1165.8000 911.1000 1167.0000 919.5000 ;
	    RECT 1292.7001 922.8000 1294.2001 924.0000 ;
	    RECT 1292.7001 916.2000 1293.9000 922.8000 ;
	    RECT 1295.4000 921.9000 1296.6000 929.7000 ;
	    RECT 1300.2001 923.7000 1301.4000 929.7000 ;
	    RECT 1305.0000 924.9000 1306.2001 929.7000 ;
	    RECT 1307.4000 925.5000 1308.6000 929.7000 ;
	    RECT 1309.8000 925.5000 1311.0000 929.7000 ;
	    RECT 1312.2001 925.5000 1313.4000 929.7000 ;
	    RECT 1314.6000 925.5000 1315.8000 929.7000 ;
	    RECT 1317.0000 926.7000 1318.2001 929.7000 ;
	    RECT 1319.4000 925.5000 1320.6000 929.7000 ;
	    RECT 1321.8000 926.7000 1323.0000 929.7000 ;
	    RECT 1324.2001 925.5000 1325.4000 929.7000 ;
	    RECT 1326.6000 925.5000 1327.8000 929.7000 ;
	    RECT 1329.0000 925.5000 1330.2001 929.7000 ;
	    RECT 1302.6000 923.7000 1306.2001 924.9000 ;
	    RECT 1331.4000 924.9000 1332.6000 929.7000 ;
	    RECT 1302.6000 922.8000 1303.8000 923.7000 ;
	    RECT 1294.8000 921.0000 1296.6000 921.9000 ;
	    RECT 1301.1000 921.9000 1303.8000 922.8000 ;
	    RECT 1309.8000 923.4000 1311.3000 924.6000 ;
	    RECT 1315.8000 923.4000 1316.1000 924.6000 ;
	    RECT 1317.0000 923.4000 1318.2001 924.6000 ;
	    RECT 1319.4000 923.7000 1326.3000 924.6000 ;
	    RECT 1331.4000 923.7000 1335.3000 924.9000 ;
	    RECT 1336.2001 923.7000 1337.4000 929.7000 ;
	    RECT 1319.4000 923.4000 1320.6000 923.7000 ;
	    RECT 1294.8000 918.0000 1295.7001 921.0000 ;
	    RECT 1301.1000 920.1000 1302.3000 921.9000 ;
	    RECT 1296.6000 918.9000 1302.3000 920.1000 ;
	    RECT 1309.8000 919.2000 1311.0000 923.4000 ;
	    RECT 1321.8000 922.5000 1323.0000 922.8000 ;
	    RECT 1319.4000 922.2000 1320.6000 922.5000 ;
	    RECT 1314.0000 921.3000 1320.6000 922.2000 ;
	    RECT 1314.0000 921.0000 1315.2001 921.3000 ;
	    RECT 1321.8000 920.4000 1323.0000 921.6000 ;
	    RECT 1325.1000 920.1000 1326.3000 923.7000 ;
	    RECT 1334.1000 922.8000 1335.3000 923.7000 ;
	    RECT 1334.1000 921.6000 1338.6000 922.8000 ;
	    RECT 1341.0000 920.7000 1342.2001 929.7000 ;
	    RECT 1367.4000 922.8000 1368.6000 929.7000 ;
	    RECT 1369.8000 923.7000 1371.0000 929.7000 ;
	    RECT 1367.4000 921.9000 1370.7001 922.8000 ;
	    RECT 1372.2001 922.5000 1373.4000 929.7000 ;
	    RECT 1386.6000 922.5000 1387.8000 929.7000 ;
	    RECT 1389.0000 926.7000 1390.2001 929.7000 ;
	    RECT 1389.0000 925.5000 1390.2001 925.8000 ;
	    RECT 1389.0000 923.4000 1390.2001 924.6000 ;
	    RECT 1408.2001 922.8000 1409.4000 929.7000 ;
	    RECT 1410.6000 923.7000 1411.8000 929.7000 ;
	    RECT 1408.2001 921.9000 1411.5000 922.8000 ;
	    RECT 1413.0000 922.5000 1414.2001 929.7000 ;
	    RECT 1427.4000 922.5000 1428.6000 929.7000 ;
	    RECT 1429.8000 926.7000 1431.0000 929.7000 ;
	    RECT 1441.8000 926.7000 1443.0000 929.7000 ;
	    RECT 1429.8000 925.5000 1431.0000 925.8000 ;
	    RECT 1441.8000 925.5000 1443.0000 925.8000 ;
	    RECT 1429.8000 923.4000 1431.0000 924.6000 ;
	    RECT 1441.8000 923.4000 1443.0000 924.6000 ;
	    RECT 1444.2001 922.5000 1445.4000 929.7000 ;
	    RECT 1456.2001 926.7000 1457.4000 929.7000 ;
	    RECT 1456.2001 925.5000 1457.4000 925.8000 ;
	    RECT 1456.2001 923.4000 1457.4000 924.6000 ;
	    RECT 1458.6000 922.5000 1459.8000 929.7000 ;
	    RECT 1482.6000 924.0000 1483.8000 929.7000 ;
	    RECT 1485.0000 924.9000 1486.2001 929.7000 ;
	    RECT 1487.4000 924.0000 1488.6000 929.7000 ;
	    RECT 1482.6000 923.7000 1488.6000 924.0000 ;
	    RECT 1489.8000 923.7000 1491.0000 929.7000 ;
	    RECT 1497.0000 924.4500 1498.2001 924.6000 ;
	    RECT 1501.8000 924.4500 1503.0000 924.6000 ;
	    RECT 1482.9000 923.1000 1488.3000 923.7000 ;
	    RECT 1489.8000 922.5000 1490.7001 923.7000 ;
	    RECT 1497.0000 923.5500 1503.0000 924.4500 ;
	    RECT 1497.0000 923.4000 1498.2001 923.5500 ;
	    RECT 1501.8000 923.4000 1503.0000 923.5500 ;
	    RECT 1504.2001 922.5000 1505.4000 929.7000 ;
	    RECT 1506.6000 926.7000 1507.8000 929.7000 ;
	    RECT 1506.6000 925.5000 1507.8000 925.8000 ;
	    RECT 1506.6000 924.4500 1507.8000 924.6000 ;
	    RECT 1530.6000 924.4500 1531.8000 924.6000 ;
	    RECT 1506.6000 923.5500 1531.8000 924.4500 ;
	    RECT 1533.0000 924.0000 1534.2001 929.7000 ;
	    RECT 1535.4000 924.9000 1536.6000 929.7000 ;
	    RECT 1537.8000 924.0000 1539.0000 929.7000 ;
	    RECT 1533.0000 923.7000 1539.0000 924.0000 ;
	    RECT 1540.2001 923.7000 1541.4000 929.7000 ;
	    RECT 1559.4000 923.7000 1560.6000 929.7000 ;
	    RECT 1563.3000 924.6000 1564.5000 929.7000 ;
	    RECT 1561.8000 923.7000 1564.5000 924.6000 ;
	    RECT 1506.6000 923.4000 1507.8000 923.5500 ;
	    RECT 1530.6000 923.4000 1531.8000 923.5500 ;
	    RECT 1533.3000 923.1000 1538.7001 923.7000 ;
	    RECT 1540.2001 922.5000 1541.1000 923.7000 ;
	    RECT 1559.4000 922.5000 1560.6000 922.8000 ;
	    RECT 1314.6000 918.9000 1319.4000 920.1000 ;
	    RECT 1325.1000 918.9000 1328.1000 920.1000 ;
	    RECT 1329.0000 919.5000 1342.2001 920.7000 ;
	    RECT 1367.4000 919.5000 1368.6000 919.8000 ;
	    RECT 1305.0000 918.0000 1306.2001 918.9000 ;
	    RECT 1294.8000 917.1000 1296.0000 918.0000 ;
	    RECT 1305.0000 917.1000 1330.5000 918.0000 ;
	    RECT 1331.4000 917.4000 1332.6000 918.6000 ;
	    RECT 1338.9000 918.0000 1340.1000 918.3000 ;
	    RECT 1333.5000 917.1000 1340.1000 918.0000 ;
	    RECT 1292.7001 915.0000 1294.2001 916.2000 ;
	    RECT 1293.0000 913.5000 1294.2001 915.0000 ;
	    RECT 1295.1000 914.4000 1296.0000 917.1000 ;
	    RECT 1296.9000 916.2000 1298.1000 916.5000 ;
	    RECT 1296.9000 915.3000 1335.3000 916.2000 ;
	    RECT 1331.1000 915.0000 1332.3000 915.3000 ;
	    RECT 1336.2001 914.4000 1337.4000 915.6000 ;
	    RECT 1295.1000 913.5000 1308.6000 914.4000 ;
	    RECT 1261.8000 912.4500 1263.0000 912.6000 ;
	    RECT 1293.0000 912.4500 1294.2001 912.6000 ;
	    RECT 1261.8000 911.5500 1294.2001 912.4500 ;
	    RECT 1261.8000 911.4000 1263.0000 911.5500 ;
	    RECT 1293.0000 911.4000 1294.2001 911.5500 ;
	    RECT 1164.0000 910.2000 1167.0000 911.1000 ;
	    RECT 1295.1000 911.1000 1296.0000 913.5000 ;
	    RECT 1307.4000 913.2000 1308.6000 913.5000 ;
	    RECT 1312.2001 913.5000 1325.1000 914.4000 ;
	    RECT 1312.2001 913.2000 1313.4000 913.5000 ;
	    RECT 1299.9000 911.4000 1303.8000 912.6000 ;
	    RECT 1151.4000 903.3000 1152.6000 907.5000 ;
	    RECT 1153.8000 903.3000 1155.0000 907.5000 ;
	    RECT 1156.2001 903.3000 1157.4000 909.3000 ;
	    RECT 1158.6000 903.3000 1159.8000 910.2000 ;
	    RECT 1164.0000 909.3000 1164.9000 910.2000 ;
	    RECT 1161.0000 902.4000 1162.2001 909.3000 ;
	    RECT 1163.4000 908.4000 1164.9000 909.3000 ;
	    RECT 1163.4000 903.3000 1164.6000 908.4000 ;
	    RECT 1165.8000 903.3000 1167.0000 909.3000 ;
	    RECT 1290.6000 903.3000 1291.8000 909.3000 ;
	    RECT 1293.0000 903.3000 1294.2001 910.5000 ;
	    RECT 1295.1000 910.2000 1299.0000 911.1000 ;
	    RECT 1295.4000 903.3000 1296.6000 909.3000 ;
	    RECT 1297.8000 903.3000 1299.0000 910.2000 ;
	    RECT 1300.2001 903.3000 1301.4000 909.3000 ;
	    RECT 1302.6000 903.3000 1303.8000 911.4000 ;
	    RECT 1304.7001 910.2000 1311.0000 911.4000 ;
	    RECT 1305.0000 903.3000 1306.2001 909.3000 ;
	    RECT 1307.4000 903.3000 1308.6000 907.5000 ;
	    RECT 1309.8000 903.3000 1311.0000 907.5000 ;
	    RECT 1312.2001 903.3000 1313.4000 907.5000 ;
	    RECT 1314.6000 903.3000 1315.8000 912.6000 ;
	    RECT 1319.4000 911.4000 1323.3000 912.6000 ;
	    RECT 1324.2001 912.3000 1325.1000 913.5000 ;
	    RECT 1326.6000 914.1000 1327.8000 914.4000 ;
	    RECT 1326.6000 913.5000 1334.7001 914.1000 ;
	    RECT 1326.6000 913.2000 1335.9000 913.5000 ;
	    RECT 1333.8000 912.3000 1335.9000 913.2000 ;
	    RECT 1324.2001 911.4000 1332.9000 912.3000 ;
	    RECT 1337.4000 912.0000 1339.8000 913.2000 ;
	    RECT 1337.4000 911.4000 1338.3000 912.0000 ;
	    RECT 1317.0000 903.3000 1318.2001 909.3000 ;
	    RECT 1319.4000 903.3000 1320.6000 910.5000 ;
	    RECT 1321.8000 903.3000 1323.0000 909.3000 ;
	    RECT 1324.2001 903.3000 1325.4000 910.5000 ;
	    RECT 1332.0000 910.2000 1338.3000 911.4000 ;
	    RECT 1341.0000 911.1000 1342.2001 919.5000 ;
	    RECT 1367.4000 917.4000 1368.6000 918.6000 ;
	    RECT 1369.8000 917.4000 1370.7001 921.9000 ;
	    RECT 1372.2001 921.4500 1373.4000 921.6000 ;
	    RECT 1374.6000 921.4500 1375.8000 921.6000 ;
	    RECT 1372.2001 920.5500 1375.8000 921.4500 ;
	    RECT 1372.2001 920.4000 1373.4000 920.5500 ;
	    RECT 1374.6000 920.4000 1375.8000 920.5500 ;
	    RECT 1377.0000 921.4500 1378.2001 921.6000 ;
	    RECT 1386.6000 921.4500 1387.8000 921.6000 ;
	    RECT 1377.0000 920.5500 1387.8000 921.4500 ;
	    RECT 1377.0000 920.4000 1378.2001 920.5500 ;
	    RECT 1386.6000 920.4000 1387.8000 920.5500 ;
	    RECT 1408.2001 919.5000 1409.4000 919.8000 ;
	    RECT 1372.2001 918.6000 1373.4000 919.5000 ;
	    RECT 1369.8000 916.2000 1371.6000 917.4000 ;
	    RECT 1369.8000 915.3000 1370.7001 916.2000 ;
	    RECT 1372.5000 915.3000 1373.4000 918.6000 ;
	    RECT 1339.2001 910.2000 1342.2001 911.1000 ;
	    RECT 1367.4000 914.4000 1370.7001 915.3000 ;
	    RECT 1326.6000 903.3000 1327.8000 907.5000 ;
	    RECT 1329.0000 903.3000 1330.2001 907.5000 ;
	    RECT 1331.4000 903.3000 1332.6000 909.3000 ;
	    RECT 1333.8000 903.3000 1335.0000 910.2000 ;
	    RECT 1339.2001 909.3000 1340.1000 910.2000 ;
	    RECT 1336.2001 902.4000 1337.4000 909.3000 ;
	    RECT 1338.6000 908.4000 1340.1000 909.3000 ;
	    RECT 1338.6000 903.3000 1339.8000 908.4000 ;
	    RECT 1341.0000 903.3000 1342.2001 909.3000 ;
	    RECT 1367.4000 903.3000 1368.6000 914.4000 ;
	    RECT 1369.8000 903.3000 1371.0000 913.5000 ;
	    RECT 1372.2001 903.3000 1373.4000 915.3000 ;
	    RECT 1386.6000 903.3000 1387.8000 919.5000 ;
	    RECT 1408.2001 917.4000 1409.4000 918.6000 ;
	    RECT 1410.6000 917.4000 1411.5000 921.9000 ;
	    RECT 1413.0000 920.4000 1414.2001 921.6000 ;
	    RECT 1417.8000 921.4500 1419.0000 921.6000 ;
	    RECT 1427.4000 921.4500 1428.6000 921.6000 ;
	    RECT 1417.8000 920.5500 1428.6000 921.4500 ;
	    RECT 1417.8000 920.4000 1419.0000 920.5500 ;
	    RECT 1427.4000 920.4000 1428.6000 920.5500 ;
	    RECT 1432.2001 921.4500 1433.4000 921.6000 ;
	    RECT 1444.2001 921.4500 1445.4000 921.6000 ;
	    RECT 1432.2001 920.5500 1445.4000 921.4500 ;
	    RECT 1432.2001 920.4000 1433.4000 920.5500 ;
	    RECT 1444.2001 920.4000 1445.4000 920.5500 ;
	    RECT 1458.6000 921.4500 1459.8000 921.6000 ;
	    RECT 1477.8000 921.4500 1479.0000 921.6000 ;
	    RECT 1458.6000 920.5500 1479.0000 921.4500 ;
	    RECT 1458.6000 920.4000 1459.8000 920.5500 ;
	    RECT 1477.8000 920.4000 1479.0000 920.5500 ;
	    RECT 1482.6000 920.4000 1483.8000 921.6000 ;
	    RECT 1484.7001 920.7000 1485.0000 922.2000 ;
	    RECT 1487.1000 920.4000 1488.9000 921.6000 ;
	    RECT 1489.8000 920.4000 1491.0000 921.6000 ;
	    RECT 1492.2001 921.4500 1493.4000 921.6000 ;
	    RECT 1504.2001 921.4500 1505.4000 921.6000 ;
	    RECT 1492.2001 920.5500 1505.4000 921.4500 ;
	    RECT 1492.2001 920.4000 1493.4000 920.5500 ;
	    RECT 1504.2001 920.4000 1505.4000 920.5500 ;
	    RECT 1518.6000 921.4500 1519.8000 921.6000 ;
	    RECT 1533.0000 921.4500 1534.2001 921.6000 ;
	    RECT 1518.6000 920.5500 1534.2001 921.4500 ;
	    RECT 1535.1000 920.7000 1535.4000 922.2000 ;
	    RECT 1518.6000 920.4000 1519.8000 920.5500 ;
	    RECT 1533.0000 920.4000 1534.2001 920.5500 ;
	    RECT 1537.5000 920.4000 1539.3000 921.6000 ;
	    RECT 1540.2001 921.4500 1541.4000 921.6000 ;
	    RECT 1542.6000 921.4500 1543.8000 921.6000 ;
	    RECT 1540.2001 920.5500 1543.8000 921.4500 ;
	    RECT 1540.2001 920.4000 1541.4000 920.5500 ;
	    RECT 1542.6000 920.4000 1543.8000 920.5500 ;
	    RECT 1559.4000 920.4000 1560.6000 921.6000 ;
	    RECT 1485.0000 919.5000 1486.2001 919.8000 ;
	    RECT 1413.0000 918.6000 1414.2001 919.5000 ;
	    RECT 1410.6000 916.2000 1412.4000 917.4000 ;
	    RECT 1410.6000 915.3000 1411.5000 916.2000 ;
	    RECT 1413.3000 915.3000 1414.2001 918.6000 ;
	    RECT 1408.2001 914.4000 1411.5000 915.3000 ;
	    RECT 1389.0000 903.3000 1390.2001 909.3000 ;
	    RECT 1408.2001 903.3000 1409.4000 914.4000 ;
	    RECT 1410.6000 903.3000 1411.8000 913.5000 ;
	    RECT 1413.0000 903.3000 1414.2001 915.3000 ;
	    RECT 1427.4000 903.3000 1428.6000 919.5000 ;
	    RECT 1429.8000 903.3000 1431.0000 909.3000 ;
	    RECT 1441.8000 903.3000 1443.0000 909.3000 ;
	    RECT 1444.2001 903.3000 1445.4000 919.5000 ;
	    RECT 1456.2001 903.3000 1457.4000 909.3000 ;
	    RECT 1458.6000 903.3000 1459.8000 919.5000 ;
	    RECT 1485.0000 917.4000 1486.2001 918.6000 ;
	    RECT 1487.1000 915.3000 1488.0000 920.4000 ;
	    RECT 1489.9501 918.4500 1490.8500 920.4000 ;
	    RECT 1535.4000 919.5000 1536.6000 919.8000 ;
	    RECT 1501.8000 918.4500 1503.0000 918.6000 ;
	    RECT 1489.9501 917.5500 1503.0000 918.4500 ;
	    RECT 1501.8000 917.4000 1503.0000 917.5500 ;
	    RECT 1482.6000 903.3000 1483.8000 915.3000 ;
	    RECT 1486.5000 914.4000 1488.0000 915.3000 ;
	    RECT 1489.8000 914.4000 1491.0000 915.6000 ;
	    RECT 1486.5000 903.3000 1487.7001 914.4000 ;
	    RECT 1488.9000 912.6000 1489.8000 913.5000 ;
	    RECT 1488.6000 911.4000 1489.8000 912.6000 ;
	    RECT 1488.9000 903.3000 1490.1000 909.3000 ;
	    RECT 1504.2001 903.3000 1505.4000 919.5000 ;
	    RECT 1521.0000 918.4500 1522.2001 918.6000 ;
	    RECT 1533.0000 918.4500 1534.2001 918.6000 ;
	    RECT 1521.0000 917.5500 1534.2001 918.4500 ;
	    RECT 1521.0000 917.4000 1522.2001 917.5500 ;
	    RECT 1533.0000 917.4000 1534.2001 917.5500 ;
	    RECT 1535.4000 917.4000 1536.6000 918.6000 ;
	    RECT 1537.5000 915.3000 1538.4000 920.4000 ;
	    RECT 1561.8000 919.5000 1563.0000 923.7000 ;
	    RECT 1561.8000 918.4500 1563.0000 918.6000 ;
	    RECT 1540.3500 917.5500 1563.0000 918.4500 ;
	    RECT 1540.3500 915.6000 1541.2500 917.5500 ;
	    RECT 1561.8000 917.4000 1563.0000 917.5500 ;
	    RECT 1506.6000 903.3000 1507.8000 909.3000 ;
	    RECT 1533.0000 903.3000 1534.2001 915.3000 ;
	    RECT 1536.9000 914.4000 1538.4000 915.3000 ;
	    RECT 1540.2001 914.4000 1541.4000 915.6000 ;
	    RECT 1536.9000 903.3000 1538.1000 914.4000 ;
	    RECT 1539.3000 912.6000 1540.2001 913.5000 ;
	    RECT 1539.0000 911.4000 1540.2001 912.6000 ;
	    RECT 1539.3000 903.3000 1540.5000 909.3000 ;
	    RECT 1559.4000 903.3000 1560.6000 909.3000 ;
	    RECT 1561.8000 903.3000 1563.0000 916.5000 ;
	    RECT 1564.2001 913.2000 1565.4000 913.5000 ;
	    RECT 1564.2001 903.3000 1565.4000 909.3000 ;
	    RECT 1.2000 900.6000 1569.0000 902.4000 ;
	    RECT 52.2000 887.7000 53.4000 899.7000 ;
	    RECT 54.6000 886.8000 55.8000 899.7000 ;
	    RECT 57.0000 887.7000 58.2000 899.7000 ;
	    RECT 59.4000 886.8000 60.6000 899.7000 ;
	    RECT 61.8000 887.7000 63.0000 899.7000 ;
	    RECT 64.2000 886.8000 65.4000 899.7000 ;
	    RECT 66.6000 887.7000 67.8000 899.7000 ;
	    RECT 69.0000 886.8000 70.2000 899.7000 ;
	    RECT 71.4000 887.7000 72.6000 899.7000 ;
	    RECT 90.6000 893.7000 91.8000 899.7000 ;
	    RECT 90.6000 889.5000 91.8000 889.8000 ;
	    RECT 85.8000 888.4500 87.0000 888.6000 ;
	    RECT 90.6000 888.4500 91.8000 888.6000 ;
	    RECT 85.8000 887.5500 91.8000 888.4500 ;
	    RECT 85.8000 887.4000 87.0000 887.5500 ;
	    RECT 90.6000 887.4000 91.8000 887.5500 ;
	    RECT 54.6000 885.6000 57.3000 886.8000 ;
	    RECT 59.4000 885.6000 62.7000 886.8000 ;
	    RECT 64.2000 885.6000 67.5000 886.8000 ;
	    RECT 69.0000 886.5000 72.6000 886.8000 ;
	    RECT 93.0000 886.5000 94.2000 899.7000 ;
	    RECT 95.4000 893.7000 96.6000 899.7000 ;
	    RECT 109.8000 893.7000 111.0000 899.7000 ;
	    RECT 69.0000 885.6000 70.5000 886.5000 ;
	    RECT 56.1000 883.5000 57.3000 885.6000 ;
	    RECT 61.5000 883.5000 62.7000 885.6000 ;
	    RECT 66.3000 883.5000 67.5000 885.6000 ;
	    RECT 71.4000 885.4500 72.6000 885.6000 ;
	    RECT 78.6000 885.4500 79.8000 885.6000 ;
	    RECT 71.4000 884.5500 79.8000 885.4500 ;
	    RECT 71.4000 884.4000 72.6000 884.5500 ;
	    RECT 78.6000 884.4000 79.8000 884.5500 ;
	    RECT 88.2000 885.4500 89.4000 885.6000 ;
	    RECT 93.0000 885.4500 94.2000 885.6000 ;
	    RECT 88.2000 884.5500 94.2000 885.4500 ;
	    RECT 88.2000 884.4000 89.4000 884.5500 ;
	    RECT 93.0000 884.4000 94.2000 884.5500 ;
	    RECT 112.2000 883.5000 113.4000 899.7000 ;
	    RECT 126.6000 893.7000 127.8000 899.7000 ;
	    RECT 129.0000 883.5000 130.2000 899.7000 ;
	    RECT 141.0000 893.7000 142.2000 899.7000 ;
	    RECT 143.4000 883.5000 144.6000 899.7000 ;
	    RECT 168.3000 893.7000 169.5000 899.7000 ;
	    RECT 168.6000 890.4000 169.8000 891.6000 ;
	    RECT 168.6000 889.5000 169.5000 890.4000 ;
	    RECT 170.7000 888.6000 171.9000 899.7000 ;
	    RECT 167.4000 887.4000 168.6000 888.6000 ;
	    RECT 170.4000 887.7000 171.9000 888.6000 ;
	    RECT 174.6000 887.7000 175.8000 899.7000 ;
	    RECT 198.6000 897.4500 199.8000 897.6000 ;
	    RECT 237.0000 897.4500 238.2000 897.6000 ;
	    RECT 198.6000 896.5500 238.2000 897.4500 ;
	    RECT 198.6000 896.4000 199.8000 896.5500 ;
	    RECT 237.0000 896.4000 238.2000 896.5500 ;
	    RECT 306.6000 893.7000 307.8000 899.7000 ;
	    RECT 309.0000 892.5000 310.2000 899.7000 ;
	    RECT 311.4000 893.7000 312.6000 899.7000 ;
	    RECT 313.8000 892.8000 315.0000 899.7000 ;
	    RECT 316.2000 893.7000 317.4000 899.7000 ;
	    RECT 311.1000 891.9000 315.0000 892.8000 ;
	    RECT 239.4000 891.4500 240.6000 891.6000 ;
	    RECT 309.0000 891.4500 310.2000 891.6000 ;
	    RECT 239.4000 890.5500 310.2000 891.4500 ;
	    RECT 239.4000 890.4000 240.6000 890.5500 ;
	    RECT 309.0000 890.4000 310.2000 890.5500 ;
	    RECT 311.1000 889.5000 312.0000 891.9000 ;
	    RECT 318.6000 891.6000 319.8000 899.7000 ;
	    RECT 321.0000 893.7000 322.2000 899.7000 ;
	    RECT 323.4000 895.5000 324.6000 899.7000 ;
	    RECT 325.8000 895.5000 327.0000 899.7000 ;
	    RECT 328.2000 895.5000 329.4000 899.7000 ;
	    RECT 320.7000 891.6000 327.0000 892.8000 ;
	    RECT 315.9000 890.4000 319.8000 891.6000 ;
	    RECT 330.6000 890.4000 331.8000 899.7000 ;
	    RECT 333.0000 893.7000 334.2000 899.7000 ;
	    RECT 335.4000 892.5000 336.6000 899.7000 ;
	    RECT 337.8000 893.7000 339.0000 899.7000 ;
	    RECT 340.2000 892.5000 341.4000 899.7000 ;
	    RECT 342.6000 895.5000 343.8000 899.7000 ;
	    RECT 345.0000 895.5000 346.2000 899.7000 ;
	    RECT 347.4000 893.7000 348.6000 899.7000 ;
	    RECT 349.8000 892.8000 351.0000 899.7000 ;
	    RECT 352.2000 893.7000 353.4000 900.6000 ;
	    RECT 354.6000 894.6000 355.8000 899.7000 ;
	    RECT 354.6000 893.7000 356.1000 894.6000 ;
	    RECT 357.0000 893.7000 358.2000 899.7000 ;
	    RECT 369.0000 893.7000 370.2000 899.7000 ;
	    RECT 355.2000 892.8000 356.1000 893.7000 ;
	    RECT 348.0000 891.6000 354.3000 892.8000 ;
	    RECT 355.2000 891.9000 358.2000 892.8000 ;
	    RECT 335.4000 890.4000 339.3000 891.6000 ;
	    RECT 340.2000 890.7000 348.9000 891.6000 ;
	    RECT 353.4000 891.0000 354.3000 891.6000 ;
	    RECT 323.4000 889.5000 324.6000 889.8000 ;
	    RECT 225.0000 888.4500 226.2000 888.6000 ;
	    RECT 304.2000 888.4500 305.4000 888.6000 ;
	    RECT 49.8000 882.4500 51.0000 882.6000 ;
	    RECT 52.2000 882.4500 53.4000 882.6000 ;
	    RECT 49.8000 881.5500 53.4000 882.4500 ;
	    RECT 54.3000 882.3000 54.9000 883.5000 ;
	    RECT 56.1000 882.3000 60.0000 883.5000 ;
	    RECT 61.5000 882.3000 65.1000 883.5000 ;
	    RECT 66.3000 882.3000 70.2000 883.5000 ;
	    RECT 49.8000 881.4000 51.0000 881.5500 ;
	    RECT 52.2000 881.4000 53.4000 881.5500 ;
	    RECT 56.1000 881.4000 57.3000 882.3000 ;
	    RECT 61.5000 881.4000 62.7000 882.3000 ;
	    RECT 66.3000 881.4000 67.5000 882.3000 ;
	    RECT 71.4000 881.4000 72.6000 883.5000 ;
	    RECT 54.6000 880.2000 57.3000 881.4000 ;
	    RECT 59.4000 880.2000 62.7000 881.4000 ;
	    RECT 64.2000 880.2000 67.5000 881.4000 ;
	    RECT 69.0000 880.2000 72.6000 881.4000 ;
	    RECT 52.2000 873.3000 53.4000 879.3000 ;
	    RECT 54.6000 873.3000 55.8000 880.2000 ;
	    RECT 57.0000 873.3000 58.2000 879.3000 ;
	    RECT 59.4000 873.3000 60.6000 880.2000 ;
	    RECT 61.8000 873.3000 63.0000 879.3000 ;
	    RECT 64.2000 873.3000 65.4000 880.2000 ;
	    RECT 66.6000 873.3000 67.8000 879.3000 ;
	    RECT 69.0000 873.3000 70.2000 880.2000 ;
	    RECT 93.0000 879.3000 94.2000 883.5000 ;
	    RECT 170.4000 882.6000 171.3000 887.7000 ;
	    RECT 225.0000 887.5500 305.4000 888.4500 ;
	    RECT 309.0000 888.0000 310.2000 889.5000 ;
	    RECT 225.0000 887.4000 226.2000 887.5500 ;
	    RECT 304.2000 887.4000 305.4000 887.5500 ;
	    RECT 308.7000 886.8000 310.2000 888.0000 ;
	    RECT 311.1000 888.6000 324.6000 889.5000 ;
	    RECT 328.2000 889.5000 329.4000 889.8000 ;
	    RECT 340.2000 889.5000 341.1000 890.7000 ;
	    RECT 349.8000 889.8000 351.9000 890.7000 ;
	    RECT 353.4000 889.8000 355.8000 891.0000 ;
	    RECT 328.2000 888.6000 341.1000 889.5000 ;
	    RECT 342.6000 889.5000 351.9000 889.8000 ;
	    RECT 342.6000 888.9000 350.7000 889.5000 ;
	    RECT 342.6000 888.6000 343.8000 888.9000 ;
	    RECT 172.2000 885.4500 173.4000 885.6000 ;
	    RECT 177.0000 885.4500 178.2000 885.6000 ;
	    RECT 172.2000 884.5500 178.2000 885.4500 ;
	    RECT 172.2000 884.4000 173.4000 884.5500 ;
	    RECT 177.0000 884.4000 178.2000 884.5500 ;
	    RECT 172.2000 883.2000 173.4000 883.5000 ;
	    RECT 95.4000 882.4500 96.6000 882.6000 ;
	    RECT 102.6000 882.4500 103.8000 882.6000 ;
	    RECT 95.4000 881.5500 103.8000 882.4500 ;
	    RECT 95.4000 881.4000 96.6000 881.5500 ;
	    RECT 102.6000 881.4000 103.8000 881.5500 ;
	    RECT 112.2000 882.4500 113.4000 882.6000 ;
	    RECT 117.0000 882.4500 118.2000 882.6000 ;
	    RECT 112.2000 881.5500 118.2000 882.4500 ;
	    RECT 112.2000 881.4000 113.4000 881.5500 ;
	    RECT 117.0000 881.4000 118.2000 881.5500 ;
	    RECT 129.0000 882.4500 130.2000 882.6000 ;
	    RECT 133.8000 882.4500 135.0000 882.6000 ;
	    RECT 129.0000 881.5500 135.0000 882.4500 ;
	    RECT 129.0000 881.4000 130.2000 881.5500 ;
	    RECT 133.8000 881.4000 135.0000 881.5500 ;
	    RECT 143.4000 882.4500 144.6000 882.6000 ;
	    RECT 155.4000 882.4500 156.6000 882.6000 ;
	    RECT 143.4000 881.5500 156.6000 882.4500 ;
	    RECT 143.4000 881.4000 144.6000 881.5500 ;
	    RECT 155.4000 881.4000 156.6000 881.5500 ;
	    RECT 167.4000 881.4000 168.6000 882.6000 ;
	    RECT 169.5000 881.4000 171.3000 882.6000 ;
	    RECT 174.6000 882.4500 175.8000 882.6000 ;
	    RECT 227.4000 882.4500 228.6000 882.6000 ;
	    RECT 173.4000 880.8000 173.7000 882.3000 ;
	    RECT 174.6000 881.5500 228.6000 882.4500 ;
	    RECT 174.6000 881.4000 175.8000 881.5500 ;
	    RECT 227.4000 881.4000 228.6000 881.5500 ;
	    RECT 95.4000 880.2000 96.6000 880.5000 ;
	    RECT 71.4000 873.3000 72.6000 879.3000 ;
	    RECT 91.5000 878.4000 94.2000 879.3000 ;
	    RECT 91.5000 873.3000 92.7000 878.4000 ;
	    RECT 95.4000 873.3000 96.6000 879.3000 ;
	    RECT 109.8000 878.4000 111.0000 879.6000 ;
	    RECT 109.8000 877.2000 111.0000 877.5000 ;
	    RECT 109.8000 873.3000 111.0000 876.3000 ;
	    RECT 112.2000 873.3000 113.4000 880.5000 ;
	    RECT 121.8000 879.4500 123.0000 879.6000 ;
	    RECT 126.6000 879.4500 127.8000 879.6000 ;
	    RECT 121.8000 878.5500 127.8000 879.4500 ;
	    RECT 121.8000 878.4000 123.0000 878.5500 ;
	    RECT 126.6000 878.4000 127.8000 878.5500 ;
	    RECT 126.6000 877.2000 127.8000 877.5000 ;
	    RECT 126.6000 873.3000 127.8000 876.3000 ;
	    RECT 129.0000 873.3000 130.2000 880.5000 ;
	    RECT 141.0000 878.4000 142.2000 879.6000 ;
	    RECT 141.0000 877.2000 142.2000 877.5000 ;
	    RECT 141.0000 873.3000 142.2000 876.3000 ;
	    RECT 143.4000 873.3000 144.6000 880.5000 ;
	    RECT 167.7000 879.3000 168.6000 880.5000 ;
	    RECT 308.7000 880.2000 309.9000 886.8000 ;
	    RECT 311.1000 885.9000 312.0000 888.6000 ;
	    RECT 347.1000 887.7000 348.3000 888.0000 ;
	    RECT 312.9000 886.8000 351.3000 887.7000 ;
	    RECT 352.2000 887.4000 353.4000 888.6000 ;
	    RECT 312.9000 886.5000 314.1000 886.8000 ;
	    RECT 310.8000 885.0000 312.0000 885.9000 ;
	    RECT 321.0000 885.0000 346.5000 885.9000 ;
	    RECT 310.8000 882.0000 311.7000 885.0000 ;
	    RECT 321.0000 884.1000 322.2000 885.0000 ;
	    RECT 347.4000 884.4000 348.6000 885.6000 ;
	    RECT 349.5000 885.0000 356.1000 885.9000 ;
	    RECT 354.9000 884.7000 356.1000 885.0000 ;
	    RECT 312.6000 882.9000 318.3000 884.1000 ;
	    RECT 310.8000 881.1000 312.6000 882.0000 ;
	    RECT 170.1000 879.3000 175.5000 879.9000 ;
	    RECT 167.4000 873.3000 168.6000 879.3000 ;
	    RECT 169.8000 879.0000 175.8000 879.3000 ;
	    RECT 308.7000 879.0000 310.2000 880.2000 ;
	    RECT 169.8000 873.3000 171.0000 879.0000 ;
	    RECT 172.2000 873.3000 173.4000 878.1000 ;
	    RECT 174.6000 873.3000 175.8000 879.0000 ;
	    RECT 306.6000 873.3000 307.8000 876.3000 ;
	    RECT 309.0000 873.3000 310.2000 879.0000 ;
	    RECT 311.4000 873.3000 312.6000 881.1000 ;
	    RECT 317.1000 881.1000 318.3000 882.9000 ;
	    RECT 317.1000 880.2000 319.8000 881.1000 ;
	    RECT 318.6000 879.3000 319.8000 880.2000 ;
	    RECT 325.8000 879.6000 327.0000 883.8000 ;
	    RECT 330.6000 882.9000 335.4000 884.1000 ;
	    RECT 341.1000 882.9000 344.1000 884.1000 ;
	    RECT 357.0000 883.5000 358.2000 891.9000 ;
	    RECT 371.4000 883.5000 372.6000 899.7000 ;
	    RECT 402.6000 887.7000 403.8000 899.7000 ;
	    RECT 406.5000 887.7000 409.5000 899.7000 ;
	    RECT 412.2000 887.7000 413.4000 899.7000 ;
	    RECT 546.6000 893.7000 547.8000 899.7000 ;
	    RECT 549.0000 892.5000 550.2000 899.7000 ;
	    RECT 551.4000 893.7000 552.6000 899.7000 ;
	    RECT 553.8000 892.8000 555.0000 899.7000 ;
	    RECT 556.2000 893.7000 557.4000 899.7000 ;
	    RECT 551.1000 891.9000 555.0000 892.8000 ;
	    RECT 450.6000 891.4500 451.8000 891.6000 ;
	    RECT 549.0000 891.4500 550.2000 891.6000 ;
	    RECT 450.6000 890.5500 550.2000 891.4500 ;
	    RECT 450.6000 890.4000 451.8000 890.5500 ;
	    RECT 549.0000 890.4000 550.2000 890.5500 ;
	    RECT 551.1000 889.5000 552.0000 891.9000 ;
	    RECT 558.6000 891.6000 559.8000 899.7000 ;
	    RECT 561.0000 893.7000 562.2000 899.7000 ;
	    RECT 563.4000 895.5000 564.6000 899.7000 ;
	    RECT 565.8000 895.5000 567.0000 899.7000 ;
	    RECT 568.2000 895.5000 569.4000 899.7000 ;
	    RECT 560.7000 891.6000 567.0000 892.8000 ;
	    RECT 555.9000 890.4000 559.8000 891.6000 ;
	    RECT 570.6000 890.4000 571.8000 899.7000 ;
	    RECT 573.0000 893.7000 574.2000 899.7000 ;
	    RECT 575.4000 892.5000 576.6000 899.7000 ;
	    RECT 577.8000 893.7000 579.0000 899.7000 ;
	    RECT 580.2000 892.5000 581.4000 899.7000 ;
	    RECT 582.6000 895.5000 583.8000 899.7000 ;
	    RECT 585.0000 895.5000 586.2000 899.7000 ;
	    RECT 587.4000 893.7000 588.6000 899.7000 ;
	    RECT 589.8000 892.8000 591.0000 899.7000 ;
	    RECT 592.2000 893.7000 593.4000 900.6000 ;
	    RECT 594.6000 894.6000 595.8000 899.7000 ;
	    RECT 594.6000 893.7000 596.1000 894.6000 ;
	    RECT 597.0000 893.7000 598.2000 899.7000 ;
	    RECT 611.4000 893.7000 612.6000 899.7000 ;
	    RECT 595.2000 892.8000 596.1000 893.7000 ;
	    RECT 588.0000 891.6000 594.3000 892.8000 ;
	    RECT 595.2000 891.9000 598.2000 892.8000 ;
	    RECT 575.4000 890.4000 579.3000 891.6000 ;
	    RECT 580.2000 890.7000 588.9000 891.6000 ;
	    RECT 593.4000 891.0000 594.3000 891.6000 ;
	    RECT 563.4000 889.5000 564.6000 889.8000 ;
	    RECT 549.0000 888.0000 550.2000 889.5000 ;
	    RECT 385.8000 885.4500 387.0000 885.6000 ;
	    RECT 405.0000 885.4500 406.2000 885.6000 ;
	    RECT 385.8000 884.5500 406.2000 885.4500 ;
	    RECT 385.8000 884.4000 387.0000 884.5500 ;
	    RECT 405.0000 884.4000 406.2000 884.5500 ;
	    RECT 407.4000 883.5000 408.3000 887.7000 ;
	    RECT 548.7000 886.8000 550.2000 888.0000 ;
	    RECT 551.1000 888.6000 564.6000 889.5000 ;
	    RECT 568.2000 889.5000 569.4000 889.8000 ;
	    RECT 580.2000 889.5000 581.1000 890.7000 ;
	    RECT 589.8000 889.8000 591.9000 890.7000 ;
	    RECT 593.4000 889.8000 595.8000 891.0000 ;
	    RECT 568.2000 888.6000 581.1000 889.5000 ;
	    RECT 582.6000 889.5000 591.9000 889.8000 ;
	    RECT 582.6000 888.9000 590.7000 889.5000 ;
	    RECT 582.6000 888.6000 583.8000 888.9000 ;
	    RECT 409.8000 884.4000 411.0000 885.6000 ;
	    RECT 412.2000 883.5000 413.4000 883.8000 ;
	    RECT 330.0000 881.7000 331.2000 882.0000 ;
	    RECT 330.0000 880.8000 336.6000 881.7000 ;
	    RECT 337.8000 881.4000 339.0000 882.6000 ;
	    RECT 335.4000 880.5000 336.6000 880.8000 ;
	    RECT 337.8000 880.2000 339.0000 880.5000 ;
	    RECT 316.2000 873.3000 317.4000 879.3000 ;
	    RECT 318.6000 878.1000 322.2000 879.3000 ;
	    RECT 325.8000 878.4000 327.3000 879.6000 ;
	    RECT 331.8000 878.4000 332.1000 879.6000 ;
	    RECT 333.0000 878.4000 334.2000 879.6000 ;
	    RECT 335.4000 879.3000 336.6000 879.6000 ;
	    RECT 341.1000 879.3000 342.3000 882.9000 ;
	    RECT 345.0000 882.3000 358.2000 883.5000 ;
	    RECT 405.0000 883.2000 406.2000 883.5000 ;
	    RECT 409.8000 883.2000 411.0000 883.5000 ;
	    RECT 350.1000 880.2000 354.6000 881.4000 ;
	    RECT 350.1000 879.3000 351.3000 880.2000 ;
	    RECT 335.4000 878.4000 342.3000 879.3000 ;
	    RECT 321.0000 873.3000 322.2000 878.1000 ;
	    RECT 347.4000 878.1000 351.3000 879.3000 ;
	    RECT 323.4000 873.3000 324.6000 877.5000 ;
	    RECT 325.8000 873.3000 327.0000 877.5000 ;
	    RECT 328.2000 873.3000 329.4000 877.5000 ;
	    RECT 330.6000 873.3000 331.8000 877.5000 ;
	    RECT 333.0000 873.3000 334.2000 876.3000 ;
	    RECT 335.4000 873.3000 336.6000 877.5000 ;
	    RECT 337.8000 873.3000 339.0000 876.3000 ;
	    RECT 340.2000 873.3000 341.4000 877.5000 ;
	    RECT 342.6000 873.3000 343.8000 877.5000 ;
	    RECT 345.0000 873.3000 346.2000 877.5000 ;
	    RECT 347.4000 873.3000 348.6000 878.1000 ;
	    RECT 352.2000 873.3000 353.4000 879.3000 ;
	    RECT 357.0000 873.3000 358.2000 882.3000 ;
	    RECT 371.4000 882.4500 372.6000 882.6000 ;
	    RECT 402.6000 882.4500 403.8000 882.6000 ;
	    RECT 371.4000 881.5500 403.8000 882.4500 ;
	    RECT 371.4000 881.4000 372.6000 881.5500 ;
	    RECT 402.6000 881.4000 403.8000 881.5500 ;
	    RECT 404.7000 880.8000 405.0000 882.3000 ;
	    RECT 407.4000 881.4000 408.6000 882.6000 ;
	    RECT 409.5000 881.4000 411.0000 882.3000 ;
	    RECT 412.2000 881.4000 413.4000 882.6000 ;
	    RECT 364.2000 879.4500 365.4000 879.6000 ;
	    RECT 369.0000 879.4500 370.2000 879.6000 ;
	    RECT 364.2000 878.5500 370.2000 879.4500 ;
	    RECT 364.2000 878.4000 365.4000 878.5500 ;
	    RECT 369.0000 878.4000 370.2000 878.5500 ;
	    RECT 369.0000 877.2000 370.2000 877.5000 ;
	    RECT 369.0000 873.3000 370.2000 876.3000 ;
	    RECT 371.4000 873.3000 372.6000 880.5000 ;
	    RECT 402.9000 879.3000 408.3000 879.9000 ;
	    RECT 410.1000 879.3000 411.0000 881.4000 ;
	    RECT 548.7000 880.2000 549.9000 886.8000 ;
	    RECT 551.1000 885.9000 552.0000 888.6000 ;
	    RECT 587.1000 887.7000 588.3000 888.0000 ;
	    RECT 552.9000 886.8000 591.3000 887.7000 ;
	    RECT 592.2000 887.4000 593.4000 888.6000 ;
	    RECT 552.9000 886.5000 554.1000 886.8000 ;
	    RECT 550.8000 885.0000 552.0000 885.9000 ;
	    RECT 561.0000 885.0000 586.5000 885.9000 ;
	    RECT 550.8000 882.0000 551.7000 885.0000 ;
	    RECT 561.0000 884.1000 562.2000 885.0000 ;
	    RECT 587.4000 884.4000 588.6000 885.6000 ;
	    RECT 589.5000 885.0000 596.1000 885.9000 ;
	    RECT 594.9000 884.7000 596.1000 885.0000 ;
	    RECT 552.6000 882.9000 558.3000 884.1000 ;
	    RECT 550.8000 881.1000 552.6000 882.0000 ;
	    RECT 402.6000 879.0000 408.6000 879.3000 ;
	    RECT 402.6000 873.3000 403.8000 879.0000 ;
	    RECT 405.0000 873.3000 406.2000 878.1000 ;
	    RECT 407.4000 874.2000 408.6000 879.0000 ;
	    RECT 409.8000 875.1000 411.0000 879.3000 ;
	    RECT 412.2000 874.2000 413.4000 879.3000 ;
	    RECT 548.7000 879.0000 550.2000 880.2000 ;
	    RECT 407.4000 873.3000 413.4000 874.2000 ;
	    RECT 546.6000 873.3000 547.8000 876.3000 ;
	    RECT 549.0000 873.3000 550.2000 879.0000 ;
	    RECT 551.4000 873.3000 552.6000 881.1000 ;
	    RECT 557.1000 881.1000 558.3000 882.9000 ;
	    RECT 557.1000 880.2000 559.8000 881.1000 ;
	    RECT 558.6000 879.3000 559.8000 880.2000 ;
	    RECT 565.8000 879.6000 567.0000 883.8000 ;
	    RECT 570.6000 882.9000 575.4000 884.1000 ;
	    RECT 581.1000 882.9000 584.1000 884.1000 ;
	    RECT 597.0000 883.5000 598.2000 891.9000 ;
	    RECT 613.8000 883.5000 615.0000 899.7000 ;
	    RECT 633.0000 893.7000 634.2000 899.7000 ;
	    RECT 633.0000 889.5000 634.2000 889.8000 ;
	    RECT 623.4000 888.4500 624.6000 888.6000 ;
	    RECT 633.0000 888.4500 634.2000 888.6000 ;
	    RECT 623.4000 887.5500 634.2000 888.4500 ;
	    RECT 623.4000 887.4000 624.6000 887.5500 ;
	    RECT 633.0000 887.4000 634.2000 887.5500 ;
	    RECT 635.4000 886.5000 636.6000 899.7000 ;
	    RECT 637.8000 893.7000 639.0000 899.7000 ;
	    RECT 633.0000 885.4500 634.2000 885.6000 ;
	    RECT 635.4000 885.4500 636.6000 885.6000 ;
	    RECT 633.0000 884.5500 636.6000 885.4500 ;
	    RECT 633.0000 884.4000 634.2000 884.5500 ;
	    RECT 635.4000 884.4000 636.6000 884.5500 ;
	    RECT 649.8000 883.5000 651.0000 899.7000 ;
	    RECT 652.2000 893.7000 653.4000 899.7000 ;
	    RECT 678.6000 893.7000 679.8000 899.7000 ;
	    RECT 678.6000 889.5000 679.8000 889.8000 ;
	    RECT 678.6000 887.4000 679.8000 888.6000 ;
	    RECT 681.0000 886.5000 682.2000 899.7000 ;
	    RECT 683.4000 893.7000 684.6000 899.7000 ;
	    RECT 731.4000 890.7000 732.6000 899.7000 ;
	    RECT 733.8000 890.7000 735.0000 899.7000 ;
	    RECT 736.2000 898.8000 742.2000 899.7000 ;
	    RECT 736.2000 890.7000 737.4000 898.8000 ;
	    RECT 738.6000 890.7000 739.8000 897.9000 ;
	    RECT 741.0000 891.0000 742.2000 898.8000 ;
	    RECT 743.7000 898.8000 749.1000 899.7000 ;
	    RECT 743.7000 898.5000 744.6000 898.8000 ;
	    RECT 731.7000 889.8000 732.6000 890.7000 ;
	    RECT 736.2000 889.8000 737.1000 890.7000 ;
	    RECT 731.7000 888.9000 737.1000 889.8000 ;
	    RECT 738.9000 890.1000 739.8000 890.7000 ;
	    RECT 743.4000 890.1000 744.6000 898.5000 ;
	    RECT 748.2000 898.5000 749.1000 898.8000 ;
	    RECT 738.9000 889.5000 744.6000 890.1000 ;
	    RECT 745.8000 889.5000 747.0000 897.9000 ;
	    RECT 748.2000 889.5000 749.4000 898.5000 ;
	    RECT 767.4000 893.7000 768.6000 899.7000 ;
	    RECT 738.9000 889.2000 744.3000 889.5000 ;
	    RECT 745.8000 888.4500 747.0000 888.6000 ;
	    RECT 767.4000 888.4500 768.6000 888.6000 ;
	    RECT 741.9000 887.4000 744.9000 888.3000 ;
	    RECT 745.8000 887.5500 768.6000 888.4500 ;
	    RECT 745.8000 887.4000 747.0000 887.5500 ;
	    RECT 767.4000 887.4000 768.6000 887.5500 ;
	    RECT 681.0000 885.4500 682.2000 885.6000 ;
	    RECT 685.8000 885.4500 687.0000 885.6000 ;
	    RECT 717.0000 885.4500 718.2000 885.6000 ;
	    RECT 681.0000 884.5500 718.2000 885.4500 ;
	    RECT 681.0000 884.4000 682.2000 884.5500 ;
	    RECT 685.8000 884.4000 687.0000 884.5500 ;
	    RECT 717.0000 884.4000 718.2000 884.5500 ;
	    RECT 738.6000 884.4000 739.8000 885.6000 ;
	    RECT 740.7000 884.4000 741.0000 885.6000 ;
	    RECT 570.0000 881.7000 571.2000 882.0000 ;
	    RECT 570.0000 880.8000 576.6000 881.7000 ;
	    RECT 577.8000 881.4000 579.0000 882.6000 ;
	    RECT 575.4000 880.5000 576.6000 880.8000 ;
	    RECT 577.8000 880.2000 579.0000 880.5000 ;
	    RECT 556.2000 873.3000 557.4000 879.3000 ;
	    RECT 558.6000 878.1000 562.2000 879.3000 ;
	    RECT 565.8000 878.4000 567.3000 879.6000 ;
	    RECT 571.8000 878.4000 572.1000 879.6000 ;
	    RECT 573.0000 878.4000 574.2000 879.6000 ;
	    RECT 575.4000 879.3000 576.6000 879.6000 ;
	    RECT 581.1000 879.3000 582.3000 882.9000 ;
	    RECT 585.0000 882.3000 598.2000 883.5000 ;
	    RECT 590.1000 880.2000 594.6000 881.4000 ;
	    RECT 590.1000 879.3000 591.3000 880.2000 ;
	    RECT 575.4000 878.4000 582.3000 879.3000 ;
	    RECT 561.0000 873.3000 562.2000 878.1000 ;
	    RECT 587.4000 878.1000 591.3000 879.3000 ;
	    RECT 563.4000 873.3000 564.6000 877.5000 ;
	    RECT 565.8000 873.3000 567.0000 877.5000 ;
	    RECT 568.2000 873.3000 569.4000 877.5000 ;
	    RECT 570.6000 873.3000 571.8000 877.5000 ;
	    RECT 573.0000 873.3000 574.2000 876.3000 ;
	    RECT 575.4000 873.3000 576.6000 877.5000 ;
	    RECT 577.8000 873.3000 579.0000 876.3000 ;
	    RECT 580.2000 873.3000 581.4000 877.5000 ;
	    RECT 582.6000 873.3000 583.8000 877.5000 ;
	    RECT 585.0000 873.3000 586.2000 877.5000 ;
	    RECT 587.4000 873.3000 588.6000 878.1000 ;
	    RECT 592.2000 873.3000 593.4000 879.3000 ;
	    RECT 597.0000 873.3000 598.2000 882.3000 ;
	    RECT 599.4000 882.4500 600.6000 882.6000 ;
	    RECT 613.8000 882.4500 615.0000 882.6000 ;
	    RECT 599.4000 881.5500 615.0000 882.4500 ;
	    RECT 599.4000 881.4000 600.6000 881.5500 ;
	    RECT 613.8000 881.4000 615.0000 881.5500 ;
	    RECT 611.4000 878.4000 612.6000 879.6000 ;
	    RECT 611.4000 877.2000 612.6000 877.5000 ;
	    RECT 611.4000 873.3000 612.6000 876.3000 ;
	    RECT 613.8000 873.3000 615.0000 880.5000 ;
	    RECT 635.4000 879.3000 636.6000 883.5000 ;
	    RECT 637.8000 881.4000 639.0000 882.6000 ;
	    RECT 642.6000 882.4500 643.8000 882.6000 ;
	    RECT 649.8000 882.4500 651.0000 882.6000 ;
	    RECT 642.6000 881.5500 651.0000 882.4500 ;
	    RECT 642.6000 881.4000 643.8000 881.5500 ;
	    RECT 649.8000 881.4000 651.0000 881.5500 ;
	    RECT 637.8000 880.2000 639.0000 880.5000 ;
	    RECT 633.9000 878.4000 636.6000 879.3000 ;
	    RECT 633.9000 873.3000 635.1000 878.4000 ;
	    RECT 637.8000 873.3000 639.0000 879.3000 ;
	    RECT 649.8000 873.3000 651.0000 880.5000 ;
	    RECT 652.2000 879.4500 653.4000 879.6000 ;
	    RECT 654.6000 879.4500 655.8000 879.6000 ;
	    RECT 652.2000 878.5500 655.8000 879.4500 ;
	    RECT 681.0000 879.3000 682.2000 883.5000 ;
	    RECT 683.4000 881.4000 684.6000 882.6000 ;
	    RECT 736.2000 881.4000 737.4000 882.6000 ;
	    RECT 738.3000 881.4000 738.6000 882.6000 ;
	    RECT 683.4000 880.2000 684.6000 880.5000 ;
	    RECT 652.2000 878.4000 653.4000 878.5500 ;
	    RECT 654.6000 878.4000 655.8000 878.5500 ;
	    RECT 679.5000 878.4000 682.2000 879.3000 ;
	    RECT 652.2000 877.2000 653.4000 877.5000 ;
	    RECT 652.2000 873.3000 653.4000 876.3000 ;
	    RECT 679.5000 873.3000 680.7000 878.4000 ;
	    RECT 683.4000 873.3000 684.6000 879.3000 ;
	    RECT 733.8000 878.4000 735.0000 879.6000 ;
	    RECT 735.9000 878.4000 736.5000 879.6000 ;
	    RECT 741.9000 877.5000 742.8000 887.4000 ;
	    RECT 769.8000 886.5000 771.0000 899.7000 ;
	    RECT 772.2000 893.7000 773.4000 899.7000 ;
	    RECT 772.2000 889.5000 773.4000 889.8000 ;
	    RECT 815.4000 888.6000 816.6000 899.7000 ;
	    RECT 817.8000 889.8000 819.3000 899.7000 ;
	    RECT 817.8000 888.6000 819.0000 888.9000 ;
	    RECT 772.2000 888.4500 773.4000 888.6000 ;
	    RECT 786.6000 888.4500 787.8000 888.6000 ;
	    RECT 772.2000 887.5500 787.8000 888.4500 ;
	    RECT 815.4000 887.7000 819.0000 888.6000 ;
	    RECT 822.0000 887.7000 824.4000 899.7000 ;
	    RECT 827.1000 889.8000 828.6000 899.7000 ;
	    RECT 827.1000 888.6000 828.3000 888.9000 ;
	    RECT 829.8000 888.6000 831.0000 899.7000 ;
	    RECT 827.1000 887.7000 831.0000 888.6000 ;
	    RECT 772.2000 887.4000 773.4000 887.5500 ;
	    RECT 786.6000 887.4000 787.8000 887.5500 ;
	    RECT 822.6000 886.5000 823.5000 887.7000 ;
	    RECT 825.3000 885.6000 826.5000 885.9000 ;
	    RECT 745.8000 885.4500 747.0000 885.6000 ;
	    RECT 769.8000 885.4500 771.0000 885.6000 ;
	    RECT 745.8000 884.5500 771.0000 885.4500 ;
	    RECT 745.8000 884.4000 747.0000 884.5500 ;
	    RECT 769.8000 884.4000 771.0000 884.5500 ;
	    RECT 813.0000 885.4500 814.2000 885.6000 ;
	    RECT 822.6000 885.4500 823.8000 885.6000 ;
	    RECT 813.0000 884.5500 823.8000 885.4500 ;
	    RECT 825.3000 884.7000 827.7000 885.6000 ;
	    RECT 813.0000 884.4000 814.2000 884.5500 ;
	    RECT 822.6000 884.4000 823.8000 884.5500 ;
	    RECT 826.5000 884.4000 827.7000 884.7000 ;
	    RECT 844.2000 883.5000 845.4000 899.7000 ;
	    RECT 846.6000 893.7000 847.8000 899.7000 ;
	    RECT 861.0000 893.7000 862.2000 899.7000 ;
	    RECT 863.4000 883.5000 864.6000 899.7000 ;
	    RECT 888.3000 893.7000 889.5000 899.7000 ;
	    RECT 888.6000 890.4000 889.8000 891.6000 ;
	    RECT 888.6000 889.5000 889.5000 890.4000 ;
	    RECT 890.7000 888.6000 891.9000 899.7000 ;
	    RECT 887.4000 887.4000 888.6000 888.6000 ;
	    RECT 890.4000 887.7000 891.9000 888.6000 ;
	    RECT 894.6000 887.7000 895.8000 899.7000 ;
	    RECT 921.0000 893.7000 922.2000 899.7000 ;
	    RECT 921.0000 889.5000 922.2000 889.8000 ;
	    RECT 767.4000 881.4000 768.6000 882.6000 ;
	    RECT 767.4000 880.2000 768.6000 880.5000 ;
	    RECT 769.8000 879.3000 771.0000 883.5000 ;
	    RECT 822.6000 882.6000 823.5000 883.5000 ;
	    RECT 815.4000 881.4000 816.6000 882.6000 ;
	    RECT 817.5000 881.4000 817.8000 882.6000 ;
	    RECT 819.6000 881.4000 820.8000 882.6000 ;
	    RECT 819.9000 880.8000 820.8000 881.4000 ;
	    RECT 822.0000 881.7000 823.5000 882.6000 ;
	    RECT 824.4000 882.9000 825.6000 883.2000 ;
	    RECT 824.4000 882.6000 828.6000 882.9000 ;
	    RECT 890.4000 882.6000 891.3000 887.7000 ;
	    RECT 921.0000 887.4000 922.2000 888.6000 ;
	    RECT 923.4000 886.5000 924.6000 899.7000 ;
	    RECT 925.8000 893.7000 927.0000 899.7000 ;
	    RECT 950.7000 893.7000 951.9000 899.7000 ;
	    RECT 951.0000 890.4000 952.2000 891.6000 ;
	    RECT 951.0000 889.5000 951.9000 890.4000 ;
	    RECT 953.1000 888.6000 954.3000 899.7000 ;
	    RECT 940.2000 888.4500 941.4000 888.6000 ;
	    RECT 949.8000 888.4500 951.0000 888.6000 ;
	    RECT 940.2000 887.5500 951.0000 888.4500 ;
	    RECT 940.2000 887.4000 941.4000 887.5500 ;
	    RECT 949.8000 887.4000 951.0000 887.5500 ;
	    RECT 952.8000 887.7000 954.3000 888.6000 ;
	    RECT 957.0000 887.7000 958.2000 899.7000 ;
	    RECT 971.4000 893.7000 972.6000 899.7000 ;
	    RECT 892.2000 884.4000 893.4000 885.6000 ;
	    RECT 894.6000 885.4500 895.8000 885.6000 ;
	    RECT 923.4000 885.4500 924.6000 885.6000 ;
	    RECT 894.6000 884.5500 924.6000 885.4500 ;
	    RECT 894.6000 884.4000 895.8000 884.5500 ;
	    RECT 923.4000 884.4000 924.6000 884.5500 ;
	    RECT 928.2000 885.4500 929.4000 885.6000 ;
	    RECT 949.8000 885.4500 951.0000 885.6000 ;
	    RECT 928.2000 884.5500 951.0000 885.4500 ;
	    RECT 928.2000 884.4000 929.4000 884.5500 ;
	    RECT 949.8000 884.4000 951.0000 884.5500 ;
	    RECT 892.2000 883.2000 893.4000 883.5000 ;
	    RECT 824.4000 882.0000 828.9000 882.6000 ;
	    RECT 827.7000 881.7000 828.9000 882.0000 ;
	    RECT 817.8000 880.2000 819.0000 880.5000 ;
	    RECT 815.4000 879.3000 819.0000 880.2000 ;
	    RECT 819.9000 879.6000 821.1000 880.8000 ;
	    RECT 736.8000 876.6000 742.8000 877.5000 ;
	    RECT 736.8000 876.3000 737.7000 876.6000 ;
	    RECT 733.8000 873.3000 735.0000 876.3000 ;
	    RECT 736.2000 875.4000 737.7000 876.3000 ;
	    RECT 741.0000 876.3000 742.8000 876.6000 ;
	    RECT 736.2000 873.3000 737.4000 875.4000 ;
	    RECT 738.6000 873.3000 739.8000 875.7000 ;
	    RECT 741.0000 873.3000 742.2000 876.3000 ;
	    RECT 767.4000 873.3000 768.6000 879.3000 ;
	    RECT 769.8000 878.4000 772.5000 879.3000 ;
	    RECT 771.3000 873.3000 772.5000 878.4000 ;
	    RECT 815.4000 873.3000 816.6000 879.3000 ;
	    RECT 822.0000 878.7000 822.9000 881.7000 ;
	    RECT 828.6000 881.4000 828.9000 881.7000 ;
	    RECT 829.8000 881.4000 831.0000 882.6000 ;
	    RECT 837.0000 882.4500 838.2000 882.6000 ;
	    RECT 844.2000 882.4500 845.4000 882.6000 ;
	    RECT 837.0000 881.5500 845.4000 882.4500 ;
	    RECT 837.0000 881.4000 838.2000 881.5500 ;
	    RECT 844.2000 881.4000 845.4000 881.5500 ;
	    RECT 863.4000 882.4500 864.6000 882.6000 ;
	    RECT 885.0000 882.4500 886.2000 882.6000 ;
	    RECT 863.4000 881.5500 886.2000 882.4500 ;
	    RECT 863.4000 881.4000 864.6000 881.5500 ;
	    RECT 885.0000 881.4000 886.2000 881.5500 ;
	    RECT 887.4000 881.4000 888.6000 882.6000 ;
	    RECT 889.5000 881.4000 891.3000 882.6000 ;
	    RECT 894.6000 882.4500 895.8000 882.6000 ;
	    RECT 899.4000 882.4500 900.6000 882.6000 ;
	    RECT 893.4000 880.8000 893.7000 882.3000 ;
	    RECT 894.6000 881.5500 900.6000 882.4500 ;
	    RECT 894.6000 881.4000 895.8000 881.5500 ;
	    RECT 899.4000 881.4000 900.6000 881.5500 ;
	    RECT 823.8000 879.6000 826.2000 880.8000 ;
	    RECT 827.1000 880.2000 828.3000 880.5000 ;
	    RECT 827.1000 879.3000 831.0000 880.2000 ;
	    RECT 817.8000 873.3000 819.3000 878.4000 ;
	    RECT 822.0000 873.3000 824.4000 878.7000 ;
	    RECT 827.1000 873.3000 828.6000 878.4000 ;
	    RECT 829.8000 873.3000 831.0000 879.3000 ;
	    RECT 844.2000 873.3000 845.4000 880.5000 ;
	    RECT 846.6000 878.4000 847.8000 879.6000 ;
	    RECT 861.0000 878.4000 862.2000 879.6000 ;
	    RECT 846.6000 877.2000 847.8000 877.5000 ;
	    RECT 861.0000 877.2000 862.2000 877.5000 ;
	    RECT 846.6000 873.3000 847.8000 876.3000 ;
	    RECT 861.0000 873.3000 862.2000 876.3000 ;
	    RECT 863.4000 873.3000 864.6000 880.5000 ;
	    RECT 887.7000 879.3000 888.6000 880.5000 ;
	    RECT 890.1000 879.3000 895.5000 879.9000 ;
	    RECT 923.4000 879.3000 924.6000 883.5000 ;
	    RECT 952.8000 882.6000 953.7000 887.7000 ;
	    RECT 954.6000 885.4500 955.8000 885.6000 ;
	    RECT 954.6000 884.5500 960.4500 885.4500 ;
	    RECT 954.6000 884.4000 955.8000 884.5500 ;
	    RECT 954.6000 883.2000 955.8000 883.5000 ;
	    RECT 925.8000 882.4500 927.0000 882.6000 ;
	    RECT 928.2000 882.4500 929.4000 882.6000 ;
	    RECT 925.8000 881.5500 929.4000 882.4500 ;
	    RECT 925.8000 881.4000 927.0000 881.5500 ;
	    RECT 928.2000 881.4000 929.4000 881.5500 ;
	    RECT 935.4000 882.4500 936.6000 882.6000 ;
	    RECT 945.0000 882.4500 946.2000 882.6000 ;
	    RECT 935.4000 881.5500 946.2000 882.4500 ;
	    RECT 935.4000 881.4000 936.6000 881.5500 ;
	    RECT 945.0000 881.4000 946.2000 881.5500 ;
	    RECT 947.4000 882.4500 948.6000 882.6000 ;
	    RECT 949.8000 882.4500 951.0000 882.6000 ;
	    RECT 947.4000 881.5500 951.0000 882.4500 ;
	    RECT 947.4000 881.4000 948.6000 881.5500 ;
	    RECT 949.8000 881.4000 951.0000 881.5500 ;
	    RECT 951.9000 881.4000 953.7000 882.6000 ;
	    RECT 955.8000 880.8000 956.1000 882.3000 ;
	    RECT 957.0000 881.4000 958.2000 882.6000 ;
	    RECT 959.5500 882.4500 960.4500 884.5500 ;
	    RECT 973.8000 883.5000 975.0000 899.7000 ;
	    RECT 978.6000 894.4500 979.8000 894.6000 ;
	    RECT 988.2000 894.4500 989.4000 894.6000 ;
	    RECT 978.6000 893.5500 989.4000 894.4500 ;
	    RECT 993.0000 893.7000 994.2000 899.7000 ;
	    RECT 978.6000 893.4000 979.8000 893.5500 ;
	    RECT 988.2000 893.4000 989.4000 893.5500 ;
	    RECT 995.4000 886.5000 996.6000 899.7000 ;
	    RECT 997.8000 893.7000 999.0000 899.7000 ;
	    RECT 997.8000 889.5000 999.0000 889.8000 ;
	    RECT 997.8000 887.4000 999.0000 888.6000 ;
	    RECT 1026.6000 887.7000 1027.8000 899.7000 ;
	    RECT 1030.5000 887.7000 1033.5000 899.7000 ;
	    RECT 1036.2001 887.7000 1037.4000 899.7000 ;
	    RECT 976.2000 885.4500 977.4000 885.6000 ;
	    RECT 995.4000 885.4500 996.6000 885.6000 ;
	    RECT 976.2000 884.5500 996.6000 885.4500 ;
	    RECT 976.2000 884.4000 977.4000 884.5500 ;
	    RECT 995.4000 884.4000 996.6000 884.5500 ;
	    RECT 1029.0000 884.4000 1030.2001 885.6000 ;
	    RECT 1026.6000 883.5000 1027.8000 883.8000 ;
	    RECT 1031.7001 883.5000 1032.6000 887.7000 ;
	    RECT 1033.8000 884.4000 1035.0000 885.6000 ;
	    RECT 1050.6000 883.5000 1051.8000 899.7000 ;
	    RECT 1053.0000 893.7000 1054.2001 899.7000 ;
	    RECT 1185.0000 893.7000 1186.2001 899.7000 ;
	    RECT 1187.4000 894.6000 1188.6000 899.7000 ;
	    RECT 1187.1000 893.7000 1188.6000 894.6000 ;
	    RECT 1189.8000 893.7000 1191.0000 900.6000 ;
	    RECT 1187.1000 892.8000 1188.0000 893.7000 ;
	    RECT 1192.2001 892.8000 1193.4000 899.7000 ;
	    RECT 1194.6000 893.7000 1195.8000 899.7000 ;
	    RECT 1197.0000 895.5000 1198.2001 899.7000 ;
	    RECT 1199.4000 895.5000 1200.6000 899.7000 ;
	    RECT 1185.0000 891.9000 1188.0000 892.8000 ;
	    RECT 1185.0000 883.5000 1186.2001 891.9000 ;
	    RECT 1188.9000 891.6000 1195.2001 892.8000 ;
	    RECT 1201.8000 892.5000 1203.0000 899.7000 ;
	    RECT 1204.2001 893.7000 1205.4000 899.7000 ;
	    RECT 1206.6000 892.5000 1207.8000 899.7000 ;
	    RECT 1209.0000 893.7000 1210.2001 899.7000 ;
	    RECT 1188.9000 891.0000 1189.8000 891.6000 ;
	    RECT 1187.4000 889.8000 1189.8000 891.0000 ;
	    RECT 1194.3000 890.7000 1203.0000 891.6000 ;
	    RECT 1191.3000 889.8000 1193.4000 890.7000 ;
	    RECT 1191.3000 889.5000 1200.6000 889.8000 ;
	    RECT 1192.5000 888.9000 1200.6000 889.5000 ;
	    RECT 1199.4000 888.6000 1200.6000 888.9000 ;
	    RECT 1202.1000 889.5000 1203.0000 890.7000 ;
	    RECT 1203.9000 890.4000 1207.8000 891.6000 ;
	    RECT 1211.4000 890.4000 1212.6000 899.7000 ;
	    RECT 1213.8000 895.5000 1215.0000 899.7000 ;
	    RECT 1216.2001 895.5000 1217.4000 899.7000 ;
	    RECT 1218.6000 895.5000 1219.8000 899.7000 ;
	    RECT 1221.0000 893.7000 1222.2001 899.7000 ;
	    RECT 1216.2001 891.6000 1222.5000 892.8000 ;
	    RECT 1223.4000 891.6000 1224.6000 899.7000 ;
	    RECT 1225.8000 893.7000 1227.0000 899.7000 ;
	    RECT 1228.2001 892.8000 1229.4000 899.7000 ;
	    RECT 1230.6000 893.7000 1231.8000 899.7000 ;
	    RECT 1228.2001 891.9000 1232.1000 892.8000 ;
	    RECT 1233.0000 892.5000 1234.2001 899.7000 ;
	    RECT 1235.4000 893.7000 1236.6000 899.7000 ;
	    RECT 1262.7001 893.7000 1263.9000 899.7000 ;
	    RECT 1223.4000 890.4000 1227.3000 891.6000 ;
	    RECT 1213.8000 889.5000 1215.0000 889.8000 ;
	    RECT 1202.1000 888.6000 1215.0000 889.5000 ;
	    RECT 1218.6000 889.5000 1219.8000 889.8000 ;
	    RECT 1231.2001 889.5000 1232.1000 891.9000 ;
	    RECT 1233.0000 891.4500 1234.2001 891.6000 ;
	    RECT 1242.6000 891.4500 1243.8000 891.6000 ;
	    RECT 1233.0000 890.5500 1243.8000 891.4500 ;
	    RECT 1233.0000 890.4000 1234.2001 890.5500 ;
	    RECT 1242.6000 890.4000 1243.8000 890.5500 ;
	    RECT 1263.0000 890.4000 1264.2001 891.6000 ;
	    RECT 1263.0000 889.5000 1263.9000 890.4000 ;
	    RECT 1218.6000 888.6000 1232.1000 889.5000 ;
	    RECT 1189.8000 887.4000 1191.0000 888.6000 ;
	    RECT 1194.9000 887.7000 1196.1000 888.0000 ;
	    RECT 1191.9000 886.8000 1230.3000 887.7000 ;
	    RECT 1229.1000 886.5000 1230.3000 886.8000 ;
	    RECT 1231.2001 885.9000 1232.1000 888.6000 ;
	    RECT 1233.0000 888.0000 1234.2001 889.5000 ;
	    RECT 1265.1000 888.6000 1266.3000 899.7000 ;
	    RECT 1235.4000 888.4500 1236.6000 888.6000 ;
	    RECT 1261.8000 888.4500 1263.0000 888.6000 ;
	    RECT 1233.0000 886.8000 1234.5000 888.0000 ;
	    RECT 1235.4000 887.5500 1263.0000 888.4500 ;
	    RECT 1235.4000 887.4000 1236.6000 887.5500 ;
	    RECT 1261.8000 887.4000 1263.0000 887.5500 ;
	    RECT 1264.8000 887.7000 1266.3000 888.6000 ;
	    RECT 1269.0000 887.7000 1270.2001 899.7000 ;
	    RECT 1290.6000 899.4000 1291.8000 900.6000 ;
	    RECT 1321.8000 887.7000 1323.0000 899.7000 ;
	    RECT 1187.1000 885.0000 1193.7001 885.9000 ;
	    RECT 1187.1000 884.7000 1188.3000 885.0000 ;
	    RECT 1194.6000 884.4000 1195.8000 885.6000 ;
	    RECT 1196.7001 885.0000 1222.2001 885.9000 ;
	    RECT 1231.2001 885.0000 1232.4000 885.9000 ;
	    RECT 1221.0000 884.1000 1222.2001 885.0000 ;
	    RECT 973.8000 882.4500 975.0000 882.6000 ;
	    RECT 959.5500 881.5500 975.0000 882.4500 ;
	    RECT 973.8000 881.4000 975.0000 881.5500 ;
	    RECT 988.2000 882.4500 989.4000 882.6000 ;
	    RECT 993.0000 882.4500 994.2000 882.6000 ;
	    RECT 988.2000 881.5500 994.2000 882.4500 ;
	    RECT 988.2000 881.4000 989.4000 881.5500 ;
	    RECT 993.0000 881.4000 994.2000 881.5500 ;
	    RECT 925.8000 880.2000 927.0000 880.5000 ;
	    RECT 950.1000 879.3000 951.0000 880.5000 ;
	    RECT 952.5000 879.3000 957.9000 879.9000 ;
	    RECT 959.4000 879.4500 960.6000 879.6000 ;
	    RECT 971.4000 879.4500 972.6000 879.6000 ;
	    RECT 887.4000 873.3000 888.6000 879.3000 ;
	    RECT 889.8000 879.0000 895.8000 879.3000 ;
	    RECT 889.8000 873.3000 891.0000 879.0000 ;
	    RECT 892.2000 873.3000 893.4000 878.1000 ;
	    RECT 894.6000 873.3000 895.8000 879.0000 ;
	    RECT 921.9000 878.4000 924.6000 879.3000 ;
	    RECT 921.9000 873.3000 923.1000 878.4000 ;
	    RECT 925.8000 873.3000 927.0000 879.3000 ;
	    RECT 949.8000 873.3000 951.0000 879.3000 ;
	    RECT 952.2000 879.0000 958.2000 879.3000 ;
	    RECT 952.2000 873.3000 953.4000 879.0000 ;
	    RECT 954.6000 873.3000 955.8000 878.1000 ;
	    RECT 957.0000 873.3000 958.2000 879.0000 ;
	    RECT 959.4000 878.5500 972.6000 879.4500 ;
	    RECT 959.4000 878.4000 960.6000 878.5500 ;
	    RECT 971.4000 878.4000 972.6000 878.5500 ;
	    RECT 971.4000 877.2000 972.6000 877.5000 ;
	    RECT 971.4000 873.3000 972.6000 876.3000 ;
	    RECT 973.8000 873.3000 975.0000 880.5000 ;
	    RECT 993.0000 880.2000 994.2000 880.5000 ;
	    RECT 995.4000 879.3000 996.6000 883.5000 ;
	    RECT 1029.0000 883.2000 1030.2001 883.5000 ;
	    RECT 1033.8000 883.2000 1035.0000 883.5000 ;
	    RECT 1026.6000 881.4000 1027.8000 882.6000 ;
	    RECT 1029.0000 881.4000 1030.5000 882.3000 ;
	    RECT 1031.4000 881.4000 1032.6000 882.6000 ;
	    RECT 1029.0000 879.3000 1029.9000 881.4000 ;
	    RECT 1035.0000 880.8000 1035.3000 882.3000 ;
	    RECT 1036.2001 881.4000 1037.4000 882.6000 ;
	    RECT 1038.6000 882.4500 1039.8000 882.6000 ;
	    RECT 1050.6000 882.4500 1051.8000 882.6000 ;
	    RECT 1038.6000 881.5500 1051.8000 882.4500 ;
	    RECT 1038.6000 881.4000 1039.8000 881.5500 ;
	    RECT 1050.6000 881.4000 1051.8000 881.5500 ;
	    RECT 1185.0000 882.3000 1198.2001 883.5000 ;
	    RECT 1199.1000 882.9000 1202.1000 884.1000 ;
	    RECT 1207.8000 882.9000 1212.6000 884.1000 ;
	    RECT 1031.7001 879.3000 1037.1000 879.9000 ;
	    RECT 993.0000 873.3000 994.2000 879.3000 ;
	    RECT 995.4000 878.4000 998.1000 879.3000 ;
	    RECT 996.9000 873.3000 998.1000 878.4000 ;
	    RECT 1026.6000 874.2000 1027.8000 879.3000 ;
	    RECT 1029.0000 875.1000 1030.2001 879.3000 ;
	    RECT 1031.4000 879.0000 1037.4000 879.3000 ;
	    RECT 1031.4000 874.2000 1032.6000 879.0000 ;
	    RECT 1026.6000 873.3000 1032.6000 874.2000 ;
	    RECT 1033.8000 873.3000 1035.0000 878.1000 ;
	    RECT 1036.2001 873.3000 1037.4000 879.0000 ;
	    RECT 1050.6000 873.3000 1051.8000 880.5000 ;
	    RECT 1053.0000 878.4000 1054.2001 879.6000 ;
	    RECT 1053.0000 877.2000 1054.2001 877.5000 ;
	    RECT 1053.0000 873.3000 1054.2001 876.3000 ;
	    RECT 1185.0000 873.3000 1186.2001 882.3000 ;
	    RECT 1188.6000 880.2000 1193.1000 881.4000 ;
	    RECT 1191.9000 879.3000 1193.1000 880.2000 ;
	    RECT 1200.9000 879.3000 1202.1000 882.9000 ;
	    RECT 1204.2001 881.4000 1205.4000 882.6000 ;
	    RECT 1212.0000 881.7000 1213.2001 882.0000 ;
	    RECT 1206.6000 880.8000 1213.2001 881.7000 ;
	    RECT 1206.6000 880.5000 1207.8000 880.8000 ;
	    RECT 1204.2001 880.2000 1205.4000 880.5000 ;
	    RECT 1216.2001 879.6000 1217.4000 883.8000 ;
	    RECT 1224.9000 882.9000 1230.6000 884.1000 ;
	    RECT 1224.9000 881.1000 1226.1000 882.9000 ;
	    RECT 1231.5000 882.0000 1232.4000 885.0000 ;
	    RECT 1206.6000 879.3000 1207.8000 879.6000 ;
	    RECT 1189.8000 873.3000 1191.0000 879.3000 ;
	    RECT 1191.9000 878.1000 1195.8000 879.3000 ;
	    RECT 1200.9000 878.4000 1207.8000 879.3000 ;
	    RECT 1209.0000 878.4000 1210.2001 879.6000 ;
	    RECT 1211.1000 878.4000 1211.4000 879.6000 ;
	    RECT 1215.9000 878.4000 1217.4000 879.6000 ;
	    RECT 1223.4000 880.2000 1226.1000 881.1000 ;
	    RECT 1230.6000 881.1000 1232.4000 882.0000 ;
	    RECT 1223.4000 879.3000 1224.6000 880.2000 ;
	    RECT 1194.6000 873.3000 1195.8000 878.1000 ;
	    RECT 1221.0000 878.1000 1224.6000 879.3000 ;
	    RECT 1197.0000 873.3000 1198.2001 877.5000 ;
	    RECT 1199.4000 873.3000 1200.6000 877.5000 ;
	    RECT 1201.8000 873.3000 1203.0000 877.5000 ;
	    RECT 1204.2001 873.3000 1205.4000 876.3000 ;
	    RECT 1206.6000 873.3000 1207.8000 877.5000 ;
	    RECT 1209.0000 873.3000 1210.2001 876.3000 ;
	    RECT 1211.4000 873.3000 1212.6000 877.5000 ;
	    RECT 1213.8000 873.3000 1215.0000 877.5000 ;
	    RECT 1216.2001 873.3000 1217.4000 877.5000 ;
	    RECT 1218.6000 873.3000 1219.8000 877.5000 ;
	    RECT 1221.0000 873.3000 1222.2001 878.1000 ;
	    RECT 1225.8000 873.3000 1227.0000 879.3000 ;
	    RECT 1230.6000 873.3000 1231.8000 881.1000 ;
	    RECT 1233.3000 880.2000 1234.5000 886.8000 ;
	    RECT 1264.8000 882.6000 1265.7001 887.7000 ;
	    RECT 1324.2001 886.8000 1325.4000 899.7000 ;
	    RECT 1326.6000 887.7000 1327.8000 899.7000 ;
	    RECT 1329.0000 886.8000 1330.2001 899.7000 ;
	    RECT 1331.4000 887.7000 1332.6000 899.7000 ;
	    RECT 1333.8000 886.8000 1335.0000 899.7000 ;
	    RECT 1336.2001 887.7000 1337.4000 899.7000 ;
	    RECT 1338.6000 886.8000 1339.8000 899.7000 ;
	    RECT 1341.0000 887.7000 1342.2001 899.7000 ;
	    RECT 1375.5000 893.7000 1376.7001 899.7000 ;
	    RECT 1375.8000 890.4000 1377.0000 891.6000 ;
	    RECT 1375.8000 889.5000 1376.7001 890.4000 ;
	    RECT 1377.9000 888.6000 1379.1000 899.7000 ;
	    RECT 1374.6000 887.4000 1375.8000 888.6000 ;
	    RECT 1377.6000 887.7000 1379.1000 888.6000 ;
	    RECT 1381.8000 887.7000 1383.0000 899.7000 ;
	    RECT 1509.0000 893.7000 1510.2001 899.7000 ;
	    RECT 1511.4000 894.6000 1512.6000 899.7000 ;
	    RECT 1511.1000 893.7000 1512.6000 894.6000 ;
	    RECT 1513.8000 893.7000 1515.0000 900.6000 ;
	    RECT 1511.1000 892.8000 1512.0000 893.7000 ;
	    RECT 1516.2001 892.8000 1517.4000 899.7000 ;
	    RECT 1518.6000 893.7000 1519.8000 899.7000 ;
	    RECT 1521.0000 895.5000 1522.2001 899.7000 ;
	    RECT 1523.4000 895.5000 1524.6000 899.7000 ;
	    RECT 1509.0000 891.9000 1512.0000 892.8000 ;
	    RECT 1321.8000 886.5000 1325.4000 886.8000 ;
	    RECT 1323.9000 885.6000 1325.4000 886.5000 ;
	    RECT 1326.9000 885.6000 1330.2001 886.8000 ;
	    RECT 1331.7001 885.6000 1335.0000 886.8000 ;
	    RECT 1337.1000 885.6000 1339.8000 886.8000 ;
	    RECT 1266.6000 884.4000 1267.8000 885.6000 ;
	    RECT 1317.0000 885.4500 1318.2001 885.6000 ;
	    RECT 1321.8000 885.4500 1323.0000 885.6000 ;
	    RECT 1317.0000 884.5500 1323.0000 885.4500 ;
	    RECT 1317.0000 884.4000 1318.2001 884.5500 ;
	    RECT 1321.8000 884.4000 1323.0000 884.5500 ;
	    RECT 1326.9000 883.5000 1328.1000 885.6000 ;
	    RECT 1331.7001 883.5000 1332.9000 885.6000 ;
	    RECT 1337.1000 883.5000 1338.3000 885.6000 ;
	    RECT 1341.0000 885.4500 1342.2001 885.6000 ;
	    RECT 1341.0000 884.5500 1344.4501 885.4500 ;
	    RECT 1341.0000 884.4000 1342.2001 884.5500 ;
	    RECT 1266.6000 883.2000 1267.8000 883.5000 ;
	    RECT 1237.8000 882.4500 1239.0000 882.6000 ;
	    RECT 1261.8000 882.4500 1263.0000 882.6000 ;
	    RECT 1237.8000 881.5500 1263.0000 882.4500 ;
	    RECT 1237.8000 881.4000 1239.0000 881.5500 ;
	    RECT 1261.8000 881.4000 1263.0000 881.5500 ;
	    RECT 1263.9000 881.4000 1265.7001 882.6000 ;
	    RECT 1269.0000 882.4500 1270.2001 882.6000 ;
	    RECT 1290.6000 882.4500 1291.8000 882.6000 ;
	    RECT 1267.8000 880.8000 1268.1000 882.3000 ;
	    RECT 1269.0000 881.5500 1291.8000 882.4500 ;
	    RECT 1269.0000 881.4000 1270.2001 881.5500 ;
	    RECT 1290.6000 881.4000 1291.8000 881.5500 ;
	    RECT 1321.8000 881.4000 1323.0000 883.5000 ;
	    RECT 1324.2001 882.3000 1328.1000 883.5000 ;
	    RECT 1329.3000 882.3000 1332.9000 883.5000 ;
	    RECT 1334.4000 882.3000 1338.3000 883.5000 ;
	    RECT 1339.5000 882.3000 1340.1000 883.5000 ;
	    RECT 1326.9000 881.4000 1328.1000 882.3000 ;
	    RECT 1331.7001 881.4000 1332.9000 882.3000 ;
	    RECT 1337.1000 881.4000 1338.3000 882.3000 ;
	    RECT 1341.0000 881.4000 1342.2001 882.6000 ;
	    RECT 1343.5500 882.4500 1344.4501 884.5500 ;
	    RECT 1377.6000 882.6000 1378.5000 887.7000 ;
	    RECT 1379.4000 885.4500 1380.6000 885.6000 ;
	    RECT 1415.4000 885.4500 1416.6000 885.6000 ;
	    RECT 1379.4000 884.5500 1416.6000 885.4500 ;
	    RECT 1379.4000 884.4000 1380.6000 884.5500 ;
	    RECT 1415.4000 884.4000 1416.6000 884.5500 ;
	    RECT 1509.0000 883.5000 1510.2001 891.9000 ;
	    RECT 1512.9000 891.6000 1519.2001 892.8000 ;
	    RECT 1525.8000 892.5000 1527.0000 899.7000 ;
	    RECT 1528.2001 893.7000 1529.4000 899.7000 ;
	    RECT 1530.6000 892.5000 1531.8000 899.7000 ;
	    RECT 1533.0000 893.7000 1534.2001 899.7000 ;
	    RECT 1512.9000 891.0000 1513.8000 891.6000 ;
	    RECT 1511.4000 889.8000 1513.8000 891.0000 ;
	    RECT 1518.3000 890.7000 1527.0000 891.6000 ;
	    RECT 1515.3000 889.8000 1517.4000 890.7000 ;
	    RECT 1515.3000 889.5000 1524.6000 889.8000 ;
	    RECT 1516.5000 888.9000 1524.6000 889.5000 ;
	    RECT 1523.4000 888.6000 1524.6000 888.9000 ;
	    RECT 1526.1000 889.5000 1527.0000 890.7000 ;
	    RECT 1527.9000 890.4000 1531.8000 891.6000 ;
	    RECT 1535.4000 890.4000 1536.6000 899.7000 ;
	    RECT 1537.8000 895.5000 1539.0000 899.7000 ;
	    RECT 1540.2001 895.5000 1541.4000 899.7000 ;
	    RECT 1542.6000 895.5000 1543.8000 899.7000 ;
	    RECT 1545.0000 893.7000 1546.2001 899.7000 ;
	    RECT 1540.2001 891.6000 1546.5000 892.8000 ;
	    RECT 1547.4000 891.6000 1548.6000 899.7000 ;
	    RECT 1549.8000 893.7000 1551.0000 899.7000 ;
	    RECT 1552.2001 892.8000 1553.4000 899.7000 ;
	    RECT 1554.6000 893.7000 1555.8000 899.7000 ;
	    RECT 1552.2001 891.9000 1556.1000 892.8000 ;
	    RECT 1557.0000 892.5000 1558.2001 899.7000 ;
	    RECT 1559.4000 893.7000 1560.6000 899.7000 ;
	    RECT 1547.4000 890.4000 1551.3000 891.6000 ;
	    RECT 1537.8000 889.5000 1539.0000 889.8000 ;
	    RECT 1526.1000 888.6000 1539.0000 889.5000 ;
	    RECT 1542.6000 889.5000 1543.8000 889.8000 ;
	    RECT 1555.2001 889.5000 1556.1000 891.9000 ;
	    RECT 1557.0000 891.4500 1558.2001 891.6000 ;
	    RECT 1559.4000 891.4500 1560.6000 891.6000 ;
	    RECT 1557.0000 890.5500 1560.6000 891.4500 ;
	    RECT 1557.0000 890.4000 1558.2001 890.5500 ;
	    RECT 1559.4000 890.4000 1560.6000 890.5500 ;
	    RECT 1542.6000 888.6000 1556.1000 889.5000 ;
	    RECT 1513.8000 887.4000 1515.0000 888.6000 ;
	    RECT 1518.9000 887.7000 1520.1000 888.0000 ;
	    RECT 1515.9000 886.8000 1554.3000 887.7000 ;
	    RECT 1553.1000 886.5000 1554.3000 886.8000 ;
	    RECT 1555.2001 885.9000 1556.1000 888.6000 ;
	    RECT 1557.0000 888.0000 1558.2001 889.5000 ;
	    RECT 1557.0000 886.8000 1558.5000 888.0000 ;
	    RECT 1511.1000 885.0000 1517.7001 885.9000 ;
	    RECT 1511.1000 884.7000 1512.3000 885.0000 ;
	    RECT 1518.6000 884.4000 1519.8000 885.6000 ;
	    RECT 1520.7001 885.0000 1546.2001 885.9000 ;
	    RECT 1555.2001 885.0000 1556.4000 885.9000 ;
	    RECT 1545.0000 884.1000 1546.2001 885.0000 ;
	    RECT 1379.4000 883.2000 1380.6000 883.5000 ;
	    RECT 1374.6000 882.4500 1375.8000 882.6000 ;
	    RECT 1343.5500 881.5500 1375.8000 882.4500 ;
	    RECT 1374.6000 881.4000 1375.8000 881.5500 ;
	    RECT 1376.7001 881.4000 1378.5000 882.6000 ;
	    RECT 1381.8000 882.4500 1383.0000 882.6000 ;
	    RECT 1441.8000 882.4500 1443.0000 882.6000 ;
	    RECT 1233.0000 879.0000 1234.5000 880.2000 ;
	    RECT 1262.1000 879.3000 1263.0000 880.5000 ;
	    RECT 1321.8000 880.2000 1325.4000 881.4000 ;
	    RECT 1326.9000 880.2000 1330.2001 881.4000 ;
	    RECT 1331.7001 880.2000 1335.0000 881.4000 ;
	    RECT 1337.1000 880.2000 1339.8000 881.4000 ;
	    RECT 1380.6000 880.8000 1380.9000 882.3000 ;
	    RECT 1381.8000 881.5500 1443.0000 882.4500 ;
	    RECT 1381.8000 881.4000 1383.0000 881.5500 ;
	    RECT 1441.8000 881.4000 1443.0000 881.5500 ;
	    RECT 1509.0000 882.3000 1522.2001 883.5000 ;
	    RECT 1523.1000 882.9000 1526.1000 884.1000 ;
	    RECT 1531.8000 882.9000 1536.6000 884.1000 ;
	    RECT 1264.5000 879.3000 1269.9000 879.9000 ;
	    RECT 1233.0000 873.3000 1234.2001 879.0000 ;
	    RECT 1235.4000 873.3000 1236.6000 876.3000 ;
	    RECT 1261.8000 873.3000 1263.0000 879.3000 ;
	    RECT 1264.2001 879.0000 1270.2001 879.3000 ;
	    RECT 1264.2001 873.3000 1265.4000 879.0000 ;
	    RECT 1266.6000 873.3000 1267.8000 878.1000 ;
	    RECT 1269.0000 873.3000 1270.2001 879.0000 ;
	    RECT 1321.8000 873.3000 1323.0000 879.3000 ;
	    RECT 1324.2001 873.3000 1325.4000 880.2000 ;
	    RECT 1326.6000 873.3000 1327.8000 879.3000 ;
	    RECT 1329.0000 873.3000 1330.2001 880.2000 ;
	    RECT 1331.4000 873.3000 1332.6000 879.3000 ;
	    RECT 1333.8000 873.3000 1335.0000 880.2000 ;
	    RECT 1336.2001 873.3000 1337.4000 879.3000 ;
	    RECT 1338.6000 873.3000 1339.8000 880.2000 ;
	    RECT 1374.9000 879.3000 1375.8000 880.5000 ;
	    RECT 1377.3000 879.3000 1382.7001 879.9000 ;
	    RECT 1341.0000 873.3000 1342.2001 879.3000 ;
	    RECT 1374.6000 873.3000 1375.8000 879.3000 ;
	    RECT 1377.0000 879.0000 1383.0000 879.3000 ;
	    RECT 1377.0000 873.3000 1378.2001 879.0000 ;
	    RECT 1379.4000 873.3000 1380.6000 878.1000 ;
	    RECT 1381.8000 873.3000 1383.0000 879.0000 ;
	    RECT 1509.0000 873.3000 1510.2001 882.3000 ;
	    RECT 1512.6000 880.2000 1517.1000 881.4000 ;
	    RECT 1515.9000 879.3000 1517.1000 880.2000 ;
	    RECT 1524.9000 879.3000 1526.1000 882.9000 ;
	    RECT 1528.2001 881.4000 1529.4000 882.6000 ;
	    RECT 1536.0000 881.7000 1537.2001 882.0000 ;
	    RECT 1530.6000 880.8000 1537.2001 881.7000 ;
	    RECT 1530.6000 880.5000 1531.8000 880.8000 ;
	    RECT 1528.2001 880.2000 1529.4000 880.5000 ;
	    RECT 1540.2001 879.6000 1541.4000 883.8000 ;
	    RECT 1548.9000 882.9000 1554.6000 884.1000 ;
	    RECT 1548.9000 881.1000 1550.1000 882.9000 ;
	    RECT 1555.5000 882.0000 1556.4000 885.0000 ;
	    RECT 1530.6000 879.3000 1531.8000 879.6000 ;
	    RECT 1513.8000 873.3000 1515.0000 879.3000 ;
	    RECT 1515.9000 878.1000 1519.8000 879.3000 ;
	    RECT 1524.9000 878.4000 1531.8000 879.3000 ;
	    RECT 1533.0000 878.4000 1534.2001 879.6000 ;
	    RECT 1535.1000 878.4000 1535.4000 879.6000 ;
	    RECT 1539.9000 878.4000 1541.4000 879.6000 ;
	    RECT 1547.4000 880.2000 1550.1000 881.1000 ;
	    RECT 1554.6000 881.1000 1556.4000 882.0000 ;
	    RECT 1547.4000 879.3000 1548.6000 880.2000 ;
	    RECT 1518.6000 873.3000 1519.8000 878.1000 ;
	    RECT 1545.0000 878.1000 1548.6000 879.3000 ;
	    RECT 1521.0000 873.3000 1522.2001 877.5000 ;
	    RECT 1523.4000 873.3000 1524.6000 877.5000 ;
	    RECT 1525.8000 873.3000 1527.0000 877.5000 ;
	    RECT 1528.2001 873.3000 1529.4000 876.3000 ;
	    RECT 1530.6000 873.3000 1531.8000 877.5000 ;
	    RECT 1533.0000 873.3000 1534.2001 876.3000 ;
	    RECT 1535.4000 873.3000 1536.6000 877.5000 ;
	    RECT 1537.8000 873.3000 1539.0000 877.5000 ;
	    RECT 1540.2001 873.3000 1541.4000 877.5000 ;
	    RECT 1542.6000 873.3000 1543.8000 877.5000 ;
	    RECT 1545.0000 873.3000 1546.2001 878.1000 ;
	    RECT 1549.8000 873.3000 1551.0000 879.3000 ;
	    RECT 1554.6000 873.3000 1555.8000 881.1000 ;
	    RECT 1557.3000 880.2000 1558.5000 886.8000 ;
	    RECT 1557.0000 879.0000 1558.5000 880.2000 ;
	    RECT 1557.0000 873.3000 1558.2001 879.0000 ;
	    RECT 1559.4000 873.3000 1560.6000 876.3000 ;
	    RECT 1.2000 870.6000 1569.0000 872.4000 ;
	    RECT 19.5000 864.6000 20.7000 869.7000 ;
	    RECT 19.5000 863.7000 22.2000 864.6000 ;
	    RECT 23.4000 863.7000 24.6000 869.7000 ;
	    RECT 47.4000 863.7000 48.6000 869.7000 ;
	    RECT 49.8000 864.0000 51.0000 869.7000 ;
	    RECT 52.2000 864.9000 53.4000 869.7000 ;
	    RECT 54.6000 864.0000 55.8000 869.7000 ;
	    RECT 49.8000 863.7000 55.8000 864.0000 ;
	    RECT 21.0000 859.5000 22.2000 863.7000 ;
	    RECT 23.4000 862.5000 24.6000 862.8000 ;
	    RECT 47.7000 862.5000 48.6000 863.7000 ;
	    RECT 50.1000 863.1000 55.5000 863.7000 ;
	    RECT 69.0000 862.5000 70.2000 869.7000 ;
	    RECT 71.4000 866.7000 72.6000 869.7000 ;
	    RECT 71.4000 865.5000 72.6000 865.8000 ;
	    RECT 91.5000 864.6000 92.7000 869.7000 ;
	    RECT 71.4000 863.4000 72.6000 864.6000 ;
	    RECT 91.5000 863.7000 94.2000 864.6000 ;
	    RECT 95.4000 863.7000 96.6000 869.7000 ;
	    RECT 119.4000 863.7000 120.6000 869.7000 ;
	    RECT 121.8000 864.0000 123.0000 869.7000 ;
	    RECT 124.2000 864.9000 125.4000 869.7000 ;
	    RECT 126.6000 864.0000 127.8000 869.7000 ;
	    RECT 121.8000 863.7000 127.8000 864.0000 ;
	    RECT 150.6000 864.0000 151.8000 869.7000 ;
	    RECT 153.0000 864.9000 154.2000 869.7000 ;
	    RECT 155.4000 864.0000 156.6000 869.7000 ;
	    RECT 150.6000 863.7000 156.6000 864.0000 ;
	    RECT 157.8000 863.7000 159.0000 869.7000 ;
	    RECT 23.4000 861.4500 24.6000 861.6000 ;
	    RECT 25.8000 861.4500 27.0000 861.6000 ;
	    RECT 23.4000 860.5500 27.0000 861.4500 ;
	    RECT 23.4000 860.4000 24.6000 860.5500 ;
	    RECT 25.8000 860.4000 27.0000 860.5500 ;
	    RECT 47.4000 860.4000 48.6000 861.6000 ;
	    RECT 49.5000 860.4000 51.3000 861.6000 ;
	    RECT 53.4000 860.7000 53.7000 862.2000 ;
	    RECT 54.6000 860.4000 55.8000 861.6000 ;
	    RECT 69.0000 861.4500 70.2000 861.6000 ;
	    RECT 57.1500 860.5500 70.2000 861.4500 ;
	    RECT 21.0000 858.4500 22.2000 858.6000 ;
	    RECT 21.0000 857.5500 48.4500 858.4500 ;
	    RECT 21.0000 857.4000 22.2000 857.5500 ;
	    RECT 18.6000 854.4000 19.8000 855.6000 ;
	    RECT 18.6000 853.2000 19.8000 853.5000 ;
	    RECT 18.6000 843.3000 19.8000 849.3000 ;
	    RECT 21.0000 843.3000 22.2000 856.5000 ;
	    RECT 47.5500 855.6000 48.4500 857.5500 ;
	    RECT 47.4000 854.4000 48.6000 855.6000 ;
	    RECT 50.4000 855.3000 51.3000 860.4000 ;
	    RECT 52.2000 859.5000 53.4000 859.8000 ;
	    RECT 52.2000 858.4500 53.4000 858.6000 ;
	    RECT 57.1500 858.4500 58.0500 860.5500 ;
	    RECT 69.0000 860.4000 70.2000 860.5500 ;
	    RECT 93.0000 859.5000 94.2000 863.7000 ;
	    RECT 95.4000 862.5000 96.6000 862.8000 ;
	    RECT 119.7000 862.5000 120.6000 863.7000 ;
	    RECT 122.1000 863.1000 127.5000 863.7000 ;
	    RECT 150.9000 863.1000 156.3000 863.7000 ;
	    RECT 157.8000 862.5000 158.7000 863.7000 ;
	    RECT 172.2000 862.5000 173.4000 869.7000 ;
	    RECT 174.6000 866.7000 175.8000 869.7000 ;
	    RECT 174.6000 865.5000 175.8000 865.8000 ;
	    RECT 174.6000 863.4000 175.8000 864.6000 ;
	    RECT 189.0000 862.5000 190.2000 869.7000 ;
	    RECT 191.4000 866.7000 192.6000 869.7000 ;
	    RECT 191.4000 865.5000 192.6000 865.8000 ;
	    RECT 191.4000 864.4500 192.6000 864.6000 ;
	    RECT 210.6000 864.4500 211.8000 864.6000 ;
	    RECT 191.4000 863.5500 211.8000 864.4500 ;
	    RECT 191.4000 863.4000 192.6000 863.5500 ;
	    RECT 210.6000 863.4000 211.8000 863.5500 ;
	    RECT 213.0000 862.5000 214.2000 869.7000 ;
	    RECT 215.4000 866.7000 216.6000 869.7000 ;
	    RECT 215.4000 865.5000 216.6000 865.8000 ;
	    RECT 215.4000 863.4000 216.6000 864.6000 ;
	    RECT 234.6000 863.7000 235.8000 869.7000 ;
	    RECT 238.5000 864.6000 239.7000 869.7000 ;
	    RECT 261.0000 867.4500 262.2000 867.6000 ;
	    RECT 337.8000 867.4500 339.0000 867.6000 ;
	    RECT 261.0000 866.5500 339.0000 867.4500 ;
	    RECT 261.0000 866.4000 262.2000 866.5500 ;
	    RECT 337.8000 866.4000 339.0000 866.5500 ;
	    RECT 237.0000 863.7000 239.7000 864.6000 ;
	    RECT 234.6000 862.5000 235.8000 862.8000 ;
	    RECT 95.4000 861.4500 96.6000 861.6000 ;
	    RECT 102.6000 861.4500 103.8000 861.6000 ;
	    RECT 95.4000 860.5500 103.8000 861.4500 ;
	    RECT 95.4000 860.4000 96.6000 860.5500 ;
	    RECT 102.6000 860.4000 103.8000 860.5500 ;
	    RECT 119.4000 860.4000 120.6000 861.6000 ;
	    RECT 121.5000 860.4000 123.3000 861.6000 ;
	    RECT 125.4000 860.7000 125.7000 862.2000 ;
	    RECT 126.6000 861.4500 127.8000 861.6000 ;
	    RECT 150.6000 861.4500 151.8000 861.6000 ;
	    RECT 126.6000 860.5500 151.8000 861.4500 ;
	    RECT 152.7000 860.7000 153.0000 862.2000 ;
	    RECT 126.6000 860.4000 127.8000 860.5500 ;
	    RECT 150.6000 860.4000 151.8000 860.5500 ;
	    RECT 155.1000 860.4000 156.9000 861.6000 ;
	    RECT 157.8000 860.4000 159.0000 861.6000 ;
	    RECT 160.2000 861.4500 161.4000 861.6000 ;
	    RECT 172.2000 861.4500 173.4000 861.6000 ;
	    RECT 160.2000 860.5500 173.4000 861.4500 ;
	    RECT 160.2000 860.4000 161.4000 860.5500 ;
	    RECT 172.2000 860.4000 173.4000 860.5500 ;
	    RECT 177.0000 861.4500 178.2000 861.6000 ;
	    RECT 189.0000 861.4500 190.2000 861.6000 ;
	    RECT 177.0000 860.5500 190.2000 861.4500 ;
	    RECT 177.0000 860.4000 178.2000 860.5500 ;
	    RECT 189.0000 860.4000 190.2000 860.5500 ;
	    RECT 213.0000 860.4000 214.2000 861.6000 ;
	    RECT 227.4000 861.4500 228.6000 861.6000 ;
	    RECT 234.6000 861.4500 235.8000 861.6000 ;
	    RECT 227.4000 860.5500 235.8000 861.4500 ;
	    RECT 227.4000 860.4000 228.6000 860.5500 ;
	    RECT 234.6000 860.4000 235.8000 860.5500 ;
	    RECT 52.2000 857.5500 58.0500 858.4500 ;
	    RECT 52.2000 857.4000 53.4000 857.5500 ;
	    RECT 50.4000 854.4000 51.9000 855.3000 ;
	    RECT 48.6000 852.6000 49.5000 853.5000 ;
	    RECT 48.6000 851.4000 49.8000 852.6000 ;
	    RECT 23.4000 843.3000 24.6000 849.3000 ;
	    RECT 48.3000 843.3000 49.5000 849.3000 ;
	    RECT 50.7000 843.3000 51.9000 854.4000 ;
	    RECT 54.6000 843.3000 55.8000 855.3000 ;
	    RECT 69.0000 843.3000 70.2000 859.5000 ;
	    RECT 93.0000 858.4500 94.2000 858.6000 ;
	    RECT 93.0000 857.5500 120.4500 858.4500 ;
	    RECT 93.0000 857.4000 94.2000 857.5500 ;
	    RECT 90.6000 854.4000 91.8000 855.6000 ;
	    RECT 90.6000 853.2000 91.8000 853.5000 ;
	    RECT 71.4000 843.3000 72.6000 849.3000 ;
	    RECT 90.6000 843.3000 91.8000 849.3000 ;
	    RECT 93.0000 843.3000 94.2000 856.5000 ;
	    RECT 119.5500 855.6000 120.4500 857.5500 ;
	    RECT 119.4000 854.4000 120.6000 855.6000 ;
	    RECT 122.4000 855.3000 123.3000 860.4000 ;
	    RECT 124.2000 859.5000 125.4000 859.8000 ;
	    RECT 153.0000 859.5000 154.2000 859.8000 ;
	    RECT 124.2000 858.4500 125.4000 858.6000 ;
	    RECT 126.6000 858.4500 127.8000 858.6000 ;
	    RECT 124.2000 857.5500 127.8000 858.4500 ;
	    RECT 124.2000 857.4000 125.4000 857.5500 ;
	    RECT 126.6000 857.4000 127.8000 857.5500 ;
	    RECT 153.0000 857.4000 154.2000 858.6000 ;
	    RECT 155.1000 855.3000 156.0000 860.4000 ;
	    RECT 157.9500 858.4500 158.8500 860.4000 ;
	    RECT 237.0000 859.5000 238.2000 863.7000 ;
	    RECT 364.2000 860.7000 365.4000 869.7000 ;
	    RECT 369.0000 863.7000 370.2000 869.7000 ;
	    RECT 373.8000 864.9000 375.0000 869.7000 ;
	    RECT 376.2000 865.5000 377.4000 869.7000 ;
	    RECT 378.6000 865.5000 379.8000 869.7000 ;
	    RECT 381.0000 865.5000 382.2000 869.7000 ;
	    RECT 383.4000 866.7000 384.6000 869.7000 ;
	    RECT 385.8000 865.5000 387.0000 869.7000 ;
	    RECT 388.2000 866.7000 389.4000 869.7000 ;
	    RECT 390.6000 865.5000 391.8000 869.7000 ;
	    RECT 393.0000 865.5000 394.2000 869.7000 ;
	    RECT 395.4000 865.5000 396.6000 869.7000 ;
	    RECT 397.8000 865.5000 399.0000 869.7000 ;
	    RECT 371.1000 863.7000 375.0000 864.9000 ;
	    RECT 400.2000 864.9000 401.4000 869.7000 ;
	    RECT 380.1000 863.7000 387.0000 864.6000 ;
	    RECT 371.1000 862.8000 372.3000 863.7000 ;
	    RECT 367.8000 861.6000 372.3000 862.8000 ;
	    RECT 364.2000 859.5000 377.4000 860.7000 ;
	    RECT 380.1000 860.1000 381.3000 863.7000 ;
	    RECT 385.8000 863.4000 387.0000 863.7000 ;
	    RECT 388.2000 863.4000 389.4000 864.6000 ;
	    RECT 390.3000 863.4000 390.6000 864.6000 ;
	    RECT 395.1000 863.4000 396.6000 864.6000 ;
	    RECT 400.2000 863.7000 403.8000 864.9000 ;
	    RECT 405.0000 863.7000 406.2000 869.7000 ;
	    RECT 383.4000 862.5000 384.6000 862.8000 ;
	    RECT 385.8000 862.2000 387.0000 862.5000 ;
	    RECT 383.4000 860.4000 384.6000 861.6000 ;
	    RECT 385.8000 861.3000 392.4000 862.2000 ;
	    RECT 391.2000 861.0000 392.4000 861.3000 ;
	    RECT 167.4000 858.4500 168.6000 858.6000 ;
	    RECT 157.9500 857.5500 168.6000 858.4500 ;
	    RECT 167.4000 857.4000 168.6000 857.5500 ;
	    RECT 122.4000 854.4000 123.9000 855.3000 ;
	    RECT 120.6000 852.6000 121.5000 853.5000 ;
	    RECT 120.6000 851.4000 121.8000 852.6000 ;
	    RECT 95.4000 843.3000 96.6000 849.3000 ;
	    RECT 120.3000 843.3000 121.5000 849.3000 ;
	    RECT 122.7000 843.3000 123.9000 854.4000 ;
	    RECT 126.6000 843.3000 127.8000 855.3000 ;
	    RECT 150.6000 843.3000 151.8000 855.3000 ;
	    RECT 154.5000 854.4000 156.0000 855.3000 ;
	    RECT 157.8000 854.4000 159.0000 855.6000 ;
	    RECT 154.5000 843.3000 155.7000 854.4000 ;
	    RECT 156.9000 852.6000 157.8000 853.5000 ;
	    RECT 156.6000 851.4000 157.8000 852.6000 ;
	    RECT 156.9000 843.3000 158.1000 849.3000 ;
	    RECT 172.2000 843.3000 173.4000 859.5000 ;
	    RECT 174.6000 843.3000 175.8000 849.3000 ;
	    RECT 189.0000 843.3000 190.2000 859.5000 ;
	    RECT 191.4000 843.3000 192.6000 849.3000 ;
	    RECT 213.0000 843.3000 214.2000 859.5000 ;
	    RECT 217.8000 858.4500 219.0000 858.6000 ;
	    RECT 237.0000 858.4500 238.2000 858.6000 ;
	    RECT 217.8000 857.5500 238.2000 858.4500 ;
	    RECT 217.8000 857.4000 219.0000 857.5500 ;
	    RECT 237.0000 857.4000 238.2000 857.5500 ;
	    RECT 215.4000 843.3000 216.6000 849.3000 ;
	    RECT 234.6000 843.3000 235.8000 849.3000 ;
	    RECT 237.0000 843.3000 238.2000 856.5000 ;
	    RECT 239.4000 854.4000 240.6000 855.6000 ;
	    RECT 239.4000 853.2000 240.6000 853.5000 ;
	    RECT 270.6000 852.4500 271.8000 852.6000 ;
	    RECT 289.8000 852.4500 291.0000 852.6000 ;
	    RECT 270.6000 851.5500 291.0000 852.4500 ;
	    RECT 270.6000 851.4000 271.8000 851.5500 ;
	    RECT 289.8000 851.4000 291.0000 851.5500 ;
	    RECT 364.2000 851.1000 365.4000 859.5000 ;
	    RECT 378.3000 858.9000 381.3000 860.1000 ;
	    RECT 387.0000 858.9000 391.8000 860.1000 ;
	    RECT 395.4000 859.2000 396.6000 863.4000 ;
	    RECT 402.6000 862.8000 403.8000 863.7000 ;
	    RECT 402.6000 861.9000 405.3000 862.8000 ;
	    RECT 404.1000 860.1000 405.3000 861.9000 ;
	    RECT 409.8000 861.9000 411.0000 869.7000 ;
	    RECT 412.2000 864.0000 413.4000 869.7000 ;
	    RECT 414.6000 866.7000 415.8000 869.7000 ;
	    RECT 412.2000 862.8000 413.7000 864.0000 ;
	    RECT 409.8000 861.0000 411.6000 861.9000 ;
	    RECT 404.1000 858.9000 409.8000 860.1000 ;
	    RECT 366.3000 858.0000 367.5000 858.3000 ;
	    RECT 366.3000 857.1000 372.9000 858.0000 ;
	    RECT 373.8000 857.4000 375.0000 858.6000 ;
	    RECT 400.2000 858.0000 401.4000 858.9000 ;
	    RECT 410.7000 858.0000 411.6000 861.0000 ;
	    RECT 375.9000 857.1000 401.4000 858.0000 ;
	    RECT 410.4000 857.1000 411.6000 858.0000 ;
	    RECT 408.3000 856.2000 409.5000 856.5000 ;
	    RECT 369.0000 854.4000 370.2000 855.6000 ;
	    RECT 371.1000 855.3000 409.5000 856.2000 ;
	    RECT 374.1000 855.0000 375.3000 855.3000 ;
	    RECT 410.4000 854.4000 411.3000 857.1000 ;
	    RECT 412.5000 856.2000 413.7000 862.8000 ;
	    RECT 426.6000 862.5000 427.8000 869.7000 ;
	    RECT 429.0000 866.7000 430.2000 869.7000 ;
	    RECT 450.6000 866.7000 451.8000 869.7000 ;
	    RECT 429.0000 865.5000 430.2000 865.8000 ;
	    RECT 450.6000 865.5000 451.8000 865.8000 ;
	    RECT 429.0000 864.4500 430.2000 864.6000 ;
	    RECT 431.4000 864.4500 432.6000 864.6000 ;
	    RECT 450.6000 864.4500 451.8000 864.6000 ;
	    RECT 429.0000 863.5500 432.6000 864.4500 ;
	    RECT 429.0000 863.4000 430.2000 863.5500 ;
	    RECT 431.4000 863.4000 432.6000 863.5500 ;
	    RECT 433.9500 863.5500 451.8000 864.4500 ;
	    RECT 426.6000 860.4000 427.8000 861.6000 ;
	    RECT 429.0000 861.4500 430.2000 861.6000 ;
	    RECT 433.9500 861.4500 434.8500 863.5500 ;
	    RECT 450.6000 863.4000 451.8000 863.5500 ;
	    RECT 453.0000 862.5000 454.2000 869.7000 ;
	    RECT 477.0000 864.0000 478.2000 869.7000 ;
	    RECT 479.4000 864.9000 480.6000 869.7000 ;
	    RECT 481.8000 864.0000 483.0000 869.7000 ;
	    RECT 477.0000 863.7000 483.0000 864.0000 ;
	    RECT 484.2000 863.7000 485.4000 869.7000 ;
	    RECT 477.3000 863.1000 482.7000 863.7000 ;
	    RECT 484.2000 862.5000 485.1000 863.7000 ;
	    RECT 498.6000 862.5000 499.8000 869.7000 ;
	    RECT 501.0000 866.7000 502.2000 869.7000 ;
	    RECT 520.2000 866.7000 521.4000 869.7000 ;
	    RECT 522.6000 866.7000 523.8000 869.7000 ;
	    RECT 525.0000 866.7000 526.2000 869.7000 ;
	    RECT 501.0000 865.5000 502.2000 865.8000 ;
	    RECT 501.0000 863.4000 502.2000 864.6000 ;
	    RECT 522.6000 862.5000 523.5000 866.7000 ;
	    RECT 525.0000 865.5000 526.2000 865.8000 ;
	    RECT 525.0000 863.4000 526.2000 864.6000 ;
	    RECT 551.4000 863.7000 552.6000 869.7000 ;
	    RECT 553.8000 864.0000 555.0000 869.7000 ;
	    RECT 556.2000 864.9000 557.4000 869.7000 ;
	    RECT 558.6000 864.0000 559.8000 869.7000 ;
	    RECT 577.8000 866.7000 579.0000 869.7000 ;
	    RECT 580.2000 866.7000 581.4000 869.7000 ;
	    RECT 582.6000 866.7000 583.8000 869.7000 ;
	    RECT 601.8000 866.7000 603.0000 869.7000 ;
	    RECT 604.2000 866.7000 605.4000 869.7000 ;
	    RECT 606.6000 866.7000 607.8000 869.7000 ;
	    RECT 618.6000 866.7000 619.8000 869.7000 ;
	    RECT 553.8000 863.7000 559.8000 864.0000 ;
	    RECT 573.0000 864.4500 574.2000 864.6000 ;
	    RECT 577.8000 864.4500 579.0000 864.6000 ;
	    RECT 551.7000 862.5000 552.6000 863.7000 ;
	    RECT 554.1000 863.1000 559.5000 863.7000 ;
	    RECT 573.0000 863.5500 579.0000 864.4500 ;
	    RECT 573.0000 863.4000 574.2000 863.5500 ;
	    RECT 577.8000 863.4000 579.0000 863.5500 ;
	    RECT 580.2000 862.5000 581.1000 866.7000 ;
	    RECT 582.6000 865.5000 583.8000 865.8000 ;
	    RECT 582.6000 864.4500 583.8000 864.6000 ;
	    RECT 599.4000 864.4500 600.6000 864.6000 ;
	    RECT 582.6000 863.5500 600.6000 864.4500 ;
	    RECT 582.6000 863.4000 583.8000 863.5500 ;
	    RECT 599.4000 863.4000 600.6000 863.5500 ;
	    RECT 604.2000 862.5000 605.1000 866.7000 ;
	    RECT 606.6000 865.5000 607.8000 865.8000 ;
	    RECT 618.6000 865.5000 619.8000 865.8000 ;
	    RECT 606.6000 863.4000 607.8000 864.6000 ;
	    RECT 618.6000 863.4000 619.8000 864.6000 ;
	    RECT 621.0000 862.5000 622.2000 869.7000 ;
	    RECT 648.3000 863.7000 649.5000 869.7000 ;
	    RECT 652.2000 863.7000 653.4000 869.7000 ;
	    RECT 654.6000 866.7000 655.8000 869.7000 ;
	    RECT 654.3000 865.5000 655.5000 865.8000 ;
	    RECT 654.6000 864.4500 655.8000 864.6000 ;
	    RECT 657.0000 864.4500 658.2000 864.6000 ;
	    RECT 429.0000 860.5500 434.8500 861.4500 ;
	    RECT 453.0000 861.4500 454.2000 861.6000 ;
	    RECT 453.0000 860.5500 475.6500 861.4500 ;
	    RECT 429.0000 860.4000 430.2000 860.5500 ;
	    RECT 453.0000 860.4000 454.2000 860.5500 ;
	    RECT 378.6000 854.1000 379.8000 854.4000 ;
	    RECT 371.7000 853.5000 379.8000 854.1000 ;
	    RECT 370.5000 853.2000 379.8000 853.5000 ;
	    RECT 381.3000 853.5000 394.2000 854.4000 ;
	    RECT 366.6000 852.0000 369.0000 853.2000 ;
	    RECT 370.5000 852.3000 372.6000 853.2000 ;
	    RECT 381.3000 852.3000 382.2000 853.5000 ;
	    RECT 393.0000 853.2000 394.2000 853.5000 ;
	    RECT 397.8000 853.5000 411.3000 854.4000 ;
	    RECT 412.2000 855.0000 413.7000 856.2000 ;
	    RECT 412.2000 853.5000 413.4000 855.0000 ;
	    RECT 397.8000 853.2000 399.0000 853.5000 ;
	    RECT 368.1000 851.4000 369.0000 852.0000 ;
	    RECT 373.5000 851.4000 382.2000 852.3000 ;
	    RECT 383.1000 851.4000 387.0000 852.6000 ;
	    RECT 364.2000 850.2000 367.2000 851.1000 ;
	    RECT 368.1000 850.2000 374.4000 851.4000 ;
	    RECT 287.4000 849.4500 288.6000 849.6000 ;
	    RECT 311.4000 849.4500 312.6000 849.6000 ;
	    RECT 239.4000 843.3000 240.6000 849.3000 ;
	    RECT 287.4000 848.5500 312.6000 849.4500 ;
	    RECT 366.3000 849.3000 367.2000 850.2000 ;
	    RECT 287.4000 848.4000 288.6000 848.5500 ;
	    RECT 311.4000 848.4000 312.6000 848.5500 ;
	    RECT 285.0000 846.4500 286.2000 846.6000 ;
	    RECT 294.6000 846.4500 295.8000 846.6000 ;
	    RECT 285.0000 845.5500 295.8000 846.4500 ;
	    RECT 285.0000 845.4000 286.2000 845.5500 ;
	    RECT 294.6000 845.4000 295.8000 845.5500 ;
	    RECT 364.2000 843.3000 365.4000 849.3000 ;
	    RECT 366.3000 848.4000 367.8000 849.3000 ;
	    RECT 366.6000 843.3000 367.8000 848.4000 ;
	    RECT 369.0000 842.4000 370.2000 849.3000 ;
	    RECT 371.4000 843.3000 372.6000 850.2000 ;
	    RECT 373.8000 843.3000 375.0000 849.3000 ;
	    RECT 376.2000 843.3000 377.4000 847.5000 ;
	    RECT 378.6000 843.3000 379.8000 847.5000 ;
	    RECT 381.0000 843.3000 382.2000 850.5000 ;
	    RECT 383.4000 843.3000 384.6000 849.3000 ;
	    RECT 385.8000 843.3000 387.0000 850.5000 ;
	    RECT 388.2000 843.3000 389.4000 849.3000 ;
	    RECT 390.6000 843.3000 391.8000 852.6000 ;
	    RECT 402.6000 851.4000 406.5000 852.6000 ;
	    RECT 395.4000 850.2000 401.7000 851.4000 ;
	    RECT 393.0000 843.3000 394.2000 847.5000 ;
	    RECT 395.4000 843.3000 396.6000 847.5000 ;
	    RECT 397.8000 843.3000 399.0000 847.5000 ;
	    RECT 400.2000 843.3000 401.4000 849.3000 ;
	    RECT 402.6000 843.3000 403.8000 851.4000 ;
	    RECT 410.4000 851.1000 411.3000 853.5000 ;
	    RECT 412.2000 851.4000 413.4000 852.6000 ;
	    RECT 407.4000 850.2000 411.3000 851.1000 ;
	    RECT 405.0000 843.3000 406.2000 849.3000 ;
	    RECT 407.4000 843.3000 408.6000 850.2000 ;
	    RECT 409.8000 843.3000 411.0000 849.3000 ;
	    RECT 412.2000 843.3000 413.4000 850.5000 ;
	    RECT 414.6000 843.3000 415.8000 849.3000 ;
	    RECT 426.6000 843.3000 427.8000 859.5000 ;
	    RECT 429.0000 843.3000 430.2000 849.3000 ;
	    RECT 450.6000 843.3000 451.8000 849.3000 ;
	    RECT 453.0000 843.3000 454.2000 859.5000 ;
	    RECT 474.7500 858.4500 475.6500 860.5500 ;
	    RECT 477.0000 860.4000 478.2000 861.6000 ;
	    RECT 479.1000 860.7000 479.4000 862.2000 ;
	    RECT 481.5000 860.4000 483.3000 861.6000 ;
	    RECT 484.2000 861.4500 485.4000 861.6000 ;
	    RECT 496.2000 861.4500 497.4000 861.6000 ;
	    RECT 484.2000 860.5500 497.4000 861.4500 ;
	    RECT 484.2000 860.4000 485.4000 860.5500 ;
	    RECT 496.2000 860.4000 497.4000 860.5500 ;
	    RECT 498.6000 861.4500 499.8000 861.6000 ;
	    RECT 517.8000 861.4500 519.0000 861.6000 ;
	    RECT 498.6000 860.5500 519.0000 861.4500 ;
	    RECT 498.6000 860.4000 499.8000 860.5500 ;
	    RECT 517.8000 860.4000 519.0000 860.5500 ;
	    RECT 522.6000 861.4500 523.8000 861.6000 ;
	    RECT 549.0000 861.4500 550.2000 861.6000 ;
	    RECT 522.6000 860.5500 550.2000 861.4500 ;
	    RECT 522.6000 860.4000 523.8000 860.5500 ;
	    RECT 549.0000 860.4000 550.2000 860.5500 ;
	    RECT 551.4000 860.4000 552.6000 861.6000 ;
	    RECT 553.5000 860.4000 555.3000 861.6000 ;
	    RECT 557.4000 860.7000 557.7000 862.2000 ;
	    RECT 558.6000 861.4500 559.8000 861.6000 ;
	    RECT 563.4000 861.4500 564.6000 861.6000 ;
	    RECT 558.6000 860.5500 564.6000 861.4500 ;
	    RECT 558.6000 860.4000 559.8000 860.5500 ;
	    RECT 563.4000 860.4000 564.6000 860.5500 ;
	    RECT 580.2000 861.4500 581.4000 861.6000 ;
	    RECT 604.2000 861.4500 605.4000 861.6000 ;
	    RECT 613.8000 861.4500 615.0000 861.6000 ;
	    RECT 580.2000 860.5500 602.8500 861.4500 ;
	    RECT 580.2000 860.4000 581.4000 860.5500 ;
	    RECT 479.4000 859.5000 480.6000 859.8000 ;
	    RECT 479.4000 858.4500 480.6000 858.6000 ;
	    RECT 474.7500 857.5500 480.6000 858.4500 ;
	    RECT 479.4000 857.4000 480.6000 857.5500 ;
	    RECT 481.5000 855.3000 482.4000 860.4000 ;
	    RECT 477.0000 843.3000 478.2000 855.3000 ;
	    RECT 480.9000 854.4000 482.4000 855.3000 ;
	    RECT 484.2000 854.4000 485.4000 855.6000 ;
	    RECT 480.9000 843.3000 482.1000 854.4000 ;
	    RECT 483.3000 852.6000 484.2000 853.5000 ;
	    RECT 483.0000 851.4000 484.2000 852.6000 ;
	    RECT 483.3000 843.3000 484.5000 849.3000 ;
	    RECT 498.6000 843.3000 499.8000 859.5000 ;
	    RECT 501.0000 858.4500 502.2000 858.6000 ;
	    RECT 520.2000 858.4500 521.4000 858.6000 ;
	    RECT 501.0000 857.5500 521.4000 858.4500 ;
	    RECT 501.0000 857.4000 502.2000 857.5500 ;
	    RECT 520.2000 857.4000 521.4000 857.5500 ;
	    RECT 520.2000 856.2000 521.4000 856.5000 ;
	    RECT 522.6000 855.3000 523.5000 859.5000 ;
	    RECT 521.1000 854.1000 523.8000 855.3000 ;
	    RECT 501.0000 843.3000 502.2000 849.3000 ;
	    RECT 521.1000 843.3000 522.3000 854.1000 ;
	    RECT 525.0000 843.3000 526.2000 855.3000 ;
	    RECT 551.4000 854.4000 552.6000 855.6000 ;
	    RECT 554.4000 855.3000 555.3000 860.4000 ;
	    RECT 556.2000 859.5000 557.4000 859.8000 ;
	    RECT 556.2000 857.4000 557.4000 858.6000 ;
	    RECT 577.8000 857.4000 579.0000 858.6000 ;
	    RECT 577.8000 856.2000 579.0000 856.5000 ;
	    RECT 580.2000 855.3000 581.1000 859.5000 ;
	    RECT 601.9500 858.6000 602.8500 860.5500 ;
	    RECT 604.2000 860.5500 615.0000 861.4500 ;
	    RECT 604.2000 860.4000 605.4000 860.5500 ;
	    RECT 613.8000 860.4000 615.0000 860.5500 ;
	    RECT 621.0000 861.4500 622.2000 861.6000 ;
	    RECT 649.8000 861.4500 651.0000 861.6000 ;
	    RECT 621.0000 860.5500 651.0000 861.4500 ;
	    RECT 621.0000 860.4000 622.2000 860.5500 ;
	    RECT 649.8000 860.4000 651.0000 860.5500 ;
	    RECT 601.8000 857.4000 603.0000 858.6000 ;
	    RECT 601.8000 856.2000 603.0000 856.5000 ;
	    RECT 604.2000 855.3000 605.1000 859.5000 ;
	    RECT 554.4000 854.4000 555.9000 855.3000 ;
	    RECT 552.6000 852.6000 553.5000 853.5000 ;
	    RECT 552.6000 851.4000 553.8000 852.6000 ;
	    RECT 552.3000 843.3000 553.5000 849.3000 ;
	    RECT 554.7000 843.3000 555.9000 854.4000 ;
	    RECT 558.6000 843.3000 559.8000 855.3000 ;
	    RECT 578.7000 854.1000 581.4000 855.3000 ;
	    RECT 578.7000 843.3000 579.9000 854.1000 ;
	    RECT 582.6000 843.3000 583.8000 855.3000 ;
	    RECT 602.7000 854.1000 605.4000 855.3000 ;
	    RECT 602.7000 843.3000 603.9000 854.1000 ;
	    RECT 606.6000 843.3000 607.8000 855.3000 ;
	    RECT 618.6000 843.3000 619.8000 849.3000 ;
	    RECT 621.0000 843.3000 622.2000 859.5000 ;
	    RECT 649.8000 859.2000 651.0000 859.5000 ;
	    RECT 647.4000 857.4000 648.6000 858.6000 ;
	    RECT 652.2000 858.3000 653.1000 863.7000 ;
	    RECT 654.6000 863.5500 658.2000 864.4500 ;
	    RECT 685.8000 864.0000 687.0000 869.7000 ;
	    RECT 688.2000 864.9000 689.4000 869.7000 ;
	    RECT 690.6000 864.0000 691.8000 869.7000 ;
	    RECT 685.8000 863.7000 691.8000 864.0000 ;
	    RECT 693.0000 863.7000 694.2000 869.7000 ;
	    RECT 707.4000 866.7000 708.6000 869.7000 ;
	    RECT 707.4000 865.5000 708.6000 865.8000 ;
	    RECT 654.6000 863.4000 655.8000 863.5500 ;
	    RECT 657.0000 863.4000 658.2000 863.5500 ;
	    RECT 686.1000 863.1000 691.5000 863.7000 ;
	    RECT 693.0000 862.5000 693.9000 863.7000 ;
	    RECT 707.4000 863.4000 708.6000 864.6000 ;
	    RECT 709.8000 862.5000 711.0000 869.7000 ;
	    RECT 729.0000 863.7000 730.2000 869.7000 ;
	    RECT 732.9000 864.6000 734.1000 869.7000 ;
	    RECT 753.0000 866.7000 754.2000 869.7000 ;
	    RECT 755.4000 866.7000 756.6000 869.7000 ;
	    RECT 757.8000 866.7000 759.0000 869.7000 ;
	    RECT 889.8000 866.7000 891.0000 869.7000 ;
	    RECT 753.0000 865.5000 754.2000 865.8000 ;
	    RECT 731.4000 863.7000 734.1000 864.6000 ;
	    RECT 729.0000 862.5000 730.2000 862.8000 ;
	    RECT 685.8000 860.4000 687.0000 861.6000 ;
	    RECT 687.9000 860.7000 688.2000 862.2000 ;
	    RECT 690.3000 860.4000 692.1000 861.6000 ;
	    RECT 693.0000 861.4500 694.2000 861.6000 ;
	    RECT 705.0000 861.4500 706.2000 861.6000 ;
	    RECT 693.0000 860.5500 706.2000 861.4500 ;
	    RECT 693.0000 860.4000 694.2000 860.5500 ;
	    RECT 705.0000 860.4000 706.2000 860.5500 ;
	    RECT 709.8000 861.4500 711.0000 861.6000 ;
	    RECT 724.2000 861.4500 725.4000 861.6000 ;
	    RECT 709.8000 860.5500 725.4000 861.4500 ;
	    RECT 709.8000 860.4000 711.0000 860.5500 ;
	    RECT 724.2000 860.4000 725.4000 860.5500 ;
	    RECT 729.0000 860.4000 730.2000 861.6000 ;
	    RECT 688.2000 859.5000 689.4000 859.8000 ;
	    RECT 654.6000 858.4500 655.8000 858.6000 ;
	    RECT 671.4000 858.4500 672.6000 858.6000 ;
	    RECT 649.5000 856.8000 649.8000 858.3000 ;
	    RECT 652.2000 857.4000 653.7000 858.3000 ;
	    RECT 654.6000 857.5500 672.6000 858.4500 ;
	    RECT 654.6000 857.4000 655.8000 857.5500 ;
	    RECT 671.4000 857.4000 672.6000 857.5500 ;
	    RECT 673.8000 858.4500 675.0000 858.6000 ;
	    RECT 688.2000 858.4500 689.4000 858.6000 ;
	    RECT 673.8000 857.5500 689.4000 858.4500 ;
	    RECT 673.8000 857.4000 675.0000 857.5500 ;
	    RECT 688.2000 857.4000 689.4000 857.5500 ;
	    RECT 654.6000 855.3000 655.5000 856.5000 ;
	    RECT 690.3000 855.3000 691.2000 860.4000 ;
	    RECT 731.4000 859.5000 732.6000 863.7000 ;
	    RECT 753.0000 863.4000 754.2000 864.6000 ;
	    RECT 755.7000 862.5000 756.6000 866.7000 ;
	    RECT 892.2000 864.0000 893.4000 869.7000 ;
	    RECT 891.9000 862.8000 893.4000 864.0000 ;
	    RECT 755.4000 861.4500 756.6000 861.6000 ;
	    RECT 784.2000 861.4500 785.4000 861.6000 ;
	    RECT 755.4000 860.5500 785.4000 861.4500 ;
	    RECT 755.4000 860.4000 756.6000 860.5500 ;
	    RECT 784.2000 860.4000 785.4000 860.5500 ;
	    RECT 647.4000 854.4000 653.4000 855.3000 ;
	    RECT 647.4000 843.3000 648.6000 854.4000 ;
	    RECT 649.8000 843.3000 651.0000 853.5000 ;
	    RECT 652.2000 843.3000 653.4000 854.4000 ;
	    RECT 654.6000 843.3000 655.8000 855.3000 ;
	    RECT 685.8000 843.3000 687.0000 855.3000 ;
	    RECT 689.7000 854.4000 691.2000 855.3000 ;
	    RECT 693.0000 855.4500 694.2000 855.6000 ;
	    RECT 707.4000 855.4500 708.6000 855.6000 ;
	    RECT 693.0000 854.5500 708.6000 855.4500 ;
	    RECT 693.0000 854.4000 694.2000 854.5500 ;
	    RECT 707.4000 854.4000 708.6000 854.5500 ;
	    RECT 689.7000 843.3000 690.9000 854.4000 ;
	    RECT 692.1000 852.6000 693.0000 853.5000 ;
	    RECT 691.8000 851.4000 693.0000 852.6000 ;
	    RECT 692.1000 843.3000 693.3000 849.3000 ;
	    RECT 707.4000 843.3000 708.6000 849.3000 ;
	    RECT 709.8000 843.3000 711.0000 859.5000 ;
	    RECT 731.4000 858.4500 732.6000 858.6000 ;
	    RECT 753.0000 858.4500 754.2000 858.6000 ;
	    RECT 731.4000 857.5500 754.2000 858.4500 ;
	    RECT 731.4000 857.4000 732.6000 857.5500 ;
	    RECT 753.0000 857.4000 754.2000 857.5500 ;
	    RECT 729.0000 843.3000 730.2000 849.3000 ;
	    RECT 731.4000 843.3000 732.6000 856.5000 ;
	    RECT 733.8000 854.4000 735.0000 855.6000 ;
	    RECT 755.7000 855.3000 756.6000 859.5000 ;
	    RECT 757.8000 857.4000 759.0000 858.6000 ;
	    RECT 757.8000 856.2000 759.0000 856.5000 ;
	    RECT 891.9000 856.2000 893.1000 862.8000 ;
	    RECT 894.6000 861.9000 895.8000 869.7000 ;
	    RECT 899.4000 863.7000 900.6000 869.7000 ;
	    RECT 904.2000 864.9000 905.4000 869.7000 ;
	    RECT 906.6000 865.5000 907.8000 869.7000 ;
	    RECT 909.0000 865.5000 910.2000 869.7000 ;
	    RECT 911.4000 865.5000 912.6000 869.7000 ;
	    RECT 913.8000 865.5000 915.0000 869.7000 ;
	    RECT 916.2000 866.7000 917.4000 869.7000 ;
	    RECT 918.6000 865.5000 919.8000 869.7000 ;
	    RECT 921.0000 866.7000 922.2000 869.7000 ;
	    RECT 923.4000 865.5000 924.6000 869.7000 ;
	    RECT 925.8000 865.5000 927.0000 869.7000 ;
	    RECT 928.2000 865.5000 929.4000 869.7000 ;
	    RECT 901.8000 863.7000 905.4000 864.9000 ;
	    RECT 930.6000 864.9000 931.8000 869.7000 ;
	    RECT 901.8000 862.8000 903.0000 863.7000 ;
	    RECT 894.0000 861.0000 895.8000 861.9000 ;
	    RECT 900.3000 861.9000 903.0000 862.8000 ;
	    RECT 909.0000 863.4000 910.5000 864.6000 ;
	    RECT 915.0000 863.4000 915.3000 864.6000 ;
	    RECT 916.2000 863.4000 917.4000 864.6000 ;
	    RECT 918.6000 863.7000 925.5000 864.6000 ;
	    RECT 930.6000 863.7000 934.5000 864.9000 ;
	    RECT 935.4000 863.7000 936.6000 869.7000 ;
	    RECT 918.6000 863.4000 919.8000 863.7000 ;
	    RECT 894.0000 858.0000 894.9000 861.0000 ;
	    RECT 900.3000 860.1000 901.5000 861.9000 ;
	    RECT 895.8000 858.9000 901.5000 860.1000 ;
	    RECT 909.0000 859.2000 910.2000 863.4000 ;
	    RECT 921.0000 862.5000 922.2000 862.8000 ;
	    RECT 918.6000 862.2000 919.8000 862.5000 ;
	    RECT 913.2000 861.3000 919.8000 862.2000 ;
	    RECT 913.2000 861.0000 914.4000 861.3000 ;
	    RECT 921.0000 860.4000 922.2000 861.6000 ;
	    RECT 924.3000 860.1000 925.5000 863.7000 ;
	    RECT 933.3000 862.8000 934.5000 863.7000 ;
	    RECT 933.3000 861.6000 937.8000 862.8000 ;
	    RECT 940.2000 860.7000 941.4000 869.7000 ;
	    RECT 954.6000 862.5000 955.8000 869.7000 ;
	    RECT 957.0000 866.7000 958.2000 869.7000 ;
	    RECT 957.0000 865.5000 958.2000 865.8000 ;
	    RECT 957.0000 864.4500 958.2000 864.6000 ;
	    RECT 969.0000 864.4500 970.2000 864.6000 ;
	    RECT 957.0000 863.5500 970.2000 864.4500 ;
	    RECT 981.0000 863.7000 982.2000 869.7000 ;
	    RECT 983.4000 864.0000 984.6000 869.7000 ;
	    RECT 985.8000 864.9000 987.0000 869.7000 ;
	    RECT 988.2000 864.0000 989.4000 869.7000 ;
	    RECT 983.4000 863.7000 989.4000 864.0000 ;
	    RECT 957.0000 863.4000 958.2000 863.5500 ;
	    RECT 969.0000 863.4000 970.2000 863.5500 ;
	    RECT 981.3000 862.5000 982.2000 863.7000 ;
	    RECT 983.7000 863.1000 989.1000 863.7000 ;
	    RECT 1002.6000 862.5000 1003.8000 869.7000 ;
	    RECT 1005.0000 866.7000 1006.2000 869.7000 ;
	    RECT 1137.0000 866.7000 1138.2001 869.7000 ;
	    RECT 1005.0000 865.5000 1006.2000 865.8000 ;
	    RECT 1005.0000 864.4500 1006.2000 864.6000 ;
	    RECT 1137.0000 864.4500 1138.2001 864.6000 ;
	    RECT 1005.0000 863.5500 1138.2001 864.4500 ;
	    RECT 1139.4000 864.0000 1140.6000 869.7000 ;
	    RECT 1005.0000 863.4000 1006.2000 863.5500 ;
	    RECT 1137.0000 863.4000 1138.2001 863.5500 ;
	    RECT 1139.1000 862.8000 1140.6000 864.0000 ;
	    RECT 913.8000 858.9000 918.6000 860.1000 ;
	    RECT 924.3000 858.9000 927.3000 860.1000 ;
	    RECT 928.2000 859.5000 941.4000 860.7000 ;
	    RECT 949.8000 861.4500 951.0000 861.6000 ;
	    RECT 954.6000 861.4500 955.8000 861.6000 ;
	    RECT 949.8000 860.5500 955.8000 861.4500 ;
	    RECT 949.8000 860.4000 951.0000 860.5500 ;
	    RECT 954.6000 860.4000 955.8000 860.5500 ;
	    RECT 981.0000 860.4000 982.2000 861.6000 ;
	    RECT 983.1000 860.4000 984.9000 861.6000 ;
	    RECT 987.0000 860.7000 987.3000 862.2000 ;
	    RECT 988.2000 860.4000 989.4000 861.6000 ;
	    RECT 1002.6000 861.4500 1003.8000 861.6000 ;
	    RECT 990.7500 860.5500 1003.8000 861.4500 ;
	    RECT 904.2000 858.0000 905.4000 858.9000 ;
	    RECT 894.0000 857.1000 895.2000 858.0000 ;
	    RECT 904.2000 857.1000 929.7000 858.0000 ;
	    RECT 930.6000 857.4000 931.8000 858.6000 ;
	    RECT 938.1000 858.0000 939.3000 858.3000 ;
	    RECT 932.7000 857.1000 939.3000 858.0000 ;
	    RECT 733.8000 853.2000 735.0000 853.5000 ;
	    RECT 733.8000 843.3000 735.0000 849.3000 ;
	    RECT 736.2000 846.4500 737.4000 846.6000 ;
	    RECT 750.6000 846.4500 751.8000 846.6000 ;
	    RECT 736.2000 845.5500 751.8000 846.4500 ;
	    RECT 736.2000 845.4000 737.4000 845.5500 ;
	    RECT 750.6000 845.4000 751.8000 845.5500 ;
	    RECT 753.0000 843.3000 754.2000 855.3000 ;
	    RECT 755.4000 854.1000 758.1000 855.3000 ;
	    RECT 891.9000 855.0000 893.4000 856.2000 ;
	    RECT 756.9000 843.3000 758.1000 854.1000 ;
	    RECT 892.2000 853.5000 893.4000 855.0000 ;
	    RECT 894.3000 854.4000 895.2000 857.1000 ;
	    RECT 896.1000 856.2000 897.3000 856.5000 ;
	    RECT 896.1000 855.3000 934.5000 856.2000 ;
	    RECT 930.3000 855.0000 931.5000 855.3000 ;
	    RECT 935.4000 854.4000 936.6000 855.6000 ;
	    RECT 894.3000 853.5000 907.8000 854.4000 ;
	    RECT 815.4000 852.4500 816.6000 852.6000 ;
	    RECT 861.0000 852.4500 862.2000 852.6000 ;
	    RECT 892.2000 852.4500 893.4000 852.6000 ;
	    RECT 815.4000 851.5500 893.4000 852.4500 ;
	    RECT 815.4000 851.4000 816.6000 851.5500 ;
	    RECT 861.0000 851.4000 862.2000 851.5500 ;
	    RECT 892.2000 851.4000 893.4000 851.5500 ;
	    RECT 894.3000 851.1000 895.2000 853.5000 ;
	    RECT 906.6000 853.2000 907.8000 853.5000 ;
	    RECT 911.4000 853.5000 924.3000 854.4000 ;
	    RECT 911.4000 853.2000 912.6000 853.5000 ;
	    RECT 899.1000 851.4000 903.0000 852.6000 ;
	    RECT 813.0000 849.4500 814.2000 849.6000 ;
	    RECT 882.6000 849.4500 883.8000 849.6000 ;
	    RECT 813.0000 848.5500 883.8000 849.4500 ;
	    RECT 813.0000 848.4000 814.2000 848.5500 ;
	    RECT 882.6000 848.4000 883.8000 848.5500 ;
	    RECT 781.8000 846.4500 783.0000 846.6000 ;
	    RECT 887.4000 846.4500 888.6000 846.6000 ;
	    RECT 781.8000 845.5500 888.6000 846.4500 ;
	    RECT 781.8000 845.4000 783.0000 845.5500 ;
	    RECT 887.4000 845.4000 888.6000 845.5500 ;
	    RECT 889.8000 843.3000 891.0000 849.3000 ;
	    RECT 892.2000 843.3000 893.4000 850.5000 ;
	    RECT 894.3000 850.2000 898.2000 851.1000 ;
	    RECT 894.6000 843.3000 895.8000 849.3000 ;
	    RECT 897.0000 843.3000 898.2000 850.2000 ;
	    RECT 899.4000 843.3000 900.6000 849.3000 ;
	    RECT 901.8000 843.3000 903.0000 851.4000 ;
	    RECT 903.9000 850.2000 910.2000 851.4000 ;
	    RECT 904.2000 843.3000 905.4000 849.3000 ;
	    RECT 906.6000 843.3000 907.8000 847.5000 ;
	    RECT 909.0000 843.3000 910.2000 847.5000 ;
	    RECT 911.4000 843.3000 912.6000 847.5000 ;
	    RECT 913.8000 843.3000 915.0000 852.6000 ;
	    RECT 918.6000 851.4000 922.5000 852.6000 ;
	    RECT 923.4000 852.3000 924.3000 853.5000 ;
	    RECT 925.8000 854.1000 927.0000 854.4000 ;
	    RECT 925.8000 853.5000 933.9000 854.1000 ;
	    RECT 925.8000 853.2000 935.1000 853.5000 ;
	    RECT 933.0000 852.3000 935.1000 853.2000 ;
	    RECT 923.4000 851.4000 932.1000 852.3000 ;
	    RECT 936.6000 852.0000 939.0000 853.2000 ;
	    RECT 936.6000 851.4000 937.5000 852.0000 ;
	    RECT 916.2000 843.3000 917.4000 849.3000 ;
	    RECT 918.6000 843.3000 919.8000 850.5000 ;
	    RECT 921.0000 843.3000 922.2000 849.3000 ;
	    RECT 923.4000 843.3000 924.6000 850.5000 ;
	    RECT 931.2000 850.2000 937.5000 851.4000 ;
	    RECT 940.2000 851.1000 941.4000 859.5000 ;
	    RECT 938.4000 850.2000 941.4000 851.1000 ;
	    RECT 925.8000 843.3000 927.0000 847.5000 ;
	    RECT 928.2000 843.3000 929.4000 847.5000 ;
	    RECT 930.6000 843.3000 931.8000 849.3000 ;
	    RECT 933.0000 843.3000 934.2000 850.2000 ;
	    RECT 938.4000 849.3000 939.3000 850.2000 ;
	    RECT 935.4000 842.4000 936.6000 849.3000 ;
	    RECT 937.8000 848.4000 939.3000 849.3000 ;
	    RECT 937.8000 843.3000 939.0000 848.4000 ;
	    RECT 940.2000 843.3000 941.4000 849.3000 ;
	    RECT 954.6000 843.3000 955.8000 859.5000 ;
	    RECT 978.6000 855.4500 979.8000 855.6000 ;
	    RECT 981.0000 855.4500 982.2000 855.6000 ;
	    RECT 978.6000 854.5500 982.2000 855.4500 ;
	    RECT 978.6000 854.4000 979.8000 854.5500 ;
	    RECT 981.0000 854.4000 982.2000 854.5500 ;
	    RECT 984.0000 855.3000 984.9000 860.4000 ;
	    RECT 985.8000 859.5000 987.0000 859.8000 ;
	    RECT 985.8000 858.4500 987.0000 858.6000 ;
	    RECT 990.7500 858.4500 991.6500 860.5500 ;
	    RECT 1002.6000 860.4000 1003.8000 860.5500 ;
	    RECT 985.8000 857.5500 991.6500 858.4500 ;
	    RECT 985.8000 857.4000 987.0000 857.5500 ;
	    RECT 984.0000 854.4000 985.5000 855.3000 ;
	    RECT 982.2000 852.6000 983.1000 853.5000 ;
	    RECT 982.2000 851.4000 983.4000 852.6000 ;
	    RECT 957.0000 843.3000 958.2000 849.3000 ;
	    RECT 981.9000 843.3000 983.1000 849.3000 ;
	    RECT 984.3000 843.3000 985.5000 854.4000 ;
	    RECT 988.2000 843.3000 989.4000 855.3000 ;
	    RECT 1002.6000 843.3000 1003.8000 859.5000 ;
	    RECT 1139.1000 856.2000 1140.3000 862.8000 ;
	    RECT 1141.8000 861.9000 1143.0000 869.7000 ;
	    RECT 1146.6000 863.7000 1147.8000 869.7000 ;
	    RECT 1151.4000 864.9000 1152.6000 869.7000 ;
	    RECT 1153.8000 865.5000 1155.0000 869.7000 ;
	    RECT 1156.2001 865.5000 1157.4000 869.7000 ;
	    RECT 1158.6000 865.5000 1159.8000 869.7000 ;
	    RECT 1161.0000 865.5000 1162.2001 869.7000 ;
	    RECT 1163.4000 866.7000 1164.6000 869.7000 ;
	    RECT 1165.8000 865.5000 1167.0000 869.7000 ;
	    RECT 1168.2001 866.7000 1169.4000 869.7000 ;
	    RECT 1170.6000 865.5000 1171.8000 869.7000 ;
	    RECT 1173.0000 865.5000 1174.2001 869.7000 ;
	    RECT 1175.4000 865.5000 1176.6000 869.7000 ;
	    RECT 1149.0000 863.7000 1152.6000 864.9000 ;
	    RECT 1177.8000 864.9000 1179.0000 869.7000 ;
	    RECT 1149.0000 862.8000 1150.2001 863.7000 ;
	    RECT 1141.2001 861.0000 1143.0000 861.9000 ;
	    RECT 1147.5000 861.9000 1150.2001 862.8000 ;
	    RECT 1156.2001 863.4000 1157.7001 864.6000 ;
	    RECT 1162.2001 863.4000 1162.5000 864.6000 ;
	    RECT 1163.4000 863.4000 1164.6000 864.6000 ;
	    RECT 1165.8000 863.7000 1172.7001 864.6000 ;
	    RECT 1177.8000 863.7000 1181.7001 864.9000 ;
	    RECT 1182.6000 863.7000 1183.8000 869.7000 ;
	    RECT 1165.8000 863.4000 1167.0000 863.7000 ;
	    RECT 1141.2001 858.0000 1142.1000 861.0000 ;
	    RECT 1147.5000 860.1000 1148.7001 861.9000 ;
	    RECT 1143.0000 858.9000 1148.7001 860.1000 ;
	    RECT 1156.2001 859.2000 1157.4000 863.4000 ;
	    RECT 1168.2001 862.5000 1169.4000 862.8000 ;
	    RECT 1165.8000 862.2000 1167.0000 862.5000 ;
	    RECT 1160.4000 861.3000 1167.0000 862.2000 ;
	    RECT 1160.4000 861.0000 1161.6000 861.3000 ;
	    RECT 1168.2001 860.4000 1169.4000 861.6000 ;
	    RECT 1171.5000 860.1000 1172.7001 863.7000 ;
	    RECT 1180.5000 862.8000 1181.7001 863.7000 ;
	    RECT 1180.5000 861.6000 1185.0000 862.8000 ;
	    RECT 1187.4000 860.7000 1188.6000 869.7000 ;
	    RECT 1206.6000 863.7000 1207.8000 869.7000 ;
	    RECT 1210.5000 864.6000 1211.7001 869.7000 ;
	    RECT 1209.0000 863.7000 1211.7001 864.6000 ;
	    RECT 1230.6000 863.7000 1231.8000 869.7000 ;
	    RECT 1234.5000 864.6000 1235.7001 869.7000 ;
	    RECT 1247.4000 866.7000 1248.6000 869.7000 ;
	    RECT 1247.4000 865.5000 1248.6000 865.8000 ;
	    RECT 1233.0000 863.7000 1235.7001 864.6000 ;
	    RECT 1242.6000 864.4500 1243.8000 864.6000 ;
	    RECT 1247.4000 864.4500 1248.6000 864.6000 ;
	    RECT 1206.6000 862.5000 1207.8000 862.8000 ;
	    RECT 1161.0000 858.9000 1165.8000 860.1000 ;
	    RECT 1171.5000 858.9000 1174.5000 860.1000 ;
	    RECT 1175.4000 859.5000 1188.6000 860.7000 ;
	    RECT 1206.6000 860.4000 1207.8000 861.6000 ;
	    RECT 1209.0000 859.5000 1210.2001 863.7000 ;
	    RECT 1230.6000 862.5000 1231.8000 862.8000 ;
	    RECT 1213.8000 861.4500 1215.0000 861.6000 ;
	    RECT 1218.6000 861.4500 1219.8000 861.6000 ;
	    RECT 1230.6000 861.4500 1231.8000 861.6000 ;
	    RECT 1213.8000 860.5500 1231.8000 861.4500 ;
	    RECT 1213.8000 860.4000 1215.0000 860.5500 ;
	    RECT 1218.6000 860.4000 1219.8000 860.5500 ;
	    RECT 1230.6000 860.4000 1231.8000 860.5500 ;
	    RECT 1233.0000 859.5000 1234.2001 863.7000 ;
	    RECT 1242.6000 863.5500 1248.6000 864.4500 ;
	    RECT 1242.6000 863.4000 1243.8000 863.5500 ;
	    RECT 1247.4000 863.4000 1248.6000 863.5500 ;
	    RECT 1249.8000 862.5000 1251.0000 869.7000 ;
	    RECT 1319.4000 862.5000 1320.6000 869.7000 ;
	    RECT 1321.8000 863.7000 1323.0000 869.7000 ;
	    RECT 1326.0000 867.6000 1327.2001 869.7000 ;
	    RECT 1324.2001 866.7000 1327.2001 867.6000 ;
	    RECT 1329.9000 866.7000 1331.4000 869.7000 ;
	    RECT 1332.6000 866.7000 1333.8000 869.7000 ;
	    RECT 1335.0000 866.7000 1336.2001 869.7000 ;
	    RECT 1338.9000 867.6000 1340.7001 869.7000 ;
	    RECT 1338.6000 866.7000 1340.7001 867.6000 ;
	    RECT 1324.2001 865.5000 1325.4000 866.7000 ;
	    RECT 1332.6000 865.8000 1333.5000 866.7000 ;
	    RECT 1326.6000 864.6000 1327.8000 865.8000 ;
	    RECT 1329.3000 864.9000 1333.5000 865.8000 ;
	    RECT 1338.6000 865.5000 1339.8000 866.7000 ;
	    RECT 1329.3000 864.6000 1330.5000 864.9000 ;
	    RECT 1249.8000 861.4500 1251.0000 861.6000 ;
	    RECT 1266.6000 861.4500 1267.8000 861.6000 ;
	    RECT 1249.8000 860.5500 1267.8000 861.4500 ;
	    RECT 1249.8000 860.4000 1251.0000 860.5500 ;
	    RECT 1266.6000 860.4000 1267.8000 860.5500 ;
	    RECT 1320.6000 860.4000 1320.9000 861.6000 ;
	    RECT 1321.8000 860.4000 1323.0000 861.6000 ;
	    RECT 1326.9000 861.3000 1327.8000 864.6000 ;
	    RECT 1343.4000 864.0000 1344.6000 869.7000 ;
	    RECT 1341.3000 863.1000 1342.5000 863.4000 ;
	    RECT 1345.8000 863.1000 1347.0000 869.7000 ;
	    RECT 1373.1000 864.6000 1374.3000 869.7000 ;
	    RECT 1373.1000 863.7000 1375.8000 864.6000 ;
	    RECT 1377.0000 863.7000 1378.2001 869.7000 ;
	    RECT 1504.2001 866.7000 1505.4000 869.7000 ;
	    RECT 1506.6000 864.0000 1507.8000 869.7000 ;
	    RECT 1341.3000 862.2000 1347.0000 863.1000 ;
	    RECT 1335.3000 861.3000 1336.5000 861.6000 ;
	    RECT 1323.9000 860.4000 1337.1000 861.3000 ;
	    RECT 1325.1000 860.1000 1326.3000 860.4000 ;
	    RECT 1151.4000 858.0000 1152.6000 858.9000 ;
	    RECT 1141.2001 857.1000 1142.4000 858.0000 ;
	    RECT 1151.4000 857.1000 1176.9000 858.0000 ;
	    RECT 1177.8000 857.4000 1179.0000 858.6000 ;
	    RECT 1185.3000 858.0000 1186.5000 858.3000 ;
	    RECT 1179.9000 857.1000 1186.5000 858.0000 ;
	    RECT 1139.1000 855.0000 1140.6000 856.2000 ;
	    RECT 1139.4000 853.5000 1140.6000 855.0000 ;
	    RECT 1141.5000 854.4000 1142.4000 857.1000 ;
	    RECT 1143.3000 856.2000 1144.5000 856.5000 ;
	    RECT 1143.3000 855.3000 1181.7001 856.2000 ;
	    RECT 1177.5000 855.0000 1178.7001 855.3000 ;
	    RECT 1182.6000 854.4000 1183.8000 855.6000 ;
	    RECT 1141.5000 853.5000 1155.0000 854.4000 ;
	    RECT 1137.0000 852.4500 1138.2001 852.6000 ;
	    RECT 1139.4000 852.4500 1140.6000 852.6000 ;
	    RECT 1137.0000 851.5500 1140.6000 852.4500 ;
	    RECT 1137.0000 851.4000 1138.2001 851.5500 ;
	    RECT 1139.4000 851.4000 1140.6000 851.5500 ;
	    RECT 1141.5000 851.1000 1142.4000 853.5000 ;
	    RECT 1153.8000 853.2000 1155.0000 853.5000 ;
	    RECT 1158.6000 853.5000 1171.5000 854.4000 ;
	    RECT 1158.6000 853.2000 1159.8000 853.5000 ;
	    RECT 1146.3000 851.4000 1150.2001 852.6000 ;
	    RECT 1005.0000 843.3000 1006.2000 849.3000 ;
	    RECT 1137.0000 843.3000 1138.2001 849.3000 ;
	    RECT 1139.4000 843.3000 1140.6000 850.5000 ;
	    RECT 1141.5000 850.2000 1145.4000 851.1000 ;
	    RECT 1141.8000 843.3000 1143.0000 849.3000 ;
	    RECT 1144.2001 843.3000 1145.4000 850.2000 ;
	    RECT 1146.6000 843.3000 1147.8000 849.3000 ;
	    RECT 1149.0000 843.3000 1150.2001 851.4000 ;
	    RECT 1151.1000 850.2000 1157.4000 851.4000 ;
	    RECT 1151.4000 843.3000 1152.6000 849.3000 ;
	    RECT 1153.8000 843.3000 1155.0000 847.5000 ;
	    RECT 1156.2001 843.3000 1157.4000 847.5000 ;
	    RECT 1158.6000 843.3000 1159.8000 847.5000 ;
	    RECT 1161.0000 843.3000 1162.2001 852.6000 ;
	    RECT 1165.8000 851.4000 1169.7001 852.6000 ;
	    RECT 1170.6000 852.3000 1171.5000 853.5000 ;
	    RECT 1173.0000 854.1000 1174.2001 854.4000 ;
	    RECT 1173.0000 853.5000 1181.1000 854.1000 ;
	    RECT 1173.0000 853.2000 1182.3000 853.5000 ;
	    RECT 1180.2001 852.3000 1182.3000 853.2000 ;
	    RECT 1170.6000 851.4000 1179.3000 852.3000 ;
	    RECT 1183.8000 852.0000 1186.2001 853.2000 ;
	    RECT 1183.8000 851.4000 1184.7001 852.0000 ;
	    RECT 1163.4000 843.3000 1164.6000 849.3000 ;
	    RECT 1165.8000 843.3000 1167.0000 850.5000 ;
	    RECT 1168.2001 843.3000 1169.4000 849.3000 ;
	    RECT 1170.6000 843.3000 1171.8000 850.5000 ;
	    RECT 1178.4000 850.2000 1184.7001 851.4000 ;
	    RECT 1187.4000 851.1000 1188.6000 859.5000 ;
	    RECT 1209.0000 858.4500 1210.2001 858.6000 ;
	    RECT 1211.4000 858.4500 1212.6000 858.6000 ;
	    RECT 1209.0000 857.5500 1212.6000 858.4500 ;
	    RECT 1209.0000 857.4000 1210.2001 857.5500 ;
	    RECT 1211.4000 857.4000 1212.6000 857.5500 ;
	    RECT 1228.2001 858.4500 1229.4000 858.6000 ;
	    RECT 1233.0000 858.4500 1234.2001 858.6000 ;
	    RECT 1228.2001 857.5500 1234.2001 858.4500 ;
	    RECT 1228.2001 857.4000 1229.4000 857.5500 ;
	    RECT 1233.0000 857.4000 1234.2001 857.5500 ;
	    RECT 1185.6000 850.2000 1188.6000 851.1000 ;
	    RECT 1173.0000 843.3000 1174.2001 847.5000 ;
	    RECT 1175.4000 843.3000 1176.6000 847.5000 ;
	    RECT 1177.8000 843.3000 1179.0000 849.3000 ;
	    RECT 1180.2001 843.3000 1181.4000 850.2000 ;
	    RECT 1185.6000 849.3000 1186.5000 850.2000 ;
	    RECT 1182.6000 842.4000 1183.8000 849.3000 ;
	    RECT 1185.0000 848.4000 1186.5000 849.3000 ;
	    RECT 1185.0000 843.3000 1186.2001 848.4000 ;
	    RECT 1187.4000 843.3000 1188.6000 849.3000 ;
	    RECT 1206.6000 843.3000 1207.8000 849.3000 ;
	    RECT 1209.0000 843.3000 1210.2001 856.5000 ;
	    RECT 1211.4000 855.4500 1212.6000 855.6000 ;
	    RECT 1223.4000 855.4500 1224.6000 855.6000 ;
	    RECT 1211.4000 854.5500 1224.6000 855.4500 ;
	    RECT 1211.4000 854.4000 1212.6000 854.5500 ;
	    RECT 1223.4000 854.4000 1224.6000 854.5500 ;
	    RECT 1211.4000 853.2000 1212.6000 853.5000 ;
	    RECT 1211.4000 843.3000 1212.6000 849.3000 ;
	    RECT 1230.6000 843.3000 1231.8000 849.3000 ;
	    RECT 1233.0000 843.3000 1234.2001 856.5000 ;
	    RECT 1235.4000 855.4500 1236.6000 855.6000 ;
	    RECT 1247.4000 855.4500 1248.6000 855.6000 ;
	    RECT 1235.4000 854.5500 1248.6000 855.4500 ;
	    RECT 1235.4000 854.4000 1236.6000 854.5500 ;
	    RECT 1247.4000 854.4000 1248.6000 854.5500 ;
	    RECT 1235.4000 853.2000 1236.6000 853.5000 ;
	    RECT 1235.4000 843.3000 1236.6000 849.3000 ;
	    RECT 1247.4000 843.3000 1248.6000 849.3000 ;
	    RECT 1249.8000 843.3000 1251.0000 859.5000 ;
	    RECT 1322.7001 858.6000 1323.9000 858.9000 ;
	    RECT 1322.7001 857.7000 1328.1000 858.6000 ;
	    RECT 1329.0000 857.4000 1330.2001 858.6000 ;
	    RECT 1319.4000 856.5000 1327.8000 856.8000 ;
	    RECT 1319.4000 856.2000 1328.1000 856.5000 ;
	    RECT 1319.4000 855.9000 1334.1000 856.2000 ;
	    RECT 1319.4000 843.3000 1320.6000 855.9000 ;
	    RECT 1326.9000 855.3000 1334.1000 855.9000 ;
	    RECT 1321.8000 843.3000 1323.0000 855.0000 ;
	    RECT 1324.2001 853.5000 1332.3000 854.4000 ;
	    RECT 1324.2001 853.2000 1325.4000 853.5000 ;
	    RECT 1331.1000 853.2000 1332.3000 853.5000 ;
	    RECT 1333.2001 853.5000 1334.1000 855.3000 ;
	    RECT 1336.2001 855.6000 1337.1000 860.4000 ;
	    RECT 1345.8000 859.5000 1347.0000 862.2000 ;
	    RECT 1374.6000 859.5000 1375.8000 863.7000 ;
	    RECT 1506.3000 862.8000 1507.8000 864.0000 ;
	    RECT 1377.0000 862.5000 1378.2001 862.8000 ;
	    RECT 1377.0000 861.4500 1378.2001 861.6000 ;
	    RECT 1437.0000 861.4500 1438.2001 861.6000 ;
	    RECT 1377.0000 860.5500 1438.2001 861.4500 ;
	    RECT 1377.0000 860.4000 1378.2001 860.5500 ;
	    RECT 1437.0000 860.4000 1438.2001 860.5500 ;
	    RECT 1338.6000 859.2000 1339.8000 859.5000 ;
	    RECT 1338.6000 858.3000 1344.3000 859.2000 ;
	    RECT 1343.1000 858.0000 1344.3000 858.3000 ;
	    RECT 1345.8000 858.4500 1347.0000 858.6000 ;
	    RECT 1365.0000 858.4500 1366.2001 858.6000 ;
	    RECT 1345.8000 857.5500 1366.2001 858.4500 ;
	    RECT 1345.8000 857.4000 1347.0000 857.5500 ;
	    RECT 1365.0000 857.4000 1366.2001 857.5500 ;
	    RECT 1374.6000 858.4500 1375.8000 858.6000 ;
	    RECT 1377.0000 858.4500 1378.2001 858.6000 ;
	    RECT 1374.6000 857.5500 1378.2001 858.4500 ;
	    RECT 1374.6000 857.4000 1375.8000 857.5500 ;
	    RECT 1377.0000 857.4000 1378.2001 857.5500 ;
	    RECT 1340.7001 857.1000 1341.9000 857.4000 ;
	    RECT 1340.7001 856.5000 1344.9000 857.1000 ;
	    RECT 1340.7001 856.2000 1347.0000 856.5000 ;
	    RECT 1336.2001 854.7000 1339.8000 855.6000 ;
	    RECT 1335.3000 853.5000 1336.5000 853.8000 ;
	    RECT 1333.2001 852.6000 1336.5000 853.5000 ;
	    RECT 1338.9000 853.2000 1339.8000 854.7000 ;
	    RECT 1338.9000 852.0000 1341.0000 853.2000 ;
	    RECT 1329.3000 851.1000 1330.5000 851.4000 ;
	    RECT 1333.5000 851.1000 1334.7001 851.4000 ;
	    RECT 1324.2001 849.3000 1325.4000 850.5000 ;
	    RECT 1329.3000 850.2000 1334.7001 851.1000 ;
	    RECT 1332.6000 849.3000 1333.5000 850.2000 ;
	    RECT 1338.6000 849.3000 1339.8000 850.5000 ;
	    RECT 1324.2001 848.4000 1327.2001 849.3000 ;
	    RECT 1326.0000 843.3000 1327.2001 848.4000 ;
	    RECT 1330.2001 843.3000 1331.4000 849.3000 ;
	    RECT 1332.6000 843.3000 1333.8000 849.3000 ;
	    RECT 1335.0000 843.3000 1336.2001 849.3000 ;
	    RECT 1338.9000 843.3000 1340.7001 849.3000 ;
	    RECT 1343.4000 843.3000 1344.6000 855.3000 ;
	    RECT 1345.8000 843.3000 1347.0000 856.2000 ;
	    RECT 1372.2001 854.4000 1373.4000 855.6000 ;
	    RECT 1372.2001 853.2000 1373.4000 853.5000 ;
	    RECT 1372.2001 843.3000 1373.4000 849.3000 ;
	    RECT 1374.6000 843.3000 1375.8000 856.5000 ;
	    RECT 1506.3000 856.2000 1507.5000 862.8000 ;
	    RECT 1509.0000 861.9000 1510.2001 869.7000 ;
	    RECT 1513.8000 863.7000 1515.0000 869.7000 ;
	    RECT 1518.6000 864.9000 1519.8000 869.7000 ;
	    RECT 1521.0000 865.5000 1522.2001 869.7000 ;
	    RECT 1523.4000 865.5000 1524.6000 869.7000 ;
	    RECT 1525.8000 865.5000 1527.0000 869.7000 ;
	    RECT 1528.2001 865.5000 1529.4000 869.7000 ;
	    RECT 1530.6000 866.7000 1531.8000 869.7000 ;
	    RECT 1533.0000 865.5000 1534.2001 869.7000 ;
	    RECT 1535.4000 866.7000 1536.6000 869.7000 ;
	    RECT 1537.8000 865.5000 1539.0000 869.7000 ;
	    RECT 1540.2001 865.5000 1541.4000 869.7000 ;
	    RECT 1542.6000 865.5000 1543.8000 869.7000 ;
	    RECT 1516.2001 863.7000 1519.8000 864.9000 ;
	    RECT 1545.0000 864.9000 1546.2001 869.7000 ;
	    RECT 1516.2001 862.8000 1517.4000 863.7000 ;
	    RECT 1508.4000 861.0000 1510.2001 861.9000 ;
	    RECT 1514.7001 861.9000 1517.4000 862.8000 ;
	    RECT 1523.4000 863.4000 1524.9000 864.6000 ;
	    RECT 1529.4000 863.4000 1529.7001 864.6000 ;
	    RECT 1530.6000 863.4000 1531.8000 864.6000 ;
	    RECT 1533.0000 863.7000 1539.9000 864.6000 ;
	    RECT 1545.0000 863.7000 1548.9000 864.9000 ;
	    RECT 1549.8000 863.7000 1551.0000 869.7000 ;
	    RECT 1533.0000 863.4000 1534.2001 863.7000 ;
	    RECT 1508.4000 858.0000 1509.3000 861.0000 ;
	    RECT 1514.7001 860.1000 1515.9000 861.9000 ;
	    RECT 1510.2001 858.9000 1515.9000 860.1000 ;
	    RECT 1523.4000 859.2000 1524.6000 863.4000 ;
	    RECT 1535.4000 862.5000 1536.6000 862.8000 ;
	    RECT 1533.0000 862.2000 1534.2001 862.5000 ;
	    RECT 1527.6000 861.3000 1534.2001 862.2000 ;
	    RECT 1527.6000 861.0000 1528.8000 861.3000 ;
	    RECT 1535.4000 860.4000 1536.6000 861.6000 ;
	    RECT 1538.7001 860.1000 1539.9000 863.7000 ;
	    RECT 1547.7001 862.8000 1548.9000 863.7000 ;
	    RECT 1547.7001 861.6000 1552.2001 862.8000 ;
	    RECT 1554.6000 860.7000 1555.8000 869.7000 ;
	    RECT 1528.2001 858.9000 1533.0000 860.1000 ;
	    RECT 1538.7001 858.9000 1541.7001 860.1000 ;
	    RECT 1542.6000 859.5000 1555.8000 860.7000 ;
	    RECT 1518.6000 858.0000 1519.8000 858.9000 ;
	    RECT 1508.4000 857.1000 1509.6000 858.0000 ;
	    RECT 1518.6000 857.1000 1544.1000 858.0000 ;
	    RECT 1545.0000 857.4000 1546.2001 858.6000 ;
	    RECT 1552.5000 858.0000 1553.7001 858.3000 ;
	    RECT 1547.1000 857.1000 1553.7001 858.0000 ;
	    RECT 1506.3000 855.0000 1507.8000 856.2000 ;
	    RECT 1506.6000 853.5000 1507.8000 855.0000 ;
	    RECT 1508.7001 854.4000 1509.6000 857.1000 ;
	    RECT 1510.5000 856.2000 1511.7001 856.5000 ;
	    RECT 1510.5000 855.3000 1548.9000 856.2000 ;
	    RECT 1549.8000 855.4500 1551.0000 855.6000 ;
	    RECT 1552.2001 855.4500 1553.4000 855.6000 ;
	    RECT 1544.7001 855.0000 1545.9000 855.3000 ;
	    RECT 1549.8000 854.5500 1553.4000 855.4500 ;
	    RECT 1549.8000 854.4000 1551.0000 854.5500 ;
	    RECT 1552.2001 854.4000 1553.4000 854.5500 ;
	    RECT 1508.7001 853.5000 1522.2001 854.4000 ;
	    RECT 1432.2001 852.4500 1433.4000 852.6000 ;
	    RECT 1506.6000 852.4500 1507.8000 852.6000 ;
	    RECT 1432.2001 851.5500 1507.8000 852.4500 ;
	    RECT 1432.2001 851.4000 1433.4000 851.5500 ;
	    RECT 1506.6000 851.4000 1507.8000 851.5500 ;
	    RECT 1508.7001 851.1000 1509.6000 853.5000 ;
	    RECT 1521.0000 853.2000 1522.2001 853.5000 ;
	    RECT 1525.8000 853.5000 1538.7001 854.4000 ;
	    RECT 1525.8000 853.2000 1527.0000 853.5000 ;
	    RECT 1513.5000 851.4000 1517.4000 852.6000 ;
	    RECT 1377.0000 843.3000 1378.2001 849.3000 ;
	    RECT 1504.2001 843.3000 1505.4000 849.3000 ;
	    RECT 1506.6000 843.3000 1507.8000 850.5000 ;
	    RECT 1508.7001 850.2000 1512.6000 851.1000 ;
	    RECT 1509.0000 843.3000 1510.2001 849.3000 ;
	    RECT 1511.4000 843.3000 1512.6000 850.2000 ;
	    RECT 1513.8000 843.3000 1515.0000 849.3000 ;
	    RECT 1516.2001 843.3000 1517.4000 851.4000 ;
	    RECT 1518.3000 850.2000 1524.6000 851.4000 ;
	    RECT 1518.6000 843.3000 1519.8000 849.3000 ;
	    RECT 1521.0000 843.3000 1522.2001 847.5000 ;
	    RECT 1523.4000 843.3000 1524.6000 847.5000 ;
	    RECT 1525.8000 843.3000 1527.0000 847.5000 ;
	    RECT 1528.2001 843.3000 1529.4000 852.6000 ;
	    RECT 1533.0000 851.4000 1536.9000 852.6000 ;
	    RECT 1537.8000 852.3000 1538.7001 853.5000 ;
	    RECT 1540.2001 854.1000 1541.4000 854.4000 ;
	    RECT 1540.2001 853.5000 1548.3000 854.1000 ;
	    RECT 1540.2001 853.2000 1549.5000 853.5000 ;
	    RECT 1547.4000 852.3000 1549.5000 853.2000 ;
	    RECT 1537.8000 851.4000 1546.5000 852.3000 ;
	    RECT 1551.0000 852.0000 1553.4000 853.2000 ;
	    RECT 1551.0000 851.4000 1551.9000 852.0000 ;
	    RECT 1530.6000 843.3000 1531.8000 849.3000 ;
	    RECT 1533.0000 843.3000 1534.2001 850.5000 ;
	    RECT 1535.4000 843.3000 1536.6000 849.3000 ;
	    RECT 1537.8000 843.3000 1539.0000 850.5000 ;
	    RECT 1545.6000 850.2000 1551.9000 851.4000 ;
	    RECT 1554.6000 851.1000 1555.8000 859.5000 ;
	    RECT 1552.8000 850.2000 1555.8000 851.1000 ;
	    RECT 1540.2001 843.3000 1541.4000 847.5000 ;
	    RECT 1542.6000 843.3000 1543.8000 847.5000 ;
	    RECT 1545.0000 843.3000 1546.2001 849.3000 ;
	    RECT 1547.4000 843.3000 1548.6000 850.2000 ;
	    RECT 1552.8000 849.3000 1553.7001 850.2000 ;
	    RECT 1549.8000 842.4000 1551.0000 849.3000 ;
	    RECT 1552.2001 848.4000 1553.7001 849.3000 ;
	    RECT 1552.2001 843.3000 1553.4000 848.4000 ;
	    RECT 1554.6000 843.3000 1555.8000 849.3000 ;
	    RECT 1566.6000 842.4000 1567.8000 843.6000 ;
	    RECT 1.2000 840.6000 1569.0000 842.4000 ;
	    RECT 124.2000 833.7000 125.4000 839.7000 ;
	    RECT 126.6000 832.5000 127.8000 839.7000 ;
	    RECT 129.0000 833.7000 130.2000 839.7000 ;
	    RECT 131.4000 832.8000 132.6000 839.7000 ;
	    RECT 133.8000 833.7000 135.0000 839.7000 ;
	    RECT 128.7000 831.9000 132.6000 832.8000 ;
	    RECT 109.8000 831.4500 111.0000 831.6000 ;
	    RECT 126.6000 831.4500 127.8000 831.6000 ;
	    RECT 109.8000 830.5500 127.8000 831.4500 ;
	    RECT 109.8000 830.4000 111.0000 830.5500 ;
	    RECT 126.6000 830.4000 127.8000 830.5500 ;
	    RECT 128.7000 829.5000 129.6000 831.9000 ;
	    RECT 136.2000 831.6000 137.4000 839.7000 ;
	    RECT 138.6000 833.7000 139.8000 839.7000 ;
	    RECT 141.0000 835.5000 142.2000 839.7000 ;
	    RECT 143.4000 835.5000 144.6000 839.7000 ;
	    RECT 145.8000 835.5000 147.0000 839.7000 ;
	    RECT 138.3000 831.6000 144.6000 832.8000 ;
	    RECT 133.5000 830.4000 137.4000 831.6000 ;
	    RECT 148.2000 830.4000 149.4000 839.7000 ;
	    RECT 150.6000 833.7000 151.8000 839.7000 ;
	    RECT 153.0000 832.5000 154.2000 839.7000 ;
	    RECT 155.4000 833.7000 156.6000 839.7000 ;
	    RECT 157.8000 832.5000 159.0000 839.7000 ;
	    RECT 160.2000 835.5000 161.4000 839.7000 ;
	    RECT 162.6000 835.5000 163.8000 839.7000 ;
	    RECT 165.0000 833.7000 166.2000 839.7000 ;
	    RECT 167.4000 832.8000 168.6000 839.7000 ;
	    RECT 169.8000 833.7000 171.0000 840.6000 ;
	    RECT 172.2000 834.6000 173.4000 839.7000 ;
	    RECT 172.2000 833.7000 173.7000 834.6000 ;
	    RECT 174.6000 833.7000 175.8000 839.7000 ;
	    RECT 172.8000 832.8000 173.7000 833.7000 ;
	    RECT 165.6000 831.6000 171.9000 832.8000 ;
	    RECT 172.8000 831.9000 175.8000 832.8000 ;
	    RECT 153.0000 830.4000 156.9000 831.6000 ;
	    RECT 157.8000 830.7000 166.5000 831.6000 ;
	    RECT 171.0000 831.0000 171.9000 831.6000 ;
	    RECT 141.0000 829.5000 142.2000 829.8000 ;
	    RECT 126.6000 828.0000 127.8000 829.5000 ;
	    RECT 126.3000 826.8000 127.8000 828.0000 ;
	    RECT 128.7000 828.6000 142.2000 829.5000 ;
	    RECT 145.8000 829.5000 147.0000 829.8000 ;
	    RECT 157.8000 829.5000 158.7000 830.7000 ;
	    RECT 167.4000 829.8000 169.5000 830.7000 ;
	    RECT 171.0000 829.8000 173.4000 831.0000 ;
	    RECT 145.8000 828.6000 158.7000 829.5000 ;
	    RECT 160.2000 829.5000 169.5000 829.8000 ;
	    RECT 160.2000 828.9000 168.3000 829.5000 ;
	    RECT 160.2000 828.6000 161.4000 828.9000 ;
	    RECT 126.3000 820.2000 127.5000 826.8000 ;
	    RECT 128.7000 825.9000 129.6000 828.6000 ;
	    RECT 164.7000 827.7000 165.9000 828.0000 ;
	    RECT 130.5000 826.8000 168.9000 827.7000 ;
	    RECT 169.8000 827.4000 171.0000 828.6000 ;
	    RECT 130.5000 826.5000 131.7000 826.8000 ;
	    RECT 128.4000 825.0000 129.6000 825.9000 ;
	    RECT 138.6000 825.0000 164.1000 825.9000 ;
	    RECT 128.4000 822.0000 129.3000 825.0000 ;
	    RECT 138.6000 824.1000 139.8000 825.0000 ;
	    RECT 165.0000 824.4000 166.2000 825.6000 ;
	    RECT 167.1000 825.0000 173.7000 825.9000 ;
	    RECT 172.5000 824.7000 173.7000 825.0000 ;
	    RECT 130.2000 822.9000 135.9000 824.1000 ;
	    RECT 128.4000 821.1000 130.2000 822.0000 ;
	    RECT 126.3000 819.0000 127.8000 820.2000 ;
	    RECT 124.2000 813.3000 125.4000 816.3000 ;
	    RECT 126.6000 813.3000 127.8000 819.0000 ;
	    RECT 129.0000 813.3000 130.2000 821.1000 ;
	    RECT 134.7000 821.1000 135.9000 822.9000 ;
	    RECT 134.7000 820.2000 137.4000 821.1000 ;
	    RECT 136.2000 819.3000 137.4000 820.2000 ;
	    RECT 143.4000 819.6000 144.6000 823.8000 ;
	    RECT 148.2000 822.9000 153.0000 824.1000 ;
	    RECT 158.7000 822.9000 161.7000 824.1000 ;
	    RECT 174.6000 823.5000 175.8000 831.9000 ;
	    RECT 213.0000 827.7000 214.2000 839.7000 ;
	    RECT 216.9000 827.7000 219.9000 839.7000 ;
	    RECT 222.6000 827.7000 223.8000 839.7000 ;
	    RECT 215.4000 824.4000 216.6000 825.6000 ;
	    RECT 217.8000 823.5000 218.7000 827.7000 ;
	    RECT 220.2000 824.4000 221.4000 825.6000 ;
	    RECT 222.6000 823.5000 223.8000 823.8000 ;
	    RECT 234.6000 823.5000 235.8000 839.7000 ;
	    RECT 237.0000 833.7000 238.2000 839.7000 ;
	    RECT 251.4000 833.7000 252.6000 839.7000 ;
	    RECT 253.8000 823.5000 255.0000 839.7000 ;
	    RECT 285.0000 827.7000 286.2000 839.7000 ;
	    RECT 288.9000 827.7000 291.9000 839.7000 ;
	    RECT 294.6000 827.7000 295.8000 839.7000 ;
	    RECT 313.8000 833.7000 315.0000 839.7000 ;
	    RECT 313.8000 829.5000 315.0000 829.8000 ;
	    RECT 301.8000 828.4500 303.0000 828.6000 ;
	    RECT 313.8000 828.4500 315.0000 828.6000 ;
	    RECT 287.4000 824.4000 288.6000 825.6000 ;
	    RECT 285.0000 823.5000 286.2000 823.8000 ;
	    RECT 290.1000 823.5000 291.0000 827.7000 ;
	    RECT 301.8000 827.5500 315.0000 828.4500 ;
	    RECT 301.8000 827.4000 303.0000 827.5500 ;
	    RECT 313.8000 827.4000 315.0000 827.5500 ;
	    RECT 316.2000 826.5000 317.4000 839.7000 ;
	    RECT 318.6000 833.7000 319.8000 839.7000 ;
	    RECT 343.5000 833.7000 344.7000 839.7000 ;
	    RECT 343.8000 830.4000 345.0000 831.6000 ;
	    RECT 343.8000 829.5000 344.7000 830.4000 ;
	    RECT 345.9000 828.6000 347.1000 839.7000 ;
	    RECT 342.6000 828.4500 343.8000 828.6000 ;
	    RECT 321.1500 827.5500 343.8000 828.4500 ;
	    RECT 292.2000 824.4000 293.4000 825.6000 ;
	    RECT 316.2000 825.4500 317.4000 825.6000 ;
	    RECT 321.1500 825.4500 322.0500 827.5500 ;
	    RECT 342.6000 827.4000 343.8000 827.5500 ;
	    RECT 345.6000 827.7000 347.1000 828.6000 ;
	    RECT 349.8000 827.7000 351.0000 839.7000 ;
	    RECT 361.8000 833.7000 363.0000 839.7000 ;
	    RECT 316.2000 824.5500 322.0500 825.4500 ;
	    RECT 316.2000 824.4000 317.4000 824.5500 ;
	    RECT 147.6000 821.7000 148.8000 822.0000 ;
	    RECT 147.6000 820.8000 154.2000 821.7000 ;
	    RECT 155.4000 821.4000 156.6000 822.6000 ;
	    RECT 153.0000 820.5000 154.2000 820.8000 ;
	    RECT 155.4000 820.2000 156.6000 820.5000 ;
	    RECT 133.8000 813.3000 135.0000 819.3000 ;
	    RECT 136.2000 818.1000 139.8000 819.3000 ;
	    RECT 143.4000 818.4000 144.9000 819.6000 ;
	    RECT 149.4000 818.4000 149.7000 819.6000 ;
	    RECT 150.6000 818.4000 151.8000 819.6000 ;
	    RECT 153.0000 819.3000 154.2000 819.6000 ;
	    RECT 158.7000 819.3000 159.9000 822.9000 ;
	    RECT 162.6000 822.3000 175.8000 823.5000 ;
	    RECT 215.4000 823.2000 216.6000 823.5000 ;
	    RECT 220.2000 823.2000 221.4000 823.5000 ;
	    RECT 287.4000 823.2000 288.6000 823.5000 ;
	    RECT 292.2000 823.2000 293.4000 823.5000 ;
	    RECT 167.7000 820.2000 172.2000 821.4000 ;
	    RECT 167.7000 819.3000 168.9000 820.2000 ;
	    RECT 153.0000 818.4000 159.9000 819.3000 ;
	    RECT 138.6000 813.3000 139.8000 818.1000 ;
	    RECT 165.0000 818.1000 168.9000 819.3000 ;
	    RECT 141.0000 813.3000 142.2000 817.5000 ;
	    RECT 143.4000 813.3000 144.6000 817.5000 ;
	    RECT 145.8000 813.3000 147.0000 817.5000 ;
	    RECT 148.2000 813.3000 149.4000 817.5000 ;
	    RECT 150.6000 813.3000 151.8000 816.3000 ;
	    RECT 153.0000 813.3000 154.2000 817.5000 ;
	    RECT 155.4000 813.3000 156.6000 816.3000 ;
	    RECT 157.8000 813.3000 159.0000 817.5000 ;
	    RECT 160.2000 813.3000 161.4000 817.5000 ;
	    RECT 162.6000 813.3000 163.8000 817.5000 ;
	    RECT 165.0000 813.3000 166.2000 818.1000 ;
	    RECT 169.8000 813.3000 171.0000 819.3000 ;
	    RECT 174.6000 813.3000 175.8000 822.3000 ;
	    RECT 213.0000 821.4000 214.2000 822.6000 ;
	    RECT 215.1000 820.8000 215.4000 822.3000 ;
	    RECT 217.8000 821.4000 219.0000 822.6000 ;
	    RECT 222.6000 822.4500 223.8000 822.6000 ;
	    RECT 234.6000 822.4500 235.8000 822.6000 ;
	    RECT 219.9000 821.4000 221.4000 822.3000 ;
	    RECT 222.6000 821.5500 235.8000 822.4500 ;
	    RECT 222.6000 821.4000 223.8000 821.5500 ;
	    RECT 234.6000 821.4000 235.8000 821.5500 ;
	    RECT 253.8000 822.4500 255.0000 822.6000 ;
	    RECT 285.0000 822.4500 286.2000 822.6000 ;
	    RECT 253.8000 821.5500 286.2000 822.4500 ;
	    RECT 253.8000 821.4000 255.0000 821.5500 ;
	    RECT 285.0000 821.4000 286.2000 821.5500 ;
	    RECT 287.4000 821.4000 288.9000 822.3000 ;
	    RECT 289.8000 821.4000 291.0000 822.6000 ;
	    RECT 213.3000 819.3000 218.7000 819.9000 ;
	    RECT 220.5000 819.3000 221.4000 821.4000 ;
	    RECT 213.0000 819.0000 219.0000 819.3000 ;
	    RECT 213.0000 813.3000 214.2000 819.0000 ;
	    RECT 215.4000 813.3000 216.6000 818.1000 ;
	    RECT 217.8000 814.2000 219.0000 819.0000 ;
	    RECT 220.2000 815.1000 221.4000 819.3000 ;
	    RECT 222.6000 814.2000 223.8000 819.3000 ;
	    RECT 217.8000 813.3000 223.8000 814.2000 ;
	    RECT 234.6000 813.3000 235.8000 820.5000 ;
	    RECT 237.0000 819.4500 238.2000 819.6000 ;
	    RECT 239.4000 819.4500 240.6000 819.6000 ;
	    RECT 237.0000 818.5500 240.6000 819.4500 ;
	    RECT 237.0000 818.4000 238.2000 818.5500 ;
	    RECT 239.4000 818.4000 240.6000 818.5500 ;
	    RECT 244.2000 819.4500 245.4000 819.6000 ;
	    RECT 251.4000 819.4500 252.6000 819.6000 ;
	    RECT 244.2000 818.5500 252.6000 819.4500 ;
	    RECT 244.2000 818.4000 245.4000 818.5500 ;
	    RECT 251.4000 818.4000 252.6000 818.5500 ;
	    RECT 237.0000 817.2000 238.2000 817.5000 ;
	    RECT 251.4000 817.2000 252.6000 817.5000 ;
	    RECT 237.0000 813.3000 238.2000 816.3000 ;
	    RECT 251.4000 813.3000 252.6000 816.3000 ;
	    RECT 253.8000 813.3000 255.0000 820.5000 ;
	    RECT 287.4000 819.3000 288.3000 821.4000 ;
	    RECT 293.4000 820.8000 293.7000 822.3000 ;
	    RECT 294.6000 821.4000 295.8000 822.6000 ;
	    RECT 290.1000 819.3000 295.5000 819.9000 ;
	    RECT 316.2000 819.3000 317.4000 823.5000 ;
	    RECT 345.6000 822.6000 346.5000 827.7000 ;
	    RECT 347.4000 824.4000 348.6000 825.6000 ;
	    RECT 364.2000 823.5000 365.4000 839.7000 ;
	    RECT 383.4000 833.7000 384.6000 839.7000 ;
	    RECT 383.4000 829.5000 384.6000 829.8000 ;
	    RECT 366.6000 828.4500 367.8000 828.6000 ;
	    RECT 383.4000 828.4500 384.6000 828.6000 ;
	    RECT 366.6000 827.5500 384.6000 828.4500 ;
	    RECT 366.6000 827.4000 367.8000 827.5500 ;
	    RECT 383.4000 827.4000 384.6000 827.5500 ;
	    RECT 385.8000 826.5000 387.0000 839.7000 ;
	    RECT 388.2000 833.7000 389.4000 839.7000 ;
	    RECT 390.6000 839.4000 391.8000 840.6000 ;
	    RECT 407.4000 833.7000 408.6000 839.7000 ;
	    RECT 407.4000 829.5000 408.6000 829.8000 ;
	    RECT 405.0000 828.4500 406.2000 828.6000 ;
	    RECT 407.4000 828.4500 408.6000 828.6000 ;
	    RECT 405.0000 827.5500 408.6000 828.4500 ;
	    RECT 405.0000 827.4000 406.2000 827.5500 ;
	    RECT 407.4000 827.4000 408.6000 827.5500 ;
	    RECT 409.8000 826.5000 411.0000 839.7000 ;
	    RECT 412.2000 833.7000 413.4000 839.7000 ;
	    RECT 474.6000 827.7000 475.8000 839.7000 ;
	    RECT 477.0000 826.8000 478.2000 839.7000 ;
	    RECT 479.4000 827.7000 480.6000 839.7000 ;
	    RECT 481.8000 826.8000 483.0000 839.7000 ;
	    RECT 484.2000 827.7000 485.4000 839.7000 ;
	    RECT 486.6000 826.8000 487.8000 839.7000 ;
	    RECT 489.0000 827.7000 490.2000 839.7000 ;
	    RECT 491.4000 826.8000 492.6000 839.7000 ;
	    RECT 493.8000 827.7000 495.0000 839.7000 ;
	    RECT 508.2000 833.7000 509.4000 839.7000 ;
	    RECT 477.0000 825.6000 479.7000 826.8000 ;
	    RECT 481.8000 825.6000 485.1000 826.8000 ;
	    RECT 486.6000 825.6000 489.9000 826.8000 ;
	    RECT 491.4000 826.5000 495.0000 826.8000 ;
	    RECT 491.4000 825.6000 492.9000 826.5000 ;
	    RECT 385.8000 825.4500 387.0000 825.6000 ;
	    RECT 402.6000 825.4500 403.8000 825.6000 ;
	    RECT 385.8000 824.5500 403.8000 825.4500 ;
	    RECT 385.8000 824.4000 387.0000 824.5500 ;
	    RECT 402.6000 824.4000 403.8000 824.5500 ;
	    RECT 409.8000 825.4500 411.0000 825.6000 ;
	    RECT 474.6000 825.4500 475.8000 825.6000 ;
	    RECT 409.8000 824.5500 475.8000 825.4500 ;
	    RECT 409.8000 824.4000 411.0000 824.5500 ;
	    RECT 474.6000 824.4000 475.8000 824.5500 ;
	    RECT 478.5000 823.5000 479.7000 825.6000 ;
	    RECT 483.9000 823.5000 485.1000 825.6000 ;
	    RECT 488.7000 823.5000 489.9000 825.6000 ;
	    RECT 493.8000 825.4500 495.0000 825.6000 ;
	    RECT 498.6000 825.4500 499.8000 825.6000 ;
	    RECT 493.8000 824.5500 499.8000 825.4500 ;
	    RECT 493.8000 824.4000 495.0000 824.5500 ;
	    RECT 498.6000 824.4000 499.8000 824.5500 ;
	    RECT 510.6000 823.5000 511.8000 839.7000 ;
	    RECT 522.6000 833.7000 523.8000 839.7000 ;
	    RECT 525.0000 823.5000 526.2000 839.7000 ;
	    RECT 551.4000 827.7000 552.6000 839.7000 ;
	    RECT 555.3000 828.6000 556.5000 839.7000 ;
	    RECT 557.7000 833.7000 558.9000 839.7000 ;
	    RECT 577.8000 833.7000 579.0000 839.7000 ;
	    RECT 557.4000 830.4000 558.6000 831.6000 ;
	    RECT 557.7000 829.5000 558.6000 830.4000 ;
	    RECT 577.8000 829.5000 579.0000 829.8000 ;
	    RECT 555.3000 827.7000 556.8000 828.6000 ;
	    RECT 553.8000 825.4500 555.0000 825.6000 ;
	    RECT 549.1500 824.5500 555.0000 825.4500 ;
	    RECT 347.4000 823.2000 348.6000 823.5000 ;
	    RECT 318.6000 821.4000 319.8000 822.6000 ;
	    RECT 323.4000 822.4500 324.6000 822.6000 ;
	    RECT 340.2000 822.4500 341.4000 822.6000 ;
	    RECT 323.4000 821.5500 341.4000 822.4500 ;
	    RECT 323.4000 821.4000 324.6000 821.5500 ;
	    RECT 340.2000 821.4000 341.4000 821.5500 ;
	    RECT 342.6000 821.4000 343.8000 822.6000 ;
	    RECT 344.7000 821.4000 346.5000 822.6000 ;
	    RECT 348.6000 820.8000 348.9000 822.3000 ;
	    RECT 349.8000 821.4000 351.0000 822.6000 ;
	    RECT 364.2000 822.4500 365.4000 822.6000 ;
	    RECT 381.0000 822.4500 382.2000 822.6000 ;
	    RECT 364.2000 821.5500 382.2000 822.4500 ;
	    RECT 364.2000 821.4000 365.4000 821.5500 ;
	    RECT 381.0000 821.4000 382.2000 821.5500 ;
	    RECT 318.6000 820.2000 319.8000 820.5000 ;
	    RECT 342.9000 819.3000 343.8000 820.5000 ;
	    RECT 345.3000 819.3000 350.7000 819.9000 ;
	    RECT 285.0000 814.2000 286.2000 819.3000 ;
	    RECT 287.4000 815.1000 288.6000 819.3000 ;
	    RECT 289.8000 819.0000 295.8000 819.3000 ;
	    RECT 289.8000 814.2000 291.0000 819.0000 ;
	    RECT 285.0000 813.3000 291.0000 814.2000 ;
	    RECT 292.2000 813.3000 293.4000 818.1000 ;
	    RECT 294.6000 813.3000 295.8000 819.0000 ;
	    RECT 314.7000 818.4000 317.4000 819.3000 ;
	    RECT 314.7000 813.3000 315.9000 818.4000 ;
	    RECT 318.6000 813.3000 319.8000 819.3000 ;
	    RECT 342.6000 813.3000 343.8000 819.3000 ;
	    RECT 345.0000 819.0000 351.0000 819.3000 ;
	    RECT 345.0000 813.3000 346.2000 819.0000 ;
	    RECT 347.4000 813.3000 348.6000 818.1000 ;
	    RECT 349.8000 813.3000 351.0000 819.0000 ;
	    RECT 361.8000 818.4000 363.0000 819.6000 ;
	    RECT 361.8000 817.2000 363.0000 817.5000 ;
	    RECT 361.8000 813.3000 363.0000 816.3000 ;
	    RECT 364.2000 813.3000 365.4000 820.5000 ;
	    RECT 385.8000 819.3000 387.0000 823.5000 ;
	    RECT 388.2000 822.4500 389.4000 822.6000 ;
	    RECT 390.6000 822.4500 391.8000 822.6000 ;
	    RECT 388.2000 821.5500 391.8000 822.4500 ;
	    RECT 388.2000 821.4000 389.4000 821.5500 ;
	    RECT 390.6000 821.4000 391.8000 821.5500 ;
	    RECT 388.2000 820.2000 389.4000 820.5000 ;
	    RECT 409.8000 819.3000 411.0000 823.5000 ;
	    RECT 412.2000 821.4000 413.4000 822.6000 ;
	    RECT 431.4000 822.4500 432.6000 822.6000 ;
	    RECT 474.6000 822.4500 475.8000 822.6000 ;
	    RECT 431.4000 821.5500 475.8000 822.4500 ;
	    RECT 476.7000 822.3000 477.3000 823.5000 ;
	    RECT 478.5000 822.3000 482.4000 823.5000 ;
	    RECT 483.9000 822.3000 487.5000 823.5000 ;
	    RECT 488.7000 822.3000 492.6000 823.5000 ;
	    RECT 431.4000 821.4000 432.6000 821.5500 ;
	    RECT 474.6000 821.4000 475.8000 821.5500 ;
	    RECT 478.5000 821.4000 479.7000 822.3000 ;
	    RECT 483.9000 821.4000 485.1000 822.3000 ;
	    RECT 488.7000 821.4000 489.9000 822.3000 ;
	    RECT 493.8000 821.4000 495.0000 823.5000 ;
	    RECT 496.2000 822.4500 497.4000 822.6000 ;
	    RECT 510.6000 822.4500 511.8000 822.6000 ;
	    RECT 496.2000 821.5500 511.8000 822.4500 ;
	    RECT 496.2000 821.4000 497.4000 821.5500 ;
	    RECT 510.6000 821.4000 511.8000 821.5500 ;
	    RECT 525.0000 822.4500 526.2000 822.6000 ;
	    RECT 549.1500 822.4500 550.0500 824.5500 ;
	    RECT 553.8000 824.4000 555.0000 824.5500 ;
	    RECT 553.8000 823.2000 555.0000 823.5000 ;
	    RECT 555.9000 822.6000 556.8000 827.7000 ;
	    RECT 558.6000 827.4000 559.8000 828.6000 ;
	    RECT 577.8000 827.4000 579.0000 828.6000 ;
	    RECT 558.7500 825.4500 559.6500 827.4000 ;
	    RECT 580.2000 826.5000 581.4000 839.7000 ;
	    RECT 582.6000 833.7000 583.8000 839.7000 ;
	    RECT 601.8000 833.7000 603.0000 839.7000 ;
	    RECT 604.2000 826.5000 605.4000 839.7000 ;
	    RECT 606.6000 833.7000 607.8000 839.7000 ;
	    RECT 631.5000 833.7000 632.7000 839.7000 ;
	    RECT 631.8000 830.4000 633.0000 831.6000 ;
	    RECT 606.6000 829.5000 607.8000 829.8000 ;
	    RECT 631.8000 829.5000 632.7000 830.4000 ;
	    RECT 633.9000 828.6000 635.1000 839.7000 ;
	    RECT 606.6000 827.4000 607.8000 828.6000 ;
	    RECT 618.6000 828.4500 619.8000 828.6000 ;
	    RECT 628.2000 828.4500 629.4000 828.6000 ;
	    RECT 630.6000 828.4500 631.8000 828.6000 ;
	    RECT 618.6000 827.5500 631.8000 828.4500 ;
	    RECT 618.6000 827.4000 619.8000 827.5500 ;
	    RECT 628.2000 827.4000 629.4000 827.5500 ;
	    RECT 630.6000 827.4000 631.8000 827.5500 ;
	    RECT 633.6000 827.7000 635.1000 828.6000 ;
	    RECT 637.8000 827.7000 639.0000 839.7000 ;
	    RECT 685.8000 828.6000 687.0000 839.7000 ;
	    RECT 688.2000 829.8000 689.7000 839.7000 ;
	    RECT 688.5000 828.6000 689.7000 828.9000 ;
	    RECT 685.8000 827.7000 689.7000 828.6000 ;
	    RECT 692.4000 827.7000 694.8000 839.7000 ;
	    RECT 697.5000 829.8000 699.0000 839.7000 ;
	    RECT 697.8000 828.6000 699.0000 828.9000 ;
	    RECT 700.2000 828.6000 701.4000 839.7000 ;
	    RECT 697.8000 827.7000 701.4000 828.6000 ;
	    RECT 731.4000 838.8000 737.4000 839.7000 ;
	    RECT 731.4000 827.7000 732.6000 838.8000 ;
	    RECT 733.8000 827.7000 735.0000 837.9000 ;
	    RECT 736.2000 828.6000 737.4000 838.8000 ;
	    RECT 738.6000 829.5000 739.8000 839.7000 ;
	    RECT 741.0000 828.6000 742.2000 839.7000 ;
	    RECT 760.2000 833.7000 761.4000 839.7000 ;
	    RECT 760.2000 829.5000 761.4000 829.8000 ;
	    RECT 736.2000 827.7000 742.2000 828.6000 ;
	    RECT 580.2000 825.4500 581.4000 825.6000 ;
	    RECT 558.7500 824.5500 581.4000 825.4500 ;
	    RECT 580.2000 824.4000 581.4000 824.5500 ;
	    RECT 582.6000 825.4500 583.8000 825.6000 ;
	    RECT 604.2000 825.4500 605.4000 825.6000 ;
	    RECT 582.6000 824.5500 605.4000 825.4500 ;
	    RECT 582.6000 824.4000 583.8000 824.5500 ;
	    RECT 604.2000 824.4000 605.4000 824.5500 ;
	    RECT 525.0000 821.5500 550.0500 822.4500 ;
	    RECT 525.0000 821.4000 526.2000 821.5500 ;
	    RECT 551.4000 821.4000 552.6000 822.6000 ;
	    RECT 412.2000 820.2000 413.4000 820.5000 ;
	    RECT 477.0000 820.2000 479.7000 821.4000 ;
	    RECT 481.8000 820.2000 485.1000 821.4000 ;
	    RECT 486.6000 820.2000 489.9000 821.4000 ;
	    RECT 491.4000 820.2000 495.0000 821.4000 ;
	    RECT 553.5000 820.8000 553.8000 822.3000 ;
	    RECT 555.9000 821.4000 557.7000 822.6000 ;
	    RECT 558.6000 822.4500 559.8000 822.6000 ;
	    RECT 570.6000 822.4500 571.8000 822.6000 ;
	    RECT 558.6000 821.5500 571.8000 822.4500 ;
	    RECT 558.6000 821.4000 559.8000 821.5500 ;
	    RECT 570.6000 821.4000 571.8000 821.5500 ;
	    RECT 384.3000 818.4000 387.0000 819.3000 ;
	    RECT 384.3000 813.3000 385.5000 818.4000 ;
	    RECT 388.2000 813.3000 389.4000 819.3000 ;
	    RECT 408.3000 818.4000 411.0000 819.3000 ;
	    RECT 408.3000 813.3000 409.5000 818.4000 ;
	    RECT 412.2000 813.3000 413.4000 819.3000 ;
	    RECT 474.6000 813.3000 475.8000 819.3000 ;
	    RECT 477.0000 813.3000 478.2000 820.2000 ;
	    RECT 479.4000 813.3000 480.6000 819.3000 ;
	    RECT 481.8000 813.3000 483.0000 820.2000 ;
	    RECT 484.2000 813.3000 485.4000 819.3000 ;
	    RECT 486.6000 813.3000 487.8000 820.2000 ;
	    RECT 489.0000 813.3000 490.2000 819.3000 ;
	    RECT 491.4000 813.3000 492.6000 820.2000 ;
	    RECT 493.8000 813.3000 495.0000 819.3000 ;
	    RECT 508.2000 818.4000 509.4000 819.6000 ;
	    RECT 508.2000 817.2000 509.4000 817.5000 ;
	    RECT 508.2000 813.3000 509.4000 816.3000 ;
	    RECT 510.6000 813.3000 511.8000 820.5000 ;
	    RECT 522.6000 818.4000 523.8000 819.6000 ;
	    RECT 522.6000 817.2000 523.8000 817.5000 ;
	    RECT 522.6000 813.3000 523.8000 816.3000 ;
	    RECT 525.0000 813.3000 526.2000 820.5000 ;
	    RECT 551.7000 819.3000 557.1000 819.9000 ;
	    RECT 558.6000 819.3000 559.5000 820.5000 ;
	    RECT 580.2000 819.3000 581.4000 823.5000 ;
	    RECT 582.6000 822.4500 583.8000 822.6000 ;
	    RECT 599.4000 822.4500 600.6000 822.6000 ;
	    RECT 601.8000 822.4500 603.0000 822.6000 ;
	    RECT 582.6000 821.5500 603.0000 822.4500 ;
	    RECT 582.6000 821.4000 583.8000 821.5500 ;
	    RECT 599.4000 821.4000 600.6000 821.5500 ;
	    RECT 601.8000 821.4000 603.0000 821.5500 ;
	    RECT 582.6000 820.2000 583.8000 820.5000 ;
	    RECT 601.8000 820.2000 603.0000 820.5000 ;
	    RECT 604.2000 819.3000 605.4000 823.5000 ;
	    RECT 633.6000 822.6000 634.5000 827.7000 ;
	    RECT 693.3000 826.5000 694.2000 827.7000 ;
	    RECT 734.1000 826.8000 735.0000 827.7000 ;
	    RECT 760.2000 827.4000 761.4000 828.6000 ;
	    RECT 731.4000 826.5000 732.6000 826.8000 ;
	    RECT 734.1000 826.5000 737.1000 826.8000 ;
	    RECT 762.6000 826.5000 763.8000 839.7000 ;
	    RECT 765.0000 833.7000 766.2000 839.7000 ;
	    RECT 785.1000 828.9000 786.3000 839.7000 ;
	    RECT 785.1000 827.7000 787.8000 828.9000 ;
	    RECT 789.0000 827.7000 790.2000 839.7000 ;
	    RECT 817.8000 827.7000 819.0000 839.7000 ;
	    RECT 821.7000 827.7000 824.7000 839.7000 ;
	    RECT 827.4000 827.7000 828.6000 839.7000 ;
	    RECT 784.2000 826.5000 785.4000 826.8000 ;
	    RECT 734.1000 825.9000 735.3000 826.5000 ;
	    RECT 690.3000 825.6000 691.5000 825.9000 ;
	    RECT 635.4000 825.4500 636.6000 825.6000 ;
	    RECT 673.8000 825.4500 675.0000 825.6000 ;
	    RECT 635.4000 824.5500 675.0000 825.4500 ;
	    RECT 635.4000 824.4000 636.6000 824.5500 ;
	    RECT 673.8000 824.4000 675.0000 824.5500 ;
	    RECT 689.1000 824.7000 691.5000 825.6000 ;
	    RECT 693.0000 825.4500 694.2000 825.6000 ;
	    RECT 705.0000 825.4500 706.2000 825.6000 ;
	    RECT 689.1000 824.4000 690.3000 824.7000 ;
	    RECT 693.0000 824.5500 706.2000 825.4500 ;
	    RECT 693.0000 824.4000 694.2000 824.5500 ;
	    RECT 705.0000 824.4000 706.2000 824.5500 ;
	    RECT 726.6000 825.4500 727.8000 825.6000 ;
	    RECT 731.4000 825.4500 732.6000 825.6000 ;
	    RECT 726.6000 824.5500 732.6000 825.4500 ;
	    RECT 726.6000 824.4000 727.8000 824.5500 ;
	    RECT 731.4000 824.4000 732.6000 824.5500 ;
	    RECT 736.2000 824.4000 737.4000 825.6000 ;
	    RECT 739.8000 824.7000 740.1000 826.2000 ;
	    RECT 741.0000 824.4000 742.2000 825.6000 ;
	    RECT 762.6000 825.4500 763.8000 825.6000 ;
	    RECT 781.8000 825.4500 783.0000 825.6000 ;
	    RECT 762.6000 824.5500 783.0000 825.4500 ;
	    RECT 762.6000 824.4000 763.8000 824.5500 ;
	    RECT 781.8000 824.4000 783.0000 824.5500 ;
	    RECT 784.2000 824.4000 785.4000 825.6000 ;
	    RECT 734.1000 823.5000 735.3000 824.4000 ;
	    RECT 738.6000 823.5000 739.8000 823.8000 ;
	    RECT 786.6000 823.5000 787.5000 827.7000 ;
	    RECT 820.2000 824.4000 821.4000 825.6000 ;
	    RECT 817.8000 823.5000 819.0000 823.8000 ;
	    RECT 822.9000 823.5000 823.8000 827.7000 ;
	    RECT 825.0000 824.4000 826.2000 825.6000 ;
	    RECT 841.8000 823.5000 843.0000 839.7000 ;
	    RECT 844.2000 833.7000 845.4000 839.7000 ;
	    RECT 858.6000 823.5000 859.8000 839.7000 ;
	    RECT 861.0000 833.7000 862.2000 839.7000 ;
	    RECT 880.2000 833.7000 881.4000 839.7000 ;
	    RECT 880.2000 829.5000 881.4000 829.8000 ;
	    RECT 875.4000 828.4500 876.6000 828.6000 ;
	    RECT 880.2000 828.4500 881.4000 828.6000 ;
	    RECT 875.4000 827.5500 881.4000 828.4500 ;
	    RECT 875.4000 827.4000 876.6000 827.5500 ;
	    RECT 880.2000 827.4000 881.4000 827.5500 ;
	    RECT 882.6000 826.5000 883.8000 839.7000 ;
	    RECT 885.0000 833.7000 886.2000 839.7000 ;
	    RECT 904.2000 833.7000 905.4000 839.7000 ;
	    RECT 868.2000 825.4500 869.4000 825.6000 ;
	    RECT 882.6000 825.4500 883.8000 825.6000 ;
	    RECT 868.2000 824.5500 883.8000 825.4500 ;
	    RECT 868.2000 824.4000 869.4000 824.5500 ;
	    RECT 882.6000 824.4000 883.8000 824.5500 ;
	    RECT 906.6000 823.5000 907.8000 839.7000 ;
	    RECT 926.7000 828.9000 927.9000 839.7000 ;
	    RECT 926.7000 827.7000 929.4000 828.9000 ;
	    RECT 930.6000 827.7000 931.8000 839.7000 ;
	    RECT 959.4000 827.7000 960.6000 839.7000 ;
	    RECT 963.3000 827.7000 966.3000 839.7000 ;
	    RECT 969.0000 827.7000 970.2000 839.7000 ;
	    RECT 973.8000 837.4500 975.0000 837.6000 ;
	    RECT 981.0000 837.4500 982.2000 837.6000 ;
	    RECT 973.8000 836.5500 982.2000 837.4500 ;
	    RECT 973.8000 836.4000 975.0000 836.5500 ;
	    RECT 981.0000 836.4000 982.2000 836.5500 ;
	    RECT 925.8000 826.5000 927.0000 826.8000 ;
	    RECT 921.0000 825.4500 922.2000 825.6000 ;
	    RECT 925.8000 825.4500 927.0000 825.6000 ;
	    RECT 921.0000 824.5500 927.0000 825.4500 ;
	    RECT 921.0000 824.4000 922.2000 824.5500 ;
	    RECT 925.8000 824.4000 927.0000 824.5500 ;
	    RECT 928.2000 823.5000 929.1000 827.7000 ;
	    RECT 961.8000 824.4000 963.0000 825.6000 ;
	    RECT 964.2000 823.5000 965.1000 827.7000 ;
	    RECT 966.6000 824.4000 967.8000 825.6000 ;
	    RECT 969.0000 823.5000 970.2000 823.8000 ;
	    RECT 983.4000 823.5000 984.6000 839.7000 ;
	    RECT 985.8000 833.7000 987.0000 839.7000 ;
	    RECT 1000.2000 823.5000 1001.4000 839.7000 ;
	    RECT 1002.6000 833.7000 1003.8000 839.7000 ;
	    RECT 1137.0000 833.7000 1138.2001 839.7000 ;
	    RECT 1139.4000 832.5000 1140.6000 839.7000 ;
	    RECT 1141.8000 833.7000 1143.0000 839.7000 ;
	    RECT 1144.2001 832.8000 1145.4000 839.7000 ;
	    RECT 1146.6000 833.7000 1147.8000 839.7000 ;
	    RECT 1141.5000 831.9000 1145.4000 832.8000 ;
	    RECT 1139.4000 830.4000 1140.6000 831.6000 ;
	    RECT 1141.5000 829.5000 1142.4000 831.9000 ;
	    RECT 1149.0000 831.6000 1150.2001 839.7000 ;
	    RECT 1151.4000 833.7000 1152.6000 839.7000 ;
	    RECT 1153.8000 835.5000 1155.0000 839.7000 ;
	    RECT 1156.2001 835.5000 1157.4000 839.7000 ;
	    RECT 1158.6000 835.5000 1159.8000 839.7000 ;
	    RECT 1151.1000 831.6000 1157.4000 832.8000 ;
	    RECT 1146.3000 830.4000 1150.2001 831.6000 ;
	    RECT 1161.0000 830.4000 1162.2001 839.7000 ;
	    RECT 1163.4000 833.7000 1164.6000 839.7000 ;
	    RECT 1165.8000 832.5000 1167.0000 839.7000 ;
	    RECT 1168.2001 833.7000 1169.4000 839.7000 ;
	    RECT 1170.6000 832.5000 1171.8000 839.7000 ;
	    RECT 1173.0000 835.5000 1174.2001 839.7000 ;
	    RECT 1175.4000 835.5000 1176.6000 839.7000 ;
	    RECT 1177.8000 833.7000 1179.0000 839.7000 ;
	    RECT 1180.2001 832.8000 1181.4000 839.7000 ;
	    RECT 1182.6000 833.7000 1183.8000 840.6000 ;
	    RECT 1185.0000 834.6000 1186.2001 839.7000 ;
	    RECT 1185.0000 833.7000 1186.5000 834.6000 ;
	    RECT 1187.4000 833.7000 1188.6000 839.7000 ;
	    RECT 1212.3000 833.7000 1213.5000 839.7000 ;
	    RECT 1185.6000 832.8000 1186.5000 833.7000 ;
	    RECT 1178.4000 831.6000 1184.7001 832.8000 ;
	    RECT 1185.6000 831.9000 1188.6000 832.8000 ;
	    RECT 1165.8000 830.4000 1169.7001 831.6000 ;
	    RECT 1170.6000 830.7000 1179.3000 831.6000 ;
	    RECT 1183.8000 831.0000 1184.7001 831.6000 ;
	    RECT 1153.8000 829.5000 1155.0000 829.8000 ;
	    RECT 1139.4000 828.0000 1140.6000 829.5000 ;
	    RECT 1139.1000 826.8000 1140.6000 828.0000 ;
	    RECT 1141.5000 828.6000 1155.0000 829.5000 ;
	    RECT 1158.6000 829.5000 1159.8000 829.8000 ;
	    RECT 1170.6000 829.5000 1171.5000 830.7000 ;
	    RECT 1180.2001 829.8000 1182.3000 830.7000 ;
	    RECT 1183.8000 829.8000 1186.2001 831.0000 ;
	    RECT 1158.6000 828.6000 1171.5000 829.5000 ;
	    RECT 1173.0000 829.5000 1182.3000 829.8000 ;
	    RECT 1173.0000 828.9000 1181.1000 829.5000 ;
	    RECT 1173.0000 828.6000 1174.2001 828.9000 ;
	    RECT 635.4000 823.2000 636.6000 823.5000 ;
	    RECT 691.2000 822.9000 692.4000 823.2000 ;
	    RECT 688.2000 822.6000 692.4000 822.9000 ;
	    RECT 630.6000 821.4000 631.8000 822.6000 ;
	    RECT 632.7000 821.4000 634.5000 822.6000 ;
	    RECT 637.8000 822.4500 639.0000 822.6000 ;
	    RECT 642.6000 822.4500 643.8000 822.6000 ;
	    RECT 636.6000 820.8000 636.9000 822.3000 ;
	    RECT 637.8000 821.5500 643.8000 822.4500 ;
	    RECT 637.8000 821.4000 639.0000 821.5500 ;
	    RECT 642.6000 821.4000 643.8000 821.5500 ;
	    RECT 685.8000 821.4000 687.0000 822.6000 ;
	    RECT 687.9000 822.0000 692.4000 822.6000 ;
	    RECT 693.3000 822.6000 694.2000 823.5000 ;
	    RECT 687.9000 821.7000 689.1000 822.0000 ;
	    RECT 693.3000 821.7000 694.8000 822.6000 ;
	    RECT 687.9000 821.4000 688.2000 821.7000 ;
	    RECT 630.9000 819.3000 631.8000 820.5000 ;
	    RECT 688.5000 820.2000 689.7000 820.5000 ;
	    RECT 633.3000 819.3000 638.7000 819.9000 ;
	    RECT 685.8000 819.3000 689.7000 820.2000 ;
	    RECT 690.6000 819.6000 693.0000 820.8000 ;
	    RECT 551.4000 819.0000 557.4000 819.3000 ;
	    RECT 551.4000 813.3000 552.6000 819.0000 ;
	    RECT 553.8000 813.3000 555.0000 818.1000 ;
	    RECT 556.2000 813.3000 557.4000 819.0000 ;
	    RECT 558.6000 813.3000 559.8000 819.3000 ;
	    RECT 578.7000 818.4000 581.4000 819.3000 ;
	    RECT 578.7000 813.3000 579.9000 818.4000 ;
	    RECT 582.6000 813.3000 583.8000 819.3000 ;
	    RECT 601.8000 813.3000 603.0000 819.3000 ;
	    RECT 604.2000 818.4000 606.9000 819.3000 ;
	    RECT 605.7000 813.3000 606.9000 818.4000 ;
	    RECT 630.6000 813.3000 631.8000 819.3000 ;
	    RECT 633.0000 819.0000 639.0000 819.3000 ;
	    RECT 633.0000 813.3000 634.2000 819.0000 ;
	    RECT 635.4000 813.3000 636.6000 818.1000 ;
	    RECT 637.8000 813.3000 639.0000 819.0000 ;
	    RECT 685.8000 813.3000 687.0000 819.3000 ;
	    RECT 693.9000 818.7000 694.8000 821.7000 ;
	    RECT 696.0000 821.4000 697.2000 822.6000 ;
	    RECT 699.0000 821.4000 699.3000 822.6000 ;
	    RECT 700.2000 821.4000 701.4000 822.6000 ;
	    RECT 707.4000 822.4500 708.6000 822.6000 ;
	    RECT 733.8000 822.4500 735.0000 822.6000 ;
	    RECT 707.4000 821.5500 735.0000 822.4500 ;
	    RECT 707.4000 821.4000 708.6000 821.5500 ;
	    RECT 733.8000 821.4000 735.0000 821.5500 ;
	    RECT 696.0000 820.8000 696.9000 821.4000 ;
	    RECT 695.7000 819.6000 696.9000 820.8000 ;
	    RECT 697.8000 820.2000 699.0000 820.5000 ;
	    RECT 697.8000 819.3000 701.4000 820.2000 ;
	    RECT 736.2000 819.3000 737.1000 823.5000 ;
	    RECT 738.6000 822.4500 739.8000 822.6000 ;
	    RECT 741.0000 822.4500 742.2000 822.6000 ;
	    RECT 738.6000 821.5500 742.2000 822.4500 ;
	    RECT 738.6000 821.4000 739.8000 821.5500 ;
	    RECT 741.0000 821.4000 742.2000 821.5500 ;
	    RECT 762.6000 819.3000 763.8000 823.5000 ;
	    RECT 820.2000 823.2000 821.4000 823.5000 ;
	    RECT 825.0000 823.2000 826.2000 823.5000 ;
	    RECT 765.0000 821.4000 766.2000 822.6000 ;
	    RECT 786.6000 822.4500 787.8000 822.6000 ;
	    RECT 815.4000 822.4500 816.6000 822.6000 ;
	    RECT 786.6000 821.5500 816.6000 822.4500 ;
	    RECT 786.6000 821.4000 787.8000 821.5500 ;
	    RECT 815.4000 821.4000 816.6000 821.5500 ;
	    RECT 817.8000 821.4000 819.0000 822.6000 ;
	    RECT 820.2000 821.4000 821.7000 822.3000 ;
	    RECT 822.6000 821.4000 823.8000 822.6000 ;
	    RECT 765.0000 820.2000 766.2000 820.5000 ;
	    RECT 688.2000 813.3000 689.7000 818.4000 ;
	    RECT 692.4000 813.3000 694.8000 818.7000 ;
	    RECT 697.5000 813.3000 699.0000 818.4000 ;
	    RECT 700.2000 813.3000 701.4000 819.3000 ;
	    RECT 731.4000 813.3000 732.6000 819.3000 ;
	    RECT 735.3000 813.3000 737.7000 819.3000 ;
	    RECT 740.4000 813.3000 741.6000 819.3000 ;
	    RECT 761.1000 818.4000 763.8000 819.3000 ;
	    RECT 761.1000 813.3000 762.3000 818.4000 ;
	    RECT 765.0000 813.3000 766.2000 819.3000 ;
	    RECT 786.6000 816.3000 787.5000 820.5000 ;
	    RECT 789.0000 818.4000 790.2000 819.6000 ;
	    RECT 820.2000 819.3000 821.1000 821.4000 ;
	    RECT 826.2000 820.8000 826.5000 822.3000 ;
	    RECT 827.4000 821.4000 828.6000 822.6000 ;
	    RECT 829.8000 822.4500 831.0000 822.6000 ;
	    RECT 841.8000 822.4500 843.0000 822.6000 ;
	    RECT 829.8000 821.5500 843.0000 822.4500 ;
	    RECT 829.8000 821.4000 831.0000 821.5500 ;
	    RECT 841.8000 821.4000 843.0000 821.5500 ;
	    RECT 844.2000 822.4500 845.4000 822.6000 ;
	    RECT 858.6000 822.4500 859.8000 822.6000 ;
	    RECT 844.2000 821.5500 859.8000 822.4500 ;
	    RECT 844.2000 821.4000 845.4000 821.5500 ;
	    RECT 858.6000 821.4000 859.8000 821.5500 ;
	    RECT 822.9000 819.3000 828.3000 819.9000 ;
	    RECT 789.0000 817.2000 790.2000 817.5000 ;
	    RECT 784.2000 813.3000 785.4000 816.3000 ;
	    RECT 786.6000 813.3000 787.8000 816.3000 ;
	    RECT 789.0000 813.3000 790.2000 816.3000 ;
	    RECT 817.8000 814.2000 819.0000 819.3000 ;
	    RECT 820.2000 815.1000 821.4000 819.3000 ;
	    RECT 822.6000 819.0000 828.6000 819.3000 ;
	    RECT 822.6000 814.2000 823.8000 819.0000 ;
	    RECT 817.8000 813.3000 823.8000 814.2000 ;
	    RECT 825.0000 813.3000 826.2000 818.1000 ;
	    RECT 827.4000 813.3000 828.6000 819.0000 ;
	    RECT 841.8000 813.3000 843.0000 820.5000 ;
	    RECT 844.2000 819.4500 845.4000 819.6000 ;
	    RECT 846.6000 819.4500 847.8000 819.6000 ;
	    RECT 844.2000 818.5500 847.8000 819.4500 ;
	    RECT 844.2000 818.4000 845.4000 818.5500 ;
	    RECT 846.6000 818.4000 847.8000 818.5500 ;
	    RECT 844.2000 817.2000 845.4000 817.5000 ;
	    RECT 844.2000 813.3000 845.4000 816.3000 ;
	    RECT 858.6000 813.3000 859.8000 820.5000 ;
	    RECT 861.0000 819.4500 862.2000 819.6000 ;
	    RECT 863.4000 819.4500 864.6000 819.6000 ;
	    RECT 861.0000 818.5500 864.6000 819.4500 ;
	    RECT 882.6000 819.3000 883.8000 823.5000 ;
	    RECT 961.8000 823.2000 963.0000 823.5000 ;
	    RECT 966.6000 823.2000 967.8000 823.5000 ;
	    RECT 885.0000 822.4500 886.2000 822.6000 ;
	    RECT 887.4000 822.4500 888.6000 822.6000 ;
	    RECT 885.0000 821.5500 888.6000 822.4500 ;
	    RECT 885.0000 821.4000 886.2000 821.5500 ;
	    RECT 887.4000 821.4000 888.6000 821.5500 ;
	    RECT 906.6000 822.4500 907.8000 822.6000 ;
	    RECT 913.8000 822.4500 915.0000 822.6000 ;
	    RECT 906.6000 821.5500 915.0000 822.4500 ;
	    RECT 906.6000 821.4000 907.8000 821.5500 ;
	    RECT 913.8000 821.4000 915.0000 821.5500 ;
	    RECT 918.6000 822.4500 919.8000 822.6000 ;
	    RECT 928.2000 822.4500 929.4000 822.6000 ;
	    RECT 918.6000 821.5500 929.4000 822.4500 ;
	    RECT 918.6000 821.4000 919.8000 821.5500 ;
	    RECT 928.2000 821.4000 929.4000 821.5500 ;
	    RECT 945.0000 822.4500 946.2000 822.6000 ;
	    RECT 959.4000 822.4500 960.6000 822.6000 ;
	    RECT 945.0000 821.5500 960.6000 822.4500 ;
	    RECT 945.0000 821.4000 946.2000 821.5500 ;
	    RECT 959.4000 821.4000 960.6000 821.5500 ;
	    RECT 961.5000 820.8000 961.8000 822.3000 ;
	    RECT 964.2000 821.4000 965.4000 822.6000 ;
	    RECT 969.0000 822.4500 970.2000 822.6000 ;
	    RECT 973.8000 822.4500 975.0000 822.6000 ;
	    RECT 966.3000 821.4000 967.8000 822.3000 ;
	    RECT 969.0000 821.5500 975.0000 822.4500 ;
	    RECT 969.0000 821.4000 970.2000 821.5500 ;
	    RECT 973.8000 821.4000 975.0000 821.5500 ;
	    RECT 983.4000 821.4000 984.6000 822.6000 ;
	    RECT 985.8000 822.4500 987.0000 822.6000 ;
	    RECT 1000.2000 822.4500 1001.4000 822.6000 ;
	    RECT 985.8000 821.5500 1001.4000 822.4500 ;
	    RECT 985.8000 821.4000 987.0000 821.5500 ;
	    RECT 1000.2000 821.4000 1001.4000 821.5500 ;
	    RECT 885.0000 820.2000 886.2000 820.5000 ;
	    RECT 887.4000 819.4500 888.6000 819.6000 ;
	    RECT 904.2000 819.4500 905.4000 819.6000 ;
	    RECT 861.0000 818.4000 862.2000 818.5500 ;
	    RECT 863.4000 818.4000 864.6000 818.5500 ;
	    RECT 881.1000 818.4000 883.8000 819.3000 ;
	    RECT 861.0000 817.2000 862.2000 817.5000 ;
	    RECT 861.0000 813.3000 862.2000 816.3000 ;
	    RECT 881.1000 813.3000 882.3000 818.4000 ;
	    RECT 885.0000 813.3000 886.2000 819.3000 ;
	    RECT 887.4000 818.5500 905.4000 819.4500 ;
	    RECT 887.4000 818.4000 888.6000 818.5500 ;
	    RECT 904.2000 818.4000 905.4000 818.5500 ;
	    RECT 904.2000 817.2000 905.4000 817.5000 ;
	    RECT 904.2000 813.3000 905.4000 816.3000 ;
	    RECT 906.6000 813.3000 907.8000 820.5000 ;
	    RECT 928.2000 816.3000 929.1000 820.5000 ;
	    RECT 930.6000 819.4500 931.8000 819.6000 ;
	    RECT 942.6000 819.4500 943.8000 819.6000 ;
	    RECT 930.6000 818.5500 943.8000 819.4500 ;
	    RECT 959.7000 819.3000 965.1000 819.9000 ;
	    RECT 966.9000 819.3000 967.8000 821.4000 ;
	    RECT 930.6000 818.4000 931.8000 818.5500 ;
	    RECT 942.6000 818.4000 943.8000 818.5500 ;
	    RECT 959.4000 819.0000 965.4000 819.3000 ;
	    RECT 930.6000 817.2000 931.8000 817.5000 ;
	    RECT 925.8000 813.3000 927.0000 816.3000 ;
	    RECT 928.2000 813.3000 929.4000 816.3000 ;
	    RECT 930.6000 813.3000 931.8000 816.3000 ;
	    RECT 959.4000 813.3000 960.6000 819.0000 ;
	    RECT 961.8000 813.3000 963.0000 818.1000 ;
	    RECT 964.2000 814.2000 965.4000 819.0000 ;
	    RECT 966.6000 815.1000 967.8000 819.3000 ;
	    RECT 969.0000 814.2000 970.2000 819.3000 ;
	    RECT 964.2000 813.3000 970.2000 814.2000 ;
	    RECT 983.4000 813.3000 984.6000 820.5000 ;
	    RECT 985.8000 819.4500 987.0000 819.6000 ;
	    RECT 988.2000 819.4500 989.4000 819.6000 ;
	    RECT 985.8000 818.5500 989.4000 819.4500 ;
	    RECT 985.8000 818.4000 987.0000 818.5500 ;
	    RECT 988.2000 818.4000 989.4000 818.5500 ;
	    RECT 985.8000 817.2000 987.0000 817.5000 ;
	    RECT 985.8000 813.3000 987.0000 816.3000 ;
	    RECT 1000.2000 813.3000 1001.4000 820.5000 ;
	    RECT 1139.1000 820.2000 1140.3000 826.8000 ;
	    RECT 1141.5000 825.9000 1142.4000 828.6000 ;
	    RECT 1177.5000 827.7000 1178.7001 828.0000 ;
	    RECT 1143.3000 826.8000 1181.7001 827.7000 ;
	    RECT 1182.6000 827.4000 1183.8000 828.6000 ;
	    RECT 1143.3000 826.5000 1144.5000 826.8000 ;
	    RECT 1141.2001 825.0000 1142.4000 825.9000 ;
	    RECT 1151.4000 825.0000 1176.9000 825.9000 ;
	    RECT 1141.2001 822.0000 1142.1000 825.0000 ;
	    RECT 1151.4000 824.1000 1152.6000 825.0000 ;
	    RECT 1177.8000 824.4000 1179.0000 825.6000 ;
	    RECT 1179.9000 825.0000 1186.5000 825.9000 ;
	    RECT 1185.3000 824.7000 1186.5000 825.0000 ;
	    RECT 1143.0000 822.9000 1148.7001 824.1000 ;
	    RECT 1141.2001 821.1000 1143.0000 822.0000 ;
	    RECT 1002.6000 819.4500 1003.8000 819.6000 ;
	    RECT 1117.8000 819.4500 1119.0000 819.6000 ;
	    RECT 1002.6000 818.5500 1119.0000 819.4500 ;
	    RECT 1139.1000 819.0000 1140.6000 820.2000 ;
	    RECT 1002.6000 818.4000 1003.8000 818.5500 ;
	    RECT 1117.8000 818.4000 1119.0000 818.5500 ;
	    RECT 1002.6000 817.2000 1003.8000 817.5000 ;
	    RECT 1002.6000 813.3000 1003.8000 816.3000 ;
	    RECT 1137.0000 813.3000 1138.2001 816.3000 ;
	    RECT 1139.4000 813.3000 1140.6000 819.0000 ;
	    RECT 1141.8000 813.3000 1143.0000 821.1000 ;
	    RECT 1147.5000 821.1000 1148.7001 822.9000 ;
	    RECT 1147.5000 820.2000 1150.2001 821.1000 ;
	    RECT 1149.0000 819.3000 1150.2001 820.2000 ;
	    RECT 1156.2001 819.6000 1157.4000 823.8000 ;
	    RECT 1161.0000 822.9000 1165.8000 824.1000 ;
	    RECT 1171.5000 822.9000 1174.5000 824.1000 ;
	    RECT 1187.4000 823.5000 1188.6000 831.9000 ;
	    RECT 1212.6000 830.4000 1213.8000 831.6000 ;
	    RECT 1212.6000 829.5000 1213.5000 830.4000 ;
	    RECT 1214.7001 828.6000 1215.9000 839.7000 ;
	    RECT 1211.4000 827.4000 1212.6000 828.6000 ;
	    RECT 1214.4000 827.7000 1215.9000 828.6000 ;
	    RECT 1218.6000 827.7000 1219.8000 839.7000 ;
	    RECT 1160.4000 821.7000 1161.6000 822.0000 ;
	    RECT 1160.4000 820.8000 1167.0000 821.7000 ;
	    RECT 1168.2001 821.4000 1169.4000 822.6000 ;
	    RECT 1165.8000 820.5000 1167.0000 820.8000 ;
	    RECT 1168.2001 820.2000 1169.4000 820.5000 ;
	    RECT 1146.6000 813.3000 1147.8000 819.3000 ;
	    RECT 1149.0000 818.1000 1152.6000 819.3000 ;
	    RECT 1156.2001 818.4000 1157.7001 819.6000 ;
	    RECT 1162.2001 818.4000 1162.5000 819.6000 ;
	    RECT 1163.4000 818.4000 1164.6000 819.6000 ;
	    RECT 1165.8000 819.3000 1167.0000 819.6000 ;
	    RECT 1171.5000 819.3000 1172.7001 822.9000 ;
	    RECT 1175.4000 822.3000 1188.6000 823.5000 ;
	    RECT 1214.4000 822.6000 1215.3000 827.7000 ;
	    RECT 1216.2001 825.4500 1217.4000 825.6000 ;
	    RECT 1216.2001 824.5500 1222.0500 825.4500 ;
	    RECT 1216.2001 824.4000 1217.4000 824.5500 ;
	    RECT 1216.2001 823.2000 1217.4000 823.5000 ;
	    RECT 1180.5000 820.2000 1185.0000 821.4000 ;
	    RECT 1180.5000 819.3000 1181.7001 820.2000 ;
	    RECT 1165.8000 818.4000 1172.7001 819.3000 ;
	    RECT 1151.4000 813.3000 1152.6000 818.1000 ;
	    RECT 1177.8000 818.1000 1181.7001 819.3000 ;
	    RECT 1153.8000 813.3000 1155.0000 817.5000 ;
	    RECT 1156.2001 813.3000 1157.4000 817.5000 ;
	    RECT 1158.6000 813.3000 1159.8000 817.5000 ;
	    RECT 1161.0000 813.3000 1162.2001 817.5000 ;
	    RECT 1163.4000 813.3000 1164.6000 816.3000 ;
	    RECT 1165.8000 813.3000 1167.0000 817.5000 ;
	    RECT 1168.2001 813.3000 1169.4000 816.3000 ;
	    RECT 1170.6000 813.3000 1171.8000 817.5000 ;
	    RECT 1173.0000 813.3000 1174.2001 817.5000 ;
	    RECT 1175.4000 813.3000 1176.6000 817.5000 ;
	    RECT 1177.8000 813.3000 1179.0000 818.1000 ;
	    RECT 1182.6000 813.3000 1183.8000 819.3000 ;
	    RECT 1187.4000 813.3000 1188.6000 822.3000 ;
	    RECT 1211.4000 821.4000 1212.6000 822.6000 ;
	    RECT 1213.5000 821.4000 1215.3000 822.6000 ;
	    RECT 1217.4000 820.8000 1217.7001 822.3000 ;
	    RECT 1218.6000 821.4000 1219.8000 822.6000 ;
	    RECT 1221.1500 822.4500 1222.0500 824.5500 ;
	    RECT 1233.0000 823.5000 1234.2001 839.7000 ;
	    RECT 1235.4000 833.7000 1236.6000 839.7000 ;
	    RECT 1329.0000 837.4500 1330.2001 837.6000 ;
	    RECT 1341.0000 837.4500 1342.2001 837.6000 ;
	    RECT 1329.0000 836.5500 1342.2001 837.4500 ;
	    RECT 1329.0000 836.4000 1330.2001 836.5500 ;
	    RECT 1341.0000 836.4000 1342.2001 836.5500 ;
	    RECT 1369.8000 833.7000 1371.0000 839.7000 ;
	    RECT 1372.2001 834.6000 1373.4000 839.7000 ;
	    RECT 1371.9000 833.7000 1373.4000 834.6000 ;
	    RECT 1374.6000 833.7000 1375.8000 840.6000 ;
	    RECT 1371.9000 832.8000 1372.8000 833.7000 ;
	    RECT 1377.0000 832.8000 1378.2001 839.7000 ;
	    RECT 1379.4000 833.7000 1380.6000 839.7000 ;
	    RECT 1381.8000 835.5000 1383.0000 839.7000 ;
	    RECT 1384.2001 835.5000 1385.4000 839.7000 ;
	    RECT 1369.8000 831.9000 1372.8000 832.8000 ;
	    RECT 1369.8000 823.5000 1371.0000 831.9000 ;
	    RECT 1373.7001 831.6000 1380.0000 832.8000 ;
	    RECT 1386.6000 832.5000 1387.8000 839.7000 ;
	    RECT 1389.0000 833.7000 1390.2001 839.7000 ;
	    RECT 1391.4000 832.5000 1392.6000 839.7000 ;
	    RECT 1393.8000 833.7000 1395.0000 839.7000 ;
	    RECT 1373.7001 831.0000 1374.6000 831.6000 ;
	    RECT 1372.2001 829.8000 1374.6000 831.0000 ;
	    RECT 1379.1000 830.7000 1387.8000 831.6000 ;
	    RECT 1376.1000 829.8000 1378.2001 830.7000 ;
	    RECT 1376.1000 829.5000 1385.4000 829.8000 ;
	    RECT 1377.3000 828.9000 1385.4000 829.5000 ;
	    RECT 1384.2001 828.6000 1385.4000 828.9000 ;
	    RECT 1386.9000 829.5000 1387.8000 830.7000 ;
	    RECT 1388.7001 830.4000 1392.6000 831.6000 ;
	    RECT 1396.2001 830.4000 1397.4000 839.7000 ;
	    RECT 1398.6000 835.5000 1399.8000 839.7000 ;
	    RECT 1401.0000 835.5000 1402.2001 839.7000 ;
	    RECT 1403.4000 835.5000 1404.6000 839.7000 ;
	    RECT 1405.8000 833.7000 1407.0000 839.7000 ;
	    RECT 1401.0000 831.6000 1407.3000 832.8000 ;
	    RECT 1408.2001 831.6000 1409.4000 839.7000 ;
	    RECT 1410.6000 833.7000 1411.8000 839.7000 ;
	    RECT 1413.0000 832.8000 1414.2001 839.7000 ;
	    RECT 1415.4000 833.7000 1416.6000 839.7000 ;
	    RECT 1413.0000 831.9000 1416.9000 832.8000 ;
	    RECT 1417.8000 832.5000 1419.0000 839.7000 ;
	    RECT 1420.2001 833.7000 1421.4000 839.7000 ;
	    RECT 1432.2001 833.7000 1433.4000 839.7000 ;
	    RECT 1408.2001 830.4000 1412.1000 831.6000 ;
	    RECT 1398.6000 829.5000 1399.8000 829.8000 ;
	    RECT 1386.9000 828.6000 1399.8000 829.5000 ;
	    RECT 1403.4000 829.5000 1404.6000 829.8000 ;
	    RECT 1416.0000 829.5000 1416.9000 831.9000 ;
	    RECT 1417.8000 831.4500 1419.0000 831.6000 ;
	    RECT 1422.6000 831.4500 1423.8000 831.6000 ;
	    RECT 1417.8000 830.5500 1423.8000 831.4500 ;
	    RECT 1417.8000 830.4000 1419.0000 830.5500 ;
	    RECT 1422.6000 830.4000 1423.8000 830.5500 ;
	    RECT 1403.4000 828.6000 1416.9000 829.5000 ;
	    RECT 1374.6000 827.4000 1375.8000 828.6000 ;
	    RECT 1379.7001 827.7000 1380.9000 828.0000 ;
	    RECT 1376.7001 826.8000 1415.1000 827.7000 ;
	    RECT 1413.9000 826.5000 1415.1000 826.8000 ;
	    RECT 1416.0000 825.9000 1416.9000 828.6000 ;
	    RECT 1417.8000 828.0000 1419.0000 829.5000 ;
	    RECT 1417.8000 826.8000 1419.3000 828.0000 ;
	    RECT 1371.9000 825.0000 1378.5000 825.9000 ;
	    RECT 1371.9000 824.7000 1373.1000 825.0000 ;
	    RECT 1379.4000 824.4000 1380.6000 825.6000 ;
	    RECT 1381.5000 825.0000 1407.0000 825.9000 ;
	    RECT 1416.0000 825.0000 1417.2001 825.9000 ;
	    RECT 1405.8000 824.1000 1407.0000 825.0000 ;
	    RECT 1233.0000 822.4500 1234.2001 822.6000 ;
	    RECT 1221.1500 821.5500 1234.2001 822.4500 ;
	    RECT 1233.0000 821.4000 1234.2001 821.5500 ;
	    RECT 1369.8000 822.3000 1383.0000 823.5000 ;
	    RECT 1383.9000 822.9000 1386.9000 824.1000 ;
	    RECT 1392.6000 822.9000 1397.4000 824.1000 ;
	    RECT 1211.7001 819.3000 1212.6000 820.5000 ;
	    RECT 1214.1000 819.3000 1219.5000 819.9000 ;
	    RECT 1211.4000 813.3000 1212.6000 819.3000 ;
	    RECT 1213.8000 819.0000 1219.8000 819.3000 ;
	    RECT 1213.8000 813.3000 1215.0000 819.0000 ;
	    RECT 1216.2001 813.3000 1217.4000 818.1000 ;
	    RECT 1218.6000 813.3000 1219.8000 819.0000 ;
	    RECT 1233.0000 813.3000 1234.2001 820.5000 ;
	    RECT 1235.4000 819.4500 1236.6000 819.6000 ;
	    RECT 1348.2001 819.4500 1349.4000 819.6000 ;
	    RECT 1235.4000 818.5500 1349.4000 819.4500 ;
	    RECT 1235.4000 818.4000 1236.6000 818.5500 ;
	    RECT 1348.2001 818.4000 1349.4000 818.5500 ;
	    RECT 1235.4000 817.2000 1236.6000 817.5000 ;
	    RECT 1235.4000 813.3000 1236.6000 816.3000 ;
	    RECT 1369.8000 813.3000 1371.0000 822.3000 ;
	    RECT 1373.4000 820.2000 1377.9000 821.4000 ;
	    RECT 1376.7001 819.3000 1377.9000 820.2000 ;
	    RECT 1385.7001 819.3000 1386.9000 822.9000 ;
	    RECT 1389.0000 821.4000 1390.2001 822.6000 ;
	    RECT 1396.8000 821.7000 1398.0000 822.0000 ;
	    RECT 1391.4000 820.8000 1398.0000 821.7000 ;
	    RECT 1391.4000 820.5000 1392.6000 820.8000 ;
	    RECT 1389.0000 820.2000 1390.2001 820.5000 ;
	    RECT 1401.0000 819.6000 1402.2001 823.8000 ;
	    RECT 1409.7001 822.9000 1415.4000 824.1000 ;
	    RECT 1409.7001 821.1000 1410.9000 822.9000 ;
	    RECT 1416.3000 822.0000 1417.2001 825.0000 ;
	    RECT 1391.4000 819.3000 1392.6000 819.6000 ;
	    RECT 1374.6000 813.3000 1375.8000 819.3000 ;
	    RECT 1376.7001 818.1000 1380.6000 819.3000 ;
	    RECT 1385.7001 818.4000 1392.6000 819.3000 ;
	    RECT 1393.8000 818.4000 1395.0000 819.6000 ;
	    RECT 1395.9000 818.4000 1396.2001 819.6000 ;
	    RECT 1400.7001 818.4000 1402.2001 819.6000 ;
	    RECT 1408.2001 820.2000 1410.9000 821.1000 ;
	    RECT 1415.4000 821.1000 1417.2001 822.0000 ;
	    RECT 1408.2001 819.3000 1409.4000 820.2000 ;
	    RECT 1379.4000 813.3000 1380.6000 818.1000 ;
	    RECT 1405.8000 818.1000 1409.4000 819.3000 ;
	    RECT 1381.8000 813.3000 1383.0000 817.5000 ;
	    RECT 1384.2001 813.3000 1385.4000 817.5000 ;
	    RECT 1386.6000 813.3000 1387.8000 817.5000 ;
	    RECT 1389.0000 813.3000 1390.2001 816.3000 ;
	    RECT 1391.4000 813.3000 1392.6000 817.5000 ;
	    RECT 1393.8000 813.3000 1395.0000 816.3000 ;
	    RECT 1396.2001 813.3000 1397.4000 817.5000 ;
	    RECT 1398.6000 813.3000 1399.8000 817.5000 ;
	    RECT 1401.0000 813.3000 1402.2001 817.5000 ;
	    RECT 1403.4000 813.3000 1404.6000 817.5000 ;
	    RECT 1405.8000 813.3000 1407.0000 818.1000 ;
	    RECT 1410.6000 813.3000 1411.8000 819.3000 ;
	    RECT 1415.4000 813.3000 1416.6000 821.1000 ;
	    RECT 1418.1000 820.2000 1419.3000 826.8000 ;
	    RECT 1434.6000 823.5000 1435.8000 839.7000 ;
	    RECT 1461.0000 827.7000 1462.2001 839.7000 ;
	    RECT 1464.9000 828.6000 1466.1000 839.7000 ;
	    RECT 1467.3000 833.7000 1468.5000 839.7000 ;
	    RECT 1467.0000 830.4000 1468.2001 831.6000 ;
	    RECT 1467.3000 829.5000 1468.2001 830.4000 ;
	    RECT 1464.9000 827.7000 1466.4000 828.6000 ;
	    RECT 1463.4000 825.4500 1464.6000 825.6000 ;
	    RECT 1458.7500 824.5500 1464.6000 825.4500 ;
	    RECT 1434.6000 822.4500 1435.8000 822.6000 ;
	    RECT 1458.7500 822.4500 1459.6500 824.5500 ;
	    RECT 1463.4000 824.4000 1464.6000 824.5500 ;
	    RECT 1463.4000 823.2000 1464.6000 823.5000 ;
	    RECT 1465.5000 822.6000 1466.4000 827.7000 ;
	    RECT 1468.2001 828.4500 1469.4000 828.6000 ;
	    RECT 1501.8000 828.4500 1503.0000 828.6000 ;
	    RECT 1468.2001 827.5500 1503.0000 828.4500 ;
	    RECT 1468.2001 827.4000 1469.4000 827.5500 ;
	    RECT 1501.8000 827.4000 1503.0000 827.5500 ;
	    RECT 1537.8000 827.1000 1539.0000 839.7000 ;
	    RECT 1540.2001 828.0000 1541.4000 839.7000 ;
	    RECT 1544.4000 834.6000 1545.6000 839.7000 ;
	    RECT 1542.6000 833.7000 1545.6000 834.6000 ;
	    RECT 1548.6000 833.7000 1549.8000 839.7000 ;
	    RECT 1551.0000 833.7000 1552.2001 839.7000 ;
	    RECT 1553.4000 833.7000 1554.6000 839.7000 ;
	    RECT 1557.3000 833.7000 1559.1000 839.7000 ;
	    RECT 1542.6000 832.5000 1543.8000 833.7000 ;
	    RECT 1551.0000 832.8000 1551.9000 833.7000 ;
	    RECT 1547.7001 831.9000 1553.1000 832.8000 ;
	    RECT 1557.0000 832.5000 1558.2001 833.7000 ;
	    RECT 1547.7001 831.6000 1548.9000 831.9000 ;
	    RECT 1551.9000 831.6000 1553.1000 831.9000 ;
	    RECT 1542.6000 829.5000 1543.8000 829.8000 ;
	    RECT 1549.5000 829.5000 1550.7001 829.8000 ;
	    RECT 1542.6000 828.6000 1550.7001 829.5000 ;
	    RECT 1551.6000 829.5000 1554.9000 830.4000 ;
	    RECT 1551.6000 827.7000 1552.5000 829.5000 ;
	    RECT 1553.7001 829.2000 1554.9000 829.5000 ;
	    RECT 1557.3000 829.8000 1559.4000 831.0000 ;
	    RECT 1557.3000 828.3000 1558.2001 829.8000 ;
	    RECT 1545.3000 827.1000 1552.5000 827.7000 ;
	    RECT 1537.8000 826.8000 1552.5000 827.1000 ;
	    RECT 1554.6000 827.4000 1558.2001 828.3000 ;
	    RECT 1561.8000 827.7000 1563.0000 839.7000 ;
	    RECT 1537.8000 826.5000 1546.5000 826.8000 ;
	    RECT 1537.8000 826.2000 1546.2001 826.5000 ;
	    RECT 1475.4000 825.4500 1476.6000 825.6000 ;
	    RECT 1533.0000 825.4500 1534.2001 825.6000 ;
	    RECT 1475.4000 824.5500 1534.2001 825.4500 ;
	    RECT 1475.4000 824.4000 1476.6000 824.5500 ;
	    RECT 1533.0000 824.4000 1534.2001 824.5500 ;
	    RECT 1541.1000 824.4000 1546.5000 825.3000 ;
	    RECT 1547.4000 824.4000 1548.6000 825.6000 ;
	    RECT 1541.1000 824.1000 1542.3000 824.4000 ;
	    RECT 1543.5000 822.6000 1544.7001 822.9000 ;
	    RECT 1554.6000 822.6000 1555.5000 827.4000 ;
	    RECT 1564.2001 826.8000 1565.4000 839.7000 ;
	    RECT 1559.1000 826.5000 1565.4000 826.8000 ;
	    RECT 1559.1000 825.9000 1563.3000 826.5000 ;
	    RECT 1559.1000 825.6000 1560.3000 825.9000 ;
	    RECT 1561.5000 824.7000 1562.7001 825.0000 ;
	    RECT 1557.0000 823.8000 1562.7001 824.7000 ;
	    RECT 1564.2001 824.4000 1565.4000 825.6000 ;
	    RECT 1557.0000 823.5000 1558.2001 823.8000 ;
	    RECT 1434.6000 821.5500 1459.6500 822.4500 ;
	    RECT 1434.6000 821.4000 1435.8000 821.5500 ;
	    RECT 1461.0000 821.4000 1462.2001 822.6000 ;
	    RECT 1463.1000 820.8000 1463.4000 822.3000 ;
	    RECT 1465.5000 821.4000 1467.3000 822.6000 ;
	    RECT 1468.2001 822.4500 1469.4000 822.6000 ;
	    RECT 1535.4000 822.4500 1536.6000 822.6000 ;
	    RECT 1468.2001 821.5500 1536.6000 822.4500 ;
	    RECT 1468.2001 821.4000 1469.4000 821.5500 ;
	    RECT 1535.4000 821.4000 1536.6000 821.5500 ;
	    RECT 1539.0000 821.4000 1539.3000 822.6000 ;
	    RECT 1540.2001 821.4000 1541.4000 822.6000 ;
	    RECT 1542.3000 821.7000 1555.5000 822.6000 ;
	    RECT 1417.8000 819.0000 1419.3000 820.2000 ;
	    RECT 1417.8000 813.3000 1419.0000 819.0000 ;
	    RECT 1432.2001 818.4000 1433.4000 819.6000 ;
	    RECT 1432.2001 817.2000 1433.4000 817.5000 ;
	    RECT 1420.2001 813.3000 1421.4000 816.3000 ;
	    RECT 1432.2001 813.3000 1433.4000 816.3000 ;
	    RECT 1434.6000 813.3000 1435.8000 820.5000 ;
	    RECT 1461.3000 819.3000 1466.7001 819.9000 ;
	    RECT 1468.2001 819.3000 1469.1000 820.5000 ;
	    RECT 1461.0000 819.0000 1467.0000 819.3000 ;
	    RECT 1461.0000 813.3000 1462.2001 819.0000 ;
	    RECT 1463.4000 813.3000 1464.6000 818.1000 ;
	    RECT 1465.8000 813.3000 1467.0000 819.0000 ;
	    RECT 1468.2001 813.3000 1469.4000 819.3000 ;
	    RECT 1537.8000 813.3000 1539.0000 820.5000 ;
	    RECT 1540.2001 813.3000 1541.4000 819.3000 ;
	    RECT 1545.3000 818.4000 1546.2001 821.7000 ;
	    RECT 1553.7001 821.4000 1554.9000 821.7000 ;
	    RECT 1564.2001 820.8000 1565.4000 823.5000 ;
	    RECT 1559.7001 819.9000 1565.4000 820.8000 ;
	    RECT 1559.7001 819.6000 1560.9000 819.9000 ;
	    RECT 1542.6000 816.3000 1543.8000 817.5000 ;
	    RECT 1545.0000 817.2000 1546.2001 818.4000 ;
	    RECT 1547.7001 818.1000 1548.9000 818.4000 ;
	    RECT 1547.7001 817.2000 1551.9000 818.1000 ;
	    RECT 1551.0000 816.3000 1551.9000 817.2000 ;
	    RECT 1557.0000 816.3000 1558.2001 817.5000 ;
	    RECT 1542.6000 815.4000 1545.6000 816.3000 ;
	    RECT 1544.4000 813.3000 1545.6000 815.4000 ;
	    RECT 1548.3000 813.3000 1549.8000 816.3000 ;
	    RECT 1551.0000 813.3000 1552.2001 816.3000 ;
	    RECT 1553.4000 813.3000 1554.6000 816.3000 ;
	    RECT 1557.0000 815.4000 1559.1000 816.3000 ;
	    RECT 1557.3000 813.3000 1559.1000 815.4000 ;
	    RECT 1561.8000 813.3000 1563.0000 819.0000 ;
	    RECT 1564.2001 813.3000 1565.4000 819.9000 ;
	    RECT 1.2000 810.6000 1569.0000 812.4000 ;
	    RECT 124.2000 806.7000 125.4000 809.7000 ;
	    RECT 126.6000 804.0000 127.8000 809.7000 ;
	    RECT 126.3000 802.8000 127.8000 804.0000 ;
	    RECT 126.3000 796.2000 127.5000 802.8000 ;
	    RECT 129.0000 801.9000 130.2000 809.7000 ;
	    RECT 133.8000 803.7000 135.0000 809.7000 ;
	    RECT 138.6000 804.9000 139.8000 809.7000 ;
	    RECT 141.0000 805.5000 142.2000 809.7000 ;
	    RECT 143.4000 805.5000 144.6000 809.7000 ;
	    RECT 145.8000 805.5000 147.0000 809.7000 ;
	    RECT 148.2000 805.5000 149.4000 809.7000 ;
	    RECT 150.6000 806.7000 151.8000 809.7000 ;
	    RECT 153.0000 805.5000 154.2000 809.7000 ;
	    RECT 155.4000 806.7000 156.6000 809.7000 ;
	    RECT 157.8000 805.5000 159.0000 809.7000 ;
	    RECT 160.2000 805.5000 161.4000 809.7000 ;
	    RECT 162.6000 805.5000 163.8000 809.7000 ;
	    RECT 136.2000 803.7000 139.8000 804.9000 ;
	    RECT 165.0000 804.9000 166.2000 809.7000 ;
	    RECT 136.2000 802.8000 137.4000 803.7000 ;
	    RECT 128.4000 801.0000 130.2000 801.9000 ;
	    RECT 134.7000 801.9000 137.4000 802.8000 ;
	    RECT 143.4000 803.4000 144.9000 804.6000 ;
	    RECT 149.4000 803.4000 149.7000 804.6000 ;
	    RECT 150.6000 803.4000 151.8000 804.6000 ;
	    RECT 153.0000 803.7000 159.9000 804.6000 ;
	    RECT 165.0000 803.7000 168.9000 804.9000 ;
	    RECT 169.8000 803.7000 171.0000 809.7000 ;
	    RECT 153.0000 803.4000 154.2000 803.7000 ;
	    RECT 128.4000 798.0000 129.3000 801.0000 ;
	    RECT 134.7000 800.1000 135.9000 801.9000 ;
	    RECT 130.2000 798.9000 135.9000 800.1000 ;
	    RECT 143.4000 799.2000 144.6000 803.4000 ;
	    RECT 155.4000 802.5000 156.6000 802.8000 ;
	    RECT 153.0000 802.2000 154.2000 802.5000 ;
	    RECT 147.6000 801.3000 154.2000 802.2000 ;
	    RECT 147.6000 801.0000 148.8000 801.3000 ;
	    RECT 155.4000 800.4000 156.6000 801.6000 ;
	    RECT 158.7000 800.1000 159.9000 803.7000 ;
	    RECT 167.7000 802.8000 168.9000 803.7000 ;
	    RECT 167.7000 801.6000 172.2000 802.8000 ;
	    RECT 174.6000 800.7000 175.8000 809.7000 ;
	    RECT 186.6000 806.7000 187.8000 809.7000 ;
	    RECT 186.6000 805.5000 187.8000 805.8000 ;
	    RECT 186.6000 803.4000 187.8000 804.6000 ;
	    RECT 189.0000 802.5000 190.2000 809.7000 ;
	    RECT 210.6000 806.7000 211.8000 809.7000 ;
	    RECT 210.6000 805.5000 211.8000 805.8000 ;
	    RECT 203.4000 804.4500 204.6000 804.6000 ;
	    RECT 210.6000 804.4500 211.8000 804.6000 ;
	    RECT 203.4000 803.5500 211.8000 804.4500 ;
	    RECT 203.4000 803.4000 204.6000 803.5500 ;
	    RECT 210.6000 803.4000 211.8000 803.5500 ;
	    RECT 213.0000 802.5000 214.2000 809.7000 ;
	    RECT 244.2000 804.0000 245.4000 809.7000 ;
	    RECT 246.6000 804.9000 247.8000 809.7000 ;
	    RECT 249.0000 808.8000 255.0000 809.7000 ;
	    RECT 249.0000 804.0000 250.2000 808.8000 ;
	    RECT 244.2000 803.7000 250.2000 804.0000 ;
	    RECT 251.4000 803.7000 252.6000 807.9000 ;
	    RECT 253.8000 803.7000 255.0000 808.8000 ;
	    RECT 244.5000 803.1000 249.9000 803.7000 ;
	    RECT 148.2000 798.9000 153.0000 800.1000 ;
	    RECT 158.7000 798.9000 161.7000 800.1000 ;
	    RECT 162.6000 799.5000 175.8000 800.7000 ;
	    RECT 189.0000 801.4500 190.2000 801.6000 ;
	    RECT 210.6000 801.4500 211.8000 801.6000 ;
	    RECT 189.0000 800.5500 211.8000 801.4500 ;
	    RECT 189.0000 800.4000 190.2000 800.5500 ;
	    RECT 210.6000 800.4000 211.8000 800.5500 ;
	    RECT 213.0000 801.4500 214.2000 801.6000 ;
	    RECT 222.6000 801.4500 223.8000 801.6000 ;
	    RECT 213.0000 800.5500 223.8000 801.4500 ;
	    RECT 213.0000 800.4000 214.2000 800.5500 ;
	    RECT 222.6000 800.4000 223.8000 800.5500 ;
	    RECT 225.0000 801.4500 226.2000 801.6000 ;
	    RECT 244.2000 801.4500 245.4000 801.6000 ;
	    RECT 225.0000 800.5500 245.4000 801.4500 ;
	    RECT 246.3000 800.7000 246.6000 802.2000 ;
	    RECT 251.7000 801.6000 252.6000 803.7000 ;
	    RECT 268.2000 802.5000 269.4000 809.7000 ;
	    RECT 270.6000 806.7000 271.8000 809.7000 ;
	    RECT 270.6000 805.5000 271.8000 805.8000 ;
	    RECT 270.6000 803.4000 271.8000 804.6000 ;
	    RECT 323.4000 803.7000 324.6000 809.7000 ;
	    RECT 325.8000 802.8000 327.0000 809.7000 ;
	    RECT 328.2000 803.7000 329.4000 809.7000 ;
	    RECT 330.6000 802.8000 331.8000 809.7000 ;
	    RECT 333.0000 803.7000 334.2000 809.7000 ;
	    RECT 335.4000 802.8000 336.6000 809.7000 ;
	    RECT 337.8000 803.7000 339.0000 809.7000 ;
	    RECT 340.2000 802.8000 341.4000 809.7000 ;
	    RECT 342.6000 803.7000 343.8000 809.7000 ;
	    RECT 325.8000 801.6000 328.5000 802.8000 ;
	    RECT 330.6000 801.6000 333.9000 802.8000 ;
	    RECT 335.4000 801.6000 338.7000 802.8000 ;
	    RECT 340.2000 801.6000 343.8000 802.8000 ;
	    RECT 357.0000 802.5000 358.2000 809.7000 ;
	    RECT 359.4000 806.7000 360.6000 809.7000 ;
	    RECT 359.4000 805.5000 360.6000 805.8000 ;
	    RECT 359.4000 804.4500 360.6000 804.6000 ;
	    RECT 383.4000 804.4500 384.6000 804.6000 ;
	    RECT 359.4000 803.5500 384.6000 804.4500 ;
	    RECT 385.8000 804.0000 387.0000 809.7000 ;
	    RECT 388.2000 804.9000 389.4000 809.7000 ;
	    RECT 390.6000 804.0000 391.8000 809.7000 ;
	    RECT 385.8000 803.7000 391.8000 804.0000 ;
	    RECT 393.0000 803.7000 394.2000 809.7000 ;
	    RECT 412.2000 803.7000 413.4000 809.7000 ;
	    RECT 416.1000 804.6000 417.3000 809.7000 ;
	    RECT 429.0000 806.7000 430.2000 809.7000 ;
	    RECT 429.0000 805.5000 430.2000 805.8000 ;
	    RECT 414.6000 803.7000 417.3000 804.6000 ;
	    RECT 359.4000 803.4000 360.6000 803.5500 ;
	    RECT 383.4000 803.4000 384.6000 803.5500 ;
	    RECT 386.1000 803.1000 391.5000 803.7000 ;
	    RECT 393.0000 802.5000 393.9000 803.7000 ;
	    RECT 412.2000 802.5000 413.4000 802.8000 ;
	    RECT 225.0000 800.4000 226.2000 800.5500 ;
	    RECT 244.2000 800.4000 245.4000 800.5500 ;
	    RECT 249.0000 800.4000 250.2000 801.6000 ;
	    RECT 251.1000 800.7000 252.6000 801.6000 ;
	    RECT 253.8000 800.4000 255.0000 801.6000 ;
	    RECT 256.2000 801.4500 257.4000 801.6000 ;
	    RECT 268.2000 801.4500 269.4000 801.6000 ;
	    RECT 256.2000 800.5500 269.4000 801.4500 ;
	    RECT 256.2000 800.4000 257.4000 800.5500 ;
	    RECT 268.2000 800.4000 269.4000 800.5500 ;
	    RECT 285.0000 801.4500 286.2000 801.6000 ;
	    RECT 323.4000 801.4500 324.6000 801.6000 ;
	    RECT 285.0000 800.5500 324.6000 801.4500 ;
	    RECT 327.3000 800.7000 328.5000 801.6000 ;
	    RECT 332.7000 800.7000 333.9000 801.6000 ;
	    RECT 337.5000 800.7000 338.7000 801.6000 ;
	    RECT 285.0000 800.4000 286.2000 800.5500 ;
	    RECT 323.4000 800.4000 324.6000 800.5500 ;
	    RECT 246.6000 799.5000 247.8000 799.8000 ;
	    RECT 251.4000 799.5000 252.6000 799.8000 ;
	    RECT 325.5000 799.5000 326.1000 800.7000 ;
	    RECT 327.3000 799.5000 331.2000 800.7000 ;
	    RECT 332.7000 799.5000 336.3000 800.7000 ;
	    RECT 337.5000 799.5000 341.4000 800.7000 ;
	    RECT 342.6000 799.5000 343.8000 801.6000 ;
	    RECT 347.4000 801.4500 348.6000 801.6000 ;
	    RECT 357.0000 801.4500 358.2000 801.6000 ;
	    RECT 347.4000 800.5500 358.2000 801.4500 ;
	    RECT 347.4000 800.4000 348.6000 800.5500 ;
	    RECT 357.0000 800.4000 358.2000 800.5500 ;
	    RECT 369.0000 801.4500 370.2000 801.6000 ;
	    RECT 385.8000 801.4500 387.0000 801.6000 ;
	    RECT 369.0000 800.5500 387.0000 801.4500 ;
	    RECT 387.9000 800.7000 388.2000 802.2000 ;
	    RECT 369.0000 800.4000 370.2000 800.5500 ;
	    RECT 385.8000 800.4000 387.0000 800.5500 ;
	    RECT 390.3000 800.4000 392.1000 801.6000 ;
	    RECT 393.0000 800.4000 394.2000 801.6000 ;
	    RECT 412.2000 800.4000 413.4000 801.6000 ;
	    RECT 388.2000 799.5000 389.4000 799.8000 ;
	    RECT 138.6000 798.0000 139.8000 798.9000 ;
	    RECT 128.4000 797.1000 129.6000 798.0000 ;
	    RECT 138.6000 797.1000 164.1000 798.0000 ;
	    RECT 165.0000 797.4000 166.2000 798.6000 ;
	    RECT 172.5000 798.0000 173.7000 798.3000 ;
	    RECT 167.1000 797.1000 173.7000 798.0000 ;
	    RECT 126.3000 795.0000 127.8000 796.2000 ;
	    RECT 126.6000 793.5000 127.8000 795.0000 ;
	    RECT 128.7000 794.4000 129.6000 797.1000 ;
	    RECT 130.5000 796.2000 131.7000 796.5000 ;
	    RECT 130.5000 795.3000 168.9000 796.2000 ;
	    RECT 164.7000 795.0000 165.9000 795.3000 ;
	    RECT 169.8000 794.4000 171.0000 795.6000 ;
	    RECT 128.7000 793.5000 142.2000 794.4000 ;
	    RECT 71.4000 792.4500 72.6000 792.6000 ;
	    RECT 126.6000 792.4500 127.8000 792.6000 ;
	    RECT 71.4000 791.5500 127.8000 792.4500 ;
	    RECT 71.4000 791.4000 72.6000 791.5500 ;
	    RECT 126.6000 791.4000 127.8000 791.5500 ;
	    RECT 128.7000 791.1000 129.6000 793.5000 ;
	    RECT 141.0000 793.2000 142.2000 793.5000 ;
	    RECT 145.8000 793.5000 158.7000 794.4000 ;
	    RECT 145.8000 793.2000 147.0000 793.5000 ;
	    RECT 133.5000 791.4000 137.4000 792.6000 ;
	    RECT 124.2000 783.3000 125.4000 789.3000 ;
	    RECT 126.6000 783.3000 127.8000 790.5000 ;
	    RECT 128.7000 790.2000 132.6000 791.1000 ;
	    RECT 129.0000 783.3000 130.2000 789.3000 ;
	    RECT 131.4000 783.3000 132.6000 790.2000 ;
	    RECT 133.8000 783.3000 135.0000 789.3000 ;
	    RECT 136.2000 783.3000 137.4000 791.4000 ;
	    RECT 138.3000 790.2000 144.6000 791.4000 ;
	    RECT 138.6000 783.3000 139.8000 789.3000 ;
	    RECT 141.0000 783.3000 142.2000 787.5000 ;
	    RECT 143.4000 783.3000 144.6000 787.5000 ;
	    RECT 145.8000 783.3000 147.0000 787.5000 ;
	    RECT 148.2000 783.3000 149.4000 792.6000 ;
	    RECT 153.0000 791.4000 156.9000 792.6000 ;
	    RECT 157.8000 792.3000 158.7000 793.5000 ;
	    RECT 160.2000 794.1000 161.4000 794.4000 ;
	    RECT 160.2000 793.5000 168.3000 794.1000 ;
	    RECT 160.2000 793.2000 169.5000 793.5000 ;
	    RECT 167.4000 792.3000 169.5000 793.2000 ;
	    RECT 157.8000 791.4000 166.5000 792.3000 ;
	    RECT 171.0000 792.0000 173.4000 793.2000 ;
	    RECT 171.0000 791.4000 171.9000 792.0000 ;
	    RECT 150.6000 783.3000 151.8000 789.3000 ;
	    RECT 153.0000 783.3000 154.2000 790.5000 ;
	    RECT 155.4000 783.3000 156.6000 789.3000 ;
	    RECT 157.8000 783.3000 159.0000 790.5000 ;
	    RECT 165.6000 790.2000 171.9000 791.4000 ;
	    RECT 174.6000 791.1000 175.8000 799.5000 ;
	    RECT 172.8000 790.2000 175.8000 791.1000 ;
	    RECT 160.2000 783.3000 161.4000 787.5000 ;
	    RECT 162.6000 783.3000 163.8000 787.5000 ;
	    RECT 165.0000 783.3000 166.2000 789.3000 ;
	    RECT 167.4000 783.3000 168.6000 790.2000 ;
	    RECT 172.8000 789.3000 173.7000 790.2000 ;
	    RECT 169.8000 782.4000 171.0000 789.3000 ;
	    RECT 172.2000 788.4000 173.7000 789.3000 ;
	    RECT 172.2000 783.3000 173.4000 788.4000 ;
	    RECT 174.6000 783.3000 175.8000 789.3000 ;
	    RECT 186.6000 783.3000 187.8000 789.3000 ;
	    RECT 189.0000 783.3000 190.2000 799.5000 ;
	    RECT 210.6000 783.3000 211.8000 789.3000 ;
	    RECT 213.0000 783.3000 214.2000 799.5000 ;
	    RECT 232.2000 798.4500 233.4000 798.6000 ;
	    RECT 246.6000 798.4500 247.8000 798.6000 ;
	    RECT 232.2000 797.5500 247.8000 798.4500 ;
	    RECT 232.2000 797.4000 233.4000 797.5500 ;
	    RECT 246.6000 797.4000 247.8000 797.5500 ;
	    RECT 249.0000 795.3000 249.9000 799.5000 ;
	    RECT 253.8000 799.2000 255.0000 799.5000 ;
	    RECT 251.4000 797.4000 252.6000 798.6000 ;
	    RECT 244.2000 783.3000 245.4000 795.3000 ;
	    RECT 248.1000 783.3000 251.1000 795.3000 ;
	    RECT 253.8000 783.3000 255.0000 795.3000 ;
	    RECT 268.2000 783.3000 269.4000 799.5000 ;
	    RECT 327.3000 797.4000 328.5000 799.5000 ;
	    RECT 332.7000 797.4000 333.9000 799.5000 ;
	    RECT 337.5000 797.4000 338.7000 799.5000 ;
	    RECT 342.6000 798.4500 343.8000 798.6000 ;
	    RECT 354.6000 798.4500 355.8000 798.6000 ;
	    RECT 342.6000 797.5500 355.8000 798.4500 ;
	    RECT 342.6000 797.4000 343.8000 797.5500 ;
	    RECT 354.6000 797.4000 355.8000 797.5500 ;
	    RECT 325.8000 796.2000 328.5000 797.4000 ;
	    RECT 330.6000 796.2000 333.9000 797.4000 ;
	    RECT 335.4000 796.2000 338.7000 797.4000 ;
	    RECT 340.2000 796.5000 341.7000 797.4000 ;
	    RECT 340.2000 796.2000 343.8000 796.5000 ;
	    RECT 270.6000 783.3000 271.8000 789.3000 ;
	    RECT 323.4000 783.3000 324.6000 795.3000 ;
	    RECT 325.8000 783.3000 327.0000 796.2000 ;
	    RECT 328.2000 783.3000 329.4000 795.3000 ;
	    RECT 330.6000 783.3000 331.8000 796.2000 ;
	    RECT 333.0000 783.3000 334.2000 795.3000 ;
	    RECT 335.4000 783.3000 336.6000 796.2000 ;
	    RECT 337.8000 783.3000 339.0000 795.3000 ;
	    RECT 340.2000 783.3000 341.4000 796.2000 ;
	    RECT 342.6000 783.3000 343.8000 795.3000 ;
	    RECT 357.0000 783.3000 358.2000 799.5000 ;
	    RECT 381.0000 798.4500 382.2000 798.6000 ;
	    RECT 388.2000 798.4500 389.4000 798.6000 ;
	    RECT 381.0000 797.5500 389.4000 798.4500 ;
	    RECT 381.0000 797.4000 382.2000 797.5500 ;
	    RECT 388.2000 797.4000 389.4000 797.5500 ;
	    RECT 390.3000 795.3000 391.2000 800.4000 ;
	    RECT 414.6000 799.5000 415.8000 803.7000 ;
	    RECT 429.0000 803.4000 430.2000 804.6000 ;
	    RECT 431.4000 802.5000 432.6000 809.7000 ;
	    RECT 419.4000 801.4500 420.6000 801.6000 ;
	    RECT 431.4000 801.4500 432.6000 801.6000 ;
	    RECT 419.4000 800.5500 432.6000 801.4500 ;
	    RECT 419.4000 800.4000 420.6000 800.5500 ;
	    RECT 431.4000 800.4000 432.6000 800.5500 ;
	    RECT 563.4000 800.7000 564.6000 809.7000 ;
	    RECT 568.2000 803.7000 569.4000 809.7000 ;
	    RECT 573.0000 804.9000 574.2000 809.7000 ;
	    RECT 575.4000 805.5000 576.6000 809.7000 ;
	    RECT 577.8000 805.5000 579.0000 809.7000 ;
	    RECT 580.2000 805.5000 581.4000 809.7000 ;
	    RECT 582.6000 806.7000 583.8000 809.7000 ;
	    RECT 585.0000 805.5000 586.2000 809.7000 ;
	    RECT 587.4000 806.7000 588.6000 809.7000 ;
	    RECT 589.8000 805.5000 591.0000 809.7000 ;
	    RECT 592.2000 805.5000 593.4000 809.7000 ;
	    RECT 594.6000 805.5000 595.8000 809.7000 ;
	    RECT 597.0000 805.5000 598.2000 809.7000 ;
	    RECT 570.3000 803.7000 574.2000 804.9000 ;
	    RECT 599.4000 804.9000 600.6000 809.7000 ;
	    RECT 579.3000 803.7000 586.2000 804.6000 ;
	    RECT 570.3000 802.8000 571.5000 803.7000 ;
	    RECT 567.0000 801.6000 571.5000 802.8000 ;
	    RECT 563.4000 799.5000 576.6000 800.7000 ;
	    RECT 579.3000 800.1000 580.5000 803.7000 ;
	    RECT 585.0000 803.4000 586.2000 803.7000 ;
	    RECT 587.4000 803.4000 588.6000 804.6000 ;
	    RECT 589.5000 803.4000 589.8000 804.6000 ;
	    RECT 594.3000 803.4000 595.8000 804.6000 ;
	    RECT 599.4000 803.7000 603.0000 804.9000 ;
	    RECT 604.2000 803.7000 605.4000 809.7000 ;
	    RECT 582.6000 802.5000 583.8000 802.8000 ;
	    RECT 585.0000 802.2000 586.2000 802.5000 ;
	    RECT 582.6000 800.4000 583.8000 801.6000 ;
	    RECT 585.0000 801.3000 591.6000 802.2000 ;
	    RECT 590.4000 801.0000 591.6000 801.3000 ;
	    RECT 414.6000 798.4500 415.8000 798.6000 ;
	    RECT 393.1500 797.5500 415.8000 798.4500 ;
	    RECT 393.1500 795.6000 394.0500 797.5500 ;
	    RECT 414.6000 797.4000 415.8000 797.5500 ;
	    RECT 359.4000 783.3000 360.6000 789.3000 ;
	    RECT 385.8000 783.3000 387.0000 795.3000 ;
	    RECT 389.7000 794.4000 391.2000 795.3000 ;
	    RECT 393.0000 794.4000 394.2000 795.6000 ;
	    RECT 389.7000 783.3000 390.9000 794.4000 ;
	    RECT 392.1000 792.6000 393.0000 793.5000 ;
	    RECT 391.8000 791.4000 393.0000 792.6000 ;
	    RECT 392.1000 783.3000 393.3000 789.3000 ;
	    RECT 412.2000 783.3000 413.4000 789.3000 ;
	    RECT 414.6000 783.3000 415.8000 796.5000 ;
	    RECT 417.0000 795.4500 418.2000 795.6000 ;
	    RECT 429.0000 795.4500 430.2000 795.6000 ;
	    RECT 417.0000 794.5500 430.2000 795.4500 ;
	    RECT 417.0000 794.4000 418.2000 794.5500 ;
	    RECT 429.0000 794.4000 430.2000 794.5500 ;
	    RECT 417.0000 793.2000 418.2000 793.5000 ;
	    RECT 417.0000 783.3000 418.2000 789.3000 ;
	    RECT 429.0000 783.3000 430.2000 789.3000 ;
	    RECT 431.4000 783.3000 432.6000 799.5000 ;
	    RECT 563.4000 791.1000 564.6000 799.5000 ;
	    RECT 577.5000 798.9000 580.5000 800.1000 ;
	    RECT 586.2000 798.9000 591.0000 800.1000 ;
	    RECT 594.6000 799.2000 595.8000 803.4000 ;
	    RECT 601.8000 802.8000 603.0000 803.7000 ;
	    RECT 601.8000 801.9000 604.5000 802.8000 ;
	    RECT 603.3000 800.1000 604.5000 801.9000 ;
	    RECT 609.0000 801.9000 610.2000 809.7000 ;
	    RECT 611.4000 804.0000 612.6000 809.7000 ;
	    RECT 613.8000 806.7000 615.0000 809.7000 ;
	    RECT 611.4000 802.8000 612.9000 804.0000 ;
	    RECT 633.0000 803.7000 634.2000 809.7000 ;
	    RECT 636.9000 804.6000 638.1000 809.7000 ;
	    RECT 635.4000 803.7000 638.1000 804.6000 ;
	    RECT 669.0000 803.7000 670.2000 809.7000 ;
	    RECT 672.9000 804.0000 674.1000 809.7000 ;
	    RECT 675.3000 805.2000 676.5000 809.7000 ;
	    RECT 690.6000 806.7000 691.8000 809.7000 ;
	    RECT 690.6000 805.5000 691.8000 805.8000 ;
	    RECT 675.3000 803.7000 677.4000 805.2000 ;
	    RECT 609.0000 801.0000 610.8000 801.9000 ;
	    RECT 603.3000 798.9000 609.0000 800.1000 ;
	    RECT 565.5000 798.0000 566.7000 798.3000 ;
	    RECT 565.5000 797.1000 572.1000 798.0000 ;
	    RECT 573.0000 797.4000 574.2000 798.6000 ;
	    RECT 599.4000 798.0000 600.6000 798.9000 ;
	    RECT 609.9000 798.0000 610.8000 801.0000 ;
	    RECT 575.1000 797.1000 600.6000 798.0000 ;
	    RECT 609.6000 797.1000 610.8000 798.0000 ;
	    RECT 607.5000 796.2000 608.7000 796.5000 ;
	    RECT 568.2000 794.4000 569.4000 795.6000 ;
	    RECT 570.3000 795.3000 608.7000 796.2000 ;
	    RECT 573.3000 795.0000 574.5000 795.3000 ;
	    RECT 609.6000 794.4000 610.5000 797.1000 ;
	    RECT 611.7000 796.2000 612.9000 802.8000 ;
	    RECT 633.0000 802.5000 634.2000 802.8000 ;
	    RECT 628.2000 801.4500 629.4000 801.6000 ;
	    RECT 633.0000 801.4500 634.2000 801.6000 ;
	    RECT 628.2000 800.5500 634.2000 801.4500 ;
	    RECT 628.2000 800.4000 629.4000 800.5500 ;
	    RECT 633.0000 800.4000 634.2000 800.5500 ;
	    RECT 635.4000 799.5000 636.6000 803.7000 ;
	    RECT 669.3000 803.4000 670.2000 803.7000 ;
	    RECT 669.3000 802.8000 672.0000 803.4000 ;
	    RECT 669.3000 802.5000 675.6000 802.8000 ;
	    RECT 671.1000 801.9000 675.6000 802.5000 ;
	    RECT 674.4000 801.6000 675.6000 801.9000 ;
	    RECT 637.8000 801.4500 639.0000 801.6000 ;
	    RECT 669.0000 801.4500 670.2000 801.6000 ;
	    RECT 637.8000 800.5500 670.2000 801.4500 ;
	    RECT 672.0000 800.7000 673.2000 801.0000 ;
	    RECT 637.8000 800.4000 639.0000 800.5500 ;
	    RECT 669.0000 800.4000 670.2000 800.5500 ;
	    RECT 671.7000 799.8000 673.2000 800.7000 ;
	    RECT 671.7000 799.5000 672.6000 799.8000 ;
	    RECT 669.0000 799.2000 670.2000 799.5000 ;
	    RECT 635.4000 798.4500 636.6000 798.6000 ;
	    RECT 642.6000 798.4500 643.8000 798.6000 ;
	    RECT 635.4000 797.5500 643.8000 798.4500 ;
	    RECT 635.4000 797.4000 636.6000 797.5500 ;
	    RECT 642.6000 797.4000 643.8000 797.5500 ;
	    RECT 671.4000 797.4000 672.6000 798.6000 ;
	    RECT 674.4000 796.5000 675.3000 801.6000 ;
	    RECT 676.5000 799.5000 677.4000 803.7000 ;
	    RECT 678.6000 804.4500 679.8000 804.6000 ;
	    RECT 690.6000 804.4500 691.8000 804.6000 ;
	    RECT 678.6000 803.5500 691.8000 804.4500 ;
	    RECT 678.6000 803.4000 679.8000 803.5500 ;
	    RECT 690.6000 803.4000 691.8000 803.5500 ;
	    RECT 693.0000 802.5000 694.2000 809.7000 ;
	    RECT 712.2000 803.7000 713.4000 809.7000 ;
	    RECT 716.1000 804.6000 717.3000 809.7000 ;
	    RECT 714.6000 803.7000 717.3000 804.6000 ;
	    RECT 736.2000 803.7000 737.4000 809.7000 ;
	    RECT 740.1000 804.6000 741.3000 809.7000 ;
	    RECT 760.2000 806.7000 761.4000 809.7000 ;
	    RECT 762.6000 806.7000 763.8000 809.7000 ;
	    RECT 765.0000 806.7000 766.2000 809.7000 ;
	    RECT 738.6000 803.7000 741.3000 804.6000 ;
	    RECT 712.2000 802.5000 713.4000 802.8000 ;
	    RECT 693.0000 801.4500 694.2000 801.6000 ;
	    RECT 709.8000 801.4500 711.0000 801.6000 ;
	    RECT 693.0000 800.5500 711.0000 801.4500 ;
	    RECT 693.0000 800.4000 694.2000 800.5500 ;
	    RECT 709.8000 800.4000 711.0000 800.5500 ;
	    RECT 712.2000 800.4000 713.4000 801.6000 ;
	    RECT 714.6000 799.5000 715.8000 803.7000 ;
	    RECT 736.2000 802.5000 737.4000 802.8000 ;
	    RECT 729.0000 801.4500 730.2000 801.6000 ;
	    RECT 736.2000 801.4500 737.4000 801.6000 ;
	    RECT 729.0000 800.5500 737.4000 801.4500 ;
	    RECT 729.0000 800.4000 730.2000 800.5500 ;
	    RECT 736.2000 800.4000 737.4000 800.5500 ;
	    RECT 738.6000 799.5000 739.8000 803.7000 ;
	    RECT 762.6000 802.5000 763.5000 806.7000 ;
	    RECT 765.0000 805.5000 766.2000 805.8000 ;
	    RECT 785.1000 804.6000 786.3000 809.7000 ;
	    RECT 765.0000 803.4000 766.2000 804.6000 ;
	    RECT 785.1000 803.7000 787.8000 804.6000 ;
	    RECT 789.0000 803.7000 790.2000 809.7000 ;
	    RECT 808.2000 806.7000 809.4000 809.7000 ;
	    RECT 810.6000 806.7000 811.8000 809.7000 ;
	    RECT 813.0000 806.7000 814.2000 809.7000 ;
	    RECT 762.6000 801.4500 763.8000 801.6000 ;
	    RECT 774.6000 801.4500 775.8000 801.6000 ;
	    RECT 762.6000 800.5500 775.8000 801.4500 ;
	    RECT 762.6000 800.4000 763.8000 800.5500 ;
	    RECT 774.6000 800.4000 775.8000 800.5500 ;
	    RECT 786.6000 799.5000 787.8000 803.7000 ;
	    RECT 789.0000 802.5000 790.2000 802.8000 ;
	    RECT 810.6000 802.5000 811.5000 806.7000 ;
	    RECT 813.0000 805.5000 814.2000 805.8000 ;
	    RECT 813.0000 804.4500 814.2000 804.6000 ;
	    RECT 822.6000 804.4500 823.8000 804.6000 ;
	    RECT 813.0000 803.5500 823.8000 804.4500 ;
	    RECT 813.0000 803.4000 814.2000 803.5500 ;
	    RECT 822.6000 803.4000 823.8000 803.5500 ;
	    RECT 789.0000 800.4000 790.2000 801.6000 ;
	    RECT 791.4000 801.4500 792.6000 801.6000 ;
	    RECT 810.6000 801.4500 811.8000 801.6000 ;
	    RECT 791.4000 800.5500 811.8000 801.4500 ;
	    RECT 838.8000 801.3000 840.0000 809.7000 ;
	    RECT 791.4000 800.4000 792.6000 800.5500 ;
	    RECT 810.6000 800.4000 811.8000 800.5500 ;
	    RECT 837.3000 800.7000 840.0000 801.3000 ;
	    RECT 844.2000 800.7000 845.4000 809.7000 ;
	    RECT 858.6000 806.7000 859.8000 809.7000 ;
	    RECT 858.6000 805.5000 859.8000 805.8000 ;
	    RECT 858.6000 803.4000 859.8000 804.6000 ;
	    RECT 861.0000 802.5000 862.2000 809.7000 ;
	    RECT 881.1000 804.6000 882.3000 809.7000 ;
	    RECT 881.1000 803.7000 883.8000 804.6000 ;
	    RECT 885.0000 803.7000 886.2000 809.7000 ;
	    RECT 1019.4000 806.7000 1020.6000 809.7000 ;
	    RECT 1021.8000 804.0000 1023.0000 809.7000 ;
	    RECT 861.0000 801.4500 862.2000 801.6000 ;
	    RECT 863.4000 801.4500 864.6000 801.6000 ;
	    RECT 837.3000 800.4000 839.7000 800.7000 ;
	    RECT 861.0000 800.5500 864.6000 801.4500 ;
	    RECT 861.0000 800.4000 862.2000 800.5500 ;
	    RECT 863.4000 800.4000 864.6000 800.5500 ;
	    RECT 676.2000 798.4500 677.4000 798.6000 ;
	    RECT 683.4000 798.4500 684.6000 798.6000 ;
	    RECT 676.2000 797.5500 684.6000 798.4500 ;
	    RECT 676.2000 797.4000 677.4000 797.5500 ;
	    RECT 683.4000 797.4000 684.6000 797.5500 ;
	    RECT 577.8000 794.1000 579.0000 794.4000 ;
	    RECT 570.9000 793.5000 579.0000 794.1000 ;
	    RECT 569.7000 793.2000 579.0000 793.5000 ;
	    RECT 580.5000 793.5000 593.4000 794.4000 ;
	    RECT 565.8000 792.0000 568.2000 793.2000 ;
	    RECT 569.7000 792.3000 571.8000 793.2000 ;
	    RECT 580.5000 792.3000 581.4000 793.5000 ;
	    RECT 592.2000 793.2000 593.4000 793.5000 ;
	    RECT 597.0000 793.5000 610.5000 794.4000 ;
	    RECT 611.4000 795.0000 612.9000 796.2000 ;
	    RECT 611.4000 793.5000 612.6000 795.0000 ;
	    RECT 597.0000 793.2000 598.2000 793.5000 ;
	    RECT 567.3000 791.4000 568.2000 792.0000 ;
	    RECT 572.7000 791.4000 581.4000 792.3000 ;
	    RECT 582.3000 791.4000 586.2000 792.6000 ;
	    RECT 563.4000 790.2000 566.4000 791.1000 ;
	    RECT 567.3000 790.2000 573.6000 791.4000 ;
	    RECT 565.5000 789.3000 566.4000 790.2000 ;
	    RECT 563.4000 783.3000 564.6000 789.3000 ;
	    RECT 565.5000 788.4000 567.0000 789.3000 ;
	    RECT 565.8000 783.3000 567.0000 788.4000 ;
	    RECT 568.2000 782.4000 569.4000 789.3000 ;
	    RECT 570.6000 783.3000 571.8000 790.2000 ;
	    RECT 573.0000 783.3000 574.2000 789.3000 ;
	    RECT 575.4000 783.3000 576.6000 787.5000 ;
	    RECT 577.8000 783.3000 579.0000 787.5000 ;
	    RECT 580.2000 783.3000 581.4000 790.5000 ;
	    RECT 582.6000 783.3000 583.8000 789.3000 ;
	    RECT 585.0000 783.3000 586.2000 790.5000 ;
	    RECT 587.4000 783.3000 588.6000 789.3000 ;
	    RECT 589.8000 783.3000 591.0000 792.6000 ;
	    RECT 601.8000 791.4000 605.7000 792.6000 ;
	    RECT 594.6000 790.2000 600.9000 791.4000 ;
	    RECT 592.2000 783.3000 593.4000 787.5000 ;
	    RECT 594.6000 783.3000 595.8000 787.5000 ;
	    RECT 597.0000 783.3000 598.2000 787.5000 ;
	    RECT 599.4000 783.3000 600.6000 789.3000 ;
	    RECT 601.8000 783.3000 603.0000 791.4000 ;
	    RECT 609.6000 791.1000 610.5000 793.5000 ;
	    RECT 611.4000 791.4000 612.6000 792.6000 ;
	    RECT 606.6000 790.2000 610.5000 791.1000 ;
	    RECT 604.2000 783.3000 605.4000 789.3000 ;
	    RECT 606.6000 783.3000 607.8000 790.2000 ;
	    RECT 609.0000 783.3000 610.2000 789.3000 ;
	    RECT 611.4000 783.3000 612.6000 790.5000 ;
	    RECT 613.8000 783.3000 615.0000 789.3000 ;
	    RECT 633.0000 783.3000 634.2000 789.3000 ;
	    RECT 635.4000 783.3000 636.6000 796.5000 ;
	    RECT 671.7000 795.6000 675.3000 796.5000 ;
	    RECT 637.8000 794.4000 639.0000 795.6000 ;
	    RECT 637.8000 793.2000 639.0000 793.5000 ;
	    RECT 671.7000 789.3000 672.6000 795.6000 ;
	    RECT 676.5000 795.3000 677.4000 796.5000 ;
	    RECT 637.8000 783.3000 639.0000 789.3000 ;
	    RECT 669.0000 783.3000 670.2000 789.3000 ;
	    RECT 671.4000 783.3000 672.6000 789.3000 ;
	    RECT 673.8000 783.3000 675.0000 794.7000 ;
	    RECT 676.2000 783.3000 677.4000 795.3000 ;
	    RECT 690.6000 783.3000 691.8000 789.3000 ;
	    RECT 693.0000 783.3000 694.2000 799.5000 ;
	    RECT 714.6000 798.4500 715.8000 798.6000 ;
	    RECT 733.8000 798.4500 735.0000 798.6000 ;
	    RECT 714.6000 797.5500 735.0000 798.4500 ;
	    RECT 714.6000 797.4000 715.8000 797.5500 ;
	    RECT 733.8000 797.4000 735.0000 797.5500 ;
	    RECT 738.6000 797.4000 739.8000 798.6000 ;
	    RECT 750.6000 798.4500 751.8000 798.6000 ;
	    RECT 760.2000 798.4500 761.4000 798.6000 ;
	    RECT 750.6000 797.5500 761.4000 798.4500 ;
	    RECT 750.6000 797.4000 751.8000 797.5500 ;
	    RECT 760.2000 797.4000 761.4000 797.5500 ;
	    RECT 712.2000 783.3000 713.4000 789.3000 ;
	    RECT 714.6000 783.3000 715.8000 796.5000 ;
	    RECT 717.0000 795.4500 718.2000 795.6000 ;
	    RECT 736.2000 795.4500 737.4000 795.6000 ;
	    RECT 717.0000 794.5500 737.4000 795.4500 ;
	    RECT 717.0000 794.4000 718.2000 794.5500 ;
	    RECT 736.2000 794.4000 737.4000 794.5500 ;
	    RECT 717.0000 793.2000 718.2000 793.5000 ;
	    RECT 717.0000 783.3000 718.2000 789.3000 ;
	    RECT 736.2000 783.3000 737.4000 789.3000 ;
	    RECT 738.6000 783.3000 739.8000 796.5000 ;
	    RECT 760.2000 796.2000 761.4000 796.5000 ;
	    RECT 741.0000 794.4000 742.2000 795.6000 ;
	    RECT 762.6000 795.3000 763.5000 799.5000 ;
	    RECT 784.2000 798.4500 785.4000 798.6000 ;
	    RECT 786.6000 798.4500 787.8000 798.6000 ;
	    RECT 784.2000 797.5500 787.8000 798.4500 ;
	    RECT 784.2000 797.4000 785.4000 797.5500 ;
	    RECT 786.6000 797.4000 787.8000 797.5500 ;
	    RECT 808.2000 797.4000 809.4000 798.6000 ;
	    RECT 761.1000 794.1000 763.8000 795.3000 ;
	    RECT 741.0000 793.2000 742.2000 793.5000 ;
	    RECT 741.0000 783.3000 742.2000 789.3000 ;
	    RECT 748.2000 786.4500 749.4000 786.6000 ;
	    RECT 753.0000 786.4500 754.2000 786.6000 ;
	    RECT 748.2000 785.5500 754.2000 786.4500 ;
	    RECT 748.2000 785.4000 749.4000 785.5500 ;
	    RECT 753.0000 785.4000 754.2000 785.5500 ;
	    RECT 761.1000 783.3000 762.3000 794.1000 ;
	    RECT 765.0000 783.3000 766.2000 795.3000 ;
	    RECT 784.2000 794.4000 785.4000 795.6000 ;
	    RECT 784.2000 793.2000 785.4000 793.5000 ;
	    RECT 784.2000 783.3000 785.4000 789.3000 ;
	    RECT 786.6000 783.3000 787.8000 796.5000 ;
	    RECT 808.2000 796.2000 809.4000 796.5000 ;
	    RECT 810.6000 795.3000 811.5000 799.5000 ;
	    RECT 837.3000 796.5000 838.2000 800.4000 ;
	    RECT 882.6000 799.5000 883.8000 803.7000 ;
	    RECT 1021.5000 802.8000 1023.0000 804.0000 ;
	    RECT 885.0000 802.5000 886.2000 802.8000 ;
	    RECT 885.0000 800.4000 886.2000 801.6000 ;
	    RECT 887.4000 801.4500 888.6000 801.6000 ;
	    RECT 966.6000 801.4500 967.8000 801.6000 ;
	    RECT 887.4000 800.5500 967.8000 801.4500 ;
	    RECT 887.4000 800.4000 888.6000 800.5500 ;
	    RECT 966.6000 800.4000 967.8000 800.5500 ;
	    RECT 840.6000 797.4000 840.9000 798.6000 ;
	    RECT 841.8000 797.4000 843.0000 798.6000 ;
	    RECT 844.2000 796.5000 845.4000 796.8000 ;
	    RECT 834.6000 795.4500 835.8000 795.6000 ;
	    RECT 837.0000 795.4500 838.2000 795.6000 ;
	    RECT 809.1000 794.1000 811.8000 795.3000 ;
	    RECT 789.0000 783.3000 790.2000 789.3000 ;
	    RECT 809.1000 783.3000 810.3000 794.1000 ;
	    RECT 813.0000 783.3000 814.2000 795.3000 ;
	    RECT 834.6000 794.5500 838.2000 795.4500 ;
	    RECT 834.6000 794.4000 835.8000 794.5500 ;
	    RECT 837.0000 794.4000 838.2000 794.5500 ;
	    RECT 844.2000 794.4000 845.4000 795.6000 ;
	    RECT 839.4000 793.5000 840.6000 793.8000 ;
	    RECT 837.3000 790.5000 838.2000 793.5000 ;
	    RECT 839.4000 791.4000 840.6000 792.6000 ;
	    RECT 841.8000 792.4500 843.0000 792.6000 ;
	    RECT 853.8000 792.4500 855.0000 792.6000 ;
	    RECT 841.8000 791.5500 855.0000 792.4500 ;
	    RECT 841.8000 791.4000 843.0000 791.5500 ;
	    RECT 853.8000 791.4000 855.0000 791.5500 ;
	    RECT 837.3000 789.6000 842.7000 790.5000 ;
	    RECT 837.3000 789.3000 838.2000 789.6000 ;
	    RECT 837.0000 783.3000 838.2000 789.3000 ;
	    RECT 841.8000 789.3000 842.7000 789.6000 ;
	    RECT 839.4000 783.3000 840.6000 788.7000 ;
	    RECT 841.8000 783.3000 843.0000 789.3000 ;
	    RECT 844.2000 783.3000 845.4000 789.3000 ;
	    RECT 858.6000 783.3000 859.8000 789.3000 ;
	    RECT 861.0000 783.3000 862.2000 799.5000 ;
	    RECT 882.6000 798.4500 883.8000 798.6000 ;
	    RECT 940.2000 798.4500 941.4000 798.6000 ;
	    RECT 882.6000 797.5500 941.4000 798.4500 ;
	    RECT 882.6000 797.4000 883.8000 797.5500 ;
	    RECT 940.2000 797.4000 941.4000 797.5500 ;
	    RECT 880.2000 794.4000 881.4000 795.6000 ;
	    RECT 880.2000 793.2000 881.4000 793.5000 ;
	    RECT 880.2000 783.3000 881.4000 789.3000 ;
	    RECT 882.6000 783.3000 883.8000 796.5000 ;
	    RECT 1021.5000 796.2000 1022.7000 802.8000 ;
	    RECT 1024.2001 801.9000 1025.4000 809.7000 ;
	    RECT 1029.0000 803.7000 1030.2001 809.7000 ;
	    RECT 1033.8000 804.9000 1035.0000 809.7000 ;
	    RECT 1036.2001 805.5000 1037.4000 809.7000 ;
	    RECT 1038.6000 805.5000 1039.8000 809.7000 ;
	    RECT 1041.0000 805.5000 1042.2001 809.7000 ;
	    RECT 1043.4000 805.5000 1044.6000 809.7000 ;
	    RECT 1045.8000 806.7000 1047.0000 809.7000 ;
	    RECT 1048.2001 805.5000 1049.4000 809.7000 ;
	    RECT 1050.6000 806.7000 1051.8000 809.7000 ;
	    RECT 1053.0000 805.5000 1054.2001 809.7000 ;
	    RECT 1055.4000 805.5000 1056.6000 809.7000 ;
	    RECT 1057.8000 805.5000 1059.0000 809.7000 ;
	    RECT 1031.4000 803.7000 1035.0000 804.9000 ;
	    RECT 1060.2001 804.9000 1061.4000 809.7000 ;
	    RECT 1031.4000 802.8000 1032.6000 803.7000 ;
	    RECT 1023.6000 801.0000 1025.4000 801.9000 ;
	    RECT 1029.9000 801.9000 1032.6000 802.8000 ;
	    RECT 1038.6000 803.4000 1040.1000 804.6000 ;
	    RECT 1044.6000 803.4000 1044.9000 804.6000 ;
	    RECT 1045.8000 803.4000 1047.0000 804.6000 ;
	    RECT 1048.2001 803.7000 1055.1000 804.6000 ;
	    RECT 1060.2001 803.7000 1064.1000 804.9000 ;
	    RECT 1065.0000 803.7000 1066.2001 809.7000 ;
	    RECT 1048.2001 803.4000 1049.4000 803.7000 ;
	    RECT 1023.6000 798.0000 1024.5000 801.0000 ;
	    RECT 1029.9000 800.1000 1031.1000 801.9000 ;
	    RECT 1025.4000 798.9000 1031.1000 800.1000 ;
	    RECT 1038.6000 799.2000 1039.8000 803.4000 ;
	    RECT 1050.6000 802.5000 1051.8000 802.8000 ;
	    RECT 1048.2001 802.2000 1049.4000 802.5000 ;
	    RECT 1042.8000 801.3000 1049.4000 802.2000 ;
	    RECT 1042.8000 801.0000 1044.0000 801.3000 ;
	    RECT 1050.6000 800.4000 1051.8000 801.6000 ;
	    RECT 1053.9000 800.1000 1055.1000 803.7000 ;
	    RECT 1062.9000 802.8000 1064.1000 803.7000 ;
	    RECT 1062.9000 801.6000 1067.4000 802.8000 ;
	    RECT 1069.8000 800.7000 1071.0000 809.7000 ;
	    RECT 1089.0000 803.7000 1090.2001 809.7000 ;
	    RECT 1092.9000 804.6000 1094.1000 809.7000 ;
	    RECT 1091.4000 803.7000 1094.1000 804.6000 ;
	    RECT 1113.0000 803.7000 1114.2001 809.7000 ;
	    RECT 1116.9000 804.6000 1118.1000 809.7000 ;
	    RECT 1115.4000 803.7000 1118.1000 804.6000 ;
	    RECT 1151.4000 803.7000 1152.6000 809.7000 ;
	    RECT 1153.8000 804.0000 1155.0000 809.7000 ;
	    RECT 1156.2001 804.9000 1157.4000 809.7000 ;
	    RECT 1158.6000 804.0000 1159.8000 809.7000 ;
	    RECT 1170.6000 806.7000 1171.8000 809.7000 ;
	    RECT 1170.6000 805.5000 1171.8000 805.8000 ;
	    RECT 1153.8000 803.7000 1159.8000 804.0000 ;
	    RECT 1089.0000 802.5000 1090.2001 802.8000 ;
	    RECT 1043.4000 798.9000 1048.2001 800.1000 ;
	    RECT 1053.9000 798.9000 1056.9000 800.1000 ;
	    RECT 1057.8000 799.5000 1071.0000 800.7000 ;
	    RECT 1089.0000 800.4000 1090.2001 801.6000 ;
	    RECT 1091.4000 799.5000 1092.6000 803.7000 ;
	    RECT 1113.0000 802.5000 1114.2001 802.8000 ;
	    RECT 1098.6000 801.4500 1099.8000 801.6000 ;
	    RECT 1113.0000 801.4500 1114.2001 801.6000 ;
	    RECT 1098.6000 800.5500 1114.2001 801.4500 ;
	    RECT 1098.6000 800.4000 1099.8000 800.5500 ;
	    RECT 1113.0000 800.4000 1114.2001 800.5500 ;
	    RECT 1115.4000 799.5000 1116.6000 803.7000 ;
	    RECT 1151.7001 802.5000 1152.6000 803.7000 ;
	    RECT 1154.1000 803.1000 1159.5000 803.7000 ;
	    RECT 1170.6000 803.4000 1171.8000 804.6000 ;
	    RECT 1173.0000 802.5000 1174.2001 809.7000 ;
	    RECT 1151.4000 800.4000 1152.6000 801.6000 ;
	    RECT 1153.5000 800.4000 1155.3000 801.6000 ;
	    RECT 1157.4000 800.7000 1157.7001 802.2000 ;
	    RECT 1158.6000 800.4000 1159.8000 801.6000 ;
	    RECT 1173.0000 801.4500 1174.2001 801.6000 ;
	    RECT 1161.1500 800.5500 1174.2001 801.4500 ;
	    RECT 1033.8000 798.0000 1035.0000 798.9000 ;
	    RECT 1023.6000 797.1000 1024.8000 798.0000 ;
	    RECT 1033.8000 797.1000 1059.3000 798.0000 ;
	    RECT 1060.2001 797.4000 1061.4000 798.6000 ;
	    RECT 1067.7001 798.0000 1068.9000 798.3000 ;
	    RECT 1062.3000 797.1000 1068.9000 798.0000 ;
	    RECT 885.0000 795.4500 886.2000 795.6000 ;
	    RECT 935.4000 795.4500 936.6000 795.6000 ;
	    RECT 885.0000 794.5500 936.6000 795.4500 ;
	    RECT 1021.5000 795.0000 1023.0000 796.2000 ;
	    RECT 885.0000 794.4000 886.2000 794.5500 ;
	    RECT 935.4000 794.4000 936.6000 794.5500 ;
	    RECT 1021.8000 793.5000 1023.0000 795.0000 ;
	    RECT 1023.9000 794.4000 1024.8000 797.1000 ;
	    RECT 1025.7001 796.2000 1026.9000 796.5000 ;
	    RECT 1025.7001 795.3000 1064.1000 796.2000 ;
	    RECT 1059.9000 795.0000 1061.1000 795.3000 ;
	    RECT 1065.0000 794.4000 1066.2001 795.6000 ;
	    RECT 1023.9000 793.5000 1037.4000 794.4000 ;
	    RECT 904.2000 792.4500 905.4000 792.6000 ;
	    RECT 1021.8000 792.4500 1023.0000 792.6000 ;
	    RECT 904.2000 791.5500 1023.0000 792.4500 ;
	    RECT 904.2000 791.4000 905.4000 791.5500 ;
	    RECT 1021.8000 791.4000 1023.0000 791.5500 ;
	    RECT 1023.9000 791.1000 1024.8000 793.5000 ;
	    RECT 1036.2001 793.2000 1037.4000 793.5000 ;
	    RECT 1041.0000 793.5000 1053.9000 794.4000 ;
	    RECT 1041.0000 793.2000 1042.2001 793.5000 ;
	    RECT 1028.7001 791.4000 1032.6000 792.6000 ;
	    RECT 885.0000 783.3000 886.2000 789.3000 ;
	    RECT 1019.4000 783.3000 1020.6000 789.3000 ;
	    RECT 1021.8000 783.3000 1023.0000 790.5000 ;
	    RECT 1023.9000 790.2000 1027.8000 791.1000 ;
	    RECT 1024.2001 783.3000 1025.4000 789.3000 ;
	    RECT 1026.6000 783.3000 1027.8000 790.2000 ;
	    RECT 1029.0000 783.3000 1030.2001 789.3000 ;
	    RECT 1031.4000 783.3000 1032.6000 791.4000 ;
	    RECT 1033.5000 790.2000 1039.8000 791.4000 ;
	    RECT 1033.8000 783.3000 1035.0000 789.3000 ;
	    RECT 1036.2001 783.3000 1037.4000 787.5000 ;
	    RECT 1038.6000 783.3000 1039.8000 787.5000 ;
	    RECT 1041.0000 783.3000 1042.2001 787.5000 ;
	    RECT 1043.4000 783.3000 1044.6000 792.6000 ;
	    RECT 1048.2001 791.4000 1052.1000 792.6000 ;
	    RECT 1053.0000 792.3000 1053.9000 793.5000 ;
	    RECT 1055.4000 794.1000 1056.6000 794.4000 ;
	    RECT 1055.4000 793.5000 1063.5000 794.1000 ;
	    RECT 1055.4000 793.2000 1064.7001 793.5000 ;
	    RECT 1062.6000 792.3000 1064.7001 793.2000 ;
	    RECT 1053.0000 791.4000 1061.7001 792.3000 ;
	    RECT 1066.2001 792.0000 1068.6000 793.2000 ;
	    RECT 1066.2001 791.4000 1067.1000 792.0000 ;
	    RECT 1045.8000 783.3000 1047.0000 789.3000 ;
	    RECT 1048.2001 783.3000 1049.4000 790.5000 ;
	    RECT 1050.6000 783.3000 1051.8000 789.3000 ;
	    RECT 1053.0000 783.3000 1054.2001 790.5000 ;
	    RECT 1060.8000 790.2000 1067.1000 791.4000 ;
	    RECT 1069.8000 791.1000 1071.0000 799.5000 ;
	    RECT 1072.2001 798.4500 1073.4000 798.6000 ;
	    RECT 1091.4000 798.4500 1092.6000 798.6000 ;
	    RECT 1072.2001 797.5500 1092.6000 798.4500 ;
	    RECT 1072.2001 797.4000 1073.4000 797.5500 ;
	    RECT 1091.4000 797.4000 1092.6000 797.5500 ;
	    RECT 1103.4000 798.4500 1104.6000 798.6000 ;
	    RECT 1115.4000 798.4500 1116.6000 798.6000 ;
	    RECT 1103.4000 797.5500 1116.6000 798.4500 ;
	    RECT 1103.4000 797.4000 1104.6000 797.5500 ;
	    RECT 1115.4000 797.4000 1116.6000 797.5500 ;
	    RECT 1068.0000 790.2000 1071.0000 791.1000 ;
	    RECT 1055.4000 783.3000 1056.6000 787.5000 ;
	    RECT 1057.8000 783.3000 1059.0000 787.5000 ;
	    RECT 1060.2001 783.3000 1061.4000 789.3000 ;
	    RECT 1062.6000 783.3000 1063.8000 790.2000 ;
	    RECT 1068.0000 789.3000 1068.9000 790.2000 ;
	    RECT 1065.0000 782.4000 1066.2001 789.3000 ;
	    RECT 1067.4000 788.4000 1068.9000 789.3000 ;
	    RECT 1067.4000 783.3000 1068.6000 788.4000 ;
	    RECT 1069.8000 783.3000 1071.0000 789.3000 ;
	    RECT 1089.0000 783.3000 1090.2001 789.3000 ;
	    RECT 1091.4000 783.3000 1092.6000 796.5000 ;
	    RECT 1093.8000 794.4000 1095.0000 795.6000 ;
	    RECT 1093.8000 793.2000 1095.0000 793.5000 ;
	    RECT 1093.8000 783.3000 1095.0000 789.3000 ;
	    RECT 1113.0000 783.3000 1114.2001 789.3000 ;
	    RECT 1115.4000 783.3000 1116.6000 796.5000 ;
	    RECT 1117.8000 794.4000 1119.0000 795.6000 ;
	    RECT 1144.2001 795.4500 1145.4000 795.6000 ;
	    RECT 1151.4000 795.4500 1152.6000 795.6000 ;
	    RECT 1144.2001 794.5500 1152.6000 795.4500 ;
	    RECT 1144.2001 794.4000 1145.4000 794.5500 ;
	    RECT 1151.4000 794.4000 1152.6000 794.5500 ;
	    RECT 1154.4000 795.3000 1155.3000 800.4000 ;
	    RECT 1156.2001 799.5000 1157.4000 799.8000 ;
	    RECT 1156.2001 798.4500 1157.4000 798.6000 ;
	    RECT 1161.1500 798.4500 1162.0500 800.5500 ;
	    RECT 1173.0000 800.4000 1174.2001 800.5500 ;
	    RECT 1300.2001 800.7000 1301.4000 809.7000 ;
	    RECT 1305.0000 803.7000 1306.2001 809.7000 ;
	    RECT 1309.8000 804.9000 1311.0000 809.7000 ;
	    RECT 1312.2001 805.5000 1313.4000 809.7000 ;
	    RECT 1314.6000 805.5000 1315.8000 809.7000 ;
	    RECT 1317.0000 805.5000 1318.2001 809.7000 ;
	    RECT 1319.4000 806.7000 1320.6000 809.7000 ;
	    RECT 1321.8000 805.5000 1323.0000 809.7000 ;
	    RECT 1324.2001 806.7000 1325.4000 809.7000 ;
	    RECT 1326.6000 805.5000 1327.8000 809.7000 ;
	    RECT 1329.0000 805.5000 1330.2001 809.7000 ;
	    RECT 1331.4000 805.5000 1332.6000 809.7000 ;
	    RECT 1333.8000 805.5000 1335.0000 809.7000 ;
	    RECT 1307.1000 803.7000 1311.0000 804.9000 ;
	    RECT 1336.2001 804.9000 1337.4000 809.7000 ;
	    RECT 1316.1000 803.7000 1323.0000 804.6000 ;
	    RECT 1307.1000 802.8000 1308.3000 803.7000 ;
	    RECT 1303.8000 801.6000 1308.3000 802.8000 ;
	    RECT 1300.2001 799.5000 1313.4000 800.7000 ;
	    RECT 1316.1000 800.1000 1317.3000 803.7000 ;
	    RECT 1321.8000 803.4000 1323.0000 803.7000 ;
	    RECT 1324.2001 803.4000 1325.4000 804.6000 ;
	    RECT 1326.3000 803.4000 1326.6000 804.6000 ;
	    RECT 1331.1000 803.4000 1332.6000 804.6000 ;
	    RECT 1336.2001 803.7000 1339.8000 804.9000 ;
	    RECT 1341.0000 803.7000 1342.2001 809.7000 ;
	    RECT 1319.4000 802.5000 1320.6000 802.8000 ;
	    RECT 1321.8000 802.2000 1323.0000 802.5000 ;
	    RECT 1319.4000 800.4000 1320.6000 801.6000 ;
	    RECT 1321.8000 801.3000 1328.4000 802.2000 ;
	    RECT 1327.2001 801.0000 1328.4000 801.3000 ;
	    RECT 1156.2001 797.5500 1162.0500 798.4500 ;
	    RECT 1156.2001 797.4000 1157.4000 797.5500 ;
	    RECT 1154.4000 794.4000 1155.9000 795.3000 ;
	    RECT 1117.8000 793.2000 1119.0000 793.5000 ;
	    RECT 1152.6000 792.6000 1153.5000 793.5000 ;
	    RECT 1152.6000 791.4000 1153.8000 792.6000 ;
	    RECT 1117.8000 783.3000 1119.0000 789.3000 ;
	    RECT 1152.3000 783.3000 1153.5000 789.3000 ;
	    RECT 1154.7001 783.3000 1155.9000 794.4000 ;
	    RECT 1158.6000 783.3000 1159.8000 795.3000 ;
	    RECT 1170.6000 783.3000 1171.8000 789.3000 ;
	    RECT 1173.0000 783.3000 1174.2001 799.5000 ;
	    RECT 1300.2001 791.1000 1301.4000 799.5000 ;
	    RECT 1314.3000 798.9000 1317.3000 800.1000 ;
	    RECT 1323.0000 798.9000 1327.8000 800.1000 ;
	    RECT 1331.4000 799.2000 1332.6000 803.4000 ;
	    RECT 1338.6000 802.8000 1339.8000 803.7000 ;
	    RECT 1338.6000 801.9000 1341.3000 802.8000 ;
	    RECT 1340.1000 800.1000 1341.3000 801.9000 ;
	    RECT 1345.8000 801.9000 1347.0000 809.7000 ;
	    RECT 1348.2001 804.0000 1349.4000 809.7000 ;
	    RECT 1350.6000 806.7000 1351.8000 809.7000 ;
	    RECT 1348.2001 802.8000 1349.7001 804.0000 ;
	    RECT 1398.6000 803.7000 1399.8000 809.7000 ;
	    RECT 1401.0000 804.6000 1402.5000 809.7000 ;
	    RECT 1405.2001 804.3000 1407.6000 809.7000 ;
	    RECT 1410.3000 804.6000 1411.8000 809.7000 ;
	    RECT 1398.6000 802.8000 1402.5000 803.7000 ;
	    RECT 1345.8000 801.0000 1347.6000 801.9000 ;
	    RECT 1340.1000 798.9000 1345.8000 800.1000 ;
	    RECT 1302.3000 798.0000 1303.5000 798.3000 ;
	    RECT 1302.3000 797.1000 1308.9000 798.0000 ;
	    RECT 1309.8000 797.4000 1311.0000 798.6000 ;
	    RECT 1336.2001 798.0000 1337.4000 798.9000 ;
	    RECT 1346.7001 798.0000 1347.6000 801.0000 ;
	    RECT 1311.9000 797.1000 1337.4000 798.0000 ;
	    RECT 1346.4000 797.1000 1347.6000 798.0000 ;
	    RECT 1344.3000 796.2000 1345.5000 796.5000 ;
	    RECT 1305.0000 794.4000 1306.2001 795.6000 ;
	    RECT 1307.1000 795.3000 1345.5000 796.2000 ;
	    RECT 1310.1000 795.0000 1311.3000 795.3000 ;
	    RECT 1346.4000 794.4000 1347.3000 797.1000 ;
	    RECT 1348.5000 796.2000 1349.7001 802.8000 ;
	    RECT 1401.3000 802.5000 1402.5000 802.8000 ;
	    RECT 1403.4000 802.2000 1405.8000 803.4000 ;
	    RECT 1377.0000 801.4500 1378.2001 801.6000 ;
	    RECT 1398.6000 801.4500 1399.8000 801.6000 ;
	    RECT 1377.0000 800.5500 1399.8000 801.4500 ;
	    RECT 1377.0000 800.4000 1378.2001 800.5500 ;
	    RECT 1398.6000 800.4000 1399.8000 800.5500 ;
	    RECT 1400.7001 801.3000 1401.0000 801.6000 ;
	    RECT 1406.7001 801.3000 1407.6000 804.3000 ;
	    RECT 1413.0000 803.7000 1414.2001 809.7000 ;
	    RECT 1408.5000 802.2000 1409.7001 803.4000 ;
	    RECT 1410.6000 802.8000 1414.2001 803.7000 ;
	    RECT 1410.6000 802.5000 1411.8000 802.8000 ;
	    RECT 1425.0000 802.5000 1426.2001 809.7000 ;
	    RECT 1427.4000 806.7000 1428.6000 809.7000 ;
	    RECT 1427.4000 805.5000 1428.6000 805.8000 ;
	    RECT 1427.4000 803.4000 1428.6000 804.6000 ;
	    RECT 1400.7001 801.0000 1401.9000 801.3000 ;
	    RECT 1400.7001 800.4000 1405.2001 801.0000 ;
	    RECT 1401.0000 800.1000 1405.2001 800.4000 ;
	    RECT 1404.0000 799.8000 1405.2001 800.1000 ;
	    RECT 1406.1000 800.4000 1407.6000 801.3000 ;
	    RECT 1408.8000 801.6000 1409.7001 802.2000 ;
	    RECT 1408.8000 800.4000 1410.0000 801.6000 ;
	    RECT 1411.8000 800.4000 1412.1000 801.6000 ;
	    RECT 1413.0000 800.4000 1414.2001 801.6000 ;
	    RECT 1415.4000 801.4500 1416.6000 801.6000 ;
	    RECT 1417.8000 801.4500 1419.0000 801.6000 ;
	    RECT 1425.0000 801.4500 1426.2001 801.6000 ;
	    RECT 1415.4000 800.5500 1426.2001 801.4500 ;
	    RECT 1455.6000 801.3000 1456.8000 809.7000 ;
	    RECT 1415.4000 800.4000 1416.6000 800.5500 ;
	    RECT 1417.8000 800.4000 1419.0000 800.5500 ;
	    RECT 1425.0000 800.4000 1426.2001 800.5500 ;
	    RECT 1454.1000 800.7000 1456.8000 801.3000 ;
	    RECT 1461.0000 800.7000 1462.2001 809.7000 ;
	    RECT 1463.4000 807.4500 1464.6000 807.6000 ;
	    RECT 1475.4000 807.4500 1476.6000 807.6000 ;
	    RECT 1463.4000 806.5500 1476.6000 807.4500 ;
	    RECT 1487.4000 806.7000 1488.6000 809.7000 ;
	    RECT 1463.4000 806.4000 1464.6000 806.5500 ;
	    RECT 1475.4000 806.4000 1476.6000 806.5500 ;
	    RECT 1487.7001 805.5000 1488.9000 805.8000 ;
	    RECT 1463.4000 804.4500 1464.6000 804.6000 ;
	    RECT 1487.4000 804.4500 1488.6000 804.6000 ;
	    RECT 1463.4000 803.5500 1488.6000 804.4500 ;
	    RECT 1489.8000 803.7000 1491.0000 809.7000 ;
	    RECT 1493.7001 803.7000 1494.9000 809.7000 ;
	    RECT 1523.4000 804.0000 1524.6000 809.7000 ;
	    RECT 1525.8000 804.9000 1527.0000 809.7000 ;
	    RECT 1528.2001 808.8000 1534.2001 809.7000 ;
	    RECT 1528.2001 804.0000 1529.4000 808.8000 ;
	    RECT 1523.4000 803.7000 1529.4000 804.0000 ;
	    RECT 1530.6000 803.7000 1531.8000 807.9000 ;
	    RECT 1533.0000 803.7000 1534.2001 808.8000 ;
	    RECT 1463.4000 803.4000 1464.6000 803.5500 ;
	    RECT 1487.4000 803.4000 1488.6000 803.5500 ;
	    RECT 1454.1000 800.4000 1456.5000 800.7000 ;
	    RECT 1406.1000 799.5000 1407.0000 800.4000 ;
	    RECT 1401.9000 798.3000 1403.1000 798.6000 ;
	    RECT 1401.9000 797.4000 1404.3000 798.3000 ;
	    RECT 1405.8000 797.4000 1407.0000 798.6000 ;
	    RECT 1403.1000 797.1000 1404.3000 797.4000 ;
	    RECT 1314.6000 794.1000 1315.8000 794.4000 ;
	    RECT 1307.7001 793.5000 1315.8000 794.1000 ;
	    RECT 1306.5000 793.2000 1315.8000 793.5000 ;
	    RECT 1317.3000 793.5000 1330.2001 794.4000 ;
	    RECT 1302.6000 792.0000 1305.0000 793.2000 ;
	    RECT 1306.5000 792.3000 1308.6000 793.2000 ;
	    RECT 1317.3000 792.3000 1318.2001 793.5000 ;
	    RECT 1329.0000 793.2000 1330.2001 793.5000 ;
	    RECT 1333.8000 793.5000 1347.3000 794.4000 ;
	    RECT 1348.2001 795.0000 1349.7001 796.2000 ;
	    RECT 1406.1000 795.3000 1407.0000 796.5000 ;
	    RECT 1348.2001 793.5000 1349.4000 795.0000 ;
	    RECT 1398.6000 794.4000 1402.5000 795.3000 ;
	    RECT 1333.8000 793.2000 1335.0000 793.5000 ;
	    RECT 1304.1000 791.4000 1305.0000 792.0000 ;
	    RECT 1309.5000 791.4000 1318.2001 792.3000 ;
	    RECT 1319.1000 791.4000 1323.0000 792.6000 ;
	    RECT 1300.2001 790.2000 1303.2001 791.1000 ;
	    RECT 1304.1000 790.2000 1310.4000 791.4000 ;
	    RECT 1302.3000 789.3000 1303.2001 790.2000 ;
	    RECT 1300.2001 783.3000 1301.4000 789.3000 ;
	    RECT 1302.3000 788.4000 1303.8000 789.3000 ;
	    RECT 1302.6000 783.3000 1303.8000 788.4000 ;
	    RECT 1305.0000 782.4000 1306.2001 789.3000 ;
	    RECT 1307.4000 783.3000 1308.6000 790.2000 ;
	    RECT 1309.8000 783.3000 1311.0000 789.3000 ;
	    RECT 1312.2001 783.3000 1313.4000 787.5000 ;
	    RECT 1314.6000 783.3000 1315.8000 787.5000 ;
	    RECT 1317.0000 783.3000 1318.2001 790.5000 ;
	    RECT 1319.4000 783.3000 1320.6000 789.3000 ;
	    RECT 1321.8000 783.3000 1323.0000 790.5000 ;
	    RECT 1324.2001 783.3000 1325.4000 789.3000 ;
	    RECT 1326.6000 783.3000 1327.8000 792.6000 ;
	    RECT 1338.6000 791.4000 1342.5000 792.6000 ;
	    RECT 1331.4000 790.2000 1337.7001 791.4000 ;
	    RECT 1329.0000 783.3000 1330.2001 787.5000 ;
	    RECT 1331.4000 783.3000 1332.6000 787.5000 ;
	    RECT 1333.8000 783.3000 1335.0000 787.5000 ;
	    RECT 1336.2001 783.3000 1337.4000 789.3000 ;
	    RECT 1338.6000 783.3000 1339.8000 791.4000 ;
	    RECT 1346.4000 791.1000 1347.3000 793.5000 ;
	    RECT 1348.2001 791.4000 1349.4000 792.6000 ;
	    RECT 1343.4000 790.2000 1347.3000 791.1000 ;
	    RECT 1341.0000 783.3000 1342.2001 789.3000 ;
	    RECT 1343.4000 783.3000 1344.6000 790.2000 ;
	    RECT 1345.8000 783.3000 1347.0000 789.3000 ;
	    RECT 1348.2001 783.3000 1349.4000 790.5000 ;
	    RECT 1350.6000 783.3000 1351.8000 789.3000 ;
	    RECT 1398.6000 783.3000 1399.8000 794.4000 ;
	    RECT 1401.3000 794.1000 1402.5000 794.4000 ;
	    RECT 1401.0000 783.3000 1402.5000 793.2000 ;
	    RECT 1405.2001 783.3000 1407.6000 795.3000 ;
	    RECT 1410.6000 794.4000 1414.2001 795.3000 ;
	    RECT 1410.6000 794.1000 1411.8000 794.4000 ;
	    RECT 1410.3000 783.3000 1411.8000 793.2000 ;
	    RECT 1413.0000 783.3000 1414.2001 794.4000 ;
	    RECT 1425.0000 783.3000 1426.2001 799.5000 ;
	    RECT 1454.1000 796.5000 1455.0000 800.4000 ;
	    RECT 1457.4000 797.4000 1457.7001 798.6000 ;
	    RECT 1458.6000 797.4000 1459.8000 798.6000 ;
	    RECT 1465.8000 798.4500 1467.0000 798.6000 ;
	    RECT 1487.4000 798.4500 1488.6000 798.6000 ;
	    RECT 1465.8000 797.5500 1488.6000 798.4500 ;
	    RECT 1490.1000 798.3000 1491.0000 803.7000 ;
	    RECT 1523.7001 803.1000 1529.1000 803.7000 ;
	    RECT 1492.2001 800.4000 1493.4000 801.6000 ;
	    RECT 1504.2001 801.4500 1505.4000 801.6000 ;
	    RECT 1523.4000 801.4500 1524.6000 801.6000 ;
	    RECT 1504.2001 800.5500 1524.6000 801.4500 ;
	    RECT 1525.5000 800.7000 1525.8000 802.2000 ;
	    RECT 1530.9000 801.6000 1531.8000 803.7000 ;
	    RECT 1504.2001 800.4000 1505.4000 800.5500 ;
	    RECT 1523.4000 800.4000 1524.6000 800.5500 ;
	    RECT 1528.2001 800.4000 1529.4000 801.6000 ;
	    RECT 1530.3000 800.7000 1531.8000 801.6000 ;
	    RECT 1533.0000 800.4000 1534.2001 801.6000 ;
	    RECT 1558.8000 801.3000 1560.0000 809.7000 ;
	    RECT 1557.3000 800.7000 1560.0000 801.3000 ;
	    RECT 1564.2001 800.7000 1565.4000 809.7000 ;
	    RECT 1557.3000 800.4000 1559.7001 800.7000 ;
	    RECT 1525.8000 799.5000 1527.0000 799.8000 ;
	    RECT 1530.6000 799.5000 1531.8000 799.8000 ;
	    RECT 1492.2001 799.2000 1493.4000 799.5000 ;
	    RECT 1465.8000 797.4000 1467.0000 797.5500 ;
	    RECT 1487.4000 797.4000 1488.6000 797.5500 ;
	    RECT 1489.5000 797.4000 1491.0000 798.3000 ;
	    RECT 1493.4000 796.8000 1493.7001 798.3000 ;
	    RECT 1494.6000 797.4000 1495.8000 798.6000 ;
	    RECT 1525.8000 797.4000 1527.0000 798.6000 ;
	    RECT 1461.0000 796.5000 1462.2001 796.8000 ;
	    RECT 1427.4000 795.4500 1428.6000 795.6000 ;
	    RECT 1437.0000 795.4500 1438.2001 795.6000 ;
	    RECT 1453.8000 795.4500 1455.0000 795.6000 ;
	    RECT 1427.4000 794.5500 1455.0000 795.4500 ;
	    RECT 1427.4000 794.4000 1428.6000 794.5500 ;
	    RECT 1437.0000 794.4000 1438.2001 794.5500 ;
	    RECT 1453.8000 794.4000 1455.0000 794.5500 ;
	    RECT 1461.0000 795.4500 1462.2001 795.6000 ;
	    RECT 1463.4000 795.4500 1464.6000 795.6000 ;
	    RECT 1461.0000 794.5500 1464.6000 795.4500 ;
	    RECT 1487.7001 795.3000 1488.6000 796.5000 ;
	    RECT 1528.2001 795.3000 1529.1000 799.5000 ;
	    RECT 1533.0000 799.2000 1534.2001 799.5000 ;
	    RECT 1530.6000 797.4000 1531.8000 798.6000 ;
	    RECT 1557.3000 796.5000 1558.2001 800.4000 ;
	    RECT 1560.6000 797.4000 1560.9000 798.6000 ;
	    RECT 1561.8000 797.4000 1563.0000 798.6000 ;
	    RECT 1564.2001 796.5000 1565.4000 796.8000 ;
	    RECT 1535.4000 795.4500 1536.6000 795.6000 ;
	    RECT 1557.0000 795.4500 1558.2001 795.6000 ;
	    RECT 1461.0000 794.4000 1462.2001 794.5500 ;
	    RECT 1463.4000 794.4000 1464.6000 794.5500 ;
	    RECT 1456.2001 793.5000 1457.4000 793.8000 ;
	    RECT 1454.1000 790.5000 1455.0000 793.5000 ;
	    RECT 1456.2001 791.4000 1457.4000 792.6000 ;
	    RECT 1454.1000 789.6000 1459.5000 790.5000 ;
	    RECT 1454.1000 789.3000 1455.0000 789.6000 ;
	    RECT 1427.4000 783.3000 1428.6000 789.3000 ;
	    RECT 1453.8000 783.3000 1455.0000 789.3000 ;
	    RECT 1458.6000 789.3000 1459.5000 789.6000 ;
	    RECT 1456.2001 783.3000 1457.4000 788.7000 ;
	    RECT 1458.6000 783.3000 1459.8000 789.3000 ;
	    RECT 1461.0000 783.3000 1462.2001 789.3000 ;
	    RECT 1487.4000 783.3000 1488.6000 795.3000 ;
	    RECT 1489.8000 794.4000 1495.8000 795.3000 ;
	    RECT 1489.8000 783.3000 1491.0000 794.4000 ;
	    RECT 1492.2001 783.3000 1493.4000 793.5000 ;
	    RECT 1494.6000 783.3000 1495.8000 794.4000 ;
	    RECT 1523.4000 783.3000 1524.6000 795.3000 ;
	    RECT 1527.3000 783.3000 1530.3000 795.3000 ;
	    RECT 1533.0000 783.3000 1534.2001 795.3000 ;
	    RECT 1535.4000 794.5500 1558.2001 795.4500 ;
	    RECT 1535.4000 794.4000 1536.6000 794.5500 ;
	    RECT 1557.0000 794.4000 1558.2001 794.5500 ;
	    RECT 1564.2001 794.4000 1565.4000 795.6000 ;
	    RECT 1559.4000 793.5000 1560.6000 793.8000 ;
	    RECT 1557.3000 790.5000 1558.2001 793.5000 ;
	    RECT 1559.4000 791.4000 1560.6000 792.6000 ;
	    RECT 1557.3000 789.6000 1562.7001 790.5000 ;
	    RECT 1557.3000 789.3000 1558.2001 789.6000 ;
	    RECT 1557.0000 783.3000 1558.2001 789.3000 ;
	    RECT 1561.8000 789.3000 1562.7001 789.6000 ;
	    RECT 1559.4000 783.3000 1560.6000 788.7000 ;
	    RECT 1561.8000 783.3000 1563.0000 789.3000 ;
	    RECT 1564.2001 783.3000 1565.4000 789.3000 ;
	    RECT 1.2000 780.6000 1569.0000 782.4000 ;
	    RECT 124.2000 773.7000 125.4000 779.7000 ;
	    RECT 126.6000 772.5000 127.8000 779.7000 ;
	    RECT 129.0000 773.7000 130.2000 779.7000 ;
	    RECT 131.4000 772.8000 132.6000 779.7000 ;
	    RECT 133.8000 773.7000 135.0000 779.7000 ;
	    RECT 128.7000 771.9000 132.6000 772.8000 ;
	    RECT 124.2000 771.4500 125.4000 771.6000 ;
	    RECT 126.6000 771.4500 127.8000 771.6000 ;
	    RECT 124.2000 770.5500 127.8000 771.4500 ;
	    RECT 124.2000 770.4000 125.4000 770.5500 ;
	    RECT 126.6000 770.4000 127.8000 770.5500 ;
	    RECT 128.7000 769.5000 129.6000 771.9000 ;
	    RECT 136.2000 771.6000 137.4000 779.7000 ;
	    RECT 138.6000 773.7000 139.8000 779.7000 ;
	    RECT 141.0000 775.5000 142.2000 779.7000 ;
	    RECT 143.4000 775.5000 144.6000 779.7000 ;
	    RECT 145.8000 775.5000 147.0000 779.7000 ;
	    RECT 138.3000 771.6000 144.6000 772.8000 ;
	    RECT 133.5000 770.4000 137.4000 771.6000 ;
	    RECT 148.2000 770.4000 149.4000 779.7000 ;
	    RECT 150.6000 773.7000 151.8000 779.7000 ;
	    RECT 153.0000 772.5000 154.2000 779.7000 ;
	    RECT 155.4000 773.7000 156.6000 779.7000 ;
	    RECT 157.8000 772.5000 159.0000 779.7000 ;
	    RECT 160.2000 775.5000 161.4000 779.7000 ;
	    RECT 162.6000 775.5000 163.8000 779.7000 ;
	    RECT 165.0000 773.7000 166.2000 779.7000 ;
	    RECT 167.4000 772.8000 168.6000 779.7000 ;
	    RECT 169.8000 773.7000 171.0000 780.6000 ;
	    RECT 172.2000 774.6000 173.4000 779.7000 ;
	    RECT 172.2000 773.7000 173.7000 774.6000 ;
	    RECT 174.6000 773.7000 175.8000 779.7000 ;
	    RECT 189.0000 773.7000 190.2000 779.7000 ;
	    RECT 172.8000 772.8000 173.7000 773.7000 ;
	    RECT 165.6000 771.6000 171.9000 772.8000 ;
	    RECT 172.8000 771.9000 175.8000 772.8000 ;
	    RECT 153.0000 770.4000 156.9000 771.6000 ;
	    RECT 157.8000 770.7000 166.5000 771.6000 ;
	    RECT 171.0000 771.0000 171.9000 771.6000 ;
	    RECT 141.0000 769.5000 142.2000 769.8000 ;
	    RECT 126.6000 768.0000 127.8000 769.5000 ;
	    RECT 126.3000 766.8000 127.8000 768.0000 ;
	    RECT 128.7000 768.6000 142.2000 769.5000 ;
	    RECT 145.8000 769.5000 147.0000 769.8000 ;
	    RECT 157.8000 769.5000 158.7000 770.7000 ;
	    RECT 167.4000 769.8000 169.5000 770.7000 ;
	    RECT 171.0000 769.8000 173.4000 771.0000 ;
	    RECT 145.8000 768.6000 158.7000 769.5000 ;
	    RECT 160.2000 769.5000 169.5000 769.8000 ;
	    RECT 160.2000 768.9000 168.3000 769.5000 ;
	    RECT 160.2000 768.6000 161.4000 768.9000 ;
	    RECT 49.8000 762.4500 51.0000 762.6000 ;
	    RECT 105.0000 762.4500 106.2000 762.6000 ;
	    RECT 49.8000 761.5500 106.2000 762.4500 ;
	    RECT 49.8000 761.4000 51.0000 761.5500 ;
	    RECT 105.0000 761.4000 106.2000 761.5500 ;
	    RECT 126.3000 760.2000 127.5000 766.8000 ;
	    RECT 128.7000 765.9000 129.6000 768.6000 ;
	    RECT 164.7000 767.7000 165.9000 768.0000 ;
	    RECT 130.5000 766.8000 168.9000 767.7000 ;
	    RECT 169.8000 767.4000 171.0000 768.6000 ;
	    RECT 130.5000 766.5000 131.7000 766.8000 ;
	    RECT 128.4000 765.0000 129.6000 765.9000 ;
	    RECT 138.6000 765.0000 164.1000 765.9000 ;
	    RECT 128.4000 762.0000 129.3000 765.0000 ;
	    RECT 138.6000 764.1000 139.8000 765.0000 ;
	    RECT 165.0000 764.4000 166.2000 765.6000 ;
	    RECT 167.1000 765.0000 173.7000 765.9000 ;
	    RECT 172.5000 764.7000 173.7000 765.0000 ;
	    RECT 130.2000 762.9000 135.9000 764.1000 ;
	    RECT 128.4000 761.1000 130.2000 762.0000 ;
	    RECT 126.3000 759.0000 127.8000 760.2000 ;
	    RECT 124.2000 753.3000 125.4000 756.3000 ;
	    RECT 126.6000 753.3000 127.8000 759.0000 ;
	    RECT 129.0000 753.3000 130.2000 761.1000 ;
	    RECT 134.7000 761.1000 135.9000 762.9000 ;
	    RECT 134.7000 760.2000 137.4000 761.1000 ;
	    RECT 136.2000 759.3000 137.4000 760.2000 ;
	    RECT 143.4000 759.6000 144.6000 763.8000 ;
	    RECT 148.2000 762.9000 153.0000 764.1000 ;
	    RECT 158.7000 762.9000 161.7000 764.1000 ;
	    RECT 174.6000 763.5000 175.8000 771.9000 ;
	    RECT 191.4000 763.5000 192.6000 779.7000 ;
	    RECT 229.8000 767.7000 231.0000 779.7000 ;
	    RECT 233.7000 767.7000 236.7000 779.7000 ;
	    RECT 239.4000 767.7000 240.6000 779.7000 ;
	    RECT 251.4000 777.4500 252.6000 777.6000 ;
	    RECT 280.2000 777.4500 281.4000 777.6000 ;
	    RECT 352.2000 777.4500 353.4000 777.6000 ;
	    RECT 251.4000 776.5500 353.4000 777.4500 ;
	    RECT 251.4000 776.4000 252.6000 776.5500 ;
	    RECT 280.2000 776.4000 281.4000 776.5500 ;
	    RECT 352.2000 776.4000 353.4000 776.5500 ;
	    RECT 364.2000 773.7000 365.4000 779.7000 ;
	    RECT 366.6000 774.6000 367.8000 779.7000 ;
	    RECT 366.3000 773.7000 367.8000 774.6000 ;
	    RECT 369.0000 773.7000 370.2000 780.6000 ;
	    RECT 366.3000 772.8000 367.2000 773.7000 ;
	    RECT 371.4000 772.8000 372.6000 779.7000 ;
	    RECT 373.8000 773.7000 375.0000 779.7000 ;
	    RECT 376.2000 775.5000 377.4000 779.7000 ;
	    RECT 378.6000 775.5000 379.8000 779.7000 ;
	    RECT 364.2000 771.9000 367.2000 772.8000 ;
	    RECT 232.2000 764.4000 233.4000 765.6000 ;
	    RECT 234.6000 763.5000 235.5000 767.7000 ;
	    RECT 237.0000 764.4000 238.2000 765.6000 ;
	    RECT 251.4000 765.4500 252.6000 765.6000 ;
	    RECT 287.4000 765.4500 288.6000 765.6000 ;
	    RECT 251.4000 764.5500 288.6000 765.4500 ;
	    RECT 251.4000 764.4000 252.6000 764.5500 ;
	    RECT 287.4000 764.4000 288.6000 764.5500 ;
	    RECT 239.4000 763.5000 240.6000 763.8000 ;
	    RECT 364.2000 763.5000 365.4000 771.9000 ;
	    RECT 368.1000 771.6000 374.4000 772.8000 ;
	    RECT 381.0000 772.5000 382.2000 779.7000 ;
	    RECT 383.4000 773.7000 384.6000 779.7000 ;
	    RECT 385.8000 772.5000 387.0000 779.7000 ;
	    RECT 388.2000 773.7000 389.4000 779.7000 ;
	    RECT 368.1000 771.0000 369.0000 771.6000 ;
	    RECT 366.6000 769.8000 369.0000 771.0000 ;
	    RECT 373.5000 770.7000 382.2000 771.6000 ;
	    RECT 370.5000 769.8000 372.6000 770.7000 ;
	    RECT 370.5000 769.5000 379.8000 769.8000 ;
	    RECT 371.7000 768.9000 379.8000 769.5000 ;
	    RECT 378.6000 768.6000 379.8000 768.9000 ;
	    RECT 381.3000 769.5000 382.2000 770.7000 ;
	    RECT 383.1000 770.4000 387.0000 771.6000 ;
	    RECT 390.6000 770.4000 391.8000 779.7000 ;
	    RECT 393.0000 775.5000 394.2000 779.7000 ;
	    RECT 395.4000 775.5000 396.6000 779.7000 ;
	    RECT 397.8000 775.5000 399.0000 779.7000 ;
	    RECT 400.2000 773.7000 401.4000 779.7000 ;
	    RECT 395.4000 771.6000 401.7000 772.8000 ;
	    RECT 402.6000 771.6000 403.8000 779.7000 ;
	    RECT 405.0000 773.7000 406.2000 779.7000 ;
	    RECT 407.4000 772.8000 408.6000 779.7000 ;
	    RECT 409.8000 773.7000 411.0000 779.7000 ;
	    RECT 407.4000 771.9000 411.3000 772.8000 ;
	    RECT 412.2000 772.5000 413.4000 779.7000 ;
	    RECT 414.6000 773.7000 415.8000 779.7000 ;
	    RECT 446.7000 773.7000 447.9000 779.7000 ;
	    RECT 402.6000 770.4000 406.5000 771.6000 ;
	    RECT 393.0000 769.5000 394.2000 769.8000 ;
	    RECT 381.3000 768.6000 394.2000 769.5000 ;
	    RECT 397.8000 769.5000 399.0000 769.8000 ;
	    RECT 410.4000 769.5000 411.3000 771.9000 ;
	    RECT 412.2000 770.4000 413.4000 771.6000 ;
	    RECT 447.0000 770.4000 448.2000 771.6000 ;
	    RECT 447.0000 769.5000 447.9000 770.4000 ;
	    RECT 397.8000 768.6000 411.3000 769.5000 ;
	    RECT 369.0000 767.4000 370.2000 768.6000 ;
	    RECT 374.1000 767.7000 375.3000 768.0000 ;
	    RECT 371.1000 766.8000 409.5000 767.7000 ;
	    RECT 408.3000 766.5000 409.5000 766.8000 ;
	    RECT 410.4000 765.9000 411.3000 768.6000 ;
	    RECT 412.2000 768.0000 413.4000 769.5000 ;
	    RECT 449.1000 768.6000 450.3000 779.7000 ;
	    RECT 431.4000 768.4500 432.6000 768.6000 ;
	    RECT 445.8000 768.4500 447.0000 768.6000 ;
	    RECT 412.2000 766.8000 413.7000 768.0000 ;
	    RECT 431.4000 767.5500 447.0000 768.4500 ;
	    RECT 431.4000 767.4000 432.6000 767.5500 ;
	    RECT 445.8000 767.4000 447.0000 767.5500 ;
	    RECT 448.8000 767.7000 450.3000 768.6000 ;
	    RECT 453.0000 767.7000 454.2000 779.7000 ;
	    RECT 563.4000 779.4000 564.6000 780.6000 ;
	    RECT 577.8000 773.7000 579.0000 779.7000 ;
	    RECT 580.2000 774.6000 581.4000 779.7000 ;
	    RECT 579.9000 773.7000 581.4000 774.6000 ;
	    RECT 582.6000 773.7000 583.8000 780.6000 ;
	    RECT 579.9000 772.8000 580.8000 773.7000 ;
	    RECT 585.0000 772.8000 586.2000 779.7000 ;
	    RECT 587.4000 773.7000 588.6000 779.7000 ;
	    RECT 589.8000 775.5000 591.0000 779.7000 ;
	    RECT 592.2000 775.5000 593.4000 779.7000 ;
	    RECT 577.8000 771.9000 580.8000 772.8000 ;
	    RECT 366.3000 765.0000 372.9000 765.9000 ;
	    RECT 366.3000 764.7000 367.5000 765.0000 ;
	    RECT 373.8000 764.4000 375.0000 765.6000 ;
	    RECT 375.9000 765.0000 401.4000 765.9000 ;
	    RECT 410.4000 765.0000 411.6000 765.9000 ;
	    RECT 400.2000 764.1000 401.4000 765.0000 ;
	    RECT 147.6000 761.7000 148.8000 762.0000 ;
	    RECT 147.6000 760.8000 154.2000 761.7000 ;
	    RECT 155.4000 761.4000 156.6000 762.6000 ;
	    RECT 153.0000 760.5000 154.2000 760.8000 ;
	    RECT 155.4000 760.2000 156.6000 760.5000 ;
	    RECT 133.8000 753.3000 135.0000 759.3000 ;
	    RECT 136.2000 758.1000 139.8000 759.3000 ;
	    RECT 143.4000 758.4000 144.9000 759.6000 ;
	    RECT 149.4000 758.4000 149.7000 759.6000 ;
	    RECT 150.6000 758.4000 151.8000 759.6000 ;
	    RECT 153.0000 759.3000 154.2000 759.6000 ;
	    RECT 158.7000 759.3000 159.9000 762.9000 ;
	    RECT 162.6000 762.3000 175.8000 763.5000 ;
	    RECT 232.2000 763.2000 233.4000 763.5000 ;
	    RECT 237.0000 763.2000 238.2000 763.5000 ;
	    RECT 167.7000 760.2000 172.2000 761.4000 ;
	    RECT 167.7000 759.3000 168.9000 760.2000 ;
	    RECT 153.0000 758.4000 159.9000 759.3000 ;
	    RECT 138.6000 753.3000 139.8000 758.1000 ;
	    RECT 165.0000 758.1000 168.9000 759.3000 ;
	    RECT 141.0000 753.3000 142.2000 757.5000 ;
	    RECT 143.4000 753.3000 144.6000 757.5000 ;
	    RECT 145.8000 753.3000 147.0000 757.5000 ;
	    RECT 148.2000 753.3000 149.4000 757.5000 ;
	    RECT 150.6000 753.3000 151.8000 756.3000 ;
	    RECT 153.0000 753.3000 154.2000 757.5000 ;
	    RECT 155.4000 753.3000 156.6000 756.3000 ;
	    RECT 157.8000 753.3000 159.0000 757.5000 ;
	    RECT 160.2000 753.3000 161.4000 757.5000 ;
	    RECT 162.6000 753.3000 163.8000 757.5000 ;
	    RECT 165.0000 753.3000 166.2000 758.1000 ;
	    RECT 169.8000 753.3000 171.0000 759.3000 ;
	    RECT 174.6000 753.3000 175.8000 762.3000 ;
	    RECT 191.4000 762.4500 192.6000 762.6000 ;
	    RECT 229.8000 762.4500 231.0000 762.6000 ;
	    RECT 191.4000 761.5500 231.0000 762.4500 ;
	    RECT 191.4000 761.4000 192.6000 761.5500 ;
	    RECT 229.8000 761.4000 231.0000 761.5500 ;
	    RECT 231.9000 760.8000 232.2000 762.3000 ;
	    RECT 234.6000 761.4000 235.8000 762.6000 ;
	    RECT 239.4000 762.4500 240.6000 762.6000 ;
	    RECT 256.2000 762.4500 257.4000 762.6000 ;
	    RECT 236.7000 761.4000 238.2000 762.3000 ;
	    RECT 239.4000 761.5500 257.4000 762.4500 ;
	    RECT 239.4000 761.4000 240.6000 761.5500 ;
	    RECT 256.2000 761.4000 257.4000 761.5500 ;
	    RECT 299.4000 762.4500 300.6000 762.6000 ;
	    RECT 359.4000 762.4500 360.6000 762.6000 ;
	    RECT 299.4000 761.5500 360.6000 762.4500 ;
	    RECT 299.4000 761.4000 300.6000 761.5500 ;
	    RECT 359.4000 761.4000 360.6000 761.5500 ;
	    RECT 364.2000 762.3000 377.4000 763.5000 ;
	    RECT 378.3000 762.9000 381.3000 764.1000 ;
	    RECT 387.0000 762.9000 391.8000 764.1000 ;
	    RECT 177.0000 759.4500 178.2000 759.6000 ;
	    RECT 181.8000 759.4500 183.0000 759.6000 ;
	    RECT 189.0000 759.4500 190.2000 759.6000 ;
	    RECT 177.0000 758.5500 190.2000 759.4500 ;
	    RECT 177.0000 758.4000 178.2000 758.5500 ;
	    RECT 181.8000 758.4000 183.0000 758.5500 ;
	    RECT 189.0000 758.4000 190.2000 758.5500 ;
	    RECT 189.0000 757.2000 190.2000 757.5000 ;
	    RECT 189.0000 753.3000 190.2000 756.3000 ;
	    RECT 191.4000 753.3000 192.6000 760.5000 ;
	    RECT 230.1000 759.3000 235.5000 759.9000 ;
	    RECT 237.3000 759.3000 238.2000 761.4000 ;
	    RECT 285.0000 759.4500 286.2000 759.6000 ;
	    RECT 361.8000 759.4500 363.0000 759.6000 ;
	    RECT 229.8000 759.0000 235.8000 759.3000 ;
	    RECT 229.8000 753.3000 231.0000 759.0000 ;
	    RECT 232.2000 753.3000 233.4000 758.1000 ;
	    RECT 234.6000 754.2000 235.8000 759.0000 ;
	    RECT 237.0000 755.1000 238.2000 759.3000 ;
	    RECT 239.4000 754.2000 240.6000 759.3000 ;
	    RECT 285.0000 758.5500 363.0000 759.4500 ;
	    RECT 285.0000 758.4000 286.2000 758.5500 ;
	    RECT 361.8000 758.4000 363.0000 758.5500 ;
	    RECT 275.4000 756.4500 276.6000 756.6000 ;
	    RECT 361.8000 756.4500 363.0000 756.6000 ;
	    RECT 275.4000 755.5500 363.0000 756.4500 ;
	    RECT 275.4000 755.4000 276.6000 755.5500 ;
	    RECT 361.8000 755.4000 363.0000 755.5500 ;
	    RECT 234.6000 753.3000 240.6000 754.2000 ;
	    RECT 364.2000 753.3000 365.4000 762.3000 ;
	    RECT 367.8000 760.2000 372.3000 761.4000 ;
	    RECT 371.1000 759.3000 372.3000 760.2000 ;
	    RECT 380.1000 759.3000 381.3000 762.9000 ;
	    RECT 383.4000 761.4000 384.6000 762.6000 ;
	    RECT 391.2000 761.7000 392.4000 762.0000 ;
	    RECT 385.8000 760.8000 392.4000 761.7000 ;
	    RECT 385.8000 760.5000 387.0000 760.8000 ;
	    RECT 383.4000 760.2000 384.6000 760.5000 ;
	    RECT 395.4000 759.6000 396.6000 763.8000 ;
	    RECT 404.1000 762.9000 409.8000 764.1000 ;
	    RECT 404.1000 761.1000 405.3000 762.9000 ;
	    RECT 410.7000 762.0000 411.6000 765.0000 ;
	    RECT 385.8000 759.3000 387.0000 759.6000 ;
	    RECT 369.0000 753.3000 370.2000 759.3000 ;
	    RECT 371.1000 758.1000 375.0000 759.3000 ;
	    RECT 380.1000 758.4000 387.0000 759.3000 ;
	    RECT 388.2000 758.4000 389.4000 759.6000 ;
	    RECT 390.3000 758.4000 390.6000 759.6000 ;
	    RECT 395.1000 758.4000 396.6000 759.6000 ;
	    RECT 402.6000 760.2000 405.3000 761.1000 ;
	    RECT 409.8000 761.1000 411.6000 762.0000 ;
	    RECT 402.6000 759.3000 403.8000 760.2000 ;
	    RECT 373.8000 753.3000 375.0000 758.1000 ;
	    RECT 400.2000 758.1000 403.8000 759.3000 ;
	    RECT 376.2000 753.3000 377.4000 757.5000 ;
	    RECT 378.6000 753.3000 379.8000 757.5000 ;
	    RECT 381.0000 753.3000 382.2000 757.5000 ;
	    RECT 383.4000 753.3000 384.6000 756.3000 ;
	    RECT 385.8000 753.3000 387.0000 757.5000 ;
	    RECT 388.2000 753.3000 389.4000 756.3000 ;
	    RECT 390.6000 753.3000 391.8000 757.5000 ;
	    RECT 393.0000 753.3000 394.2000 757.5000 ;
	    RECT 395.4000 753.3000 396.6000 757.5000 ;
	    RECT 397.8000 753.3000 399.0000 757.5000 ;
	    RECT 400.2000 753.3000 401.4000 758.1000 ;
	    RECT 405.0000 753.3000 406.2000 759.3000 ;
	    RECT 409.8000 753.3000 411.0000 761.1000 ;
	    RECT 412.5000 760.2000 413.7000 766.8000 ;
	    RECT 448.8000 762.6000 449.7000 767.7000 ;
	    RECT 450.6000 765.4500 451.8000 765.6000 ;
	    RECT 496.2000 765.4500 497.4000 765.6000 ;
	    RECT 450.6000 764.5500 497.4000 765.4500 ;
	    RECT 450.6000 764.4000 451.8000 764.5500 ;
	    RECT 496.2000 764.4000 497.4000 764.5500 ;
	    RECT 577.8000 763.5000 579.0000 771.9000 ;
	    RECT 581.7000 771.6000 588.0000 772.8000 ;
	    RECT 594.6000 772.5000 595.8000 779.7000 ;
	    RECT 597.0000 773.7000 598.2000 779.7000 ;
	    RECT 599.4000 772.5000 600.6000 779.7000 ;
	    RECT 601.8000 773.7000 603.0000 779.7000 ;
	    RECT 581.7000 771.0000 582.6000 771.6000 ;
	    RECT 580.2000 769.8000 582.6000 771.0000 ;
	    RECT 587.1000 770.7000 595.8000 771.6000 ;
	    RECT 584.1000 769.8000 586.2000 770.7000 ;
	    RECT 584.1000 769.5000 593.4000 769.8000 ;
	    RECT 585.3000 768.9000 593.4000 769.5000 ;
	    RECT 592.2000 768.6000 593.4000 768.9000 ;
	    RECT 594.9000 769.5000 595.8000 770.7000 ;
	    RECT 596.7000 770.4000 600.6000 771.6000 ;
	    RECT 604.2000 770.4000 605.4000 779.7000 ;
	    RECT 606.6000 775.5000 607.8000 779.7000 ;
	    RECT 609.0000 775.5000 610.2000 779.7000 ;
	    RECT 611.4000 775.5000 612.6000 779.7000 ;
	    RECT 613.8000 773.7000 615.0000 779.7000 ;
	    RECT 609.0000 771.6000 615.3000 772.8000 ;
	    RECT 616.2000 771.6000 617.4000 779.7000 ;
	    RECT 618.6000 773.7000 619.8000 779.7000 ;
	    RECT 621.0000 772.8000 622.2000 779.7000 ;
	    RECT 623.4000 773.7000 624.6000 779.7000 ;
	    RECT 621.0000 771.9000 624.9000 772.8000 ;
	    RECT 625.8000 772.5000 627.0000 779.7000 ;
	    RECT 628.2000 773.7000 629.4000 779.7000 ;
	    RECT 616.2000 770.4000 620.1000 771.6000 ;
	    RECT 606.6000 769.5000 607.8000 769.8000 ;
	    RECT 594.9000 768.6000 607.8000 769.5000 ;
	    RECT 611.4000 769.5000 612.6000 769.8000 ;
	    RECT 624.0000 769.5000 624.9000 771.9000 ;
	    RECT 625.8000 770.4000 627.0000 771.6000 ;
	    RECT 611.4000 768.6000 624.9000 769.5000 ;
	    RECT 582.6000 767.4000 583.8000 768.6000 ;
	    RECT 587.7000 767.7000 588.9000 768.0000 ;
	    RECT 584.7000 766.8000 623.1000 767.7000 ;
	    RECT 621.9000 766.5000 623.1000 766.8000 ;
	    RECT 624.0000 765.9000 624.9000 768.6000 ;
	    RECT 625.8000 768.0000 627.0000 769.5000 ;
	    RECT 654.6000 768.6000 655.8000 779.7000 ;
	    RECT 657.0000 769.5000 658.2000 779.7000 ;
	    RECT 659.4000 768.6000 660.6000 779.7000 ;
	    RECT 625.8000 766.8000 627.3000 768.0000 ;
	    RECT 654.6000 767.7000 660.6000 768.6000 ;
	    RECT 661.8000 767.7000 663.0000 779.7000 ;
	    RECT 688.2000 773.7000 689.4000 779.7000 ;
	    RECT 579.9000 765.0000 586.5000 765.9000 ;
	    RECT 579.9000 764.7000 581.1000 765.0000 ;
	    RECT 587.4000 764.4000 588.6000 765.6000 ;
	    RECT 589.5000 765.0000 615.0000 765.9000 ;
	    RECT 624.0000 765.0000 625.2000 765.9000 ;
	    RECT 613.8000 764.1000 615.0000 765.0000 ;
	    RECT 450.6000 763.2000 451.8000 763.5000 ;
	    RECT 445.8000 761.4000 447.0000 762.6000 ;
	    RECT 447.9000 761.4000 449.7000 762.6000 ;
	    RECT 453.0000 762.4500 454.2000 762.6000 ;
	    RECT 493.8000 762.4500 495.0000 762.6000 ;
	    RECT 451.8000 760.8000 452.1000 762.3000 ;
	    RECT 453.0000 761.5500 495.0000 762.4500 ;
	    RECT 453.0000 761.4000 454.2000 761.5500 ;
	    RECT 493.8000 761.4000 495.0000 761.5500 ;
	    RECT 577.8000 762.3000 591.0000 763.5000 ;
	    RECT 591.9000 762.9000 594.9000 764.1000 ;
	    RECT 600.6000 762.9000 605.4000 764.1000 ;
	    RECT 412.2000 759.0000 413.7000 760.2000 ;
	    RECT 446.1000 759.3000 447.0000 760.5000 ;
	    RECT 448.5000 759.3000 453.9000 759.9000 ;
	    RECT 412.2000 753.3000 413.4000 759.0000 ;
	    RECT 414.6000 753.3000 415.8000 756.3000 ;
	    RECT 445.8000 753.3000 447.0000 759.3000 ;
	    RECT 448.2000 759.0000 454.2000 759.3000 ;
	    RECT 448.2000 753.3000 449.4000 759.0000 ;
	    RECT 450.6000 753.3000 451.8000 758.1000 ;
	    RECT 453.0000 753.3000 454.2000 759.0000 ;
	    RECT 577.8000 753.3000 579.0000 762.3000 ;
	    RECT 581.4000 760.2000 585.9000 761.4000 ;
	    RECT 584.7000 759.3000 585.9000 760.2000 ;
	    RECT 593.7000 759.3000 594.9000 762.9000 ;
	    RECT 597.0000 761.4000 598.2000 762.6000 ;
	    RECT 604.8000 761.7000 606.0000 762.0000 ;
	    RECT 599.4000 760.8000 606.0000 761.7000 ;
	    RECT 599.4000 760.5000 600.6000 760.8000 ;
	    RECT 597.0000 760.2000 598.2000 760.5000 ;
	    RECT 609.0000 759.6000 610.2000 763.8000 ;
	    RECT 617.7000 762.9000 623.4000 764.1000 ;
	    RECT 617.7000 761.1000 618.9000 762.9000 ;
	    RECT 624.3000 762.0000 625.2000 765.0000 ;
	    RECT 599.4000 759.3000 600.6000 759.6000 ;
	    RECT 582.6000 753.3000 583.8000 759.3000 ;
	    RECT 584.7000 758.1000 588.6000 759.3000 ;
	    RECT 593.7000 758.4000 600.6000 759.3000 ;
	    RECT 601.8000 758.4000 603.0000 759.6000 ;
	    RECT 603.9000 758.4000 604.2000 759.6000 ;
	    RECT 608.7000 758.4000 610.2000 759.6000 ;
	    RECT 616.2000 760.2000 618.9000 761.1000 ;
	    RECT 623.4000 761.1000 625.2000 762.0000 ;
	    RECT 616.2000 759.3000 617.4000 760.2000 ;
	    RECT 587.4000 753.3000 588.6000 758.1000 ;
	    RECT 613.8000 758.1000 617.4000 759.3000 ;
	    RECT 589.8000 753.3000 591.0000 757.5000 ;
	    RECT 592.2000 753.3000 593.4000 757.5000 ;
	    RECT 594.6000 753.3000 595.8000 757.5000 ;
	    RECT 597.0000 753.3000 598.2000 756.3000 ;
	    RECT 599.4000 753.3000 600.6000 757.5000 ;
	    RECT 601.8000 753.3000 603.0000 756.3000 ;
	    RECT 604.2000 753.3000 605.4000 757.5000 ;
	    RECT 606.6000 753.3000 607.8000 757.5000 ;
	    RECT 609.0000 753.3000 610.2000 757.5000 ;
	    RECT 611.4000 753.3000 612.6000 757.5000 ;
	    RECT 613.8000 753.3000 615.0000 758.1000 ;
	    RECT 618.6000 753.3000 619.8000 759.3000 ;
	    RECT 623.4000 753.3000 624.6000 761.1000 ;
	    RECT 626.1000 760.2000 627.3000 766.8000 ;
	    RECT 661.8000 766.5000 662.7000 767.7000 ;
	    RECT 690.6000 766.5000 691.8000 779.7000 ;
	    RECT 693.0000 773.7000 694.2000 779.7000 ;
	    RECT 705.0000 773.7000 706.2000 779.7000 ;
	    RECT 693.0000 769.5000 694.2000 769.8000 ;
	    RECT 693.0000 767.4000 694.2000 768.6000 ;
	    RECT 645.0000 765.4500 646.2000 765.6000 ;
	    RECT 654.6000 765.4500 655.8000 765.6000 ;
	    RECT 645.0000 764.5500 655.8000 765.4500 ;
	    RECT 656.7000 764.7000 657.0000 766.2000 ;
	    RECT 659.4000 764.7000 660.9000 765.6000 ;
	    RECT 645.0000 764.4000 646.2000 764.5500 ;
	    RECT 654.6000 764.4000 655.8000 764.5500 ;
	    RECT 657.0000 763.5000 658.2000 763.8000 ;
	    RECT 657.0000 761.4000 658.2000 762.6000 ;
	    RECT 625.8000 759.0000 627.3000 760.2000 ;
	    RECT 659.4000 759.3000 660.3000 764.7000 ;
	    RECT 661.8000 764.4000 663.0000 765.6000 ;
	    RECT 664.2000 765.4500 665.4000 765.6000 ;
	    RECT 690.6000 765.4500 691.8000 765.6000 ;
	    RECT 664.2000 764.5500 691.8000 765.4500 ;
	    RECT 664.2000 764.4000 665.4000 764.5500 ;
	    RECT 690.6000 764.4000 691.8000 764.5500 ;
	    RECT 707.4000 763.5000 708.6000 779.7000 ;
	    RECT 719.4000 773.7000 720.6000 779.7000 ;
	    RECT 721.8000 763.5000 723.0000 779.7000 ;
	    RECT 745.8000 773.7000 747.0000 779.7000 ;
	    RECT 748.2000 773.7000 749.4000 779.7000 ;
	    RECT 750.6000 774.3000 751.8000 779.7000 ;
	    RECT 748.5000 773.4000 749.4000 773.7000 ;
	    RECT 753.0000 773.7000 754.2000 779.7000 ;
	    RECT 777.0000 773.7000 778.2000 779.7000 ;
	    RECT 779.4000 773.7000 780.6000 779.7000 ;
	    RECT 781.8000 774.3000 783.0000 779.7000 ;
	    RECT 753.0000 773.4000 753.9000 773.7000 ;
	    RECT 748.5000 772.5000 753.9000 773.4000 ;
	    RECT 779.7000 773.4000 780.6000 773.7000 ;
	    RECT 784.2000 773.7000 785.4000 779.7000 ;
	    RECT 784.2000 773.4000 785.1000 773.7000 ;
	    RECT 779.7000 772.5000 785.1000 773.4000 ;
	    RECT 750.6000 770.4000 751.8000 771.6000 ;
	    RECT 753.0000 769.5000 753.9000 772.5000 ;
	    RECT 781.8000 770.4000 783.0000 771.6000 ;
	    RECT 784.2000 769.5000 785.1000 772.5000 ;
	    RECT 750.6000 769.2000 751.8000 769.5000 ;
	    RECT 781.8000 769.2000 783.0000 769.5000 ;
	    RECT 804.3000 768.9000 805.5000 779.7000 ;
	    RECT 738.6000 768.4500 739.8000 768.6000 ;
	    RECT 745.8000 768.4500 747.0000 768.6000 ;
	    RECT 738.6000 767.5500 747.0000 768.4500 ;
	    RECT 738.6000 767.4000 739.8000 767.5500 ;
	    RECT 745.8000 767.4000 747.0000 767.5500 ;
	    RECT 753.0000 768.4500 754.2000 768.6000 ;
	    RECT 760.2000 768.4500 761.4000 768.6000 ;
	    RECT 765.0000 768.4500 766.2000 768.6000 ;
	    RECT 777.0000 768.4500 778.2000 768.6000 ;
	    RECT 753.0000 767.5500 758.8500 768.4500 ;
	    RECT 753.0000 767.4000 754.2000 767.5500 ;
	    RECT 745.8000 766.2000 747.0000 766.5000 ;
	    RECT 748.2000 764.4000 749.4000 765.6000 ;
	    RECT 750.3000 764.4000 750.6000 765.6000 ;
	    RECT 688.2000 761.4000 689.4000 762.6000 ;
	    RECT 688.2000 760.2000 689.4000 760.5000 ;
	    RECT 625.8000 753.3000 627.0000 759.0000 ;
	    RECT 628.2000 753.3000 629.4000 756.3000 ;
	    RECT 655.5000 753.3000 656.7000 759.3000 ;
	    RECT 659.4000 753.3000 660.6000 759.3000 ;
	    RECT 661.8000 758.4000 663.0000 759.6000 ;
	    RECT 690.6000 759.3000 691.8000 763.5000 ;
	    RECT 753.0000 762.6000 753.9000 766.5000 ;
	    RECT 757.9500 765.4500 758.8500 767.5500 ;
	    RECT 760.2000 767.5500 778.2000 768.4500 ;
	    RECT 760.2000 767.4000 761.4000 767.5500 ;
	    RECT 765.0000 767.4000 766.2000 767.5500 ;
	    RECT 777.0000 767.4000 778.2000 767.5500 ;
	    RECT 784.2000 768.4500 785.4000 768.6000 ;
	    RECT 801.0000 768.4500 802.2000 768.6000 ;
	    RECT 784.2000 767.5500 802.2000 768.4500 ;
	    RECT 804.3000 767.7000 807.0000 768.9000 ;
	    RECT 808.2000 767.7000 809.4000 779.7000 ;
	    RECT 822.6000 773.7000 823.8000 779.7000 ;
	    RECT 784.2000 767.4000 785.4000 767.5500 ;
	    RECT 801.0000 767.4000 802.2000 767.5500 ;
	    RECT 803.4000 766.5000 804.6000 766.8000 ;
	    RECT 777.0000 766.2000 778.2000 766.5000 ;
	    RECT 769.8000 765.4500 771.0000 765.6000 ;
	    RECT 757.9500 764.5500 771.0000 765.4500 ;
	    RECT 769.8000 764.4000 771.0000 764.5500 ;
	    RECT 779.4000 764.4000 780.6000 765.6000 ;
	    RECT 781.5000 764.4000 781.8000 765.6000 ;
	    RECT 784.2000 762.6000 785.1000 766.5000 ;
	    RECT 803.4000 764.4000 804.6000 765.6000 ;
	    RECT 805.8000 763.5000 806.7000 767.7000 ;
	    RECT 808.2000 765.4500 809.4000 765.6000 ;
	    RECT 822.6000 765.4500 823.8000 765.6000 ;
	    RECT 808.2000 764.5500 823.8000 765.4500 ;
	    RECT 808.2000 764.4000 809.4000 764.5500 ;
	    RECT 822.6000 764.4000 823.8000 764.5500 ;
	    RECT 825.0000 763.5000 826.2000 779.7000 ;
	    RECT 853.8000 767.7000 855.0000 779.7000 ;
	    RECT 857.7000 767.7000 860.7000 779.7000 ;
	    RECT 863.4000 767.7000 864.6000 779.7000 ;
	    RECT 899.4000 767.7000 900.6000 779.7000 ;
	    RECT 903.3000 767.7000 906.3000 779.7000 ;
	    RECT 909.0000 767.7000 910.2000 779.7000 ;
	    RECT 935.4000 767.7000 936.6000 779.7000 ;
	    RECT 939.3000 768.6000 940.5000 779.7000 ;
	    RECT 941.7000 773.7000 942.9000 779.7000 ;
	    RECT 941.4000 770.4000 942.6000 771.6000 ;
	    RECT 941.7000 769.5000 942.6000 770.4000 ;
	    RECT 939.3000 767.7000 940.8000 768.6000 ;
	    RECT 827.4000 765.4500 828.6000 765.6000 ;
	    RECT 853.8000 765.4500 855.0000 765.6000 ;
	    RECT 827.4000 764.5500 855.0000 765.4500 ;
	    RECT 827.4000 764.4000 828.6000 764.5500 ;
	    RECT 853.8000 764.4000 855.0000 764.5500 ;
	    RECT 856.2000 764.4000 857.4000 765.6000 ;
	    RECT 858.6000 763.5000 859.5000 767.7000 ;
	    RECT 861.0000 764.4000 862.2000 765.6000 ;
	    RECT 873.0000 765.4500 874.2000 765.6000 ;
	    RECT 899.4000 765.4500 900.6000 765.6000 ;
	    RECT 873.0000 764.5500 900.6000 765.4500 ;
	    RECT 873.0000 764.4000 874.2000 764.5500 ;
	    RECT 899.4000 764.4000 900.6000 764.5500 ;
	    RECT 901.8000 764.4000 903.0000 765.6000 ;
	    RECT 863.4000 763.5000 864.6000 763.8000 ;
	    RECT 904.2000 763.5000 905.1000 767.7000 ;
	    RECT 906.6000 764.4000 907.8000 765.6000 ;
	    RECT 913.8000 765.4500 915.0000 765.6000 ;
	    RECT 937.8000 765.4500 939.0000 765.6000 ;
	    RECT 913.8000 764.5500 939.0000 765.4500 ;
	    RECT 913.8000 764.4000 915.0000 764.5500 ;
	    RECT 937.8000 764.4000 939.0000 764.5500 ;
	    RECT 909.0000 763.5000 910.2000 763.8000 ;
	    RECT 856.2000 763.2000 857.4000 763.5000 ;
	    RECT 861.0000 763.2000 862.2000 763.5000 ;
	    RECT 901.8000 763.2000 903.0000 763.5000 ;
	    RECT 906.6000 763.2000 907.8000 763.5000 ;
	    RECT 937.8000 763.2000 939.0000 763.5000 ;
	    RECT 939.9000 762.6000 940.8000 767.7000 ;
	    RECT 942.6000 767.4000 943.8000 768.6000 ;
	    RECT 957.0000 763.5000 958.2000 779.7000 ;
	    RECT 959.4000 773.7000 960.6000 779.7000 ;
	    RECT 973.8000 773.7000 975.0000 779.7000 ;
	    RECT 976.2000 763.5000 977.4000 779.7000 ;
	    RECT 1000.2000 767.7000 1001.4000 779.7000 ;
	    RECT 1004.1000 768.6000 1005.3000 779.7000 ;
	    RECT 1006.5000 773.7000 1007.7000 779.7000 ;
	    RECT 1006.2000 770.4000 1007.4000 771.6000 ;
	    RECT 1006.5000 769.5000 1007.4000 770.4000 ;
	    RECT 1004.1000 767.7000 1005.6000 768.6000 ;
	    RECT 1002.6000 765.4500 1003.8000 765.6000 ;
	    RECT 997.9500 764.5500 1003.8000 765.4500 ;
	    RECT 707.4000 762.4500 708.6000 762.6000 ;
	    RECT 719.4000 762.4500 720.6000 762.6000 ;
	    RECT 707.4000 761.5500 720.6000 762.4500 ;
	    RECT 707.4000 761.4000 708.6000 761.5500 ;
	    RECT 719.4000 761.4000 720.6000 761.5500 ;
	    RECT 721.8000 762.4500 723.0000 762.6000 ;
	    RECT 741.0000 762.4500 742.2000 762.6000 ;
	    RECT 721.8000 761.5500 742.2000 762.4500 ;
	    RECT 751.5000 762.3000 753.9000 762.6000 ;
	    RECT 782.7000 762.3000 785.1000 762.6000 ;
	    RECT 721.8000 761.4000 723.0000 761.5500 ;
	    RECT 741.0000 761.4000 742.2000 761.5500 ;
	    RECT 700.2000 759.4500 701.4000 759.6000 ;
	    RECT 705.0000 759.4500 706.2000 759.6000 ;
	    RECT 661.5000 757.2000 662.7000 757.5000 ;
	    RECT 661.8000 753.3000 663.0000 756.3000 ;
	    RECT 688.2000 753.3000 689.4000 759.3000 ;
	    RECT 690.6000 758.4000 693.3000 759.3000 ;
	    RECT 700.2000 758.5500 706.2000 759.4500 ;
	    RECT 700.2000 758.4000 701.4000 758.5500 ;
	    RECT 705.0000 758.4000 706.2000 758.5500 ;
	    RECT 692.1000 753.3000 693.3000 758.4000 ;
	    RECT 705.0000 757.2000 706.2000 757.5000 ;
	    RECT 705.0000 753.3000 706.2000 756.3000 ;
	    RECT 707.4000 753.3000 708.6000 760.5000 ;
	    RECT 712.2000 759.4500 713.4000 759.6000 ;
	    RECT 719.4000 759.4500 720.6000 759.6000 ;
	    RECT 712.2000 758.5500 720.6000 759.4500 ;
	    RECT 712.2000 758.4000 713.4000 758.5500 ;
	    RECT 719.4000 758.4000 720.6000 758.5500 ;
	    RECT 719.4000 757.2000 720.6000 757.5000 ;
	    RECT 719.4000 753.3000 720.6000 756.3000 ;
	    RECT 721.8000 753.3000 723.0000 760.5000 ;
	    RECT 745.8000 753.3000 747.0000 762.3000 ;
	    RECT 751.2000 761.7000 753.9000 762.3000 ;
	    RECT 751.2000 753.3000 752.4000 761.7000 ;
	    RECT 760.2000 756.4500 761.4000 756.6000 ;
	    RECT 774.6000 756.4500 775.8000 756.6000 ;
	    RECT 760.2000 755.5500 775.8000 756.4500 ;
	    RECT 760.2000 755.4000 761.4000 755.5500 ;
	    RECT 774.6000 755.4000 775.8000 755.5500 ;
	    RECT 777.0000 753.3000 778.2000 762.3000 ;
	    RECT 782.4000 761.7000 785.1000 762.3000 ;
	    RECT 786.6000 762.4500 787.8000 762.6000 ;
	    RECT 805.8000 762.4500 807.0000 762.6000 ;
	    RECT 782.4000 753.3000 783.6000 761.7000 ;
	    RECT 786.6000 761.5500 807.0000 762.4500 ;
	    RECT 786.6000 761.4000 787.8000 761.5500 ;
	    RECT 805.8000 761.4000 807.0000 761.5500 ;
	    RECT 825.0000 762.4500 826.2000 762.6000 ;
	    RECT 853.8000 762.4500 855.0000 762.6000 ;
	    RECT 825.0000 761.5500 855.0000 762.4500 ;
	    RECT 825.0000 761.4000 826.2000 761.5500 ;
	    RECT 853.8000 761.4000 855.0000 761.5500 ;
	    RECT 855.9000 760.8000 856.2000 762.3000 ;
	    RECT 858.6000 761.4000 859.8000 762.6000 ;
	    RECT 860.7000 761.4000 862.2000 762.3000 ;
	    RECT 863.4000 761.4000 864.6000 762.6000 ;
	    RECT 885.0000 762.4500 886.2000 762.6000 ;
	    RECT 899.4000 762.4500 900.6000 762.6000 ;
	    RECT 885.0000 761.5500 900.6000 762.4500 ;
	    RECT 885.0000 761.4000 886.2000 761.5500 ;
	    RECT 899.4000 761.4000 900.6000 761.5500 ;
	    RECT 805.8000 756.3000 806.7000 760.5000 ;
	    RECT 808.2000 758.4000 809.4000 759.6000 ;
	    RECT 822.6000 758.4000 823.8000 759.6000 ;
	    RECT 808.2000 757.2000 809.4000 757.5000 ;
	    RECT 822.6000 757.2000 823.8000 757.5000 ;
	    RECT 803.4000 753.3000 804.6000 756.3000 ;
	    RECT 805.8000 753.3000 807.0000 756.3000 ;
	    RECT 808.2000 753.3000 809.4000 756.3000 ;
	    RECT 822.6000 753.3000 823.8000 756.3000 ;
	    RECT 825.0000 753.3000 826.2000 760.5000 ;
	    RECT 854.1000 759.3000 859.5000 759.9000 ;
	    RECT 861.3000 759.3000 862.2000 761.4000 ;
	    RECT 901.5000 760.8000 901.8000 762.3000 ;
	    RECT 904.2000 761.4000 905.4000 762.6000 ;
	    RECT 909.0000 762.4500 910.2000 762.6000 ;
	    RECT 911.4000 762.4500 912.6000 762.6000 ;
	    RECT 906.3000 761.4000 907.8000 762.3000 ;
	    RECT 909.0000 761.5500 912.6000 762.4500 ;
	    RECT 909.0000 761.4000 910.2000 761.5500 ;
	    RECT 911.4000 761.4000 912.6000 761.5500 ;
	    RECT 935.4000 761.4000 936.6000 762.6000 ;
	    RECT 899.7000 759.3000 905.1000 759.9000 ;
	    RECT 906.9000 759.3000 907.8000 761.4000 ;
	    RECT 937.5000 760.8000 937.8000 762.3000 ;
	    RECT 939.9000 761.4000 941.7000 762.6000 ;
	    RECT 942.6000 762.4500 943.8000 762.6000 ;
	    RECT 947.4000 762.4500 948.6000 762.6000 ;
	    RECT 942.6000 761.5500 948.6000 762.4500 ;
	    RECT 942.6000 761.4000 943.8000 761.5500 ;
	    RECT 947.4000 761.4000 948.6000 761.5500 ;
	    RECT 949.8000 762.4500 951.0000 762.6000 ;
	    RECT 957.0000 762.4500 958.2000 762.6000 ;
	    RECT 949.8000 761.5500 958.2000 762.4500 ;
	    RECT 949.8000 761.4000 951.0000 761.5500 ;
	    RECT 957.0000 761.4000 958.2000 761.5500 ;
	    RECT 976.2000 762.4500 977.4000 762.6000 ;
	    RECT 997.9500 762.4500 998.8500 764.5500 ;
	    RECT 1002.6000 764.4000 1003.8000 764.5500 ;
	    RECT 1002.6000 763.2000 1003.8000 763.5000 ;
	    RECT 1004.7000 762.6000 1005.6000 767.7000 ;
	    RECT 1007.4000 768.4500 1008.6000 768.6000 ;
	    RECT 1065.0000 768.4500 1066.2001 768.6000 ;
	    RECT 1007.4000 767.5500 1066.2001 768.4500 ;
	    RECT 1007.4000 767.4000 1008.6000 767.5500 ;
	    RECT 1065.0000 767.4000 1066.2001 767.5500 ;
	    RECT 1077.0000 766.8000 1078.2001 779.7000 ;
	    RECT 1079.4000 767.7000 1080.6000 779.7000 ;
	    RECT 1083.3000 773.7000 1085.1000 779.7000 ;
	    RECT 1087.8000 773.7000 1089.0000 779.7000 ;
	    RECT 1090.2001 773.7000 1091.4000 779.7000 ;
	    RECT 1092.6000 773.7000 1093.8000 779.7000 ;
	    RECT 1096.8000 774.6000 1098.0000 779.7000 ;
	    RECT 1096.8000 773.7000 1099.8000 774.6000 ;
	    RECT 1084.2001 772.5000 1085.4000 773.7000 ;
	    RECT 1090.5000 772.8000 1091.4000 773.7000 ;
	    RECT 1089.3000 771.9000 1094.7001 772.8000 ;
	    RECT 1098.6000 772.5000 1099.8000 773.7000 ;
	    RECT 1089.3000 771.6000 1090.5000 771.9000 ;
	    RECT 1093.5000 771.6000 1094.7001 771.9000 ;
	    RECT 1083.0000 769.8000 1085.1000 771.0000 ;
	    RECT 1084.2001 768.3000 1085.1000 769.8000 ;
	    RECT 1087.5000 769.5000 1090.8000 770.4000 ;
	    RECT 1087.5000 769.2000 1088.7001 769.5000 ;
	    RECT 1084.2001 767.4000 1087.8000 768.3000 ;
	    RECT 1077.0000 766.5000 1083.3000 766.8000 ;
	    RECT 1079.1000 765.9000 1083.3000 766.5000 ;
	    RECT 1082.1000 765.6000 1083.3000 765.9000 ;
	    RECT 1055.4000 765.4500 1056.6000 765.6000 ;
	    RECT 1077.0000 765.4500 1078.2001 765.6000 ;
	    RECT 1055.4000 764.5500 1078.2001 765.4500 ;
	    RECT 1055.4000 764.4000 1056.6000 764.5500 ;
	    RECT 1077.0000 764.4000 1078.2001 764.5500 ;
	    RECT 1079.7001 764.7000 1080.9000 765.0000 ;
	    RECT 1079.7001 763.8000 1085.4000 764.7000 ;
	    RECT 1084.2001 763.5000 1085.4000 763.8000 ;
	    RECT 976.2000 761.5500 998.8500 762.4500 ;
	    RECT 976.2000 761.4000 977.4000 761.5500 ;
	    RECT 1000.2000 761.4000 1001.4000 762.6000 ;
	    RECT 1002.3000 760.8000 1002.6000 762.3000 ;
	    RECT 1004.7000 761.4000 1006.5000 762.6000 ;
	    RECT 1007.4000 762.4500 1008.6000 762.6000 ;
	    RECT 1043.4000 762.4500 1044.6000 762.6000 ;
	    RECT 1007.4000 761.5500 1044.6000 762.4500 ;
	    RECT 1007.4000 761.4000 1008.6000 761.5500 ;
	    RECT 1043.4000 761.4000 1044.6000 761.5500 ;
	    RECT 1077.0000 760.8000 1078.2001 763.5000 ;
	    RECT 1086.9000 762.6000 1087.8000 767.4000 ;
	    RECT 1089.9000 767.7000 1090.8000 769.5000 ;
	    RECT 1091.7001 769.5000 1092.9000 769.8000 ;
	    RECT 1098.6000 769.5000 1099.8000 769.8000 ;
	    RECT 1091.7001 768.6000 1099.8000 769.5000 ;
	    RECT 1101.0000 768.0000 1102.2001 779.7000 ;
	    RECT 1089.9000 767.1000 1097.1000 767.7000 ;
	    RECT 1103.4000 767.1000 1104.6000 779.7000 ;
	    RECT 1122.6000 773.7000 1123.8000 779.7000 ;
	    RECT 1122.6000 769.5000 1123.8000 769.8000 ;
	    RECT 1117.8000 768.4500 1119.0000 768.6000 ;
	    RECT 1122.6000 768.4500 1123.8000 768.6000 ;
	    RECT 1117.8000 767.5500 1123.8000 768.4500 ;
	    RECT 1117.8000 767.4000 1119.0000 767.5500 ;
	    RECT 1122.6000 767.4000 1123.8000 767.5500 ;
	    RECT 1089.9000 766.8000 1104.6000 767.1000 ;
	    RECT 1095.9000 766.5000 1104.6000 766.8000 ;
	    RECT 1125.0000 766.5000 1126.2001 779.7000 ;
	    RECT 1127.4000 773.7000 1128.6000 779.7000 ;
	    RECT 1151.4000 779.4000 1152.6000 780.6000 ;
	    RECT 1158.6000 767.7000 1159.8000 779.7000 ;
	    RECT 1162.5000 768.6000 1163.7001 779.7000 ;
	    RECT 1164.9000 773.7000 1166.1000 779.7000 ;
	    RECT 1185.0000 773.7000 1186.2001 779.7000 ;
	    RECT 1164.6000 770.4000 1165.8000 771.6000 ;
	    RECT 1164.9000 769.5000 1165.8000 770.4000 ;
	    RECT 1185.0000 769.5000 1186.2001 769.8000 ;
	    RECT 1162.5000 767.7000 1164.0000 768.6000 ;
	    RECT 1096.2001 766.2000 1104.6000 766.5000 ;
	    RECT 1093.8000 764.4000 1095.0000 765.6000 ;
	    RECT 1125.0000 765.4500 1126.2001 765.6000 ;
	    RECT 1144.2001 765.4500 1145.4000 765.6000 ;
	    RECT 1095.9000 764.4000 1101.3000 765.3000 ;
	    RECT 1125.0000 764.5500 1145.4000 765.4500 ;
	    RECT 1125.0000 764.4000 1126.2001 764.5500 ;
	    RECT 1144.2001 764.4000 1145.4000 764.5500 ;
	    RECT 1161.0000 764.4000 1162.2001 765.6000 ;
	    RECT 1100.1000 764.1000 1101.3000 764.4000 ;
	    RECT 1097.7001 762.6000 1098.9000 762.9000 ;
	    RECT 1086.9000 761.7000 1100.1000 762.6000 ;
	    RECT 1087.5000 761.4000 1088.7001 761.7000 ;
	    RECT 935.7000 759.3000 941.1000 759.9000 ;
	    RECT 942.6000 759.3000 943.5000 760.5000 ;
	    RECT 853.8000 759.0000 859.8000 759.3000 ;
	    RECT 853.8000 753.3000 855.0000 759.0000 ;
	    RECT 856.2000 753.3000 857.4000 758.1000 ;
	    RECT 858.6000 754.2000 859.8000 759.0000 ;
	    RECT 861.0000 755.1000 862.2000 759.3000 ;
	    RECT 863.4000 754.2000 864.6000 759.3000 ;
	    RECT 899.4000 759.0000 905.4000 759.3000 ;
	    RECT 875.4000 756.4500 876.6000 756.6000 ;
	    RECT 889.8000 756.4500 891.0000 756.6000 ;
	    RECT 875.4000 755.5500 891.0000 756.4500 ;
	    RECT 875.4000 755.4000 876.6000 755.5500 ;
	    RECT 889.8000 755.4000 891.0000 755.5500 ;
	    RECT 858.6000 753.3000 864.6000 754.2000 ;
	    RECT 899.4000 753.3000 900.6000 759.0000 ;
	    RECT 901.8000 753.3000 903.0000 758.1000 ;
	    RECT 904.2000 754.2000 905.4000 759.0000 ;
	    RECT 906.6000 755.1000 907.8000 759.3000 ;
	    RECT 909.0000 754.2000 910.2000 759.3000 ;
	    RECT 904.2000 753.3000 910.2000 754.2000 ;
	    RECT 935.4000 759.0000 941.4000 759.3000 ;
	    RECT 935.4000 753.3000 936.6000 759.0000 ;
	    RECT 937.8000 753.3000 939.0000 758.1000 ;
	    RECT 940.2000 753.3000 941.4000 759.0000 ;
	    RECT 942.6000 753.3000 943.8000 759.3000 ;
	    RECT 957.0000 753.3000 958.2000 760.5000 ;
	    RECT 959.4000 758.4000 960.6000 759.6000 ;
	    RECT 969.0000 759.4500 970.2000 759.6000 ;
	    RECT 973.8000 759.4500 975.0000 759.6000 ;
	    RECT 969.0000 758.5500 975.0000 759.4500 ;
	    RECT 969.0000 758.4000 970.2000 758.5500 ;
	    RECT 973.8000 758.4000 975.0000 758.5500 ;
	    RECT 959.4000 757.2000 960.6000 757.5000 ;
	    RECT 973.8000 757.2000 975.0000 757.5000 ;
	    RECT 959.4000 753.3000 960.6000 756.3000 ;
	    RECT 973.8000 753.3000 975.0000 756.3000 ;
	    RECT 976.2000 753.3000 977.4000 760.5000 ;
	    RECT 1000.5000 759.3000 1005.9000 759.9000 ;
	    RECT 1007.4000 759.3000 1008.3000 760.5000 ;
	    RECT 1077.0000 759.9000 1082.7001 760.8000 ;
	    RECT 1000.2000 759.0000 1006.2000 759.3000 ;
	    RECT 1000.2000 753.3000 1001.4000 759.0000 ;
	    RECT 1002.6000 753.3000 1003.8000 758.1000 ;
	    RECT 1005.0000 753.3000 1006.2000 759.0000 ;
	    RECT 1007.4000 753.3000 1008.6000 759.3000 ;
	    RECT 1077.0000 753.3000 1078.2001 759.9000 ;
	    RECT 1081.5000 759.6000 1082.7001 759.9000 ;
	    RECT 1079.4000 753.3000 1080.6000 759.0000 ;
	    RECT 1096.2001 758.4000 1097.1000 761.7000 ;
	    RECT 1101.0000 761.4000 1102.2001 762.6000 ;
	    RECT 1103.1000 761.4000 1103.4000 762.6000 ;
	    RECT 1093.5000 758.1000 1094.7001 758.4000 ;
	    RECT 1084.2001 756.3000 1085.4000 757.5000 ;
	    RECT 1090.5000 757.2000 1094.7001 758.1000 ;
	    RECT 1096.2001 757.2000 1097.4000 758.4000 ;
	    RECT 1090.5000 756.3000 1091.4000 757.2000 ;
	    RECT 1098.6000 756.3000 1099.8000 757.5000 ;
	    RECT 1083.3000 755.4000 1085.4000 756.3000 ;
	    RECT 1083.3000 753.3000 1085.1000 755.4000 ;
	    RECT 1087.8000 753.3000 1089.0000 756.3000 ;
	    RECT 1090.2001 753.3000 1091.4000 756.3000 ;
	    RECT 1092.6000 753.3000 1094.1000 756.3000 ;
	    RECT 1096.8000 755.4000 1099.8000 756.3000 ;
	    RECT 1096.8000 753.3000 1098.0000 755.4000 ;
	    RECT 1101.0000 753.3000 1102.2001 759.3000 ;
	    RECT 1103.4000 753.3000 1104.6000 760.5000 ;
	    RECT 1125.0000 759.3000 1126.2001 763.5000 ;
	    RECT 1161.0000 763.2000 1162.2001 763.5000 ;
	    RECT 1163.1000 762.6000 1164.0000 767.7000 ;
	    RECT 1165.8000 767.4000 1167.0000 768.6000 ;
	    RECT 1170.6000 768.4500 1171.8000 768.6000 ;
	    RECT 1185.0000 768.4500 1186.2001 768.6000 ;
	    RECT 1170.6000 767.5500 1186.2001 768.4500 ;
	    RECT 1170.6000 767.4000 1171.8000 767.5500 ;
	    RECT 1185.0000 767.4000 1186.2001 767.5500 ;
	    RECT 1165.9501 765.4500 1166.8500 767.4000 ;
	    RECT 1187.4000 766.5000 1188.6000 779.7000 ;
	    RECT 1189.8000 773.7000 1191.0000 779.7000 ;
	    RECT 1201.8000 773.7000 1203.0000 779.7000 ;
	    RECT 1187.4000 765.4500 1188.6000 765.6000 ;
	    RECT 1165.9501 764.5500 1188.6000 765.4500 ;
	    RECT 1187.4000 764.4000 1188.6000 764.5500 ;
	    RECT 1204.2001 763.5000 1205.4000 779.7000 ;
	    RECT 1230.6000 767.7000 1231.8000 779.7000 ;
	    RECT 1234.5000 768.6000 1235.7001 779.7000 ;
	    RECT 1236.9000 773.7000 1238.1000 779.7000 ;
	    RECT 1236.6000 770.4000 1237.8000 771.6000 ;
	    RECT 1236.9000 769.5000 1237.8000 770.4000 ;
	    RECT 1234.5000 767.7000 1236.0000 768.6000 ;
	    RECT 1233.0000 765.4500 1234.2001 765.6000 ;
	    RECT 1209.1500 764.5500 1234.2001 765.4500 ;
	    RECT 1127.4000 762.4500 1128.6000 762.6000 ;
	    RECT 1151.4000 762.4500 1152.6000 762.6000 ;
	    RECT 1158.6000 762.4500 1159.8000 762.6000 ;
	    RECT 1127.4000 761.5500 1159.8000 762.4500 ;
	    RECT 1127.4000 761.4000 1128.6000 761.5500 ;
	    RECT 1151.4000 761.4000 1152.6000 761.5500 ;
	    RECT 1158.6000 761.4000 1159.8000 761.5500 ;
	    RECT 1160.7001 760.8000 1161.0000 762.3000 ;
	    RECT 1163.1000 761.4000 1164.9000 762.6000 ;
	    RECT 1165.8000 762.4500 1167.0000 762.6000 ;
	    RECT 1180.2001 762.4500 1181.4000 762.6000 ;
	    RECT 1165.8000 761.5500 1181.4000 762.4500 ;
	    RECT 1165.8000 761.4000 1167.0000 761.5500 ;
	    RECT 1180.2001 761.4000 1181.4000 761.5500 ;
	    RECT 1127.4000 760.2000 1128.6000 760.5000 ;
	    RECT 1158.9000 759.3000 1164.3000 759.9000 ;
	    RECT 1165.8000 759.3000 1166.7001 760.5000 ;
	    RECT 1187.4000 759.3000 1188.6000 763.5000 ;
	    RECT 1189.8000 762.4500 1191.0000 762.6000 ;
	    RECT 1199.4000 762.4500 1200.6000 762.6000 ;
	    RECT 1189.8000 761.5500 1200.6000 762.4500 ;
	    RECT 1189.8000 761.4000 1191.0000 761.5500 ;
	    RECT 1199.4000 761.4000 1200.6000 761.5500 ;
	    RECT 1204.2001 762.4500 1205.4000 762.6000 ;
	    RECT 1209.1500 762.4500 1210.0500 764.5500 ;
	    RECT 1233.0000 764.4000 1234.2001 764.5500 ;
	    RECT 1233.0000 763.2000 1234.2001 763.5000 ;
	    RECT 1235.1000 762.6000 1236.0000 767.7000 ;
	    RECT 1237.8000 768.4500 1239.0000 768.6000 ;
	    RECT 1240.2001 768.4500 1241.4000 768.6000 ;
	    RECT 1237.8000 767.5500 1241.4000 768.4500 ;
	    RECT 1237.8000 767.4000 1239.0000 767.5500 ;
	    RECT 1240.2001 767.4000 1241.4000 767.5500 ;
	    RECT 1307.4000 767.1000 1308.6000 779.7000 ;
	    RECT 1309.8000 768.0000 1311.0000 779.7000 ;
	    RECT 1314.0000 774.6000 1315.2001 779.7000 ;
	    RECT 1312.2001 773.7000 1315.2001 774.6000 ;
	    RECT 1318.2001 773.7000 1319.4000 779.7000 ;
	    RECT 1320.6000 773.7000 1321.8000 779.7000 ;
	    RECT 1323.0000 773.7000 1324.2001 779.7000 ;
	    RECT 1326.9000 773.7000 1328.7001 779.7000 ;
	    RECT 1312.2001 772.5000 1313.4000 773.7000 ;
	    RECT 1320.6000 772.8000 1321.5000 773.7000 ;
	    RECT 1317.3000 771.9000 1322.7001 772.8000 ;
	    RECT 1326.6000 772.5000 1327.8000 773.7000 ;
	    RECT 1317.3000 771.6000 1318.5000 771.9000 ;
	    RECT 1321.5000 771.6000 1322.7001 771.9000 ;
	    RECT 1312.2001 769.5000 1313.4000 769.8000 ;
	    RECT 1319.1000 769.5000 1320.3000 769.8000 ;
	    RECT 1312.2001 768.6000 1320.3000 769.5000 ;
	    RECT 1321.2001 769.5000 1324.5000 770.4000 ;
	    RECT 1321.2001 767.7000 1322.1000 769.5000 ;
	    RECT 1323.3000 769.2000 1324.5000 769.5000 ;
	    RECT 1326.9000 769.8000 1329.0000 771.0000 ;
	    RECT 1326.9000 768.3000 1327.8000 769.8000 ;
	    RECT 1314.9000 767.1000 1322.1000 767.7000 ;
	    RECT 1307.4000 766.8000 1322.1000 767.1000 ;
	    RECT 1324.2001 767.4000 1327.8000 768.3000 ;
	    RECT 1331.4000 767.7000 1332.6000 779.7000 ;
	    RECT 1307.4000 766.5000 1316.1000 766.8000 ;
	    RECT 1307.4000 766.2000 1315.8000 766.5000 ;
	    RECT 1310.7001 764.4000 1316.1000 765.3000 ;
	    RECT 1317.0000 764.4000 1318.2001 765.6000 ;
	    RECT 1310.7001 764.1000 1311.9000 764.4000 ;
	    RECT 1313.1000 762.6000 1314.3000 762.9000 ;
	    RECT 1324.2001 762.6000 1325.1000 767.4000 ;
	    RECT 1333.8000 766.8000 1335.0000 779.7000 ;
	    RECT 1328.7001 766.5000 1335.0000 766.8000 ;
	    RECT 1410.6000 767.1000 1411.8000 779.7000 ;
	    RECT 1413.0000 768.0000 1414.2001 779.7000 ;
	    RECT 1417.2001 774.6000 1418.4000 779.7000 ;
	    RECT 1415.4000 773.7000 1418.4000 774.6000 ;
	    RECT 1421.4000 773.7000 1422.6000 779.7000 ;
	    RECT 1423.8000 773.7000 1425.0000 779.7000 ;
	    RECT 1426.2001 773.7000 1427.4000 779.7000 ;
	    RECT 1430.1000 773.7000 1431.9000 779.7000 ;
	    RECT 1415.4000 772.5000 1416.6000 773.7000 ;
	    RECT 1423.8000 772.8000 1424.7001 773.7000 ;
	    RECT 1420.5000 771.9000 1425.9000 772.8000 ;
	    RECT 1429.8000 772.5000 1431.0000 773.7000 ;
	    RECT 1420.5000 771.6000 1421.7001 771.9000 ;
	    RECT 1424.7001 771.6000 1425.9000 771.9000 ;
	    RECT 1415.4000 769.5000 1416.6000 769.8000 ;
	    RECT 1422.3000 769.5000 1423.5000 769.8000 ;
	    RECT 1415.4000 768.6000 1423.5000 769.5000 ;
	    RECT 1424.4000 769.5000 1427.7001 770.4000 ;
	    RECT 1424.4000 767.7000 1425.3000 769.5000 ;
	    RECT 1426.5000 769.2000 1427.7001 769.5000 ;
	    RECT 1430.1000 769.8000 1432.2001 771.0000 ;
	    RECT 1430.1000 768.3000 1431.0000 769.8000 ;
	    RECT 1418.1000 767.1000 1425.3000 767.7000 ;
	    RECT 1410.6000 766.8000 1425.3000 767.1000 ;
	    RECT 1427.4000 767.4000 1431.0000 768.3000 ;
	    RECT 1434.6000 767.7000 1435.8000 779.7000 ;
	    RECT 1410.6000 766.5000 1419.3000 766.8000 ;
	    RECT 1328.7001 765.9000 1332.9000 766.5000 ;
	    RECT 1410.6000 766.2000 1419.0000 766.5000 ;
	    RECT 1328.7001 765.6000 1329.9000 765.9000 ;
	    RECT 1333.8000 765.4500 1335.0000 765.6000 ;
	    RECT 1374.6000 765.4500 1375.8000 765.6000 ;
	    RECT 1331.1000 764.7000 1332.3000 765.0000 ;
	    RECT 1326.6000 763.8000 1332.3000 764.7000 ;
	    RECT 1333.8000 764.5500 1375.8000 765.4500 ;
	    RECT 1333.8000 764.4000 1335.0000 764.5500 ;
	    RECT 1374.6000 764.4000 1375.8000 764.5500 ;
	    RECT 1413.9000 764.4000 1419.3000 765.3000 ;
	    RECT 1420.2001 764.4000 1421.4000 765.6000 ;
	    RECT 1413.9000 764.1000 1415.1000 764.4000 ;
	    RECT 1326.6000 763.5000 1327.8000 763.8000 ;
	    RECT 1204.2001 761.5500 1210.0500 762.4500 ;
	    RECT 1211.4000 762.4500 1212.6000 762.6000 ;
	    RECT 1230.6000 762.4500 1231.8000 762.6000 ;
	    RECT 1211.4000 761.5500 1231.8000 762.4500 ;
	    RECT 1204.2001 761.4000 1205.4000 761.5500 ;
	    RECT 1211.4000 761.4000 1212.6000 761.5500 ;
	    RECT 1230.6000 761.4000 1231.8000 761.5500 ;
	    RECT 1232.7001 760.8000 1233.0000 762.3000 ;
	    RECT 1235.1000 761.4000 1236.9000 762.6000 ;
	    RECT 1237.8000 762.4500 1239.0000 762.6000 ;
	    RECT 1249.8000 762.4500 1251.0000 762.6000 ;
	    RECT 1237.8000 761.5500 1251.0000 762.4500 ;
	    RECT 1237.8000 761.4000 1239.0000 761.5500 ;
	    RECT 1249.8000 761.4000 1251.0000 761.5500 ;
	    RECT 1308.6000 761.4000 1308.9000 762.6000 ;
	    RECT 1309.8000 761.4000 1311.0000 762.6000 ;
	    RECT 1311.9000 761.7000 1325.1000 762.6000 ;
	    RECT 1189.8000 760.2000 1191.0000 760.5000 ;
	    RECT 1123.5000 758.4000 1126.2001 759.3000 ;
	    RECT 1123.5000 753.3000 1124.7001 758.4000 ;
	    RECT 1127.4000 753.3000 1128.6000 759.3000 ;
	    RECT 1158.6000 759.0000 1164.6000 759.3000 ;
	    RECT 1158.6000 753.3000 1159.8000 759.0000 ;
	    RECT 1161.0000 753.3000 1162.2001 758.1000 ;
	    RECT 1163.4000 753.3000 1164.6000 759.0000 ;
	    RECT 1165.8000 753.3000 1167.0000 759.3000 ;
	    RECT 1185.9000 758.4000 1188.6000 759.3000 ;
	    RECT 1185.9000 753.3000 1187.1000 758.4000 ;
	    RECT 1189.8000 753.3000 1191.0000 759.3000 ;
	    RECT 1201.8000 758.4000 1203.0000 759.6000 ;
	    RECT 1201.8000 757.2000 1203.0000 757.5000 ;
	    RECT 1201.8000 753.3000 1203.0000 756.3000 ;
	    RECT 1204.2001 753.3000 1205.4000 760.5000 ;
	    RECT 1230.9000 759.3000 1236.3000 759.9000 ;
	    RECT 1237.8000 759.3000 1238.7001 760.5000 ;
	    RECT 1230.6000 759.0000 1236.6000 759.3000 ;
	    RECT 1230.6000 753.3000 1231.8000 759.0000 ;
	    RECT 1233.0000 753.3000 1234.2001 758.1000 ;
	    RECT 1235.4000 753.3000 1236.6000 759.0000 ;
	    RECT 1237.8000 753.3000 1239.0000 759.3000 ;
	    RECT 1307.4000 753.3000 1308.6000 760.5000 ;
	    RECT 1309.8000 753.3000 1311.0000 759.3000 ;
	    RECT 1314.9000 758.4000 1315.8000 761.7000 ;
	    RECT 1323.3000 761.4000 1324.5000 761.7000 ;
	    RECT 1333.8000 760.8000 1335.0000 763.5000 ;
	    RECT 1416.3000 762.6000 1417.5000 762.9000 ;
	    RECT 1427.4000 762.6000 1428.3000 767.4000 ;
	    RECT 1437.0000 766.8000 1438.2001 779.7000 ;
	    RECT 1431.9000 766.5000 1438.2001 766.8000 ;
	    RECT 1431.9000 765.9000 1436.1000 766.5000 ;
	    RECT 1431.9000 765.6000 1433.1000 765.9000 ;
	    RECT 1437.0000 765.4500 1438.2001 765.6000 ;
	    RECT 1439.4000 765.4500 1440.6000 765.6000 ;
	    RECT 1434.3000 764.7000 1435.5000 765.0000 ;
	    RECT 1429.8000 763.8000 1435.5000 764.7000 ;
	    RECT 1437.0000 764.5500 1440.6000 765.4500 ;
	    RECT 1437.0000 764.4000 1438.2001 764.5500 ;
	    RECT 1439.4000 764.4000 1440.6000 764.5500 ;
	    RECT 1429.8000 763.5000 1431.0000 763.8000 ;
	    RECT 1451.4000 763.5000 1452.6000 779.7000 ;
	    RECT 1453.8000 773.7000 1455.0000 779.7000 ;
	    RECT 1458.6000 779.4000 1459.8000 780.6000 ;
	    RECT 1480.2001 767.7000 1481.4000 779.7000 ;
	    RECT 1484.1000 768.6000 1485.3000 779.7000 ;
	    RECT 1486.5000 773.7000 1487.7001 779.7000 ;
	    RECT 1486.2001 770.4000 1487.4000 771.6000 ;
	    RECT 1486.5000 769.5000 1487.4000 770.4000 ;
	    RECT 1484.1000 767.7000 1485.6000 768.6000 ;
	    RECT 1482.6000 765.4500 1483.8000 765.6000 ;
	    RECT 1477.9501 764.5500 1483.8000 765.4500 ;
	    RECT 1411.8000 761.4000 1412.1000 762.6000 ;
	    RECT 1413.0000 761.4000 1414.2001 762.6000 ;
	    RECT 1415.1000 761.7000 1428.3000 762.6000 ;
	    RECT 1329.3000 759.9000 1335.0000 760.8000 ;
	    RECT 1329.3000 759.6000 1330.5000 759.9000 ;
	    RECT 1312.2001 756.3000 1313.4000 757.5000 ;
	    RECT 1314.6000 757.2000 1315.8000 758.4000 ;
	    RECT 1317.3000 758.1000 1318.5000 758.4000 ;
	    RECT 1317.3000 757.2000 1321.5000 758.1000 ;
	    RECT 1320.6000 756.3000 1321.5000 757.2000 ;
	    RECT 1326.6000 756.3000 1327.8000 757.5000 ;
	    RECT 1312.2001 755.4000 1315.2001 756.3000 ;
	    RECT 1314.0000 753.3000 1315.2001 755.4000 ;
	    RECT 1317.9000 753.3000 1319.4000 756.3000 ;
	    RECT 1320.6000 753.3000 1321.8000 756.3000 ;
	    RECT 1323.0000 753.3000 1324.2001 756.3000 ;
	    RECT 1326.6000 755.4000 1328.7001 756.3000 ;
	    RECT 1326.9000 753.3000 1328.7001 755.4000 ;
	    RECT 1331.4000 753.3000 1332.6000 759.0000 ;
	    RECT 1333.8000 753.3000 1335.0000 759.9000 ;
	    RECT 1410.6000 753.3000 1411.8000 760.5000 ;
	    RECT 1413.0000 753.3000 1414.2001 759.3000 ;
	    RECT 1418.1000 758.4000 1419.0000 761.7000 ;
	    RECT 1426.5000 761.4000 1427.7001 761.7000 ;
	    RECT 1437.0000 760.8000 1438.2001 763.5000 ;
	    RECT 1451.4000 762.4500 1452.6000 762.6000 ;
	    RECT 1477.9501 762.4500 1478.8500 764.5500 ;
	    RECT 1482.6000 764.4000 1483.8000 764.5500 ;
	    RECT 1482.6000 763.2000 1483.8000 763.5000 ;
	    RECT 1484.7001 762.6000 1485.6000 767.7000 ;
	    RECT 1487.4000 768.4500 1488.6000 768.6000 ;
	    RECT 1499.4000 768.4500 1500.6000 768.6000 ;
	    RECT 1487.4000 767.5500 1500.6000 768.4500 ;
	    RECT 1511.4000 767.7000 1512.6000 779.7000 ;
	    RECT 1513.8000 768.6000 1515.0000 779.7000 ;
	    RECT 1516.2001 769.5000 1517.4000 779.7000 ;
	    RECT 1518.6000 768.6000 1519.8000 779.7000 ;
	    RECT 1545.9000 773.7000 1547.1000 779.7000 ;
	    RECT 1546.2001 770.4000 1547.4000 771.6000 ;
	    RECT 1546.2001 769.5000 1547.1000 770.4000 ;
	    RECT 1548.3000 768.6000 1549.5000 779.7000 ;
	    RECT 1513.8000 767.7000 1519.8000 768.6000 ;
	    RECT 1523.4000 768.4500 1524.6000 768.6000 ;
	    RECT 1533.0000 768.4500 1534.2001 768.6000 ;
	    RECT 1545.0000 768.4500 1546.2001 768.6000 ;
	    RECT 1487.4000 767.4000 1488.6000 767.5500 ;
	    RECT 1499.4000 767.4000 1500.6000 767.5500 ;
	    RECT 1511.7001 766.5000 1512.6000 767.7000 ;
	    RECT 1523.4000 767.5500 1546.2001 768.4500 ;
	    RECT 1523.4000 767.4000 1524.6000 767.5500 ;
	    RECT 1533.0000 767.4000 1534.2001 767.5500 ;
	    RECT 1545.0000 767.4000 1546.2001 767.5500 ;
	    RECT 1548.0000 767.7000 1549.5000 768.6000 ;
	    RECT 1552.2001 767.7000 1553.4000 779.7000 ;
	    RECT 1511.4000 764.4000 1512.6000 765.6000 ;
	    RECT 1513.5000 764.7000 1515.0000 765.6000 ;
	    RECT 1517.4000 764.7000 1517.7001 766.2000 ;
	    RECT 1451.4000 761.5500 1478.8500 762.4500 ;
	    RECT 1451.4000 761.4000 1452.6000 761.5500 ;
	    RECT 1480.2001 761.4000 1481.4000 762.6000 ;
	    RECT 1482.3000 760.8000 1482.6000 762.3000 ;
	    RECT 1484.7001 761.4000 1486.5000 762.6000 ;
	    RECT 1487.4000 762.4500 1488.6000 762.6000 ;
	    RECT 1504.2001 762.4500 1505.4000 762.6000 ;
	    RECT 1487.4000 761.5500 1505.4000 762.4500 ;
	    RECT 1487.4000 761.4000 1488.6000 761.5500 ;
	    RECT 1504.2001 761.4000 1505.4000 761.5500 ;
	    RECT 1432.5000 759.9000 1438.2001 760.8000 ;
	    RECT 1432.5000 759.6000 1433.7001 759.9000 ;
	    RECT 1415.4000 756.3000 1416.6000 757.5000 ;
	    RECT 1417.8000 757.2000 1419.0000 758.4000 ;
	    RECT 1420.5000 758.1000 1421.7001 758.4000 ;
	    RECT 1420.5000 757.2000 1424.7001 758.1000 ;
	    RECT 1423.8000 756.3000 1424.7001 757.2000 ;
	    RECT 1429.8000 756.3000 1431.0000 757.5000 ;
	    RECT 1415.4000 755.4000 1418.4000 756.3000 ;
	    RECT 1417.2001 753.3000 1418.4000 755.4000 ;
	    RECT 1421.1000 753.3000 1422.6000 756.3000 ;
	    RECT 1423.8000 753.3000 1425.0000 756.3000 ;
	    RECT 1426.2001 753.3000 1427.4000 756.3000 ;
	    RECT 1429.8000 755.4000 1431.9000 756.3000 ;
	    RECT 1430.1000 753.3000 1431.9000 755.4000 ;
	    RECT 1434.6000 753.3000 1435.8000 759.0000 ;
	    RECT 1437.0000 753.3000 1438.2001 759.9000 ;
	    RECT 1451.4000 753.3000 1452.6000 760.5000 ;
	    RECT 1453.8000 759.4500 1455.0000 759.6000 ;
	    RECT 1461.0000 759.4500 1462.2001 759.6000 ;
	    RECT 1453.8000 758.5500 1462.2001 759.4500 ;
	    RECT 1480.5000 759.3000 1485.9000 759.9000 ;
	    RECT 1487.4000 759.3000 1488.3000 760.5000 ;
	    RECT 1492.2001 759.4500 1493.4000 759.6000 ;
	    RECT 1511.4000 759.4500 1512.6000 759.6000 ;
	    RECT 1453.8000 758.4000 1455.0000 758.5500 ;
	    RECT 1461.0000 758.4000 1462.2001 758.5500 ;
	    RECT 1480.2001 759.0000 1486.2001 759.3000 ;
	    RECT 1453.8000 757.2000 1455.0000 757.5000 ;
	    RECT 1453.8000 753.3000 1455.0000 756.3000 ;
	    RECT 1480.2001 753.3000 1481.4000 759.0000 ;
	    RECT 1482.6000 753.3000 1483.8000 758.1000 ;
	    RECT 1485.0000 753.3000 1486.2001 759.0000 ;
	    RECT 1487.4000 753.3000 1488.6000 759.3000 ;
	    RECT 1492.2001 758.5500 1512.6000 759.4500 ;
	    RECT 1514.1000 759.3000 1515.0000 764.7000 ;
	    RECT 1518.6000 764.4000 1519.8000 765.6000 ;
	    RECT 1516.2001 763.5000 1517.4000 763.8000 ;
	    RECT 1548.0000 762.6000 1548.9000 767.7000 ;
	    RECT 1549.8000 764.4000 1551.0000 765.6000 ;
	    RECT 1549.8000 763.2000 1551.0000 763.5000 ;
	    RECT 1516.2001 761.4000 1517.4000 762.6000 ;
	    RECT 1530.6000 762.4500 1531.8000 762.6000 ;
	    RECT 1545.0000 762.4500 1546.2001 762.6000 ;
	    RECT 1530.6000 761.5500 1546.2001 762.4500 ;
	    RECT 1530.6000 761.4000 1531.8000 761.5500 ;
	    RECT 1545.0000 761.4000 1546.2001 761.5500 ;
	    RECT 1547.1000 761.4000 1548.9000 762.6000 ;
	    RECT 1551.0000 760.8000 1551.3000 762.3000 ;
	    RECT 1552.2001 761.4000 1553.4000 762.6000 ;
	    RECT 1545.3000 759.3000 1546.2001 760.5000 ;
	    RECT 1547.7001 759.3000 1553.1000 759.9000 ;
	    RECT 1492.2001 758.4000 1493.4000 758.5500 ;
	    RECT 1511.4000 758.4000 1512.6000 758.5500 ;
	    RECT 1511.7001 757.2000 1512.9000 757.5000 ;
	    RECT 1511.4000 753.3000 1512.6000 756.3000 ;
	    RECT 1513.8000 753.3000 1515.0000 759.3000 ;
	    RECT 1517.7001 753.3000 1518.9000 759.3000 ;
	    RECT 1545.0000 753.3000 1546.2001 759.3000 ;
	    RECT 1547.4000 759.0000 1553.4000 759.3000 ;
	    RECT 1547.4000 753.3000 1548.6000 759.0000 ;
	    RECT 1549.8000 753.3000 1551.0000 758.1000 ;
	    RECT 1552.2001 753.3000 1553.4000 759.0000 ;
	    RECT 1.2000 750.6000 1569.0000 752.4000 ;
	    RECT 124.2000 746.7000 125.4000 749.7000 ;
	    RECT 126.6000 744.0000 127.8000 749.7000 ;
	    RECT 126.3000 742.8000 127.8000 744.0000 ;
	    RECT 126.3000 736.2000 127.5000 742.8000 ;
	    RECT 129.0000 741.9000 130.2000 749.7000 ;
	    RECT 133.8000 743.7000 135.0000 749.7000 ;
	    RECT 138.6000 744.9000 139.8000 749.7000 ;
	    RECT 141.0000 745.5000 142.2000 749.7000 ;
	    RECT 143.4000 745.5000 144.6000 749.7000 ;
	    RECT 145.8000 745.5000 147.0000 749.7000 ;
	    RECT 148.2000 745.5000 149.4000 749.7000 ;
	    RECT 150.6000 746.7000 151.8000 749.7000 ;
	    RECT 153.0000 745.5000 154.2000 749.7000 ;
	    RECT 155.4000 746.7000 156.6000 749.7000 ;
	    RECT 157.8000 745.5000 159.0000 749.7000 ;
	    RECT 160.2000 745.5000 161.4000 749.7000 ;
	    RECT 162.6000 745.5000 163.8000 749.7000 ;
	    RECT 136.2000 743.7000 139.8000 744.9000 ;
	    RECT 165.0000 744.9000 166.2000 749.7000 ;
	    RECT 136.2000 742.8000 137.4000 743.7000 ;
	    RECT 128.4000 741.0000 130.2000 741.9000 ;
	    RECT 134.7000 741.9000 137.4000 742.8000 ;
	    RECT 143.4000 743.4000 144.9000 744.6000 ;
	    RECT 149.4000 743.4000 149.7000 744.6000 ;
	    RECT 150.6000 743.4000 151.8000 744.6000 ;
	    RECT 153.0000 743.7000 159.9000 744.6000 ;
	    RECT 165.0000 743.7000 168.9000 744.9000 ;
	    RECT 169.8000 743.7000 171.0000 749.7000 ;
	    RECT 153.0000 743.4000 154.2000 743.7000 ;
	    RECT 128.4000 738.0000 129.3000 741.0000 ;
	    RECT 134.7000 740.1000 135.9000 741.9000 ;
	    RECT 130.2000 738.9000 135.9000 740.1000 ;
	    RECT 143.4000 739.2000 144.6000 743.4000 ;
	    RECT 155.4000 742.5000 156.6000 742.8000 ;
	    RECT 153.0000 742.2000 154.2000 742.5000 ;
	    RECT 147.6000 741.3000 154.2000 742.2000 ;
	    RECT 147.6000 741.0000 148.8000 741.3000 ;
	    RECT 155.4000 740.4000 156.6000 741.6000 ;
	    RECT 158.7000 740.1000 159.9000 743.7000 ;
	    RECT 167.7000 742.8000 168.9000 743.7000 ;
	    RECT 167.7000 741.6000 172.2000 742.8000 ;
	    RECT 174.6000 740.7000 175.8000 749.7000 ;
	    RECT 193.8000 746.7000 195.0000 749.7000 ;
	    RECT 196.2000 746.7000 197.4000 749.7000 ;
	    RECT 198.6000 746.7000 199.8000 749.7000 ;
	    RECT 193.8000 745.5000 195.0000 745.8000 ;
	    RECT 193.8000 743.4000 195.0000 744.6000 ;
	    RECT 196.5000 742.5000 197.4000 746.7000 ;
	    RECT 225.0000 743.7000 226.2000 749.7000 ;
	    RECT 228.9000 744.6000 230.1000 749.7000 ;
	    RECT 244.2000 746.7000 245.4000 749.7000 ;
	    RECT 244.2000 745.5000 245.4000 745.8000 ;
	    RECT 227.4000 743.7000 230.1000 744.6000 ;
	    RECT 239.4000 744.4500 240.6000 744.6000 ;
	    RECT 244.2000 744.4500 245.4000 744.6000 ;
	    RECT 225.0000 742.5000 226.2000 742.8000 ;
	    RECT 148.2000 738.9000 153.0000 740.1000 ;
	    RECT 158.7000 738.9000 161.7000 740.1000 ;
	    RECT 162.6000 739.5000 175.8000 740.7000 ;
	    RECT 196.2000 741.4500 197.4000 741.6000 ;
	    RECT 225.0000 741.4500 226.2000 741.6000 ;
	    RECT 196.2000 740.5500 226.2000 741.4500 ;
	    RECT 196.2000 740.4000 197.4000 740.5500 ;
	    RECT 225.0000 740.4000 226.2000 740.5500 ;
	    RECT 227.4000 739.5000 228.6000 743.7000 ;
	    RECT 239.4000 743.5500 245.4000 744.4500 ;
	    RECT 239.4000 743.4000 240.6000 743.5500 ;
	    RECT 244.2000 743.4000 245.4000 743.5500 ;
	    RECT 246.6000 742.5000 247.8000 749.7000 ;
	    RECT 266.7000 744.6000 267.9000 749.7000 ;
	    RECT 266.7000 743.7000 269.4000 744.6000 ;
	    RECT 270.6000 743.7000 271.8000 749.7000 ;
	    RECT 244.2000 741.4500 245.4000 741.6000 ;
	    RECT 246.6000 741.4500 247.8000 741.6000 ;
	    RECT 244.2000 740.5500 247.8000 741.4500 ;
	    RECT 244.2000 740.4000 245.4000 740.5500 ;
	    RECT 246.6000 740.4000 247.8000 740.5500 ;
	    RECT 268.2000 739.5000 269.4000 743.7000 ;
	    RECT 270.6000 742.5000 271.8000 742.8000 ;
	    RECT 282.6000 742.5000 283.8000 749.7000 ;
	    RECT 285.0000 746.7000 286.2000 749.7000 ;
	    RECT 299.4000 746.7000 300.6000 749.7000 ;
	    RECT 285.0000 745.5000 286.2000 745.8000 ;
	    RECT 299.4000 745.5000 300.6000 745.8000 ;
	    RECT 285.0000 743.4000 286.2000 744.6000 ;
	    RECT 299.4000 743.4000 300.6000 744.6000 ;
	    RECT 301.8000 742.5000 303.0000 749.7000 ;
	    RECT 316.2000 746.7000 317.4000 749.7000 ;
	    RECT 316.2000 745.5000 317.4000 745.8000 ;
	    RECT 316.2000 743.4000 317.4000 744.6000 ;
	    RECT 318.6000 742.5000 319.8000 749.7000 ;
	    RECT 349.8000 748.8000 355.8000 749.7000 ;
	    RECT 349.8000 743.7000 351.0000 748.8000 ;
	    RECT 352.2000 743.7000 353.4000 747.9000 ;
	    RECT 354.6000 744.0000 355.8000 748.8000 ;
	    RECT 357.0000 744.9000 358.2000 749.7000 ;
	    RECT 359.4000 744.0000 360.6000 749.7000 ;
	    RECT 354.6000 743.7000 360.6000 744.0000 ;
	    RECT 352.2000 741.6000 353.1000 743.7000 ;
	    RECT 354.9000 743.1000 360.3000 743.7000 ;
	    RECT 270.6000 740.4000 271.8000 741.6000 ;
	    RECT 282.6000 741.4500 283.8000 741.6000 ;
	    RECT 285.0000 741.4500 286.2000 741.6000 ;
	    RECT 282.6000 740.5500 286.2000 741.4500 ;
	    RECT 282.6000 740.4000 283.8000 740.5500 ;
	    RECT 285.0000 740.4000 286.2000 740.5500 ;
	    RECT 287.4000 741.4500 288.6000 741.6000 ;
	    RECT 301.8000 741.4500 303.0000 741.6000 ;
	    RECT 287.4000 740.5500 303.0000 741.4500 ;
	    RECT 287.4000 740.4000 288.6000 740.5500 ;
	    RECT 301.8000 740.4000 303.0000 740.5500 ;
	    RECT 318.6000 741.4500 319.8000 741.6000 ;
	    RECT 349.8000 741.4500 351.0000 741.6000 ;
	    RECT 318.6000 740.5500 351.0000 741.4500 ;
	    RECT 352.2000 740.7000 353.7000 741.6000 ;
	    RECT 318.6000 740.4000 319.8000 740.5500 ;
	    RECT 349.8000 740.4000 351.0000 740.5500 ;
	    RECT 354.6000 740.4000 355.8000 741.6000 ;
	    RECT 358.2000 740.7000 358.5000 742.2000 ;
	    RECT 359.4000 741.4500 360.6000 741.6000 ;
	    RECT 419.4000 741.4500 420.6000 741.6000 ;
	    RECT 359.4000 740.5500 420.6000 741.4500 ;
	    RECT 359.4000 740.4000 360.6000 740.5500 ;
	    RECT 419.4000 740.4000 420.6000 740.5500 ;
	    RECT 491.4000 740.7000 492.6000 749.7000 ;
	    RECT 496.2000 743.7000 497.4000 749.7000 ;
	    RECT 501.0000 744.9000 502.2000 749.7000 ;
	    RECT 503.4000 745.5000 504.6000 749.7000 ;
	    RECT 505.8000 745.5000 507.0000 749.7000 ;
	    RECT 508.2000 745.5000 509.4000 749.7000 ;
	    RECT 510.6000 746.7000 511.8000 749.7000 ;
	    RECT 513.0000 745.5000 514.2000 749.7000 ;
	    RECT 515.4000 746.7000 516.6000 749.7000 ;
	    RECT 517.8000 745.5000 519.0000 749.7000 ;
	    RECT 520.2000 745.5000 521.4000 749.7000 ;
	    RECT 522.6000 745.5000 523.8000 749.7000 ;
	    RECT 525.0000 745.5000 526.2000 749.7000 ;
	    RECT 498.3000 743.7000 502.2000 744.9000 ;
	    RECT 527.4000 744.9000 528.6000 749.7000 ;
	    RECT 507.3000 743.7000 514.2000 744.6000 ;
	    RECT 498.3000 742.8000 499.5000 743.7000 ;
	    RECT 495.0000 741.6000 499.5000 742.8000 ;
	    RECT 352.2000 739.5000 353.4000 739.8000 ;
	    RECT 357.0000 739.5000 358.2000 739.8000 ;
	    RECT 491.4000 739.5000 504.6000 740.7000 ;
	    RECT 507.3000 740.1000 508.5000 743.7000 ;
	    RECT 513.0000 743.4000 514.2000 743.7000 ;
	    RECT 515.4000 743.4000 516.6000 744.6000 ;
	    RECT 517.5000 743.4000 517.8000 744.6000 ;
	    RECT 522.3000 743.4000 523.8000 744.6000 ;
	    RECT 527.4000 743.7000 531.0000 744.9000 ;
	    RECT 532.2000 743.7000 533.4000 749.7000 ;
	    RECT 510.6000 742.5000 511.8000 742.8000 ;
	    RECT 513.0000 742.2000 514.2000 742.5000 ;
	    RECT 510.6000 740.4000 511.8000 741.6000 ;
	    RECT 513.0000 741.3000 519.6000 742.2000 ;
	    RECT 518.4000 741.0000 519.6000 741.3000 ;
	    RECT 138.6000 738.0000 139.8000 738.9000 ;
	    RECT 128.4000 737.1000 129.6000 738.0000 ;
	    RECT 138.6000 737.1000 164.1000 738.0000 ;
	    RECT 165.0000 737.4000 166.2000 738.6000 ;
	    RECT 172.5000 738.0000 173.7000 738.3000 ;
	    RECT 167.1000 737.1000 173.7000 738.0000 ;
	    RECT 126.3000 735.0000 127.8000 736.2000 ;
	    RECT 126.6000 733.5000 127.8000 735.0000 ;
	    RECT 128.7000 734.4000 129.6000 737.1000 ;
	    RECT 130.5000 736.2000 131.7000 736.5000 ;
	    RECT 130.5000 735.3000 168.9000 736.2000 ;
	    RECT 164.7000 735.0000 165.9000 735.3000 ;
	    RECT 169.8000 734.4000 171.0000 735.6000 ;
	    RECT 128.7000 733.5000 142.2000 734.4000 ;
	    RECT 90.6000 732.4500 91.8000 732.6000 ;
	    RECT 97.8000 732.4500 99.0000 732.6000 ;
	    RECT 126.6000 732.4500 127.8000 732.6000 ;
	    RECT 90.6000 731.5500 127.8000 732.4500 ;
	    RECT 90.6000 731.4000 91.8000 731.5500 ;
	    RECT 97.8000 731.4000 99.0000 731.5500 ;
	    RECT 126.6000 731.4000 127.8000 731.5500 ;
	    RECT 128.7000 731.1000 129.6000 733.5000 ;
	    RECT 141.0000 733.2000 142.2000 733.5000 ;
	    RECT 145.8000 733.5000 158.7000 734.4000 ;
	    RECT 145.8000 733.2000 147.0000 733.5000 ;
	    RECT 133.5000 731.4000 137.4000 732.6000 ;
	    RECT 124.2000 723.3000 125.4000 729.3000 ;
	    RECT 126.6000 723.3000 127.8000 730.5000 ;
	    RECT 128.7000 730.2000 132.6000 731.1000 ;
	    RECT 129.0000 723.3000 130.2000 729.3000 ;
	    RECT 131.4000 723.3000 132.6000 730.2000 ;
	    RECT 133.8000 723.3000 135.0000 729.3000 ;
	    RECT 136.2000 723.3000 137.4000 731.4000 ;
	    RECT 138.3000 730.2000 144.6000 731.4000 ;
	    RECT 138.6000 723.3000 139.8000 729.3000 ;
	    RECT 141.0000 723.3000 142.2000 727.5000 ;
	    RECT 143.4000 723.3000 144.6000 727.5000 ;
	    RECT 145.8000 723.3000 147.0000 727.5000 ;
	    RECT 148.2000 723.3000 149.4000 732.6000 ;
	    RECT 153.0000 731.4000 156.9000 732.6000 ;
	    RECT 157.8000 732.3000 158.7000 733.5000 ;
	    RECT 160.2000 734.1000 161.4000 734.4000 ;
	    RECT 160.2000 733.5000 168.3000 734.1000 ;
	    RECT 160.2000 733.2000 169.5000 733.5000 ;
	    RECT 167.4000 732.3000 169.5000 733.2000 ;
	    RECT 157.8000 731.4000 166.5000 732.3000 ;
	    RECT 171.0000 732.0000 173.4000 733.2000 ;
	    RECT 171.0000 731.4000 171.9000 732.0000 ;
	    RECT 150.6000 723.3000 151.8000 729.3000 ;
	    RECT 153.0000 723.3000 154.2000 730.5000 ;
	    RECT 155.4000 723.3000 156.6000 729.3000 ;
	    RECT 157.8000 723.3000 159.0000 730.5000 ;
	    RECT 165.6000 730.2000 171.9000 731.4000 ;
	    RECT 174.6000 731.1000 175.8000 739.5000 ;
	    RECT 196.5000 735.3000 197.4000 739.5000 ;
	    RECT 198.6000 738.4500 199.8000 738.6000 ;
	    RECT 215.4000 738.4500 216.6000 738.6000 ;
	    RECT 198.6000 737.5500 216.6000 738.4500 ;
	    RECT 198.6000 737.4000 199.8000 737.5500 ;
	    RECT 215.4000 737.4000 216.6000 737.5500 ;
	    RECT 227.4000 737.4000 228.6000 738.6000 ;
	    RECT 198.6000 736.2000 199.8000 736.5000 ;
	    RECT 172.8000 730.2000 175.8000 731.1000 ;
	    RECT 160.2000 723.3000 161.4000 727.5000 ;
	    RECT 162.6000 723.3000 163.8000 727.5000 ;
	    RECT 165.0000 723.3000 166.2000 729.3000 ;
	    RECT 167.4000 723.3000 168.6000 730.2000 ;
	    RECT 172.8000 729.3000 173.7000 730.2000 ;
	    RECT 169.8000 722.4000 171.0000 729.3000 ;
	    RECT 172.2000 728.4000 173.7000 729.3000 ;
	    RECT 172.2000 723.3000 173.4000 728.4000 ;
	    RECT 174.6000 723.3000 175.8000 729.3000 ;
	    RECT 193.8000 723.3000 195.0000 735.3000 ;
	    RECT 196.2000 734.1000 198.9000 735.3000 ;
	    RECT 197.7000 723.3000 198.9000 734.1000 ;
	    RECT 225.0000 723.3000 226.2000 729.3000 ;
	    RECT 227.4000 723.3000 228.6000 736.5000 ;
	    RECT 229.8000 734.4000 231.0000 735.6000 ;
	    RECT 229.8000 733.2000 231.0000 733.5000 ;
	    RECT 229.8000 723.3000 231.0000 729.3000 ;
	    RECT 244.2000 723.3000 245.4000 729.3000 ;
	    RECT 246.6000 723.3000 247.8000 739.5000 ;
	    RECT 268.2000 738.4500 269.4000 738.6000 ;
	    RECT 275.4000 738.4500 276.6000 738.6000 ;
	    RECT 268.2000 737.5500 276.6000 738.4500 ;
	    RECT 268.2000 737.4000 269.4000 737.5500 ;
	    RECT 275.4000 737.4000 276.6000 737.5500 ;
	    RECT 249.0000 735.4500 250.2000 735.6000 ;
	    RECT 265.8000 735.4500 267.0000 735.6000 ;
	    RECT 249.0000 734.5500 267.0000 735.4500 ;
	    RECT 249.0000 734.4000 250.2000 734.5500 ;
	    RECT 265.8000 734.4000 267.0000 734.5500 ;
	    RECT 265.8000 733.2000 267.0000 733.5000 ;
	    RECT 265.8000 723.3000 267.0000 729.3000 ;
	    RECT 268.2000 723.3000 269.4000 736.5000 ;
	    RECT 270.6000 723.3000 271.8000 729.3000 ;
	    RECT 282.6000 723.3000 283.8000 739.5000 ;
	    RECT 285.0000 723.3000 286.2000 729.3000 ;
	    RECT 299.4000 723.3000 300.6000 729.3000 ;
	    RECT 301.8000 723.3000 303.0000 739.5000 ;
	    RECT 316.2000 723.3000 317.4000 729.3000 ;
	    RECT 318.6000 723.3000 319.8000 739.5000 ;
	    RECT 349.8000 739.2000 351.0000 739.5000 ;
	    RECT 352.2000 737.4000 353.4000 738.6000 ;
	    RECT 354.9000 735.3000 355.8000 739.5000 ;
	    RECT 357.0000 737.4000 358.2000 738.6000 ;
	    RECT 349.8000 723.3000 351.0000 735.3000 ;
	    RECT 353.7000 723.3000 356.7000 735.3000 ;
	    RECT 359.4000 723.3000 360.6000 735.3000 ;
	    RECT 491.4000 731.1000 492.6000 739.5000 ;
	    RECT 505.5000 738.9000 508.5000 740.1000 ;
	    RECT 514.2000 738.9000 519.0000 740.1000 ;
	    RECT 522.6000 739.2000 523.8000 743.4000 ;
	    RECT 529.8000 742.8000 531.0000 743.7000 ;
	    RECT 529.8000 741.9000 532.5000 742.8000 ;
	    RECT 531.3000 740.1000 532.5000 741.9000 ;
	    RECT 537.0000 741.9000 538.2000 749.7000 ;
	    RECT 539.4000 744.0000 540.6000 749.7000 ;
	    RECT 541.8000 746.7000 543.0000 749.7000 ;
	    RECT 556.2000 746.7000 557.4000 749.7000 ;
	    RECT 556.2000 745.5000 557.4000 745.8000 ;
	    RECT 546.6000 744.4500 547.8000 744.6000 ;
	    RECT 556.2000 744.4500 557.4000 744.6000 ;
	    RECT 539.4000 742.8000 540.9000 744.0000 ;
	    RECT 546.6000 743.5500 557.4000 744.4500 ;
	    RECT 546.6000 743.4000 547.8000 743.5500 ;
	    RECT 556.2000 743.4000 557.4000 743.5500 ;
	    RECT 537.0000 741.0000 538.8000 741.9000 ;
	    RECT 531.3000 738.9000 537.0000 740.1000 ;
	    RECT 493.5000 738.0000 494.7000 738.3000 ;
	    RECT 493.5000 737.1000 500.1000 738.0000 ;
	    RECT 501.0000 737.4000 502.2000 738.6000 ;
	    RECT 527.4000 738.0000 528.6000 738.9000 ;
	    RECT 537.9000 738.0000 538.8000 741.0000 ;
	    RECT 503.1000 737.1000 528.6000 738.0000 ;
	    RECT 537.6000 737.1000 538.8000 738.0000 ;
	    RECT 535.5000 736.2000 536.7000 736.5000 ;
	    RECT 496.2000 734.4000 497.4000 735.6000 ;
	    RECT 498.3000 735.3000 536.7000 736.2000 ;
	    RECT 501.3000 735.0000 502.5000 735.3000 ;
	    RECT 537.6000 734.4000 538.5000 737.1000 ;
	    RECT 539.7000 736.2000 540.9000 742.8000 ;
	    RECT 558.6000 742.5000 559.8000 749.7000 ;
	    RECT 578.7000 744.6000 579.9000 749.7000 ;
	    RECT 578.7000 743.7000 581.4000 744.6000 ;
	    RECT 582.6000 743.7000 583.8000 749.7000 ;
	    RECT 594.6000 746.7000 595.8000 749.7000 ;
	    RECT 594.6000 745.5000 595.8000 745.8000 ;
	    RECT 592.2000 744.4500 593.4000 744.6000 ;
	    RECT 594.6000 744.4500 595.8000 744.6000 ;
	    RECT 558.6000 741.4500 559.8000 741.6000 ;
	    RECT 577.8000 741.4500 579.0000 741.6000 ;
	    RECT 558.6000 740.5500 579.0000 741.4500 ;
	    RECT 558.6000 740.4000 559.8000 740.5500 ;
	    RECT 577.8000 740.4000 579.0000 740.5500 ;
	    RECT 580.2000 739.5000 581.4000 743.7000 ;
	    RECT 592.2000 743.5500 595.8000 744.4500 ;
	    RECT 592.2000 743.4000 593.4000 743.5500 ;
	    RECT 594.6000 743.4000 595.8000 743.5500 ;
	    RECT 582.6000 742.5000 583.8000 742.8000 ;
	    RECT 597.0000 742.5000 598.2000 749.7000 ;
	    RECT 616.2000 743.7000 617.4000 749.7000 ;
	    RECT 620.1000 744.6000 621.3000 749.7000 ;
	    RECT 618.6000 743.7000 621.3000 744.6000 ;
	    RECT 616.2000 742.5000 617.4000 742.8000 ;
	    RECT 582.6000 741.4500 583.8000 741.6000 ;
	    RECT 592.2000 741.4500 593.4000 741.6000 ;
	    RECT 582.6000 740.5500 593.4000 741.4500 ;
	    RECT 582.6000 740.4000 583.8000 740.5500 ;
	    RECT 592.2000 740.4000 593.4000 740.5500 ;
	    RECT 597.0000 741.4500 598.2000 741.6000 ;
	    RECT 616.2000 741.4500 617.4000 741.6000 ;
	    RECT 597.0000 740.5500 617.4000 741.4500 ;
	    RECT 597.0000 740.4000 598.2000 740.5500 ;
	    RECT 616.2000 740.4000 617.4000 740.5500 ;
	    RECT 618.6000 739.5000 619.8000 743.7000 ;
	    RECT 646.8000 741.3000 648.0000 749.7000 ;
	    RECT 645.3000 740.7000 648.0000 741.3000 ;
	    RECT 652.2000 740.7000 653.4000 749.7000 ;
	    RECT 673.8000 746.7000 675.0000 749.7000 ;
	    RECT 673.8000 745.5000 675.0000 745.8000 ;
	    RECT 673.8000 743.4000 675.0000 744.6000 ;
	    RECT 676.2000 742.5000 677.4000 749.7000 ;
	    RECT 696.3000 744.6000 697.5000 749.7000 ;
	    RECT 696.3000 743.7000 699.0000 744.6000 ;
	    RECT 700.2000 743.7000 701.4000 749.7000 ;
	    RECT 714.6000 746.7000 715.8000 749.7000 ;
	    RECT 714.6000 745.5000 715.8000 745.8000 ;
	    RECT 712.2000 744.4500 713.4000 744.6000 ;
	    RECT 714.6000 744.4500 715.8000 744.6000 ;
	    RECT 654.6000 741.4500 655.8000 741.6000 ;
	    RECT 676.2000 741.4500 677.4000 741.6000 ;
	    RECT 645.3000 740.4000 647.7000 740.7000 ;
	    RECT 654.6000 740.5500 677.4000 741.4500 ;
	    RECT 654.6000 740.4000 655.8000 740.5500 ;
	    RECT 676.2000 740.4000 677.4000 740.5500 ;
	    RECT 505.8000 734.1000 507.0000 734.4000 ;
	    RECT 498.9000 733.5000 507.0000 734.1000 ;
	    RECT 497.7000 733.2000 507.0000 733.5000 ;
	    RECT 508.5000 733.5000 521.4000 734.4000 ;
	    RECT 493.8000 732.0000 496.2000 733.2000 ;
	    RECT 497.7000 732.3000 499.8000 733.2000 ;
	    RECT 508.5000 732.3000 509.4000 733.5000 ;
	    RECT 520.2000 733.2000 521.4000 733.5000 ;
	    RECT 525.0000 733.5000 538.5000 734.4000 ;
	    RECT 539.4000 735.0000 540.9000 736.2000 ;
	    RECT 539.4000 733.5000 540.6000 735.0000 ;
	    RECT 525.0000 733.2000 526.2000 733.5000 ;
	    RECT 495.3000 731.4000 496.2000 732.0000 ;
	    RECT 500.7000 731.4000 509.4000 732.3000 ;
	    RECT 510.3000 731.4000 514.2000 732.6000 ;
	    RECT 491.4000 730.2000 494.4000 731.1000 ;
	    RECT 495.3000 730.2000 501.6000 731.4000 ;
	    RECT 493.5000 729.3000 494.4000 730.2000 ;
	    RECT 491.4000 723.3000 492.6000 729.3000 ;
	    RECT 493.5000 728.4000 495.0000 729.3000 ;
	    RECT 493.8000 723.3000 495.0000 728.4000 ;
	    RECT 496.2000 722.4000 497.4000 729.3000 ;
	    RECT 498.6000 723.3000 499.8000 730.2000 ;
	    RECT 501.0000 723.3000 502.2000 729.3000 ;
	    RECT 503.4000 723.3000 504.6000 727.5000 ;
	    RECT 505.8000 723.3000 507.0000 727.5000 ;
	    RECT 508.2000 723.3000 509.4000 730.5000 ;
	    RECT 510.6000 723.3000 511.8000 729.3000 ;
	    RECT 513.0000 723.3000 514.2000 730.5000 ;
	    RECT 515.4000 723.3000 516.6000 729.3000 ;
	    RECT 517.8000 723.3000 519.0000 732.6000 ;
	    RECT 529.8000 731.4000 533.7000 732.6000 ;
	    RECT 522.6000 730.2000 528.9000 731.4000 ;
	    RECT 520.2000 723.3000 521.4000 727.5000 ;
	    RECT 522.6000 723.3000 523.8000 727.5000 ;
	    RECT 525.0000 723.3000 526.2000 727.5000 ;
	    RECT 527.4000 723.3000 528.6000 729.3000 ;
	    RECT 529.8000 723.3000 531.0000 731.4000 ;
	    RECT 537.6000 731.1000 538.5000 733.5000 ;
	    RECT 539.4000 731.4000 540.6000 732.6000 ;
	    RECT 534.6000 730.2000 538.5000 731.1000 ;
	    RECT 532.2000 723.3000 533.4000 729.3000 ;
	    RECT 534.6000 723.3000 535.8000 730.2000 ;
	    RECT 537.0000 723.3000 538.2000 729.3000 ;
	    RECT 539.4000 723.3000 540.6000 730.5000 ;
	    RECT 541.8000 723.3000 543.0000 729.3000 ;
	    RECT 556.2000 723.3000 557.4000 729.3000 ;
	    RECT 558.6000 723.3000 559.8000 739.5000 ;
	    RECT 580.2000 738.4500 581.4000 738.6000 ;
	    RECT 594.6000 738.4500 595.8000 738.6000 ;
	    RECT 580.2000 737.5500 595.8000 738.4500 ;
	    RECT 580.2000 737.4000 581.4000 737.5500 ;
	    RECT 594.6000 737.4000 595.8000 737.5500 ;
	    RECT 568.2000 735.4500 569.4000 735.6000 ;
	    RECT 577.8000 735.4500 579.0000 735.6000 ;
	    RECT 568.2000 734.5500 579.0000 735.4500 ;
	    RECT 568.2000 734.4000 569.4000 734.5500 ;
	    RECT 577.8000 734.4000 579.0000 734.5500 ;
	    RECT 577.8000 733.2000 579.0000 733.5000 ;
	    RECT 577.8000 723.3000 579.0000 729.3000 ;
	    RECT 580.2000 723.3000 581.4000 736.5000 ;
	    RECT 582.6000 723.3000 583.8000 729.3000 ;
	    RECT 594.6000 723.3000 595.8000 729.3000 ;
	    RECT 597.0000 723.3000 598.2000 739.5000 ;
	    RECT 618.6000 738.4500 619.8000 738.6000 ;
	    RECT 637.8000 738.4500 639.0000 738.6000 ;
	    RECT 618.6000 737.5500 639.0000 738.4500 ;
	    RECT 618.6000 737.4000 619.8000 737.5500 ;
	    RECT 637.8000 737.4000 639.0000 737.5500 ;
	    RECT 645.3000 736.5000 646.2000 740.4000 ;
	    RECT 697.8000 739.5000 699.0000 743.7000 ;
	    RECT 712.2000 743.5500 715.8000 744.4500 ;
	    RECT 712.2000 743.4000 713.4000 743.5500 ;
	    RECT 714.6000 743.4000 715.8000 743.5500 ;
	    RECT 700.2000 742.5000 701.4000 742.8000 ;
	    RECT 717.0000 742.5000 718.2000 749.7000 ;
	    RECT 700.2000 741.4500 701.4000 741.6000 ;
	    RECT 714.6000 741.4500 715.8000 741.6000 ;
	    RECT 700.2000 740.5500 715.8000 741.4500 ;
	    RECT 700.2000 740.4000 701.4000 740.5500 ;
	    RECT 714.6000 740.4000 715.8000 740.5500 ;
	    RECT 717.0000 741.4500 718.2000 741.6000 ;
	    RECT 733.8000 741.4500 735.0000 741.6000 ;
	    RECT 717.0000 740.5500 735.0000 741.4500 ;
	    RECT 741.0000 740.7000 742.2000 749.7000 ;
	    RECT 746.4000 741.3000 747.6000 749.7000 ;
	    RECT 762.6000 742.5000 763.8000 749.7000 ;
	    RECT 765.0000 746.7000 766.2000 749.7000 ;
	    RECT 765.0000 745.5000 766.2000 745.8000 ;
	    RECT 765.0000 744.4500 766.2000 744.6000 ;
	    RECT 786.6000 744.4500 787.8000 744.6000 ;
	    RECT 765.0000 743.5500 787.8000 744.4500 ;
	    RECT 765.0000 743.4000 766.2000 743.5500 ;
	    RECT 786.6000 743.4000 787.8000 743.5500 ;
	    RECT 750.6000 741.4500 751.8000 741.6000 ;
	    RECT 762.6000 741.4500 763.8000 741.6000 ;
	    RECT 746.4000 740.7000 749.1000 741.3000 ;
	    RECT 717.0000 740.4000 718.2000 740.5500 ;
	    RECT 733.8000 740.4000 735.0000 740.5500 ;
	    RECT 746.7000 740.4000 749.1000 740.7000 ;
	    RECT 750.6000 740.5500 763.8000 741.4500 ;
	    RECT 793.2000 741.3000 794.4000 749.7000 ;
	    RECT 750.6000 740.4000 751.8000 740.5500 ;
	    RECT 762.6000 740.4000 763.8000 740.5500 ;
	    RECT 791.7000 740.7000 794.4000 741.3000 ;
	    RECT 798.6000 740.7000 799.8000 749.7000 ;
	    RECT 827.4000 744.0000 828.6000 749.7000 ;
	    RECT 829.8000 744.9000 831.0000 749.7000 ;
	    RECT 832.2000 748.8000 838.2000 749.7000 ;
	    RECT 832.2000 744.0000 833.4000 748.8000 ;
	    RECT 827.4000 743.7000 833.4000 744.0000 ;
	    RECT 834.6000 743.7000 835.8000 747.9000 ;
	    RECT 837.0000 743.7000 838.2000 748.8000 ;
	    RECT 857.1000 744.6000 858.3000 749.7000 ;
	    RECT 857.1000 743.7000 859.8000 744.6000 ;
	    RECT 861.0000 743.7000 862.2000 749.7000 ;
	    RECT 875.4000 746.7000 876.6000 749.7000 ;
	    RECT 875.4000 745.5000 876.6000 745.8000 ;
	    RECT 827.7000 743.1000 833.1000 743.7000 ;
	    RECT 791.7000 740.4000 794.1000 740.7000 ;
	    RECT 827.4000 740.4000 828.6000 741.6000 ;
	    RECT 829.5000 740.7000 829.8000 742.2000 ;
	    RECT 834.9000 741.6000 835.8000 743.7000 ;
	    RECT 832.2000 740.4000 833.4000 741.6000 ;
	    RECT 834.3000 740.7000 835.8000 741.6000 ;
	    RECT 837.0000 740.4000 838.2000 741.6000 ;
	    RECT 648.6000 737.4000 648.9000 738.6000 ;
	    RECT 649.8000 737.4000 651.0000 738.6000 ;
	    RECT 652.2000 736.5000 653.4000 736.8000 ;
	    RECT 616.2000 723.3000 617.4000 729.3000 ;
	    RECT 618.6000 723.3000 619.8000 736.5000 ;
	    RECT 621.0000 734.4000 622.2000 735.6000 ;
	    RECT 645.0000 734.4000 646.2000 735.6000 ;
	    RECT 652.2000 734.4000 653.4000 735.6000 ;
	    RECT 647.4000 733.5000 648.6000 733.8000 ;
	    RECT 621.0000 733.2000 622.2000 733.5000 ;
	    RECT 645.3000 730.5000 646.2000 733.5000 ;
	    RECT 647.4000 732.4500 648.6000 732.6000 ;
	    RECT 654.6000 732.4500 655.8000 732.6000 ;
	    RECT 647.4000 731.5500 655.8000 732.4500 ;
	    RECT 647.4000 731.4000 648.6000 731.5500 ;
	    RECT 654.6000 731.4000 655.8000 731.5500 ;
	    RECT 645.3000 729.6000 650.7000 730.5000 ;
	    RECT 645.3000 729.3000 646.2000 729.6000 ;
	    RECT 621.0000 723.3000 622.2000 729.3000 ;
	    RECT 645.0000 723.3000 646.2000 729.3000 ;
	    RECT 649.8000 729.3000 650.7000 729.6000 ;
	    RECT 647.4000 723.3000 648.6000 728.7000 ;
	    RECT 649.8000 723.3000 651.0000 729.3000 ;
	    RECT 652.2000 723.3000 653.4000 729.3000 ;
	    RECT 673.8000 723.3000 675.0000 729.3000 ;
	    RECT 676.2000 723.3000 677.4000 739.5000 ;
	    RECT 693.0000 738.4500 694.2000 738.6000 ;
	    RECT 697.8000 738.4500 699.0000 738.6000 ;
	    RECT 693.0000 737.5500 699.0000 738.4500 ;
	    RECT 693.0000 737.4000 694.2000 737.5500 ;
	    RECT 697.8000 737.4000 699.0000 737.5500 ;
	    RECT 690.6000 735.4500 691.8000 735.6000 ;
	    RECT 695.4000 735.4500 696.6000 735.6000 ;
	    RECT 690.6000 734.5500 696.6000 735.4500 ;
	    RECT 690.6000 734.4000 691.8000 734.5500 ;
	    RECT 695.4000 734.4000 696.6000 734.5500 ;
	    RECT 695.4000 733.2000 696.6000 733.5000 ;
	    RECT 695.4000 723.3000 696.6000 729.3000 ;
	    RECT 697.8000 723.3000 699.0000 736.5000 ;
	    RECT 700.2000 723.3000 701.4000 729.3000 ;
	    RECT 714.6000 723.3000 715.8000 729.3000 ;
	    RECT 717.0000 723.3000 718.2000 739.5000 ;
	    RECT 743.4000 737.4000 744.6000 738.6000 ;
	    RECT 745.5000 737.4000 745.8000 738.6000 ;
	    RECT 741.0000 736.5000 742.2000 736.8000 ;
	    RECT 748.2000 736.5000 749.1000 740.4000 ;
	    RECT 733.8000 735.4500 735.0000 735.6000 ;
	    RECT 741.0000 735.4500 742.2000 735.6000 ;
	    RECT 733.8000 734.5500 742.2000 735.4500 ;
	    RECT 733.8000 734.4000 735.0000 734.5500 ;
	    RECT 741.0000 734.4000 742.2000 734.5500 ;
	    RECT 748.2000 734.4000 749.4000 735.6000 ;
	    RECT 745.8000 733.5000 747.0000 733.8000 ;
	    RECT 745.8000 731.4000 747.0000 732.6000 ;
	    RECT 748.2000 730.5000 749.1000 733.5000 ;
	    RECT 743.7000 729.6000 749.1000 730.5000 ;
	    RECT 743.7000 729.3000 744.6000 729.6000 ;
	    RECT 741.0000 723.3000 742.2000 729.3000 ;
	    RECT 743.4000 723.3000 744.6000 729.3000 ;
	    RECT 748.2000 729.3000 749.1000 729.6000 ;
	    RECT 745.8000 723.3000 747.0000 728.7000 ;
	    RECT 748.2000 723.3000 749.4000 729.3000 ;
	    RECT 762.6000 723.3000 763.8000 739.5000 ;
	    RECT 791.7000 736.5000 792.6000 740.4000 ;
	    RECT 829.8000 739.5000 831.0000 739.8000 ;
	    RECT 834.6000 739.5000 835.8000 739.8000 ;
	    RECT 858.6000 739.5000 859.8000 743.7000 ;
	    RECT 875.4000 743.4000 876.6000 744.6000 ;
	    RECT 861.0000 742.5000 862.2000 742.8000 ;
	    RECT 877.8000 742.5000 879.0000 749.7000 ;
	    RECT 889.8000 747.4500 891.0000 747.6000 ;
	    RECT 1005.0000 747.4500 1006.2000 747.6000 ;
	    RECT 889.8000 746.5500 1006.2000 747.4500 ;
	    RECT 1012.2000 746.7000 1013.4000 749.7000 ;
	    RECT 889.8000 746.4000 891.0000 746.5500 ;
	    RECT 1005.0000 746.4000 1006.2000 746.5500 ;
	    RECT 1014.6000 744.0000 1015.8000 749.7000 ;
	    RECT 1014.3000 742.8000 1015.8000 744.0000 ;
	    RECT 861.0000 740.4000 862.2000 741.6000 ;
	    RECT 877.8000 741.4500 879.0000 741.6000 ;
	    RECT 885.0000 741.4500 886.2000 741.6000 ;
	    RECT 877.8000 740.5500 886.2000 741.4500 ;
	    RECT 877.8000 740.4000 879.0000 740.5500 ;
	    RECT 885.0000 740.4000 886.2000 740.5500 ;
	    RECT 795.0000 737.4000 795.3000 738.6000 ;
	    RECT 796.2000 737.4000 797.4000 738.6000 ;
	    RECT 820.2000 738.4500 821.4000 738.6000 ;
	    RECT 829.8000 738.4500 831.0000 738.6000 ;
	    RECT 820.2000 737.5500 831.0000 738.4500 ;
	    RECT 820.2000 737.4000 821.4000 737.5500 ;
	    RECT 829.8000 737.4000 831.0000 737.5500 ;
	    RECT 798.6000 736.5000 799.8000 736.8000 ;
	    RECT 791.4000 734.4000 792.6000 735.6000 ;
	    RECT 798.6000 735.4500 799.8000 735.6000 ;
	    RECT 805.8000 735.4500 807.0000 735.6000 ;
	    RECT 798.6000 734.5500 807.0000 735.4500 ;
	    RECT 832.2000 735.3000 833.1000 739.5000 ;
	    RECT 837.0000 739.2000 838.2000 739.5000 ;
	    RECT 834.6000 737.4000 835.8000 738.6000 ;
	    RECT 858.6000 738.4500 859.8000 738.6000 ;
	    RECT 873.0000 738.4500 874.2000 738.6000 ;
	    RECT 858.6000 737.5500 874.2000 738.4500 ;
	    RECT 858.6000 737.4000 859.8000 737.5500 ;
	    RECT 873.0000 737.4000 874.2000 737.5500 ;
	    RECT 798.6000 734.4000 799.8000 734.5500 ;
	    RECT 805.8000 734.4000 807.0000 734.5500 ;
	    RECT 793.8000 733.5000 795.0000 733.8000 ;
	    RECT 791.7000 730.5000 792.6000 733.5000 ;
	    RECT 793.8000 731.4000 795.0000 732.6000 ;
	    RECT 791.7000 729.6000 797.1000 730.5000 ;
	    RECT 791.7000 729.3000 792.6000 729.6000 ;
	    RECT 765.0000 723.3000 766.2000 729.3000 ;
	    RECT 791.4000 723.3000 792.6000 729.3000 ;
	    RECT 796.2000 729.3000 797.1000 729.6000 ;
	    RECT 793.8000 723.3000 795.0000 728.7000 ;
	    RECT 796.2000 723.3000 797.4000 729.3000 ;
	    RECT 798.6000 723.3000 799.8000 729.3000 ;
	    RECT 827.4000 723.3000 828.6000 735.3000 ;
	    RECT 831.3000 723.3000 834.3000 735.3000 ;
	    RECT 837.0000 723.3000 838.2000 735.3000 ;
	    RECT 856.2000 734.4000 857.4000 735.6000 ;
	    RECT 856.2000 733.2000 857.4000 733.5000 ;
	    RECT 856.2000 723.3000 857.4000 729.3000 ;
	    RECT 858.6000 723.3000 859.8000 736.5000 ;
	    RECT 861.0000 723.3000 862.2000 729.3000 ;
	    RECT 875.4000 723.3000 876.6000 729.3000 ;
	    RECT 877.8000 723.3000 879.0000 739.5000 ;
	    RECT 930.6000 738.4500 931.8000 738.6000 ;
	    RECT 1012.2000 738.4500 1013.4000 738.6000 ;
	    RECT 930.6000 737.5500 1013.4000 738.4500 ;
	    RECT 930.6000 737.4000 931.8000 737.5500 ;
	    RECT 1012.2000 737.4000 1013.4000 737.5500 ;
	    RECT 1014.3000 736.2000 1015.5000 742.8000 ;
	    RECT 1017.0000 741.9000 1018.2000 749.7000 ;
	    RECT 1021.8000 743.7000 1023.0000 749.7000 ;
	    RECT 1026.6000 744.9000 1027.8000 749.7000 ;
	    RECT 1029.0000 745.5000 1030.2001 749.7000 ;
	    RECT 1031.4000 745.5000 1032.6000 749.7000 ;
	    RECT 1033.8000 745.5000 1035.0000 749.7000 ;
	    RECT 1036.2001 745.5000 1037.4000 749.7000 ;
	    RECT 1038.6000 746.7000 1039.8000 749.7000 ;
	    RECT 1041.0000 745.5000 1042.2001 749.7000 ;
	    RECT 1043.4000 746.7000 1044.6000 749.7000 ;
	    RECT 1045.8000 745.5000 1047.0000 749.7000 ;
	    RECT 1048.2001 745.5000 1049.4000 749.7000 ;
	    RECT 1050.6000 745.5000 1051.8000 749.7000 ;
	    RECT 1024.2001 743.7000 1027.8000 744.9000 ;
	    RECT 1053.0000 744.9000 1054.2001 749.7000 ;
	    RECT 1024.2001 742.8000 1025.4000 743.7000 ;
	    RECT 1016.4000 741.0000 1018.2000 741.9000 ;
	    RECT 1022.7000 741.9000 1025.4000 742.8000 ;
	    RECT 1031.4000 743.4000 1032.9000 744.6000 ;
	    RECT 1037.4000 743.4000 1037.7001 744.6000 ;
	    RECT 1038.6000 743.4000 1039.8000 744.6000 ;
	    RECT 1041.0000 743.7000 1047.9000 744.6000 ;
	    RECT 1053.0000 743.7000 1056.9000 744.9000 ;
	    RECT 1057.8000 743.7000 1059.0000 749.7000 ;
	    RECT 1041.0000 743.4000 1042.2001 743.7000 ;
	    RECT 1016.4000 738.0000 1017.3000 741.0000 ;
	    RECT 1022.7000 740.1000 1023.9000 741.9000 ;
	    RECT 1018.2000 738.9000 1023.9000 740.1000 ;
	    RECT 1031.4000 739.2000 1032.6000 743.4000 ;
	    RECT 1043.4000 742.5000 1044.6000 742.8000 ;
	    RECT 1041.0000 742.2000 1042.2001 742.5000 ;
	    RECT 1035.6000 741.3000 1042.2001 742.2000 ;
	    RECT 1035.6000 741.0000 1036.8000 741.3000 ;
	    RECT 1043.4000 740.4000 1044.6000 741.6000 ;
	    RECT 1046.7001 740.1000 1047.9000 743.7000 ;
	    RECT 1055.7001 742.8000 1056.9000 743.7000 ;
	    RECT 1055.7001 741.6000 1060.2001 742.8000 ;
	    RECT 1062.6000 740.7000 1063.8000 749.7000 ;
	    RECT 1082.7001 744.6000 1083.9000 749.7000 ;
	    RECT 1082.7001 743.7000 1085.4000 744.6000 ;
	    RECT 1086.6000 743.7000 1087.8000 749.7000 ;
	    RECT 1218.6000 746.7000 1219.8000 749.7000 ;
	    RECT 1221.0000 744.0000 1222.2001 749.7000 ;
	    RECT 1036.2001 738.9000 1041.0000 740.1000 ;
	    RECT 1046.7001 738.9000 1049.7001 740.1000 ;
	    RECT 1050.6000 739.5000 1063.8000 740.7000 ;
	    RECT 1084.2001 739.5000 1085.4000 743.7000 ;
	    RECT 1220.7001 742.8000 1222.2001 744.0000 ;
	    RECT 1086.6000 742.5000 1087.8000 742.8000 ;
	    RECT 1086.6000 740.4000 1087.8000 741.6000 ;
	    RECT 1026.6000 738.0000 1027.8000 738.9000 ;
	    RECT 1016.4000 737.1000 1017.6000 738.0000 ;
	    RECT 1026.6000 737.1000 1052.1000 738.0000 ;
	    RECT 1053.0000 737.4000 1054.2001 738.6000 ;
	    RECT 1060.5000 738.0000 1061.7001 738.3000 ;
	    RECT 1055.1000 737.1000 1061.7001 738.0000 ;
	    RECT 882.6000 735.4500 883.8000 735.6000 ;
	    RECT 971.4000 735.4500 972.6000 735.6000 ;
	    RECT 882.6000 734.5500 972.6000 735.4500 ;
	    RECT 1014.3000 735.0000 1015.8000 736.2000 ;
	    RECT 882.6000 734.4000 883.8000 734.5500 ;
	    RECT 971.4000 734.4000 972.6000 734.5500 ;
	    RECT 1014.6000 733.5000 1015.8000 735.0000 ;
	    RECT 1016.7000 734.4000 1017.6000 737.1000 ;
	    RECT 1018.5000 736.2000 1019.7000 736.5000 ;
	    RECT 1018.5000 735.3000 1056.9000 736.2000 ;
	    RECT 1052.7001 735.0000 1053.9000 735.3000 ;
	    RECT 1057.8000 734.4000 1059.0000 735.6000 ;
	    RECT 1016.7000 733.5000 1030.2001 734.4000 ;
	    RECT 925.8000 732.4500 927.0000 732.6000 ;
	    RECT 973.8000 732.4500 975.0000 732.6000 ;
	    RECT 1014.6000 732.4500 1015.8000 732.6000 ;
	    RECT 925.8000 731.5500 1015.8000 732.4500 ;
	    RECT 925.8000 731.4000 927.0000 731.5500 ;
	    RECT 973.8000 731.4000 975.0000 731.5500 ;
	    RECT 1014.6000 731.4000 1015.8000 731.5500 ;
	    RECT 1016.7000 731.1000 1017.6000 733.5000 ;
	    RECT 1029.0000 733.2000 1030.2001 733.5000 ;
	    RECT 1033.8000 733.5000 1046.7001 734.4000 ;
	    RECT 1033.8000 733.2000 1035.0000 733.5000 ;
	    RECT 1021.5000 731.4000 1025.4000 732.6000 ;
	    RECT 889.8000 729.4500 891.0000 729.6000 ;
	    RECT 1007.4000 729.4500 1008.6000 729.6000 ;
	    RECT 889.8000 728.5500 1008.6000 729.4500 ;
	    RECT 889.8000 728.4000 891.0000 728.5500 ;
	    RECT 1007.4000 728.4000 1008.6000 728.5500 ;
	    RECT 880.2000 726.4500 881.4000 726.6000 ;
	    RECT 949.8000 726.4500 951.0000 726.6000 ;
	    RECT 880.2000 725.5500 951.0000 726.4500 ;
	    RECT 880.2000 725.4000 881.4000 725.5500 ;
	    RECT 949.8000 725.4000 951.0000 725.5500 ;
	    RECT 1012.2000 723.3000 1013.4000 729.3000 ;
	    RECT 1014.6000 723.3000 1015.8000 730.5000 ;
	    RECT 1016.7000 730.2000 1020.6000 731.1000 ;
	    RECT 1017.0000 723.3000 1018.2000 729.3000 ;
	    RECT 1019.4000 723.3000 1020.6000 730.2000 ;
	    RECT 1021.8000 723.3000 1023.0000 729.3000 ;
	    RECT 1024.2001 723.3000 1025.4000 731.4000 ;
	    RECT 1026.3000 730.2000 1032.6000 731.4000 ;
	    RECT 1026.6000 723.3000 1027.8000 729.3000 ;
	    RECT 1029.0000 723.3000 1030.2001 727.5000 ;
	    RECT 1031.4000 723.3000 1032.6000 727.5000 ;
	    RECT 1033.8000 723.3000 1035.0000 727.5000 ;
	    RECT 1036.2001 723.3000 1037.4000 732.6000 ;
	    RECT 1041.0000 731.4000 1044.9000 732.6000 ;
	    RECT 1045.8000 732.3000 1046.7001 733.5000 ;
	    RECT 1048.2001 734.1000 1049.4000 734.4000 ;
	    RECT 1048.2001 733.5000 1056.3000 734.1000 ;
	    RECT 1048.2001 733.2000 1057.5000 733.5000 ;
	    RECT 1055.4000 732.3000 1057.5000 733.2000 ;
	    RECT 1045.8000 731.4000 1054.5000 732.3000 ;
	    RECT 1059.0000 732.0000 1061.4000 733.2000 ;
	    RECT 1059.0000 731.4000 1059.9000 732.0000 ;
	    RECT 1038.6000 723.3000 1039.8000 729.3000 ;
	    RECT 1041.0000 723.3000 1042.2001 730.5000 ;
	    RECT 1043.4000 723.3000 1044.6000 729.3000 ;
	    RECT 1045.8000 723.3000 1047.0000 730.5000 ;
	    RECT 1053.6000 730.2000 1059.9000 731.4000 ;
	    RECT 1062.6000 731.1000 1063.8000 739.5000 ;
	    RECT 1069.8000 738.4500 1071.0000 738.6000 ;
	    RECT 1084.2001 738.4500 1085.4000 738.6000 ;
	    RECT 1069.8000 737.5500 1085.4000 738.4500 ;
	    RECT 1069.8000 737.4000 1071.0000 737.5500 ;
	    RECT 1084.2001 737.4000 1085.4000 737.5500 ;
	    RECT 1081.8000 734.4000 1083.0000 735.6000 ;
	    RECT 1081.8000 733.2000 1083.0000 733.5000 ;
	    RECT 1060.8000 730.2000 1063.8000 731.1000 ;
	    RECT 1048.2001 723.3000 1049.4000 727.5000 ;
	    RECT 1050.6000 723.3000 1051.8000 727.5000 ;
	    RECT 1053.0000 723.3000 1054.2001 729.3000 ;
	    RECT 1055.4000 723.3000 1056.6000 730.2000 ;
	    RECT 1060.8000 729.3000 1061.7001 730.2000 ;
	    RECT 1057.8000 722.4000 1059.0000 729.3000 ;
	    RECT 1060.2001 728.4000 1061.7001 729.3000 ;
	    RECT 1060.2001 723.3000 1061.4000 728.4000 ;
	    RECT 1062.6000 723.3000 1063.8000 729.3000 ;
	    RECT 1081.8000 723.3000 1083.0000 729.3000 ;
	    RECT 1084.2001 723.3000 1085.4000 736.5000 ;
	    RECT 1220.7001 736.2000 1221.9000 742.8000 ;
	    RECT 1223.4000 741.9000 1224.6000 749.7000 ;
	    RECT 1228.2001 743.7000 1229.4000 749.7000 ;
	    RECT 1233.0000 744.9000 1234.2001 749.7000 ;
	    RECT 1235.4000 745.5000 1236.6000 749.7000 ;
	    RECT 1237.8000 745.5000 1239.0000 749.7000 ;
	    RECT 1240.2001 745.5000 1241.4000 749.7000 ;
	    RECT 1242.6000 745.5000 1243.8000 749.7000 ;
	    RECT 1245.0000 746.7000 1246.2001 749.7000 ;
	    RECT 1247.4000 745.5000 1248.6000 749.7000 ;
	    RECT 1249.8000 746.7000 1251.0000 749.7000 ;
	    RECT 1252.2001 745.5000 1253.4000 749.7000 ;
	    RECT 1254.6000 745.5000 1255.8000 749.7000 ;
	    RECT 1257.0000 745.5000 1258.2001 749.7000 ;
	    RECT 1230.6000 743.7000 1234.2001 744.9000 ;
	    RECT 1259.4000 744.9000 1260.6000 749.7000 ;
	    RECT 1230.6000 742.8000 1231.8000 743.7000 ;
	    RECT 1222.8000 741.0000 1224.6000 741.9000 ;
	    RECT 1229.1000 741.9000 1231.8000 742.8000 ;
	    RECT 1237.8000 743.4000 1239.3000 744.6000 ;
	    RECT 1243.8000 743.4000 1244.1000 744.6000 ;
	    RECT 1245.0000 743.4000 1246.2001 744.6000 ;
	    RECT 1247.4000 743.7000 1254.3000 744.6000 ;
	    RECT 1259.4000 743.7000 1263.3000 744.9000 ;
	    RECT 1264.2001 743.7000 1265.4000 749.7000 ;
	    RECT 1247.4000 743.4000 1248.6000 743.7000 ;
	    RECT 1222.8000 738.0000 1223.7001 741.0000 ;
	    RECT 1229.1000 740.1000 1230.3000 741.9000 ;
	    RECT 1224.6000 738.9000 1230.3000 740.1000 ;
	    RECT 1237.8000 739.2000 1239.0000 743.4000 ;
	    RECT 1249.8000 742.5000 1251.0000 742.8000 ;
	    RECT 1247.4000 742.2000 1248.6000 742.5000 ;
	    RECT 1242.0000 741.3000 1248.6000 742.2000 ;
	    RECT 1242.0000 741.0000 1243.2001 741.3000 ;
	    RECT 1249.8000 740.4000 1251.0000 741.6000 ;
	    RECT 1253.1000 740.1000 1254.3000 743.7000 ;
	    RECT 1262.1000 742.8000 1263.3000 743.7000 ;
	    RECT 1262.1000 741.6000 1266.6000 742.8000 ;
	    RECT 1269.0000 740.7000 1270.2001 749.7000 ;
	    RECT 1293.0000 743.7000 1294.2001 749.7000 ;
	    RECT 1295.4000 744.0000 1296.6000 749.7000 ;
	    RECT 1297.8000 744.9000 1299.0000 749.7000 ;
	    RECT 1300.2001 744.0000 1301.4000 749.7000 ;
	    RECT 1295.4000 743.7000 1301.4000 744.0000 ;
	    RECT 1326.6000 743.7000 1327.8000 749.7000 ;
	    RECT 1329.0000 744.0000 1330.2001 749.7000 ;
	    RECT 1331.4000 744.9000 1332.6000 749.7000 ;
	    RECT 1333.8000 744.0000 1335.0000 749.7000 ;
	    RECT 1329.0000 743.7000 1335.0000 744.0000 ;
	    RECT 1365.0000 743.7000 1366.2001 749.7000 ;
	    RECT 1367.4000 744.0000 1368.6000 749.7000 ;
	    RECT 1369.8000 744.9000 1371.0000 749.7000 ;
	    RECT 1372.2001 744.0000 1373.4000 749.7000 ;
	    RECT 1367.4000 743.7000 1373.4000 744.0000 ;
	    RECT 1293.3000 742.5000 1294.2001 743.7000 ;
	    RECT 1295.7001 743.1000 1301.1000 743.7000 ;
	    RECT 1326.9000 742.5000 1327.8000 743.7000 ;
	    RECT 1329.3000 743.1000 1334.7001 743.7000 ;
	    RECT 1365.3000 742.5000 1366.2001 743.7000 ;
	    RECT 1367.7001 743.1000 1373.1000 743.7000 ;
	    RECT 1384.2001 742.5000 1385.4000 749.7000 ;
	    RECT 1386.6000 746.7000 1387.8000 749.7000 ;
	    RECT 1386.6000 745.5000 1387.8000 745.8000 ;
	    RECT 1386.6000 743.4000 1387.8000 744.6000 ;
	    RECT 1410.6000 743.7000 1411.8000 749.7000 ;
	    RECT 1413.0000 744.0000 1414.2001 749.7000 ;
	    RECT 1415.4000 744.9000 1416.6000 749.7000 ;
	    RECT 1417.8000 744.0000 1419.0000 749.7000 ;
	    RECT 1432.2001 746.7000 1433.4000 749.7000 ;
	    RECT 1432.2001 745.5000 1433.4000 745.8000 ;
	    RECT 1413.0000 743.7000 1419.0000 744.0000 ;
	    RECT 1410.9000 742.5000 1411.8000 743.7000 ;
	    RECT 1413.3000 743.1000 1418.7001 743.7000 ;
	    RECT 1432.2001 743.4000 1433.4000 744.6000 ;
	    RECT 1434.6000 742.5000 1435.8000 749.7000 ;
	    RECT 1453.8000 743.7000 1455.0000 749.7000 ;
	    RECT 1457.7001 744.6000 1458.9000 749.7000 ;
	    RECT 1456.2001 743.7000 1458.9000 744.6000 ;
	    RECT 1485.0000 744.0000 1486.2001 749.7000 ;
	    RECT 1487.4000 744.9000 1488.6000 749.7000 ;
	    RECT 1489.8000 744.0000 1491.0000 749.7000 ;
	    RECT 1485.0000 743.7000 1491.0000 744.0000 ;
	    RECT 1492.2001 743.7000 1493.4000 749.7000 ;
	    RECT 1517.1000 743.7000 1518.3000 749.7000 ;
	    RECT 1521.0000 743.7000 1522.2001 749.7000 ;
	    RECT 1523.4000 746.7000 1524.6000 749.7000 ;
	    RECT 1523.1000 745.5000 1524.3000 745.8000 ;
	    RECT 1453.8000 742.5000 1455.0000 742.8000 ;
	    RECT 1242.6000 738.9000 1247.4000 740.1000 ;
	    RECT 1253.1000 738.9000 1256.1000 740.1000 ;
	    RECT 1257.0000 739.5000 1270.2001 740.7000 ;
	    RECT 1288.2001 741.4500 1289.4000 741.6000 ;
	    RECT 1293.0000 741.4500 1294.2001 741.6000 ;
	    RECT 1288.2001 740.5500 1294.2001 741.4500 ;
	    RECT 1288.2001 740.4000 1289.4000 740.5500 ;
	    RECT 1293.0000 740.4000 1294.2001 740.5500 ;
	    RECT 1295.1000 740.4000 1296.9000 741.6000 ;
	    RECT 1299.0000 740.7000 1299.3000 742.2000 ;
	    RECT 1300.2001 741.4500 1301.4000 741.6000 ;
	    RECT 1312.2001 741.4500 1313.4000 741.6000 ;
	    RECT 1300.2001 740.5500 1313.4000 741.4500 ;
	    RECT 1300.2001 740.4000 1301.4000 740.5500 ;
	    RECT 1312.2001 740.4000 1313.4000 740.5500 ;
	    RECT 1317.0000 741.4500 1318.2001 741.6000 ;
	    RECT 1326.6000 741.4500 1327.8000 741.6000 ;
	    RECT 1317.0000 740.5500 1327.8000 741.4500 ;
	    RECT 1317.0000 740.4000 1318.2001 740.5500 ;
	    RECT 1326.6000 740.4000 1327.8000 740.5500 ;
	    RECT 1328.7001 740.4000 1330.5000 741.6000 ;
	    RECT 1332.6000 740.7000 1332.9000 742.2000 ;
	    RECT 1333.8000 740.4000 1335.0000 741.6000 ;
	    RECT 1343.4000 741.4500 1344.6000 741.6000 ;
	    RECT 1365.0000 741.4500 1366.2001 741.6000 ;
	    RECT 1343.4000 740.5500 1366.2001 741.4500 ;
	    RECT 1343.4000 740.4000 1344.6000 740.5500 ;
	    RECT 1365.0000 740.4000 1366.2001 740.5500 ;
	    RECT 1367.1000 740.4000 1368.9000 741.6000 ;
	    RECT 1371.0000 740.7000 1371.3000 742.2000 ;
	    RECT 1372.2001 741.4500 1373.4000 741.6000 ;
	    RECT 1384.2001 741.4500 1385.4000 741.6000 ;
	    RECT 1401.0000 741.4500 1402.2001 741.6000 ;
	    RECT 1372.2001 740.5500 1402.2001 741.4500 ;
	    RECT 1372.2001 740.4000 1373.4000 740.5500 ;
	    RECT 1384.2001 740.4000 1385.4000 740.5500 ;
	    RECT 1401.0000 740.4000 1402.2001 740.5500 ;
	    RECT 1410.6000 740.4000 1411.8000 741.6000 ;
	    RECT 1412.7001 740.4000 1414.5000 741.6000 ;
	    RECT 1416.6000 740.7000 1416.9000 742.2000 ;
	    RECT 1417.8000 741.4500 1419.0000 741.6000 ;
	    RECT 1425.0000 741.4500 1426.2001 741.6000 ;
	    RECT 1417.8000 740.5500 1426.2001 741.4500 ;
	    RECT 1417.8000 740.4000 1419.0000 740.5500 ;
	    RECT 1425.0000 740.4000 1426.2001 740.5500 ;
	    RECT 1434.6000 741.4500 1435.8000 741.6000 ;
	    RECT 1453.8000 741.4500 1455.0000 741.6000 ;
	    RECT 1434.6000 740.5500 1455.0000 741.4500 ;
	    RECT 1434.6000 740.4000 1435.8000 740.5500 ;
	    RECT 1453.8000 740.4000 1455.0000 740.5500 ;
	    RECT 1233.0000 738.0000 1234.2001 738.9000 ;
	    RECT 1222.8000 737.1000 1224.0000 738.0000 ;
	    RECT 1233.0000 737.1000 1258.5000 738.0000 ;
	    RECT 1259.4000 737.4000 1260.6000 738.6000 ;
	    RECT 1266.9000 738.0000 1268.1000 738.3000 ;
	    RECT 1261.5000 737.1000 1268.1000 738.0000 ;
	    RECT 1220.7001 735.0000 1222.2001 736.2000 ;
	    RECT 1221.0000 733.5000 1222.2001 735.0000 ;
	    RECT 1223.1000 734.4000 1224.0000 737.1000 ;
	    RECT 1224.9000 736.2000 1226.1000 736.5000 ;
	    RECT 1224.9000 735.3000 1263.3000 736.2000 ;
	    RECT 1259.1000 735.0000 1260.3000 735.3000 ;
	    RECT 1264.2001 734.4000 1265.4000 735.6000 ;
	    RECT 1223.1000 733.5000 1236.6000 734.4000 ;
	    RECT 1201.8000 732.4500 1203.0000 732.6000 ;
	    RECT 1221.0000 732.4500 1222.2001 732.6000 ;
	    RECT 1201.8000 731.5500 1222.2001 732.4500 ;
	    RECT 1201.8000 731.4000 1203.0000 731.5500 ;
	    RECT 1221.0000 731.4000 1222.2001 731.5500 ;
	    RECT 1223.1000 731.1000 1224.0000 733.5000 ;
	    RECT 1235.4000 733.2000 1236.6000 733.5000 ;
	    RECT 1240.2001 733.5000 1253.1000 734.4000 ;
	    RECT 1240.2001 733.2000 1241.4000 733.5000 ;
	    RECT 1227.9000 731.4000 1231.8000 732.6000 ;
	    RECT 1086.6000 723.3000 1087.8000 729.3000 ;
	    RECT 1218.6000 723.3000 1219.8000 729.3000 ;
	    RECT 1221.0000 723.3000 1222.2001 730.5000 ;
	    RECT 1223.1000 730.2000 1227.0000 731.1000 ;
	    RECT 1223.4000 723.3000 1224.6000 729.3000 ;
	    RECT 1225.8000 723.3000 1227.0000 730.2000 ;
	    RECT 1228.2001 723.3000 1229.4000 729.3000 ;
	    RECT 1230.6000 723.3000 1231.8000 731.4000 ;
	    RECT 1232.7001 730.2000 1239.0000 731.4000 ;
	    RECT 1233.0000 723.3000 1234.2001 729.3000 ;
	    RECT 1235.4000 723.3000 1236.6000 727.5000 ;
	    RECT 1237.8000 723.3000 1239.0000 727.5000 ;
	    RECT 1240.2001 723.3000 1241.4000 727.5000 ;
	    RECT 1242.6000 723.3000 1243.8000 732.6000 ;
	    RECT 1247.4000 731.4000 1251.3000 732.6000 ;
	    RECT 1252.2001 732.3000 1253.1000 733.5000 ;
	    RECT 1254.6000 734.1000 1255.8000 734.4000 ;
	    RECT 1254.6000 733.5000 1262.7001 734.1000 ;
	    RECT 1254.6000 733.2000 1263.9000 733.5000 ;
	    RECT 1261.8000 732.3000 1263.9000 733.2000 ;
	    RECT 1252.2001 731.4000 1260.9000 732.3000 ;
	    RECT 1265.4000 732.0000 1267.8000 733.2000 ;
	    RECT 1265.4000 731.4000 1266.3000 732.0000 ;
	    RECT 1245.0000 723.3000 1246.2001 729.3000 ;
	    RECT 1247.4000 723.3000 1248.6000 730.5000 ;
	    RECT 1249.8000 723.3000 1251.0000 729.3000 ;
	    RECT 1252.2001 723.3000 1253.4000 730.5000 ;
	    RECT 1260.0000 730.2000 1266.3000 731.4000 ;
	    RECT 1269.0000 731.1000 1270.2001 739.5000 ;
	    RECT 1276.2001 735.4500 1277.4000 735.6000 ;
	    RECT 1293.0000 735.4500 1294.2001 735.6000 ;
	    RECT 1276.2001 734.5500 1294.2001 735.4500 ;
	    RECT 1276.2001 734.4000 1277.4000 734.5500 ;
	    RECT 1293.0000 734.4000 1294.2001 734.5500 ;
	    RECT 1296.0000 735.3000 1296.9000 740.4000 ;
	    RECT 1297.8000 739.5000 1299.0000 739.8000 ;
	    RECT 1297.8000 738.4500 1299.0000 738.6000 ;
	    RECT 1326.6000 738.4500 1327.8000 738.6000 ;
	    RECT 1297.8000 737.5500 1327.8000 738.4500 ;
	    RECT 1297.8000 737.4000 1299.0000 737.5500 ;
	    RECT 1326.6000 737.4000 1327.8000 737.5500 ;
	    RECT 1317.0000 735.4500 1318.2001 735.6000 ;
	    RECT 1326.6000 735.4500 1327.8000 735.6000 ;
	    RECT 1296.0000 734.4000 1297.5000 735.3000 ;
	    RECT 1294.2001 732.6000 1295.1000 733.5000 ;
	    RECT 1294.2001 731.4000 1295.4000 732.6000 ;
	    RECT 1267.2001 730.2000 1270.2001 731.1000 ;
	    RECT 1254.6000 723.3000 1255.8000 727.5000 ;
	    RECT 1257.0000 723.3000 1258.2001 727.5000 ;
	    RECT 1259.4000 723.3000 1260.6000 729.3000 ;
	    RECT 1261.8000 723.3000 1263.0000 730.2000 ;
	    RECT 1267.2001 729.3000 1268.1000 730.2000 ;
	    RECT 1264.2001 722.4000 1265.4000 729.3000 ;
	    RECT 1266.6000 728.4000 1268.1000 729.3000 ;
	    RECT 1266.6000 723.3000 1267.8000 728.4000 ;
	    RECT 1269.0000 723.3000 1270.2001 729.3000 ;
	    RECT 1293.9000 723.3000 1295.1000 729.3000 ;
	    RECT 1296.3000 723.3000 1297.5000 734.4000 ;
	    RECT 1300.2001 723.3000 1301.4000 735.3000 ;
	    RECT 1317.0000 734.5500 1327.8000 735.4500 ;
	    RECT 1317.0000 734.4000 1318.2001 734.5500 ;
	    RECT 1326.6000 734.4000 1327.8000 734.5500 ;
	    RECT 1329.6000 735.3000 1330.5000 740.4000 ;
	    RECT 1331.4000 739.5000 1332.6000 739.8000 ;
	    RECT 1331.4000 737.4000 1332.6000 738.6000 ;
	    RECT 1350.6000 735.4500 1351.8000 735.6000 ;
	    RECT 1365.0000 735.4500 1366.2001 735.6000 ;
	    RECT 1329.6000 734.4000 1331.1000 735.3000 ;
	    RECT 1327.8000 732.6000 1328.7001 733.5000 ;
	    RECT 1327.8000 731.4000 1329.0000 732.6000 ;
	    RECT 1327.5000 723.3000 1328.7001 729.3000 ;
	    RECT 1329.9000 723.3000 1331.1000 734.4000 ;
	    RECT 1333.8000 723.3000 1335.0000 735.3000 ;
	    RECT 1350.6000 734.5500 1366.2001 735.4500 ;
	    RECT 1350.6000 734.4000 1351.8000 734.5500 ;
	    RECT 1365.0000 734.4000 1366.2001 734.5500 ;
	    RECT 1368.0000 735.3000 1368.9000 740.4000 ;
	    RECT 1369.8000 739.5000 1371.0000 739.8000 ;
	    RECT 1369.8000 737.4000 1371.0000 738.6000 ;
	    RECT 1368.0000 734.4000 1369.5000 735.3000 ;
	    RECT 1366.2001 732.6000 1367.1000 733.5000 ;
	    RECT 1366.2001 731.4000 1367.4000 732.6000 ;
	    RECT 1365.9000 723.3000 1367.1000 729.3000 ;
	    RECT 1368.3000 723.3000 1369.5000 734.4000 ;
	    RECT 1372.2001 723.3000 1373.4000 735.3000 ;
	    RECT 1384.2001 723.3000 1385.4000 739.5000 ;
	    RECT 1405.8000 735.4500 1407.0000 735.6000 ;
	    RECT 1410.6000 735.4500 1411.8000 735.6000 ;
	    RECT 1405.8000 734.5500 1411.8000 735.4500 ;
	    RECT 1405.8000 734.4000 1407.0000 734.5500 ;
	    RECT 1410.6000 734.4000 1411.8000 734.5500 ;
	    RECT 1413.6000 735.3000 1414.5000 740.4000 ;
	    RECT 1415.4000 739.5000 1416.6000 739.8000 ;
	    RECT 1456.2001 739.5000 1457.4000 743.7000 ;
	    RECT 1485.3000 743.1000 1490.7001 743.7000 ;
	    RECT 1492.2001 742.5000 1493.1000 743.7000 ;
	    RECT 1477.8000 741.4500 1479.0000 741.6000 ;
	    RECT 1480.2001 741.4500 1481.4000 741.6000 ;
	    RECT 1485.0000 741.4500 1486.2001 741.6000 ;
	    RECT 1477.8000 740.5500 1486.2001 741.4500 ;
	    RECT 1487.1000 740.7000 1487.4000 742.2000 ;
	    RECT 1477.8000 740.4000 1479.0000 740.5500 ;
	    RECT 1480.2001 740.4000 1481.4000 740.5500 ;
	    RECT 1485.0000 740.4000 1486.2001 740.5500 ;
	    RECT 1489.5000 740.4000 1491.3000 741.6000 ;
	    RECT 1492.2001 741.4500 1493.4000 741.6000 ;
	    RECT 1504.2001 741.4500 1505.4000 741.6000 ;
	    RECT 1492.2001 740.5500 1505.4000 741.4500 ;
	    RECT 1492.2001 740.4000 1493.4000 740.5500 ;
	    RECT 1504.2001 740.4000 1505.4000 740.5500 ;
	    RECT 1506.6000 741.4500 1507.8000 741.6000 ;
	    RECT 1518.6000 741.4500 1519.8000 741.6000 ;
	    RECT 1506.6000 740.5500 1519.8000 741.4500 ;
	    RECT 1506.6000 740.4000 1507.8000 740.5500 ;
	    RECT 1518.6000 740.4000 1519.8000 740.5500 ;
	    RECT 1487.4000 739.5000 1488.6000 739.8000 ;
	    RECT 1415.4000 737.4000 1416.6000 738.6000 ;
	    RECT 1413.6000 734.4000 1415.1000 735.3000 ;
	    RECT 1411.8000 732.6000 1412.7001 733.5000 ;
	    RECT 1411.8000 731.4000 1413.0000 732.6000 ;
	    RECT 1386.6000 723.3000 1387.8000 729.3000 ;
	    RECT 1411.5000 723.3000 1412.7001 729.3000 ;
	    RECT 1413.9000 723.3000 1415.1000 734.4000 ;
	    RECT 1417.8000 723.3000 1419.0000 735.3000 ;
	    RECT 1432.2001 723.3000 1433.4000 729.3000 ;
	    RECT 1434.6000 723.3000 1435.8000 739.5000 ;
	    RECT 1456.2001 738.4500 1457.4000 738.6000 ;
	    RECT 1485.0000 738.4500 1486.2001 738.6000 ;
	    RECT 1456.2001 737.5500 1486.2001 738.4500 ;
	    RECT 1456.2001 737.4000 1457.4000 737.5500 ;
	    RECT 1485.0000 737.4000 1486.2001 737.5500 ;
	    RECT 1487.4000 737.4000 1488.6000 738.6000 ;
	    RECT 1453.8000 723.3000 1455.0000 729.3000 ;
	    RECT 1456.2001 723.3000 1457.4000 736.5000 ;
	    RECT 1458.6000 734.4000 1459.8000 735.6000 ;
	    RECT 1489.5000 735.3000 1490.4000 740.4000 ;
	    RECT 1518.6000 739.2000 1519.8000 739.5000 ;
	    RECT 1506.6000 738.4500 1507.8000 738.6000 ;
	    RECT 1509.0000 738.4500 1510.2001 738.6000 ;
	    RECT 1516.2001 738.4500 1517.4000 738.6000 ;
	    RECT 1506.6000 737.5500 1517.4000 738.4500 ;
	    RECT 1521.0000 738.3000 1521.9000 743.7000 ;
	    RECT 1523.4000 743.4000 1524.6000 744.6000 ;
	    RECT 1549.2001 741.3000 1550.4000 749.7000 ;
	    RECT 1547.7001 740.7000 1550.4000 741.3000 ;
	    RECT 1554.6000 740.7000 1555.8000 749.7000 ;
	    RECT 1547.7001 740.4000 1550.1000 740.7000 ;
	    RECT 1523.4000 738.4500 1524.6000 738.6000 ;
	    RECT 1528.2001 738.4500 1529.4000 738.6000 ;
	    RECT 1506.6000 737.4000 1507.8000 737.5500 ;
	    RECT 1509.0000 737.4000 1510.2001 737.5500 ;
	    RECT 1516.2001 737.4000 1517.4000 737.5500 ;
	    RECT 1518.3000 736.8000 1518.6000 738.3000 ;
	    RECT 1521.0000 737.4000 1522.5000 738.3000 ;
	    RECT 1523.4000 737.5500 1529.4000 738.4500 ;
	    RECT 1523.4000 737.4000 1524.6000 737.5500 ;
	    RECT 1528.2001 737.4000 1529.4000 737.5500 ;
	    RECT 1547.7001 736.5000 1548.6000 740.4000 ;
	    RECT 1551.0000 737.4000 1551.3000 738.6000 ;
	    RECT 1552.2001 737.4000 1553.4000 738.6000 ;
	    RECT 1554.6000 736.5000 1555.8000 736.8000 ;
	    RECT 1458.6000 733.2000 1459.8000 733.5000 ;
	    RECT 1458.6000 723.3000 1459.8000 729.3000 ;
	    RECT 1485.0000 723.3000 1486.2001 735.3000 ;
	    RECT 1488.9000 734.4000 1490.4000 735.3000 ;
	    RECT 1492.2001 734.4000 1493.4000 735.6000 ;
	    RECT 1523.4000 735.3000 1524.3000 736.5000 ;
	    RECT 1516.2001 734.4000 1522.2001 735.3000 ;
	    RECT 1488.9000 723.3000 1490.1000 734.4000 ;
	    RECT 1491.3000 732.6000 1492.2001 733.5000 ;
	    RECT 1491.0000 731.4000 1492.2001 732.6000 ;
	    RECT 1491.3000 723.3000 1492.5000 729.3000 ;
	    RECT 1516.2001 723.3000 1517.4000 734.4000 ;
	    RECT 1518.6000 723.3000 1519.8000 733.5000 ;
	    RECT 1521.0000 723.3000 1522.2001 734.4000 ;
	    RECT 1523.4000 723.3000 1524.6000 735.3000 ;
	    RECT 1547.4000 734.4000 1548.6000 735.6000 ;
	    RECT 1554.6000 734.4000 1555.8000 735.6000 ;
	    RECT 1549.8000 733.5000 1551.0000 733.8000 ;
	    RECT 1547.7001 730.5000 1548.6000 733.5000 ;
	    RECT 1549.8000 731.4000 1551.0000 732.6000 ;
	    RECT 1547.7001 729.6000 1553.1000 730.5000 ;
	    RECT 1547.7001 729.3000 1548.6000 729.6000 ;
	    RECT 1547.4000 723.3000 1548.6000 729.3000 ;
	    RECT 1552.2001 729.3000 1553.1000 729.6000 ;
	    RECT 1549.8000 723.3000 1551.0000 728.7000 ;
	    RECT 1552.2001 723.3000 1553.4000 729.3000 ;
	    RECT 1554.6000 723.3000 1555.8000 729.3000 ;
	    RECT 1566.6000 722.4000 1567.8000 723.6000 ;
	    RECT 1.2000 720.6000 1569.0000 722.4000 ;
	    RECT 49.8000 707.7000 51.0000 719.7000 ;
	    RECT 52.2000 706.8000 53.4000 719.7000 ;
	    RECT 54.6000 707.7000 55.8000 719.7000 ;
	    RECT 57.0000 706.8000 58.2000 719.7000 ;
	    RECT 59.4000 707.7000 60.6000 719.7000 ;
	    RECT 61.8000 706.8000 63.0000 719.7000 ;
	    RECT 64.2000 707.7000 65.4000 719.7000 ;
	    RECT 66.6000 706.8000 67.8000 719.7000 ;
	    RECT 69.0000 707.7000 70.2000 719.7000 ;
	    RECT 81.0000 713.7000 82.2000 719.7000 ;
	    RECT 52.2000 705.6000 54.9000 706.8000 ;
	    RECT 57.0000 705.6000 60.3000 706.8000 ;
	    RECT 61.8000 705.6000 65.1000 706.8000 ;
	    RECT 66.6000 706.5000 70.2000 706.8000 ;
	    RECT 66.6000 705.6000 68.1000 706.5000 ;
	    RECT 53.7000 703.5000 54.9000 705.6000 ;
	    RECT 59.1000 703.5000 60.3000 705.6000 ;
	    RECT 63.9000 703.5000 65.1000 705.6000 ;
	    RECT 69.0000 705.4500 70.2000 705.6000 ;
	    RECT 81.0000 705.4500 82.2000 705.6000 ;
	    RECT 69.0000 704.5500 82.2000 705.4500 ;
	    RECT 69.0000 704.4000 70.2000 704.5500 ;
	    RECT 81.0000 704.4000 82.2000 704.5500 ;
	    RECT 83.4000 703.5000 84.6000 719.7000 ;
	    RECT 97.8000 713.7000 99.0000 719.7000 ;
	    RECT 100.2000 703.5000 101.4000 719.7000 ;
	    RECT 124.2000 707.7000 125.4000 719.7000 ;
	    RECT 128.1000 708.6000 129.3000 719.7000 ;
	    RECT 130.5000 713.7000 131.7000 719.7000 ;
	    RECT 130.2000 710.4000 131.4000 711.6000 ;
	    RECT 130.5000 709.5000 131.4000 710.4000 ;
	    RECT 128.1000 707.7000 129.6000 708.6000 ;
	    RECT 126.6000 705.4500 127.8000 705.6000 ;
	    RECT 121.9500 704.5500 127.8000 705.4500 ;
	    RECT 49.8000 701.4000 51.0000 702.6000 ;
	    RECT 51.9000 702.3000 52.5000 703.5000 ;
	    RECT 53.7000 702.3000 57.6000 703.5000 ;
	    RECT 59.1000 702.3000 62.7000 703.5000 ;
	    RECT 63.9000 702.3000 67.8000 703.5000 ;
	    RECT 53.7000 701.4000 54.9000 702.3000 ;
	    RECT 59.1000 701.4000 60.3000 702.3000 ;
	    RECT 63.9000 701.4000 65.1000 702.3000 ;
	    RECT 69.0000 701.4000 70.2000 703.5000 ;
	    RECT 83.4000 702.4500 84.6000 702.6000 ;
	    RECT 95.4000 702.4500 96.6000 702.6000 ;
	    RECT 83.4000 701.5500 96.6000 702.4500 ;
	    RECT 83.4000 701.4000 84.6000 701.5500 ;
	    RECT 95.4000 701.4000 96.6000 701.5500 ;
	    RECT 100.2000 702.4500 101.4000 702.6000 ;
	    RECT 121.9500 702.4500 122.8500 704.5500 ;
	    RECT 126.6000 704.4000 127.8000 704.5500 ;
	    RECT 126.6000 703.2000 127.8000 703.5000 ;
	    RECT 128.7000 702.6000 129.6000 707.7000 ;
	    RECT 131.4000 708.4500 132.6000 708.6000 ;
	    RECT 141.0000 708.4500 142.2000 708.6000 ;
	    RECT 131.4000 707.5500 142.2000 708.4500 ;
	    RECT 162.6000 707.7000 163.8000 719.7000 ;
	    RECT 166.5000 707.7000 169.5000 719.7000 ;
	    RECT 172.2000 707.7000 173.4000 719.7000 ;
	    RECT 192.3000 708.9000 193.5000 719.7000 ;
	    RECT 192.3000 707.7000 195.0000 708.9000 ;
	    RECT 196.2000 707.7000 197.4000 719.7000 ;
	    RECT 222.6000 707.7000 223.8000 719.7000 ;
	    RECT 226.5000 708.9000 227.7000 719.7000 ;
	    RECT 246.6000 713.7000 247.8000 719.7000 ;
	    RECT 225.0000 707.7000 227.7000 708.9000 ;
	    RECT 131.4000 707.4000 132.6000 707.5500 ;
	    RECT 141.0000 707.4000 142.2000 707.5500 ;
	    RECT 136.2000 705.4500 137.4000 705.6000 ;
	    RECT 136.2000 704.5500 161.2500 705.4500 ;
	    RECT 136.2000 704.4000 137.4000 704.5500 ;
	    RECT 100.2000 701.5500 122.8500 702.4500 ;
	    RECT 100.2000 701.4000 101.4000 701.5500 ;
	    RECT 124.2000 701.4000 125.4000 702.6000 ;
	    RECT 52.2000 700.2000 54.9000 701.4000 ;
	    RECT 57.0000 700.2000 60.3000 701.4000 ;
	    RECT 61.8000 700.2000 65.1000 701.4000 ;
	    RECT 66.6000 700.2000 70.2000 701.4000 ;
	    RECT 126.3000 700.8000 126.6000 702.3000 ;
	    RECT 128.7000 701.4000 130.5000 702.6000 ;
	    RECT 131.4000 702.4500 132.6000 702.6000 ;
	    RECT 155.4000 702.4500 156.6000 702.6000 ;
	    RECT 131.4000 701.5500 156.6000 702.4500 ;
	    RECT 160.3500 702.4500 161.2500 704.5500 ;
	    RECT 165.0000 704.4000 166.2000 705.6000 ;
	    RECT 162.6000 703.5000 163.8000 703.8000 ;
	    RECT 167.7000 703.5000 168.6000 707.7000 ;
	    RECT 191.4000 706.5000 192.6000 706.8000 ;
	    RECT 169.8000 704.4000 171.0000 705.6000 ;
	    RECT 172.2000 705.4500 173.4000 705.6000 ;
	    RECT 191.4000 705.4500 192.6000 705.6000 ;
	    RECT 172.2000 704.5500 192.6000 705.4500 ;
	    RECT 172.2000 704.4000 173.4000 704.5500 ;
	    RECT 191.4000 704.4000 192.6000 704.5500 ;
	    RECT 193.8000 703.5000 194.7000 707.7000 ;
	    RECT 225.3000 703.5000 226.2000 707.7000 ;
	    RECT 227.4000 706.5000 228.6000 706.8000 ;
	    RECT 249.0000 706.5000 250.2000 719.7000 ;
	    RECT 251.4000 713.7000 252.6000 719.7000 ;
	    RECT 268.2000 719.4000 269.4000 720.6000 ;
	    RECT 270.6000 713.7000 271.8000 719.7000 ;
	    RECT 251.4000 709.5000 252.6000 709.8000 ;
	    RECT 251.4000 707.4000 252.6000 708.6000 ;
	    RECT 265.8000 708.4500 267.0000 708.6000 ;
	    RECT 253.9500 707.5500 267.0000 708.4500 ;
	    RECT 227.4000 705.4500 228.6000 705.6000 ;
	    RECT 232.2000 705.4500 233.4000 705.6000 ;
	    RECT 227.4000 704.5500 233.4000 705.4500 ;
	    RECT 227.4000 704.4000 228.6000 704.5500 ;
	    RECT 232.2000 704.4000 233.4000 704.5500 ;
	    RECT 249.0000 705.4500 250.2000 705.6000 ;
	    RECT 253.9500 705.4500 254.8500 707.5500 ;
	    RECT 265.8000 707.4000 267.0000 707.5500 ;
	    RECT 273.0000 706.5000 274.2000 719.7000 ;
	    RECT 275.4000 713.7000 276.6000 719.7000 ;
	    RECT 275.4000 709.5000 276.6000 709.8000 ;
	    RECT 275.4000 708.4500 276.6000 708.6000 ;
	    RECT 301.8000 708.4500 303.0000 708.6000 ;
	    RECT 275.4000 707.5500 303.0000 708.4500 ;
	    RECT 306.6000 707.7000 307.8000 719.7000 ;
	    RECT 310.5000 707.7000 313.5000 719.7000 ;
	    RECT 316.2000 707.7000 317.4000 719.7000 ;
	    RECT 335.4000 707.7000 336.6000 719.7000 ;
	    RECT 339.3000 708.9000 340.5000 719.7000 ;
	    RECT 359.4000 713.7000 360.6000 719.7000 ;
	    RECT 337.8000 707.7000 340.5000 708.9000 ;
	    RECT 354.6000 708.4500 355.8000 708.6000 ;
	    RECT 275.4000 707.4000 276.6000 707.5500 ;
	    RECT 301.8000 707.4000 303.0000 707.5500 ;
	    RECT 249.0000 704.5500 254.8500 705.4500 ;
	    RECT 256.2000 705.4500 257.4000 705.6000 ;
	    RECT 273.0000 705.4500 274.2000 705.6000 ;
	    RECT 256.2000 704.5500 274.2000 705.4500 ;
	    RECT 249.0000 704.4000 250.2000 704.5500 ;
	    RECT 256.2000 704.4000 257.4000 704.5500 ;
	    RECT 273.0000 704.4000 274.2000 704.5500 ;
	    RECT 309.0000 704.4000 310.2000 705.6000 ;
	    RECT 306.6000 703.5000 307.8000 703.8000 ;
	    RECT 311.7000 703.5000 312.6000 707.7000 ;
	    RECT 313.8000 704.4000 315.0000 705.6000 ;
	    RECT 338.1000 703.5000 339.0000 707.7000 ;
	    RECT 342.7500 707.5500 355.8000 708.4500 ;
	    RECT 340.2000 706.5000 341.4000 706.8000 ;
	    RECT 340.2000 705.4500 341.4000 705.6000 ;
	    RECT 342.7500 705.4500 343.6500 707.5500 ;
	    RECT 354.6000 707.4000 355.8000 707.5500 ;
	    RECT 361.8000 706.5000 363.0000 719.7000 ;
	    RECT 364.2000 713.7000 365.4000 719.7000 ;
	    RECT 383.4000 713.7000 384.6000 719.7000 ;
	    RECT 364.2000 709.5000 365.4000 709.8000 ;
	    RECT 383.4000 709.5000 384.6000 709.8000 ;
	    RECT 364.2000 708.4500 365.4000 708.6000 ;
	    RECT 366.6000 708.4500 367.8000 708.6000 ;
	    RECT 364.2000 707.5500 367.8000 708.4500 ;
	    RECT 364.2000 707.4000 365.4000 707.5500 ;
	    RECT 366.6000 707.4000 367.8000 707.5500 ;
	    RECT 369.0000 708.4500 370.2000 708.6000 ;
	    RECT 383.4000 708.4500 384.6000 708.6000 ;
	    RECT 369.0000 707.5500 384.6000 708.4500 ;
	    RECT 369.0000 707.4000 370.2000 707.5500 ;
	    RECT 383.4000 707.4000 384.6000 707.5500 ;
	    RECT 385.8000 706.5000 387.0000 719.7000 ;
	    RECT 388.2000 713.7000 389.4000 719.7000 ;
	    RECT 412.2000 707.7000 413.4000 719.7000 ;
	    RECT 416.1000 708.6000 417.3000 719.7000 ;
	    RECT 418.5000 713.7000 419.7000 719.7000 ;
	    RECT 418.2000 710.4000 419.4000 711.6000 ;
	    RECT 418.5000 709.5000 419.4000 710.4000 ;
	    RECT 416.1000 707.7000 417.6000 708.6000 ;
	    RECT 340.2000 704.5500 343.6500 705.4500 ;
	    RECT 352.2000 705.4500 353.4000 705.6000 ;
	    RECT 361.8000 705.4500 363.0000 705.6000 ;
	    RECT 352.2000 704.5500 363.0000 705.4500 ;
	    RECT 340.2000 704.4000 341.4000 704.5500 ;
	    RECT 352.2000 704.4000 353.4000 704.5500 ;
	    RECT 361.8000 704.4000 363.0000 704.5500 ;
	    RECT 385.8000 705.4500 387.0000 705.6000 ;
	    RECT 412.2000 705.4500 413.4000 705.6000 ;
	    RECT 385.8000 704.5500 413.4000 705.4500 ;
	    RECT 385.8000 704.4000 387.0000 704.5500 ;
	    RECT 412.2000 704.4000 413.4000 704.5500 ;
	    RECT 414.6000 704.4000 415.8000 705.6000 ;
	    RECT 165.0000 703.2000 166.2000 703.5000 ;
	    RECT 169.8000 703.2000 171.0000 703.5000 ;
	    RECT 162.6000 702.4500 163.8000 702.6000 ;
	    RECT 160.3500 701.5500 163.8000 702.4500 ;
	    RECT 131.4000 701.4000 132.6000 701.5500 ;
	    RECT 155.4000 701.4000 156.6000 701.5500 ;
	    RECT 162.6000 701.4000 163.8000 701.5500 ;
	    RECT 165.0000 701.4000 166.5000 702.3000 ;
	    RECT 167.4000 701.4000 168.6000 702.6000 ;
	    RECT 49.8000 693.3000 51.0000 699.3000 ;
	    RECT 52.2000 693.3000 53.4000 700.2000 ;
	    RECT 54.6000 693.3000 55.8000 699.3000 ;
	    RECT 57.0000 693.3000 58.2000 700.2000 ;
	    RECT 59.4000 693.3000 60.6000 699.3000 ;
	    RECT 61.8000 693.3000 63.0000 700.2000 ;
	    RECT 64.2000 693.3000 65.4000 699.3000 ;
	    RECT 66.6000 693.3000 67.8000 700.2000 ;
	    RECT 71.4000 699.4500 72.6000 699.6000 ;
	    RECT 81.0000 699.4500 82.2000 699.6000 ;
	    RECT 69.0000 693.3000 70.2000 699.3000 ;
	    RECT 71.4000 698.5500 82.2000 699.4500 ;
	    RECT 71.4000 698.4000 72.6000 698.5500 ;
	    RECT 81.0000 698.4000 82.2000 698.5500 ;
	    RECT 81.0000 697.2000 82.2000 697.5000 ;
	    RECT 81.0000 693.3000 82.2000 696.3000 ;
	    RECT 83.4000 693.3000 84.6000 700.5000 ;
	    RECT 97.8000 698.4000 99.0000 699.6000 ;
	    RECT 97.8000 697.2000 99.0000 697.5000 ;
	    RECT 97.8000 693.3000 99.0000 696.3000 ;
	    RECT 100.2000 693.3000 101.4000 700.5000 ;
	    RECT 124.5000 699.3000 129.9000 699.9000 ;
	    RECT 131.4000 699.3000 132.3000 700.5000 ;
	    RECT 165.0000 699.3000 165.9000 701.4000 ;
	    RECT 171.0000 700.8000 171.3000 702.3000 ;
	    RECT 172.2000 701.4000 173.4000 702.6000 ;
	    RECT 189.0000 702.4500 190.2000 702.6000 ;
	    RECT 193.8000 702.4500 195.0000 702.6000 ;
	    RECT 189.0000 701.5500 195.0000 702.4500 ;
	    RECT 189.0000 701.4000 190.2000 701.5500 ;
	    RECT 193.8000 701.4000 195.0000 701.5500 ;
	    RECT 196.2000 702.4500 197.4000 702.6000 ;
	    RECT 225.0000 702.4500 226.2000 702.6000 ;
	    RECT 239.4000 702.4500 240.6000 702.6000 ;
	    RECT 196.2000 701.5500 223.6500 702.4500 ;
	    RECT 196.2000 701.4000 197.4000 701.5500 ;
	    RECT 167.7000 699.3000 173.1000 699.9000 ;
	    RECT 124.2000 699.0000 130.2000 699.3000 ;
	    RECT 124.2000 693.3000 125.4000 699.0000 ;
	    RECT 126.6000 693.3000 127.8000 698.1000 ;
	    RECT 129.0000 693.3000 130.2000 699.0000 ;
	    RECT 131.4000 693.3000 132.6000 699.3000 ;
	    RECT 162.6000 694.2000 163.8000 699.3000 ;
	    RECT 165.0000 695.1000 166.2000 699.3000 ;
	    RECT 167.4000 699.0000 173.4000 699.3000 ;
	    RECT 167.4000 694.2000 168.6000 699.0000 ;
	    RECT 162.6000 693.3000 168.6000 694.2000 ;
	    RECT 169.8000 693.3000 171.0000 698.1000 ;
	    RECT 172.2000 693.3000 173.4000 699.0000 ;
	    RECT 193.8000 696.3000 194.7000 700.5000 ;
	    RECT 222.7500 699.6000 223.6500 701.5500 ;
	    RECT 225.0000 701.5500 240.6000 702.4500 ;
	    RECT 225.0000 701.4000 226.2000 701.5500 ;
	    RECT 239.4000 701.4000 240.6000 701.5500 ;
	    RECT 246.6000 701.4000 247.8000 702.6000 ;
	    RECT 196.2000 698.4000 197.4000 699.6000 ;
	    RECT 222.6000 698.4000 223.8000 699.6000 ;
	    RECT 196.2000 697.2000 197.4000 697.5000 ;
	    RECT 222.6000 697.2000 223.8000 697.5000 ;
	    RECT 198.6000 696.4500 199.8000 696.6000 ;
	    RECT 220.2000 696.4500 221.4000 696.6000 ;
	    RECT 191.4000 693.3000 192.6000 696.3000 ;
	    RECT 193.8000 693.3000 195.0000 696.3000 ;
	    RECT 196.2000 693.3000 197.4000 696.3000 ;
	    RECT 198.6000 695.5500 221.4000 696.4500 ;
	    RECT 225.3000 696.3000 226.2000 700.5000 ;
	    RECT 246.6000 700.2000 247.8000 700.5000 ;
	    RECT 249.0000 699.3000 250.2000 703.5000 ;
	    RECT 270.6000 701.4000 271.8000 702.6000 ;
	    RECT 270.6000 700.2000 271.8000 700.5000 ;
	    RECT 273.0000 699.3000 274.2000 703.5000 ;
	    RECT 309.0000 703.2000 310.2000 703.5000 ;
	    RECT 313.8000 703.2000 315.0000 703.5000 ;
	    RECT 285.0000 702.4500 286.2000 702.6000 ;
	    RECT 306.6000 702.4500 307.8000 702.6000 ;
	    RECT 285.0000 701.5500 307.8000 702.4500 ;
	    RECT 285.0000 701.4000 286.2000 701.5500 ;
	    RECT 306.6000 701.4000 307.8000 701.5500 ;
	    RECT 309.0000 701.4000 310.5000 702.3000 ;
	    RECT 311.4000 701.4000 312.6000 702.6000 ;
	    RECT 309.0000 699.3000 309.9000 701.4000 ;
	    RECT 315.0000 700.8000 315.3000 702.3000 ;
	    RECT 316.2000 701.4000 317.4000 702.6000 ;
	    RECT 325.8000 702.4500 327.0000 702.6000 ;
	    RECT 337.8000 702.4500 339.0000 702.6000 ;
	    RECT 325.8000 701.5500 339.0000 702.4500 ;
	    RECT 325.8000 701.4000 327.0000 701.5500 ;
	    RECT 337.8000 701.4000 339.0000 701.5500 ;
	    RECT 340.2000 702.4500 341.4000 702.6000 ;
	    RECT 349.8000 702.4500 351.0000 702.6000 ;
	    RECT 354.6000 702.4500 355.8000 702.6000 ;
	    RECT 359.4000 702.4500 360.6000 702.6000 ;
	    RECT 340.2000 701.5500 360.6000 702.4500 ;
	    RECT 340.2000 701.4000 341.4000 701.5500 ;
	    RECT 349.8000 701.4000 351.0000 701.5500 ;
	    RECT 354.6000 701.4000 355.8000 701.5500 ;
	    RECT 359.4000 701.4000 360.6000 701.5500 ;
	    RECT 311.7000 699.3000 317.1000 699.9000 ;
	    RECT 318.6000 699.4500 319.8000 699.6000 ;
	    RECT 335.4000 699.4500 336.6000 699.6000 ;
	    RECT 198.6000 695.4000 199.8000 695.5500 ;
	    RECT 220.2000 695.4000 221.4000 695.5500 ;
	    RECT 222.6000 693.3000 223.8000 696.3000 ;
	    RECT 225.0000 693.3000 226.2000 696.3000 ;
	    RECT 227.4000 693.3000 228.6000 696.3000 ;
	    RECT 246.6000 693.3000 247.8000 699.3000 ;
	    RECT 249.0000 698.4000 251.7000 699.3000 ;
	    RECT 250.5000 693.3000 251.7000 698.4000 ;
	    RECT 270.6000 693.3000 271.8000 699.3000 ;
	    RECT 273.0000 698.4000 275.7000 699.3000 ;
	    RECT 274.5000 693.3000 275.7000 698.4000 ;
	    RECT 306.6000 694.2000 307.8000 699.3000 ;
	    RECT 309.0000 695.1000 310.2000 699.3000 ;
	    RECT 311.4000 699.0000 317.4000 699.3000 ;
	    RECT 311.4000 694.2000 312.6000 699.0000 ;
	    RECT 306.6000 693.3000 312.6000 694.2000 ;
	    RECT 313.8000 693.3000 315.0000 698.1000 ;
	    RECT 316.2000 693.3000 317.4000 699.0000 ;
	    RECT 318.6000 698.5500 336.6000 699.4500 ;
	    RECT 318.6000 698.4000 319.8000 698.5500 ;
	    RECT 335.4000 698.4000 336.6000 698.5500 ;
	    RECT 335.4000 697.2000 336.6000 697.5000 ;
	    RECT 338.1000 696.3000 339.0000 700.5000 ;
	    RECT 359.4000 700.2000 360.6000 700.5000 ;
	    RECT 361.8000 699.3000 363.0000 703.5000 ;
	    RECT 385.8000 699.3000 387.0000 703.5000 ;
	    RECT 414.6000 703.2000 415.8000 703.5000 ;
	    RECT 416.7000 702.6000 417.6000 707.7000 ;
	    RECT 419.4000 707.4000 420.6000 708.6000 ;
	    RECT 441.0000 703.5000 442.2000 719.7000 ;
	    RECT 443.4000 713.7000 444.6000 719.7000 ;
	    RECT 462.6000 708.6000 463.8000 719.7000 ;
	    RECT 465.0000 709.5000 466.2000 719.7000 ;
	    RECT 462.6000 707.7000 465.9000 708.6000 ;
	    RECT 467.4000 707.7000 468.6000 719.7000 ;
	    RECT 594.6000 713.7000 595.8000 719.7000 ;
	    RECT 597.0000 714.6000 598.2000 719.7000 ;
	    RECT 596.7000 713.7000 598.2000 714.6000 ;
	    RECT 599.4000 713.7000 600.6000 720.6000 ;
	    RECT 596.7000 712.8000 597.6000 713.7000 ;
	    RECT 601.8000 712.8000 603.0000 719.7000 ;
	    RECT 604.2000 713.7000 605.4000 719.7000 ;
	    RECT 606.6000 715.5000 607.8000 719.7000 ;
	    RECT 609.0000 715.5000 610.2000 719.7000 ;
	    RECT 465.0000 706.8000 465.9000 707.7000 ;
	    RECT 465.0000 705.6000 466.8000 706.8000 ;
	    RECT 462.6000 703.2000 463.8000 703.5000 ;
	    RECT 388.2000 702.4500 389.4000 702.6000 ;
	    RECT 405.0000 702.4500 406.2000 702.6000 ;
	    RECT 388.2000 701.5500 406.2000 702.4500 ;
	    RECT 388.2000 701.4000 389.4000 701.5500 ;
	    RECT 405.0000 701.4000 406.2000 701.5500 ;
	    RECT 412.2000 701.4000 413.4000 702.6000 ;
	    RECT 414.3000 700.8000 414.6000 702.3000 ;
	    RECT 416.7000 701.4000 418.5000 702.6000 ;
	    RECT 419.4000 701.4000 420.6000 702.6000 ;
	    RECT 421.8000 702.4500 423.0000 702.6000 ;
	    RECT 441.0000 702.4500 442.2000 702.6000 ;
	    RECT 421.8000 701.5500 442.2000 702.4500 ;
	    RECT 421.8000 701.4000 423.0000 701.5500 ;
	    RECT 441.0000 701.4000 442.2000 701.5500 ;
	    RECT 465.0000 701.1000 465.9000 705.6000 ;
	    RECT 467.7000 704.4000 468.6000 707.7000 ;
	    RECT 467.4000 703.5000 468.6000 704.4000 ;
	    RECT 594.6000 711.9000 597.6000 712.8000 ;
	    RECT 594.6000 703.5000 595.8000 711.9000 ;
	    RECT 598.5000 711.6000 604.8000 712.8000 ;
	    RECT 611.4000 712.5000 612.6000 719.7000 ;
	    RECT 613.8000 713.7000 615.0000 719.7000 ;
	    RECT 616.2000 712.5000 617.4000 719.7000 ;
	    RECT 618.6000 713.7000 619.8000 719.7000 ;
	    RECT 598.5000 711.0000 599.4000 711.6000 ;
	    RECT 597.0000 709.8000 599.4000 711.0000 ;
	    RECT 603.9000 710.7000 612.6000 711.6000 ;
	    RECT 600.9000 709.8000 603.0000 710.7000 ;
	    RECT 600.9000 709.5000 610.2000 709.8000 ;
	    RECT 602.1000 708.9000 610.2000 709.5000 ;
	    RECT 609.0000 708.6000 610.2000 708.9000 ;
	    RECT 611.7000 709.5000 612.6000 710.7000 ;
	    RECT 613.5000 710.4000 617.4000 711.6000 ;
	    RECT 621.0000 710.4000 622.2000 719.7000 ;
	    RECT 623.4000 715.5000 624.6000 719.7000 ;
	    RECT 625.8000 715.5000 627.0000 719.7000 ;
	    RECT 628.2000 715.5000 629.4000 719.7000 ;
	    RECT 630.6000 713.7000 631.8000 719.7000 ;
	    RECT 625.8000 711.6000 632.1000 712.8000 ;
	    RECT 633.0000 711.6000 634.2000 719.7000 ;
	    RECT 635.4000 713.7000 636.6000 719.7000 ;
	    RECT 637.8000 712.8000 639.0000 719.7000 ;
	    RECT 640.2000 713.7000 641.4000 719.7000 ;
	    RECT 637.8000 711.9000 641.7000 712.8000 ;
	    RECT 642.6000 712.5000 643.8000 719.7000 ;
	    RECT 645.0000 713.7000 646.2000 719.7000 ;
	    RECT 671.4000 713.7000 672.6000 719.7000 ;
	    RECT 633.0000 710.4000 636.9000 711.6000 ;
	    RECT 623.4000 709.5000 624.6000 709.8000 ;
	    RECT 611.7000 708.6000 624.6000 709.5000 ;
	    RECT 628.2000 709.5000 629.4000 709.8000 ;
	    RECT 640.8000 709.5000 641.7000 711.9000 ;
	    RECT 642.6000 710.4000 643.8000 711.6000 ;
	    RECT 628.2000 708.6000 641.7000 709.5000 ;
	    RECT 599.4000 707.4000 600.6000 708.6000 ;
	    RECT 604.5000 707.7000 605.7000 708.0000 ;
	    RECT 601.5000 706.8000 639.9000 707.7000 ;
	    RECT 638.7000 706.5000 639.9000 706.8000 ;
	    RECT 640.8000 705.9000 641.7000 708.6000 ;
	    RECT 642.6000 708.0000 643.8000 709.5000 ;
	    RECT 642.6000 706.8000 644.1000 708.0000 ;
	    RECT 596.7000 705.0000 603.3000 705.9000 ;
	    RECT 596.7000 704.7000 597.9000 705.0000 ;
	    RECT 604.2000 704.4000 605.4000 705.6000 ;
	    RECT 606.3000 705.0000 631.8000 705.9000 ;
	    RECT 640.8000 705.0000 642.0000 705.9000 ;
	    RECT 630.6000 704.1000 631.8000 705.0000 ;
	    RECT 467.4000 702.4500 468.6000 702.6000 ;
	    RECT 479.4000 702.4500 480.6000 702.6000 ;
	    RECT 467.4000 701.5500 480.6000 702.4500 ;
	    RECT 467.4000 701.4000 468.6000 701.5500 ;
	    RECT 479.4000 701.4000 480.6000 701.5500 ;
	    RECT 594.6000 702.3000 607.8000 703.5000 ;
	    RECT 608.7000 702.9000 611.7000 704.1000 ;
	    RECT 617.4000 702.9000 622.2000 704.1000 ;
	    RECT 388.2000 700.2000 389.4000 700.5000 ;
	    RECT 412.5000 699.3000 417.9000 699.9000 ;
	    RECT 419.4000 699.3000 420.3000 700.5000 ;
	    RECT 335.4000 693.3000 336.6000 696.3000 ;
	    RECT 337.8000 693.3000 339.0000 696.3000 ;
	    RECT 340.2000 693.3000 341.4000 696.3000 ;
	    RECT 359.4000 693.3000 360.6000 699.3000 ;
	    RECT 361.8000 698.4000 364.5000 699.3000 ;
	    RECT 363.3000 693.3000 364.5000 698.4000 ;
	    RECT 384.3000 698.4000 387.0000 699.3000 ;
	    RECT 384.3000 693.3000 385.5000 698.4000 ;
	    RECT 388.2000 693.3000 389.4000 699.3000 ;
	    RECT 412.2000 699.0000 418.2000 699.3000 ;
	    RECT 412.2000 693.3000 413.4000 699.0000 ;
	    RECT 414.6000 693.3000 415.8000 698.1000 ;
	    RECT 417.0000 693.3000 418.2000 699.0000 ;
	    RECT 419.4000 693.3000 420.6000 699.3000 ;
	    RECT 441.0000 693.3000 442.2000 700.5000 ;
	    RECT 462.6000 700.2000 465.9000 701.1000 ;
	    RECT 443.4000 699.4500 444.6000 699.6000 ;
	    RECT 460.2000 699.4500 461.4000 699.6000 ;
	    RECT 443.4000 698.5500 461.4000 699.4500 ;
	    RECT 443.4000 698.4000 444.6000 698.5500 ;
	    RECT 460.2000 698.4000 461.4000 698.5500 ;
	    RECT 443.4000 697.2000 444.6000 697.5000 ;
	    RECT 443.4000 693.3000 444.6000 696.3000 ;
	    RECT 462.6000 693.3000 463.8000 700.2000 ;
	    RECT 465.0000 693.3000 466.2000 699.3000 ;
	    RECT 467.4000 693.3000 468.6000 700.5000 ;
	    RECT 594.6000 693.3000 595.8000 702.3000 ;
	    RECT 598.2000 700.2000 602.7000 701.4000 ;
	    RECT 601.5000 699.3000 602.7000 700.2000 ;
	    RECT 610.5000 699.3000 611.7000 702.9000 ;
	    RECT 613.8000 701.4000 615.0000 702.6000 ;
	    RECT 621.6000 701.7000 622.8000 702.0000 ;
	    RECT 616.2000 700.8000 622.8000 701.7000 ;
	    RECT 616.2000 700.5000 617.4000 700.8000 ;
	    RECT 613.8000 700.2000 615.0000 700.5000 ;
	    RECT 625.8000 699.6000 627.0000 703.8000 ;
	    RECT 634.5000 702.9000 640.2000 704.1000 ;
	    RECT 634.5000 701.1000 635.7000 702.9000 ;
	    RECT 641.1000 702.0000 642.0000 705.0000 ;
	    RECT 616.2000 699.3000 617.4000 699.6000 ;
	    RECT 599.4000 693.3000 600.6000 699.3000 ;
	    RECT 601.5000 698.1000 605.4000 699.3000 ;
	    RECT 610.5000 698.4000 617.4000 699.3000 ;
	    RECT 618.6000 698.4000 619.8000 699.6000 ;
	    RECT 620.7000 698.4000 621.0000 699.6000 ;
	    RECT 625.5000 698.4000 627.0000 699.6000 ;
	    RECT 633.0000 700.2000 635.7000 701.1000 ;
	    RECT 640.2000 701.1000 642.0000 702.0000 ;
	    RECT 633.0000 699.3000 634.2000 700.2000 ;
	    RECT 604.2000 693.3000 605.4000 698.1000 ;
	    RECT 630.6000 698.1000 634.2000 699.3000 ;
	    RECT 606.6000 693.3000 607.8000 697.5000 ;
	    RECT 609.0000 693.3000 610.2000 697.5000 ;
	    RECT 611.4000 693.3000 612.6000 697.5000 ;
	    RECT 613.8000 693.3000 615.0000 696.3000 ;
	    RECT 616.2000 693.3000 617.4000 697.5000 ;
	    RECT 618.6000 693.3000 619.8000 696.3000 ;
	    RECT 621.0000 693.3000 622.2000 697.5000 ;
	    RECT 623.4000 693.3000 624.6000 697.5000 ;
	    RECT 625.8000 693.3000 627.0000 697.5000 ;
	    RECT 628.2000 693.3000 629.4000 697.5000 ;
	    RECT 630.6000 693.3000 631.8000 698.1000 ;
	    RECT 635.4000 693.3000 636.6000 699.3000 ;
	    RECT 640.2000 693.3000 641.4000 701.1000 ;
	    RECT 642.9000 700.2000 644.1000 706.8000 ;
	    RECT 673.8000 706.5000 675.0000 719.7000 ;
	    RECT 676.2000 713.7000 677.4000 719.7000 ;
	    RECT 676.2000 709.5000 677.4000 709.8000 ;
	    RECT 696.3000 708.9000 697.5000 719.7000 ;
	    RECT 676.2000 707.4000 677.4000 708.6000 ;
	    RECT 696.3000 707.7000 699.0000 708.9000 ;
	    RECT 700.2000 707.7000 701.4000 719.7000 ;
	    RECT 714.6000 713.7000 715.8000 719.7000 ;
	    RECT 695.4000 706.5000 696.6000 706.8000 ;
	    RECT 654.6000 705.4500 655.8000 705.6000 ;
	    RECT 673.8000 705.4500 675.0000 705.6000 ;
	    RECT 654.6000 704.5500 675.0000 705.4500 ;
	    RECT 654.6000 704.4000 655.8000 704.5500 ;
	    RECT 673.8000 704.4000 675.0000 704.5500 ;
	    RECT 695.4000 704.4000 696.6000 705.6000 ;
	    RECT 697.8000 703.5000 698.7000 707.7000 ;
	    RECT 717.0000 703.5000 718.2000 719.7000 ;
	    RECT 741.0000 713.7000 742.2000 719.7000 ;
	    RECT 743.4000 713.7000 744.6000 719.7000 ;
	    RECT 745.8000 714.3000 747.0000 719.7000 ;
	    RECT 743.7000 713.4000 744.6000 713.7000 ;
	    RECT 748.2000 713.7000 749.4000 719.7000 ;
	    RECT 772.2000 713.7000 773.4000 719.7000 ;
	    RECT 774.6000 713.7000 775.8000 719.7000 ;
	    RECT 777.0000 714.3000 778.2000 719.7000 ;
	    RECT 748.2000 713.4000 749.1000 713.7000 ;
	    RECT 743.7000 712.5000 749.1000 713.4000 ;
	    RECT 774.9000 713.4000 775.8000 713.7000 ;
	    RECT 779.4000 713.7000 780.6000 719.7000 ;
	    RECT 798.6000 713.7000 799.8000 719.7000 ;
	    RECT 779.4000 713.4000 780.3000 713.7000 ;
	    RECT 774.9000 712.5000 780.3000 713.4000 ;
	    RECT 733.8000 711.4500 735.0000 711.6000 ;
	    RECT 743.4000 711.4500 744.6000 711.6000 ;
	    RECT 733.8000 710.5500 744.6000 711.4500 ;
	    RECT 733.8000 710.4000 735.0000 710.5500 ;
	    RECT 743.4000 710.4000 744.6000 710.5500 ;
	    RECT 745.8000 710.4000 747.0000 711.6000 ;
	    RECT 748.2000 709.5000 749.1000 712.5000 ;
	    RECT 750.6000 711.4500 751.8000 711.6000 ;
	    RECT 777.0000 711.4500 778.2000 711.6000 ;
	    RECT 750.6000 710.5500 778.2000 711.4500 ;
	    RECT 750.6000 710.4000 751.8000 710.5500 ;
	    RECT 777.0000 710.4000 778.2000 710.5500 ;
	    RECT 779.4000 709.5000 780.3000 712.5000 ;
	    RECT 781.8000 711.4500 783.0000 711.6000 ;
	    RECT 798.6000 711.4500 799.8000 711.6000 ;
	    RECT 781.8000 710.5500 799.8000 711.4500 ;
	    RECT 781.8000 710.4000 783.0000 710.5500 ;
	    RECT 798.6000 710.4000 799.8000 710.5500 ;
	    RECT 745.8000 709.2000 747.0000 709.5000 ;
	    RECT 777.0000 709.2000 778.2000 709.5000 ;
	    RECT 721.8000 708.4500 723.0000 708.6000 ;
	    RECT 741.0000 708.4500 742.2000 708.6000 ;
	    RECT 721.8000 707.5500 742.2000 708.4500 ;
	    RECT 721.8000 707.4000 723.0000 707.5500 ;
	    RECT 741.0000 707.4000 742.2000 707.5500 ;
	    RECT 748.2000 708.4500 749.4000 708.6000 ;
	    RECT 765.0000 708.4500 766.2000 708.6000 ;
	    RECT 748.2000 707.5500 766.2000 708.4500 ;
	    RECT 748.2000 707.4000 749.4000 707.5500 ;
	    RECT 765.0000 707.4000 766.2000 707.5500 ;
	    RECT 772.2000 707.4000 773.4000 708.6000 ;
	    RECT 779.4000 708.4500 780.6000 708.6000 ;
	    RECT 784.2000 708.4500 785.4000 708.6000 ;
	    RECT 779.4000 707.5500 785.4000 708.4500 ;
	    RECT 779.4000 707.4000 780.6000 707.5500 ;
	    RECT 784.2000 707.4000 785.4000 707.5500 ;
	    RECT 801.0000 706.5000 802.2000 719.7000 ;
	    RECT 803.4000 713.7000 804.6000 719.7000 ;
	    RECT 803.4000 709.5000 804.6000 709.8000 ;
	    RECT 823.5000 708.9000 824.7000 719.7000 ;
	    RECT 803.4000 708.4500 804.6000 708.6000 ;
	    RECT 808.2000 708.4500 809.4000 708.6000 ;
	    RECT 803.4000 707.5500 809.4000 708.4500 ;
	    RECT 823.5000 707.7000 826.2000 708.9000 ;
	    RECT 827.4000 707.7000 828.6000 719.7000 ;
	    RECT 846.6000 707.7000 847.8000 719.7000 ;
	    RECT 850.5000 708.9000 851.7000 719.7000 ;
	    RECT 858.6000 719.4000 859.8000 720.6000 ;
	    RECT 870.6000 713.7000 871.8000 719.7000 ;
	    RECT 849.0000 707.7000 851.7000 708.9000 ;
	    RECT 853.8000 708.4500 855.0000 708.6000 ;
	    RECT 870.6000 708.4500 871.8000 708.6000 ;
	    RECT 803.4000 707.4000 804.6000 707.5500 ;
	    RECT 808.2000 707.4000 809.4000 707.5500 ;
	    RECT 822.6000 706.5000 823.8000 706.8000 ;
	    RECT 741.0000 706.2000 742.2000 706.5000 ;
	    RECT 743.4000 704.4000 744.6000 705.6000 ;
	    RECT 745.5000 704.4000 745.8000 705.6000 ;
	    RECT 671.4000 701.4000 672.6000 702.6000 ;
	    RECT 671.4000 700.2000 672.6000 700.5000 ;
	    RECT 642.6000 699.0000 644.1000 700.2000 ;
	    RECT 673.8000 699.3000 675.0000 703.5000 ;
	    RECT 748.2000 702.6000 749.1000 706.5000 ;
	    RECT 772.2000 706.2000 773.4000 706.5000 ;
	    RECT 774.6000 704.4000 775.8000 705.6000 ;
	    RECT 776.7000 704.4000 777.0000 705.6000 ;
	    RECT 779.4000 702.6000 780.3000 706.5000 ;
	    RECT 801.0000 704.4000 802.2000 705.6000 ;
	    RECT 822.6000 704.4000 823.8000 705.6000 ;
	    RECT 825.0000 703.5000 825.9000 707.7000 ;
	    RECT 832.2000 705.4500 833.4000 705.6000 ;
	    RECT 846.6000 705.4500 847.8000 705.6000 ;
	    RECT 832.2000 704.5500 847.8000 705.4500 ;
	    RECT 832.2000 704.4000 833.4000 704.5500 ;
	    RECT 846.6000 704.4000 847.8000 704.5500 ;
	    RECT 849.3000 703.5000 850.2000 707.7000 ;
	    RECT 853.8000 707.5500 871.8000 708.4500 ;
	    RECT 853.8000 707.4000 855.0000 707.5500 ;
	    RECT 870.6000 707.4000 871.8000 707.5500 ;
	    RECT 851.4000 706.5000 852.6000 706.8000 ;
	    RECT 873.0000 706.5000 874.2000 719.7000 ;
	    RECT 875.4000 713.7000 876.6000 719.7000 ;
	    RECT 875.4000 709.5000 876.6000 709.8000 ;
	    RECT 875.4000 708.4500 876.6000 708.6000 ;
	    RECT 877.8000 708.4500 879.0000 708.6000 ;
	    RECT 904.2000 708.4500 905.4000 708.6000 ;
	    RECT 875.4000 707.5500 905.4000 708.4500 ;
	    RECT 911.4000 707.7000 912.6000 719.7000 ;
	    RECT 915.3000 707.7000 918.3000 719.7000 ;
	    RECT 921.0000 707.7000 922.2000 719.7000 ;
	    RECT 945.9000 713.7000 947.1000 719.7000 ;
	    RECT 946.2000 710.4000 947.4000 711.6000 ;
	    RECT 946.2000 709.5000 947.1000 710.4000 ;
	    RECT 948.3000 708.6000 949.5000 719.7000 ;
	    RECT 875.4000 707.4000 876.6000 707.5500 ;
	    RECT 877.8000 707.4000 879.0000 707.5500 ;
	    RECT 904.2000 707.4000 905.4000 707.5500 ;
	    RECT 851.4000 705.4500 852.6000 705.6000 ;
	    RECT 868.2000 705.4500 869.4000 705.6000 ;
	    RECT 851.4000 704.5500 869.4000 705.4500 ;
	    RECT 851.4000 704.4000 852.6000 704.5500 ;
	    RECT 868.2000 704.4000 869.4000 704.5500 ;
	    RECT 873.0000 705.4500 874.2000 705.6000 ;
	    RECT 880.2000 705.4500 881.4000 705.6000 ;
	    RECT 873.0000 704.5500 881.4000 705.4500 ;
	    RECT 873.0000 704.4000 874.2000 704.5500 ;
	    RECT 880.2000 704.4000 881.4000 704.5500 ;
	    RECT 913.8000 704.4000 915.0000 705.6000 ;
	    RECT 911.4000 703.5000 912.6000 703.8000 ;
	    RECT 916.5000 703.5000 917.4000 707.7000 ;
	    RECT 945.0000 707.4000 946.2000 708.6000 ;
	    RECT 948.0000 707.7000 949.5000 708.6000 ;
	    RECT 952.2000 707.7000 953.4000 719.7000 ;
	    RECT 918.6000 704.4000 919.8000 705.6000 ;
	    RECT 676.2000 702.4500 677.4000 702.6000 ;
	    RECT 697.8000 702.4500 699.0000 702.6000 ;
	    RECT 676.2000 701.5500 699.0000 702.4500 ;
	    RECT 676.2000 701.4000 677.4000 701.5500 ;
	    RECT 697.8000 701.4000 699.0000 701.5500 ;
	    RECT 717.0000 702.4500 718.2000 702.6000 ;
	    RECT 733.8000 702.4500 735.0000 702.6000 ;
	    RECT 717.0000 701.5500 735.0000 702.4500 ;
	    RECT 746.7000 702.3000 749.1000 702.6000 ;
	    RECT 777.9000 702.3000 780.3000 702.6000 ;
	    RECT 717.0000 701.4000 718.2000 701.5500 ;
	    RECT 733.8000 701.4000 735.0000 701.5500 ;
	    RECT 642.6000 693.3000 643.8000 699.0000 ;
	    RECT 645.0000 693.3000 646.2000 696.3000 ;
	    RECT 671.4000 693.3000 672.6000 699.3000 ;
	    RECT 673.8000 698.4000 676.5000 699.3000 ;
	    RECT 675.3000 693.3000 676.5000 698.4000 ;
	    RECT 697.8000 696.3000 698.7000 700.5000 ;
	    RECT 700.2000 699.4500 701.4000 699.6000 ;
	    RECT 709.8000 699.4500 711.0000 699.6000 ;
	    RECT 700.2000 698.5500 711.0000 699.4500 ;
	    RECT 700.2000 698.4000 701.4000 698.5500 ;
	    RECT 709.8000 698.4000 711.0000 698.5500 ;
	    RECT 714.6000 698.4000 715.8000 699.6000 ;
	    RECT 700.2000 697.2000 701.4000 697.5000 ;
	    RECT 714.6000 697.2000 715.8000 697.5000 ;
	    RECT 695.4000 693.3000 696.6000 696.3000 ;
	    RECT 697.8000 693.3000 699.0000 696.3000 ;
	    RECT 700.2000 693.3000 701.4000 696.3000 ;
	    RECT 714.6000 693.3000 715.8000 696.3000 ;
	    RECT 717.0000 693.3000 718.2000 700.5000 ;
	    RECT 741.0000 693.3000 742.2000 702.3000 ;
	    RECT 746.4000 701.7000 749.1000 702.3000 ;
	    RECT 746.4000 693.3000 747.6000 701.7000 ;
	    RECT 772.2000 693.3000 773.4000 702.3000 ;
	    RECT 777.6000 701.7000 780.3000 702.3000 ;
	    RECT 777.6000 693.3000 778.8000 701.7000 ;
	    RECT 798.6000 701.4000 799.8000 702.6000 ;
	    RECT 798.6000 700.2000 799.8000 700.5000 ;
	    RECT 801.0000 699.3000 802.2000 703.5000 ;
	    RECT 803.4000 702.4500 804.6000 702.6000 ;
	    RECT 825.0000 702.4500 826.2000 702.6000 ;
	    RECT 803.4000 701.5500 826.2000 702.4500 ;
	    RECT 803.4000 701.4000 804.6000 701.5500 ;
	    RECT 825.0000 701.4000 826.2000 701.5500 ;
	    RECT 829.8000 702.4500 831.0000 702.6000 ;
	    RECT 849.0000 702.4500 850.2000 702.6000 ;
	    RECT 829.8000 701.5500 850.2000 702.4500 ;
	    RECT 829.8000 701.4000 831.0000 701.5500 ;
	    RECT 849.0000 701.4000 850.2000 701.5500 ;
	    RECT 858.6000 702.4500 859.8000 702.6000 ;
	    RECT 870.6000 702.4500 871.8000 702.6000 ;
	    RECT 858.6000 701.5500 871.8000 702.4500 ;
	    RECT 858.6000 701.4000 859.8000 701.5500 ;
	    RECT 870.6000 701.4000 871.8000 701.5500 ;
	    RECT 798.6000 693.3000 799.8000 699.3000 ;
	    RECT 801.0000 698.4000 803.7000 699.3000 ;
	    RECT 802.5000 693.3000 803.7000 698.4000 ;
	    RECT 825.0000 696.3000 825.9000 700.5000 ;
	    RECT 827.4000 698.4000 828.6000 699.6000 ;
	    RECT 846.6000 698.4000 847.8000 699.6000 ;
	    RECT 827.4000 697.2000 828.6000 697.5000 ;
	    RECT 846.6000 697.2000 847.8000 697.5000 ;
	    RECT 849.3000 696.3000 850.2000 700.5000 ;
	    RECT 870.6000 700.2000 871.8000 700.5000 ;
	    RECT 873.0000 699.3000 874.2000 703.5000 ;
	    RECT 913.8000 703.2000 915.0000 703.5000 ;
	    RECT 918.6000 703.2000 919.8000 703.5000 ;
	    RECT 948.0000 702.6000 948.9000 707.7000 ;
	    RECT 949.8000 705.4500 951.0000 705.6000 ;
	    RECT 949.8000 704.5500 960.4500 705.4500 ;
	    RECT 949.8000 704.4000 951.0000 704.5500 ;
	    RECT 949.8000 703.2000 951.0000 703.5000 ;
	    RECT 875.4000 702.4500 876.6000 702.6000 ;
	    RECT 901.8000 702.4500 903.0000 702.6000 ;
	    RECT 875.4000 701.5500 903.0000 702.4500 ;
	    RECT 875.4000 701.4000 876.6000 701.5500 ;
	    RECT 901.8000 701.4000 903.0000 701.5500 ;
	    RECT 911.4000 701.4000 912.6000 702.6000 ;
	    RECT 913.8000 701.4000 915.3000 702.3000 ;
	    RECT 916.2000 701.4000 917.4000 702.6000 ;
	    RECT 913.8000 699.3000 914.7000 701.4000 ;
	    RECT 919.8000 700.8000 920.1000 702.3000 ;
	    RECT 921.0000 701.4000 922.2000 702.6000 ;
	    RECT 945.0000 701.4000 946.2000 702.6000 ;
	    RECT 947.1000 701.4000 948.9000 702.6000 ;
	    RECT 952.2000 702.4500 953.4000 702.6000 ;
	    RECT 954.6000 702.4500 955.8000 702.6000 ;
	    RECT 951.0000 700.8000 951.3000 702.3000 ;
	    RECT 952.2000 701.5500 955.8000 702.4500 ;
	    RECT 959.5500 702.4500 960.4500 704.5500 ;
	    RECT 966.6000 703.5000 967.8000 719.7000 ;
	    RECT 969.0000 713.7000 970.2000 719.7000 ;
	    RECT 983.4000 703.5000 984.6000 719.7000 ;
	    RECT 985.8000 713.7000 987.0000 719.7000 ;
	    RECT 1000.2000 713.7000 1001.4000 719.7000 ;
	    RECT 1002.6000 703.5000 1003.8000 719.7000 ;
	    RECT 1026.6000 707.7000 1027.8000 719.7000 ;
	    RECT 1030.5000 708.6000 1031.7001 719.7000 ;
	    RECT 1032.9000 713.7000 1034.1000 719.7000 ;
	    RECT 1165.8000 713.7000 1167.0000 719.7000 ;
	    RECT 1168.2001 712.5000 1169.4000 719.7000 ;
	    RECT 1170.6000 713.7000 1171.8000 719.7000 ;
	    RECT 1173.0000 712.8000 1174.2001 719.7000 ;
	    RECT 1175.4000 713.7000 1176.6000 719.7000 ;
	    RECT 1170.3000 711.9000 1174.2001 712.8000 ;
	    RECT 1032.6000 710.4000 1033.8000 711.6000 ;
	    RECT 1081.8000 711.4500 1083.0000 711.6000 ;
	    RECT 1151.4000 711.4500 1152.6000 711.6000 ;
	    RECT 1168.2001 711.4500 1169.4000 711.6000 ;
	    RECT 1081.8000 710.5500 1169.4000 711.4500 ;
	    RECT 1081.8000 710.4000 1083.0000 710.5500 ;
	    RECT 1151.4000 710.4000 1152.6000 710.5500 ;
	    RECT 1168.2001 710.4000 1169.4000 710.5500 ;
	    RECT 1032.9000 709.5000 1033.8000 710.4000 ;
	    RECT 1170.3000 709.5000 1171.2001 711.9000 ;
	    RECT 1177.8000 711.6000 1179.0000 719.7000 ;
	    RECT 1180.2001 713.7000 1181.4000 719.7000 ;
	    RECT 1182.6000 715.5000 1183.8000 719.7000 ;
	    RECT 1185.0000 715.5000 1186.2001 719.7000 ;
	    RECT 1187.4000 715.5000 1188.6000 719.7000 ;
	    RECT 1179.9000 711.6000 1186.2001 712.8000 ;
	    RECT 1175.1000 710.4000 1179.0000 711.6000 ;
	    RECT 1189.8000 710.4000 1191.0000 719.7000 ;
	    RECT 1192.2001 713.7000 1193.4000 719.7000 ;
	    RECT 1194.6000 712.5000 1195.8000 719.7000 ;
	    RECT 1197.0000 713.7000 1198.2001 719.7000 ;
	    RECT 1199.4000 712.5000 1200.6000 719.7000 ;
	    RECT 1201.8000 715.5000 1203.0000 719.7000 ;
	    RECT 1204.2001 715.5000 1205.4000 719.7000 ;
	    RECT 1206.6000 713.7000 1207.8000 719.7000 ;
	    RECT 1209.0000 712.8000 1210.2001 719.7000 ;
	    RECT 1211.4000 713.7000 1212.6000 720.6000 ;
	    RECT 1213.8000 714.6000 1215.0000 719.7000 ;
	    RECT 1213.8000 713.7000 1215.3000 714.6000 ;
	    RECT 1216.2001 713.7000 1217.4000 719.7000 ;
	    RECT 1242.6000 713.7000 1243.8000 719.7000 ;
	    RECT 1245.0000 714.3000 1246.2001 719.7000 ;
	    RECT 1214.4000 712.8000 1215.3000 713.7000 ;
	    RECT 1242.9000 713.4000 1243.8000 713.7000 ;
	    RECT 1247.4000 713.7000 1248.6000 719.7000 ;
	    RECT 1249.8000 713.7000 1251.0000 719.7000 ;
	    RECT 1247.4000 713.4000 1248.3000 713.7000 ;
	    RECT 1207.2001 711.6000 1213.5000 712.8000 ;
	    RECT 1214.4000 711.9000 1217.4000 712.8000 ;
	    RECT 1194.6000 710.4000 1198.5000 711.6000 ;
	    RECT 1199.4000 710.7000 1208.1000 711.6000 ;
	    RECT 1212.6000 711.0000 1213.5000 711.6000 ;
	    RECT 1182.6000 709.5000 1183.8000 709.8000 ;
	    RECT 1030.5000 707.7000 1032.0000 708.6000 ;
	    RECT 1029.0000 705.4500 1030.2001 705.6000 ;
	    RECT 1024.3500 704.5500 1030.2001 705.4500 ;
	    RECT 966.6000 702.4500 967.8000 702.6000 ;
	    RECT 959.5500 701.5500 967.8000 702.4500 ;
	    RECT 952.2000 701.4000 953.4000 701.5500 ;
	    RECT 954.6000 701.4000 955.8000 701.5500 ;
	    RECT 966.6000 701.4000 967.8000 701.5500 ;
	    RECT 969.0000 702.4500 970.2000 702.6000 ;
	    RECT 983.4000 702.4500 984.6000 702.6000 ;
	    RECT 969.0000 701.5500 984.6000 702.4500 ;
	    RECT 969.0000 701.4000 970.2000 701.5500 ;
	    RECT 983.4000 701.4000 984.6000 701.5500 ;
	    RECT 1002.6000 702.4500 1003.8000 702.6000 ;
	    RECT 1024.3500 702.4500 1025.2500 704.5500 ;
	    RECT 1029.0000 704.4000 1030.2001 704.5500 ;
	    RECT 1029.0000 703.2000 1030.2001 703.5000 ;
	    RECT 1031.1000 702.6000 1032.0000 707.7000 ;
	    RECT 1033.8000 708.4500 1035.0000 708.6000 ;
	    RECT 1072.2001 708.4500 1073.4000 708.6000 ;
	    RECT 1033.8000 707.5500 1073.4000 708.4500 ;
	    RECT 1168.2001 708.0000 1169.4000 709.5000 ;
	    RECT 1033.8000 707.4000 1035.0000 707.5500 ;
	    RECT 1072.2001 707.4000 1073.4000 707.5500 ;
	    RECT 1167.9000 706.8000 1169.4000 708.0000 ;
	    RECT 1170.3000 708.6000 1183.8000 709.5000 ;
	    RECT 1187.4000 709.5000 1188.6000 709.8000 ;
	    RECT 1199.4000 709.5000 1200.3000 710.7000 ;
	    RECT 1209.0000 709.8000 1211.1000 710.7000 ;
	    RECT 1212.6000 709.8000 1215.0000 711.0000 ;
	    RECT 1187.4000 708.6000 1200.3000 709.5000 ;
	    RECT 1201.8000 709.5000 1211.1000 709.8000 ;
	    RECT 1201.8000 708.9000 1209.9000 709.5000 ;
	    RECT 1201.8000 708.6000 1203.0000 708.9000 ;
	    RECT 1002.6000 701.5500 1025.2500 702.4500 ;
	    RECT 1002.6000 701.4000 1003.8000 701.5500 ;
	    RECT 1026.6000 701.4000 1027.8000 702.6000 ;
	    RECT 1028.7001 700.8000 1029.0000 702.3000 ;
	    RECT 1031.1000 701.4000 1032.9000 702.6000 ;
	    RECT 1033.8000 702.4500 1035.0000 702.6000 ;
	    RECT 1110.6000 702.4500 1111.8000 702.6000 ;
	    RECT 1033.8000 701.5500 1111.8000 702.4500 ;
	    RECT 1033.8000 701.4000 1035.0000 701.5500 ;
	    RECT 1110.6000 701.4000 1111.8000 701.5500 ;
	    RECT 916.5000 699.3000 921.9000 699.9000 ;
	    RECT 945.3000 699.3000 946.2000 700.5000 ;
	    RECT 947.7000 699.3000 953.1000 699.9000 ;
	    RECT 822.6000 693.3000 823.8000 696.3000 ;
	    RECT 825.0000 693.3000 826.2000 696.3000 ;
	    RECT 827.4000 693.3000 828.6000 696.3000 ;
	    RECT 846.6000 693.3000 847.8000 696.3000 ;
	    RECT 849.0000 693.3000 850.2000 696.3000 ;
	    RECT 851.4000 693.3000 852.6000 696.3000 ;
	    RECT 870.6000 693.3000 871.8000 699.3000 ;
	    RECT 873.0000 698.4000 875.7000 699.3000 ;
	    RECT 874.5000 693.3000 875.7000 698.4000 ;
	    RECT 911.4000 694.2000 912.6000 699.3000 ;
	    RECT 913.8000 695.1000 915.0000 699.3000 ;
	    RECT 916.2000 699.0000 922.2000 699.3000 ;
	    RECT 916.2000 694.2000 917.4000 699.0000 ;
	    RECT 911.4000 693.3000 917.4000 694.2000 ;
	    RECT 918.6000 693.3000 919.8000 698.1000 ;
	    RECT 921.0000 693.3000 922.2000 699.0000 ;
	    RECT 945.0000 693.3000 946.2000 699.3000 ;
	    RECT 947.4000 699.0000 953.4000 699.3000 ;
	    RECT 947.4000 693.3000 948.6000 699.0000 ;
	    RECT 949.8000 693.3000 951.0000 698.1000 ;
	    RECT 952.2000 693.3000 953.4000 699.0000 ;
	    RECT 966.6000 693.3000 967.8000 700.5000 ;
	    RECT 969.0000 699.4500 970.2000 699.6000 ;
	    RECT 978.6000 699.4500 979.8000 699.6000 ;
	    RECT 969.0000 698.5500 979.8000 699.4500 ;
	    RECT 969.0000 698.4000 970.2000 698.5500 ;
	    RECT 978.6000 698.4000 979.8000 698.5500 ;
	    RECT 969.0000 697.2000 970.2000 697.5000 ;
	    RECT 969.0000 693.3000 970.2000 696.3000 ;
	    RECT 983.4000 693.3000 984.6000 700.5000 ;
	    RECT 985.8000 698.4000 987.0000 699.6000 ;
	    RECT 988.2000 699.4500 989.4000 699.6000 ;
	    RECT 1000.2000 699.4500 1001.4000 699.6000 ;
	    RECT 988.2000 698.5500 1001.4000 699.4500 ;
	    RECT 988.2000 698.4000 989.4000 698.5500 ;
	    RECT 1000.2000 698.4000 1001.4000 698.5500 ;
	    RECT 985.8000 697.2000 987.0000 697.5000 ;
	    RECT 1000.2000 697.2000 1001.4000 697.5000 ;
	    RECT 985.8000 693.3000 987.0000 696.3000 ;
	    RECT 1000.2000 693.3000 1001.4000 696.3000 ;
	    RECT 1002.6000 693.3000 1003.8000 700.5000 ;
	    RECT 1026.9000 699.3000 1032.3000 699.9000 ;
	    RECT 1033.8000 699.3000 1034.7001 700.5000 ;
	    RECT 1167.9000 700.2000 1169.1000 706.8000 ;
	    RECT 1170.3000 705.9000 1171.2001 708.6000 ;
	    RECT 1206.3000 707.7000 1207.5000 708.0000 ;
	    RECT 1172.1000 706.8000 1210.5000 707.7000 ;
	    RECT 1211.4000 707.4000 1212.6000 708.6000 ;
	    RECT 1172.1000 706.5000 1173.3000 706.8000 ;
	    RECT 1170.0000 705.0000 1171.2001 705.9000 ;
	    RECT 1180.2001 705.0000 1205.7001 705.9000 ;
	    RECT 1170.0000 702.0000 1170.9000 705.0000 ;
	    RECT 1180.2001 704.1000 1181.4000 705.0000 ;
	    RECT 1206.6000 704.4000 1207.8000 705.6000 ;
	    RECT 1208.7001 705.0000 1215.3000 705.9000 ;
	    RECT 1214.1000 704.7000 1215.3000 705.0000 ;
	    RECT 1171.8000 702.9000 1177.5000 704.1000 ;
	    RECT 1170.0000 701.1000 1171.8000 702.0000 ;
	    RECT 1026.6000 699.0000 1032.6000 699.3000 ;
	    RECT 1026.6000 693.3000 1027.8000 699.0000 ;
	    RECT 1029.0000 693.3000 1030.2001 698.1000 ;
	    RECT 1031.4000 693.3000 1032.6000 699.0000 ;
	    RECT 1033.8000 693.3000 1035.0000 699.3000 ;
	    RECT 1167.9000 699.0000 1169.4000 700.2000 ;
	    RECT 1165.8000 693.3000 1167.0000 696.3000 ;
	    RECT 1168.2001 693.3000 1169.4000 699.0000 ;
	    RECT 1170.6000 693.3000 1171.8000 701.1000 ;
	    RECT 1176.3000 701.1000 1177.5000 702.9000 ;
	    RECT 1176.3000 700.2000 1179.0000 701.1000 ;
	    RECT 1177.8000 699.3000 1179.0000 700.2000 ;
	    RECT 1185.0000 699.6000 1186.2001 703.8000 ;
	    RECT 1189.8000 702.9000 1194.6000 704.1000 ;
	    RECT 1200.3000 702.9000 1203.3000 704.1000 ;
	    RECT 1216.2001 703.5000 1217.4000 711.9000 ;
	    RECT 1242.9000 712.5000 1248.3000 713.4000 ;
	    RECT 1242.9000 709.5000 1243.8000 712.5000 ;
	    RECT 1245.0000 710.4000 1246.2001 711.6000 ;
	    RECT 1245.0000 709.2000 1246.2001 709.5000 ;
	    RECT 1242.6000 707.4000 1243.8000 708.6000 ;
	    RECT 1249.8000 708.4500 1251.0000 708.6000 ;
	    RECT 1249.8000 707.5500 1253.2500 708.4500 ;
	    RECT 1269.0000 707.7000 1270.2001 719.7000 ;
	    RECT 1272.9000 708.9000 1274.1000 719.7000 ;
	    RECT 1297.8000 713.7000 1299.0000 719.7000 ;
	    RECT 1300.2001 713.7000 1301.4000 719.7000 ;
	    RECT 1302.6000 714.3000 1303.8000 719.7000 ;
	    RECT 1300.5000 713.4000 1301.4000 713.7000 ;
	    RECT 1305.0000 713.7000 1306.2001 719.7000 ;
	    RECT 1305.0000 713.4000 1305.9000 713.7000 ;
	    RECT 1300.5000 712.5000 1305.9000 713.4000 ;
	    RECT 1302.6000 710.4000 1303.8000 711.6000 ;
	    RECT 1305.0000 709.5000 1305.9000 712.5000 ;
	    RECT 1302.6000 709.2000 1303.8000 709.5000 ;
	    RECT 1271.4000 707.7000 1274.1000 708.9000 ;
	    RECT 1329.9000 708.6000 1331.1000 719.7000 ;
	    RECT 1249.8000 707.4000 1251.0000 707.5500 ;
	    RECT 1189.2001 701.7000 1190.4000 702.0000 ;
	    RECT 1189.2001 700.8000 1195.8000 701.7000 ;
	    RECT 1197.0000 701.4000 1198.2001 702.6000 ;
	    RECT 1194.6000 700.5000 1195.8000 700.8000 ;
	    RECT 1197.0000 700.2000 1198.2001 700.5000 ;
	    RECT 1175.4000 693.3000 1176.6000 699.3000 ;
	    RECT 1177.8000 698.1000 1181.4000 699.3000 ;
	    RECT 1185.0000 698.4000 1186.5000 699.6000 ;
	    RECT 1191.0000 698.4000 1191.3000 699.6000 ;
	    RECT 1192.2001 698.4000 1193.4000 699.6000 ;
	    RECT 1194.6000 699.3000 1195.8000 699.6000 ;
	    RECT 1200.3000 699.3000 1201.5000 702.9000 ;
	    RECT 1204.2001 702.3000 1217.4000 703.5000 ;
	    RECT 1209.3000 700.2000 1213.8000 701.4000 ;
	    RECT 1209.3000 699.3000 1210.5000 700.2000 ;
	    RECT 1194.6000 698.4000 1201.5000 699.3000 ;
	    RECT 1180.2001 693.3000 1181.4000 698.1000 ;
	    RECT 1206.6000 698.1000 1210.5000 699.3000 ;
	    RECT 1182.6000 693.3000 1183.8000 697.5000 ;
	    RECT 1185.0000 693.3000 1186.2001 697.5000 ;
	    RECT 1187.4000 693.3000 1188.6000 697.5000 ;
	    RECT 1189.8000 693.3000 1191.0000 697.5000 ;
	    RECT 1192.2001 693.3000 1193.4000 696.3000 ;
	    RECT 1194.6000 693.3000 1195.8000 697.5000 ;
	    RECT 1197.0000 693.3000 1198.2001 696.3000 ;
	    RECT 1199.4000 693.3000 1200.6000 697.5000 ;
	    RECT 1201.8000 693.3000 1203.0000 697.5000 ;
	    RECT 1204.2001 693.3000 1205.4000 697.5000 ;
	    RECT 1206.6000 693.3000 1207.8000 698.1000 ;
	    RECT 1211.4000 693.3000 1212.6000 699.3000 ;
	    RECT 1216.2001 693.3000 1217.4000 702.3000 ;
	    RECT 1242.9000 702.6000 1243.8000 706.5000 ;
	    RECT 1249.8000 706.2000 1251.0000 706.5000 ;
	    RECT 1246.2001 704.4000 1246.5000 705.6000 ;
	    RECT 1247.4000 704.4000 1248.6000 705.6000 ;
	    RECT 1242.9000 702.3000 1245.3000 702.6000 ;
	    RECT 1252.3500 702.4500 1253.2500 707.5500 ;
	    RECT 1271.7001 703.5000 1272.6000 707.7000 ;
	    RECT 1297.8000 707.4000 1299.0000 708.6000 ;
	    RECT 1305.0000 708.4500 1306.2001 708.6000 ;
	    RECT 1317.0000 708.4500 1318.2001 708.6000 ;
	    RECT 1305.0000 707.5500 1318.2001 708.4500 ;
	    RECT 1305.0000 707.4000 1306.2001 707.5500 ;
	    RECT 1317.0000 707.4000 1318.2001 707.5500 ;
	    RECT 1329.0000 707.7000 1331.1000 708.6000 ;
	    RECT 1332.3000 707.7000 1333.5000 719.7000 ;
	    RECT 1273.8000 706.5000 1275.0000 706.8000 ;
	    RECT 1329.0000 706.5000 1329.9000 707.7000 ;
	    RECT 1336.2001 706.8000 1337.4000 719.7000 ;
	    RECT 1386.6000 708.6000 1387.8000 719.7000 ;
	    RECT 1389.0000 709.8000 1390.5000 719.7000 ;
	    RECT 1389.3000 708.6000 1390.5000 708.9000 ;
	    RECT 1386.6000 707.7000 1390.5000 708.6000 ;
	    RECT 1393.2001 707.7000 1395.6000 719.7000 ;
	    RECT 1398.3000 709.8000 1399.8000 719.7000 ;
	    RECT 1398.6000 708.6000 1399.8000 708.9000 ;
	    RECT 1401.0000 708.6000 1402.2001 719.7000 ;
	    RECT 1420.2001 713.7000 1421.4000 719.7000 ;
	    RECT 1420.2001 709.5000 1421.4000 709.8000 ;
	    RECT 1398.6000 707.7000 1402.2001 708.6000 ;
	    RECT 1297.8000 706.2000 1299.0000 706.5000 ;
	    RECT 1273.8000 704.4000 1275.0000 705.6000 ;
	    RECT 1300.2001 704.4000 1301.4000 705.6000 ;
	    RECT 1302.3000 704.4000 1302.6000 705.6000 ;
	    RECT 1305.0000 702.6000 1305.9000 706.5000 ;
	    RECT 1331.4000 706.2000 1337.4000 706.8000 ;
	    RECT 1394.1000 706.5000 1395.0000 707.7000 ;
	    RECT 1420.2001 707.4000 1421.4000 708.6000 ;
	    RECT 1422.6000 706.5000 1423.8000 719.7000 ;
	    RECT 1425.0000 713.7000 1426.2001 719.7000 ;
	    RECT 1449.0000 708.6000 1450.2001 719.7000 ;
	    RECT 1451.4000 709.5000 1452.6000 719.7000 ;
	    RECT 1453.8000 708.6000 1455.0000 719.7000 ;
	    RECT 1449.0000 707.7000 1455.0000 708.6000 ;
	    RECT 1456.2001 707.7000 1457.4000 719.7000 ;
	    RECT 1480.2001 713.7000 1481.4000 719.7000 ;
	    RECT 1482.6000 713.7000 1483.8000 719.7000 ;
	    RECT 1485.0000 714.3000 1486.2001 719.7000 ;
	    RECT 1482.9000 713.4000 1483.8000 713.7000 ;
	    RECT 1487.4000 713.7000 1488.6000 719.7000 ;
	    RECT 1506.6000 713.7000 1507.8000 719.7000 ;
	    RECT 1487.4000 713.4000 1488.3000 713.7000 ;
	    RECT 1482.9000 712.5000 1488.3000 713.4000 ;
	    RECT 1480.2001 711.4500 1481.4000 711.6000 ;
	    RECT 1485.0000 711.4500 1486.2001 711.6000 ;
	    RECT 1480.2001 710.5500 1486.2001 711.4500 ;
	    RECT 1480.2001 710.4000 1481.4000 710.5500 ;
	    RECT 1485.0000 710.4000 1486.2001 710.5500 ;
	    RECT 1487.4000 709.5000 1488.3000 712.5000 ;
	    RECT 1485.0000 709.2000 1486.2001 709.5000 ;
	    RECT 1475.4000 708.4500 1476.6000 708.6000 ;
	    RECT 1480.2001 708.4500 1481.4000 708.6000 ;
	    RECT 1456.2001 706.5000 1457.1000 707.7000 ;
	    RECT 1475.4000 707.5500 1481.4000 708.4500 ;
	    RECT 1475.4000 707.4000 1476.6000 707.5500 ;
	    RECT 1480.2001 707.4000 1481.4000 707.5500 ;
	    RECT 1487.4000 708.4500 1488.6000 708.6000 ;
	    RECT 1506.6000 708.4500 1507.8000 708.6000 ;
	    RECT 1487.4000 707.5500 1507.8000 708.4500 ;
	    RECT 1487.4000 707.4000 1488.6000 707.5500 ;
	    RECT 1506.6000 707.4000 1507.8000 707.5500 ;
	    RECT 1509.0000 706.5000 1510.2001 719.7000 ;
	    RECT 1511.4000 713.7000 1512.6000 719.7000 ;
	    RECT 1511.4000 709.5000 1512.6000 709.8000 ;
	    RECT 1511.4000 707.4000 1512.6000 708.6000 ;
	    RECT 1535.4000 707.7000 1536.6000 719.7000 ;
	    RECT 1539.3000 708.6000 1540.5000 719.7000 ;
	    RECT 1541.7001 713.7000 1542.9000 719.7000 ;
	    RECT 1561.8000 713.7000 1563.0000 719.7000 ;
	    RECT 1541.4000 710.4000 1542.6000 711.6000 ;
	    RECT 1541.7001 709.5000 1542.6000 710.4000 ;
	    RECT 1539.3000 707.7000 1540.8000 708.6000 ;
	    RECT 1480.2001 706.2000 1481.4000 706.5000 ;
	    RECT 1331.1000 705.9000 1337.4000 706.2000 ;
	    RECT 1309.8000 705.4500 1311.0000 705.6000 ;
	    RECT 1329.0000 705.4500 1330.2001 705.6000 ;
	    RECT 1309.8000 704.5500 1330.2001 705.4500 ;
	    RECT 1309.8000 704.4000 1311.0000 704.5500 ;
	    RECT 1329.0000 704.4000 1330.2001 704.5500 ;
	    RECT 1331.1000 705.0000 1332.3000 705.9000 ;
	    RECT 1391.1000 705.6000 1392.3000 705.9000 ;
	    RECT 1271.4000 702.4500 1272.6000 702.6000 ;
	    RECT 1242.9000 701.7000 1245.6000 702.3000 ;
	    RECT 1244.4000 693.3000 1245.6000 701.7000 ;
	    RECT 1249.8000 693.3000 1251.0000 702.3000 ;
	    RECT 1252.3500 701.5500 1272.6000 702.4500 ;
	    RECT 1303.5000 702.3000 1305.9000 702.6000 ;
	    RECT 1271.4000 701.4000 1272.6000 701.5500 ;
	    RECT 1269.0000 698.4000 1270.2001 699.6000 ;
	    RECT 1269.0000 697.2000 1270.2001 697.5000 ;
	    RECT 1271.7001 696.3000 1272.6000 700.5000 ;
	    RECT 1269.0000 693.3000 1270.2001 696.3000 ;
	    RECT 1271.4000 693.3000 1272.6000 696.3000 ;
	    RECT 1273.8000 693.3000 1275.0000 696.3000 ;
	    RECT 1297.8000 693.3000 1299.0000 702.3000 ;
	    RECT 1303.2001 701.7000 1305.9000 702.3000 ;
	    RECT 1303.2001 693.3000 1304.4000 701.7000 ;
	    RECT 1329.0000 699.3000 1329.9000 703.5000 ;
	    RECT 1331.1000 700.5000 1332.0000 705.0000 ;
	    RECT 1389.9000 704.7000 1392.3000 705.6000 ;
	    RECT 1389.9000 704.4000 1391.1000 704.7000 ;
	    RECT 1393.8000 704.4000 1395.0000 705.6000 ;
	    RECT 1415.4000 705.4500 1416.6000 705.6000 ;
	    RECT 1422.6000 705.4500 1423.8000 705.6000 ;
	    RECT 1415.4000 704.5500 1423.8000 705.4500 ;
	    RECT 1415.4000 704.4000 1416.6000 704.5500 ;
	    RECT 1422.6000 704.4000 1423.8000 704.5500 ;
	    RECT 1449.0000 704.4000 1450.2001 705.6000 ;
	    RECT 1451.1000 704.7000 1451.4000 706.2000 ;
	    RECT 1453.8000 704.7000 1455.3000 705.6000 ;
	    RECT 1456.2001 705.4500 1457.4000 705.6000 ;
	    RECT 1477.8000 705.4500 1479.0000 705.6000 ;
	    RECT 1333.2001 703.5000 1334.4000 703.8000 ;
	    RECT 1451.4000 703.5000 1452.6000 703.8000 ;
	    RECT 1392.0000 702.9000 1393.2001 703.2000 ;
	    RECT 1389.0000 702.6000 1393.2001 702.9000 ;
	    RECT 1333.8000 702.4500 1335.0000 702.6000 ;
	    RECT 1345.8000 702.4500 1347.0000 702.6000 ;
	    RECT 1333.8000 701.5500 1347.0000 702.4500 ;
	    RECT 1333.8000 701.4000 1335.0000 701.5500 ;
	    RECT 1345.8000 701.4000 1347.0000 701.5500 ;
	    RECT 1369.8000 702.4500 1371.0000 702.6000 ;
	    RECT 1386.6000 702.4500 1387.8000 702.6000 ;
	    RECT 1369.8000 701.5500 1387.8000 702.4500 ;
	    RECT 1369.8000 701.4000 1371.0000 701.5500 ;
	    RECT 1386.6000 701.4000 1387.8000 701.5500 ;
	    RECT 1388.7001 702.0000 1393.2001 702.6000 ;
	    RECT 1394.1000 702.6000 1395.0000 703.5000 ;
	    RECT 1388.7001 701.7000 1389.9000 702.0000 ;
	    RECT 1394.1000 701.7000 1395.6000 702.6000 ;
	    RECT 1388.7001 701.4000 1389.0000 701.7000 ;
	    RECT 1331.1000 699.6000 1334.7001 700.5000 ;
	    RECT 1389.3000 700.2000 1390.5000 700.5000 ;
	    RECT 1329.0000 693.3000 1330.2001 699.3000 ;
	    RECT 1331.4000 693.3000 1332.6000 698.7000 ;
	    RECT 1333.8000 696.3000 1334.7001 699.6000 ;
	    RECT 1336.2001 699.4500 1337.4000 699.6000 ;
	    RECT 1369.8000 699.4500 1371.0000 699.6000 ;
	    RECT 1384.2001 699.4500 1385.4000 699.6000 ;
	    RECT 1336.2001 698.5500 1385.4000 699.4500 ;
	    RECT 1336.2001 698.4000 1337.4000 698.5500 ;
	    RECT 1369.8000 698.4000 1371.0000 698.5500 ;
	    RECT 1384.2001 698.4000 1385.4000 698.5500 ;
	    RECT 1386.6000 699.3000 1390.5000 700.2000 ;
	    RECT 1391.4000 699.6000 1393.8000 700.8000 ;
	    RECT 1336.2001 697.2000 1337.4000 697.5000 ;
	    RECT 1333.8000 693.3000 1335.0000 696.3000 ;
	    RECT 1336.2001 693.3000 1337.4000 696.3000 ;
	    RECT 1386.6000 693.3000 1387.8000 699.3000 ;
	    RECT 1394.7001 698.7000 1395.6000 701.7000 ;
	    RECT 1396.8000 701.4000 1398.0000 702.6000 ;
	    RECT 1399.8000 701.4000 1400.1000 702.6000 ;
	    RECT 1401.0000 701.4000 1402.2001 702.6000 ;
	    RECT 1396.8000 700.8000 1397.7001 701.4000 ;
	    RECT 1396.5000 699.6000 1397.7001 700.8000 ;
	    RECT 1398.6000 700.2000 1399.8000 700.5000 ;
	    RECT 1398.6000 699.3000 1402.2001 700.2000 ;
	    RECT 1422.6000 699.3000 1423.8000 703.5000 ;
	    RECT 1425.0000 702.4500 1426.2001 702.6000 ;
	    RECT 1449.0000 702.4500 1450.2001 702.6000 ;
	    RECT 1425.0000 701.5500 1450.2001 702.4500 ;
	    RECT 1425.0000 701.4000 1426.2001 701.5500 ;
	    RECT 1449.0000 701.4000 1450.2001 701.5500 ;
	    RECT 1451.4000 701.4000 1452.6000 702.6000 ;
	    RECT 1425.0000 700.2000 1426.2001 700.5000 ;
	    RECT 1453.8000 699.3000 1454.7001 704.7000 ;
	    RECT 1456.2001 704.5500 1479.0000 705.4500 ;
	    RECT 1456.2001 704.4000 1457.4000 704.5500 ;
	    RECT 1477.8000 704.4000 1479.0000 704.5500 ;
	    RECT 1482.6000 704.4000 1483.8000 705.6000 ;
	    RECT 1484.7001 704.4000 1485.0000 705.6000 ;
	    RECT 1487.4000 702.6000 1488.3000 706.5000 ;
	    RECT 1509.0000 705.4500 1510.2001 705.6000 ;
	    RECT 1525.8000 705.4500 1527.0000 705.6000 ;
	    RECT 1509.0000 704.5500 1527.0000 705.4500 ;
	    RECT 1509.0000 704.4000 1510.2001 704.5500 ;
	    RECT 1525.8000 704.4000 1527.0000 704.5500 ;
	    RECT 1537.8000 704.4000 1539.0000 705.6000 ;
	    RECT 1485.9000 702.3000 1488.3000 702.6000 ;
	    RECT 1389.0000 693.3000 1390.5000 698.4000 ;
	    RECT 1393.2001 693.3000 1395.6000 698.7000 ;
	    RECT 1398.3000 693.3000 1399.8000 698.4000 ;
	    RECT 1401.0000 693.3000 1402.2001 699.3000 ;
	    RECT 1421.1000 698.4000 1423.8000 699.3000 ;
	    RECT 1421.1000 693.3000 1422.3000 698.4000 ;
	    RECT 1425.0000 693.3000 1426.2001 699.3000 ;
	    RECT 1449.9000 693.3000 1451.1000 699.3000 ;
	    RECT 1453.8000 693.3000 1455.0000 699.3000 ;
	    RECT 1456.2001 698.4000 1457.4000 699.6000 ;
	    RECT 1455.9000 697.2000 1457.1000 697.5000 ;
	    RECT 1456.2001 693.3000 1457.4000 696.3000 ;
	    RECT 1480.2001 693.3000 1481.4000 702.3000 ;
	    RECT 1485.6000 701.7000 1488.3000 702.3000 ;
	    RECT 1489.8000 702.4500 1491.0000 702.6000 ;
	    RECT 1506.6000 702.4500 1507.8000 702.6000 ;
	    RECT 1485.6000 693.3000 1486.8000 701.7000 ;
	    RECT 1489.8000 701.5500 1507.8000 702.4500 ;
	    RECT 1489.8000 701.4000 1491.0000 701.5500 ;
	    RECT 1506.6000 701.4000 1507.8000 701.5500 ;
	    RECT 1506.6000 700.2000 1507.8000 700.5000 ;
	    RECT 1509.0000 699.3000 1510.2001 703.5000 ;
	    RECT 1537.8000 703.2000 1539.0000 703.5000 ;
	    RECT 1539.9000 702.6000 1540.8000 707.7000 ;
	    RECT 1542.6000 707.4000 1543.8000 708.6000 ;
	    RECT 1564.2001 706.5000 1565.4000 719.7000 ;
	    RECT 1566.6000 713.7000 1567.8000 719.7000 ;
	    RECT 1566.6000 709.5000 1567.8000 709.8000 ;
	    RECT 1545.0000 705.4500 1546.2001 705.6000 ;
	    RECT 1564.2001 705.4500 1565.4000 705.6000 ;
	    RECT 1545.0000 704.5500 1565.4000 705.4500 ;
	    RECT 1545.0000 704.4000 1546.2001 704.5500 ;
	    RECT 1564.2001 704.4000 1565.4000 704.5500 ;
	    RECT 1523.4000 702.4500 1524.6000 702.6000 ;
	    RECT 1535.4000 702.4500 1536.6000 702.6000 ;
	    RECT 1523.4000 701.5500 1536.6000 702.4500 ;
	    RECT 1523.4000 701.4000 1524.6000 701.5500 ;
	    RECT 1535.4000 701.4000 1536.6000 701.5500 ;
	    RECT 1537.5000 700.8000 1537.8000 702.3000 ;
	    RECT 1539.9000 701.4000 1541.7001 702.6000 ;
	    RECT 1542.6000 702.4500 1543.8000 702.6000 ;
	    RECT 1554.6000 702.4500 1555.8000 702.6000 ;
	    RECT 1542.6000 701.5500 1555.8000 702.4500 ;
	    RECT 1542.6000 701.4000 1543.8000 701.5500 ;
	    RECT 1554.6000 701.4000 1555.8000 701.5500 ;
	    RECT 1561.8000 701.4000 1563.0000 702.6000 ;
	    RECT 1535.7001 699.3000 1541.1000 699.9000 ;
	    RECT 1542.6000 699.3000 1543.5000 700.5000 ;
	    RECT 1561.8000 700.2000 1563.0000 700.5000 ;
	    RECT 1564.2001 699.3000 1565.4000 703.5000 ;
	    RECT 1506.6000 693.3000 1507.8000 699.3000 ;
	    RECT 1509.0000 698.4000 1511.7001 699.3000 ;
	    RECT 1510.5000 693.3000 1511.7001 698.4000 ;
	    RECT 1535.4000 699.0000 1541.4000 699.3000 ;
	    RECT 1535.4000 693.3000 1536.6000 699.0000 ;
	    RECT 1537.8000 693.3000 1539.0000 698.1000 ;
	    RECT 1540.2001 693.3000 1541.4000 699.0000 ;
	    RECT 1542.6000 693.3000 1543.8000 699.3000 ;
	    RECT 1561.8000 693.3000 1563.0000 699.3000 ;
	    RECT 1564.2001 698.4000 1566.9000 699.3000 ;
	    RECT 1565.7001 693.3000 1566.9000 698.4000 ;
	    RECT 1.2000 690.6000 1569.0000 692.4000 ;
	    RECT 52.2000 683.7000 53.4000 689.7000 ;
	    RECT 54.6000 682.8000 55.8000 689.7000 ;
	    RECT 57.0000 683.7000 58.2000 689.7000 ;
	    RECT 59.4000 682.8000 60.6000 689.7000 ;
	    RECT 61.8000 683.7000 63.0000 689.7000 ;
	    RECT 64.2000 682.8000 65.4000 689.7000 ;
	    RECT 66.6000 683.7000 67.8000 689.7000 ;
	    RECT 69.0000 682.8000 70.2000 689.7000 ;
	    RECT 71.4000 683.7000 72.6000 689.7000 ;
	    RECT 95.4000 683.7000 96.6000 689.7000 ;
	    RECT 97.8000 684.0000 99.0000 689.7000 ;
	    RECT 100.2000 684.9000 101.4000 689.7000 ;
	    RECT 102.6000 684.0000 103.8000 689.7000 ;
	    RECT 97.8000 683.7000 103.8000 684.0000 ;
	    RECT 54.6000 681.6000 57.3000 682.8000 ;
	    RECT 59.4000 681.6000 62.7000 682.8000 ;
	    RECT 64.2000 681.6000 67.5000 682.8000 ;
	    RECT 69.0000 681.6000 72.6000 682.8000 ;
	    RECT 95.7000 682.5000 96.6000 683.7000 ;
	    RECT 98.1000 683.1000 103.5000 683.7000 ;
	    RECT 117.0000 682.5000 118.2000 689.7000 ;
	    RECT 119.4000 686.7000 120.6000 689.7000 ;
	    RECT 119.4000 685.5000 120.6000 685.8000 ;
	    RECT 119.4000 684.4500 120.6000 684.6000 ;
	    RECT 121.8000 684.4500 123.0000 684.6000 ;
	    RECT 133.8000 684.4500 135.0000 684.6000 ;
	    RECT 119.4000 683.5500 135.0000 684.4500 ;
	    RECT 150.6000 684.0000 151.8000 689.7000 ;
	    RECT 153.0000 684.9000 154.2000 689.7000 ;
	    RECT 155.4000 688.8000 161.4000 689.7000 ;
	    RECT 155.4000 684.0000 156.6000 688.8000 ;
	    RECT 150.6000 683.7000 156.6000 684.0000 ;
	    RECT 157.8000 683.7000 159.0000 687.9000 ;
	    RECT 160.2000 683.7000 161.4000 688.8000 ;
	    RECT 174.6000 686.7000 175.8000 689.7000 ;
	    RECT 174.6000 685.5000 175.8000 685.8000 ;
	    RECT 162.6000 684.4500 163.8000 684.6000 ;
	    RECT 174.6000 684.4500 175.8000 684.6000 ;
	    RECT 119.4000 683.4000 120.6000 683.5500 ;
	    RECT 121.8000 683.4000 123.0000 683.5500 ;
	    RECT 133.8000 683.4000 135.0000 683.5500 ;
	    RECT 150.9000 683.1000 156.3000 683.7000 ;
	    RECT 49.8000 681.4500 51.0000 681.6000 ;
	    RECT 52.2000 681.4500 53.4000 681.6000 ;
	    RECT 49.8000 680.5500 53.4000 681.4500 ;
	    RECT 56.1000 680.7000 57.3000 681.6000 ;
	    RECT 61.5000 680.7000 62.7000 681.6000 ;
	    RECT 66.3000 680.7000 67.5000 681.6000 ;
	    RECT 49.8000 680.4000 51.0000 680.5500 ;
	    RECT 52.2000 680.4000 53.4000 680.5500 ;
	    RECT 54.3000 679.5000 54.9000 680.7000 ;
	    RECT 56.1000 679.5000 60.0000 680.7000 ;
	    RECT 61.5000 679.5000 65.1000 680.7000 ;
	    RECT 66.3000 679.5000 70.2000 680.7000 ;
	    RECT 71.4000 679.5000 72.6000 681.6000 ;
	    RECT 95.4000 680.4000 96.6000 681.6000 ;
	    RECT 97.5000 680.4000 99.3000 681.6000 ;
	    RECT 101.4000 680.7000 101.7000 682.2000 ;
	    RECT 102.6000 680.4000 103.8000 681.6000 ;
	    RECT 117.0000 681.4500 118.2000 681.6000 ;
	    RECT 105.1500 680.5500 118.2000 681.4500 ;
	    RECT 56.1000 677.4000 57.3000 679.5000 ;
	    RECT 61.5000 677.4000 62.7000 679.5000 ;
	    RECT 66.3000 677.4000 67.5000 679.5000 ;
	    RECT 71.4000 678.4500 72.6000 678.6000 ;
	    RECT 93.0000 678.4500 94.2000 678.6000 ;
	    RECT 71.4000 677.5500 94.2000 678.4500 ;
	    RECT 71.4000 677.4000 72.6000 677.5500 ;
	    RECT 93.0000 677.4000 94.2000 677.5500 ;
	    RECT 54.6000 676.2000 57.3000 677.4000 ;
	    RECT 59.4000 676.2000 62.7000 677.4000 ;
	    RECT 64.2000 676.2000 67.5000 677.4000 ;
	    RECT 69.0000 676.5000 70.5000 677.4000 ;
	    RECT 69.0000 676.2000 72.6000 676.5000 ;
	    RECT 52.2000 663.3000 53.4000 675.3000 ;
	    RECT 54.6000 663.3000 55.8000 676.2000 ;
	    RECT 57.0000 663.3000 58.2000 675.3000 ;
	    RECT 59.4000 663.3000 60.6000 676.2000 ;
	    RECT 61.8000 663.3000 63.0000 675.3000 ;
	    RECT 64.2000 663.3000 65.4000 676.2000 ;
	    RECT 66.6000 663.3000 67.8000 675.3000 ;
	    RECT 69.0000 663.3000 70.2000 676.2000 ;
	    RECT 88.2000 675.4500 89.4000 675.6000 ;
	    RECT 95.4000 675.4500 96.6000 675.6000 ;
	    RECT 71.4000 663.3000 72.6000 675.3000 ;
	    RECT 88.2000 674.5500 96.6000 675.4500 ;
	    RECT 88.2000 674.4000 89.4000 674.5500 ;
	    RECT 95.4000 674.4000 96.6000 674.5500 ;
	    RECT 98.4000 675.3000 99.3000 680.4000 ;
	    RECT 100.2000 679.5000 101.4000 679.8000 ;
	    RECT 100.2000 678.4500 101.4000 678.6000 ;
	    RECT 105.1500 678.4500 106.0500 680.5500 ;
	    RECT 117.0000 680.4000 118.2000 680.5500 ;
	    RECT 129.0000 681.4500 130.2000 681.6000 ;
	    RECT 150.6000 681.4500 151.8000 681.6000 ;
	    RECT 129.0000 680.5500 151.8000 681.4500 ;
	    RECT 152.7000 680.7000 153.0000 682.2000 ;
	    RECT 158.1000 681.6000 159.0000 683.7000 ;
	    RECT 162.6000 683.5500 175.8000 684.4500 ;
	    RECT 162.6000 683.4000 163.8000 683.5500 ;
	    RECT 174.6000 683.4000 175.8000 683.5500 ;
	    RECT 177.0000 682.5000 178.2000 689.7000 ;
	    RECT 215.4000 688.8000 221.4000 689.7000 ;
	    RECT 189.0000 687.4500 190.2000 687.6000 ;
	    RECT 213.0000 687.4500 214.2000 687.6000 ;
	    RECT 189.0000 686.5500 214.2000 687.4500 ;
	    RECT 189.0000 686.4000 190.2000 686.5500 ;
	    RECT 213.0000 686.4000 214.2000 686.5500 ;
	    RECT 179.4000 684.4500 180.6000 684.6000 ;
	    RECT 213.0000 684.4500 214.2000 684.6000 ;
	    RECT 179.4000 683.5500 214.2000 684.4500 ;
	    RECT 215.4000 683.7000 216.6000 688.8000 ;
	    RECT 217.8000 683.7000 219.0000 687.9000 ;
	    RECT 220.2000 684.0000 221.4000 688.8000 ;
	    RECT 222.6000 684.9000 223.8000 689.7000 ;
	    RECT 225.0000 684.0000 226.2000 689.7000 ;
	    RECT 220.2000 683.7000 226.2000 684.0000 ;
	    RECT 249.0000 684.0000 250.2000 689.7000 ;
	    RECT 251.4000 684.9000 252.6000 689.7000 ;
	    RECT 253.8000 684.0000 255.0000 689.7000 ;
	    RECT 249.0000 683.7000 255.0000 684.0000 ;
	    RECT 256.2000 683.7000 257.4000 689.7000 ;
	    RECT 275.4000 683.7000 276.6000 689.7000 ;
	    RECT 279.3000 684.6000 280.5000 689.7000 ;
	    RECT 405.0000 686.7000 406.2000 689.7000 ;
	    RECT 277.8000 683.7000 280.5000 684.6000 ;
	    RECT 407.4000 684.0000 408.6000 689.7000 ;
	    RECT 179.4000 683.4000 180.6000 683.5500 ;
	    RECT 213.0000 683.4000 214.2000 683.5500 ;
	    RECT 217.8000 681.6000 218.7000 683.7000 ;
	    RECT 220.5000 683.1000 225.9000 683.7000 ;
	    RECT 249.3000 683.1000 254.7000 683.7000 ;
	    RECT 256.2000 682.5000 257.1000 683.7000 ;
	    RECT 275.4000 682.5000 276.6000 682.8000 ;
	    RECT 129.0000 680.4000 130.2000 680.5500 ;
	    RECT 150.6000 680.4000 151.8000 680.5500 ;
	    RECT 155.4000 680.4000 156.6000 681.6000 ;
	    RECT 157.5000 680.7000 159.0000 681.6000 ;
	    RECT 160.2000 681.4500 161.4000 681.6000 ;
	    RECT 174.6000 681.4500 175.8000 681.6000 ;
	    RECT 160.2000 680.5500 175.8000 681.4500 ;
	    RECT 160.2000 680.4000 161.4000 680.5500 ;
	    RECT 174.6000 680.4000 175.8000 680.5500 ;
	    RECT 177.0000 681.4500 178.2000 681.6000 ;
	    RECT 215.4000 681.4500 216.6000 681.6000 ;
	    RECT 177.0000 680.5500 216.6000 681.4500 ;
	    RECT 217.8000 680.7000 219.3000 681.6000 ;
	    RECT 177.0000 680.4000 178.2000 680.5500 ;
	    RECT 215.4000 680.4000 216.6000 680.5500 ;
	    RECT 220.2000 680.4000 221.4000 681.6000 ;
	    RECT 223.8000 680.7000 224.1000 682.2000 ;
	    RECT 225.0000 681.4500 226.2000 681.6000 ;
	    RECT 227.4000 681.4500 228.6000 681.6000 ;
	    RECT 225.0000 680.5500 228.6000 681.4500 ;
	    RECT 225.0000 680.4000 226.2000 680.5500 ;
	    RECT 227.4000 680.4000 228.6000 680.5500 ;
	    RECT 249.0000 680.4000 250.2000 681.6000 ;
	    RECT 251.1000 680.7000 251.4000 682.2000 ;
	    RECT 253.5000 680.4000 255.3000 681.6000 ;
	    RECT 256.2000 681.4500 257.4000 681.6000 ;
	    RECT 261.0000 681.4500 262.2000 681.6000 ;
	    RECT 256.2000 680.5500 262.2000 681.4500 ;
	    RECT 256.2000 680.4000 257.4000 680.5500 ;
	    RECT 261.0000 680.4000 262.2000 680.5500 ;
	    RECT 275.4000 680.4000 276.6000 681.6000 ;
	    RECT 153.0000 679.5000 154.2000 679.8000 ;
	    RECT 157.8000 679.5000 159.0000 679.8000 ;
	    RECT 217.8000 679.5000 219.0000 679.8000 ;
	    RECT 222.6000 679.5000 223.8000 679.8000 ;
	    RECT 251.4000 679.5000 252.6000 679.8000 ;
	    RECT 100.2000 677.5500 106.0500 678.4500 ;
	    RECT 100.2000 677.4000 101.4000 677.5500 ;
	    RECT 98.4000 674.4000 99.9000 675.3000 ;
	    RECT 96.6000 672.6000 97.5000 673.5000 ;
	    RECT 96.6000 671.4000 97.8000 672.6000 ;
	    RECT 96.3000 663.3000 97.5000 669.3000 ;
	    RECT 98.7000 663.3000 99.9000 674.4000 ;
	    RECT 102.6000 663.3000 103.8000 675.3000 ;
	    RECT 117.0000 663.3000 118.2000 679.5000 ;
	    RECT 153.0000 677.4000 154.2000 678.6000 ;
	    RECT 155.4000 675.3000 156.3000 679.5000 ;
	    RECT 160.2000 679.2000 161.4000 679.5000 ;
	    RECT 157.8000 677.4000 159.0000 678.6000 ;
	    RECT 119.4000 663.3000 120.6000 669.3000 ;
	    RECT 150.6000 663.3000 151.8000 675.3000 ;
	    RECT 154.5000 663.3000 157.5000 675.3000 ;
	    RECT 160.2000 663.3000 161.4000 675.3000 ;
	    RECT 174.6000 663.3000 175.8000 669.3000 ;
	    RECT 177.0000 663.3000 178.2000 679.5000 ;
	    RECT 215.4000 679.2000 216.6000 679.5000 ;
	    RECT 217.8000 677.4000 219.0000 678.6000 ;
	    RECT 220.5000 675.3000 221.4000 679.5000 ;
	    RECT 222.6000 678.4500 223.8000 678.6000 ;
	    RECT 239.4000 678.4500 240.6000 678.6000 ;
	    RECT 222.6000 677.5500 240.6000 678.4500 ;
	    RECT 222.6000 677.4000 223.8000 677.5500 ;
	    RECT 239.4000 677.4000 240.6000 677.5500 ;
	    RECT 244.2000 678.4500 245.4000 678.6000 ;
	    RECT 251.4000 678.4500 252.6000 678.6000 ;
	    RECT 244.2000 677.5500 252.6000 678.4500 ;
	    RECT 244.2000 677.4000 245.4000 677.5500 ;
	    RECT 251.4000 677.4000 252.6000 677.5500 ;
	    RECT 253.5000 675.3000 254.4000 680.4000 ;
	    RECT 277.8000 679.5000 279.0000 683.7000 ;
	    RECT 407.1000 682.8000 408.6000 684.0000 ;
	    RECT 277.8000 677.4000 279.0000 678.6000 ;
	    RECT 215.4000 663.3000 216.6000 675.3000 ;
	    RECT 219.3000 663.3000 222.3000 675.3000 ;
	    RECT 225.0000 663.3000 226.2000 675.3000 ;
	    RECT 249.0000 663.3000 250.2000 675.3000 ;
	    RECT 252.9000 674.4000 254.4000 675.3000 ;
	    RECT 256.2000 674.4000 257.4000 675.6000 ;
	    RECT 252.9000 663.3000 254.1000 674.4000 ;
	    RECT 255.3000 672.6000 256.2000 673.5000 ;
	    RECT 255.0000 671.4000 256.2000 672.6000 ;
	    RECT 255.3000 663.3000 256.5000 669.3000 ;
	    RECT 275.4000 663.3000 276.6000 669.3000 ;
	    RECT 277.8000 663.3000 279.0000 676.5000 ;
	    RECT 407.1000 676.2000 408.3000 682.8000 ;
	    RECT 409.8000 681.9000 411.0000 689.7000 ;
	    RECT 414.6000 683.7000 415.8000 689.7000 ;
	    RECT 419.4000 684.9000 420.6000 689.7000 ;
	    RECT 421.8000 685.5000 423.0000 689.7000 ;
	    RECT 424.2000 685.5000 425.4000 689.7000 ;
	    RECT 426.6000 685.5000 427.8000 689.7000 ;
	    RECT 429.0000 685.5000 430.2000 689.7000 ;
	    RECT 431.4000 686.7000 432.6000 689.7000 ;
	    RECT 433.8000 685.5000 435.0000 689.7000 ;
	    RECT 436.2000 686.7000 437.4000 689.7000 ;
	    RECT 438.6000 685.5000 439.8000 689.7000 ;
	    RECT 441.0000 685.5000 442.2000 689.7000 ;
	    RECT 443.4000 685.5000 444.6000 689.7000 ;
	    RECT 417.0000 683.7000 420.6000 684.9000 ;
	    RECT 445.8000 684.9000 447.0000 689.7000 ;
	    RECT 417.0000 682.8000 418.2000 683.7000 ;
	    RECT 409.2000 681.0000 411.0000 681.9000 ;
	    RECT 415.5000 681.9000 418.2000 682.8000 ;
	    RECT 424.2000 683.4000 425.7000 684.6000 ;
	    RECT 430.2000 683.4000 430.5000 684.6000 ;
	    RECT 431.4000 683.4000 432.6000 684.6000 ;
	    RECT 433.8000 683.7000 440.7000 684.6000 ;
	    RECT 445.8000 683.7000 449.7000 684.9000 ;
	    RECT 450.6000 683.7000 451.8000 689.7000 ;
	    RECT 433.8000 683.4000 435.0000 683.7000 ;
	    RECT 409.2000 678.0000 410.1000 681.0000 ;
	    RECT 415.5000 680.1000 416.7000 681.9000 ;
	    RECT 411.0000 678.9000 416.7000 680.1000 ;
	    RECT 424.2000 679.2000 425.4000 683.4000 ;
	    RECT 436.2000 682.5000 437.4000 682.8000 ;
	    RECT 433.8000 682.2000 435.0000 682.5000 ;
	    RECT 428.4000 681.3000 435.0000 682.2000 ;
	    RECT 428.4000 681.0000 429.6000 681.3000 ;
	    RECT 436.2000 680.4000 437.4000 681.6000 ;
	    RECT 439.5000 680.1000 440.7000 683.7000 ;
	    RECT 448.5000 682.8000 449.7000 683.7000 ;
	    RECT 448.5000 681.6000 453.0000 682.8000 ;
	    RECT 455.4000 680.7000 456.6000 689.7000 ;
	    RECT 429.0000 678.9000 433.8000 680.1000 ;
	    RECT 439.5000 678.9000 442.5000 680.1000 ;
	    RECT 443.4000 679.5000 456.6000 680.7000 ;
	    RECT 419.4000 678.0000 420.6000 678.9000 ;
	    RECT 409.2000 677.1000 410.4000 678.0000 ;
	    RECT 419.4000 677.1000 444.9000 678.0000 ;
	    RECT 445.8000 677.4000 447.0000 678.6000 ;
	    RECT 453.3000 678.0000 454.5000 678.3000 ;
	    RECT 447.9000 677.1000 454.5000 678.0000 ;
	    RECT 280.2000 675.4500 281.4000 675.6000 ;
	    RECT 364.2000 675.4500 365.4000 675.6000 ;
	    RECT 280.2000 674.5500 365.4000 675.4500 ;
	    RECT 407.1000 675.0000 408.6000 676.2000 ;
	    RECT 280.2000 674.4000 281.4000 674.5500 ;
	    RECT 364.2000 674.4000 365.4000 674.5500 ;
	    RECT 407.4000 673.5000 408.6000 675.0000 ;
	    RECT 409.5000 674.4000 410.4000 677.1000 ;
	    RECT 411.3000 676.2000 412.5000 676.5000 ;
	    RECT 411.3000 675.3000 449.7000 676.2000 ;
	    RECT 445.5000 675.0000 446.7000 675.3000 ;
	    RECT 450.6000 674.4000 451.8000 675.6000 ;
	    RECT 409.5000 673.5000 423.0000 674.4000 ;
	    RECT 280.2000 673.2000 281.4000 673.5000 ;
	    RECT 340.2000 672.4500 341.4000 672.6000 ;
	    RECT 381.0000 672.4500 382.2000 672.6000 ;
	    RECT 407.4000 672.4500 408.6000 672.6000 ;
	    RECT 340.2000 671.5500 408.6000 672.4500 ;
	    RECT 340.2000 671.4000 341.4000 671.5500 ;
	    RECT 381.0000 671.4000 382.2000 671.5500 ;
	    RECT 407.4000 671.4000 408.6000 671.5500 ;
	    RECT 409.5000 671.1000 410.4000 673.5000 ;
	    RECT 421.8000 673.2000 423.0000 673.5000 ;
	    RECT 426.6000 673.5000 439.5000 674.4000 ;
	    RECT 426.6000 673.2000 427.8000 673.5000 ;
	    RECT 414.3000 671.4000 418.2000 672.6000 ;
	    RECT 280.2000 663.3000 281.4000 669.3000 ;
	    RECT 405.0000 663.3000 406.2000 669.3000 ;
	    RECT 407.4000 663.3000 408.6000 670.5000 ;
	    RECT 409.5000 670.2000 413.4000 671.1000 ;
	    RECT 409.8000 663.3000 411.0000 669.3000 ;
	    RECT 412.2000 663.3000 413.4000 670.2000 ;
	    RECT 414.6000 663.3000 415.8000 669.3000 ;
	    RECT 417.0000 663.3000 418.2000 671.4000 ;
	    RECT 419.1000 670.2000 425.4000 671.4000 ;
	    RECT 419.4000 663.3000 420.6000 669.3000 ;
	    RECT 421.8000 663.3000 423.0000 667.5000 ;
	    RECT 424.2000 663.3000 425.4000 667.5000 ;
	    RECT 426.6000 663.3000 427.8000 667.5000 ;
	    RECT 429.0000 663.3000 430.2000 672.6000 ;
	    RECT 433.8000 671.4000 437.7000 672.6000 ;
	    RECT 438.6000 672.3000 439.5000 673.5000 ;
	    RECT 441.0000 674.1000 442.2000 674.4000 ;
	    RECT 441.0000 673.5000 449.1000 674.1000 ;
	    RECT 441.0000 673.2000 450.3000 673.5000 ;
	    RECT 448.2000 672.3000 450.3000 673.2000 ;
	    RECT 438.6000 671.4000 447.3000 672.3000 ;
	    RECT 451.8000 672.0000 454.2000 673.2000 ;
	    RECT 451.8000 671.4000 452.7000 672.0000 ;
	    RECT 431.4000 663.3000 432.6000 669.3000 ;
	    RECT 433.8000 663.3000 435.0000 670.5000 ;
	    RECT 436.2000 663.3000 437.4000 669.3000 ;
	    RECT 438.6000 663.3000 439.8000 670.5000 ;
	    RECT 446.4000 670.2000 452.7000 671.4000 ;
	    RECT 455.4000 671.1000 456.6000 679.5000 ;
	    RECT 587.4000 680.7000 588.6000 689.7000 ;
	    RECT 592.2000 683.7000 593.4000 689.7000 ;
	    RECT 597.0000 684.9000 598.2000 689.7000 ;
	    RECT 599.4000 685.5000 600.6000 689.7000 ;
	    RECT 601.8000 685.5000 603.0000 689.7000 ;
	    RECT 604.2000 685.5000 605.4000 689.7000 ;
	    RECT 606.6000 686.7000 607.8000 689.7000 ;
	    RECT 609.0000 685.5000 610.2000 689.7000 ;
	    RECT 611.4000 686.7000 612.6000 689.7000 ;
	    RECT 613.8000 685.5000 615.0000 689.7000 ;
	    RECT 616.2000 685.5000 617.4000 689.7000 ;
	    RECT 618.6000 685.5000 619.8000 689.7000 ;
	    RECT 621.0000 685.5000 622.2000 689.7000 ;
	    RECT 594.3000 683.7000 598.2000 684.9000 ;
	    RECT 623.4000 684.9000 624.6000 689.7000 ;
	    RECT 603.3000 683.7000 610.2000 684.6000 ;
	    RECT 594.3000 682.8000 595.5000 683.7000 ;
	    RECT 591.0000 681.6000 595.5000 682.8000 ;
	    RECT 587.4000 679.5000 600.6000 680.7000 ;
	    RECT 603.3000 680.1000 604.5000 683.7000 ;
	    RECT 609.0000 683.4000 610.2000 683.7000 ;
	    RECT 611.4000 683.4000 612.6000 684.6000 ;
	    RECT 613.5000 683.4000 613.8000 684.6000 ;
	    RECT 618.3000 683.4000 619.8000 684.6000 ;
	    RECT 623.4000 683.7000 627.0000 684.9000 ;
	    RECT 628.2000 683.7000 629.4000 689.7000 ;
	    RECT 606.6000 682.5000 607.8000 682.8000 ;
	    RECT 609.0000 682.2000 610.2000 682.5000 ;
	    RECT 606.6000 680.4000 607.8000 681.6000 ;
	    RECT 609.0000 681.3000 615.6000 682.2000 ;
	    RECT 614.4000 681.0000 615.6000 681.3000 ;
	    RECT 508.2000 678.4500 509.4000 678.6000 ;
	    RECT 582.6000 678.4500 583.8000 678.6000 ;
	    RECT 508.2000 677.5500 583.8000 678.4500 ;
	    RECT 508.2000 677.4000 509.4000 677.5500 ;
	    RECT 582.6000 677.4000 583.8000 677.5500 ;
	    RECT 453.6000 670.2000 456.6000 671.1000 ;
	    RECT 587.4000 671.1000 588.6000 679.5000 ;
	    RECT 601.5000 678.9000 604.5000 680.1000 ;
	    RECT 610.2000 678.9000 615.0000 680.1000 ;
	    RECT 618.6000 679.2000 619.8000 683.4000 ;
	    RECT 625.8000 682.8000 627.0000 683.7000 ;
	    RECT 625.8000 681.9000 628.5000 682.8000 ;
	    RECT 627.3000 680.1000 628.5000 681.9000 ;
	    RECT 633.0000 681.9000 634.2000 689.7000 ;
	    RECT 635.4000 684.0000 636.6000 689.7000 ;
	    RECT 637.8000 686.7000 639.0000 689.7000 ;
	    RECT 635.4000 682.8000 636.9000 684.0000 ;
	    RECT 669.0000 683.7000 670.2000 689.7000 ;
	    RECT 671.4000 684.0000 672.6000 689.7000 ;
	    RECT 673.8000 684.9000 675.0000 689.7000 ;
	    RECT 676.2000 684.0000 677.4000 689.7000 ;
	    RECT 671.4000 683.7000 677.4000 684.0000 ;
	    RECT 633.0000 681.0000 634.8000 681.9000 ;
	    RECT 627.3000 678.9000 633.0000 680.1000 ;
	    RECT 589.5000 678.0000 590.7000 678.3000 ;
	    RECT 589.5000 677.1000 596.1000 678.0000 ;
	    RECT 597.0000 677.4000 598.2000 678.6000 ;
	    RECT 623.4000 678.0000 624.6000 678.9000 ;
	    RECT 633.9000 678.0000 634.8000 681.0000 ;
	    RECT 599.1000 677.1000 624.6000 678.0000 ;
	    RECT 633.6000 677.1000 634.8000 678.0000 ;
	    RECT 631.5000 676.2000 632.7000 676.5000 ;
	    RECT 589.8000 675.4500 591.0000 675.6000 ;
	    RECT 592.2000 675.4500 593.4000 675.6000 ;
	    RECT 589.8000 674.5500 593.4000 675.4500 ;
	    RECT 594.3000 675.3000 632.7000 676.2000 ;
	    RECT 597.3000 675.0000 598.5000 675.3000 ;
	    RECT 589.8000 674.4000 591.0000 674.5500 ;
	    RECT 592.2000 674.4000 593.4000 674.5500 ;
	    RECT 633.6000 674.4000 634.5000 677.1000 ;
	    RECT 635.7000 676.2000 636.9000 682.8000 ;
	    RECT 669.3000 682.5000 670.2000 683.7000 ;
	    RECT 671.7000 683.1000 677.1000 683.7000 ;
	    RECT 690.6000 682.5000 691.8000 689.7000 ;
	    RECT 693.0000 686.7000 694.2000 689.7000 ;
	    RECT 693.0000 685.5000 694.2000 685.8000 ;
	    RECT 693.0000 684.4500 694.2000 684.6000 ;
	    RECT 707.4000 684.4500 708.6000 684.6000 ;
	    RECT 693.0000 683.5500 708.6000 684.4500 ;
	    RECT 712.2000 683.7000 713.4000 689.7000 ;
	    RECT 716.1000 684.6000 717.3000 689.7000 ;
	    RECT 731.4000 686.7000 732.6000 689.7000 ;
	    RECT 731.4000 685.5000 732.6000 685.8000 ;
	    RECT 714.6000 683.7000 717.3000 684.6000 ;
	    RECT 693.0000 683.4000 694.2000 683.5500 ;
	    RECT 707.4000 683.4000 708.6000 683.5500 ;
	    RECT 712.2000 682.5000 713.4000 682.8000 ;
	    RECT 637.8000 681.4500 639.0000 681.6000 ;
	    RECT 669.0000 681.4500 670.2000 681.6000 ;
	    RECT 637.8000 680.5500 670.2000 681.4500 ;
	    RECT 637.8000 680.4000 639.0000 680.5500 ;
	    RECT 669.0000 680.4000 670.2000 680.5500 ;
	    RECT 671.1000 680.4000 672.9000 681.6000 ;
	    RECT 675.0000 680.7000 675.3000 682.2000 ;
	    RECT 676.2000 680.4000 677.4000 681.6000 ;
	    RECT 690.6000 681.4500 691.8000 681.6000 ;
	    RECT 678.7500 680.5500 691.8000 681.4500 ;
	    RECT 601.8000 674.1000 603.0000 674.4000 ;
	    RECT 594.9000 673.5000 603.0000 674.1000 ;
	    RECT 593.7000 673.2000 603.0000 673.5000 ;
	    RECT 604.5000 673.5000 617.4000 674.4000 ;
	    RECT 589.8000 672.0000 592.2000 673.2000 ;
	    RECT 593.7000 672.3000 595.8000 673.2000 ;
	    RECT 604.5000 672.3000 605.4000 673.5000 ;
	    RECT 616.2000 673.2000 617.4000 673.5000 ;
	    RECT 621.0000 673.5000 634.5000 674.4000 ;
	    RECT 635.4000 675.0000 636.9000 676.2000 ;
	    RECT 642.6000 675.4500 643.8000 675.6000 ;
	    RECT 669.0000 675.4500 670.2000 675.6000 ;
	    RECT 635.4000 673.5000 636.6000 675.0000 ;
	    RECT 642.6000 674.5500 670.2000 675.4500 ;
	    RECT 642.6000 674.4000 643.8000 674.5500 ;
	    RECT 669.0000 674.4000 670.2000 674.5500 ;
	    RECT 672.0000 675.3000 672.9000 680.4000 ;
	    RECT 673.8000 679.5000 675.0000 679.8000 ;
	    RECT 673.8000 678.4500 675.0000 678.6000 ;
	    RECT 678.7500 678.4500 679.6500 680.5500 ;
	    RECT 690.6000 680.4000 691.8000 680.5500 ;
	    RECT 695.4000 681.4500 696.6000 681.6000 ;
	    RECT 712.2000 681.4500 713.4000 681.6000 ;
	    RECT 695.4000 680.5500 713.4000 681.4500 ;
	    RECT 695.4000 680.4000 696.6000 680.5500 ;
	    RECT 712.2000 680.4000 713.4000 680.5500 ;
	    RECT 714.6000 679.5000 715.8000 683.7000 ;
	    RECT 731.4000 683.4000 732.6000 684.6000 ;
	    RECT 733.8000 682.5000 735.0000 689.7000 ;
	    RECT 762.6000 684.0000 763.8000 689.7000 ;
	    RECT 765.0000 684.9000 766.2000 689.7000 ;
	    RECT 767.4000 688.8000 773.4000 689.7000 ;
	    RECT 767.4000 684.0000 768.6000 688.8000 ;
	    RECT 762.6000 683.7000 768.6000 684.0000 ;
	    RECT 769.8000 683.7000 771.0000 687.9000 ;
	    RECT 772.2000 683.7000 773.4000 688.8000 ;
	    RECT 791.4000 686.7000 792.6000 689.7000 ;
	    RECT 793.8000 686.7000 795.0000 689.7000 ;
	    RECT 796.2000 686.7000 797.4000 689.7000 ;
	    RECT 810.6000 686.7000 811.8000 689.7000 ;
	    RECT 791.4000 685.5000 792.6000 685.8000 ;
	    RECT 781.8000 684.4500 783.0000 684.6000 ;
	    RECT 791.4000 684.4500 792.6000 684.6000 ;
	    RECT 762.9000 683.1000 768.3000 683.7000 ;
	    RECT 733.8000 681.4500 735.0000 681.6000 ;
	    RECT 762.6000 681.4500 763.8000 681.6000 ;
	    RECT 733.8000 680.5500 763.8000 681.4500 ;
	    RECT 764.7000 680.7000 765.0000 682.2000 ;
	    RECT 770.1000 681.6000 771.0000 683.7000 ;
	    RECT 781.8000 683.5500 792.6000 684.4500 ;
	    RECT 781.8000 683.4000 783.0000 683.5500 ;
	    RECT 791.4000 683.4000 792.6000 683.5500 ;
	    RECT 794.1000 682.5000 795.0000 686.7000 ;
	    RECT 810.6000 685.5000 811.8000 685.8000 ;
	    RECT 810.6000 683.4000 811.8000 684.6000 ;
	    RECT 813.0000 682.5000 814.2000 689.7000 ;
	    RECT 833.1000 684.6000 834.3000 689.7000 ;
	    RECT 833.1000 683.7000 835.8000 684.6000 ;
	    RECT 837.0000 683.7000 838.2000 689.7000 ;
	    RECT 858.6000 684.4500 859.8000 684.6000 ;
	    RECT 733.8000 680.4000 735.0000 680.5500 ;
	    RECT 762.6000 680.4000 763.8000 680.5500 ;
	    RECT 767.4000 680.4000 768.6000 681.6000 ;
	    RECT 769.5000 680.7000 771.0000 681.6000 ;
	    RECT 772.2000 680.4000 773.4000 681.6000 ;
	    RECT 789.0000 681.4500 790.2000 681.6000 ;
	    RECT 793.8000 681.4500 795.0000 681.6000 ;
	    RECT 789.0000 680.5500 795.0000 681.4500 ;
	    RECT 789.0000 680.4000 790.2000 680.5500 ;
	    RECT 793.8000 680.4000 795.0000 680.5500 ;
	    RECT 813.0000 681.4500 814.2000 681.6000 ;
	    RECT 822.6000 681.4500 823.8000 681.6000 ;
	    RECT 813.0000 680.5500 823.8000 681.4500 ;
	    RECT 813.0000 680.4000 814.2000 680.5500 ;
	    RECT 822.6000 680.4000 823.8000 680.5500 ;
	    RECT 765.0000 679.5000 766.2000 679.8000 ;
	    RECT 769.8000 679.5000 771.0000 679.8000 ;
	    RECT 834.6000 679.5000 835.8000 683.7000 ;
	    RECT 849.1500 683.5500 859.8000 684.4500 ;
	    RECT 865.8000 684.0000 867.0000 689.7000 ;
	    RECT 868.2000 684.9000 869.4000 689.7000 ;
	    RECT 870.6000 688.8000 876.6000 689.7000 ;
	    RECT 870.6000 684.0000 871.8000 688.8000 ;
	    RECT 865.8000 683.7000 871.8000 684.0000 ;
	    RECT 873.0000 683.7000 874.2000 687.9000 ;
	    RECT 875.4000 683.7000 876.6000 688.8000 ;
	    RECT 837.0000 682.5000 838.2000 682.8000 ;
	    RECT 837.0000 681.4500 838.2000 681.6000 ;
	    RECT 849.1500 681.4500 850.0500 683.5500 ;
	    RECT 858.6000 683.4000 859.8000 683.5500 ;
	    RECT 866.1000 683.1000 871.5000 683.7000 ;
	    RECT 837.0000 680.5500 850.0500 681.4500 ;
	    RECT 851.4000 681.4500 852.6000 681.6000 ;
	    RECT 865.8000 681.4500 867.0000 681.6000 ;
	    RECT 851.4000 680.5500 867.0000 681.4500 ;
	    RECT 867.9000 680.7000 868.2000 682.2000 ;
	    RECT 873.3000 681.6000 874.2000 683.7000 ;
	    RECT 889.8000 682.5000 891.0000 689.7000 ;
	    RECT 892.2000 686.7000 893.4000 689.7000 ;
	    RECT 913.8000 686.7000 915.0000 689.7000 ;
	    RECT 892.2000 685.5000 893.4000 685.8000 ;
	    RECT 913.8000 685.5000 915.0000 685.8000 ;
	    RECT 892.2000 684.4500 893.4000 684.6000 ;
	    RECT 904.2000 684.4500 905.4000 684.6000 ;
	    RECT 892.2000 683.5500 905.4000 684.4500 ;
	    RECT 892.2000 683.4000 893.4000 683.5500 ;
	    RECT 904.2000 683.4000 905.4000 683.5500 ;
	    RECT 913.8000 683.4000 915.0000 684.6000 ;
	    RECT 916.2000 682.5000 917.4000 689.7000 ;
	    RECT 945.0000 684.0000 946.2000 689.7000 ;
	    RECT 947.4000 684.9000 948.6000 689.7000 ;
	    RECT 949.8000 688.8000 955.8000 689.7000 ;
	    RECT 949.8000 684.0000 951.0000 688.8000 ;
	    RECT 945.0000 683.7000 951.0000 684.0000 ;
	    RECT 952.2000 683.7000 953.4000 687.9000 ;
	    RECT 954.6000 683.7000 955.8000 688.8000 ;
	    RECT 1079.4000 686.7000 1080.6000 689.7000 ;
	    RECT 1081.8000 684.0000 1083.0000 689.7000 ;
	    RECT 945.3000 683.1000 950.7000 683.7000 ;
	    RECT 837.0000 680.4000 838.2000 680.5500 ;
	    RECT 851.4000 680.4000 852.6000 680.5500 ;
	    RECT 865.8000 680.4000 867.0000 680.5500 ;
	    RECT 870.6000 680.4000 871.8000 681.6000 ;
	    RECT 872.7000 680.7000 874.2000 681.6000 ;
	    RECT 875.4000 681.4500 876.6000 681.6000 ;
	    RECT 889.8000 681.4500 891.0000 681.6000 ;
	    RECT 875.4000 680.5500 891.0000 681.4500 ;
	    RECT 875.4000 680.4000 876.6000 680.5500 ;
	    RECT 889.8000 680.4000 891.0000 680.5500 ;
	    RECT 916.2000 681.4500 917.4000 681.6000 ;
	    RECT 921.0000 681.4500 922.2000 681.6000 ;
	    RECT 916.2000 680.5500 922.2000 681.4500 ;
	    RECT 916.2000 680.4000 917.4000 680.5500 ;
	    RECT 921.0000 680.4000 922.2000 680.5500 ;
	    RECT 933.0000 681.4500 934.2000 681.6000 ;
	    RECT 945.0000 681.4500 946.2000 681.6000 ;
	    RECT 933.0000 680.5500 946.2000 681.4500 ;
	    RECT 947.1000 680.7000 947.4000 682.2000 ;
	    RECT 952.5000 681.6000 953.4000 683.7000 ;
	    RECT 1081.5000 682.8000 1083.0000 684.0000 ;
	    RECT 933.0000 680.4000 934.2000 680.5500 ;
	    RECT 945.0000 680.4000 946.2000 680.5500 ;
	    RECT 949.8000 680.4000 951.0000 681.6000 ;
	    RECT 951.9000 680.7000 953.4000 681.6000 ;
	    RECT 954.6000 681.4500 955.8000 681.6000 ;
	    RECT 1009.8000 681.4500 1011.0000 681.6000 ;
	    RECT 954.6000 680.5500 1011.0000 681.4500 ;
	    RECT 954.6000 680.4000 955.8000 680.5500 ;
	    RECT 1009.8000 680.4000 1011.0000 680.5500 ;
	    RECT 868.2000 679.5000 869.4000 679.8000 ;
	    RECT 873.0000 679.5000 874.2000 679.8000 ;
	    RECT 947.4000 679.5000 948.6000 679.8000 ;
	    RECT 952.2000 679.5000 953.4000 679.8000 ;
	    RECT 673.8000 677.5500 679.6500 678.4500 ;
	    RECT 673.8000 677.4000 675.0000 677.5500 ;
	    RECT 672.0000 674.4000 673.5000 675.3000 ;
	    RECT 621.0000 673.2000 622.2000 673.5000 ;
	    RECT 591.3000 671.4000 592.2000 672.0000 ;
	    RECT 596.7000 671.4000 605.4000 672.3000 ;
	    RECT 606.3000 671.4000 610.2000 672.6000 ;
	    RECT 587.4000 670.2000 590.4000 671.1000 ;
	    RECT 591.3000 670.2000 597.6000 671.4000 ;
	    RECT 441.0000 663.3000 442.2000 667.5000 ;
	    RECT 443.4000 663.3000 444.6000 667.5000 ;
	    RECT 445.8000 663.3000 447.0000 669.3000 ;
	    RECT 448.2000 663.3000 449.4000 670.2000 ;
	    RECT 453.6000 669.3000 454.5000 670.2000 ;
	    RECT 589.5000 669.3000 590.4000 670.2000 ;
	    RECT 450.6000 662.4000 451.8000 669.3000 ;
	    RECT 453.0000 668.4000 454.5000 669.3000 ;
	    RECT 453.0000 663.3000 454.2000 668.4000 ;
	    RECT 455.4000 663.3000 456.6000 669.3000 ;
	    RECT 587.4000 663.3000 588.6000 669.3000 ;
	    RECT 589.5000 668.4000 591.0000 669.3000 ;
	    RECT 589.8000 663.3000 591.0000 668.4000 ;
	    RECT 592.2000 662.4000 593.4000 669.3000 ;
	    RECT 594.6000 663.3000 595.8000 670.2000 ;
	    RECT 597.0000 663.3000 598.2000 669.3000 ;
	    RECT 599.4000 663.3000 600.6000 667.5000 ;
	    RECT 601.8000 663.3000 603.0000 667.5000 ;
	    RECT 604.2000 663.3000 605.4000 670.5000 ;
	    RECT 606.6000 663.3000 607.8000 669.3000 ;
	    RECT 609.0000 663.3000 610.2000 670.5000 ;
	    RECT 611.4000 663.3000 612.6000 669.3000 ;
	    RECT 613.8000 663.3000 615.0000 672.6000 ;
	    RECT 625.8000 671.4000 629.7000 672.6000 ;
	    RECT 618.6000 670.2000 624.9000 671.4000 ;
	    RECT 616.2000 663.3000 617.4000 667.5000 ;
	    RECT 618.6000 663.3000 619.8000 667.5000 ;
	    RECT 621.0000 663.3000 622.2000 667.5000 ;
	    RECT 623.4000 663.3000 624.6000 669.3000 ;
	    RECT 625.8000 663.3000 627.0000 671.4000 ;
	    RECT 633.6000 671.1000 634.5000 673.5000 ;
	    RECT 670.2000 672.6000 671.1000 673.5000 ;
	    RECT 635.4000 671.4000 636.6000 672.6000 ;
	    RECT 670.2000 671.4000 671.4000 672.6000 ;
	    RECT 630.6000 670.2000 634.5000 671.1000 ;
	    RECT 628.2000 663.3000 629.4000 669.3000 ;
	    RECT 630.6000 663.3000 631.8000 670.2000 ;
	    RECT 633.0000 663.3000 634.2000 669.3000 ;
	    RECT 635.4000 663.3000 636.6000 670.5000 ;
	    RECT 637.8000 663.3000 639.0000 669.3000 ;
	    RECT 669.9000 663.3000 671.1000 669.3000 ;
	    RECT 672.3000 663.3000 673.5000 674.4000 ;
	    RECT 676.2000 663.3000 677.4000 675.3000 ;
	    RECT 690.6000 663.3000 691.8000 679.5000 ;
	    RECT 693.0000 678.4500 694.2000 678.6000 ;
	    RECT 714.6000 678.4500 715.8000 678.6000 ;
	    RECT 693.0000 677.5500 715.8000 678.4500 ;
	    RECT 693.0000 677.4000 694.2000 677.5500 ;
	    RECT 714.6000 677.4000 715.8000 677.5500 ;
	    RECT 693.0000 663.3000 694.2000 669.3000 ;
	    RECT 712.2000 663.3000 713.4000 669.3000 ;
	    RECT 714.6000 663.3000 715.8000 676.5000 ;
	    RECT 717.0000 674.4000 718.2000 675.6000 ;
	    RECT 717.0000 673.2000 718.2000 673.5000 ;
	    RECT 717.0000 663.3000 718.2000 669.3000 ;
	    RECT 731.4000 663.3000 732.6000 669.3000 ;
	    RECT 733.8000 663.3000 735.0000 679.5000 ;
	    RECT 765.0000 677.4000 766.2000 678.6000 ;
	    RECT 767.4000 675.3000 768.3000 679.5000 ;
	    RECT 772.2000 679.2000 773.4000 679.5000 ;
	    RECT 769.8000 677.4000 771.0000 678.6000 ;
	    RECT 794.1000 675.3000 795.0000 679.5000 ;
	    RECT 796.2000 677.4000 797.4000 678.6000 ;
	    RECT 796.2000 676.2000 797.4000 676.5000 ;
	    RECT 762.6000 663.3000 763.8000 675.3000 ;
	    RECT 766.5000 663.3000 769.5000 675.3000 ;
	    RECT 772.2000 663.3000 773.4000 675.3000 ;
	    RECT 791.4000 663.3000 792.6000 675.3000 ;
	    RECT 793.8000 674.1000 796.5000 675.3000 ;
	    RECT 795.3000 663.3000 796.5000 674.1000 ;
	    RECT 810.6000 663.3000 811.8000 669.3000 ;
	    RECT 813.0000 663.3000 814.2000 679.5000 ;
	    RECT 825.0000 678.4500 826.2000 678.6000 ;
	    RECT 834.6000 678.4500 835.8000 678.6000 ;
	    RECT 825.0000 677.5500 835.8000 678.4500 ;
	    RECT 825.0000 677.4000 826.2000 677.5500 ;
	    RECT 834.6000 677.4000 835.8000 677.5500 ;
	    RECT 868.2000 677.4000 869.4000 678.6000 ;
	    RECT 832.2000 674.4000 833.4000 675.6000 ;
	    RECT 832.2000 673.2000 833.4000 673.5000 ;
	    RECT 832.2000 663.3000 833.4000 669.3000 ;
	    RECT 834.6000 663.3000 835.8000 676.5000 ;
	    RECT 870.6000 675.3000 871.5000 679.5000 ;
	    RECT 875.4000 679.2000 876.6000 679.5000 ;
	    RECT 873.0000 677.4000 874.2000 678.6000 ;
	    RECT 837.0000 663.3000 838.2000 669.3000 ;
	    RECT 865.8000 663.3000 867.0000 675.3000 ;
	    RECT 869.7000 663.3000 872.7000 675.3000 ;
	    RECT 875.4000 663.3000 876.6000 675.3000 ;
	    RECT 889.8000 663.3000 891.0000 679.5000 ;
	    RECT 892.2000 663.3000 893.4000 669.3000 ;
	    RECT 913.8000 663.3000 915.0000 669.3000 ;
	    RECT 916.2000 663.3000 917.4000 679.5000 ;
	    RECT 947.4000 677.4000 948.6000 678.6000 ;
	    RECT 949.8000 675.3000 950.7000 679.5000 ;
	    RECT 954.6000 679.2000 955.8000 679.5000 ;
	    RECT 952.2000 677.4000 953.4000 678.6000 ;
	    RECT 1081.5000 676.2000 1082.7001 682.8000 ;
	    RECT 1084.2001 681.9000 1085.4000 689.7000 ;
	    RECT 1089.0000 683.7000 1090.2001 689.7000 ;
	    RECT 1093.8000 684.9000 1095.0000 689.7000 ;
	    RECT 1096.2001 685.5000 1097.4000 689.7000 ;
	    RECT 1098.6000 685.5000 1099.8000 689.7000 ;
	    RECT 1101.0000 685.5000 1102.2001 689.7000 ;
	    RECT 1103.4000 685.5000 1104.6000 689.7000 ;
	    RECT 1105.8000 686.7000 1107.0000 689.7000 ;
	    RECT 1108.2001 685.5000 1109.4000 689.7000 ;
	    RECT 1110.6000 686.7000 1111.8000 689.7000 ;
	    RECT 1113.0000 685.5000 1114.2001 689.7000 ;
	    RECT 1115.4000 685.5000 1116.6000 689.7000 ;
	    RECT 1117.8000 685.5000 1119.0000 689.7000 ;
	    RECT 1091.4000 683.7000 1095.0000 684.9000 ;
	    RECT 1120.2001 684.9000 1121.4000 689.7000 ;
	    RECT 1091.4000 682.8000 1092.6000 683.7000 ;
	    RECT 1083.6000 681.0000 1085.4000 681.9000 ;
	    RECT 1089.9000 681.9000 1092.6000 682.8000 ;
	    RECT 1098.6000 683.4000 1100.1000 684.6000 ;
	    RECT 1104.6000 683.4000 1104.9000 684.6000 ;
	    RECT 1105.8000 683.4000 1107.0000 684.6000 ;
	    RECT 1108.2001 683.7000 1115.1000 684.6000 ;
	    RECT 1120.2001 683.7000 1124.1000 684.9000 ;
	    RECT 1125.0000 683.7000 1126.2001 689.7000 ;
	    RECT 1108.2001 683.4000 1109.4000 683.7000 ;
	    RECT 1083.6000 678.0000 1084.5000 681.0000 ;
	    RECT 1089.9000 680.1000 1091.1000 681.9000 ;
	    RECT 1085.4000 678.9000 1091.1000 680.1000 ;
	    RECT 1098.6000 679.2000 1099.8000 683.4000 ;
	    RECT 1110.6000 682.5000 1111.8000 682.8000 ;
	    RECT 1108.2001 682.2000 1109.4000 682.5000 ;
	    RECT 1102.8000 681.3000 1109.4000 682.2000 ;
	    RECT 1102.8000 681.0000 1104.0000 681.3000 ;
	    RECT 1110.6000 680.4000 1111.8000 681.6000 ;
	    RECT 1113.9000 680.1000 1115.1000 683.7000 ;
	    RECT 1122.9000 682.8000 1124.1000 683.7000 ;
	    RECT 1122.9000 681.6000 1127.4000 682.8000 ;
	    RECT 1129.8000 680.7000 1131.0000 689.7000 ;
	    RECT 1151.4000 686.7000 1152.6000 689.7000 ;
	    RECT 1151.4000 685.5000 1152.6000 685.8000 ;
	    RECT 1151.4000 683.4000 1152.6000 684.6000 ;
	    RECT 1153.8000 682.5000 1155.0000 689.7000 ;
	    RECT 1173.9000 684.6000 1175.1000 689.7000 ;
	    RECT 1173.9000 683.7000 1176.6000 684.6000 ;
	    RECT 1177.8000 683.7000 1179.0000 689.7000 ;
	    RECT 1192.2001 687.4500 1193.4000 687.6000 ;
	    RECT 1197.0000 687.4500 1198.2001 687.6000 ;
	    RECT 1192.2001 686.5500 1198.2001 687.4500 ;
	    RECT 1192.2001 686.4000 1193.4000 686.5500 ;
	    RECT 1197.0000 686.4000 1198.2001 686.5500 ;
	    RECT 1230.6000 683.7000 1231.8000 689.7000 ;
	    RECT 1103.4000 678.9000 1108.2001 680.1000 ;
	    RECT 1113.9000 678.9000 1116.9000 680.1000 ;
	    RECT 1117.8000 679.5000 1131.0000 680.7000 ;
	    RECT 1153.8000 681.4500 1155.0000 681.6000 ;
	    RECT 1161.0000 681.4500 1162.2001 681.6000 ;
	    RECT 1153.8000 680.5500 1162.2001 681.4500 ;
	    RECT 1153.8000 680.4000 1155.0000 680.5500 ;
	    RECT 1161.0000 680.4000 1162.2001 680.5500 ;
	    RECT 1175.4000 679.5000 1176.6000 683.7000 ;
	    RECT 1233.0000 682.8000 1234.2001 689.7000 ;
	    RECT 1235.4000 683.7000 1236.6000 689.7000 ;
	    RECT 1237.8000 682.8000 1239.0000 689.7000 ;
	    RECT 1240.2001 683.7000 1241.4000 689.7000 ;
	    RECT 1242.6000 682.8000 1243.8000 689.7000 ;
	    RECT 1245.0000 683.7000 1246.2001 689.7000 ;
	    RECT 1247.4000 682.8000 1248.6000 689.7000 ;
	    RECT 1249.8000 683.7000 1251.0000 689.7000 ;
	    RECT 1269.9000 684.6000 1271.1000 689.7000 ;
	    RECT 1269.9000 683.7000 1272.6000 684.6000 ;
	    RECT 1273.8000 683.7000 1275.0000 689.7000 ;
	    RECT 1293.9000 684.6000 1295.1000 689.7000 ;
	    RECT 1293.9000 683.7000 1296.6000 684.6000 ;
	    RECT 1297.8000 683.7000 1299.0000 689.7000 ;
	    RECT 1324.2001 684.0000 1325.4000 689.7000 ;
	    RECT 1326.6000 684.9000 1327.8000 689.7000 ;
	    RECT 1329.0000 684.0000 1330.2001 689.7000 ;
	    RECT 1324.2001 683.7000 1330.2001 684.0000 ;
	    RECT 1331.4000 683.7000 1332.6000 689.7000 ;
	    RECT 1350.6000 683.7000 1351.8000 689.7000 ;
	    RECT 1354.5000 684.6000 1355.7001 689.7000 ;
	    RECT 1353.0000 683.7000 1355.7001 684.6000 ;
	    RECT 1177.8000 682.5000 1179.0000 682.8000 ;
	    RECT 1233.0000 681.6000 1235.7001 682.8000 ;
	    RECT 1237.8000 681.6000 1241.1000 682.8000 ;
	    RECT 1242.6000 681.6000 1245.9000 682.8000 ;
	    RECT 1247.4000 681.6000 1251.0000 682.8000 ;
	    RECT 1177.8000 681.4500 1179.0000 681.6000 ;
	    RECT 1180.2001 681.4500 1181.4000 681.6000 ;
	    RECT 1177.8000 680.5500 1181.4000 681.4500 ;
	    RECT 1177.8000 680.4000 1179.0000 680.5500 ;
	    RECT 1180.2001 680.4000 1181.4000 680.5500 ;
	    RECT 1230.6000 680.4000 1231.8000 681.6000 ;
	    RECT 1234.5000 680.7000 1235.7001 681.6000 ;
	    RECT 1239.9000 680.7000 1241.1000 681.6000 ;
	    RECT 1244.7001 680.7000 1245.9000 681.6000 ;
	    RECT 1093.8000 678.0000 1095.0000 678.9000 ;
	    RECT 1083.6000 677.1000 1084.8000 678.0000 ;
	    RECT 1093.8000 677.1000 1119.3000 678.0000 ;
	    RECT 1120.2001 677.4000 1121.4000 678.6000 ;
	    RECT 1127.7001 678.0000 1128.9000 678.3000 ;
	    RECT 1122.3000 677.1000 1128.9000 678.0000 ;
	    RECT 945.0000 663.3000 946.2000 675.3000 ;
	    RECT 948.9000 663.3000 951.9000 675.3000 ;
	    RECT 954.6000 663.3000 955.8000 675.3000 ;
	    RECT 1081.5000 675.0000 1083.0000 676.2000 ;
	    RECT 1081.8000 673.5000 1083.0000 675.0000 ;
	    RECT 1083.9000 674.4000 1084.8000 677.1000 ;
	    RECT 1085.7001 676.2000 1086.9000 676.5000 ;
	    RECT 1085.7001 675.3000 1124.1000 676.2000 ;
	    RECT 1119.9000 675.0000 1121.1000 675.3000 ;
	    RECT 1125.0000 674.4000 1126.2001 675.6000 ;
	    RECT 1083.9000 673.5000 1097.4000 674.4000 ;
	    RECT 1000.2000 672.4500 1001.4000 672.6000 ;
	    RECT 1007.4000 672.4500 1008.6000 672.6000 ;
	    RECT 1081.8000 672.4500 1083.0000 672.6000 ;
	    RECT 1000.2000 671.5500 1083.0000 672.4500 ;
	    RECT 1000.2000 671.4000 1001.4000 671.5500 ;
	    RECT 1007.4000 671.4000 1008.6000 671.5500 ;
	    RECT 1081.8000 671.4000 1083.0000 671.5500 ;
	    RECT 1083.9000 671.1000 1084.8000 673.5000 ;
	    RECT 1096.2001 673.2000 1097.4000 673.5000 ;
	    RECT 1101.0000 673.5000 1113.9000 674.4000 ;
	    RECT 1101.0000 673.2000 1102.2001 673.5000 ;
	    RECT 1088.7001 671.4000 1092.6000 672.6000 ;
	    RECT 1079.4000 663.3000 1080.6000 669.3000 ;
	    RECT 1081.8000 663.3000 1083.0000 670.5000 ;
	    RECT 1083.9000 670.2000 1087.8000 671.1000 ;
	    RECT 1084.2001 663.3000 1085.4000 669.3000 ;
	    RECT 1086.6000 663.3000 1087.8000 670.2000 ;
	    RECT 1089.0000 663.3000 1090.2001 669.3000 ;
	    RECT 1091.4000 663.3000 1092.6000 671.4000 ;
	    RECT 1093.5000 670.2000 1099.8000 671.4000 ;
	    RECT 1093.8000 663.3000 1095.0000 669.3000 ;
	    RECT 1096.2001 663.3000 1097.4000 667.5000 ;
	    RECT 1098.6000 663.3000 1099.8000 667.5000 ;
	    RECT 1101.0000 663.3000 1102.2001 667.5000 ;
	    RECT 1103.4000 663.3000 1104.6000 672.6000 ;
	    RECT 1108.2001 671.4000 1112.1000 672.6000 ;
	    RECT 1113.0000 672.3000 1113.9000 673.5000 ;
	    RECT 1115.4000 674.1000 1116.6000 674.4000 ;
	    RECT 1115.4000 673.5000 1123.5000 674.1000 ;
	    RECT 1115.4000 673.2000 1124.7001 673.5000 ;
	    RECT 1122.6000 672.3000 1124.7001 673.2000 ;
	    RECT 1113.0000 671.4000 1121.7001 672.3000 ;
	    RECT 1126.2001 672.0000 1128.6000 673.2000 ;
	    RECT 1126.2001 671.4000 1127.1000 672.0000 ;
	    RECT 1105.8000 663.3000 1107.0000 669.3000 ;
	    RECT 1108.2001 663.3000 1109.4000 670.5000 ;
	    RECT 1110.6000 663.3000 1111.8000 669.3000 ;
	    RECT 1113.0000 663.3000 1114.2001 670.5000 ;
	    RECT 1120.8000 670.2000 1127.1000 671.4000 ;
	    RECT 1129.8000 671.1000 1131.0000 679.5000 ;
	    RECT 1128.0000 670.2000 1131.0000 671.1000 ;
	    RECT 1115.4000 663.3000 1116.6000 667.5000 ;
	    RECT 1117.8000 663.3000 1119.0000 667.5000 ;
	    RECT 1120.2001 663.3000 1121.4000 669.3000 ;
	    RECT 1122.6000 663.3000 1123.8000 670.2000 ;
	    RECT 1128.0000 669.3000 1128.9000 670.2000 ;
	    RECT 1125.0000 662.4000 1126.2001 669.3000 ;
	    RECT 1127.4000 668.4000 1128.9000 669.3000 ;
	    RECT 1127.4000 663.3000 1128.6000 668.4000 ;
	    RECT 1129.8000 663.3000 1131.0000 669.3000 ;
	    RECT 1151.4000 663.3000 1152.6000 669.3000 ;
	    RECT 1153.8000 663.3000 1155.0000 679.5000 ;
	    RECT 1175.4000 677.4000 1176.6000 678.6000 ;
	    RECT 1177.8000 678.4500 1179.0000 678.6000 ;
	    RECT 1225.8000 678.4500 1227.0000 678.6000 ;
	    RECT 1230.7500 678.4500 1231.6500 680.4000 ;
	    RECT 1232.7001 679.5000 1233.3000 680.7000 ;
	    RECT 1234.5000 679.5000 1238.4000 680.7000 ;
	    RECT 1239.9000 679.5000 1243.5000 680.7000 ;
	    RECT 1244.7001 679.5000 1248.6000 680.7000 ;
	    RECT 1249.8000 679.5000 1251.0000 681.6000 ;
	    RECT 1271.4000 679.5000 1272.6000 683.7000 ;
	    RECT 1273.8000 682.5000 1275.0000 682.8000 ;
	    RECT 1273.8000 680.4000 1275.0000 681.6000 ;
	    RECT 1295.4000 679.5000 1296.6000 683.7000 ;
	    RECT 1324.5000 683.1000 1329.9000 683.7000 ;
	    RECT 1297.8000 682.5000 1299.0000 682.8000 ;
	    RECT 1331.4000 682.5000 1332.3000 683.7000 ;
	    RECT 1350.6000 682.5000 1351.8000 682.8000 ;
	    RECT 1297.8000 680.4000 1299.0000 681.6000 ;
	    RECT 1309.8000 681.4500 1311.0000 681.6000 ;
	    RECT 1324.2001 681.4500 1325.4000 681.6000 ;
	    RECT 1309.8000 680.5500 1325.4000 681.4500 ;
	    RECT 1326.3000 680.7000 1326.6000 682.2000 ;
	    RECT 1309.8000 680.4000 1311.0000 680.5500 ;
	    RECT 1324.2001 680.4000 1325.4000 680.5500 ;
	    RECT 1328.7001 680.4000 1330.5000 681.6000 ;
	    RECT 1331.4000 680.4000 1332.6000 681.6000 ;
	    RECT 1345.8000 681.4500 1347.0000 681.6000 ;
	    RECT 1350.6000 681.4500 1351.8000 681.6000 ;
	    RECT 1345.8000 680.5500 1351.8000 681.4500 ;
	    RECT 1345.8000 680.4000 1347.0000 680.5500 ;
	    RECT 1350.6000 680.4000 1351.8000 680.5500 ;
	    RECT 1326.6000 679.5000 1327.8000 679.8000 ;
	    RECT 1177.8000 677.5500 1231.6500 678.4500 ;
	    RECT 1177.8000 677.4000 1179.0000 677.5500 ;
	    RECT 1225.8000 677.4000 1227.0000 677.5500 ;
	    RECT 1234.5000 677.4000 1235.7001 679.5000 ;
	    RECT 1239.9000 677.4000 1241.1000 679.5000 ;
	    RECT 1244.7001 677.4000 1245.9000 679.5000 ;
	    RECT 1249.8000 678.4500 1251.0000 678.6000 ;
	    RECT 1266.6000 678.4500 1267.8000 678.6000 ;
	    RECT 1249.8000 677.5500 1267.8000 678.4500 ;
	    RECT 1249.8000 677.4000 1251.0000 677.5500 ;
	    RECT 1266.6000 677.4000 1267.8000 677.5500 ;
	    RECT 1271.4000 678.4500 1272.6000 678.6000 ;
	    RECT 1276.2001 678.4500 1277.4000 678.6000 ;
	    RECT 1271.4000 677.5500 1277.4000 678.4500 ;
	    RECT 1271.4000 677.4000 1272.6000 677.5500 ;
	    RECT 1276.2001 677.4000 1277.4000 677.5500 ;
	    RECT 1278.6000 678.4500 1279.8000 678.6000 ;
	    RECT 1295.4000 678.4500 1296.6000 678.6000 ;
	    RECT 1278.6000 677.5500 1296.6000 678.4500 ;
	    RECT 1278.6000 677.4000 1279.8000 677.5500 ;
	    RECT 1295.4000 677.4000 1296.6000 677.5500 ;
	    RECT 1326.6000 677.4000 1327.8000 678.6000 ;
	    RECT 1165.8000 675.4500 1167.0000 675.6000 ;
	    RECT 1173.0000 675.4500 1174.2001 675.6000 ;
	    RECT 1165.8000 674.5500 1174.2001 675.4500 ;
	    RECT 1165.8000 674.4000 1167.0000 674.5500 ;
	    RECT 1173.0000 674.4000 1174.2001 674.5500 ;
	    RECT 1173.0000 673.2000 1174.2001 673.5000 ;
	    RECT 1173.0000 663.3000 1174.2001 669.3000 ;
	    RECT 1175.4000 663.3000 1176.6000 676.5000 ;
	    RECT 1233.0000 676.2000 1235.7001 677.4000 ;
	    RECT 1237.8000 676.2000 1241.1000 677.4000 ;
	    RECT 1242.6000 676.2000 1245.9000 677.4000 ;
	    RECT 1247.4000 676.5000 1248.9000 677.4000 ;
	    RECT 1247.4000 676.2000 1251.0000 676.5000 ;
	    RECT 1177.8000 663.3000 1179.0000 669.3000 ;
	    RECT 1230.6000 663.3000 1231.8000 675.3000 ;
	    RECT 1233.0000 663.3000 1234.2001 676.2000 ;
	    RECT 1235.4000 663.3000 1236.6000 675.3000 ;
	    RECT 1237.8000 663.3000 1239.0000 676.2000 ;
	    RECT 1240.2001 663.3000 1241.4000 675.3000 ;
	    RECT 1242.6000 663.3000 1243.8000 676.2000 ;
	    RECT 1245.0000 663.3000 1246.2001 675.3000 ;
	    RECT 1247.4000 663.3000 1248.6000 676.2000 ;
	    RECT 1266.6000 675.4500 1267.8000 675.6000 ;
	    RECT 1269.0000 675.4500 1270.2001 675.6000 ;
	    RECT 1249.8000 663.3000 1251.0000 675.3000 ;
	    RECT 1266.6000 674.5500 1270.2001 675.4500 ;
	    RECT 1266.6000 674.4000 1267.8000 674.5500 ;
	    RECT 1269.0000 674.4000 1270.2001 674.5500 ;
	    RECT 1269.0000 673.2000 1270.2001 673.5000 ;
	    RECT 1269.0000 663.3000 1270.2001 669.3000 ;
	    RECT 1271.4000 663.3000 1272.6000 676.5000 ;
	    RECT 1293.0000 674.4000 1294.2001 675.6000 ;
	    RECT 1293.0000 673.2000 1294.2001 673.5000 ;
	    RECT 1273.8000 663.3000 1275.0000 669.3000 ;
	    RECT 1293.0000 663.3000 1294.2001 669.3000 ;
	    RECT 1295.4000 663.3000 1296.6000 676.5000 ;
	    RECT 1328.7001 675.3000 1329.6000 680.4000 ;
	    RECT 1353.0000 679.5000 1354.2001 683.7000 ;
	    RECT 1381.8000 682.8000 1383.0000 689.7000 ;
	    RECT 1384.2001 683.7000 1385.4000 689.7000 ;
	    RECT 1381.8000 681.9000 1385.1000 682.8000 ;
	    RECT 1386.6000 682.5000 1387.8000 689.7000 ;
	    RECT 1405.8000 683.7000 1407.0000 689.7000 ;
	    RECT 1409.7001 684.6000 1410.9000 689.7000 ;
	    RECT 1425.0000 686.7000 1426.2001 689.7000 ;
	    RECT 1425.0000 685.5000 1426.2001 685.8000 ;
	    RECT 1408.2001 683.7000 1410.9000 684.6000 ;
	    RECT 1422.6000 684.4500 1423.8000 684.6000 ;
	    RECT 1425.0000 684.4500 1426.2001 684.6000 ;
	    RECT 1405.8000 682.5000 1407.0000 682.8000 ;
	    RECT 1381.8000 679.5000 1383.0000 679.8000 ;
	    RECT 1350.6000 678.4500 1351.8000 678.6000 ;
	    RECT 1353.0000 678.4500 1354.2001 678.6000 ;
	    RECT 1350.6000 677.5500 1354.2001 678.4500 ;
	    RECT 1350.6000 677.4000 1351.8000 677.5500 ;
	    RECT 1353.0000 677.4000 1354.2001 677.5500 ;
	    RECT 1367.4000 678.4500 1368.6000 678.6000 ;
	    RECT 1381.8000 678.4500 1383.0000 678.6000 ;
	    RECT 1367.4000 677.5500 1383.0000 678.4500 ;
	    RECT 1367.4000 677.4000 1368.6000 677.5500 ;
	    RECT 1381.8000 677.4000 1383.0000 677.5500 ;
	    RECT 1384.2001 677.4000 1385.1000 681.9000 ;
	    RECT 1386.6000 681.4500 1387.8000 681.6000 ;
	    RECT 1405.8000 681.4500 1407.0000 681.6000 ;
	    RECT 1386.6000 680.5500 1407.0000 681.4500 ;
	    RECT 1386.6000 680.4000 1387.8000 680.5500 ;
	    RECT 1405.8000 680.4000 1407.0000 680.5500 ;
	    RECT 1408.2001 679.5000 1409.4000 683.7000 ;
	    RECT 1422.6000 683.5500 1426.2001 684.4500 ;
	    RECT 1422.6000 683.4000 1423.8000 683.5500 ;
	    RECT 1425.0000 683.4000 1426.2001 683.5500 ;
	    RECT 1427.4000 682.5000 1428.6000 689.7000 ;
	    RECT 1427.4000 681.4500 1428.6000 681.6000 ;
	    RECT 1439.4000 681.4500 1440.6000 681.6000 ;
	    RECT 1427.4000 680.5500 1440.6000 681.4500 ;
	    RECT 1451.4000 680.7000 1452.6000 689.7000 ;
	    RECT 1456.8000 681.3000 1458.0000 689.7000 ;
	    RECT 1482.6000 684.0000 1483.8000 689.7000 ;
	    RECT 1485.0000 684.9000 1486.2001 689.7000 ;
	    RECT 1487.4000 684.0000 1488.6000 689.7000 ;
	    RECT 1482.6000 683.7000 1488.6000 684.0000 ;
	    RECT 1489.8000 683.7000 1491.0000 689.7000 ;
	    RECT 1514.7001 683.7000 1515.9000 689.7000 ;
	    RECT 1518.6000 683.7000 1519.8000 689.7000 ;
	    RECT 1521.0000 686.7000 1522.2001 689.7000 ;
	    RECT 1547.4000 686.7000 1548.6000 689.7000 ;
	    RECT 1520.7001 685.5000 1521.9000 685.8000 ;
	    RECT 1547.7001 685.5000 1548.9000 685.8000 ;
	    RECT 1482.9000 683.1000 1488.3000 683.7000 ;
	    RECT 1489.8000 682.5000 1490.7001 683.7000 ;
	    RECT 1456.8000 680.7000 1459.5000 681.3000 ;
	    RECT 1427.4000 680.4000 1428.6000 680.5500 ;
	    RECT 1439.4000 680.4000 1440.6000 680.5500 ;
	    RECT 1457.1000 680.4000 1459.5000 680.7000 ;
	    RECT 1482.6000 680.4000 1483.8000 681.6000 ;
	    RECT 1484.7001 680.7000 1485.0000 682.2000 ;
	    RECT 1487.1000 680.4000 1488.9000 681.6000 ;
	    RECT 1489.8000 680.4000 1491.0000 681.6000 ;
	    RECT 1511.4000 681.4500 1512.6000 681.6000 ;
	    RECT 1516.2001 681.4500 1517.4000 681.6000 ;
	    RECT 1511.4000 680.5500 1517.4000 681.4500 ;
	    RECT 1511.4000 680.4000 1512.6000 680.5500 ;
	    RECT 1516.2001 680.4000 1517.4000 680.5500 ;
	    RECT 1386.6000 678.6000 1387.8000 679.5000 ;
	    RECT 1297.8000 663.3000 1299.0000 669.3000 ;
	    RECT 1324.2001 663.3000 1325.4000 675.3000 ;
	    RECT 1328.1000 674.4000 1329.6000 675.3000 ;
	    RECT 1331.4000 674.4000 1332.6000 675.6000 ;
	    RECT 1328.1000 663.3000 1329.3000 674.4000 ;
	    RECT 1330.5000 672.6000 1331.4000 673.5000 ;
	    RECT 1330.2001 671.4000 1331.4000 672.6000 ;
	    RECT 1330.5000 663.3000 1331.7001 669.3000 ;
	    RECT 1350.6000 663.3000 1351.8000 669.3000 ;
	    RECT 1353.0000 663.3000 1354.2001 676.5000 ;
	    RECT 1384.2001 676.2000 1386.0000 677.4000 ;
	    RECT 1355.4000 675.4500 1356.6000 675.6000 ;
	    RECT 1369.8000 675.4500 1371.0000 675.6000 ;
	    RECT 1355.4000 674.5500 1371.0000 675.4500 ;
	    RECT 1384.2001 675.3000 1385.1000 676.2000 ;
	    RECT 1386.9000 675.3000 1387.8000 678.6000 ;
	    RECT 1408.2001 678.4500 1409.4000 678.6000 ;
	    RECT 1413.0000 678.4500 1414.2001 678.6000 ;
	    RECT 1408.2001 677.5500 1414.2001 678.4500 ;
	    RECT 1408.2001 677.4000 1409.4000 677.5500 ;
	    RECT 1413.0000 677.4000 1414.2001 677.5500 ;
	    RECT 1355.4000 674.4000 1356.6000 674.5500 ;
	    RECT 1369.8000 674.4000 1371.0000 674.5500 ;
	    RECT 1381.8000 674.4000 1385.1000 675.3000 ;
	    RECT 1355.4000 673.2000 1356.6000 673.5000 ;
	    RECT 1355.4000 663.3000 1356.6000 669.3000 ;
	    RECT 1381.8000 663.3000 1383.0000 674.4000 ;
	    RECT 1384.2001 663.3000 1385.4000 673.5000 ;
	    RECT 1386.6000 663.3000 1387.8000 675.3000 ;
	    RECT 1405.8000 663.3000 1407.0000 669.3000 ;
	    RECT 1408.2001 663.3000 1409.4000 676.5000 ;
	    RECT 1410.6000 675.4500 1411.8000 675.6000 ;
	    RECT 1425.0000 675.4500 1426.2001 675.6000 ;
	    RECT 1410.6000 674.5500 1426.2001 675.4500 ;
	    RECT 1410.6000 674.4000 1411.8000 674.5500 ;
	    RECT 1425.0000 674.4000 1426.2001 674.5500 ;
	    RECT 1410.6000 673.2000 1411.8000 673.5000 ;
	    RECT 1410.6000 663.3000 1411.8000 669.3000 ;
	    RECT 1425.0000 663.3000 1426.2001 669.3000 ;
	    RECT 1427.4000 663.3000 1428.6000 679.5000 ;
	    RECT 1453.8000 677.4000 1455.0000 678.6000 ;
	    RECT 1455.9000 677.4000 1456.2001 678.6000 ;
	    RECT 1451.4000 676.5000 1452.6000 676.8000 ;
	    RECT 1458.6000 676.5000 1459.5000 680.4000 ;
	    RECT 1485.0000 679.5000 1486.2001 679.8000 ;
	    RECT 1485.0000 677.4000 1486.2001 678.6000 ;
	    RECT 1432.2001 675.4500 1433.4000 675.6000 ;
	    RECT 1451.4000 675.4500 1452.6000 675.6000 ;
	    RECT 1432.2001 674.5500 1452.6000 675.4500 ;
	    RECT 1432.2001 674.4000 1433.4000 674.5500 ;
	    RECT 1451.4000 674.4000 1452.6000 674.5500 ;
	    RECT 1458.6000 675.4500 1459.8000 675.6000 ;
	    RECT 1461.0000 675.4500 1462.2001 675.6000 ;
	    RECT 1458.6000 674.5500 1462.2001 675.4500 ;
	    RECT 1487.1000 675.3000 1488.0000 680.4000 ;
	    RECT 1516.2001 679.2000 1517.4000 679.5000 ;
	    RECT 1506.6000 678.4500 1507.8000 678.6000 ;
	    RECT 1513.8000 678.4500 1515.0000 678.6000 ;
	    RECT 1506.6000 677.5500 1515.0000 678.4500 ;
	    RECT 1518.6000 678.3000 1519.5000 683.7000 ;
	    RECT 1521.0000 683.4000 1522.2001 684.6000 ;
	    RECT 1525.8000 684.4500 1527.0000 684.6000 ;
	    RECT 1547.4000 684.4500 1548.6000 684.6000 ;
	    RECT 1525.8000 683.5500 1548.6000 684.4500 ;
	    RECT 1549.8000 683.7000 1551.0000 689.7000 ;
	    RECT 1553.7001 683.7000 1554.9000 689.7000 ;
	    RECT 1525.8000 683.4000 1527.0000 683.5500 ;
	    RECT 1547.4000 683.4000 1548.6000 683.5500 ;
	    RECT 1521.0000 678.4500 1522.2001 678.6000 ;
	    RECT 1523.4000 678.4500 1524.6000 678.6000 ;
	    RECT 1506.6000 677.4000 1507.8000 677.5500 ;
	    RECT 1513.8000 677.4000 1515.0000 677.5500 ;
	    RECT 1515.9000 676.8000 1516.2001 678.3000 ;
	    RECT 1518.6000 677.4000 1520.1000 678.3000 ;
	    RECT 1521.0000 677.5500 1524.6000 678.4500 ;
	    RECT 1521.0000 677.4000 1522.2001 677.5500 ;
	    RECT 1523.4000 677.4000 1524.6000 677.5500 ;
	    RECT 1525.8000 678.4500 1527.0000 678.6000 ;
	    RECT 1547.4000 678.4500 1548.6000 678.6000 ;
	    RECT 1525.8000 677.5500 1548.6000 678.4500 ;
	    RECT 1550.1000 678.3000 1551.0000 683.7000 ;
	    RECT 1552.2001 681.4500 1553.4000 681.6000 ;
	    RECT 1557.0000 681.4500 1558.2001 681.6000 ;
	    RECT 1552.2001 680.5500 1558.2001 681.4500 ;
	    RECT 1552.2001 680.4000 1553.4000 680.5500 ;
	    RECT 1557.0000 680.4000 1558.2001 680.5500 ;
	    RECT 1552.2001 679.2000 1553.4000 679.5000 ;
	    RECT 1525.8000 677.4000 1527.0000 677.5500 ;
	    RECT 1547.4000 677.4000 1548.6000 677.5500 ;
	    RECT 1549.5000 677.4000 1551.0000 678.3000 ;
	    RECT 1553.4000 676.8000 1553.7001 678.3000 ;
	    RECT 1554.6000 677.4000 1555.8000 678.6000 ;
	    RECT 1458.6000 674.4000 1459.8000 674.5500 ;
	    RECT 1461.0000 674.4000 1462.2001 674.5500 ;
	    RECT 1456.2001 673.5000 1457.4000 673.8000 ;
	    RECT 1441.8000 672.4500 1443.0000 672.6000 ;
	    RECT 1451.4000 672.4500 1452.6000 672.6000 ;
	    RECT 1456.2001 672.4500 1457.4000 672.6000 ;
	    RECT 1441.8000 671.5500 1457.4000 672.4500 ;
	    RECT 1441.8000 671.4000 1443.0000 671.5500 ;
	    RECT 1451.4000 671.4000 1452.6000 671.5500 ;
	    RECT 1456.2001 671.4000 1457.4000 671.5500 ;
	    RECT 1458.6000 670.5000 1459.5000 673.5000 ;
	    RECT 1454.1000 669.6000 1459.5000 670.5000 ;
	    RECT 1454.1000 669.3000 1455.0000 669.6000 ;
	    RECT 1451.4000 663.3000 1452.6000 669.3000 ;
	    RECT 1453.8000 663.3000 1455.0000 669.3000 ;
	    RECT 1458.6000 669.3000 1459.5000 669.6000 ;
	    RECT 1456.2001 663.3000 1457.4000 668.7000 ;
	    RECT 1458.6000 663.3000 1459.8000 669.3000 ;
	    RECT 1482.6000 663.3000 1483.8000 675.3000 ;
	    RECT 1486.5000 674.4000 1488.0000 675.3000 ;
	    RECT 1489.8000 675.4500 1491.0000 675.6000 ;
	    RECT 1497.0000 675.4500 1498.2001 675.6000 ;
	    RECT 1489.8000 674.5500 1498.2001 675.4500 ;
	    RECT 1521.0000 675.3000 1521.9000 676.5000 ;
	    RECT 1547.7001 675.3000 1548.6000 676.5000 ;
	    RECT 1489.8000 674.4000 1491.0000 674.5500 ;
	    RECT 1497.0000 674.4000 1498.2001 674.5500 ;
	    RECT 1513.8000 674.4000 1519.8000 675.3000 ;
	    RECT 1486.5000 663.3000 1487.7001 674.4000 ;
	    RECT 1488.9000 672.6000 1489.8000 673.5000 ;
	    RECT 1488.6000 671.4000 1489.8000 672.6000 ;
	    RECT 1488.9000 663.3000 1490.1000 669.3000 ;
	    RECT 1513.8000 663.3000 1515.0000 674.4000 ;
	    RECT 1516.2001 663.3000 1517.4000 673.5000 ;
	    RECT 1518.6000 663.3000 1519.8000 674.4000 ;
	    RECT 1521.0000 663.3000 1522.2001 675.3000 ;
	    RECT 1547.4000 663.3000 1548.6000 675.3000 ;
	    RECT 1549.8000 674.4000 1555.8000 675.3000 ;
	    RECT 1549.8000 663.3000 1551.0000 674.4000 ;
	    RECT 1552.2001 663.3000 1553.4000 673.5000 ;
	    RECT 1554.6000 663.3000 1555.8000 674.4000 ;
	    RECT 1.2000 660.6000 1569.0000 662.4000 ;
	    RECT 18.6000 653.7000 19.8000 659.7000 ;
	    RECT 18.6000 649.5000 19.8000 649.8000 ;
	    RECT 18.6000 647.4000 19.8000 648.6000 ;
	    RECT 21.0000 646.5000 22.2000 659.7000 ;
	    RECT 23.4000 653.7000 24.6000 659.7000 ;
	    RECT 42.6000 653.7000 43.8000 659.7000 ;
	    RECT 42.6000 649.5000 43.8000 649.8000 ;
	    RECT 40.2000 648.4500 41.4000 648.6000 ;
	    RECT 42.6000 648.4500 43.8000 648.6000 ;
	    RECT 40.2000 647.5500 43.8000 648.4500 ;
	    RECT 40.2000 647.4000 41.4000 647.5500 ;
	    RECT 42.6000 647.4000 43.8000 647.5500 ;
	    RECT 45.0000 646.5000 46.2000 659.7000 ;
	    RECT 47.4000 653.7000 48.6000 659.7000 ;
	    RECT 72.3000 653.7000 73.5000 659.7000 ;
	    RECT 72.6000 650.4000 73.8000 651.6000 ;
	    RECT 72.6000 649.5000 73.5000 650.4000 ;
	    RECT 74.7000 648.6000 75.9000 659.7000 ;
	    RECT 66.6000 648.4500 67.8000 648.6000 ;
	    RECT 71.4000 648.4500 72.6000 648.6000 ;
	    RECT 66.6000 647.5500 72.6000 648.4500 ;
	    RECT 66.6000 647.4000 67.8000 647.5500 ;
	    RECT 71.4000 647.4000 72.6000 647.5500 ;
	    RECT 74.4000 647.7000 75.9000 648.6000 ;
	    RECT 78.6000 647.7000 79.8000 659.7000 ;
	    RECT 21.0000 645.4500 22.2000 645.6000 ;
	    RECT 42.6000 645.4500 43.8000 645.6000 ;
	    RECT 21.0000 644.5500 43.8000 645.4500 ;
	    RECT 21.0000 644.4000 22.2000 644.5500 ;
	    RECT 42.6000 644.4000 43.8000 644.5500 ;
	    RECT 45.0000 645.4500 46.2000 645.6000 ;
	    RECT 47.4000 645.4500 48.6000 645.6000 ;
	    RECT 45.0000 644.5500 48.6000 645.4500 ;
	    RECT 45.0000 644.4000 46.2000 644.5500 ;
	    RECT 47.4000 644.4000 48.6000 644.5500 ;
	    RECT 21.0000 639.3000 22.2000 643.5000 ;
	    RECT 23.4000 642.4500 24.6000 642.6000 ;
	    RECT 40.2000 642.4500 41.4000 642.6000 ;
	    RECT 23.4000 641.5500 41.4000 642.4500 ;
	    RECT 23.4000 641.4000 24.6000 641.5500 ;
	    RECT 40.2000 641.4000 41.4000 641.5500 ;
	    RECT 23.4000 640.2000 24.6000 640.5000 ;
	    RECT 45.0000 639.3000 46.2000 643.5000 ;
	    RECT 74.4000 642.6000 75.3000 647.7000 ;
	    RECT 76.2000 645.4500 77.4000 645.6000 ;
	    RECT 76.2000 644.5500 82.0500 645.4500 ;
	    RECT 76.2000 644.4000 77.4000 644.5500 ;
	    RECT 76.2000 643.2000 77.4000 643.5000 ;
	    RECT 47.4000 642.4500 48.6000 642.6000 ;
	    RECT 52.2000 642.4500 53.4000 642.6000 ;
	    RECT 47.4000 641.5500 53.4000 642.4500 ;
	    RECT 47.4000 641.4000 48.6000 641.5500 ;
	    RECT 52.2000 641.4000 53.4000 641.5500 ;
	    RECT 71.4000 641.4000 72.6000 642.6000 ;
	    RECT 73.5000 641.4000 75.3000 642.6000 ;
	    RECT 77.4000 640.8000 77.7000 642.3000 ;
	    RECT 78.6000 641.4000 79.8000 642.6000 ;
	    RECT 81.1500 642.4500 82.0500 644.5500 ;
	    RECT 93.0000 643.5000 94.2000 659.7000 ;
	    RECT 95.4000 653.7000 96.6000 659.7000 ;
	    RECT 114.6000 653.7000 115.8000 659.7000 ;
	    RECT 114.6000 649.5000 115.8000 649.8000 ;
	    RECT 114.6000 647.4000 115.8000 648.6000 ;
	    RECT 117.0000 646.5000 118.2000 659.7000 ;
	    RECT 119.4000 653.7000 120.6000 659.7000 ;
	    RECT 131.4000 653.7000 132.6000 659.7000 ;
	    RECT 117.0000 645.4500 118.2000 645.6000 ;
	    RECT 121.8000 645.4500 123.0000 645.6000 ;
	    RECT 117.0000 644.5500 123.0000 645.4500 ;
	    RECT 117.0000 644.4000 118.2000 644.5500 ;
	    RECT 121.8000 644.4000 123.0000 644.5500 ;
	    RECT 133.8000 643.5000 135.0000 659.7000 ;
	    RECT 138.6000 657.4500 139.8000 657.6000 ;
	    RECT 162.6000 657.4500 163.8000 657.6000 ;
	    RECT 138.6000 656.5500 163.8000 657.4500 ;
	    RECT 138.6000 656.4000 139.8000 656.5500 ;
	    RECT 162.6000 656.4000 163.8000 656.5500 ;
	    RECT 165.0000 647.7000 166.2000 659.7000 ;
	    RECT 168.9000 647.7000 171.9000 659.7000 ;
	    RECT 174.6000 647.7000 175.8000 659.7000 ;
	    RECT 213.0000 647.7000 214.2000 659.7000 ;
	    RECT 216.9000 647.7000 219.9000 659.7000 ;
	    RECT 222.6000 647.7000 223.8000 659.7000 ;
	    RECT 241.8000 647.7000 243.0000 659.7000 ;
	    RECT 245.7000 648.9000 246.9000 659.7000 ;
	    RECT 244.2000 647.7000 246.9000 648.9000 ;
	    RECT 277.8000 647.7000 279.0000 659.7000 ;
	    RECT 281.7000 647.7000 284.7000 659.7000 ;
	    RECT 287.4000 647.7000 288.6000 659.7000 ;
	    RECT 167.4000 644.4000 168.6000 645.6000 ;
	    RECT 165.0000 643.5000 166.2000 643.8000 ;
	    RECT 170.1000 643.5000 171.0000 647.7000 ;
	    RECT 172.2000 645.4500 173.4000 645.6000 ;
	    RECT 179.4000 645.4500 180.6000 645.6000 ;
	    RECT 172.2000 644.5500 180.6000 645.4500 ;
	    RECT 172.2000 644.4000 173.4000 644.5500 ;
	    RECT 179.4000 644.4000 180.6000 644.5500 ;
	    RECT 215.4000 644.4000 216.6000 645.6000 ;
	    RECT 217.8000 643.5000 218.7000 647.7000 ;
	    RECT 220.2000 644.4000 221.4000 645.6000 ;
	    RECT 222.6000 643.5000 223.8000 643.8000 ;
	    RECT 244.5000 643.5000 245.4000 647.7000 ;
	    RECT 246.6000 646.5000 247.8000 646.8000 ;
	    RECT 246.6000 645.4500 247.8000 645.6000 ;
	    RECT 253.8000 645.4500 255.0000 645.6000 ;
	    RECT 246.6000 644.5500 255.0000 645.4500 ;
	    RECT 246.6000 644.4000 247.8000 644.5500 ;
	    RECT 253.8000 644.4000 255.0000 644.5500 ;
	    RECT 280.2000 644.4000 281.4000 645.6000 ;
	    RECT 277.8000 643.5000 279.0000 643.8000 ;
	    RECT 282.9000 643.5000 283.8000 647.7000 ;
	    RECT 285.0000 644.4000 286.2000 645.6000 ;
	    RECT 299.4000 643.5000 300.6000 659.7000 ;
	    RECT 301.8000 653.7000 303.0000 659.7000 ;
	    RECT 304.2000 657.4500 305.4000 657.6000 ;
	    RECT 311.4000 657.4500 312.6000 657.6000 ;
	    RECT 304.2000 656.5500 312.6000 657.4500 ;
	    RECT 304.2000 656.4000 305.4000 656.5500 ;
	    RECT 311.4000 656.4000 312.6000 656.5500 ;
	    RECT 321.0000 653.7000 322.2000 659.7000 ;
	    RECT 323.4000 646.5000 324.6000 659.7000 ;
	    RECT 325.8000 653.7000 327.0000 659.7000 ;
	    RECT 340.2000 653.7000 341.4000 659.7000 ;
	    RECT 325.8000 649.5000 327.0000 649.8000 ;
	    RECT 325.8000 647.4000 327.0000 648.6000 ;
	    RECT 323.4000 644.4000 324.6000 645.6000 ;
	    RECT 342.6000 643.5000 343.8000 659.7000 ;
	    RECT 361.8000 653.7000 363.0000 659.7000 ;
	    RECT 361.8000 649.5000 363.0000 649.8000 ;
	    RECT 345.0000 648.4500 346.2000 648.6000 ;
	    RECT 361.8000 648.4500 363.0000 648.6000 ;
	    RECT 345.0000 647.5500 363.0000 648.4500 ;
	    RECT 345.0000 647.4000 346.2000 647.5500 ;
	    RECT 361.8000 647.4000 363.0000 647.5500 ;
	    RECT 364.2000 646.5000 365.4000 659.7000 ;
	    RECT 366.6000 653.7000 367.8000 659.7000 ;
	    RECT 405.0000 659.4000 406.2000 660.6000 ;
	    RECT 412.2000 659.4000 413.4000 660.6000 ;
	    RECT 424.2000 657.4500 425.4000 657.6000 ;
	    RECT 445.8000 657.4500 447.0000 657.6000 ;
	    RECT 424.2000 656.5500 447.0000 657.4500 ;
	    RECT 424.2000 656.4000 425.4000 656.5500 ;
	    RECT 445.8000 656.4000 447.0000 656.5500 ;
	    RECT 419.4000 654.4500 420.6000 654.6000 ;
	    RECT 450.6000 654.4500 451.8000 654.6000 ;
	    RECT 419.4000 653.5500 451.8000 654.4500 ;
	    RECT 498.6000 653.7000 499.8000 659.7000 ;
	    RECT 501.0000 654.6000 502.2000 659.7000 ;
	    RECT 500.7000 653.7000 502.2000 654.6000 ;
	    RECT 503.4000 653.7000 504.6000 660.6000 ;
	    RECT 419.4000 653.4000 420.6000 653.5500 ;
	    RECT 450.6000 653.4000 451.8000 653.5500 ;
	    RECT 500.7000 652.8000 501.6000 653.7000 ;
	    RECT 505.8000 652.8000 507.0000 659.7000 ;
	    RECT 508.2000 653.7000 509.4000 659.7000 ;
	    RECT 510.6000 655.5000 511.8000 659.7000 ;
	    RECT 513.0000 655.5000 514.2000 659.7000 ;
	    RECT 498.6000 651.9000 501.6000 652.8000 ;
	    RECT 364.2000 645.4500 365.4000 645.6000 ;
	    RECT 429.0000 645.4500 430.2000 645.6000 ;
	    RECT 364.2000 644.5500 430.2000 645.4500 ;
	    RECT 364.2000 644.4000 365.4000 644.5500 ;
	    RECT 429.0000 644.4000 430.2000 644.5500 ;
	    RECT 498.6000 643.5000 499.8000 651.9000 ;
	    RECT 502.5000 651.6000 508.8000 652.8000 ;
	    RECT 515.4000 652.5000 516.6000 659.7000 ;
	    RECT 517.8000 653.7000 519.0000 659.7000 ;
	    RECT 520.2000 652.5000 521.4000 659.7000 ;
	    RECT 522.6000 653.7000 523.8000 659.7000 ;
	    RECT 502.5000 651.0000 503.4000 651.6000 ;
	    RECT 501.0000 649.8000 503.4000 651.0000 ;
	    RECT 507.9000 650.7000 516.6000 651.6000 ;
	    RECT 504.9000 649.8000 507.0000 650.7000 ;
	    RECT 504.9000 649.5000 514.2000 649.8000 ;
	    RECT 506.1000 648.9000 514.2000 649.5000 ;
	    RECT 513.0000 648.6000 514.2000 648.9000 ;
	    RECT 515.7000 649.5000 516.6000 650.7000 ;
	    RECT 517.5000 650.4000 521.4000 651.6000 ;
	    RECT 525.0000 650.4000 526.2000 659.7000 ;
	    RECT 527.4000 655.5000 528.6000 659.7000 ;
	    RECT 529.8000 655.5000 531.0000 659.7000 ;
	    RECT 532.2000 655.5000 533.4000 659.7000 ;
	    RECT 534.6000 653.7000 535.8000 659.7000 ;
	    RECT 529.8000 651.6000 536.1000 652.8000 ;
	    RECT 537.0000 651.6000 538.2000 659.7000 ;
	    RECT 539.4000 653.7000 540.6000 659.7000 ;
	    RECT 541.8000 652.8000 543.0000 659.7000 ;
	    RECT 544.2000 653.7000 545.4000 659.7000 ;
	    RECT 541.8000 651.9000 545.7000 652.8000 ;
	    RECT 546.6000 652.5000 547.8000 659.7000 ;
	    RECT 549.0000 653.7000 550.2000 659.7000 ;
	    RECT 563.4000 653.7000 564.6000 659.7000 ;
	    RECT 537.0000 650.4000 540.9000 651.6000 ;
	    RECT 527.4000 649.5000 528.6000 649.8000 ;
	    RECT 515.7000 648.6000 528.6000 649.5000 ;
	    RECT 532.2000 649.5000 533.4000 649.8000 ;
	    RECT 544.8000 649.5000 545.7000 651.9000 ;
	    RECT 546.6000 650.4000 547.8000 651.6000 ;
	    RECT 532.2000 648.6000 545.7000 649.5000 ;
	    RECT 503.4000 647.4000 504.6000 648.6000 ;
	    RECT 508.5000 647.7000 509.7000 648.0000 ;
	    RECT 505.5000 646.8000 543.9000 647.7000 ;
	    RECT 542.7000 646.5000 543.9000 646.8000 ;
	    RECT 544.8000 645.9000 545.7000 648.6000 ;
	    RECT 546.6000 648.0000 547.8000 649.5000 ;
	    RECT 546.6000 646.8000 548.1000 648.0000 ;
	    RECT 500.7000 645.0000 507.3000 645.9000 ;
	    RECT 500.7000 644.7000 501.9000 645.0000 ;
	    RECT 508.2000 644.4000 509.4000 645.6000 ;
	    RECT 510.3000 645.0000 535.8000 645.9000 ;
	    RECT 544.8000 645.0000 546.0000 645.9000 ;
	    RECT 534.6000 644.1000 535.8000 645.0000 ;
	    RECT 93.0000 642.4500 94.2000 642.6000 ;
	    RECT 81.1500 641.5500 94.2000 642.4500 ;
	    RECT 93.0000 641.4000 94.2000 641.5500 ;
	    RECT 47.4000 640.2000 48.6000 640.5000 ;
	    RECT 71.7000 639.3000 72.6000 640.5000 ;
	    RECT 74.1000 639.3000 79.5000 639.9000 ;
	    RECT 19.5000 638.4000 22.2000 639.3000 ;
	    RECT 19.5000 633.3000 20.7000 638.4000 ;
	    RECT 23.4000 633.3000 24.6000 639.3000 ;
	    RECT 43.5000 638.4000 46.2000 639.3000 ;
	    RECT 43.5000 633.3000 44.7000 638.4000 ;
	    RECT 47.4000 633.3000 48.6000 639.3000 ;
	    RECT 71.4000 633.3000 72.6000 639.3000 ;
	    RECT 73.8000 639.0000 79.8000 639.3000 ;
	    RECT 73.8000 633.3000 75.0000 639.0000 ;
	    RECT 76.2000 633.3000 77.4000 638.1000 ;
	    RECT 78.6000 633.3000 79.8000 639.0000 ;
	    RECT 93.0000 633.3000 94.2000 640.5000 ;
	    RECT 95.4000 639.4500 96.6000 639.6000 ;
	    RECT 112.2000 639.4500 113.4000 639.6000 ;
	    RECT 95.4000 638.5500 113.4000 639.4500 ;
	    RECT 117.0000 639.3000 118.2000 643.5000 ;
	    RECT 167.4000 643.2000 168.6000 643.5000 ;
	    RECT 172.2000 643.2000 173.4000 643.5000 ;
	    RECT 215.4000 643.2000 216.6000 643.5000 ;
	    RECT 220.2000 643.2000 221.4000 643.5000 ;
	    RECT 280.2000 643.2000 281.4000 643.5000 ;
	    RECT 285.0000 643.2000 286.2000 643.5000 ;
	    RECT 119.4000 641.4000 120.6000 642.6000 ;
	    RECT 133.8000 642.4500 135.0000 642.6000 ;
	    RECT 165.0000 642.4500 166.2000 642.6000 ;
	    RECT 133.8000 641.5500 166.2000 642.4500 ;
	    RECT 133.8000 641.4000 135.0000 641.5500 ;
	    RECT 165.0000 641.4000 166.2000 641.5500 ;
	    RECT 167.4000 641.4000 168.9000 642.3000 ;
	    RECT 169.8000 641.4000 171.0000 642.6000 ;
	    RECT 174.6000 642.4500 175.8000 642.6000 ;
	    RECT 177.0000 642.4500 178.2000 642.6000 ;
	    RECT 119.4000 640.2000 120.6000 640.5000 ;
	    RECT 124.2000 639.4500 125.4000 639.6000 ;
	    RECT 131.4000 639.4500 132.6000 639.6000 ;
	    RECT 95.4000 638.4000 96.6000 638.5500 ;
	    RECT 112.2000 638.4000 113.4000 638.5500 ;
	    RECT 115.5000 638.4000 118.2000 639.3000 ;
	    RECT 95.4000 637.2000 96.6000 637.5000 ;
	    RECT 95.4000 633.3000 96.6000 636.3000 ;
	    RECT 115.5000 633.3000 116.7000 638.4000 ;
	    RECT 119.4000 633.3000 120.6000 639.3000 ;
	    RECT 124.2000 638.5500 132.6000 639.4500 ;
	    RECT 124.2000 638.4000 125.4000 638.5500 ;
	    RECT 131.4000 638.4000 132.6000 638.5500 ;
	    RECT 131.4000 637.2000 132.6000 637.5000 ;
	    RECT 131.4000 633.3000 132.6000 636.3000 ;
	    RECT 133.8000 633.3000 135.0000 640.5000 ;
	    RECT 167.4000 639.3000 168.3000 641.4000 ;
	    RECT 173.4000 640.8000 173.7000 642.3000 ;
	    RECT 174.6000 641.5500 178.2000 642.4500 ;
	    RECT 174.6000 641.4000 175.8000 641.5500 ;
	    RECT 177.0000 641.4000 178.2000 641.5500 ;
	    RECT 189.0000 642.4500 190.2000 642.6000 ;
	    RECT 213.0000 642.4500 214.2000 642.6000 ;
	    RECT 189.0000 641.5500 214.2000 642.4500 ;
	    RECT 189.0000 641.4000 190.2000 641.5500 ;
	    RECT 213.0000 641.4000 214.2000 641.5500 ;
	    RECT 215.1000 640.8000 215.4000 642.3000 ;
	    RECT 217.8000 641.4000 219.0000 642.6000 ;
	    RECT 219.9000 641.4000 221.4000 642.3000 ;
	    RECT 222.6000 641.4000 223.8000 642.6000 ;
	    RECT 244.2000 642.4500 245.4000 642.6000 ;
	    RECT 270.6000 642.4500 271.8000 642.6000 ;
	    RECT 244.2000 641.5500 271.8000 642.4500 ;
	    RECT 244.2000 641.4000 245.4000 641.5500 ;
	    RECT 270.6000 641.4000 271.8000 641.5500 ;
	    RECT 275.4000 642.4500 276.6000 642.6000 ;
	    RECT 277.8000 642.4500 279.0000 642.6000 ;
	    RECT 275.4000 641.5500 279.0000 642.4500 ;
	    RECT 275.4000 641.4000 276.6000 641.5500 ;
	    RECT 277.8000 641.4000 279.0000 641.5500 ;
	    RECT 280.2000 641.4000 281.7000 642.3000 ;
	    RECT 282.6000 641.4000 283.8000 642.6000 ;
	    RECT 170.1000 639.3000 175.5000 639.9000 ;
	    RECT 213.3000 639.3000 218.7000 639.9000 ;
	    RECT 220.5000 639.3000 221.4000 641.4000 ;
	    RECT 239.4000 639.4500 240.6000 639.6000 ;
	    RECT 241.8000 639.4500 243.0000 639.6000 ;
	    RECT 165.0000 634.2000 166.2000 639.3000 ;
	    RECT 167.4000 635.1000 168.6000 639.3000 ;
	    RECT 169.8000 639.0000 175.8000 639.3000 ;
	    RECT 169.8000 634.2000 171.0000 639.0000 ;
	    RECT 165.0000 633.3000 171.0000 634.2000 ;
	    RECT 172.2000 633.3000 173.4000 638.1000 ;
	    RECT 174.6000 633.3000 175.8000 639.0000 ;
	    RECT 213.0000 639.0000 219.0000 639.3000 ;
	    RECT 213.0000 633.3000 214.2000 639.0000 ;
	    RECT 215.4000 633.3000 216.6000 638.1000 ;
	    RECT 217.8000 634.2000 219.0000 639.0000 ;
	    RECT 220.2000 635.1000 221.4000 639.3000 ;
	    RECT 222.6000 634.2000 223.8000 639.3000 ;
	    RECT 239.4000 638.5500 243.0000 639.4500 ;
	    RECT 239.4000 638.4000 240.6000 638.5500 ;
	    RECT 241.8000 638.4000 243.0000 638.5500 ;
	    RECT 241.8000 637.2000 243.0000 637.5000 ;
	    RECT 244.5000 636.3000 245.4000 640.5000 ;
	    RECT 280.2000 639.3000 281.1000 641.4000 ;
	    RECT 286.2000 640.8000 286.5000 642.3000 ;
	    RECT 287.4000 641.4000 288.6000 642.6000 ;
	    RECT 289.8000 642.4500 291.0000 642.6000 ;
	    RECT 299.4000 642.4500 300.6000 642.6000 ;
	    RECT 289.8000 641.5500 300.6000 642.4500 ;
	    RECT 289.8000 641.4000 291.0000 641.5500 ;
	    RECT 299.4000 641.4000 300.6000 641.5500 ;
	    RECT 321.0000 641.4000 322.2000 642.6000 ;
	    RECT 282.9000 639.3000 288.3000 639.9000 ;
	    RECT 217.8000 633.3000 223.8000 634.2000 ;
	    RECT 241.8000 633.3000 243.0000 636.3000 ;
	    RECT 244.2000 633.3000 245.4000 636.3000 ;
	    RECT 246.6000 633.3000 247.8000 636.3000 ;
	    RECT 277.8000 634.2000 279.0000 639.3000 ;
	    RECT 280.2000 635.1000 281.4000 639.3000 ;
	    RECT 282.6000 639.0000 288.6000 639.3000 ;
	    RECT 282.6000 634.2000 283.8000 639.0000 ;
	    RECT 277.8000 633.3000 283.8000 634.2000 ;
	    RECT 285.0000 633.3000 286.2000 638.1000 ;
	    RECT 287.4000 633.3000 288.6000 639.0000 ;
	    RECT 299.4000 633.3000 300.6000 640.5000 ;
	    RECT 321.0000 640.2000 322.2000 640.5000 ;
	    RECT 301.8000 639.4500 303.0000 639.6000 ;
	    RECT 306.6000 639.4500 307.8000 639.6000 ;
	    RECT 301.8000 638.5500 307.8000 639.4500 ;
	    RECT 323.4000 639.3000 324.6000 643.5000 ;
	    RECT 342.6000 642.4500 343.8000 642.6000 ;
	    RECT 361.8000 642.4500 363.0000 642.6000 ;
	    RECT 342.6000 641.5500 363.0000 642.4500 ;
	    RECT 342.6000 641.4000 343.8000 641.5500 ;
	    RECT 361.8000 641.4000 363.0000 641.5500 ;
	    RECT 301.8000 638.4000 303.0000 638.5500 ;
	    RECT 306.6000 638.4000 307.8000 638.5500 ;
	    RECT 301.8000 637.2000 303.0000 637.5000 ;
	    RECT 301.8000 633.3000 303.0000 636.3000 ;
	    RECT 321.0000 633.3000 322.2000 639.3000 ;
	    RECT 323.4000 638.4000 326.1000 639.3000 ;
	    RECT 340.2000 638.4000 341.4000 639.6000 ;
	    RECT 324.9000 633.3000 326.1000 638.4000 ;
	    RECT 340.2000 637.2000 341.4000 637.5000 ;
	    RECT 340.2000 633.3000 341.4000 636.3000 ;
	    RECT 342.6000 633.3000 343.8000 640.5000 ;
	    RECT 364.2000 639.3000 365.4000 643.5000 ;
	    RECT 366.6000 642.4500 367.8000 642.6000 ;
	    RECT 450.6000 642.4500 451.8000 642.6000 ;
	    RECT 366.6000 641.5500 451.8000 642.4500 ;
	    RECT 366.6000 641.4000 367.8000 641.5500 ;
	    RECT 450.6000 641.4000 451.8000 641.5500 ;
	    RECT 498.6000 642.3000 511.8000 643.5000 ;
	    RECT 512.7000 642.9000 515.7000 644.1000 ;
	    RECT 521.4000 642.9000 526.2000 644.1000 ;
	    RECT 366.6000 640.2000 367.8000 640.5000 ;
	    RECT 362.7000 638.4000 365.4000 639.3000 ;
	    RECT 362.7000 633.3000 363.9000 638.4000 ;
	    RECT 366.6000 633.3000 367.8000 639.3000 ;
	    RECT 498.6000 633.3000 499.8000 642.3000 ;
	    RECT 502.2000 640.2000 506.7000 641.4000 ;
	    RECT 505.5000 639.3000 506.7000 640.2000 ;
	    RECT 514.5000 639.3000 515.7000 642.9000 ;
	    RECT 517.8000 641.4000 519.0000 642.6000 ;
	    RECT 525.6000 641.7000 526.8000 642.0000 ;
	    RECT 520.2000 640.8000 526.8000 641.7000 ;
	    RECT 520.2000 640.5000 521.4000 640.8000 ;
	    RECT 517.8000 640.2000 519.0000 640.5000 ;
	    RECT 529.8000 639.6000 531.0000 643.8000 ;
	    RECT 538.5000 642.9000 544.2000 644.1000 ;
	    RECT 538.5000 641.1000 539.7000 642.9000 ;
	    RECT 545.1000 642.0000 546.0000 645.0000 ;
	    RECT 520.2000 639.3000 521.4000 639.6000 ;
	    RECT 503.4000 633.3000 504.6000 639.3000 ;
	    RECT 505.5000 638.1000 509.4000 639.3000 ;
	    RECT 514.5000 638.4000 521.4000 639.3000 ;
	    RECT 522.6000 638.4000 523.8000 639.6000 ;
	    RECT 524.7000 638.4000 525.0000 639.6000 ;
	    RECT 529.5000 638.4000 531.0000 639.6000 ;
	    RECT 537.0000 640.2000 539.7000 641.1000 ;
	    RECT 544.2000 641.1000 546.0000 642.0000 ;
	    RECT 537.0000 639.3000 538.2000 640.2000 ;
	    RECT 508.2000 633.3000 509.4000 638.1000 ;
	    RECT 534.6000 638.1000 538.2000 639.3000 ;
	    RECT 510.6000 633.3000 511.8000 637.5000 ;
	    RECT 513.0000 633.3000 514.2000 637.5000 ;
	    RECT 515.4000 633.3000 516.6000 637.5000 ;
	    RECT 517.8000 633.3000 519.0000 636.3000 ;
	    RECT 520.2000 633.3000 521.4000 637.5000 ;
	    RECT 522.6000 633.3000 523.8000 636.3000 ;
	    RECT 525.0000 633.3000 526.2000 637.5000 ;
	    RECT 527.4000 633.3000 528.6000 637.5000 ;
	    RECT 529.8000 633.3000 531.0000 637.5000 ;
	    RECT 532.2000 633.3000 533.4000 637.5000 ;
	    RECT 534.6000 633.3000 535.8000 638.1000 ;
	    RECT 539.4000 633.3000 540.6000 639.3000 ;
	    RECT 544.2000 633.3000 545.4000 641.1000 ;
	    RECT 546.9000 640.2000 548.1000 646.8000 ;
	    RECT 565.8000 643.5000 567.0000 659.7000 ;
	    RECT 593.1000 653.7000 594.3000 659.7000 ;
	    RECT 593.4000 650.4000 594.6000 651.6000 ;
	    RECT 593.4000 649.5000 594.3000 650.4000 ;
	    RECT 595.5000 648.6000 596.7000 659.7000 ;
	    RECT 592.2000 647.4000 593.4000 648.6000 ;
	    RECT 595.2000 647.7000 596.7000 648.6000 ;
	    RECT 599.4000 647.7000 600.6000 659.7000 ;
	    RECT 601.8000 659.4000 603.0000 660.6000 ;
	    RECT 595.2000 642.6000 596.1000 647.7000 ;
	    RECT 597.0000 645.4500 598.2000 645.6000 ;
	    RECT 597.0000 644.5500 602.8500 645.4500 ;
	    RECT 597.0000 644.4000 598.2000 644.5500 ;
	    RECT 597.0000 643.2000 598.2000 643.5000 ;
	    RECT 565.8000 642.4500 567.0000 642.6000 ;
	    RECT 589.8000 642.4500 591.0000 642.6000 ;
	    RECT 565.8000 641.5500 591.0000 642.4500 ;
	    RECT 565.8000 641.4000 567.0000 641.5500 ;
	    RECT 589.8000 641.4000 591.0000 641.5500 ;
	    RECT 592.2000 641.4000 593.4000 642.6000 ;
	    RECT 594.3000 641.4000 596.1000 642.6000 ;
	    RECT 598.2000 640.8000 598.5000 642.3000 ;
	    RECT 599.4000 641.4000 600.6000 642.6000 ;
	    RECT 601.9500 642.4500 602.8500 644.5500 ;
	    RECT 611.4000 643.5000 612.6000 659.7000 ;
	    RECT 613.8000 653.7000 615.0000 659.7000 ;
	    RECT 628.2000 653.7000 629.4000 659.7000 ;
	    RECT 630.6000 643.5000 631.8000 659.7000 ;
	    RECT 657.0000 653.7000 658.2000 659.7000 ;
	    RECT 659.4000 653.7000 660.6000 659.7000 ;
	    RECT 661.8000 654.3000 663.0000 659.7000 ;
	    RECT 659.7000 653.4000 660.6000 653.7000 ;
	    RECT 664.2000 653.7000 665.4000 659.7000 ;
	    RECT 673.8000 659.4000 675.0000 660.6000 ;
	    RECT 676.2000 657.4500 677.4000 657.6000 ;
	    RECT 695.4000 657.4500 696.6000 657.6000 ;
	    RECT 676.2000 656.5500 696.6000 657.4500 ;
	    RECT 676.2000 656.4000 677.4000 656.5500 ;
	    RECT 695.4000 656.4000 696.6000 656.5500 ;
	    RECT 664.2000 653.4000 665.1000 653.7000 ;
	    RECT 659.7000 652.5000 665.1000 653.4000 ;
	    RECT 647.4000 651.4500 648.6000 651.6000 ;
	    RECT 657.0000 651.4500 658.2000 651.6000 ;
	    RECT 647.4000 650.5500 658.2000 651.4500 ;
	    RECT 647.4000 650.4000 648.6000 650.5500 ;
	    RECT 657.0000 650.4000 658.2000 650.5500 ;
	    RECT 661.8000 650.4000 663.0000 651.6000 ;
	    RECT 664.2000 649.5000 665.1000 652.5000 ;
	    RECT 661.8000 649.2000 663.0000 649.5000 ;
	    RECT 657.0000 648.4500 658.2000 648.6000 ;
	    RECT 659.4000 648.4500 660.6000 648.6000 ;
	    RECT 657.0000 647.5500 660.6000 648.4500 ;
	    RECT 657.0000 647.4000 658.2000 647.5500 ;
	    RECT 659.4000 647.4000 660.6000 647.5500 ;
	    RECT 664.2000 648.4500 665.4000 648.6000 ;
	    RECT 697.8000 648.4500 699.0000 648.6000 ;
	    RECT 664.2000 647.5500 699.0000 648.4500 ;
	    RECT 700.2000 647.7000 701.4000 659.7000 ;
	    RECT 704.1000 647.7000 707.1000 659.7000 ;
	    RECT 709.8000 647.7000 711.0000 659.7000 ;
	    RECT 717.0000 654.4500 718.2000 654.6000 ;
	    RECT 762.6000 654.4500 763.8000 654.6000 ;
	    RECT 717.0000 653.5500 763.8000 654.4500 ;
	    RECT 717.0000 653.4000 718.2000 653.5500 ;
	    RECT 762.6000 653.4000 763.8000 653.5500 ;
	    RECT 765.0000 647.7000 766.2000 659.7000 ;
	    RECT 664.2000 647.4000 665.4000 647.5500 ;
	    RECT 697.8000 647.4000 699.0000 647.5500 ;
	    RECT 657.0000 646.2000 658.2000 646.5000 ;
	    RECT 659.4000 644.4000 660.6000 645.6000 ;
	    RECT 661.5000 644.4000 661.8000 645.6000 ;
	    RECT 664.2000 642.6000 665.1000 646.5000 ;
	    RECT 702.6000 644.4000 703.8000 645.6000 ;
	    RECT 700.2000 643.5000 701.4000 643.8000 ;
	    RECT 705.3000 643.5000 706.2000 647.7000 ;
	    RECT 767.4000 646.8000 768.6000 659.7000 ;
	    RECT 769.8000 647.7000 771.0000 659.7000 ;
	    RECT 772.2000 646.8000 773.4000 659.7000 ;
	    RECT 774.6000 647.7000 775.8000 659.7000 ;
	    RECT 777.0000 646.8000 778.2000 659.7000 ;
	    RECT 779.4000 647.7000 780.6000 659.7000 ;
	    RECT 781.8000 646.8000 783.0000 659.7000 ;
	    RECT 784.2000 647.7000 785.4000 659.7000 ;
	    RECT 813.0000 647.7000 814.2000 659.7000 ;
	    RECT 816.9000 647.7000 819.9000 659.7000 ;
	    RECT 822.6000 647.7000 823.8000 659.7000 ;
	    RECT 837.0000 653.7000 838.2000 659.7000 ;
	    RECT 765.0000 646.5000 768.6000 646.8000 ;
	    RECT 767.1000 645.6000 768.6000 646.5000 ;
	    RECT 770.1000 645.6000 773.4000 646.8000 ;
	    RECT 774.9000 645.6000 778.2000 646.8000 ;
	    RECT 780.3000 645.6000 783.0000 646.8000 ;
	    RECT 707.4000 644.4000 708.6000 645.6000 ;
	    RECT 709.8000 645.4500 711.0000 645.6000 ;
	    RECT 755.4000 645.4500 756.6000 645.6000 ;
	    RECT 709.8000 644.5500 756.6000 645.4500 ;
	    RECT 709.8000 644.4000 711.0000 644.5500 ;
	    RECT 755.4000 644.4000 756.6000 644.5500 ;
	    RECT 760.2000 645.4500 761.4000 645.6000 ;
	    RECT 765.0000 645.4500 766.2000 645.6000 ;
	    RECT 760.2000 644.5500 766.2000 645.4500 ;
	    RECT 760.2000 644.4000 761.4000 644.5500 ;
	    RECT 765.0000 644.4000 766.2000 644.5500 ;
	    RECT 770.1000 643.5000 771.3000 645.6000 ;
	    RECT 774.9000 643.5000 776.1000 645.6000 ;
	    RECT 780.3000 643.5000 781.5000 645.6000 ;
	    RECT 815.4000 644.4000 816.6000 645.6000 ;
	    RECT 813.0000 643.5000 814.2000 643.8000 ;
	    RECT 818.1000 643.5000 819.0000 647.7000 ;
	    RECT 820.2000 644.4000 821.4000 645.6000 ;
	    RECT 839.4000 643.5000 840.6000 659.7000 ;
	    RECT 882.6000 657.4500 883.8000 657.6000 ;
	    RECT 966.6000 657.4500 967.8000 657.6000 ;
	    RECT 882.6000 656.5500 967.8000 657.4500 ;
	    RECT 882.6000 656.4000 883.8000 656.5500 ;
	    RECT 966.6000 656.4000 967.8000 656.5500 ;
	    RECT 868.2000 654.4500 869.4000 654.6000 ;
	    RECT 961.8000 654.4500 963.0000 654.6000 ;
	    RECT 868.2000 653.5500 963.0000 654.4500 ;
	    RECT 971.4000 653.7000 972.6000 659.7000 ;
	    RECT 973.8000 654.6000 975.0000 659.7000 ;
	    RECT 973.5000 653.7000 975.0000 654.6000 ;
	    RECT 976.2000 653.7000 977.4000 660.6000 ;
	    RECT 868.2000 653.4000 869.4000 653.5500 ;
	    RECT 961.8000 653.4000 963.0000 653.5500 ;
	    RECT 973.5000 652.8000 974.4000 653.7000 ;
	    RECT 978.6000 652.8000 979.8000 659.7000 ;
	    RECT 981.0000 653.7000 982.2000 659.7000 ;
	    RECT 983.4000 655.5000 984.6000 659.7000 ;
	    RECT 985.8000 655.5000 987.0000 659.7000 ;
	    RECT 971.4000 651.9000 974.4000 652.8000 ;
	    RECT 971.4000 643.5000 972.6000 651.9000 ;
	    RECT 975.3000 651.6000 981.6000 652.8000 ;
	    RECT 988.2000 652.5000 989.4000 659.7000 ;
	    RECT 990.6000 653.7000 991.8000 659.7000 ;
	    RECT 993.0000 652.5000 994.2000 659.7000 ;
	    RECT 995.4000 653.7000 996.6000 659.7000 ;
	    RECT 975.3000 651.0000 976.2000 651.6000 ;
	    RECT 973.8000 649.8000 976.2000 651.0000 ;
	    RECT 980.7000 650.7000 989.4000 651.6000 ;
	    RECT 977.7000 649.8000 979.8000 650.7000 ;
	    RECT 977.7000 649.5000 987.0000 649.8000 ;
	    RECT 978.9000 648.9000 987.0000 649.5000 ;
	    RECT 985.8000 648.6000 987.0000 648.9000 ;
	    RECT 988.5000 649.5000 989.4000 650.7000 ;
	    RECT 990.3000 650.4000 994.2000 651.6000 ;
	    RECT 997.8000 650.4000 999.0000 659.7000 ;
	    RECT 1000.2000 655.5000 1001.4000 659.7000 ;
	    RECT 1002.6000 655.5000 1003.8000 659.7000 ;
	    RECT 1005.0000 655.5000 1006.2000 659.7000 ;
	    RECT 1007.4000 653.7000 1008.6000 659.7000 ;
	    RECT 1002.6000 651.6000 1008.9000 652.8000 ;
	    RECT 1009.8000 651.6000 1011.0000 659.7000 ;
	    RECT 1012.2000 653.7000 1013.4000 659.7000 ;
	    RECT 1014.6000 652.8000 1015.8000 659.7000 ;
	    RECT 1017.0000 653.7000 1018.2000 659.7000 ;
	    RECT 1014.6000 651.9000 1018.5000 652.8000 ;
	    RECT 1019.4000 652.5000 1020.6000 659.7000 ;
	    RECT 1021.8000 653.7000 1023.0000 659.7000 ;
	    RECT 1036.2001 653.7000 1037.4000 659.7000 ;
	    RECT 1009.8000 650.4000 1013.7000 651.6000 ;
	    RECT 1000.2000 649.5000 1001.4000 649.8000 ;
	    RECT 988.5000 648.6000 1001.4000 649.5000 ;
	    RECT 1005.0000 649.5000 1006.2000 649.8000 ;
	    RECT 1017.6000 649.5000 1018.5000 651.9000 ;
	    RECT 1019.4000 650.4000 1020.6000 651.6000 ;
	    RECT 1005.0000 648.6000 1018.5000 649.5000 ;
	    RECT 976.2000 647.4000 977.4000 648.6000 ;
	    RECT 981.3000 647.7000 982.5000 648.0000 ;
	    RECT 978.3000 646.8000 1016.7000 647.7000 ;
	    RECT 1015.5000 646.5000 1016.7000 646.8000 ;
	    RECT 1017.6000 645.9000 1018.5000 648.6000 ;
	    RECT 1019.4000 648.0000 1020.6000 649.5000 ;
	    RECT 1019.4000 646.8000 1020.9000 648.0000 ;
	    RECT 973.5000 645.0000 980.1000 645.9000 ;
	    RECT 973.5000 644.7000 974.7000 645.0000 ;
	    RECT 981.0000 644.4000 982.2000 645.6000 ;
	    RECT 983.1000 645.0000 1008.6000 645.9000 ;
	    RECT 1017.6000 645.0000 1018.8000 645.9000 ;
	    RECT 1007.4000 644.1000 1008.6000 645.0000 ;
	    RECT 702.6000 643.2000 703.8000 643.5000 ;
	    RECT 707.4000 643.2000 708.6000 643.5000 ;
	    RECT 611.4000 642.4500 612.6000 642.6000 ;
	    RECT 601.9500 641.5500 612.6000 642.4500 ;
	    RECT 611.4000 641.4000 612.6000 641.5500 ;
	    RECT 630.6000 642.4500 631.8000 642.6000 ;
	    RECT 649.8000 642.4500 651.0000 642.6000 ;
	    RECT 630.6000 641.5500 651.0000 642.4500 ;
	    RECT 662.7000 642.3000 665.1000 642.6000 ;
	    RECT 630.6000 641.4000 631.8000 641.5500 ;
	    RECT 649.8000 641.4000 651.0000 641.5500 ;
	    RECT 546.6000 639.0000 548.1000 640.2000 ;
	    RECT 546.6000 633.3000 547.8000 639.0000 ;
	    RECT 563.4000 638.4000 564.6000 639.6000 ;
	    RECT 563.4000 637.2000 564.6000 637.5000 ;
	    RECT 549.0000 633.3000 550.2000 636.3000 ;
	    RECT 563.4000 633.3000 564.6000 636.3000 ;
	    RECT 565.8000 633.3000 567.0000 640.5000 ;
	    RECT 592.5000 639.3000 593.4000 640.5000 ;
	    RECT 594.9000 639.3000 600.3000 639.9000 ;
	    RECT 592.2000 633.3000 593.4000 639.3000 ;
	    RECT 594.6000 639.0000 600.6000 639.3000 ;
	    RECT 594.6000 633.3000 595.8000 639.0000 ;
	    RECT 597.0000 633.3000 598.2000 638.1000 ;
	    RECT 599.4000 633.3000 600.6000 639.0000 ;
	    RECT 611.4000 633.3000 612.6000 640.5000 ;
	    RECT 613.8000 639.4500 615.0000 639.6000 ;
	    RECT 628.2000 639.4500 629.4000 639.6000 ;
	    RECT 613.8000 638.5500 629.4000 639.4500 ;
	    RECT 613.8000 638.4000 615.0000 638.5500 ;
	    RECT 628.2000 638.4000 629.4000 638.5500 ;
	    RECT 613.8000 637.2000 615.0000 637.5000 ;
	    RECT 628.2000 637.2000 629.4000 637.5000 ;
	    RECT 613.8000 633.3000 615.0000 636.3000 ;
	    RECT 628.2000 633.3000 629.4000 636.3000 ;
	    RECT 630.6000 633.3000 631.8000 640.5000 ;
	    RECT 657.0000 633.3000 658.2000 642.3000 ;
	    RECT 662.4000 641.7000 665.1000 642.3000 ;
	    RECT 685.8000 642.4500 687.0000 642.6000 ;
	    RECT 700.2000 642.4500 701.4000 642.6000 ;
	    RECT 662.4000 633.3000 663.6000 641.7000 ;
	    RECT 685.8000 641.5500 701.4000 642.4500 ;
	    RECT 685.8000 641.4000 687.0000 641.5500 ;
	    RECT 700.2000 641.4000 701.4000 641.5500 ;
	    RECT 702.6000 641.4000 704.1000 642.3000 ;
	    RECT 705.0000 641.4000 706.2000 642.6000 ;
	    RECT 709.8000 642.4500 711.0000 642.6000 ;
	    RECT 712.2000 642.4500 713.4000 642.6000 ;
	    RECT 702.6000 639.3000 703.5000 641.4000 ;
	    RECT 708.6000 640.8000 708.9000 642.3000 ;
	    RECT 709.8000 641.5500 713.4000 642.4500 ;
	    RECT 709.8000 641.4000 711.0000 641.5500 ;
	    RECT 712.2000 641.4000 713.4000 641.5500 ;
	    RECT 714.6000 642.4500 715.8000 642.6000 ;
	    RECT 760.2000 642.4500 761.4000 642.6000 ;
	    RECT 714.6000 641.5500 761.4000 642.4500 ;
	    RECT 714.6000 641.4000 715.8000 641.5500 ;
	    RECT 760.2000 641.4000 761.4000 641.5500 ;
	    RECT 765.0000 641.4000 766.2000 643.5000 ;
	    RECT 767.4000 642.3000 771.3000 643.5000 ;
	    RECT 772.5000 642.3000 776.1000 643.5000 ;
	    RECT 777.6000 642.3000 781.5000 643.5000 ;
	    RECT 782.7000 642.3000 783.3000 643.5000 ;
	    RECT 815.4000 643.2000 816.6000 643.5000 ;
	    RECT 820.2000 643.2000 821.4000 643.5000 ;
	    RECT 770.1000 641.4000 771.3000 642.3000 ;
	    RECT 774.9000 641.4000 776.1000 642.3000 ;
	    RECT 780.3000 641.4000 781.5000 642.3000 ;
	    RECT 784.2000 641.4000 785.4000 642.6000 ;
	    RECT 786.6000 642.4500 787.8000 642.6000 ;
	    RECT 813.0000 642.4500 814.2000 642.6000 ;
	    RECT 786.6000 641.5500 814.2000 642.4500 ;
	    RECT 786.6000 641.4000 787.8000 641.5500 ;
	    RECT 813.0000 641.4000 814.2000 641.5500 ;
	    RECT 815.4000 641.4000 816.9000 642.3000 ;
	    RECT 817.8000 641.4000 819.0000 642.6000 ;
	    RECT 765.0000 640.2000 768.6000 641.4000 ;
	    RECT 770.1000 640.2000 773.4000 641.4000 ;
	    RECT 774.9000 640.2000 778.2000 641.4000 ;
	    RECT 780.3000 640.2000 783.0000 641.4000 ;
	    RECT 705.3000 639.3000 710.7000 639.9000 ;
	    RECT 700.2000 634.2000 701.4000 639.3000 ;
	    RECT 702.6000 635.1000 703.8000 639.3000 ;
	    RECT 705.0000 639.0000 711.0000 639.3000 ;
	    RECT 705.0000 634.2000 706.2000 639.0000 ;
	    RECT 700.2000 633.3000 706.2000 634.2000 ;
	    RECT 707.4000 633.3000 708.6000 638.1000 ;
	    RECT 709.8000 633.3000 711.0000 639.0000 ;
	    RECT 753.0000 636.4500 754.2000 636.6000 ;
	    RECT 762.6000 636.4500 763.8000 636.6000 ;
	    RECT 753.0000 635.5500 763.8000 636.4500 ;
	    RECT 753.0000 635.4000 754.2000 635.5500 ;
	    RECT 762.6000 635.4000 763.8000 635.5500 ;
	    RECT 765.0000 633.3000 766.2000 639.3000 ;
	    RECT 767.4000 633.3000 768.6000 640.2000 ;
	    RECT 769.8000 633.3000 771.0000 639.3000 ;
	    RECT 772.2000 633.3000 773.4000 640.2000 ;
	    RECT 774.6000 633.3000 775.8000 639.3000 ;
	    RECT 777.0000 633.3000 778.2000 640.2000 ;
	    RECT 779.4000 633.3000 780.6000 639.3000 ;
	    RECT 781.8000 633.3000 783.0000 640.2000 ;
	    RECT 815.4000 639.3000 816.3000 641.4000 ;
	    RECT 821.4000 640.8000 821.7000 642.3000 ;
	    RECT 822.6000 641.4000 823.8000 642.6000 ;
	    RECT 839.4000 642.4500 840.6000 642.6000 ;
	    RECT 942.6000 642.4500 943.8000 642.6000 ;
	    RECT 839.4000 641.5500 943.8000 642.4500 ;
	    RECT 839.4000 641.4000 840.6000 641.5500 ;
	    RECT 942.6000 641.4000 943.8000 641.5500 ;
	    RECT 971.4000 642.3000 984.6000 643.5000 ;
	    RECT 985.5000 642.9000 988.5000 644.1000 ;
	    RECT 994.2000 642.9000 999.0000 644.1000 ;
	    RECT 818.1000 639.3000 823.5000 639.9000 ;
	    RECT 832.2000 639.4500 833.4000 639.6000 ;
	    RECT 837.0000 639.4500 838.2000 639.6000 ;
	    RECT 784.2000 633.3000 785.4000 639.3000 ;
	    RECT 813.0000 634.2000 814.2000 639.3000 ;
	    RECT 815.4000 635.1000 816.6000 639.3000 ;
	    RECT 817.8000 639.0000 823.8000 639.3000 ;
	    RECT 817.8000 634.2000 819.0000 639.0000 ;
	    RECT 813.0000 633.3000 819.0000 634.2000 ;
	    RECT 820.2000 633.3000 821.4000 638.1000 ;
	    RECT 822.6000 633.3000 823.8000 639.0000 ;
	    RECT 832.2000 638.5500 838.2000 639.4500 ;
	    RECT 832.2000 638.4000 833.4000 638.5500 ;
	    RECT 837.0000 638.4000 838.2000 638.5500 ;
	    RECT 837.0000 637.2000 838.2000 637.5000 ;
	    RECT 837.0000 633.3000 838.2000 636.3000 ;
	    RECT 839.4000 633.3000 840.6000 640.5000 ;
	    RECT 849.0000 639.4500 850.2000 639.6000 ;
	    RECT 942.6000 639.4500 943.8000 639.6000 ;
	    RECT 849.0000 638.5500 943.8000 639.4500 ;
	    RECT 849.0000 638.4000 850.2000 638.5500 ;
	    RECT 942.6000 638.4000 943.8000 638.5500 ;
	    RECT 971.4000 633.3000 972.6000 642.3000 ;
	    RECT 975.0000 640.2000 979.5000 641.4000 ;
	    RECT 978.3000 639.3000 979.5000 640.2000 ;
	    RECT 987.3000 639.3000 988.5000 642.9000 ;
	    RECT 990.6000 641.4000 991.8000 642.6000 ;
	    RECT 998.4000 641.7000 999.6000 642.0000 ;
	    RECT 993.0000 640.8000 999.6000 641.7000 ;
	    RECT 993.0000 640.5000 994.2000 640.8000 ;
	    RECT 990.6000 640.2000 991.8000 640.5000 ;
	    RECT 1002.6000 639.6000 1003.8000 643.8000 ;
	    RECT 1011.3000 642.9000 1017.0000 644.1000 ;
	    RECT 1011.3000 641.1000 1012.5000 642.9000 ;
	    RECT 1017.9000 642.0000 1018.8000 645.0000 ;
	    RECT 993.0000 639.3000 994.2000 639.6000 ;
	    RECT 976.2000 633.3000 977.4000 639.3000 ;
	    RECT 978.3000 638.1000 982.2000 639.3000 ;
	    RECT 987.3000 638.4000 994.2000 639.3000 ;
	    RECT 995.4000 638.4000 996.6000 639.6000 ;
	    RECT 997.5000 638.4000 997.8000 639.6000 ;
	    RECT 1002.3000 638.4000 1003.8000 639.6000 ;
	    RECT 1009.8000 640.2000 1012.5000 641.1000 ;
	    RECT 1017.0000 641.1000 1018.8000 642.0000 ;
	    RECT 1009.8000 639.3000 1011.0000 640.2000 ;
	    RECT 981.0000 633.3000 982.2000 638.1000 ;
	    RECT 1007.4000 638.1000 1011.0000 639.3000 ;
	    RECT 983.4000 633.3000 984.6000 637.5000 ;
	    RECT 985.8000 633.3000 987.0000 637.5000 ;
	    RECT 988.2000 633.3000 989.4000 637.5000 ;
	    RECT 990.6000 633.3000 991.8000 636.3000 ;
	    RECT 993.0000 633.3000 994.2000 637.5000 ;
	    RECT 995.4000 633.3000 996.6000 636.3000 ;
	    RECT 997.8000 633.3000 999.0000 637.5000 ;
	    RECT 1000.2000 633.3000 1001.4000 637.5000 ;
	    RECT 1002.6000 633.3000 1003.8000 637.5000 ;
	    RECT 1005.0000 633.3000 1006.2000 637.5000 ;
	    RECT 1007.4000 633.3000 1008.6000 638.1000 ;
	    RECT 1012.2000 633.3000 1013.4000 639.3000 ;
	    RECT 1017.0000 633.3000 1018.2000 641.1000 ;
	    RECT 1019.7000 640.2000 1020.9000 646.8000 ;
	    RECT 1038.6000 643.5000 1039.8000 659.7000 ;
	    RECT 1062.6000 647.7000 1063.8000 659.7000 ;
	    RECT 1066.5000 648.6000 1067.7001 659.7000 ;
	    RECT 1068.9000 653.7000 1070.1000 659.7000 ;
	    RECT 1081.8000 653.7000 1083.0000 659.7000 ;
	    RECT 1068.6000 650.4000 1069.8000 651.6000 ;
	    RECT 1068.9000 649.5000 1069.8000 650.4000 ;
	    RECT 1066.5000 647.7000 1068.0000 648.6000 ;
	    RECT 1065.0000 645.4500 1066.2001 645.6000 ;
	    RECT 1055.5500 644.5500 1066.2001 645.4500 ;
	    RECT 1038.6000 642.4500 1039.8000 642.6000 ;
	    RECT 1055.5500 642.4500 1056.4501 644.5500 ;
	    RECT 1065.0000 644.4000 1066.2001 644.5500 ;
	    RECT 1065.0000 643.2000 1066.2001 643.5000 ;
	    RECT 1067.1000 642.6000 1068.0000 647.7000 ;
	    RECT 1069.8000 647.4000 1071.0000 648.6000 ;
	    RECT 1084.2001 643.5000 1085.4000 659.7000 ;
	    RECT 1110.6000 647.7000 1111.8000 659.7000 ;
	    RECT 1114.5000 648.6000 1115.7001 659.7000 ;
	    RECT 1116.9000 653.7000 1118.1000 659.7000 ;
	    RECT 1116.6000 650.4000 1117.8000 651.6000 ;
	    RECT 1116.9000 649.5000 1117.8000 650.4000 ;
	    RECT 1114.5000 647.7000 1116.0000 648.6000 ;
	    RECT 1113.0000 645.4500 1114.2001 645.6000 ;
	    RECT 1108.3500 644.5500 1114.2001 645.4500 ;
	    RECT 1038.6000 641.5500 1056.4501 642.4500 ;
	    RECT 1057.8000 642.4500 1059.0000 642.6000 ;
	    RECT 1062.6000 642.4500 1063.8000 642.6000 ;
	    RECT 1057.8000 641.5500 1063.8000 642.4500 ;
	    RECT 1038.6000 641.4000 1039.8000 641.5500 ;
	    RECT 1057.8000 641.4000 1059.0000 641.5500 ;
	    RECT 1062.6000 641.4000 1063.8000 641.5500 ;
	    RECT 1064.7001 640.8000 1065.0000 642.3000 ;
	    RECT 1067.1000 641.4000 1068.9000 642.6000 ;
	    RECT 1069.8000 642.4500 1071.0000 642.6000 ;
	    RECT 1081.8000 642.4500 1083.0000 642.6000 ;
	    RECT 1069.8000 641.5500 1083.0000 642.4500 ;
	    RECT 1069.8000 641.4000 1071.0000 641.5500 ;
	    RECT 1081.8000 641.4000 1083.0000 641.5500 ;
	    RECT 1084.2001 642.4500 1085.4000 642.6000 ;
	    RECT 1108.3500 642.4500 1109.2500 644.5500 ;
	    RECT 1113.0000 644.4000 1114.2001 644.5500 ;
	    RECT 1113.0000 643.2000 1114.2001 643.5000 ;
	    RECT 1115.1000 642.6000 1116.0000 647.7000 ;
	    RECT 1117.8000 648.4500 1119.0000 648.6000 ;
	    RECT 1134.6000 648.4500 1135.8000 648.6000 ;
	    RECT 1117.8000 647.5500 1135.8000 648.4500 ;
	    RECT 1177.8000 647.7000 1179.0000 659.7000 ;
	    RECT 1117.8000 647.4000 1119.0000 647.5500 ;
	    RECT 1134.6000 647.4000 1135.8000 647.5500 ;
	    RECT 1180.2001 646.8000 1181.4000 659.7000 ;
	    RECT 1182.6000 647.7000 1183.8000 659.7000 ;
	    RECT 1185.0000 646.8000 1186.2001 659.7000 ;
	    RECT 1187.4000 647.7000 1188.6000 659.7000 ;
	    RECT 1189.8000 646.8000 1191.0000 659.7000 ;
	    RECT 1192.2001 647.7000 1193.4000 659.7000 ;
	    RECT 1194.6000 646.8000 1195.8000 659.7000 ;
	    RECT 1197.0000 647.7000 1198.2001 659.7000 ;
	    RECT 1217.1000 648.9000 1218.3000 659.7000 ;
	    RECT 1217.1000 647.7000 1219.8000 648.9000 ;
	    RECT 1221.0000 647.7000 1222.2001 659.7000 ;
	    RECT 1245.9000 653.7000 1247.1000 659.7000 ;
	    RECT 1246.2001 650.4000 1247.4000 651.6000 ;
	    RECT 1246.2001 649.5000 1247.1000 650.4000 ;
	    RECT 1248.3000 648.6000 1249.5000 659.7000 ;
	    RECT 1228.2001 648.4500 1229.4000 648.6000 ;
	    RECT 1245.0000 648.4500 1246.2001 648.6000 ;
	    RECT 1180.2001 645.6000 1182.9000 646.8000 ;
	    RECT 1185.0000 645.6000 1188.3000 646.8000 ;
	    RECT 1189.8000 645.6000 1193.1000 646.8000 ;
	    RECT 1194.6000 646.5000 1198.2001 646.8000 ;
	    RECT 1216.2001 646.5000 1217.4000 646.8000 ;
	    RECT 1194.6000 645.6000 1196.1000 646.5000 ;
	    RECT 1181.7001 643.5000 1182.9000 645.6000 ;
	    RECT 1187.1000 643.5000 1188.3000 645.6000 ;
	    RECT 1191.9000 643.5000 1193.1000 645.6000 ;
	    RECT 1197.0000 644.4000 1198.2001 645.6000 ;
	    RECT 1216.2001 644.4000 1217.4000 645.6000 ;
	    RECT 1218.6000 643.5000 1219.5000 647.7000 ;
	    RECT 1228.2001 647.5500 1246.2001 648.4500 ;
	    RECT 1228.2001 647.4000 1229.4000 647.5500 ;
	    RECT 1245.0000 647.4000 1246.2001 647.5500 ;
	    RECT 1248.0000 647.7000 1249.5000 648.6000 ;
	    RECT 1252.2001 647.7000 1253.4000 659.7000 ;
	    RECT 1271.4000 653.7000 1272.6000 659.7000 ;
	    RECT 1084.2001 641.5500 1109.2500 642.4500 ;
	    RECT 1084.2001 641.4000 1085.4000 641.5500 ;
	    RECT 1110.6000 641.4000 1111.8000 642.6000 ;
	    RECT 1112.7001 640.8000 1113.0000 642.3000 ;
	    RECT 1115.1000 641.4000 1116.9000 642.6000 ;
	    RECT 1117.8000 641.4000 1119.0000 642.6000 ;
	    RECT 1177.8000 641.4000 1179.0000 642.6000 ;
	    RECT 1179.9000 642.3000 1180.5000 643.5000 ;
	    RECT 1181.7001 642.3000 1185.6000 643.5000 ;
	    RECT 1187.1000 642.3000 1190.7001 643.5000 ;
	    RECT 1191.9000 642.3000 1195.8000 643.5000 ;
	    RECT 1181.7001 641.4000 1182.9000 642.3000 ;
	    RECT 1187.1000 641.4000 1188.3000 642.3000 ;
	    RECT 1191.9000 641.4000 1193.1000 642.3000 ;
	    RECT 1197.0000 641.4000 1198.2001 643.5000 ;
	    RECT 1248.0000 642.6000 1248.9000 647.7000 ;
	    RECT 1273.8000 646.5000 1275.0000 659.7000 ;
	    RECT 1276.2001 653.7000 1277.4000 659.7000 ;
	    RECT 1300.2001 653.7000 1301.4000 659.7000 ;
	    RECT 1302.6000 653.7000 1303.8000 659.7000 ;
	    RECT 1305.0000 654.3000 1306.2001 659.7000 ;
	    RECT 1302.9000 653.4000 1303.8000 653.7000 ;
	    RECT 1307.4000 653.7000 1308.6000 659.7000 ;
	    RECT 1321.8000 653.7000 1323.0000 659.7000 ;
	    RECT 1307.4000 653.4000 1308.3000 653.7000 ;
	    RECT 1302.9000 652.5000 1308.3000 653.4000 ;
	    RECT 1305.0000 650.4000 1306.2001 651.6000 ;
	    RECT 1276.2001 649.5000 1277.4000 649.8000 ;
	    RECT 1307.4000 649.5000 1308.3000 652.5000 ;
	    RECT 1305.0000 649.2000 1306.2001 649.5000 ;
	    RECT 1276.2001 647.4000 1277.4000 648.6000 ;
	    RECT 1297.8000 648.4500 1299.0000 648.6000 ;
	    RECT 1300.2001 648.4500 1301.4000 648.6000 ;
	    RECT 1297.8000 647.5500 1301.4000 648.4500 ;
	    RECT 1297.8000 647.4000 1299.0000 647.5500 ;
	    RECT 1300.2001 647.4000 1301.4000 647.5500 ;
	    RECT 1307.4000 648.4500 1308.6000 648.6000 ;
	    RECT 1319.4000 648.4500 1320.6000 648.6000 ;
	    RECT 1307.4000 647.5500 1320.6000 648.4500 ;
	    RECT 1307.4000 647.4000 1308.6000 647.5500 ;
	    RECT 1319.4000 647.4000 1320.6000 647.5500 ;
	    RECT 1300.2001 646.2000 1301.4000 646.5000 ;
	    RECT 1249.8000 644.4000 1251.0000 645.6000 ;
	    RECT 1269.0000 645.4500 1270.2001 645.6000 ;
	    RECT 1273.8000 645.4500 1275.0000 645.6000 ;
	    RECT 1269.0000 644.5500 1275.0000 645.4500 ;
	    RECT 1269.0000 644.4000 1270.2001 644.5500 ;
	    RECT 1273.8000 644.4000 1275.0000 644.5500 ;
	    RECT 1302.6000 644.4000 1303.8000 645.6000 ;
	    RECT 1304.7001 644.4000 1305.0000 645.6000 ;
	    RECT 1249.8000 643.2000 1251.0000 643.5000 ;
	    RECT 1213.8000 642.4500 1215.0000 642.6000 ;
	    RECT 1218.6000 642.4500 1219.8000 642.6000 ;
	    RECT 1237.8000 642.4500 1239.0000 642.6000 ;
	    RECT 1213.8000 641.5500 1239.0000 642.4500 ;
	    RECT 1213.8000 641.4000 1215.0000 641.5500 ;
	    RECT 1218.6000 641.4000 1219.8000 641.5500 ;
	    RECT 1237.8000 641.4000 1239.0000 641.5500 ;
	    RECT 1245.0000 641.4000 1246.2001 642.6000 ;
	    RECT 1247.1000 641.4000 1248.9000 642.6000 ;
	    RECT 1019.4000 639.0000 1020.9000 640.2000 ;
	    RECT 1019.4000 633.3000 1020.6000 639.0000 ;
	    RECT 1036.2001 638.4000 1037.4000 639.6000 ;
	    RECT 1036.2001 637.2000 1037.4000 637.5000 ;
	    RECT 1021.8000 633.3000 1023.0000 636.3000 ;
	    RECT 1036.2001 633.3000 1037.4000 636.3000 ;
	    RECT 1038.6000 633.3000 1039.8000 640.5000 ;
	    RECT 1062.9000 639.3000 1068.3000 639.9000 ;
	    RECT 1069.8000 639.3000 1070.7001 640.5000 ;
	    RECT 1074.6000 639.4500 1075.8000 639.6000 ;
	    RECT 1081.8000 639.4500 1083.0000 639.6000 ;
	    RECT 1062.6000 639.0000 1068.6000 639.3000 ;
	    RECT 1062.6000 633.3000 1063.8000 639.0000 ;
	    RECT 1065.0000 633.3000 1066.2001 638.1000 ;
	    RECT 1067.4000 633.3000 1068.6000 639.0000 ;
	    RECT 1069.8000 633.3000 1071.0000 639.3000 ;
	    RECT 1074.6000 638.5500 1083.0000 639.4500 ;
	    RECT 1074.6000 638.4000 1075.8000 638.5500 ;
	    RECT 1081.8000 638.4000 1083.0000 638.5500 ;
	    RECT 1081.8000 637.2000 1083.0000 637.5000 ;
	    RECT 1081.8000 633.3000 1083.0000 636.3000 ;
	    RECT 1084.2001 633.3000 1085.4000 640.5000 ;
	    RECT 1110.9000 639.3000 1116.3000 639.9000 ;
	    RECT 1117.8000 639.3000 1118.7001 640.5000 ;
	    RECT 1180.2001 640.2000 1182.9000 641.4000 ;
	    RECT 1185.0000 640.2000 1188.3000 641.4000 ;
	    RECT 1189.8000 640.2000 1193.1000 641.4000 ;
	    RECT 1194.6000 640.2000 1198.2001 641.4000 ;
	    RECT 1251.0000 640.8000 1251.3000 642.3000 ;
	    RECT 1252.2001 641.4000 1253.4000 642.6000 ;
	    RECT 1271.4000 641.4000 1272.6000 642.6000 ;
	    RECT 1110.6000 639.0000 1116.6000 639.3000 ;
	    RECT 1110.6000 633.3000 1111.8000 639.0000 ;
	    RECT 1113.0000 633.3000 1114.2001 638.1000 ;
	    RECT 1115.4000 633.3000 1116.6000 639.0000 ;
	    RECT 1117.8000 633.3000 1119.0000 639.3000 ;
	    RECT 1177.8000 633.3000 1179.0000 639.3000 ;
	    RECT 1180.2001 633.3000 1181.4000 640.2000 ;
	    RECT 1182.6000 633.3000 1183.8000 639.3000 ;
	    RECT 1185.0000 633.3000 1186.2001 640.2000 ;
	    RECT 1187.4000 633.3000 1188.6000 639.3000 ;
	    RECT 1189.8000 633.3000 1191.0000 640.2000 ;
	    RECT 1192.2001 633.3000 1193.4000 639.3000 ;
	    RECT 1194.6000 633.3000 1195.8000 640.2000 ;
	    RECT 1197.0000 633.3000 1198.2001 639.3000 ;
	    RECT 1218.6000 636.3000 1219.5000 640.5000 ;
	    RECT 1221.0000 638.4000 1222.2001 639.6000 ;
	    RECT 1245.3000 639.3000 1246.2001 640.5000 ;
	    RECT 1271.4000 640.2000 1272.6000 640.5000 ;
	    RECT 1247.7001 639.3000 1253.1000 639.9000 ;
	    RECT 1273.8000 639.3000 1275.0000 643.5000 ;
	    RECT 1307.4000 642.6000 1308.3000 646.5000 ;
	    RECT 1324.2001 643.5000 1325.4000 659.7000 ;
	    RECT 1348.2001 653.7000 1349.4000 659.7000 ;
	    RECT 1350.6000 653.7000 1351.8000 659.7000 ;
	    RECT 1353.0000 654.3000 1354.2001 659.7000 ;
	    RECT 1350.9000 653.4000 1351.8000 653.7000 ;
	    RECT 1355.4000 653.7000 1356.6000 659.7000 ;
	    RECT 1393.8000 658.8000 1399.8000 659.7000 ;
	    RECT 1355.4000 653.4000 1356.3000 653.7000 ;
	    RECT 1350.9000 652.5000 1356.3000 653.4000 ;
	    RECT 1338.6000 651.4500 1339.8000 651.6000 ;
	    RECT 1353.0000 651.4500 1354.2001 651.6000 ;
	    RECT 1338.6000 650.5500 1354.2001 651.4500 ;
	    RECT 1338.6000 650.4000 1339.8000 650.5500 ;
	    RECT 1353.0000 650.4000 1354.2001 650.5500 ;
	    RECT 1355.4000 649.5000 1356.3000 652.5000 ;
	    RECT 1353.0000 649.2000 1354.2001 649.5000 ;
	    RECT 1348.2001 647.4000 1349.4000 648.6000 ;
	    RECT 1355.4000 648.4500 1356.6000 648.6000 ;
	    RECT 1391.4000 648.4500 1392.6000 648.6000 ;
	    RECT 1355.4000 647.5500 1392.6000 648.4500 ;
	    RECT 1393.8000 647.7000 1395.0000 658.8000 ;
	    RECT 1396.2001 647.7000 1397.4000 657.9000 ;
	    RECT 1398.6000 648.6000 1399.8000 658.8000 ;
	    RECT 1401.0000 649.5000 1402.2001 659.7000 ;
	    RECT 1403.4000 648.6000 1404.6000 659.7000 ;
	    RECT 1398.6000 647.7000 1404.6000 648.6000 ;
	    RECT 1427.4000 647.7000 1428.6000 659.7000 ;
	    RECT 1431.3000 648.6000 1432.5000 659.7000 ;
	    RECT 1433.7001 653.7000 1434.9000 659.7000 ;
	    RECT 1458.6000 653.7000 1459.8000 659.7000 ;
	    RECT 1461.0000 653.7000 1462.2001 659.7000 ;
	    RECT 1463.4000 654.3000 1464.6000 659.7000 ;
	    RECT 1461.3000 653.4000 1462.2001 653.7000 ;
	    RECT 1465.8000 653.7000 1467.0000 659.7000 ;
	    RECT 1465.8000 653.4000 1466.7001 653.7000 ;
	    RECT 1461.3000 652.5000 1466.7001 653.4000 ;
	    RECT 1433.4000 650.4000 1434.6000 651.6000 ;
	    RECT 1463.4000 650.4000 1464.6000 651.6000 ;
	    RECT 1433.7001 649.5000 1434.6000 650.4000 ;
	    RECT 1465.8000 649.5000 1466.7001 652.5000 ;
	    RECT 1463.4000 649.2000 1464.6000 649.5000 ;
	    RECT 1492.2001 648.6000 1493.4000 659.7000 ;
	    RECT 1494.6000 649.5000 1495.8000 659.7000 ;
	    RECT 1497.0000 648.6000 1498.2001 659.7000 ;
	    RECT 1431.3000 647.7000 1432.8000 648.6000 ;
	    RECT 1355.4000 647.4000 1356.6000 647.5500 ;
	    RECT 1391.4000 647.4000 1392.6000 647.5500 ;
	    RECT 1396.5000 646.8000 1397.4000 647.7000 ;
	    RECT 1393.8000 646.5000 1395.0000 646.8000 ;
	    RECT 1396.5000 646.5000 1399.5000 646.8000 ;
	    RECT 1348.2001 646.2000 1349.4000 646.5000 ;
	    RECT 1350.6000 644.4000 1351.8000 645.6000 ;
	    RECT 1352.7001 644.4000 1353.0000 645.6000 ;
	    RECT 1355.4000 642.6000 1356.3000 646.5000 ;
	    RECT 1396.5000 645.9000 1397.7001 646.5000 ;
	    RECT 1381.8000 645.4500 1383.0000 645.6000 ;
	    RECT 1393.8000 645.4500 1395.0000 645.6000 ;
	    RECT 1381.8000 644.5500 1395.0000 645.4500 ;
	    RECT 1381.8000 644.4000 1383.0000 644.5500 ;
	    RECT 1393.8000 644.4000 1395.0000 644.5500 ;
	    RECT 1398.6000 644.4000 1399.8000 645.6000 ;
	    RECT 1402.2001 644.7000 1402.5000 646.2000 ;
	    RECT 1403.4000 644.4000 1404.6000 645.6000 ;
	    RECT 1429.8000 644.4000 1431.0000 645.6000 ;
	    RECT 1396.5000 643.5000 1397.7001 644.4000 ;
	    RECT 1401.0000 643.5000 1402.2001 643.8000 ;
	    RECT 1305.9000 642.3000 1308.3000 642.6000 ;
	    RECT 1221.0000 637.2000 1222.2001 637.5000 ;
	    RECT 1216.2001 633.3000 1217.4000 636.3000 ;
	    RECT 1218.6000 633.3000 1219.8000 636.3000 ;
	    RECT 1221.0000 633.3000 1222.2001 636.3000 ;
	    RECT 1245.0000 633.3000 1246.2001 639.3000 ;
	    RECT 1247.4000 639.0000 1253.4000 639.3000 ;
	    RECT 1247.4000 633.3000 1248.6000 639.0000 ;
	    RECT 1249.8000 633.3000 1251.0000 638.1000 ;
	    RECT 1252.2001 633.3000 1253.4000 639.0000 ;
	    RECT 1271.4000 633.3000 1272.6000 639.3000 ;
	    RECT 1273.8000 638.4000 1276.5000 639.3000 ;
	    RECT 1275.3000 633.3000 1276.5000 638.4000 ;
	    RECT 1300.2001 633.3000 1301.4000 642.3000 ;
	    RECT 1305.6000 641.7000 1308.3000 642.3000 ;
	    RECT 1324.2001 642.4500 1325.4000 642.6000 ;
	    RECT 1345.8000 642.4500 1347.0000 642.6000 ;
	    RECT 1305.6000 633.3000 1306.8000 641.7000 ;
	    RECT 1324.2001 641.5500 1347.0000 642.4500 ;
	    RECT 1353.9000 642.3000 1356.3000 642.6000 ;
	    RECT 1324.2001 641.4000 1325.4000 641.5500 ;
	    RECT 1345.8000 641.4000 1347.0000 641.5500 ;
	    RECT 1319.4000 639.4500 1320.6000 639.6000 ;
	    RECT 1321.8000 639.4500 1323.0000 639.6000 ;
	    RECT 1319.4000 638.5500 1323.0000 639.4500 ;
	    RECT 1319.4000 638.4000 1320.6000 638.5500 ;
	    RECT 1321.8000 638.4000 1323.0000 638.5500 ;
	    RECT 1321.8000 637.2000 1323.0000 637.5000 ;
	    RECT 1321.8000 633.3000 1323.0000 636.3000 ;
	    RECT 1324.2001 633.3000 1325.4000 640.5000 ;
	    RECT 1348.2001 633.3000 1349.4000 642.3000 ;
	    RECT 1353.6000 641.7000 1356.3000 642.3000 ;
	    RECT 1369.8000 642.4500 1371.0000 642.6000 ;
	    RECT 1396.2001 642.4500 1397.4000 642.6000 ;
	    RECT 1353.6000 633.3000 1354.8000 641.7000 ;
	    RECT 1369.8000 641.5500 1397.4000 642.4500 ;
	    RECT 1369.8000 641.4000 1371.0000 641.5500 ;
	    RECT 1396.2001 641.4000 1397.4000 641.5500 ;
	    RECT 1398.6000 639.3000 1399.5000 643.5000 ;
	    RECT 1429.8000 643.2000 1431.0000 643.5000 ;
	    RECT 1431.9000 642.6000 1432.8000 647.7000 ;
	    RECT 1434.6000 648.4500 1435.8000 648.6000 ;
	    RECT 1437.0000 648.4500 1438.2001 648.6000 ;
	    RECT 1434.6000 647.5500 1438.2001 648.4500 ;
	    RECT 1434.6000 647.4000 1435.8000 647.5500 ;
	    RECT 1437.0000 647.4000 1438.2001 647.5500 ;
	    RECT 1449.0000 648.4500 1450.2001 648.6000 ;
	    RECT 1453.8000 648.4500 1455.0000 648.6000 ;
	    RECT 1458.6000 648.4500 1459.8000 648.6000 ;
	    RECT 1449.0000 647.5500 1459.8000 648.4500 ;
	    RECT 1449.0000 647.4000 1450.2001 647.5500 ;
	    RECT 1453.8000 647.4000 1455.0000 647.5500 ;
	    RECT 1458.6000 647.4000 1459.8000 647.5500 ;
	    RECT 1465.8000 648.4500 1467.0000 648.6000 ;
	    RECT 1480.2001 648.4500 1481.4000 648.6000 ;
	    RECT 1465.8000 647.5500 1481.4000 648.4500 ;
	    RECT 1492.2001 647.7000 1498.2001 648.6000 ;
	    RECT 1499.4000 647.7000 1500.6000 659.7000 ;
	    RECT 1523.4000 647.7000 1524.6000 659.7000 ;
	    RECT 1525.8000 648.6000 1527.0000 659.7000 ;
	    RECT 1528.2001 649.5000 1529.4000 659.7000 ;
	    RECT 1530.6000 648.6000 1531.8000 659.7000 ;
	    RECT 1545.0000 653.7000 1546.2001 659.7000 ;
	    RECT 1525.8000 647.7000 1531.8000 648.6000 ;
	    RECT 1465.8000 647.4000 1467.0000 647.5500 ;
	    RECT 1480.2001 647.4000 1481.4000 647.5500 ;
	    RECT 1499.4000 646.5000 1500.3000 647.7000 ;
	    RECT 1523.7001 646.5000 1524.6000 647.7000 ;
	    RECT 1458.6000 646.2000 1459.8000 646.5000 ;
	    RECT 1461.0000 644.4000 1462.2001 645.6000 ;
	    RECT 1463.1000 644.4000 1463.4000 645.6000 ;
	    RECT 1465.8000 642.6000 1466.7001 646.5000 ;
	    RECT 1492.2001 644.4000 1493.4000 645.6000 ;
	    RECT 1494.3000 644.7000 1494.6000 646.2000 ;
	    RECT 1497.0000 644.7000 1498.5000 645.6000 ;
	    RECT 1499.4000 645.4500 1500.6000 645.6000 ;
	    RECT 1501.8000 645.4500 1503.0000 645.6000 ;
	    RECT 1494.6000 643.5000 1495.8000 643.8000 ;
	    RECT 1401.0000 642.4500 1402.2001 642.6000 ;
	    RECT 1408.2001 642.4500 1409.4000 642.6000 ;
	    RECT 1401.0000 641.5500 1409.4000 642.4500 ;
	    RECT 1401.0000 641.4000 1402.2001 641.5500 ;
	    RECT 1408.2001 641.4000 1409.4000 641.5500 ;
	    RECT 1420.2001 642.4500 1421.4000 642.6000 ;
	    RECT 1427.4000 642.4500 1428.6000 642.6000 ;
	    RECT 1420.2001 641.5500 1428.6000 642.4500 ;
	    RECT 1420.2001 641.4000 1421.4000 641.5500 ;
	    RECT 1427.4000 641.4000 1428.6000 641.5500 ;
	    RECT 1429.5000 640.8000 1429.8000 642.3000 ;
	    RECT 1431.9000 641.4000 1433.7001 642.6000 ;
	    RECT 1434.6000 642.4500 1435.8000 642.6000 ;
	    RECT 1444.2001 642.4500 1445.4000 642.6000 ;
	    RECT 1434.6000 641.5500 1445.4000 642.4500 ;
	    RECT 1464.3000 642.3000 1466.7001 642.6000 ;
	    RECT 1434.6000 641.4000 1435.8000 641.5500 ;
	    RECT 1444.2001 641.4000 1445.4000 641.5500 ;
	    RECT 1427.7001 639.3000 1433.1000 639.9000 ;
	    RECT 1434.6000 639.3000 1435.5000 640.5000 ;
	    RECT 1393.8000 633.3000 1395.0000 639.3000 ;
	    RECT 1397.7001 633.3000 1400.1000 639.3000 ;
	    RECT 1402.8000 633.3000 1404.0000 639.3000 ;
	    RECT 1427.4000 639.0000 1433.4000 639.3000 ;
	    RECT 1427.4000 633.3000 1428.6000 639.0000 ;
	    RECT 1429.8000 633.3000 1431.0000 638.1000 ;
	    RECT 1432.2001 633.3000 1433.4000 639.0000 ;
	    RECT 1434.6000 633.3000 1435.8000 639.3000 ;
	    RECT 1458.6000 633.3000 1459.8000 642.3000 ;
	    RECT 1464.0000 641.7000 1466.7001 642.3000 ;
	    RECT 1464.0000 633.3000 1465.2001 641.7000 ;
	    RECT 1494.6000 641.4000 1495.8000 642.6000 ;
	    RECT 1497.0000 639.3000 1497.9000 644.7000 ;
	    RECT 1499.4000 644.5500 1503.0000 645.4500 ;
	    RECT 1499.4000 644.4000 1500.6000 644.5500 ;
	    RECT 1501.8000 644.4000 1503.0000 644.5500 ;
	    RECT 1504.2001 645.4500 1505.4000 645.6000 ;
	    RECT 1523.4000 645.4500 1524.6000 645.6000 ;
	    RECT 1504.2001 644.5500 1524.6000 645.4500 ;
	    RECT 1525.5000 644.7000 1527.0000 645.6000 ;
	    RECT 1529.4000 644.7000 1529.7001 646.2000 ;
	    RECT 1504.2001 644.4000 1505.4000 644.5500 ;
	    RECT 1523.4000 644.4000 1524.6000 644.5500 ;
	    RECT 1499.4000 639.4500 1500.6000 639.6000 ;
	    RECT 1504.2001 639.4500 1505.4000 639.6000 ;
	    RECT 1493.1000 633.3000 1494.3000 639.3000 ;
	    RECT 1497.0000 633.3000 1498.2001 639.3000 ;
	    RECT 1499.4000 638.5500 1505.4000 639.4500 ;
	    RECT 1499.4000 638.4000 1500.6000 638.5500 ;
	    RECT 1504.2001 638.4000 1505.4000 638.5500 ;
	    RECT 1523.4000 638.4000 1524.6000 639.6000 ;
	    RECT 1526.1000 639.3000 1527.0000 644.7000 ;
	    RECT 1530.6000 644.4000 1531.8000 645.6000 ;
	    RECT 1528.2001 643.5000 1529.4000 643.8000 ;
	    RECT 1547.4000 643.5000 1548.6000 659.7000 ;
	    RECT 1528.2001 641.4000 1529.4000 642.6000 ;
	    RECT 1547.4000 641.4000 1548.6000 642.6000 ;
	    RECT 1535.4000 639.4500 1536.6000 639.6000 ;
	    RECT 1545.0000 639.4500 1546.2001 639.6000 ;
	    RECT 1499.1000 637.2000 1500.3000 637.5000 ;
	    RECT 1523.7001 637.2000 1524.9000 637.5000 ;
	    RECT 1499.4000 633.3000 1500.6000 636.3000 ;
	    RECT 1523.4000 633.3000 1524.6000 636.3000 ;
	    RECT 1525.8000 633.3000 1527.0000 639.3000 ;
	    RECT 1529.7001 633.3000 1530.9000 639.3000 ;
	    RECT 1535.4000 638.5500 1546.2001 639.4500 ;
	    RECT 1535.4000 638.4000 1536.6000 638.5500 ;
	    RECT 1545.0000 638.4000 1546.2001 638.5500 ;
	    RECT 1545.0000 637.2000 1546.2001 637.5000 ;
	    RECT 1545.0000 633.3000 1546.2001 636.3000 ;
	    RECT 1547.4000 633.3000 1548.6000 640.5000 ;
	    RECT 1.2000 630.6000 1569.0000 632.4000 ;
	    RECT 126.6000 620.7000 127.8000 629.7000 ;
	    RECT 131.4000 623.7000 132.6000 629.7000 ;
	    RECT 136.2000 624.9000 137.4000 629.7000 ;
	    RECT 138.6000 625.5000 139.8000 629.7000 ;
	    RECT 141.0000 625.5000 142.2000 629.7000 ;
	    RECT 143.4000 625.5000 144.6000 629.7000 ;
	    RECT 145.8000 626.7000 147.0000 629.7000 ;
	    RECT 148.2000 625.5000 149.4000 629.7000 ;
	    RECT 150.6000 626.7000 151.8000 629.7000 ;
	    RECT 153.0000 625.5000 154.2000 629.7000 ;
	    RECT 155.4000 625.5000 156.6000 629.7000 ;
	    RECT 157.8000 625.5000 159.0000 629.7000 ;
	    RECT 160.2000 625.5000 161.4000 629.7000 ;
	    RECT 133.5000 623.7000 137.4000 624.9000 ;
	    RECT 162.6000 624.9000 163.8000 629.7000 ;
	    RECT 142.5000 623.7000 149.4000 624.6000 ;
	    RECT 133.5000 622.8000 134.7000 623.7000 ;
	    RECT 130.2000 621.6000 134.7000 622.8000 ;
	    RECT 126.6000 619.5000 139.8000 620.7000 ;
	    RECT 142.5000 620.1000 143.7000 623.7000 ;
	    RECT 148.2000 623.4000 149.4000 623.7000 ;
	    RECT 150.6000 623.4000 151.8000 624.6000 ;
	    RECT 152.7000 623.4000 153.0000 624.6000 ;
	    RECT 157.5000 623.4000 159.0000 624.6000 ;
	    RECT 162.6000 623.7000 166.2000 624.9000 ;
	    RECT 167.4000 623.7000 168.6000 629.7000 ;
	    RECT 145.8000 622.5000 147.0000 622.8000 ;
	    RECT 148.2000 622.2000 149.4000 622.5000 ;
	    RECT 145.8000 620.4000 147.0000 621.6000 ;
	    RECT 148.2000 621.3000 154.8000 622.2000 ;
	    RECT 153.6000 621.0000 154.8000 621.3000 ;
	    RECT 126.6000 611.1000 127.8000 619.5000 ;
	    RECT 140.7000 618.9000 143.7000 620.1000 ;
	    RECT 149.4000 618.9000 154.2000 620.1000 ;
	    RECT 157.8000 619.2000 159.0000 623.4000 ;
	    RECT 165.0000 622.8000 166.2000 623.7000 ;
	    RECT 165.0000 621.9000 167.7000 622.8000 ;
	    RECT 166.5000 620.1000 167.7000 621.9000 ;
	    RECT 172.2000 621.9000 173.4000 629.7000 ;
	    RECT 174.6000 624.0000 175.8000 629.7000 ;
	    RECT 177.0000 626.7000 178.2000 629.7000 ;
	    RECT 174.6000 622.8000 176.1000 624.0000 ;
	    RECT 172.2000 621.0000 174.0000 621.9000 ;
	    RECT 166.5000 618.9000 172.2000 620.1000 ;
	    RECT 128.7000 618.0000 129.9000 618.3000 ;
	    RECT 128.7000 617.1000 135.3000 618.0000 ;
	    RECT 136.2000 617.4000 137.4000 618.6000 ;
	    RECT 162.6000 618.0000 163.8000 618.9000 ;
	    RECT 173.1000 618.0000 174.0000 621.0000 ;
	    RECT 138.3000 617.1000 163.8000 618.0000 ;
	    RECT 172.8000 617.1000 174.0000 618.0000 ;
	    RECT 170.7000 616.2000 171.9000 616.5000 ;
	    RECT 131.4000 614.4000 132.6000 615.6000 ;
	    RECT 133.5000 615.3000 171.9000 616.2000 ;
	    RECT 136.5000 615.0000 137.7000 615.3000 ;
	    RECT 172.8000 614.4000 173.7000 617.1000 ;
	    RECT 174.9000 616.2000 176.1000 622.8000 ;
	    RECT 191.4000 622.5000 192.6000 629.7000 ;
	    RECT 193.8000 626.7000 195.0000 629.7000 ;
	    RECT 193.8000 625.5000 195.0000 625.8000 ;
	    RECT 193.8000 624.4500 195.0000 624.6000 ;
	    RECT 196.2000 624.4500 197.4000 624.6000 ;
	    RECT 193.8000 623.5500 197.4000 624.4500 ;
	    RECT 193.8000 623.4000 195.0000 623.5500 ;
	    RECT 196.2000 623.4000 197.4000 623.5500 ;
	    RECT 213.0000 622.5000 214.2000 629.7000 ;
	    RECT 215.4000 626.7000 216.6000 629.7000 ;
	    RECT 234.6000 626.7000 235.8000 629.7000 ;
	    RECT 237.0000 626.7000 238.2000 629.7000 ;
	    RECT 239.4000 626.7000 240.6000 629.7000 ;
	    RECT 258.6000 626.7000 259.8000 629.7000 ;
	    RECT 261.0000 626.7000 262.2000 629.7000 ;
	    RECT 263.4000 626.7000 264.6000 629.7000 ;
	    RECT 215.4000 625.5000 216.6000 625.8000 ;
	    RECT 234.6000 625.5000 235.8000 625.8000 ;
	    RECT 215.4000 623.4000 216.6000 624.6000 ;
	    RECT 234.6000 623.4000 235.8000 624.6000 ;
	    RECT 237.3000 622.5000 238.2000 626.7000 ;
	    RECT 258.6000 625.5000 259.8000 625.8000 ;
	    RECT 258.6000 623.4000 259.8000 624.6000 ;
	    RECT 261.3000 622.5000 262.2000 626.7000 ;
	    RECT 289.8000 623.7000 291.0000 629.7000 ;
	    RECT 292.2000 624.0000 293.4000 629.7000 ;
	    RECT 294.6000 624.9000 295.8000 629.7000 ;
	    RECT 297.0000 624.0000 298.2000 629.7000 ;
	    RECT 292.2000 623.7000 298.2000 624.0000 ;
	    RECT 290.1000 622.5000 291.0000 623.7000 ;
	    RECT 292.5000 623.1000 297.9000 623.7000 ;
	    RECT 309.0000 622.5000 310.2000 629.7000 ;
	    RECT 311.4000 626.7000 312.6000 629.7000 ;
	    RECT 330.6000 626.7000 331.8000 629.7000 ;
	    RECT 333.0000 626.7000 334.2000 629.7000 ;
	    RECT 335.4000 626.7000 336.6000 629.7000 ;
	    RECT 311.4000 625.5000 312.6000 625.8000 ;
	    RECT 311.4000 624.4500 312.6000 624.6000 ;
	    RECT 316.2000 624.4500 317.4000 624.6000 ;
	    RECT 311.4000 623.5500 317.4000 624.4500 ;
	    RECT 311.4000 623.4000 312.6000 623.5500 ;
	    RECT 316.2000 623.4000 317.4000 623.5500 ;
	    RECT 333.0000 622.5000 333.9000 626.7000 ;
	    RECT 335.4000 625.5000 336.6000 625.8000 ;
	    RECT 335.4000 624.4500 336.6000 624.6000 ;
	    RECT 340.2000 624.4500 341.4000 624.6000 ;
	    RECT 335.4000 623.5500 341.4000 624.4500 ;
	    RECT 359.4000 623.7000 360.6000 629.7000 ;
	    RECT 361.8000 624.0000 363.0000 629.7000 ;
	    RECT 364.2000 624.9000 365.4000 629.7000 ;
	    RECT 366.6000 624.0000 367.8000 629.7000 ;
	    RECT 361.8000 623.7000 367.8000 624.0000 ;
	    RECT 386.7000 624.6000 387.9000 629.7000 ;
	    RECT 386.7000 623.7000 389.4000 624.6000 ;
	    RECT 390.6000 623.7000 391.8000 629.7000 ;
	    RECT 335.4000 623.4000 336.6000 623.5500 ;
	    RECT 340.2000 623.4000 341.4000 623.5500 ;
	    RECT 359.7000 622.5000 360.6000 623.7000 ;
	    RECT 362.1000 623.1000 367.5000 623.7000 ;
	    RECT 177.0000 621.4500 178.2000 621.6000 ;
	    RECT 191.4000 621.4500 192.6000 621.6000 ;
	    RECT 177.0000 620.5500 192.6000 621.4500 ;
	    RECT 177.0000 620.4000 178.2000 620.5500 ;
	    RECT 191.4000 620.4000 192.6000 620.5500 ;
	    RECT 213.0000 621.4500 214.2000 621.6000 ;
	    RECT 227.4000 621.4500 228.6000 621.6000 ;
	    RECT 213.0000 620.5500 228.6000 621.4500 ;
	    RECT 213.0000 620.4000 214.2000 620.5500 ;
	    RECT 227.4000 620.4000 228.6000 620.5500 ;
	    RECT 237.0000 620.4000 238.2000 621.6000 ;
	    RECT 251.4000 621.4500 252.6000 621.6000 ;
	    RECT 261.0000 621.4500 262.2000 621.6000 ;
	    RECT 251.4000 620.5500 262.2000 621.4500 ;
	    RECT 251.4000 620.4000 252.6000 620.5500 ;
	    RECT 261.0000 620.4000 262.2000 620.5500 ;
	    RECT 285.0000 621.4500 286.2000 621.6000 ;
	    RECT 289.8000 621.4500 291.0000 621.6000 ;
	    RECT 285.0000 620.5500 291.0000 621.4500 ;
	    RECT 285.0000 620.4000 286.2000 620.5500 ;
	    RECT 289.8000 620.4000 291.0000 620.5500 ;
	    RECT 291.9000 620.4000 293.7000 621.6000 ;
	    RECT 295.8000 620.7000 296.1000 622.2000 ;
	    RECT 297.0000 620.4000 298.2000 621.6000 ;
	    RECT 309.0000 621.4500 310.2000 621.6000 ;
	    RECT 299.5500 620.5500 310.2000 621.4500 ;
	    RECT 141.0000 614.1000 142.2000 614.4000 ;
	    RECT 134.1000 613.5000 142.2000 614.1000 ;
	    RECT 132.9000 613.2000 142.2000 613.5000 ;
	    RECT 143.7000 613.5000 156.6000 614.4000 ;
	    RECT 129.0000 612.0000 131.4000 613.2000 ;
	    RECT 132.9000 612.3000 135.0000 613.2000 ;
	    RECT 143.7000 612.3000 144.6000 613.5000 ;
	    RECT 155.4000 613.2000 156.6000 613.5000 ;
	    RECT 160.2000 613.5000 173.7000 614.4000 ;
	    RECT 174.6000 615.0000 176.1000 616.2000 ;
	    RECT 174.6000 613.5000 175.8000 615.0000 ;
	    RECT 160.2000 613.2000 161.4000 613.5000 ;
	    RECT 130.5000 611.4000 131.4000 612.0000 ;
	    RECT 135.9000 611.4000 144.6000 612.3000 ;
	    RECT 145.5000 611.4000 149.4000 612.6000 ;
	    RECT 126.6000 610.2000 129.6000 611.1000 ;
	    RECT 130.5000 610.2000 136.8000 611.4000 ;
	    RECT 128.7000 609.3000 129.6000 610.2000 ;
	    RECT 126.6000 603.3000 127.8000 609.3000 ;
	    RECT 128.7000 608.4000 130.2000 609.3000 ;
	    RECT 129.0000 603.3000 130.2000 608.4000 ;
	    RECT 131.4000 602.4000 132.6000 609.3000 ;
	    RECT 133.8000 603.3000 135.0000 610.2000 ;
	    RECT 136.2000 603.3000 137.4000 609.3000 ;
	    RECT 138.6000 603.3000 139.8000 607.5000 ;
	    RECT 141.0000 603.3000 142.2000 607.5000 ;
	    RECT 143.4000 603.3000 144.6000 610.5000 ;
	    RECT 145.8000 603.3000 147.0000 609.3000 ;
	    RECT 148.2000 603.3000 149.4000 610.5000 ;
	    RECT 150.6000 603.3000 151.8000 609.3000 ;
	    RECT 153.0000 603.3000 154.2000 612.6000 ;
	    RECT 165.0000 611.4000 168.9000 612.6000 ;
	    RECT 157.8000 610.2000 164.1000 611.4000 ;
	    RECT 155.4000 603.3000 156.6000 607.5000 ;
	    RECT 157.8000 603.3000 159.0000 607.5000 ;
	    RECT 160.2000 603.3000 161.4000 607.5000 ;
	    RECT 162.6000 603.3000 163.8000 609.3000 ;
	    RECT 165.0000 603.3000 166.2000 611.4000 ;
	    RECT 172.8000 611.1000 173.7000 613.5000 ;
	    RECT 174.6000 611.4000 175.8000 612.6000 ;
	    RECT 169.8000 610.2000 173.7000 611.1000 ;
	    RECT 167.4000 603.3000 168.6000 609.3000 ;
	    RECT 169.8000 603.3000 171.0000 610.2000 ;
	    RECT 172.2000 603.3000 173.4000 609.3000 ;
	    RECT 174.6000 603.3000 175.8000 610.5000 ;
	    RECT 177.0000 603.3000 178.2000 609.3000 ;
	    RECT 191.4000 603.3000 192.6000 619.5000 ;
	    RECT 193.8000 603.3000 195.0000 609.3000 ;
	    RECT 213.0000 603.3000 214.2000 619.5000 ;
	    RECT 237.3000 615.3000 238.2000 619.5000 ;
	    RECT 239.4000 617.4000 240.6000 618.6000 ;
	    RECT 241.8000 618.4500 243.0000 618.6000 ;
	    RECT 249.0000 618.4500 250.2000 618.6000 ;
	    RECT 241.8000 617.5500 250.2000 618.4500 ;
	    RECT 241.8000 617.4000 243.0000 617.5500 ;
	    RECT 249.0000 617.4000 250.2000 617.5500 ;
	    RECT 239.4000 616.2000 240.6000 616.5000 ;
	    RECT 261.3000 615.3000 262.2000 619.5000 ;
	    RECT 263.4000 618.4500 264.6000 618.6000 ;
	    RECT 282.6000 618.4500 283.8000 618.6000 ;
	    RECT 263.4000 617.5500 283.8000 618.4500 ;
	    RECT 263.4000 617.4000 264.6000 617.5500 ;
	    RECT 282.6000 617.4000 283.8000 617.5500 ;
	    RECT 263.4000 616.2000 264.6000 616.5000 ;
	    RECT 277.8000 615.4500 279.0000 615.6000 ;
	    RECT 289.8000 615.4500 291.0000 615.6000 ;
	    RECT 215.4000 603.3000 216.6000 609.3000 ;
	    RECT 234.6000 603.3000 235.8000 615.3000 ;
	    RECT 237.0000 614.1000 239.7000 615.3000 ;
	    RECT 238.5000 603.3000 239.7000 614.1000 ;
	    RECT 258.6000 603.3000 259.8000 615.3000 ;
	    RECT 261.0000 614.1000 263.7000 615.3000 ;
	    RECT 277.8000 614.5500 291.0000 615.4500 ;
	    RECT 277.8000 614.4000 279.0000 614.5500 ;
	    RECT 289.8000 614.4000 291.0000 614.5500 ;
	    RECT 292.8000 615.3000 293.7000 620.4000 ;
	    RECT 294.6000 619.5000 295.8000 619.8000 ;
	    RECT 294.6000 618.4500 295.8000 618.6000 ;
	    RECT 299.5500 618.4500 300.4500 620.5500 ;
	    RECT 309.0000 620.4000 310.2000 620.5500 ;
	    RECT 333.0000 621.4500 334.2000 621.6000 ;
	    RECT 357.0000 621.4500 358.2000 621.6000 ;
	    RECT 333.0000 620.5500 358.2000 621.4500 ;
	    RECT 333.0000 620.4000 334.2000 620.5500 ;
	    RECT 357.0000 620.4000 358.2000 620.5500 ;
	    RECT 359.4000 620.4000 360.6000 621.6000 ;
	    RECT 361.5000 620.4000 363.3000 621.6000 ;
	    RECT 365.4000 620.7000 365.7000 622.2000 ;
	    RECT 366.6000 620.4000 367.8000 621.6000 ;
	    RECT 294.6000 617.5500 300.4500 618.4500 ;
	    RECT 294.6000 617.4000 295.8000 617.5500 ;
	    RECT 292.8000 614.4000 294.3000 615.3000 ;
	    RECT 262.5000 603.3000 263.7000 614.1000 ;
	    RECT 291.0000 612.6000 291.9000 613.5000 ;
	    RECT 291.0000 611.4000 292.2000 612.6000 ;
	    RECT 290.7000 603.3000 291.9000 609.3000 ;
	    RECT 293.1000 603.3000 294.3000 614.4000 ;
	    RECT 297.0000 603.3000 298.2000 615.3000 ;
	    RECT 309.0000 603.3000 310.2000 619.5000 ;
	    RECT 330.6000 617.4000 331.8000 618.6000 ;
	    RECT 330.6000 616.2000 331.8000 616.5000 ;
	    RECT 333.0000 615.3000 333.9000 619.5000 ;
	    RECT 331.5000 614.1000 334.2000 615.3000 ;
	    RECT 311.4000 603.3000 312.6000 609.3000 ;
	    RECT 331.5000 603.3000 332.7000 614.1000 ;
	    RECT 335.4000 603.3000 336.6000 615.3000 ;
	    RECT 359.4000 614.4000 360.6000 615.6000 ;
	    RECT 362.4000 615.3000 363.3000 620.4000 ;
	    RECT 364.2000 619.5000 365.4000 619.8000 ;
	    RECT 388.2000 619.5000 389.4000 623.7000 ;
	    RECT 390.6000 622.5000 391.8000 622.8000 ;
	    RECT 405.0000 622.5000 406.2000 629.7000 ;
	    RECT 407.4000 626.7000 408.6000 629.7000 ;
	    RECT 407.4000 625.5000 408.6000 625.8000 ;
	    RECT 407.4000 624.4500 408.6000 624.6000 ;
	    RECT 426.6000 624.4500 427.8000 624.6000 ;
	    RECT 407.4000 623.5500 427.8000 624.4500 ;
	    RECT 438.6000 623.7000 439.8000 629.7000 ;
	    RECT 441.0000 624.0000 442.2000 629.7000 ;
	    RECT 443.4000 624.9000 444.6000 629.7000 ;
	    RECT 445.8000 624.0000 447.0000 629.7000 ;
	    RECT 441.0000 623.7000 447.0000 624.0000 ;
	    RECT 407.4000 623.4000 408.6000 623.5500 ;
	    RECT 426.6000 623.4000 427.8000 623.5500 ;
	    RECT 438.9000 622.5000 439.8000 623.7000 ;
	    RECT 441.3000 623.1000 446.7000 623.7000 ;
	    RECT 460.2000 622.5000 461.4000 629.7000 ;
	    RECT 462.6000 626.7000 463.8000 629.7000 ;
	    RECT 462.6000 625.5000 463.8000 625.8000 ;
	    RECT 462.6000 624.4500 463.8000 624.6000 ;
	    RECT 474.6000 624.4500 475.8000 624.6000 ;
	    RECT 462.6000 623.5500 475.8000 624.4500 ;
	    RECT 462.6000 623.4000 463.8000 623.5500 ;
	    RECT 474.6000 623.4000 475.8000 623.5500 ;
	    RECT 477.0000 622.5000 478.2000 629.7000 ;
	    RECT 479.4000 626.7000 480.6000 629.7000 ;
	    RECT 479.4000 625.5000 480.6000 625.8000 ;
	    RECT 479.4000 624.4500 480.6000 624.6000 ;
	    RECT 491.4000 624.4500 492.6000 624.6000 ;
	    RECT 479.4000 623.5500 492.6000 624.4500 ;
	    RECT 479.4000 623.4000 480.6000 623.5500 ;
	    RECT 491.4000 623.4000 492.6000 623.5500 ;
	    RECT 493.8000 622.5000 495.0000 629.7000 ;
	    RECT 496.2000 626.7000 497.4000 629.7000 ;
	    RECT 496.2000 625.5000 497.4000 625.8000 ;
	    RECT 496.2000 624.4500 497.4000 624.6000 ;
	    RECT 618.6000 624.4500 619.8000 624.6000 ;
	    RECT 496.2000 623.5500 619.8000 624.4500 ;
	    RECT 496.2000 623.4000 497.4000 623.5500 ;
	    RECT 618.6000 623.4000 619.8000 623.5500 ;
	    RECT 390.6000 620.4000 391.8000 621.6000 ;
	    RECT 405.0000 621.4500 406.2000 621.6000 ;
	    RECT 424.2000 621.4500 425.4000 621.6000 ;
	    RECT 405.0000 620.5500 425.4000 621.4500 ;
	    RECT 405.0000 620.4000 406.2000 620.5500 ;
	    RECT 424.2000 620.4000 425.4000 620.5500 ;
	    RECT 431.4000 621.4500 432.6000 621.6000 ;
	    RECT 438.6000 621.4500 439.8000 621.6000 ;
	    RECT 431.4000 620.5500 439.8000 621.4500 ;
	    RECT 431.4000 620.4000 432.6000 620.5500 ;
	    RECT 438.6000 620.4000 439.8000 620.5500 ;
	    RECT 440.7000 620.4000 442.5000 621.6000 ;
	    RECT 444.6000 620.7000 444.9000 622.2000 ;
	    RECT 445.8000 621.4500 447.0000 621.6000 ;
	    RECT 450.6000 621.4500 451.8000 621.6000 ;
	    RECT 445.8000 620.5500 451.8000 621.4500 ;
	    RECT 445.8000 620.4000 447.0000 620.5500 ;
	    RECT 450.6000 620.4000 451.8000 620.5500 ;
	    RECT 460.2000 621.4500 461.4000 621.6000 ;
	    RECT 462.6000 621.4500 463.8000 621.6000 ;
	    RECT 460.2000 620.5500 463.8000 621.4500 ;
	    RECT 460.2000 620.4000 461.4000 620.5500 ;
	    RECT 462.6000 620.4000 463.8000 620.5500 ;
	    RECT 465.0000 621.4500 466.2000 621.6000 ;
	    RECT 477.0000 621.4500 478.2000 621.6000 ;
	    RECT 465.0000 620.5500 478.2000 621.4500 ;
	    RECT 465.0000 620.4000 466.2000 620.5500 ;
	    RECT 477.0000 620.4000 478.2000 620.5500 ;
	    RECT 493.8000 621.4500 495.0000 621.6000 ;
	    RECT 508.2000 621.4500 509.4000 621.6000 ;
	    RECT 522.6000 621.4500 523.8000 621.6000 ;
	    RECT 493.8000 620.5500 523.8000 621.4500 ;
	    RECT 493.8000 620.4000 495.0000 620.5500 ;
	    RECT 508.2000 620.4000 509.4000 620.5500 ;
	    RECT 522.6000 620.4000 523.8000 620.5500 ;
	    RECT 623.4000 620.7000 624.6000 629.7000 ;
	    RECT 628.2000 623.7000 629.4000 629.7000 ;
	    RECT 633.0000 624.9000 634.2000 629.7000 ;
	    RECT 635.4000 625.5000 636.6000 629.7000 ;
	    RECT 637.8000 625.5000 639.0000 629.7000 ;
	    RECT 640.2000 625.5000 641.4000 629.7000 ;
	    RECT 642.6000 626.7000 643.8000 629.7000 ;
	    RECT 645.0000 625.5000 646.2000 629.7000 ;
	    RECT 647.4000 626.7000 648.6000 629.7000 ;
	    RECT 649.8000 625.5000 651.0000 629.7000 ;
	    RECT 652.2000 625.5000 653.4000 629.7000 ;
	    RECT 654.6000 625.5000 655.8000 629.7000 ;
	    RECT 657.0000 625.5000 658.2000 629.7000 ;
	    RECT 630.3000 623.7000 634.2000 624.9000 ;
	    RECT 659.4000 624.9000 660.6000 629.7000 ;
	    RECT 639.3000 623.7000 646.2000 624.6000 ;
	    RECT 630.3000 622.8000 631.5000 623.7000 ;
	    RECT 627.0000 621.6000 631.5000 622.8000 ;
	    RECT 364.2000 617.4000 365.4000 618.6000 ;
	    RECT 388.2000 617.4000 389.4000 618.6000 ;
	    RECT 362.4000 614.4000 363.9000 615.3000 ;
	    RECT 360.6000 612.6000 361.5000 613.5000 ;
	    RECT 360.6000 611.4000 361.8000 612.6000 ;
	    RECT 360.3000 603.3000 361.5000 609.3000 ;
	    RECT 362.7000 603.3000 363.9000 614.4000 ;
	    RECT 366.6000 603.3000 367.8000 615.3000 ;
	    RECT 385.8000 614.4000 387.0000 615.6000 ;
	    RECT 385.8000 613.2000 387.0000 613.5000 ;
	    RECT 385.8000 603.3000 387.0000 609.3000 ;
	    RECT 388.2000 603.3000 389.4000 616.5000 ;
	    RECT 390.6000 603.3000 391.8000 609.3000 ;
	    RECT 405.0000 603.3000 406.2000 619.5000 ;
	    RECT 429.0000 615.4500 430.2000 615.6000 ;
	    RECT 438.6000 615.4500 439.8000 615.6000 ;
	    RECT 429.0000 614.5500 439.8000 615.4500 ;
	    RECT 429.0000 614.4000 430.2000 614.5500 ;
	    RECT 438.6000 614.4000 439.8000 614.5500 ;
	    RECT 441.6000 615.3000 442.5000 620.4000 ;
	    RECT 443.4000 619.5000 444.6000 619.8000 ;
	    RECT 623.4000 619.5000 636.6000 620.7000 ;
	    RECT 639.3000 620.1000 640.5000 623.7000 ;
	    RECT 645.0000 623.4000 646.2000 623.7000 ;
	    RECT 647.4000 623.4000 648.6000 624.6000 ;
	    RECT 649.5000 623.4000 649.8000 624.6000 ;
	    RECT 654.3000 623.4000 655.8000 624.6000 ;
	    RECT 659.4000 623.7000 663.0000 624.9000 ;
	    RECT 664.2000 623.7000 665.4000 629.7000 ;
	    RECT 642.6000 622.5000 643.8000 622.8000 ;
	    RECT 645.0000 622.2000 646.2000 622.5000 ;
	    RECT 642.6000 620.4000 643.8000 621.6000 ;
	    RECT 645.0000 621.3000 651.6000 622.2000 ;
	    RECT 650.4000 621.0000 651.6000 621.3000 ;
	    RECT 443.4000 618.4500 444.6000 618.6000 ;
	    RECT 445.8000 618.4500 447.0000 618.6000 ;
	    RECT 443.4000 617.5500 447.0000 618.4500 ;
	    RECT 443.4000 617.4000 444.6000 617.5500 ;
	    RECT 445.8000 617.4000 447.0000 617.5500 ;
	    RECT 441.6000 614.4000 443.1000 615.3000 ;
	    RECT 439.8000 612.6000 440.7000 613.5000 ;
	    RECT 439.8000 611.4000 441.0000 612.6000 ;
	    RECT 407.4000 603.3000 408.6000 609.3000 ;
	    RECT 439.5000 603.3000 440.7000 609.3000 ;
	    RECT 441.9000 603.3000 443.1000 614.4000 ;
	    RECT 445.8000 603.3000 447.0000 615.3000 ;
	    RECT 460.2000 603.3000 461.4000 619.5000 ;
	    RECT 462.6000 603.3000 463.8000 609.3000 ;
	    RECT 477.0000 603.3000 478.2000 619.5000 ;
	    RECT 479.4000 603.3000 480.6000 609.3000 ;
	    RECT 493.8000 603.3000 495.0000 619.5000 ;
	    RECT 623.4000 611.1000 624.6000 619.5000 ;
	    RECT 637.5000 618.9000 640.5000 620.1000 ;
	    RECT 646.2000 618.9000 651.0000 620.1000 ;
	    RECT 654.6000 619.2000 655.8000 623.4000 ;
	    RECT 661.8000 622.8000 663.0000 623.7000 ;
	    RECT 661.8000 621.9000 664.5000 622.8000 ;
	    RECT 663.3000 620.1000 664.5000 621.9000 ;
	    RECT 669.0000 621.9000 670.2000 629.7000 ;
	    RECT 671.4000 624.0000 672.6000 629.7000 ;
	    RECT 673.8000 626.7000 675.0000 629.7000 ;
	    RECT 695.4000 626.7000 696.6000 629.7000 ;
	    RECT 695.4000 625.5000 696.6000 625.8000 ;
	    RECT 671.4000 622.8000 672.9000 624.0000 ;
	    RECT 695.4000 623.4000 696.6000 624.6000 ;
	    RECT 669.0000 621.0000 670.8000 621.9000 ;
	    RECT 663.3000 618.9000 669.0000 620.1000 ;
	    RECT 625.5000 618.0000 626.7000 618.3000 ;
	    RECT 625.5000 617.1000 632.1000 618.0000 ;
	    RECT 633.0000 617.4000 634.2000 618.6000 ;
	    RECT 659.4000 618.0000 660.6000 618.9000 ;
	    RECT 669.9000 618.0000 670.8000 621.0000 ;
	    RECT 635.1000 617.1000 660.6000 618.0000 ;
	    RECT 669.6000 617.1000 670.8000 618.0000 ;
	    RECT 667.5000 616.2000 668.7000 616.5000 ;
	    RECT 628.2000 614.4000 629.4000 615.6000 ;
	    RECT 630.3000 615.3000 668.7000 616.2000 ;
	    RECT 633.3000 615.0000 634.5000 615.3000 ;
	    RECT 669.6000 614.4000 670.5000 617.1000 ;
	    RECT 671.7000 616.2000 672.9000 622.8000 ;
	    RECT 697.8000 622.5000 699.0000 629.7000 ;
	    RECT 712.2000 622.5000 713.4000 629.7000 ;
	    RECT 714.6000 626.7000 715.8000 629.7000 ;
	    RECT 743.4000 628.8000 749.4000 629.7000 ;
	    RECT 714.6000 625.5000 715.8000 625.8000 ;
	    RECT 714.6000 623.4000 715.8000 624.6000 ;
	    RECT 743.4000 623.7000 744.6000 628.8000 ;
	    RECT 745.8000 623.7000 747.0000 627.9000 ;
	    RECT 748.2000 624.0000 749.4000 628.8000 ;
	    RECT 750.6000 624.9000 751.8000 629.7000 ;
	    RECT 753.0000 624.0000 754.2000 629.7000 ;
	    RECT 755.4000 627.4500 756.6000 627.6000 ;
	    RECT 817.8000 627.4500 819.0000 627.6000 ;
	    RECT 755.4000 626.5500 819.0000 627.4500 ;
	    RECT 755.4000 626.4000 756.6000 626.5500 ;
	    RECT 817.8000 626.4000 819.0000 626.5500 ;
	    RECT 748.2000 623.7000 754.2000 624.0000 ;
	    RECT 745.8000 621.6000 746.7000 623.7000 ;
	    RECT 748.5000 623.1000 753.9000 623.7000 ;
	    RECT 697.8000 621.4500 699.0000 621.6000 ;
	    RECT 709.8000 621.4500 711.0000 621.6000 ;
	    RECT 697.8000 620.5500 711.0000 621.4500 ;
	    RECT 697.8000 620.4000 699.0000 620.5500 ;
	    RECT 709.8000 620.4000 711.0000 620.5500 ;
	    RECT 712.2000 620.4000 713.4000 621.6000 ;
	    RECT 731.4000 621.4500 732.6000 621.6000 ;
	    RECT 743.4000 621.4500 744.6000 621.6000 ;
	    RECT 731.4000 620.5500 744.6000 621.4500 ;
	    RECT 745.8000 620.7000 747.3000 621.6000 ;
	    RECT 731.4000 620.4000 732.6000 620.5500 ;
	    RECT 743.4000 620.4000 744.6000 620.5500 ;
	    RECT 748.2000 620.4000 749.4000 621.6000 ;
	    RECT 751.8000 620.7000 752.1000 622.2000 ;
	    RECT 753.0000 620.4000 754.2000 621.6000 ;
	    RECT 779.4000 621.4500 780.6000 621.6000 ;
	    RECT 882.6000 621.4500 883.8000 621.6000 ;
	    RECT 779.4000 620.5500 883.8000 621.4500 ;
	    RECT 779.4000 620.4000 780.6000 620.5500 ;
	    RECT 882.6000 620.4000 883.8000 620.5500 ;
	    RECT 887.4000 620.7000 888.6000 629.7000 ;
	    RECT 892.2000 623.7000 893.4000 629.7000 ;
	    RECT 897.0000 624.9000 898.2000 629.7000 ;
	    RECT 899.4000 625.5000 900.6000 629.7000 ;
	    RECT 901.8000 625.5000 903.0000 629.7000 ;
	    RECT 904.2000 625.5000 905.4000 629.7000 ;
	    RECT 906.6000 626.7000 907.8000 629.7000 ;
	    RECT 909.0000 625.5000 910.2000 629.7000 ;
	    RECT 911.4000 626.7000 912.6000 629.7000 ;
	    RECT 913.8000 625.5000 915.0000 629.7000 ;
	    RECT 916.2000 625.5000 917.4000 629.7000 ;
	    RECT 918.6000 625.5000 919.8000 629.7000 ;
	    RECT 921.0000 625.5000 922.2000 629.7000 ;
	    RECT 894.3000 623.7000 898.2000 624.9000 ;
	    RECT 923.4000 624.9000 924.6000 629.7000 ;
	    RECT 903.3000 623.7000 910.2000 624.6000 ;
	    RECT 894.3000 622.8000 895.5000 623.7000 ;
	    RECT 891.0000 621.6000 895.5000 622.8000 ;
	    RECT 745.8000 619.5000 747.0000 619.8000 ;
	    RECT 750.6000 619.5000 751.8000 619.8000 ;
	    RECT 887.4000 619.5000 900.6000 620.7000 ;
	    RECT 903.3000 620.1000 904.5000 623.7000 ;
	    RECT 909.0000 623.4000 910.2000 623.7000 ;
	    RECT 911.4000 623.4000 912.6000 624.6000 ;
	    RECT 913.5000 623.4000 913.8000 624.6000 ;
	    RECT 918.3000 623.4000 919.8000 624.6000 ;
	    RECT 923.4000 623.7000 927.0000 624.9000 ;
	    RECT 928.2000 623.7000 929.4000 629.7000 ;
	    RECT 906.6000 622.5000 907.8000 622.8000 ;
	    RECT 909.0000 622.2000 910.2000 622.5000 ;
	    RECT 906.6000 620.4000 907.8000 621.6000 ;
	    RECT 909.0000 621.3000 915.6000 622.2000 ;
	    RECT 914.4000 621.0000 915.6000 621.3000 ;
	    RECT 637.8000 614.1000 639.0000 614.4000 ;
	    RECT 630.9000 613.5000 639.0000 614.1000 ;
	    RECT 629.7000 613.2000 639.0000 613.5000 ;
	    RECT 640.5000 613.5000 653.4000 614.4000 ;
	    RECT 625.8000 612.0000 628.2000 613.2000 ;
	    RECT 629.7000 612.3000 631.8000 613.2000 ;
	    RECT 640.5000 612.3000 641.4000 613.5000 ;
	    RECT 652.2000 613.2000 653.4000 613.5000 ;
	    RECT 657.0000 613.5000 670.5000 614.4000 ;
	    RECT 671.4000 615.0000 672.9000 616.2000 ;
	    RECT 671.4000 613.5000 672.6000 615.0000 ;
	    RECT 657.0000 613.2000 658.2000 613.5000 ;
	    RECT 627.3000 611.4000 628.2000 612.0000 ;
	    RECT 632.7000 611.4000 641.4000 612.3000 ;
	    RECT 642.3000 611.4000 646.2000 612.6000 ;
	    RECT 623.4000 610.2000 626.4000 611.1000 ;
	    RECT 627.3000 610.2000 633.6000 611.4000 ;
	    RECT 498.6000 609.4500 499.8000 609.6000 ;
	    RECT 520.2000 609.4500 521.4000 609.6000 ;
	    RECT 496.2000 603.3000 497.4000 609.3000 ;
	    RECT 498.6000 608.5500 521.4000 609.4500 ;
	    RECT 625.5000 609.3000 626.4000 610.2000 ;
	    RECT 498.6000 608.4000 499.8000 608.5500 ;
	    RECT 520.2000 608.4000 521.4000 608.5500 ;
	    RECT 623.4000 603.3000 624.6000 609.3000 ;
	    RECT 625.5000 608.4000 627.0000 609.3000 ;
	    RECT 625.8000 603.3000 627.0000 608.4000 ;
	    RECT 628.2000 602.4000 629.4000 609.3000 ;
	    RECT 630.6000 603.3000 631.8000 610.2000 ;
	    RECT 633.0000 603.3000 634.2000 609.3000 ;
	    RECT 635.4000 603.3000 636.6000 607.5000 ;
	    RECT 637.8000 603.3000 639.0000 607.5000 ;
	    RECT 640.2000 603.3000 641.4000 610.5000 ;
	    RECT 642.6000 603.3000 643.8000 609.3000 ;
	    RECT 645.0000 603.3000 646.2000 610.5000 ;
	    RECT 647.4000 603.3000 648.6000 609.3000 ;
	    RECT 649.8000 603.3000 651.0000 612.6000 ;
	    RECT 661.8000 611.4000 665.7000 612.6000 ;
	    RECT 654.6000 610.2000 660.9000 611.4000 ;
	    RECT 652.2000 603.3000 653.4000 607.5000 ;
	    RECT 654.6000 603.3000 655.8000 607.5000 ;
	    RECT 657.0000 603.3000 658.2000 607.5000 ;
	    RECT 659.4000 603.3000 660.6000 609.3000 ;
	    RECT 661.8000 603.3000 663.0000 611.4000 ;
	    RECT 669.6000 611.1000 670.5000 613.5000 ;
	    RECT 671.4000 611.4000 672.6000 612.6000 ;
	    RECT 666.6000 610.2000 670.5000 611.1000 ;
	    RECT 664.2000 603.3000 665.4000 609.3000 ;
	    RECT 666.6000 603.3000 667.8000 610.2000 ;
	    RECT 669.0000 603.3000 670.2000 609.3000 ;
	    RECT 671.4000 603.3000 672.6000 610.5000 ;
	    RECT 676.2000 609.4500 677.4000 609.6000 ;
	    RECT 683.4000 609.4500 684.6000 609.6000 ;
	    RECT 673.8000 603.3000 675.0000 609.3000 ;
	    RECT 676.2000 608.5500 684.6000 609.4500 ;
	    RECT 676.2000 608.4000 677.4000 608.5500 ;
	    RECT 683.4000 608.4000 684.6000 608.5500 ;
	    RECT 695.4000 603.3000 696.6000 609.3000 ;
	    RECT 697.8000 603.3000 699.0000 619.5000 ;
	    RECT 712.2000 603.3000 713.4000 619.5000 ;
	    RECT 743.4000 619.2000 744.6000 619.5000 ;
	    RECT 745.8000 617.4000 747.0000 618.6000 ;
	    RECT 748.5000 615.3000 749.4000 619.5000 ;
	    RECT 750.6000 618.4500 751.8000 618.6000 ;
	    RECT 820.2000 618.4500 821.4000 618.6000 ;
	    RECT 750.6000 617.5500 821.4000 618.4500 ;
	    RECT 750.6000 617.4000 751.8000 617.5500 ;
	    RECT 820.2000 617.4000 821.4000 617.5500 ;
	    RECT 714.6000 603.3000 715.8000 609.3000 ;
	    RECT 743.4000 603.3000 744.6000 615.3000 ;
	    RECT 747.3000 603.3000 750.3000 615.3000 ;
	    RECT 753.0000 603.3000 754.2000 615.3000 ;
	    RECT 887.4000 611.1000 888.6000 619.5000 ;
	    RECT 901.5000 618.9000 904.5000 620.1000 ;
	    RECT 910.2000 618.9000 915.0000 620.1000 ;
	    RECT 918.6000 619.2000 919.8000 623.4000 ;
	    RECT 925.8000 622.8000 927.0000 623.7000 ;
	    RECT 925.8000 621.9000 928.5000 622.8000 ;
	    RECT 927.3000 620.1000 928.5000 621.9000 ;
	    RECT 933.0000 621.9000 934.2000 629.7000 ;
	    RECT 935.4000 624.0000 936.6000 629.7000 ;
	    RECT 937.8000 626.7000 939.0000 629.7000 ;
	    RECT 949.8000 626.7000 951.0000 629.7000 ;
	    RECT 949.8000 625.5000 951.0000 625.8000 ;
	    RECT 937.8000 624.4500 939.0000 624.6000 ;
	    RECT 949.8000 624.4500 951.0000 624.6000 ;
	    RECT 935.4000 622.8000 936.9000 624.0000 ;
	    RECT 937.8000 623.5500 951.0000 624.4500 ;
	    RECT 937.8000 623.4000 939.0000 623.5500 ;
	    RECT 949.8000 623.4000 951.0000 623.5500 ;
	    RECT 933.0000 621.0000 934.8000 621.9000 ;
	    RECT 927.3000 618.9000 933.0000 620.1000 ;
	    RECT 889.5000 618.0000 890.7000 618.3000 ;
	    RECT 889.5000 617.1000 896.1000 618.0000 ;
	    RECT 897.0000 617.4000 898.2000 618.6000 ;
	    RECT 923.4000 618.0000 924.6000 618.9000 ;
	    RECT 933.9000 618.0000 934.8000 621.0000 ;
	    RECT 899.1000 617.1000 924.6000 618.0000 ;
	    RECT 933.6000 617.1000 934.8000 618.0000 ;
	    RECT 931.5000 616.2000 932.7000 616.5000 ;
	    RECT 892.2000 614.4000 893.4000 615.6000 ;
	    RECT 894.3000 615.3000 932.7000 616.2000 ;
	    RECT 897.3000 615.0000 898.5000 615.3000 ;
	    RECT 933.6000 614.4000 934.5000 617.1000 ;
	    RECT 935.7000 616.2000 936.9000 622.8000 ;
	    RECT 952.2000 622.5000 953.4000 629.7000 ;
	    RECT 1077.0000 626.7000 1078.2001 629.7000 ;
	    RECT 1079.4000 624.0000 1080.6000 629.7000 ;
	    RECT 1079.1000 622.8000 1080.6000 624.0000 ;
	    RECT 952.2000 621.4500 953.4000 621.6000 ;
	    RECT 959.4000 621.4500 960.6000 621.6000 ;
	    RECT 952.2000 620.5500 960.6000 621.4500 ;
	    RECT 952.2000 620.4000 953.4000 620.5500 ;
	    RECT 959.4000 620.4000 960.6000 620.5500 ;
	    RECT 901.8000 614.1000 903.0000 614.4000 ;
	    RECT 894.9000 613.5000 903.0000 614.1000 ;
	    RECT 893.7000 613.2000 903.0000 613.5000 ;
	    RECT 904.5000 613.5000 917.4000 614.4000 ;
	    RECT 889.8000 612.0000 892.2000 613.2000 ;
	    RECT 893.7000 612.3000 895.8000 613.2000 ;
	    RECT 904.5000 612.3000 905.4000 613.5000 ;
	    RECT 916.2000 613.2000 917.4000 613.5000 ;
	    RECT 921.0000 613.5000 934.5000 614.4000 ;
	    RECT 935.4000 615.0000 936.9000 616.2000 ;
	    RECT 935.4000 613.5000 936.6000 615.0000 ;
	    RECT 921.0000 613.2000 922.2000 613.5000 ;
	    RECT 891.3000 611.4000 892.2000 612.0000 ;
	    RECT 896.7000 611.4000 905.4000 612.3000 ;
	    RECT 906.3000 611.4000 910.2000 612.6000 ;
	    RECT 887.4000 610.2000 890.4000 611.1000 ;
	    RECT 891.3000 610.2000 897.6000 611.4000 ;
	    RECT 889.5000 609.3000 890.4000 610.2000 ;
	    RECT 887.4000 603.3000 888.6000 609.3000 ;
	    RECT 889.5000 608.4000 891.0000 609.3000 ;
	    RECT 889.8000 603.3000 891.0000 608.4000 ;
	    RECT 892.2000 602.4000 893.4000 609.3000 ;
	    RECT 894.6000 603.3000 895.8000 610.2000 ;
	    RECT 897.0000 603.3000 898.2000 609.3000 ;
	    RECT 899.4000 603.3000 900.6000 607.5000 ;
	    RECT 901.8000 603.3000 903.0000 607.5000 ;
	    RECT 904.2000 603.3000 905.4000 610.5000 ;
	    RECT 906.6000 603.3000 907.8000 609.3000 ;
	    RECT 909.0000 603.3000 910.2000 610.5000 ;
	    RECT 911.4000 603.3000 912.6000 609.3000 ;
	    RECT 913.8000 603.3000 915.0000 612.6000 ;
	    RECT 925.8000 611.4000 929.7000 612.6000 ;
	    RECT 918.6000 610.2000 924.9000 611.4000 ;
	    RECT 916.2000 603.3000 917.4000 607.5000 ;
	    RECT 918.6000 603.3000 919.8000 607.5000 ;
	    RECT 921.0000 603.3000 922.2000 607.5000 ;
	    RECT 923.4000 603.3000 924.6000 609.3000 ;
	    RECT 925.8000 603.3000 927.0000 611.4000 ;
	    RECT 933.6000 611.1000 934.5000 613.5000 ;
	    RECT 935.4000 612.4500 936.6000 612.6000 ;
	    RECT 937.8000 612.4500 939.0000 612.6000 ;
	    RECT 935.4000 611.5500 939.0000 612.4500 ;
	    RECT 935.4000 611.4000 936.6000 611.5500 ;
	    RECT 937.8000 611.4000 939.0000 611.5500 ;
	    RECT 930.6000 610.2000 934.5000 611.1000 ;
	    RECT 928.2000 603.3000 929.4000 609.3000 ;
	    RECT 930.6000 603.3000 931.8000 610.2000 ;
	    RECT 933.0000 603.3000 934.2000 609.3000 ;
	    RECT 935.4000 603.3000 936.6000 610.5000 ;
	    RECT 937.8000 603.3000 939.0000 609.3000 ;
	    RECT 949.8000 603.3000 951.0000 609.3000 ;
	    RECT 952.2000 603.3000 953.4000 619.5000 ;
	    RECT 1079.1000 616.2000 1080.3000 622.8000 ;
	    RECT 1081.8000 621.9000 1083.0000 629.7000 ;
	    RECT 1086.6000 623.7000 1087.8000 629.7000 ;
	    RECT 1091.4000 624.9000 1092.6000 629.7000 ;
	    RECT 1093.8000 625.5000 1095.0000 629.7000 ;
	    RECT 1096.2001 625.5000 1097.4000 629.7000 ;
	    RECT 1098.6000 625.5000 1099.8000 629.7000 ;
	    RECT 1101.0000 625.5000 1102.2001 629.7000 ;
	    RECT 1103.4000 626.7000 1104.6000 629.7000 ;
	    RECT 1105.8000 625.5000 1107.0000 629.7000 ;
	    RECT 1108.2001 626.7000 1109.4000 629.7000 ;
	    RECT 1110.6000 625.5000 1111.8000 629.7000 ;
	    RECT 1113.0000 625.5000 1114.2001 629.7000 ;
	    RECT 1115.4000 625.5000 1116.6000 629.7000 ;
	    RECT 1089.0000 623.7000 1092.6000 624.9000 ;
	    RECT 1117.8000 624.9000 1119.0000 629.7000 ;
	    RECT 1089.0000 622.8000 1090.2001 623.7000 ;
	    RECT 1081.2001 621.0000 1083.0000 621.9000 ;
	    RECT 1087.5000 621.9000 1090.2001 622.8000 ;
	    RECT 1096.2001 623.4000 1097.7001 624.6000 ;
	    RECT 1102.2001 623.4000 1102.5000 624.6000 ;
	    RECT 1103.4000 623.4000 1104.6000 624.6000 ;
	    RECT 1105.8000 623.7000 1112.7001 624.6000 ;
	    RECT 1117.8000 623.7000 1121.7001 624.9000 ;
	    RECT 1122.6000 623.7000 1123.8000 629.7000 ;
	    RECT 1105.8000 623.4000 1107.0000 623.7000 ;
	    RECT 1081.2001 618.0000 1082.1000 621.0000 ;
	    RECT 1087.5000 620.1000 1088.7001 621.9000 ;
	    RECT 1083.0000 618.9000 1088.7001 620.1000 ;
	    RECT 1096.2001 619.2000 1097.4000 623.4000 ;
	    RECT 1108.2001 622.5000 1109.4000 622.8000 ;
	    RECT 1105.8000 622.2000 1107.0000 622.5000 ;
	    RECT 1100.4000 621.3000 1107.0000 622.2000 ;
	    RECT 1100.4000 621.0000 1101.6000 621.3000 ;
	    RECT 1108.2001 620.4000 1109.4000 621.6000 ;
	    RECT 1111.5000 620.1000 1112.7001 623.7000 ;
	    RECT 1120.5000 622.8000 1121.7001 623.7000 ;
	    RECT 1120.5000 621.6000 1125.0000 622.8000 ;
	    RECT 1127.4000 620.7000 1128.6000 629.7000 ;
	    RECT 1146.6000 626.7000 1147.8000 629.7000 ;
	    RECT 1146.6000 625.5000 1147.8000 625.8000 ;
	    RECT 1146.6000 623.4000 1147.8000 624.6000 ;
	    RECT 1149.0000 622.5000 1150.2001 629.7000 ;
	    RECT 1101.0000 618.9000 1105.8000 620.1000 ;
	    RECT 1111.5000 618.9000 1114.5000 620.1000 ;
	    RECT 1115.4000 619.5000 1128.6000 620.7000 ;
	    RECT 1149.0000 621.4500 1150.2001 621.6000 ;
	    RECT 1173.0000 621.4500 1174.2001 621.6000 ;
	    RECT 1149.0000 620.5500 1174.2001 621.4500 ;
	    RECT 1175.4000 620.7000 1176.6000 629.7000 ;
	    RECT 1180.8000 621.3000 1182.0000 629.7000 ;
	    RECT 1207.5000 623.7000 1208.7001 629.7000 ;
	    RECT 1211.4000 623.7000 1212.6000 629.7000 ;
	    RECT 1213.8000 626.7000 1215.0000 629.7000 ;
	    RECT 1213.5000 625.5000 1214.7001 625.8000 ;
	    RECT 1180.8000 620.7000 1183.5000 621.3000 ;
	    RECT 1149.0000 620.4000 1150.2001 620.5500 ;
	    RECT 1173.0000 620.4000 1174.2001 620.5500 ;
	    RECT 1181.1000 620.4000 1183.5000 620.7000 ;
	    RECT 1209.0000 620.4000 1210.2001 621.6000 ;
	    RECT 1091.4000 618.0000 1092.6000 618.9000 ;
	    RECT 1081.2001 617.1000 1082.4000 618.0000 ;
	    RECT 1091.4000 617.1000 1116.9000 618.0000 ;
	    RECT 1117.8000 617.4000 1119.0000 618.6000 ;
	    RECT 1125.3000 618.0000 1126.5000 618.3000 ;
	    RECT 1119.9000 617.1000 1126.5000 618.0000 ;
	    RECT 1079.1000 615.0000 1080.6000 616.2000 ;
	    RECT 1079.4000 613.5000 1080.6000 615.0000 ;
	    RECT 1081.5000 614.4000 1082.4000 617.1000 ;
	    RECT 1083.3000 616.2000 1084.5000 616.5000 ;
	    RECT 1083.3000 615.3000 1121.7001 616.2000 ;
	    RECT 1117.5000 615.0000 1118.7001 615.3000 ;
	    RECT 1122.6000 614.4000 1123.8000 615.6000 ;
	    RECT 1081.5000 613.5000 1095.0000 614.4000 ;
	    RECT 1036.2001 612.4500 1037.4000 612.6000 ;
	    RECT 1079.4000 612.4500 1080.6000 612.6000 ;
	    RECT 1036.2001 611.5500 1080.6000 612.4500 ;
	    RECT 1036.2001 611.4000 1037.4000 611.5500 ;
	    RECT 1079.4000 611.4000 1080.6000 611.5500 ;
	    RECT 1081.5000 611.1000 1082.4000 613.5000 ;
	    RECT 1093.8000 613.2000 1095.0000 613.5000 ;
	    RECT 1098.6000 613.5000 1111.5000 614.4000 ;
	    RECT 1098.6000 613.2000 1099.8000 613.5000 ;
	    RECT 1086.3000 611.4000 1090.2001 612.6000 ;
	    RECT 1077.0000 603.3000 1078.2001 609.3000 ;
	    RECT 1079.4000 603.3000 1080.6000 610.5000 ;
	    RECT 1081.5000 610.2000 1085.4000 611.1000 ;
	    RECT 1081.8000 603.3000 1083.0000 609.3000 ;
	    RECT 1084.2001 603.3000 1085.4000 610.2000 ;
	    RECT 1086.6000 603.3000 1087.8000 609.3000 ;
	    RECT 1089.0000 603.3000 1090.2001 611.4000 ;
	    RECT 1091.1000 610.2000 1097.4000 611.4000 ;
	    RECT 1091.4000 603.3000 1092.6000 609.3000 ;
	    RECT 1093.8000 603.3000 1095.0000 607.5000 ;
	    RECT 1096.2001 603.3000 1097.4000 607.5000 ;
	    RECT 1098.6000 603.3000 1099.8000 607.5000 ;
	    RECT 1101.0000 603.3000 1102.2001 612.6000 ;
	    RECT 1105.8000 611.4000 1109.7001 612.6000 ;
	    RECT 1110.6000 612.3000 1111.5000 613.5000 ;
	    RECT 1113.0000 614.1000 1114.2001 614.4000 ;
	    RECT 1113.0000 613.5000 1121.1000 614.1000 ;
	    RECT 1113.0000 613.2000 1122.3000 613.5000 ;
	    RECT 1120.2001 612.3000 1122.3000 613.2000 ;
	    RECT 1110.6000 611.4000 1119.3000 612.3000 ;
	    RECT 1123.8000 612.0000 1126.2001 613.2000 ;
	    RECT 1123.8000 611.4000 1124.7001 612.0000 ;
	    RECT 1103.4000 603.3000 1104.6000 609.3000 ;
	    RECT 1105.8000 603.3000 1107.0000 610.5000 ;
	    RECT 1108.2001 603.3000 1109.4000 609.3000 ;
	    RECT 1110.6000 603.3000 1111.8000 610.5000 ;
	    RECT 1118.4000 610.2000 1124.7001 611.4000 ;
	    RECT 1127.4000 611.1000 1128.6000 619.5000 ;
	    RECT 1125.6000 610.2000 1128.6000 611.1000 ;
	    RECT 1113.0000 603.3000 1114.2001 607.5000 ;
	    RECT 1115.4000 603.3000 1116.6000 607.5000 ;
	    RECT 1117.8000 603.3000 1119.0000 609.3000 ;
	    RECT 1120.2001 603.3000 1121.4000 610.2000 ;
	    RECT 1125.6000 609.3000 1126.5000 610.2000 ;
	    RECT 1122.6000 602.4000 1123.8000 609.3000 ;
	    RECT 1125.0000 608.4000 1126.5000 609.3000 ;
	    RECT 1125.0000 603.3000 1126.2001 608.4000 ;
	    RECT 1127.4000 603.3000 1128.6000 609.3000 ;
	    RECT 1146.6000 603.3000 1147.8000 609.3000 ;
	    RECT 1149.0000 603.3000 1150.2001 619.5000 ;
	    RECT 1177.8000 617.4000 1179.0000 618.6000 ;
	    RECT 1179.9000 617.4000 1180.2001 618.6000 ;
	    RECT 1175.4000 616.5000 1176.6000 616.8000 ;
	    RECT 1182.6000 616.5000 1183.5000 620.4000 ;
	    RECT 1209.0000 619.2000 1210.2001 619.5000 ;
	    RECT 1206.6000 617.4000 1207.8000 618.6000 ;
	    RECT 1211.4000 618.3000 1212.3000 623.7000 ;
	    RECT 1213.8000 623.4000 1215.0000 624.6000 ;
	    RECT 1225.8000 622.5000 1227.0000 629.7000 ;
	    RECT 1228.2001 626.7000 1229.4000 629.7000 ;
	    RECT 1228.2001 625.5000 1229.4000 625.8000 ;
	    RECT 1248.3000 624.6000 1249.5000 629.7000 ;
	    RECT 1228.2001 623.4000 1229.4000 624.6000 ;
	    RECT 1248.3000 623.7000 1251.0000 624.6000 ;
	    RECT 1252.2001 623.7000 1253.4000 629.7000 ;
	    RECT 1279.5000 623.7000 1280.7001 629.7000 ;
	    RECT 1283.4000 623.7000 1284.6000 629.7000 ;
	    RECT 1285.8000 626.7000 1287.0000 629.7000 ;
	    RECT 1285.5000 625.5000 1286.7001 625.8000 ;
	    RECT 1285.8000 624.4500 1287.0000 624.6000 ;
	    RECT 1302.6000 624.4500 1303.8000 624.6000 ;
	    RECT 1213.8000 621.4500 1215.0000 621.6000 ;
	    RECT 1225.8000 621.4500 1227.0000 621.6000 ;
	    RECT 1213.8000 620.5500 1227.0000 621.4500 ;
	    RECT 1213.8000 620.4000 1215.0000 620.5500 ;
	    RECT 1225.8000 620.4000 1227.0000 620.5500 ;
	    RECT 1249.8000 619.5000 1251.0000 623.7000 ;
	    RECT 1252.2001 622.5000 1253.4000 622.8000 ;
	    RECT 1252.2001 621.4500 1253.4000 621.6000 ;
	    RECT 1276.2001 621.4500 1277.4000 621.6000 ;
	    RECT 1252.2001 620.5500 1277.4000 621.4500 ;
	    RECT 1252.2001 620.4000 1253.4000 620.5500 ;
	    RECT 1276.2001 620.4000 1277.4000 620.5500 ;
	    RECT 1281.0000 620.4000 1282.2001 621.6000 ;
	    RECT 1213.8000 618.4500 1215.0000 618.6000 ;
	    RECT 1223.4000 618.4500 1224.6000 618.6000 ;
	    RECT 1208.7001 616.8000 1209.0000 618.3000 ;
	    RECT 1211.4000 617.4000 1212.9000 618.3000 ;
	    RECT 1213.8000 617.5500 1224.6000 618.4500 ;
	    RECT 1213.8000 617.4000 1215.0000 617.5500 ;
	    RECT 1223.4000 617.4000 1224.6000 617.5500 ;
	    RECT 1175.4000 614.4000 1176.6000 615.6000 ;
	    RECT 1182.6000 615.4500 1183.8000 615.6000 ;
	    RECT 1204.2001 615.4500 1205.4000 615.6000 ;
	    RECT 1182.6000 614.5500 1205.4000 615.4500 ;
	    RECT 1213.8000 615.3000 1214.7001 616.5000 ;
	    RECT 1182.6000 614.4000 1183.8000 614.5500 ;
	    RECT 1204.2001 614.4000 1205.4000 614.5500 ;
	    RECT 1206.6000 614.4000 1212.6000 615.3000 ;
	    RECT 1180.2001 613.5000 1181.4000 613.8000 ;
	    RECT 1177.8000 612.4500 1179.0000 612.6000 ;
	    RECT 1180.2001 612.4500 1181.4000 612.6000 ;
	    RECT 1177.8000 611.5500 1181.4000 612.4500 ;
	    RECT 1177.8000 611.4000 1179.0000 611.5500 ;
	    RECT 1180.2001 611.4000 1181.4000 611.5500 ;
	    RECT 1182.6000 610.5000 1183.5000 613.5000 ;
	    RECT 1178.1000 609.6000 1183.5000 610.5000 ;
	    RECT 1178.1000 609.3000 1179.0000 609.6000 ;
	    RECT 1175.4000 603.3000 1176.6000 609.3000 ;
	    RECT 1177.8000 603.3000 1179.0000 609.3000 ;
	    RECT 1182.6000 609.3000 1183.5000 609.6000 ;
	    RECT 1180.2001 603.3000 1181.4000 608.7000 ;
	    RECT 1182.6000 603.3000 1183.8000 609.3000 ;
	    RECT 1206.6000 603.3000 1207.8000 614.4000 ;
	    RECT 1209.0000 603.3000 1210.2001 613.5000 ;
	    RECT 1211.4000 603.3000 1212.6000 614.4000 ;
	    RECT 1213.8000 603.3000 1215.0000 615.3000 ;
	    RECT 1225.8000 603.3000 1227.0000 619.5000 ;
	    RECT 1281.0000 619.2000 1282.2001 619.5000 ;
	    RECT 1228.2001 618.4500 1229.4000 618.6000 ;
	    RECT 1242.6000 618.4500 1243.8000 618.6000 ;
	    RECT 1249.8000 618.4500 1251.0000 618.6000 ;
	    RECT 1228.2001 617.5500 1251.0000 618.4500 ;
	    RECT 1228.2001 617.4000 1229.4000 617.5500 ;
	    RECT 1242.6000 617.4000 1243.8000 617.5500 ;
	    RECT 1249.8000 617.4000 1251.0000 617.5500 ;
	    RECT 1278.6000 617.4000 1279.8000 618.6000 ;
	    RECT 1283.4000 618.3000 1284.3000 623.7000 ;
	    RECT 1285.8000 623.5500 1303.8000 624.4500 ;
	    RECT 1285.8000 623.4000 1287.0000 623.5500 ;
	    RECT 1302.6000 623.4000 1303.8000 623.5500 ;
	    RECT 1309.8000 620.7000 1311.0000 629.7000 ;
	    RECT 1315.2001 621.3000 1316.4000 629.7000 ;
	    RECT 1341.0000 626.7000 1342.2001 629.7000 ;
	    RECT 1341.3000 625.5000 1342.5000 625.8000 ;
	    RECT 1341.0000 623.4000 1342.2001 624.6000 ;
	    RECT 1343.4000 623.7000 1344.6000 629.7000 ;
	    RECT 1347.3000 623.7000 1348.5000 629.7000 ;
	    RECT 1315.2001 620.7000 1317.9000 621.3000 ;
	    RECT 1315.5000 620.4000 1317.9000 620.7000 ;
	    RECT 1285.8000 618.4500 1287.0000 618.6000 ;
	    RECT 1305.0000 618.4500 1306.2001 618.6000 ;
	    RECT 1280.7001 616.8000 1281.0000 618.3000 ;
	    RECT 1283.4000 617.4000 1284.9000 618.3000 ;
	    RECT 1285.8000 617.5500 1306.2001 618.4500 ;
	    RECT 1285.8000 617.4000 1287.0000 617.5500 ;
	    RECT 1305.0000 617.4000 1306.2001 617.5500 ;
	    RECT 1312.2001 617.4000 1313.4000 618.6000 ;
	    RECT 1314.3000 617.4000 1314.6000 618.6000 ;
	    RECT 1309.8000 616.5000 1311.0000 616.8000 ;
	    RECT 1317.0000 616.5000 1317.9000 620.4000 ;
	    RECT 1336.2001 618.4500 1337.4000 618.6000 ;
	    RECT 1341.0000 618.4500 1342.2001 618.6000 ;
	    RECT 1336.2001 617.5500 1342.2001 618.4500 ;
	    RECT 1343.7001 618.3000 1344.6000 623.7000 ;
	    RECT 1345.8000 620.4000 1347.0000 621.6000 ;
	    RECT 1379.4000 620.7000 1380.6000 629.7000 ;
	    RECT 1384.8000 621.3000 1386.0000 629.7000 ;
	    RECT 1389.0000 621.4500 1390.2001 621.6000 ;
	    RECT 1398.6000 621.4500 1399.8000 621.6000 ;
	    RECT 1384.8000 620.7000 1387.5000 621.3000 ;
	    RECT 1385.1000 620.4000 1387.5000 620.7000 ;
	    RECT 1389.0000 620.5500 1399.8000 621.4500 ;
	    RECT 1413.0000 620.7000 1414.2001 629.7000 ;
	    RECT 1418.4000 621.3000 1419.6000 629.7000 ;
	    RECT 1473.0000 626.7000 1474.2001 629.7000 ;
	    RECT 1475.4000 627.3000 1476.6000 629.7000 ;
	    RECT 1477.8000 627.6000 1479.0000 629.7000 ;
	    RECT 1472.4000 626.4000 1474.2001 626.7000 ;
	    RECT 1477.5000 626.7000 1479.0000 627.6000 ;
	    RECT 1480.2001 626.7000 1481.4000 629.7000 ;
	    RECT 1477.5000 626.4000 1478.4000 626.7000 ;
	    RECT 1472.4000 625.5000 1478.4000 626.4000 ;
	    RECT 1418.4000 620.7000 1421.1000 621.3000 ;
	    RECT 1389.0000 620.4000 1390.2001 620.5500 ;
	    RECT 1398.6000 620.4000 1399.8000 620.5500 ;
	    RECT 1418.7001 620.4000 1421.1000 620.7000 ;
	    RECT 1345.8000 619.2000 1347.0000 619.5000 ;
	    RECT 1336.2001 617.4000 1337.4000 617.5500 ;
	    RECT 1341.0000 617.4000 1342.2001 617.5500 ;
	    RECT 1343.1000 617.4000 1344.6000 618.3000 ;
	    RECT 1347.0000 616.8000 1347.3000 618.3000 ;
	    RECT 1348.2001 617.4000 1349.4000 618.6000 ;
	    RECT 1381.8000 617.4000 1383.0000 618.6000 ;
	    RECT 1383.9000 617.4000 1384.2001 618.6000 ;
	    RECT 1379.4000 616.5000 1380.6000 616.8000 ;
	    RECT 1386.6000 616.5000 1387.5000 620.4000 ;
	    RECT 1415.4000 617.4000 1416.6000 618.6000 ;
	    RECT 1417.5000 617.4000 1417.8000 618.6000 ;
	    RECT 1413.0000 616.5000 1414.2001 616.8000 ;
	    RECT 1420.2001 616.5000 1421.1000 620.4000 ;
	    RECT 1247.4000 614.4000 1248.6000 615.6000 ;
	    RECT 1247.4000 613.2000 1248.6000 613.5000 ;
	    RECT 1228.2001 603.3000 1229.4000 609.3000 ;
	    RECT 1247.4000 603.3000 1248.6000 609.3000 ;
	    RECT 1249.8000 603.3000 1251.0000 616.5000 ;
	    RECT 1285.8000 615.3000 1286.7001 616.5000 ;
	    RECT 1300.2001 615.4500 1301.4000 615.6000 ;
	    RECT 1309.8000 615.4500 1311.0000 615.6000 ;
	    RECT 1278.6000 614.4000 1284.6000 615.3000 ;
	    RECT 1252.2001 603.3000 1253.4000 609.3000 ;
	    RECT 1278.6000 603.3000 1279.8000 614.4000 ;
	    RECT 1281.0000 603.3000 1282.2001 613.5000 ;
	    RECT 1283.4000 603.3000 1284.6000 614.4000 ;
	    RECT 1285.8000 603.3000 1287.0000 615.3000 ;
	    RECT 1300.2001 614.5500 1311.0000 615.4500 ;
	    RECT 1300.2001 614.4000 1301.4000 614.5500 ;
	    RECT 1309.8000 614.4000 1311.0000 614.5500 ;
	    RECT 1317.0000 615.4500 1318.2001 615.6000 ;
	    RECT 1338.6000 615.4500 1339.8000 615.6000 ;
	    RECT 1317.0000 614.5500 1339.8000 615.4500 ;
	    RECT 1341.3000 615.3000 1342.2001 616.5000 ;
	    RECT 1472.4000 615.6000 1473.3000 625.5000 ;
	    RECT 1478.7001 623.4000 1479.3000 624.6000 ;
	    RECT 1480.2001 623.4000 1481.4000 624.6000 ;
	    RECT 1476.6000 620.4000 1476.9000 621.6000 ;
	    RECT 1477.8000 620.4000 1479.0000 621.6000 ;
	    RECT 1506.6000 620.7000 1507.8000 629.7000 ;
	    RECT 1512.0000 621.3000 1513.2001 629.7000 ;
	    RECT 1542.0000 621.3000 1543.2001 629.7000 ;
	    RECT 1512.0000 620.7000 1514.7001 621.3000 ;
	    RECT 1512.3000 620.4000 1514.7001 620.7000 ;
	    RECT 1474.2001 617.4000 1474.5000 618.6000 ;
	    RECT 1475.4000 617.4000 1476.6000 618.6000 ;
	    RECT 1509.0000 617.4000 1510.2001 618.6000 ;
	    RECT 1511.1000 617.4000 1511.4000 618.6000 ;
	    RECT 1506.6000 616.5000 1507.8000 616.8000 ;
	    RECT 1513.8000 616.5000 1514.7001 620.4000 ;
	    RECT 1540.5000 620.7000 1543.2001 621.3000 ;
	    RECT 1547.4000 620.7000 1548.6000 629.7000 ;
	    RECT 1540.5000 620.4000 1542.9000 620.7000 ;
	    RECT 1540.5000 616.5000 1541.4000 620.4000 ;
	    RECT 1543.8000 617.4000 1544.1000 618.6000 ;
	    RECT 1545.0000 617.4000 1546.2001 618.6000 ;
	    RECT 1547.4000 616.5000 1548.6000 616.8000 ;
	    RECT 1369.8000 615.4500 1371.0000 615.6000 ;
	    RECT 1379.4000 615.4500 1380.6000 615.6000 ;
	    RECT 1317.0000 614.4000 1318.2001 614.5500 ;
	    RECT 1338.6000 614.4000 1339.8000 614.5500 ;
	    RECT 1314.6000 613.5000 1315.8000 613.8000 ;
	    RECT 1302.6000 612.4500 1303.8000 612.6000 ;
	    RECT 1314.6000 612.4500 1315.8000 612.6000 ;
	    RECT 1302.6000 611.5500 1315.8000 612.4500 ;
	    RECT 1302.6000 611.4000 1303.8000 611.5500 ;
	    RECT 1314.6000 611.4000 1315.8000 611.5500 ;
	    RECT 1317.0000 610.5000 1317.9000 613.5000 ;
	    RECT 1312.5000 609.6000 1317.9000 610.5000 ;
	    RECT 1312.5000 609.3000 1313.4000 609.6000 ;
	    RECT 1309.8000 603.3000 1311.0000 609.3000 ;
	    RECT 1312.2001 603.3000 1313.4000 609.3000 ;
	    RECT 1317.0000 609.3000 1317.9000 609.6000 ;
	    RECT 1314.6000 603.3000 1315.8000 608.7000 ;
	    RECT 1317.0000 603.3000 1318.2001 609.3000 ;
	    RECT 1341.0000 603.3000 1342.2001 615.3000 ;
	    RECT 1343.4000 614.4000 1349.4000 615.3000 ;
	    RECT 1369.8000 614.5500 1380.6000 615.4500 ;
	    RECT 1369.8000 614.4000 1371.0000 614.5500 ;
	    RECT 1379.4000 614.4000 1380.6000 614.5500 ;
	    RECT 1386.6000 615.4500 1387.8000 615.6000 ;
	    RECT 1408.2001 615.4500 1409.4000 615.6000 ;
	    RECT 1386.6000 614.5500 1409.4000 615.4500 ;
	    RECT 1386.6000 614.4000 1387.8000 614.5500 ;
	    RECT 1408.2001 614.4000 1409.4000 614.5500 ;
	    RECT 1413.0000 615.4500 1414.2001 615.6000 ;
	    RECT 1415.4000 615.4500 1416.6000 615.6000 ;
	    RECT 1413.0000 614.5500 1416.6000 615.4500 ;
	    RECT 1413.0000 614.4000 1414.2001 614.5500 ;
	    RECT 1415.4000 614.4000 1416.6000 614.5500 ;
	    RECT 1420.2001 615.4500 1421.4000 615.6000 ;
	    RECT 1427.4000 615.4500 1428.6000 615.6000 ;
	    RECT 1420.2001 614.5500 1428.6000 615.4500 ;
	    RECT 1420.2001 614.4000 1421.4000 614.5500 ;
	    RECT 1427.4000 614.4000 1428.6000 614.5500 ;
	    RECT 1437.0000 615.4500 1438.2001 615.6000 ;
	    RECT 1468.2001 615.4500 1469.4000 615.6000 ;
	    RECT 1437.0000 614.5500 1469.4000 615.4500 ;
	    RECT 1470.3000 614.7000 1473.3000 615.6000 ;
	    RECT 1497.0000 615.4500 1498.2001 615.6000 ;
	    RECT 1506.6000 615.4500 1507.8000 615.6000 ;
	    RECT 1437.0000 614.4000 1438.2001 614.5500 ;
	    RECT 1468.2001 614.4000 1469.4000 614.5500 ;
	    RECT 1497.0000 614.5500 1507.8000 615.4500 ;
	    RECT 1497.0000 614.4000 1498.2001 614.5500 ;
	    RECT 1506.6000 614.4000 1507.8000 614.5500 ;
	    RECT 1513.8000 615.4500 1515.0000 615.6000 ;
	    RECT 1518.6000 615.4500 1519.8000 615.6000 ;
	    RECT 1513.8000 614.5500 1519.8000 615.4500 ;
	    RECT 1513.8000 614.4000 1515.0000 614.5500 ;
	    RECT 1518.6000 614.4000 1519.8000 614.5500 ;
	    RECT 1521.0000 615.4500 1522.2001 615.6000 ;
	    RECT 1540.2001 615.4500 1541.4000 615.6000 ;
	    RECT 1521.0000 614.5500 1541.4000 615.4500 ;
	    RECT 1521.0000 614.4000 1522.2001 614.5500 ;
	    RECT 1540.2001 614.4000 1541.4000 614.5500 ;
	    RECT 1547.4000 614.4000 1548.6000 615.6000 ;
	    RECT 1343.4000 603.3000 1344.6000 614.4000 ;
	    RECT 1345.8000 603.3000 1347.0000 613.5000 ;
	    RECT 1348.2001 603.3000 1349.4000 614.4000 ;
	    RECT 1384.2001 613.5000 1385.4000 613.8000 ;
	    RECT 1417.8000 613.5000 1419.0000 613.8000 ;
	    RECT 1470.9000 613.5000 1476.3000 613.8000 ;
	    RECT 1384.2001 611.4000 1385.4000 612.6000 ;
	    RECT 1386.6000 610.5000 1387.5000 613.5000 ;
	    RECT 1417.8000 611.4000 1419.0000 612.6000 ;
	    RECT 1420.2001 610.5000 1421.1000 613.5000 ;
	    RECT 1382.1000 609.6000 1387.5000 610.5000 ;
	    RECT 1382.1000 609.3000 1383.0000 609.6000 ;
	    RECT 1379.4000 603.3000 1380.6000 609.3000 ;
	    RECT 1381.8000 603.3000 1383.0000 609.3000 ;
	    RECT 1386.6000 609.3000 1387.5000 609.6000 ;
	    RECT 1415.7001 609.6000 1421.1000 610.5000 ;
	    RECT 1415.7001 609.3000 1416.6000 609.6000 ;
	    RECT 1384.2001 603.3000 1385.4000 608.7000 ;
	    RECT 1386.6000 603.3000 1387.8000 609.3000 ;
	    RECT 1413.0000 603.3000 1414.2001 609.3000 ;
	    RECT 1415.4000 603.3000 1416.6000 609.3000 ;
	    RECT 1420.2001 609.3000 1421.1000 609.6000 ;
	    RECT 1417.8000 603.3000 1419.0000 608.7000 ;
	    RECT 1420.2001 603.3000 1421.4000 609.3000 ;
	    RECT 1465.8000 604.5000 1467.0000 613.5000 ;
	    RECT 1468.2001 605.1000 1469.4000 613.5000 ;
	    RECT 1470.6000 612.9000 1476.3000 613.5000 ;
	    RECT 1466.1000 604.2000 1467.0000 604.5000 ;
	    RECT 1470.6000 604.5000 1471.8000 612.9000 ;
	    RECT 1475.4000 612.3000 1476.3000 612.9000 ;
	    RECT 1478.1000 613.2000 1483.5000 614.1000 ;
	    RECT 1511.4000 613.5000 1512.6000 613.8000 ;
	    RECT 1542.6000 613.5000 1543.8000 613.8000 ;
	    RECT 1478.1000 612.3000 1479.0000 613.2000 ;
	    RECT 1482.6000 612.3000 1483.5000 613.2000 ;
	    RECT 1485.0000 612.4500 1486.2001 612.6000 ;
	    RECT 1511.4000 612.4500 1512.6000 612.6000 ;
	    RECT 1470.6000 604.2000 1471.5000 604.5000 ;
	    RECT 1466.1000 603.3000 1471.5000 604.2000 ;
	    RECT 1473.0000 604.2000 1474.2001 612.0000 ;
	    RECT 1475.4000 605.1000 1476.6000 612.3000 ;
	    RECT 1477.8000 604.2000 1479.0000 612.3000 ;
	    RECT 1473.0000 603.3000 1479.0000 604.2000 ;
	    RECT 1480.2001 603.3000 1481.4000 612.3000 ;
	    RECT 1482.6000 603.3000 1483.8000 612.3000 ;
	    RECT 1485.0000 611.5500 1512.6000 612.4500 ;
	    RECT 1485.0000 611.4000 1486.2001 611.5500 ;
	    RECT 1511.4000 611.4000 1512.6000 611.5500 ;
	    RECT 1513.8000 610.5000 1514.7001 613.5000 ;
	    RECT 1509.3000 609.6000 1514.7001 610.5000 ;
	    RECT 1509.3000 609.3000 1510.2001 609.6000 ;
	    RECT 1506.6000 603.3000 1507.8000 609.3000 ;
	    RECT 1509.0000 603.3000 1510.2001 609.3000 ;
	    RECT 1513.8000 609.3000 1514.7001 609.6000 ;
	    RECT 1540.5000 610.5000 1541.4000 613.5000 ;
	    RECT 1542.6000 611.4000 1543.8000 612.6000 ;
	    RECT 1540.5000 609.6000 1545.9000 610.5000 ;
	    RECT 1540.5000 609.3000 1541.4000 609.6000 ;
	    RECT 1511.4000 603.3000 1512.6000 608.7000 ;
	    RECT 1513.8000 603.3000 1515.0000 609.3000 ;
	    RECT 1540.2001 603.3000 1541.4000 609.3000 ;
	    RECT 1545.0000 609.3000 1545.9000 609.6000 ;
	    RECT 1542.6000 603.3000 1543.8000 608.7000 ;
	    RECT 1545.0000 603.3000 1546.2001 609.3000 ;
	    RECT 1547.4000 603.3000 1548.6000 609.3000 ;
	    RECT 1.2000 600.6000 1569.0000 602.4000 ;
	    RECT 126.6000 593.7000 127.8000 599.7000 ;
	    RECT 129.0000 594.6000 130.2000 599.7000 ;
	    RECT 128.7000 593.7000 130.2000 594.6000 ;
	    RECT 131.4000 593.7000 132.6000 600.6000 ;
	    RECT 128.7000 592.8000 129.6000 593.7000 ;
	    RECT 133.8000 592.8000 135.0000 599.7000 ;
	    RECT 136.2000 593.7000 137.4000 599.7000 ;
	    RECT 138.6000 595.5000 139.8000 599.7000 ;
	    RECT 141.0000 595.5000 142.2000 599.7000 ;
	    RECT 126.6000 591.9000 129.6000 592.8000 ;
	    RECT 126.6000 583.5000 127.8000 591.9000 ;
	    RECT 130.5000 591.6000 136.8000 592.8000 ;
	    RECT 143.4000 592.5000 144.6000 599.7000 ;
	    RECT 145.8000 593.7000 147.0000 599.7000 ;
	    RECT 148.2000 592.5000 149.4000 599.7000 ;
	    RECT 150.6000 593.7000 151.8000 599.7000 ;
	    RECT 130.5000 591.0000 131.4000 591.6000 ;
	    RECT 129.0000 589.8000 131.4000 591.0000 ;
	    RECT 135.9000 590.7000 144.6000 591.6000 ;
	    RECT 132.9000 589.8000 135.0000 590.7000 ;
	    RECT 132.9000 589.5000 142.2000 589.8000 ;
	    RECT 134.1000 588.9000 142.2000 589.5000 ;
	    RECT 141.0000 588.6000 142.2000 588.9000 ;
	    RECT 143.7000 589.5000 144.6000 590.7000 ;
	    RECT 145.5000 590.4000 149.4000 591.6000 ;
	    RECT 153.0000 590.4000 154.2000 599.7000 ;
	    RECT 155.4000 595.5000 156.6000 599.7000 ;
	    RECT 157.8000 595.5000 159.0000 599.7000 ;
	    RECT 160.2000 595.5000 161.4000 599.7000 ;
	    RECT 162.6000 593.7000 163.8000 599.7000 ;
	    RECT 157.8000 591.6000 164.1000 592.8000 ;
	    RECT 165.0000 591.6000 166.2000 599.7000 ;
	    RECT 167.4000 593.7000 168.6000 599.7000 ;
	    RECT 169.8000 592.8000 171.0000 599.7000 ;
	    RECT 172.2000 593.7000 173.4000 599.7000 ;
	    RECT 169.8000 591.9000 173.7000 592.8000 ;
	    RECT 174.6000 592.5000 175.8000 599.7000 ;
	    RECT 177.0000 593.7000 178.2000 599.7000 ;
	    RECT 165.0000 590.4000 168.9000 591.6000 ;
	    RECT 155.4000 589.5000 156.6000 589.8000 ;
	    RECT 143.7000 588.6000 156.6000 589.5000 ;
	    RECT 160.2000 589.5000 161.4000 589.8000 ;
	    RECT 172.8000 589.5000 173.7000 591.9000 ;
	    RECT 174.6000 590.4000 175.8000 591.6000 ;
	    RECT 160.2000 588.6000 173.7000 589.5000 ;
	    RECT 131.4000 587.4000 132.6000 588.6000 ;
	    RECT 136.5000 587.7000 137.7000 588.0000 ;
	    RECT 133.5000 586.8000 171.9000 587.7000 ;
	    RECT 170.7000 586.5000 171.9000 586.8000 ;
	    RECT 172.8000 585.9000 173.7000 588.6000 ;
	    RECT 174.6000 588.0000 175.8000 589.5000 ;
	    RECT 174.6000 586.8000 176.1000 588.0000 ;
	    RECT 128.7000 585.0000 135.3000 585.9000 ;
	    RECT 128.7000 584.7000 129.9000 585.0000 ;
	    RECT 136.2000 584.4000 137.4000 585.6000 ;
	    RECT 138.3000 585.0000 163.8000 585.9000 ;
	    RECT 172.8000 585.0000 174.0000 585.9000 ;
	    RECT 162.6000 584.1000 163.8000 585.0000 ;
	    RECT 126.6000 582.3000 139.8000 583.5000 ;
	    RECT 140.7000 582.9000 143.7000 584.1000 ;
	    RECT 149.4000 582.9000 154.2000 584.1000 ;
	    RECT 126.6000 573.3000 127.8000 582.3000 ;
	    RECT 130.2000 580.2000 134.7000 581.4000 ;
	    RECT 133.5000 579.3000 134.7000 580.2000 ;
	    RECT 142.5000 579.3000 143.7000 582.9000 ;
	    RECT 145.8000 581.4000 147.0000 582.6000 ;
	    RECT 153.6000 581.7000 154.8000 582.0000 ;
	    RECT 148.2000 580.8000 154.8000 581.7000 ;
	    RECT 148.2000 580.5000 149.4000 580.8000 ;
	    RECT 145.8000 580.2000 147.0000 580.5000 ;
	    RECT 157.8000 579.6000 159.0000 583.8000 ;
	    RECT 166.5000 582.9000 172.2000 584.1000 ;
	    RECT 166.5000 581.1000 167.7000 582.9000 ;
	    RECT 173.1000 582.0000 174.0000 585.0000 ;
	    RECT 148.2000 579.3000 149.4000 579.6000 ;
	    RECT 131.4000 573.3000 132.6000 579.3000 ;
	    RECT 133.5000 578.1000 137.4000 579.3000 ;
	    RECT 142.5000 578.4000 149.4000 579.3000 ;
	    RECT 150.6000 578.4000 151.8000 579.6000 ;
	    RECT 152.7000 578.4000 153.0000 579.6000 ;
	    RECT 157.5000 578.4000 159.0000 579.6000 ;
	    RECT 165.0000 580.2000 167.7000 581.1000 ;
	    RECT 172.2000 581.1000 174.0000 582.0000 ;
	    RECT 165.0000 579.3000 166.2000 580.2000 ;
	    RECT 136.2000 573.3000 137.4000 578.1000 ;
	    RECT 162.6000 578.1000 166.2000 579.3000 ;
	    RECT 138.6000 573.3000 139.8000 577.5000 ;
	    RECT 141.0000 573.3000 142.2000 577.5000 ;
	    RECT 143.4000 573.3000 144.6000 577.5000 ;
	    RECT 145.8000 573.3000 147.0000 576.3000 ;
	    RECT 148.2000 573.3000 149.4000 577.5000 ;
	    RECT 150.6000 573.3000 151.8000 576.3000 ;
	    RECT 153.0000 573.3000 154.2000 577.5000 ;
	    RECT 155.4000 573.3000 156.6000 577.5000 ;
	    RECT 157.8000 573.3000 159.0000 577.5000 ;
	    RECT 160.2000 573.3000 161.4000 577.5000 ;
	    RECT 162.6000 573.3000 163.8000 578.1000 ;
	    RECT 167.4000 573.3000 168.6000 579.3000 ;
	    RECT 172.2000 573.3000 173.4000 581.1000 ;
	    RECT 174.9000 580.2000 176.1000 586.8000 ;
	    RECT 191.4000 583.5000 192.6000 599.7000 ;
	    RECT 193.8000 593.7000 195.0000 599.7000 ;
	    RECT 213.0000 583.5000 214.2000 599.7000 ;
	    RECT 215.4000 593.7000 216.6000 599.7000 ;
	    RECT 246.6000 587.7000 247.8000 599.7000 ;
	    RECT 250.5000 587.7000 253.5000 599.7000 ;
	    RECT 256.2000 587.7000 257.4000 599.7000 ;
	    RECT 261.1500 597.4500 262.0500 600.6000 ;
	    RECT 270.6000 597.4500 271.8000 597.6000 ;
	    RECT 261.1500 596.5500 271.8000 597.4500 ;
	    RECT 270.6000 596.4000 271.8000 596.5500 ;
	    RECT 275.4000 593.7000 276.6000 599.7000 ;
	    RECT 258.6000 591.4500 259.8000 591.6000 ;
	    RECT 268.2000 591.4500 269.4000 591.6000 ;
	    RECT 258.6000 590.5500 269.4000 591.4500 ;
	    RECT 258.6000 590.4000 259.8000 590.5500 ;
	    RECT 268.2000 590.4000 269.4000 590.5500 ;
	    RECT 232.2000 585.4500 233.4000 585.6000 ;
	    RECT 249.0000 585.4500 250.2000 585.6000 ;
	    RECT 232.2000 584.5500 250.2000 585.4500 ;
	    RECT 232.2000 584.4000 233.4000 584.5500 ;
	    RECT 249.0000 584.4000 250.2000 584.5500 ;
	    RECT 251.4000 583.5000 252.3000 587.7000 ;
	    RECT 277.8000 586.5000 279.0000 599.7000 ;
	    RECT 280.2000 593.7000 281.4000 599.7000 ;
	    RECT 299.4000 593.7000 300.6000 599.7000 ;
	    RECT 280.2000 589.5000 281.4000 589.8000 ;
	    RECT 280.2000 587.4000 281.4000 588.6000 ;
	    RECT 301.8000 586.5000 303.0000 599.7000 ;
	    RECT 304.2000 593.7000 305.4000 599.7000 ;
	    RECT 304.2000 589.5000 305.4000 589.8000 ;
	    RECT 304.2000 588.4500 305.4000 588.6000 ;
	    RECT 306.6000 588.4500 307.8000 588.6000 ;
	    RECT 304.2000 587.5500 307.8000 588.4500 ;
	    RECT 335.4000 587.7000 336.6000 599.7000 ;
	    RECT 339.3000 587.7000 342.3000 599.7000 ;
	    RECT 345.0000 587.7000 346.2000 599.7000 ;
	    RECT 304.2000 587.4000 305.4000 587.5500 ;
	    RECT 306.6000 587.4000 307.8000 587.5500 ;
	    RECT 253.8000 584.4000 255.0000 585.6000 ;
	    RECT 277.8000 584.4000 279.0000 585.6000 ;
	    RECT 280.2000 585.4500 281.4000 585.6000 ;
	    RECT 301.8000 585.4500 303.0000 585.6000 ;
	    RECT 280.2000 584.5500 303.0000 585.4500 ;
	    RECT 280.2000 584.4000 281.4000 584.5500 ;
	    RECT 301.8000 584.4000 303.0000 584.5500 ;
	    RECT 337.8000 584.4000 339.0000 585.6000 ;
	    RECT 256.2000 583.5000 257.4000 583.8000 ;
	    RECT 335.4000 583.5000 336.6000 583.8000 ;
	    RECT 340.5000 583.5000 341.4000 587.7000 ;
	    RECT 342.6000 584.4000 343.8000 585.6000 ;
	    RECT 359.4000 583.5000 360.6000 599.7000 ;
	    RECT 361.8000 593.7000 363.0000 599.7000 ;
	    RECT 364.2000 599.4000 365.4000 600.6000 ;
	    RECT 381.0000 593.7000 382.2000 599.7000 ;
	    RECT 383.4000 586.5000 384.6000 599.7000 ;
	    RECT 385.8000 593.7000 387.0000 599.7000 ;
	    RECT 388.3500 597.4500 389.2500 600.6000 ;
	    RECT 393.0000 597.4500 394.2000 597.6000 ;
	    RECT 388.3500 596.5500 394.2000 597.4500 ;
	    RECT 393.0000 596.4000 394.2000 596.5500 ;
	    RECT 405.0000 593.7000 406.2000 599.7000 ;
	    RECT 385.8000 589.5000 387.0000 589.8000 ;
	    RECT 385.8000 588.4500 387.0000 588.6000 ;
	    RECT 393.0000 588.4500 394.2000 588.6000 ;
	    RECT 385.8000 587.5500 394.2000 588.4500 ;
	    RECT 385.8000 587.4000 387.0000 587.5500 ;
	    RECT 393.0000 587.4000 394.2000 587.5500 ;
	    RECT 407.4000 586.5000 408.6000 599.7000 ;
	    RECT 409.8000 593.7000 411.0000 599.7000 ;
	    RECT 409.8000 589.5000 411.0000 589.8000 ;
	    RECT 409.8000 588.4500 411.0000 588.6000 ;
	    RECT 419.4000 588.4500 420.6000 588.6000 ;
	    RECT 409.8000 587.5500 420.6000 588.4500 ;
	    RECT 409.8000 587.4000 411.0000 587.5500 ;
	    RECT 419.4000 587.4000 420.6000 587.5500 ;
	    RECT 383.4000 585.4500 384.6000 585.6000 ;
	    RECT 405.0000 585.4500 406.2000 585.6000 ;
	    RECT 383.4000 584.5500 406.2000 585.4500 ;
	    RECT 383.4000 584.4000 384.6000 584.5500 ;
	    RECT 405.0000 584.4000 406.2000 584.5500 ;
	    RECT 407.4000 585.4500 408.6000 585.6000 ;
	    RECT 421.8000 585.4500 423.0000 585.6000 ;
	    RECT 407.4000 584.5500 423.0000 585.4500 ;
	    RECT 407.4000 584.4000 408.6000 584.5500 ;
	    RECT 421.8000 584.4000 423.0000 584.5500 ;
	    RECT 424.2000 583.5000 425.4000 599.7000 ;
	    RECT 426.6000 593.7000 427.8000 599.7000 ;
	    RECT 458.7000 593.7000 459.9000 599.7000 ;
	    RECT 459.0000 590.4000 460.2000 591.6000 ;
	    RECT 459.0000 589.5000 459.9000 590.4000 ;
	    RECT 461.1000 588.6000 462.3000 599.7000 ;
	    RECT 457.8000 587.4000 459.0000 588.6000 ;
	    RECT 460.8000 587.7000 462.3000 588.6000 ;
	    RECT 465.0000 587.7000 466.2000 599.7000 ;
	    RECT 489.9000 593.7000 491.1000 599.7000 ;
	    RECT 490.2000 590.4000 491.4000 591.6000 ;
	    RECT 490.2000 589.5000 491.1000 590.4000 ;
	    RECT 492.3000 588.6000 493.5000 599.7000 ;
	    RECT 249.0000 583.2000 250.2000 583.5000 ;
	    RECT 253.8000 583.2000 255.0000 583.5000 ;
	    RECT 177.0000 582.4500 178.2000 582.6000 ;
	    RECT 191.4000 582.4500 192.6000 582.6000 ;
	    RECT 177.0000 581.5500 192.6000 582.4500 ;
	    RECT 177.0000 581.4000 178.2000 581.5500 ;
	    RECT 191.4000 581.4000 192.6000 581.5500 ;
	    RECT 213.0000 582.4500 214.2000 582.6000 ;
	    RECT 222.6000 582.4500 223.8000 582.6000 ;
	    RECT 213.0000 581.5500 223.8000 582.4500 ;
	    RECT 213.0000 581.4000 214.2000 581.5500 ;
	    RECT 222.6000 581.4000 223.8000 581.5500 ;
	    RECT 225.0000 582.4500 226.2000 582.6000 ;
	    RECT 246.6000 582.4500 247.8000 582.6000 ;
	    RECT 225.0000 581.5500 247.8000 582.4500 ;
	    RECT 225.0000 581.4000 226.2000 581.5500 ;
	    RECT 246.6000 581.4000 247.8000 581.5500 ;
	    RECT 248.7000 580.8000 249.0000 582.3000 ;
	    RECT 251.4000 581.4000 252.6000 582.6000 ;
	    RECT 256.2000 582.4500 257.4000 582.6000 ;
	    RECT 258.6000 582.4500 259.8000 582.6000 ;
	    RECT 253.5000 581.4000 255.0000 582.3000 ;
	    RECT 256.2000 581.5500 259.8000 582.4500 ;
	    RECT 256.2000 581.4000 257.4000 581.5500 ;
	    RECT 258.6000 581.4000 259.8000 581.5500 ;
	    RECT 275.4000 581.4000 276.6000 582.6000 ;
	    RECT 174.6000 579.0000 176.1000 580.2000 ;
	    RECT 174.6000 573.3000 175.8000 579.0000 ;
	    RECT 177.0000 573.3000 178.2000 576.3000 ;
	    RECT 191.4000 573.3000 192.6000 580.5000 ;
	    RECT 193.8000 579.4500 195.0000 579.6000 ;
	    RECT 210.6000 579.4500 211.8000 579.6000 ;
	    RECT 193.8000 578.5500 211.8000 579.4500 ;
	    RECT 193.8000 578.4000 195.0000 578.5500 ;
	    RECT 210.6000 578.4000 211.8000 578.5500 ;
	    RECT 193.8000 577.2000 195.0000 577.5000 ;
	    RECT 193.8000 573.3000 195.0000 576.3000 ;
	    RECT 213.0000 573.3000 214.2000 580.5000 ;
	    RECT 215.4000 578.4000 216.6000 579.6000 ;
	    RECT 246.9000 579.3000 252.3000 579.9000 ;
	    RECT 254.1000 579.3000 255.0000 581.4000 ;
	    RECT 275.4000 580.2000 276.6000 580.5000 ;
	    RECT 277.8000 579.3000 279.0000 583.5000 ;
	    RECT 297.0000 582.4500 298.2000 582.6000 ;
	    RECT 299.4000 582.4500 300.6000 582.6000 ;
	    RECT 297.0000 581.5500 300.6000 582.4500 ;
	    RECT 297.0000 581.4000 298.2000 581.5500 ;
	    RECT 299.4000 581.4000 300.6000 581.5500 ;
	    RECT 299.4000 580.2000 300.6000 580.5000 ;
	    RECT 301.8000 579.3000 303.0000 583.5000 ;
	    RECT 337.8000 583.2000 339.0000 583.5000 ;
	    RECT 342.6000 583.2000 343.8000 583.5000 ;
	    RECT 335.4000 581.4000 336.6000 582.6000 ;
	    RECT 337.8000 581.4000 339.3000 582.3000 ;
	    RECT 340.2000 581.4000 341.4000 582.6000 ;
	    RECT 337.8000 579.3000 338.7000 581.4000 ;
	    RECT 343.8000 580.8000 344.1000 582.3000 ;
	    RECT 345.0000 581.4000 346.2000 582.6000 ;
	    RECT 349.8000 582.4500 351.0000 582.6000 ;
	    RECT 359.4000 582.4500 360.6000 582.6000 ;
	    RECT 349.8000 581.5500 360.6000 582.4500 ;
	    RECT 349.8000 581.4000 351.0000 581.5500 ;
	    RECT 359.4000 581.4000 360.6000 581.5500 ;
	    RECT 381.0000 581.4000 382.2000 582.6000 ;
	    RECT 340.5000 579.3000 345.9000 579.9000 ;
	    RECT 246.6000 579.0000 252.6000 579.3000 ;
	    RECT 215.4000 577.2000 216.6000 577.5000 ;
	    RECT 215.4000 573.3000 216.6000 576.3000 ;
	    RECT 246.6000 573.3000 247.8000 579.0000 ;
	    RECT 249.0000 573.3000 250.2000 578.1000 ;
	    RECT 251.4000 574.2000 252.6000 579.0000 ;
	    RECT 253.8000 575.1000 255.0000 579.3000 ;
	    RECT 256.2000 574.2000 257.4000 579.3000 ;
	    RECT 251.4000 573.3000 257.4000 574.2000 ;
	    RECT 275.4000 573.3000 276.6000 579.3000 ;
	    RECT 277.8000 578.4000 280.5000 579.3000 ;
	    RECT 279.3000 573.3000 280.5000 578.4000 ;
	    RECT 299.4000 573.3000 300.6000 579.3000 ;
	    RECT 301.8000 578.4000 304.5000 579.3000 ;
	    RECT 303.3000 573.3000 304.5000 578.4000 ;
	    RECT 335.4000 574.2000 336.6000 579.3000 ;
	    RECT 337.8000 575.1000 339.0000 579.3000 ;
	    RECT 340.2000 579.0000 346.2000 579.3000 ;
	    RECT 340.2000 574.2000 341.4000 579.0000 ;
	    RECT 335.4000 573.3000 341.4000 574.2000 ;
	    RECT 342.6000 573.3000 343.8000 578.1000 ;
	    RECT 345.0000 573.3000 346.2000 579.0000 ;
	    RECT 359.4000 573.3000 360.6000 580.5000 ;
	    RECT 381.0000 580.2000 382.2000 580.5000 ;
	    RECT 361.8000 578.4000 363.0000 579.6000 ;
	    RECT 383.4000 579.3000 384.6000 583.5000 ;
	    RECT 385.8000 582.4500 387.0000 582.6000 ;
	    RECT 405.0000 582.4500 406.2000 582.6000 ;
	    RECT 385.8000 581.5500 406.2000 582.4500 ;
	    RECT 385.8000 581.4000 387.0000 581.5500 ;
	    RECT 405.0000 581.4000 406.2000 581.5500 ;
	    RECT 405.0000 580.2000 406.2000 580.5000 ;
	    RECT 407.4000 579.3000 408.6000 583.5000 ;
	    RECT 460.8000 582.6000 461.7000 587.7000 ;
	    RECT 489.0000 587.4000 490.2000 588.6000 ;
	    RECT 492.0000 587.7000 493.5000 588.6000 ;
	    RECT 496.2000 587.7000 497.4000 599.7000 ;
	    RECT 462.6000 584.4000 463.8000 585.6000 ;
	    RECT 462.6000 583.2000 463.8000 583.5000 ;
	    RECT 492.0000 582.6000 492.9000 587.7000 ;
	    RECT 493.8000 585.4500 495.0000 585.6000 ;
	    RECT 493.8000 584.5500 506.8500 585.4500 ;
	    RECT 493.8000 584.4000 495.0000 584.5500 ;
	    RECT 493.8000 583.2000 495.0000 583.5000 ;
	    RECT 409.8000 582.4500 411.0000 582.6000 ;
	    RECT 424.2000 582.4500 425.4000 582.6000 ;
	    RECT 409.8000 581.5500 425.4000 582.4500 ;
	    RECT 409.8000 581.4000 411.0000 581.5500 ;
	    RECT 424.2000 581.4000 425.4000 581.5500 ;
	    RECT 457.8000 581.4000 459.0000 582.6000 ;
	    RECT 459.9000 581.4000 461.7000 582.6000 ;
	    RECT 465.0000 582.4500 466.2000 582.6000 ;
	    RECT 486.6000 582.4500 487.8000 582.6000 ;
	    RECT 463.8000 580.8000 464.1000 582.3000 ;
	    RECT 465.0000 581.5500 487.8000 582.4500 ;
	    RECT 465.0000 581.4000 466.2000 581.5500 ;
	    RECT 486.6000 581.4000 487.8000 581.5500 ;
	    RECT 489.0000 581.4000 490.2000 582.6000 ;
	    RECT 491.1000 581.4000 492.9000 582.6000 ;
	    RECT 496.2000 582.4500 497.4000 582.6000 ;
	    RECT 503.4000 582.4500 504.6000 582.6000 ;
	    RECT 495.0000 580.8000 495.3000 582.3000 ;
	    RECT 496.2000 581.5500 504.6000 582.4500 ;
	    RECT 505.9500 582.4500 506.8500 584.5500 ;
	    RECT 510.6000 583.5000 511.8000 599.7000 ;
	    RECT 513.0000 593.7000 514.2000 599.7000 ;
	    RECT 532.2000 593.7000 533.4000 599.7000 ;
	    RECT 534.6000 586.5000 535.8000 599.7000 ;
	    RECT 537.0000 593.7000 538.2000 599.7000 ;
	    RECT 537.0000 589.5000 538.2000 589.8000 ;
	    RECT 577.8000 588.6000 579.0000 599.7000 ;
	    RECT 580.2000 589.8000 581.7000 599.7000 ;
	    RECT 580.2000 588.6000 581.4000 588.9000 ;
	    RECT 537.0000 588.4500 538.2000 588.6000 ;
	    RECT 563.4000 588.4500 564.6000 588.6000 ;
	    RECT 537.0000 587.5500 564.6000 588.4500 ;
	    RECT 577.8000 587.7000 581.4000 588.6000 ;
	    RECT 584.4000 587.7000 586.8000 599.7000 ;
	    RECT 589.5000 589.8000 591.0000 599.7000 ;
	    RECT 589.5000 588.6000 590.7000 588.9000 ;
	    RECT 592.2000 588.6000 593.4000 599.7000 ;
	    RECT 712.2000 599.4000 713.4000 600.6000 ;
	    RECT 609.0000 597.4500 610.2000 597.6000 ;
	    RECT 721.8000 597.4500 723.0000 597.6000 ;
	    RECT 609.0000 596.5500 723.0000 597.4500 ;
	    RECT 609.0000 596.4000 610.2000 596.5500 ;
	    RECT 721.8000 596.4000 723.0000 596.5500 ;
	    RECT 724.2000 593.7000 725.4000 599.7000 ;
	    RECT 726.6000 594.6000 727.8000 599.7000 ;
	    RECT 726.3000 593.7000 727.8000 594.6000 ;
	    RECT 729.0000 593.7000 730.2000 600.6000 ;
	    RECT 726.3000 592.8000 727.2000 593.7000 ;
	    RECT 731.4000 592.8000 732.6000 599.7000 ;
	    RECT 733.8000 593.7000 735.0000 599.7000 ;
	    RECT 736.2000 595.5000 737.4000 599.7000 ;
	    RECT 738.6000 595.5000 739.8000 599.7000 ;
	    RECT 589.5000 587.7000 593.4000 588.6000 ;
	    RECT 724.2000 591.9000 727.2000 592.8000 ;
	    RECT 537.0000 587.4000 538.2000 587.5500 ;
	    RECT 563.4000 587.4000 564.6000 587.5500 ;
	    RECT 585.0000 586.5000 585.9000 587.7000 ;
	    RECT 587.7000 585.6000 588.9000 585.9000 ;
	    RECT 534.6000 585.4500 535.8000 585.6000 ;
	    RECT 577.8000 585.4500 579.0000 585.6000 ;
	    RECT 534.6000 584.5500 579.0000 585.4500 ;
	    RECT 534.6000 584.4000 535.8000 584.5500 ;
	    RECT 577.8000 584.4000 579.0000 584.5500 ;
	    RECT 585.0000 584.4000 586.2000 585.6000 ;
	    RECT 587.7000 584.7000 590.1000 585.6000 ;
	    RECT 588.9000 584.4000 590.1000 584.7000 ;
	    RECT 724.2000 583.5000 725.4000 591.9000 ;
	    RECT 728.1000 591.6000 734.4000 592.8000 ;
	    RECT 741.0000 592.5000 742.2000 599.7000 ;
	    RECT 743.4000 593.7000 744.6000 599.7000 ;
	    RECT 745.8000 592.5000 747.0000 599.7000 ;
	    RECT 748.2000 593.7000 749.4000 599.7000 ;
	    RECT 728.1000 591.0000 729.0000 591.6000 ;
	    RECT 726.6000 589.8000 729.0000 591.0000 ;
	    RECT 733.5000 590.7000 742.2000 591.6000 ;
	    RECT 730.5000 589.8000 732.6000 590.7000 ;
	    RECT 730.5000 589.5000 739.8000 589.8000 ;
	    RECT 731.7000 588.9000 739.8000 589.5000 ;
	    RECT 738.6000 588.6000 739.8000 588.9000 ;
	    RECT 741.3000 589.5000 742.2000 590.7000 ;
	    RECT 743.1000 590.4000 747.0000 591.6000 ;
	    RECT 750.6000 590.4000 751.8000 599.7000 ;
	    RECT 753.0000 595.5000 754.2000 599.7000 ;
	    RECT 755.4000 595.5000 756.6000 599.7000 ;
	    RECT 757.8000 595.5000 759.0000 599.7000 ;
	    RECT 760.2000 593.7000 761.4000 599.7000 ;
	    RECT 755.4000 591.6000 761.7000 592.8000 ;
	    RECT 762.6000 591.6000 763.8000 599.7000 ;
	    RECT 765.0000 593.7000 766.2000 599.7000 ;
	    RECT 767.4000 592.8000 768.6000 599.7000 ;
	    RECT 769.8000 593.7000 771.0000 599.7000 ;
	    RECT 767.4000 591.9000 771.3000 592.8000 ;
	    RECT 772.2000 592.5000 773.4000 599.7000 ;
	    RECT 774.6000 593.7000 775.8000 599.7000 ;
	    RECT 762.6000 590.4000 766.5000 591.6000 ;
	    RECT 753.0000 589.5000 754.2000 589.8000 ;
	    RECT 741.3000 588.6000 754.2000 589.5000 ;
	    RECT 757.8000 589.5000 759.0000 589.8000 ;
	    RECT 770.4000 589.5000 771.3000 591.9000 ;
	    RECT 772.2000 590.4000 773.4000 591.6000 ;
	    RECT 757.8000 588.6000 771.3000 589.5000 ;
	    RECT 726.6000 588.4500 727.8000 588.6000 ;
	    RECT 729.0000 588.4500 730.2000 588.6000 ;
	    RECT 726.6000 587.5500 730.2000 588.4500 ;
	    RECT 734.1000 587.7000 735.3000 588.0000 ;
	    RECT 726.6000 587.4000 727.8000 587.5500 ;
	    RECT 729.0000 587.4000 730.2000 587.5500 ;
	    RECT 731.1000 586.8000 769.5000 587.7000 ;
	    RECT 768.3000 586.5000 769.5000 586.8000 ;
	    RECT 770.4000 585.9000 771.3000 588.6000 ;
	    RECT 772.2000 588.0000 773.4000 589.5000 ;
	    RECT 817.8000 588.6000 819.0000 599.7000 ;
	    RECT 820.2000 589.8000 821.7000 599.7000 ;
	    RECT 820.2000 588.6000 821.4000 588.9000 ;
	    RECT 772.2000 586.8000 773.7000 588.0000 ;
	    RECT 817.8000 587.7000 821.4000 588.6000 ;
	    RECT 824.4000 587.7000 826.8000 599.7000 ;
	    RECT 829.5000 589.8000 831.0000 599.7000 ;
	    RECT 829.5000 588.6000 830.7000 588.9000 ;
	    RECT 832.2000 588.6000 833.4000 599.7000 ;
	    RECT 846.6000 593.7000 847.8000 599.7000 ;
	    RECT 829.5000 587.7000 833.4000 588.6000 ;
	    RECT 726.3000 585.0000 732.9000 585.9000 ;
	    RECT 726.3000 584.7000 727.5000 585.0000 ;
	    RECT 733.8000 584.4000 735.0000 585.6000 ;
	    RECT 735.9000 585.0000 761.4000 585.9000 ;
	    RECT 770.4000 585.0000 771.6000 585.9000 ;
	    RECT 760.2000 584.1000 761.4000 585.0000 ;
	    RECT 510.6000 582.4500 511.8000 582.6000 ;
	    RECT 505.9500 581.5500 511.8000 582.4500 ;
	    RECT 496.2000 581.4000 497.4000 581.5500 ;
	    RECT 503.4000 581.4000 504.6000 581.5500 ;
	    RECT 510.6000 581.4000 511.8000 581.5500 ;
	    RECT 515.4000 582.4500 516.6000 582.6000 ;
	    RECT 532.2000 582.4500 533.4000 582.6000 ;
	    RECT 515.4000 581.5500 533.4000 582.4500 ;
	    RECT 515.4000 581.4000 516.6000 581.5500 ;
	    RECT 532.2000 581.4000 533.4000 581.5500 ;
	    RECT 361.8000 577.2000 363.0000 577.5000 ;
	    RECT 361.8000 573.3000 363.0000 576.3000 ;
	    RECT 381.0000 573.3000 382.2000 579.3000 ;
	    RECT 383.4000 578.4000 386.1000 579.3000 ;
	    RECT 384.9000 573.3000 386.1000 578.4000 ;
	    RECT 405.0000 573.3000 406.2000 579.3000 ;
	    RECT 407.4000 578.4000 410.1000 579.3000 ;
	    RECT 408.9000 573.3000 410.1000 578.4000 ;
	    RECT 424.2000 573.3000 425.4000 580.5000 ;
	    RECT 426.6000 579.4500 427.8000 579.6000 ;
	    RECT 453.0000 579.4500 454.2000 579.6000 ;
	    RECT 426.6000 578.5500 454.2000 579.4500 ;
	    RECT 458.1000 579.3000 459.0000 580.5000 ;
	    RECT 460.5000 579.3000 465.9000 579.9000 ;
	    RECT 489.3000 579.3000 490.2000 580.5000 ;
	    RECT 491.7000 579.3000 497.1000 579.9000 ;
	    RECT 426.6000 578.4000 427.8000 578.5500 ;
	    RECT 453.0000 578.4000 454.2000 578.5500 ;
	    RECT 426.6000 577.2000 427.8000 577.5000 ;
	    RECT 426.6000 573.3000 427.8000 576.3000 ;
	    RECT 457.8000 573.3000 459.0000 579.3000 ;
	    RECT 460.2000 579.0000 466.2000 579.3000 ;
	    RECT 460.2000 573.3000 461.4000 579.0000 ;
	    RECT 462.6000 573.3000 463.8000 578.1000 ;
	    RECT 465.0000 573.3000 466.2000 579.0000 ;
	    RECT 489.0000 573.3000 490.2000 579.3000 ;
	    RECT 491.4000 579.0000 497.4000 579.3000 ;
	    RECT 491.4000 573.3000 492.6000 579.0000 ;
	    RECT 493.8000 573.3000 495.0000 578.1000 ;
	    RECT 496.2000 573.3000 497.4000 579.0000 ;
	    RECT 510.6000 573.3000 511.8000 580.5000 ;
	    RECT 532.2000 580.2000 533.4000 580.5000 ;
	    RECT 513.0000 579.4500 514.2000 579.6000 ;
	    RECT 520.2000 579.4500 521.4000 579.6000 ;
	    RECT 513.0000 578.5500 521.4000 579.4500 ;
	    RECT 534.6000 579.3000 535.8000 583.5000 ;
	    RECT 585.0000 582.6000 585.9000 583.5000 ;
	    RECT 563.4000 582.4500 564.6000 582.6000 ;
	    RECT 575.4000 582.4500 576.6000 582.6000 ;
	    RECT 577.8000 582.4500 579.0000 582.6000 ;
	    RECT 563.4000 581.5500 579.0000 582.4500 ;
	    RECT 563.4000 581.4000 564.6000 581.5500 ;
	    RECT 575.4000 581.4000 576.6000 581.5500 ;
	    RECT 577.8000 581.4000 579.0000 581.5500 ;
	    RECT 579.9000 581.4000 580.2000 582.6000 ;
	    RECT 582.0000 581.4000 583.2000 582.6000 ;
	    RECT 582.3000 580.8000 583.2000 581.4000 ;
	    RECT 584.4000 581.7000 585.9000 582.6000 ;
	    RECT 586.8000 582.9000 588.0000 583.2000 ;
	    RECT 586.8000 582.6000 591.0000 582.9000 ;
	    RECT 586.8000 582.0000 591.3000 582.6000 ;
	    RECT 590.1000 581.7000 591.3000 582.0000 ;
	    RECT 580.2000 580.2000 581.4000 580.5000 ;
	    RECT 577.8000 579.3000 581.4000 580.2000 ;
	    RECT 582.3000 579.6000 583.5000 580.8000 ;
	    RECT 513.0000 578.4000 514.2000 578.5500 ;
	    RECT 520.2000 578.4000 521.4000 578.5500 ;
	    RECT 513.0000 577.2000 514.2000 577.5000 ;
	    RECT 513.0000 573.3000 514.2000 576.3000 ;
	    RECT 532.2000 573.3000 533.4000 579.3000 ;
	    RECT 534.6000 578.4000 537.3000 579.3000 ;
	    RECT 536.1000 573.3000 537.3000 578.4000 ;
	    RECT 577.8000 573.3000 579.0000 579.3000 ;
	    RECT 584.4000 578.7000 585.3000 581.7000 ;
	    RECT 591.0000 581.4000 591.3000 581.7000 ;
	    RECT 592.2000 582.4500 593.4000 582.6000 ;
	    RECT 630.6000 582.4500 631.8000 582.6000 ;
	    RECT 592.2000 581.5500 631.8000 582.4500 ;
	    RECT 592.2000 581.4000 593.4000 581.5500 ;
	    RECT 630.6000 581.4000 631.8000 581.5500 ;
	    RECT 724.2000 582.3000 737.4000 583.5000 ;
	    RECT 738.3000 582.9000 741.3000 584.1000 ;
	    RECT 747.0000 582.9000 751.8000 584.1000 ;
	    RECT 586.2000 579.6000 588.6000 580.8000 ;
	    RECT 589.5000 580.2000 590.7000 580.5000 ;
	    RECT 589.5000 579.3000 593.4000 580.2000 ;
	    RECT 580.2000 573.3000 581.7000 578.4000 ;
	    RECT 584.4000 573.3000 586.8000 578.7000 ;
	    RECT 589.5000 573.3000 591.0000 578.4000 ;
	    RECT 592.2000 573.3000 593.4000 579.3000 ;
	    RECT 724.2000 573.3000 725.4000 582.3000 ;
	    RECT 727.8000 580.2000 732.3000 581.4000 ;
	    RECT 731.1000 579.3000 732.3000 580.2000 ;
	    RECT 740.1000 579.3000 741.3000 582.9000 ;
	    RECT 743.4000 581.4000 744.6000 582.6000 ;
	    RECT 751.2000 581.7000 752.4000 582.0000 ;
	    RECT 745.8000 580.8000 752.4000 581.7000 ;
	    RECT 745.8000 580.5000 747.0000 580.8000 ;
	    RECT 743.4000 580.2000 744.6000 580.5000 ;
	    RECT 755.4000 579.6000 756.6000 583.8000 ;
	    RECT 764.1000 582.9000 769.8000 584.1000 ;
	    RECT 764.1000 581.1000 765.3000 582.9000 ;
	    RECT 770.7000 582.0000 771.6000 585.0000 ;
	    RECT 745.8000 579.3000 747.0000 579.6000 ;
	    RECT 729.0000 573.3000 730.2000 579.3000 ;
	    RECT 731.1000 578.1000 735.0000 579.3000 ;
	    RECT 740.1000 578.4000 747.0000 579.3000 ;
	    RECT 748.2000 578.4000 749.4000 579.6000 ;
	    RECT 750.3000 578.4000 750.6000 579.6000 ;
	    RECT 755.1000 578.4000 756.6000 579.6000 ;
	    RECT 762.6000 580.2000 765.3000 581.1000 ;
	    RECT 769.8000 581.1000 771.6000 582.0000 ;
	    RECT 762.6000 579.3000 763.8000 580.2000 ;
	    RECT 733.8000 573.3000 735.0000 578.1000 ;
	    RECT 760.2000 578.1000 763.8000 579.3000 ;
	    RECT 736.2000 573.3000 737.4000 577.5000 ;
	    RECT 738.6000 573.3000 739.8000 577.5000 ;
	    RECT 741.0000 573.3000 742.2000 577.5000 ;
	    RECT 743.4000 573.3000 744.6000 576.3000 ;
	    RECT 745.8000 573.3000 747.0000 577.5000 ;
	    RECT 748.2000 573.3000 749.4000 576.3000 ;
	    RECT 750.6000 573.3000 751.8000 577.5000 ;
	    RECT 753.0000 573.3000 754.2000 577.5000 ;
	    RECT 755.4000 573.3000 756.6000 577.5000 ;
	    RECT 757.8000 573.3000 759.0000 577.5000 ;
	    RECT 760.2000 573.3000 761.4000 578.1000 ;
	    RECT 765.0000 573.3000 766.2000 579.3000 ;
	    RECT 769.8000 573.3000 771.0000 581.1000 ;
	    RECT 772.5000 580.2000 773.7000 586.8000 ;
	    RECT 825.0000 586.5000 825.9000 587.7000 ;
	    RECT 827.7000 585.6000 828.9000 585.9000 ;
	    RECT 774.6000 585.4500 775.8000 585.6000 ;
	    RECT 825.0000 585.4500 826.2000 585.6000 ;
	    RECT 774.6000 584.5500 826.2000 585.4500 ;
	    RECT 827.7000 584.7000 830.1000 585.6000 ;
	    RECT 774.6000 584.4000 775.8000 584.5500 ;
	    RECT 825.0000 584.4000 826.2000 584.5500 ;
	    RECT 828.9000 584.4000 830.1000 584.7000 ;
	    RECT 849.0000 583.5000 850.2000 599.7000 ;
	    RECT 873.0000 593.7000 874.2000 599.7000 ;
	    RECT 875.4000 593.7000 876.6000 599.7000 ;
	    RECT 877.8000 594.3000 879.0000 599.7000 ;
	    RECT 875.7000 593.4000 876.6000 593.7000 ;
	    RECT 880.2000 593.7000 881.4000 599.7000 ;
	    RECT 906.6000 593.7000 907.8000 599.7000 ;
	    RECT 880.2000 593.4000 881.1000 593.7000 ;
	    RECT 875.7000 592.5000 881.1000 593.4000 ;
	    RECT 870.6000 591.4500 871.8000 591.6000 ;
	    RECT 877.8000 591.4500 879.0000 591.6000 ;
	    RECT 870.6000 590.5500 879.0000 591.4500 ;
	    RECT 870.6000 590.4000 871.8000 590.5500 ;
	    RECT 877.8000 590.4000 879.0000 590.5500 ;
	    RECT 880.2000 589.5000 881.1000 592.5000 ;
	    RECT 906.6000 589.5000 907.8000 589.8000 ;
	    RECT 877.8000 589.2000 879.0000 589.5000 ;
	    RECT 861.0000 588.4500 862.2000 588.6000 ;
	    RECT 873.0000 588.4500 874.2000 588.6000 ;
	    RECT 861.0000 587.5500 874.2000 588.4500 ;
	    RECT 861.0000 587.4000 862.2000 587.5500 ;
	    RECT 873.0000 587.4000 874.2000 587.5500 ;
	    RECT 880.2000 588.4500 881.4000 588.6000 ;
	    RECT 906.6000 588.4500 907.8000 588.6000 ;
	    RECT 880.2000 587.5500 907.8000 588.4500 ;
	    RECT 880.2000 587.4000 881.4000 587.5500 ;
	    RECT 906.6000 587.4000 907.8000 587.5500 ;
	    RECT 909.0000 586.5000 910.2000 599.7000 ;
	    RECT 911.4000 593.7000 912.6000 599.7000 ;
	    RECT 873.0000 586.2000 874.2000 586.5000 ;
	    RECT 875.4000 584.4000 876.6000 585.6000 ;
	    RECT 877.5000 584.4000 877.8000 585.6000 ;
	    RECT 825.0000 582.6000 825.9000 583.5000 ;
	    RECT 786.6000 582.4500 787.8000 582.6000 ;
	    RECT 805.8000 582.4500 807.0000 582.6000 ;
	    RECT 817.8000 582.4500 819.0000 582.6000 ;
	    RECT 786.6000 581.5500 819.0000 582.4500 ;
	    RECT 786.6000 581.4000 787.8000 581.5500 ;
	    RECT 805.8000 581.4000 807.0000 581.5500 ;
	    RECT 817.8000 581.4000 819.0000 581.5500 ;
	    RECT 819.9000 581.4000 820.2000 582.6000 ;
	    RECT 822.0000 581.4000 823.2000 582.6000 ;
	    RECT 822.3000 580.8000 823.2000 581.4000 ;
	    RECT 824.4000 581.7000 825.9000 582.6000 ;
	    RECT 826.8000 582.9000 828.0000 583.2000 ;
	    RECT 826.8000 582.6000 831.0000 582.9000 ;
	    RECT 880.2000 582.6000 881.1000 586.5000 ;
	    RECT 909.0000 585.4500 910.2000 585.6000 ;
	    RECT 913.8000 585.4500 915.0000 585.6000 ;
	    RECT 909.0000 584.5500 915.0000 585.4500 ;
	    RECT 909.0000 584.4000 910.2000 584.5500 ;
	    RECT 913.8000 584.4000 915.0000 584.5500 ;
	    RECT 925.8000 583.5000 927.0000 599.7000 ;
	    RECT 928.2000 593.7000 929.4000 599.7000 ;
	    RECT 949.8000 599.4000 951.0000 600.6000 ;
	    RECT 955.5000 593.7000 956.7000 599.7000 ;
	    RECT 955.8000 590.4000 957.0000 591.6000 ;
	    RECT 955.8000 589.5000 956.7000 590.4000 ;
	    RECT 957.9000 588.6000 959.1000 599.7000 ;
	    RECT 954.6000 587.4000 955.8000 588.6000 ;
	    RECT 957.6000 587.7000 959.1000 588.6000 ;
	    RECT 961.8000 587.7000 963.0000 599.7000 ;
	    RECT 981.0000 593.7000 982.2000 599.7000 ;
	    RECT 981.0000 589.5000 982.2000 589.8000 ;
	    RECT 978.6000 588.4500 979.8000 588.6000 ;
	    RECT 981.0000 588.4500 982.2000 588.6000 ;
	    RECT 826.8000 582.0000 831.3000 582.6000 ;
	    RECT 830.1000 581.7000 831.3000 582.0000 ;
	    RECT 820.2000 580.2000 821.4000 580.5000 ;
	    RECT 772.2000 579.0000 773.7000 580.2000 ;
	    RECT 817.8000 579.3000 821.4000 580.2000 ;
	    RECT 822.3000 579.6000 823.5000 580.8000 ;
	    RECT 772.2000 573.3000 773.4000 579.0000 ;
	    RECT 774.6000 573.3000 775.8000 576.3000 ;
	    RECT 817.8000 573.3000 819.0000 579.3000 ;
	    RECT 824.4000 578.7000 825.3000 581.7000 ;
	    RECT 831.0000 581.4000 831.3000 581.7000 ;
	    RECT 832.2000 582.4500 833.4000 582.6000 ;
	    RECT 837.0000 582.4500 838.2000 582.6000 ;
	    RECT 832.2000 581.5500 838.2000 582.4500 ;
	    RECT 832.2000 581.4000 833.4000 581.5500 ;
	    RECT 837.0000 581.4000 838.2000 581.5500 ;
	    RECT 849.0000 582.4500 850.2000 582.6000 ;
	    RECT 870.6000 582.4500 871.8000 582.6000 ;
	    RECT 849.0000 581.5500 871.8000 582.4500 ;
	    RECT 878.7000 582.3000 881.1000 582.6000 ;
	    RECT 849.0000 581.4000 850.2000 581.5500 ;
	    RECT 870.6000 581.4000 871.8000 581.5500 ;
	    RECT 826.2000 579.6000 828.6000 580.8000 ;
	    RECT 829.5000 580.2000 830.7000 580.5000 ;
	    RECT 829.5000 579.3000 833.4000 580.2000 ;
	    RECT 820.2000 573.3000 821.7000 578.4000 ;
	    RECT 824.4000 573.3000 826.8000 578.7000 ;
	    RECT 829.5000 573.3000 831.0000 578.4000 ;
	    RECT 832.2000 573.3000 833.4000 579.3000 ;
	    RECT 841.8000 579.4500 843.0000 579.6000 ;
	    RECT 846.6000 579.4500 847.8000 579.6000 ;
	    RECT 841.8000 578.5500 847.8000 579.4500 ;
	    RECT 841.8000 578.4000 843.0000 578.5500 ;
	    RECT 846.6000 578.4000 847.8000 578.5500 ;
	    RECT 846.6000 577.2000 847.8000 577.5000 ;
	    RECT 846.6000 573.3000 847.8000 576.3000 ;
	    RECT 849.0000 573.3000 850.2000 580.5000 ;
	    RECT 873.0000 573.3000 874.2000 582.3000 ;
	    RECT 878.4000 581.7000 881.1000 582.3000 ;
	    RECT 878.4000 573.3000 879.6000 581.7000 ;
	    RECT 909.0000 579.3000 910.2000 583.5000 ;
	    RECT 957.6000 582.6000 958.5000 587.7000 ;
	    RECT 978.6000 587.5500 982.2000 588.4500 ;
	    RECT 978.6000 587.4000 979.8000 587.5500 ;
	    RECT 981.0000 587.4000 982.2000 587.5500 ;
	    RECT 983.4000 586.5000 984.6000 599.7000 ;
	    RECT 985.8000 593.7000 987.0000 599.7000 ;
	    RECT 1120.2001 593.7000 1121.4000 599.7000 ;
	    RECT 1122.6000 594.6000 1123.8000 599.7000 ;
	    RECT 1122.3000 593.7000 1123.8000 594.6000 ;
	    RECT 1125.0000 593.7000 1126.2001 600.6000 ;
	    RECT 1122.3000 592.8000 1123.2001 593.7000 ;
	    RECT 1127.4000 592.8000 1128.6000 599.7000 ;
	    RECT 1129.8000 593.7000 1131.0000 599.7000 ;
	    RECT 1132.2001 595.5000 1133.4000 599.7000 ;
	    RECT 1134.6000 595.5000 1135.8000 599.7000 ;
	    RECT 1120.2001 591.9000 1123.2001 592.8000 ;
	    RECT 959.4000 584.4000 960.6000 585.6000 ;
	    RECT 964.2000 585.4500 965.4000 585.6000 ;
	    RECT 983.4000 585.4500 984.6000 585.6000 ;
	    RECT 964.2000 584.5500 984.6000 585.4500 ;
	    RECT 964.2000 584.4000 965.4000 584.5500 ;
	    RECT 983.4000 584.4000 984.6000 584.5500 ;
	    RECT 1120.2001 583.5000 1121.4000 591.9000 ;
	    RECT 1124.1000 591.6000 1130.4000 592.8000 ;
	    RECT 1137.0000 592.5000 1138.2001 599.7000 ;
	    RECT 1139.4000 593.7000 1140.6000 599.7000 ;
	    RECT 1141.8000 592.5000 1143.0000 599.7000 ;
	    RECT 1144.2001 593.7000 1145.4000 599.7000 ;
	    RECT 1124.1000 591.0000 1125.0000 591.6000 ;
	    RECT 1122.6000 589.8000 1125.0000 591.0000 ;
	    RECT 1129.5000 590.7000 1138.2001 591.6000 ;
	    RECT 1126.5000 589.8000 1128.6000 590.7000 ;
	    RECT 1126.5000 589.5000 1135.8000 589.8000 ;
	    RECT 1127.7001 588.9000 1135.8000 589.5000 ;
	    RECT 1134.6000 588.6000 1135.8000 588.9000 ;
	    RECT 1137.3000 589.5000 1138.2001 590.7000 ;
	    RECT 1139.1000 590.4000 1143.0000 591.6000 ;
	    RECT 1146.6000 590.4000 1147.8000 599.7000 ;
	    RECT 1149.0000 595.5000 1150.2001 599.7000 ;
	    RECT 1151.4000 595.5000 1152.6000 599.7000 ;
	    RECT 1153.8000 595.5000 1155.0000 599.7000 ;
	    RECT 1156.2001 593.7000 1157.4000 599.7000 ;
	    RECT 1151.4000 591.6000 1157.7001 592.8000 ;
	    RECT 1158.6000 591.6000 1159.8000 599.7000 ;
	    RECT 1161.0000 593.7000 1162.2001 599.7000 ;
	    RECT 1163.4000 592.8000 1164.6000 599.7000 ;
	    RECT 1165.8000 593.7000 1167.0000 599.7000 ;
	    RECT 1163.4000 591.9000 1167.3000 592.8000 ;
	    RECT 1168.2001 592.5000 1169.4000 599.7000 ;
	    RECT 1170.6000 593.7000 1171.8000 599.7000 ;
	    RECT 1189.8000 593.7000 1191.0000 599.7000 ;
	    RECT 1158.6000 590.4000 1162.5000 591.6000 ;
	    RECT 1149.0000 589.5000 1150.2001 589.8000 ;
	    RECT 1137.3000 588.6000 1150.2001 589.5000 ;
	    RECT 1153.8000 589.5000 1155.0000 589.8000 ;
	    RECT 1166.4000 589.5000 1167.3000 591.9000 ;
	    RECT 1168.2001 590.4000 1169.4000 591.6000 ;
	    RECT 1153.8000 588.6000 1167.3000 589.5000 ;
	    RECT 1125.0000 587.4000 1126.2001 588.6000 ;
	    RECT 1130.1000 587.7000 1131.3000 588.0000 ;
	    RECT 1127.1000 586.8000 1165.5000 587.7000 ;
	    RECT 1164.3000 586.5000 1165.5000 586.8000 ;
	    RECT 1166.4000 585.9000 1167.3000 588.6000 ;
	    RECT 1168.2001 588.0000 1169.4000 589.5000 ;
	    RECT 1168.2001 586.8000 1169.7001 588.0000 ;
	    RECT 1122.3000 585.0000 1128.9000 585.9000 ;
	    RECT 1122.3000 584.7000 1123.5000 585.0000 ;
	    RECT 1129.8000 584.4000 1131.0000 585.6000 ;
	    RECT 1131.9000 585.0000 1157.4000 585.9000 ;
	    RECT 1166.4000 585.0000 1167.6000 585.9000 ;
	    RECT 1156.2001 584.1000 1157.4000 585.0000 ;
	    RECT 959.4000 583.2000 960.6000 583.5000 ;
	    RECT 911.4000 581.4000 912.6000 582.6000 ;
	    RECT 925.8000 582.4500 927.0000 582.6000 ;
	    RECT 933.0000 582.4500 934.2000 582.6000 ;
	    RECT 925.8000 581.5500 934.2000 582.4500 ;
	    RECT 925.8000 581.4000 927.0000 581.5500 ;
	    RECT 933.0000 581.4000 934.2000 581.5500 ;
	    RECT 935.4000 582.4500 936.6000 582.6000 ;
	    RECT 954.6000 582.4500 955.8000 582.6000 ;
	    RECT 935.4000 581.5500 955.8000 582.4500 ;
	    RECT 935.4000 581.4000 936.6000 581.5500 ;
	    RECT 954.6000 581.4000 955.8000 581.5500 ;
	    RECT 956.7000 581.4000 958.5000 582.6000 ;
	    RECT 960.6000 580.8000 960.9000 582.3000 ;
	    RECT 961.8000 581.4000 963.0000 582.6000 ;
	    RECT 911.4000 580.2000 912.6000 580.5000 ;
	    RECT 907.5000 578.4000 910.2000 579.3000 ;
	    RECT 907.5000 573.3000 908.7000 578.4000 ;
	    RECT 911.4000 573.3000 912.6000 579.3000 ;
	    RECT 925.8000 573.3000 927.0000 580.5000 ;
	    RECT 928.2000 578.4000 929.4000 579.6000 ;
	    RECT 954.9000 579.3000 955.8000 580.5000 ;
	    RECT 957.3000 579.3000 962.7000 579.9000 ;
	    RECT 983.4000 579.3000 984.6000 583.5000 ;
	    RECT 985.8000 582.4500 987.0000 582.6000 ;
	    RECT 1007.4000 582.4500 1008.6000 582.6000 ;
	    RECT 985.8000 581.5500 1008.6000 582.4500 ;
	    RECT 985.8000 581.4000 987.0000 581.5500 ;
	    RECT 1007.4000 581.4000 1008.6000 581.5500 ;
	    RECT 1120.2001 582.3000 1133.4000 583.5000 ;
	    RECT 1134.3000 582.9000 1137.3000 584.1000 ;
	    RECT 1143.0000 582.9000 1147.8000 584.1000 ;
	    RECT 985.8000 580.2000 987.0000 580.5000 ;
	    RECT 928.2000 577.2000 929.4000 577.5000 ;
	    RECT 928.2000 573.3000 929.4000 576.3000 ;
	    RECT 954.6000 573.3000 955.8000 579.3000 ;
	    RECT 957.0000 579.0000 963.0000 579.3000 ;
	    RECT 957.0000 573.3000 958.2000 579.0000 ;
	    RECT 959.4000 573.3000 960.6000 578.1000 ;
	    RECT 961.8000 573.3000 963.0000 579.0000 ;
	    RECT 981.9000 578.4000 984.6000 579.3000 ;
	    RECT 981.9000 573.3000 983.1000 578.4000 ;
	    RECT 985.8000 573.3000 987.0000 579.3000 ;
	    RECT 1120.2001 573.3000 1121.4000 582.3000 ;
	    RECT 1123.8000 580.2000 1128.3000 581.4000 ;
	    RECT 1127.1000 579.3000 1128.3000 580.2000 ;
	    RECT 1136.1000 579.3000 1137.3000 582.9000 ;
	    RECT 1139.4000 581.4000 1140.6000 582.6000 ;
	    RECT 1147.2001 581.7000 1148.4000 582.0000 ;
	    RECT 1141.8000 580.8000 1148.4000 581.7000 ;
	    RECT 1141.8000 580.5000 1143.0000 580.8000 ;
	    RECT 1139.4000 580.2000 1140.6000 580.5000 ;
	    RECT 1151.4000 579.6000 1152.6000 583.8000 ;
	    RECT 1160.1000 582.9000 1165.8000 584.1000 ;
	    RECT 1160.1000 581.1000 1161.3000 582.9000 ;
	    RECT 1166.7001 582.0000 1167.6000 585.0000 ;
	    RECT 1141.8000 579.3000 1143.0000 579.6000 ;
	    RECT 1125.0000 573.3000 1126.2001 579.3000 ;
	    RECT 1127.1000 578.1000 1131.0000 579.3000 ;
	    RECT 1136.1000 578.4000 1143.0000 579.3000 ;
	    RECT 1144.2001 578.4000 1145.4000 579.6000 ;
	    RECT 1146.3000 578.4000 1146.6000 579.6000 ;
	    RECT 1151.1000 578.4000 1152.6000 579.6000 ;
	    RECT 1158.6000 580.2000 1161.3000 581.1000 ;
	    RECT 1165.8000 581.1000 1167.6000 582.0000 ;
	    RECT 1158.6000 579.3000 1159.8000 580.2000 ;
	    RECT 1129.8000 573.3000 1131.0000 578.1000 ;
	    RECT 1156.2001 578.1000 1159.8000 579.3000 ;
	    RECT 1132.2001 573.3000 1133.4000 577.5000 ;
	    RECT 1134.6000 573.3000 1135.8000 577.5000 ;
	    RECT 1137.0000 573.3000 1138.2001 577.5000 ;
	    RECT 1139.4000 573.3000 1140.6000 576.3000 ;
	    RECT 1141.8000 573.3000 1143.0000 577.5000 ;
	    RECT 1144.2001 573.3000 1145.4000 576.3000 ;
	    RECT 1146.6000 573.3000 1147.8000 577.5000 ;
	    RECT 1149.0000 573.3000 1150.2001 577.5000 ;
	    RECT 1151.4000 573.3000 1152.6000 577.5000 ;
	    RECT 1153.8000 573.3000 1155.0000 577.5000 ;
	    RECT 1156.2001 573.3000 1157.4000 578.1000 ;
	    RECT 1161.0000 573.3000 1162.2001 579.3000 ;
	    RECT 1165.8000 573.3000 1167.0000 581.1000 ;
	    RECT 1168.5000 580.2000 1169.7001 586.8000 ;
	    RECT 1192.2001 586.5000 1193.4000 599.7000 ;
	    RECT 1194.6000 593.7000 1195.8000 599.7000 ;
	    RECT 1213.8000 593.7000 1215.0000 599.7000 ;
	    RECT 1194.6000 589.5000 1195.8000 589.8000 ;
	    RECT 1213.8000 589.5000 1215.0000 589.8000 ;
	    RECT 1194.6000 588.4500 1195.8000 588.6000 ;
	    RECT 1199.4000 588.4500 1200.6000 588.6000 ;
	    RECT 1194.6000 587.5500 1200.6000 588.4500 ;
	    RECT 1194.6000 587.4000 1195.8000 587.5500 ;
	    RECT 1199.4000 587.4000 1200.6000 587.5500 ;
	    RECT 1204.2001 588.4500 1205.4000 588.6000 ;
	    RECT 1213.8000 588.4500 1215.0000 588.6000 ;
	    RECT 1204.2001 587.5500 1215.0000 588.4500 ;
	    RECT 1204.2001 587.4000 1205.4000 587.5500 ;
	    RECT 1213.8000 587.4000 1215.0000 587.5500 ;
	    RECT 1216.2001 586.5000 1217.4000 599.7000 ;
	    RECT 1218.6000 593.7000 1219.8000 599.7000 ;
	    RECT 1242.6000 587.7000 1243.8000 599.7000 ;
	    RECT 1246.5000 588.6000 1247.7001 599.7000 ;
	    RECT 1248.9000 593.7000 1250.1000 599.7000 ;
	    RECT 1269.0000 593.7000 1270.2001 599.7000 ;
	    RECT 1248.6000 590.4000 1249.8000 591.6000 ;
	    RECT 1248.9000 589.5000 1249.8000 590.4000 ;
	    RECT 1246.5000 587.7000 1248.0000 588.6000 ;
	    RECT 1182.6000 585.4500 1183.8000 585.6000 ;
	    RECT 1192.2001 585.4500 1193.4000 585.6000 ;
	    RECT 1182.6000 584.5500 1193.4000 585.4500 ;
	    RECT 1182.6000 584.4000 1183.8000 584.5500 ;
	    RECT 1192.2001 584.4000 1193.4000 584.5500 ;
	    RECT 1216.2001 584.4000 1217.4000 585.6000 ;
	    RECT 1245.0000 584.4000 1246.2001 585.6000 ;
	    RECT 1170.6000 582.4500 1171.8000 582.6000 ;
	    RECT 1189.8000 582.4500 1191.0000 582.6000 ;
	    RECT 1170.6000 581.5500 1191.0000 582.4500 ;
	    RECT 1170.6000 581.4000 1171.8000 581.5500 ;
	    RECT 1189.8000 581.4000 1191.0000 581.5500 ;
	    RECT 1189.8000 580.2000 1191.0000 580.5000 ;
	    RECT 1168.2001 579.0000 1169.7001 580.2000 ;
	    RECT 1192.2001 579.3000 1193.4000 583.5000 ;
	    RECT 1216.2001 579.3000 1217.4000 583.5000 ;
	    RECT 1245.0000 583.2000 1246.2001 583.5000 ;
	    RECT 1247.1000 582.6000 1248.0000 587.7000 ;
	    RECT 1249.8000 587.4000 1251.0000 588.6000 ;
	    RECT 1271.4000 586.5000 1272.6000 599.7000 ;
	    RECT 1273.8000 593.7000 1275.0000 599.7000 ;
	    RECT 1297.8000 593.7000 1299.0000 599.7000 ;
	    RECT 1300.2001 593.7000 1301.4000 599.7000 ;
	    RECT 1302.6000 594.3000 1303.8000 599.7000 ;
	    RECT 1300.5000 593.4000 1301.4000 593.7000 ;
	    RECT 1305.0000 593.7000 1306.2001 599.7000 ;
	    RECT 1331.4000 593.7000 1332.6000 599.7000 ;
	    RECT 1333.8000 593.7000 1335.0000 599.7000 ;
	    RECT 1336.2001 594.3000 1337.4000 599.7000 ;
	    RECT 1305.0000 593.4000 1305.9000 593.7000 ;
	    RECT 1300.5000 592.5000 1305.9000 593.4000 ;
	    RECT 1334.1000 593.4000 1335.0000 593.7000 ;
	    RECT 1338.6000 593.7000 1339.8000 599.7000 ;
	    RECT 1372.2001 593.7000 1373.4000 599.7000 ;
	    RECT 1374.6000 593.7000 1375.8000 599.7000 ;
	    RECT 1377.0000 594.3000 1378.2001 599.7000 ;
	    RECT 1338.6000 593.4000 1339.5000 593.7000 ;
	    RECT 1334.1000 592.5000 1339.5000 593.4000 ;
	    RECT 1374.9000 593.4000 1375.8000 593.7000 ;
	    RECT 1379.4000 593.7000 1380.6000 599.7000 ;
	    RECT 1403.4000 593.7000 1404.6000 599.7000 ;
	    RECT 1405.8000 593.7000 1407.0000 599.7000 ;
	    RECT 1408.2001 594.3000 1409.4000 599.7000 ;
	    RECT 1379.4000 593.4000 1380.3000 593.7000 ;
	    RECT 1374.9000 592.5000 1380.3000 593.4000 ;
	    RECT 1406.1000 593.4000 1407.0000 593.7000 ;
	    RECT 1410.6000 593.7000 1411.8000 599.7000 ;
	    RECT 1417.8000 599.4000 1419.0000 600.6000 ;
	    RECT 1429.8000 593.7000 1431.0000 599.7000 ;
	    RECT 1410.6000 593.4000 1411.5000 593.7000 ;
	    RECT 1406.1000 592.5000 1411.5000 593.4000 ;
	    RECT 1281.0000 591.4500 1282.2001 591.6000 ;
	    RECT 1302.6000 591.4500 1303.8000 591.6000 ;
	    RECT 1281.0000 590.5500 1303.8000 591.4500 ;
	    RECT 1281.0000 590.4000 1282.2001 590.5500 ;
	    RECT 1302.6000 590.4000 1303.8000 590.5500 ;
	    RECT 1273.8000 589.5000 1275.0000 589.8000 ;
	    RECT 1305.0000 589.5000 1305.9000 592.5000 ;
	    RECT 1312.2001 591.4500 1313.4000 591.6000 ;
	    RECT 1336.2001 591.4500 1337.4000 591.6000 ;
	    RECT 1312.2001 590.5500 1337.4000 591.4500 ;
	    RECT 1312.2001 590.4000 1313.4000 590.5500 ;
	    RECT 1336.2001 590.4000 1337.4000 590.5500 ;
	    RECT 1338.6000 589.5000 1339.5000 592.5000 ;
	    RECT 1377.0000 590.4000 1378.2001 591.6000 ;
	    RECT 1379.4000 589.5000 1380.3000 592.5000 ;
	    RECT 1408.2001 591.4500 1409.4000 591.6000 ;
	    RECT 1401.1500 590.5500 1409.4000 591.4500 ;
	    RECT 1302.6000 589.2000 1303.8000 589.5000 ;
	    RECT 1336.2001 589.2000 1337.4000 589.5000 ;
	    RECT 1377.0000 589.2000 1378.2001 589.5000 ;
	    RECT 1273.8000 588.4500 1275.0000 588.6000 ;
	    RECT 1276.2001 588.4500 1277.4000 588.6000 ;
	    RECT 1273.8000 587.5500 1277.4000 588.4500 ;
	    RECT 1273.8000 587.4000 1275.0000 587.5500 ;
	    RECT 1276.2001 587.4000 1277.4000 587.5500 ;
	    RECT 1278.6000 588.4500 1279.8000 588.6000 ;
	    RECT 1285.8000 588.4500 1287.0000 588.6000 ;
	    RECT 1297.8000 588.4500 1299.0000 588.6000 ;
	    RECT 1300.2001 588.4500 1301.4000 588.6000 ;
	    RECT 1278.6000 587.5500 1301.4000 588.4500 ;
	    RECT 1278.6000 587.4000 1279.8000 587.5500 ;
	    RECT 1285.8000 587.4000 1287.0000 587.5500 ;
	    RECT 1297.8000 587.4000 1299.0000 587.5500 ;
	    RECT 1300.2001 587.4000 1301.4000 587.5500 ;
	    RECT 1305.0000 588.4500 1306.2001 588.6000 ;
	    RECT 1329.0000 588.4500 1330.2001 588.6000 ;
	    RECT 1305.0000 587.5500 1330.2001 588.4500 ;
	    RECT 1305.0000 587.4000 1306.2001 587.5500 ;
	    RECT 1329.0000 587.4000 1330.2001 587.5500 ;
	    RECT 1331.4000 587.4000 1332.6000 588.6000 ;
	    RECT 1338.6000 588.4500 1339.8000 588.6000 ;
	    RECT 1343.4000 588.4500 1344.6000 588.6000 ;
	    RECT 1338.6000 587.5500 1344.6000 588.4500 ;
	    RECT 1338.6000 587.4000 1339.8000 587.5500 ;
	    RECT 1343.4000 587.4000 1344.6000 587.5500 ;
	    RECT 1348.2001 588.4500 1349.4000 588.6000 ;
	    RECT 1372.2001 588.4500 1373.4000 588.6000 ;
	    RECT 1348.2001 587.5500 1373.4000 588.4500 ;
	    RECT 1348.2001 587.4000 1349.4000 587.5500 ;
	    RECT 1372.2001 587.4000 1373.4000 587.5500 ;
	    RECT 1379.4000 588.4500 1380.6000 588.6000 ;
	    RECT 1401.1500 588.4500 1402.0500 590.5500 ;
	    RECT 1408.2001 590.4000 1409.4000 590.5500 ;
	    RECT 1410.6000 589.5000 1411.5000 592.5000 ;
	    RECT 1408.2001 589.2000 1409.4000 589.5000 ;
	    RECT 1379.4000 587.5500 1402.0500 588.4500 ;
	    RECT 1379.4000 587.4000 1380.6000 587.5500 ;
	    RECT 1403.4000 587.4000 1404.6000 588.6000 ;
	    RECT 1410.6000 587.4000 1411.8000 588.6000 ;
	    RECT 1432.2001 586.5000 1433.4000 599.7000 ;
	    RECT 1434.6000 593.7000 1435.8000 599.7000 ;
	    RECT 1458.6000 593.7000 1459.8000 599.7000 ;
	    RECT 1461.0000 593.7000 1462.2001 599.7000 ;
	    RECT 1463.4000 594.3000 1464.6000 599.7000 ;
	    RECT 1461.3000 593.4000 1462.2001 593.7000 ;
	    RECT 1465.8000 593.7000 1467.0000 599.7000 ;
	    RECT 1489.8000 593.7000 1491.0000 599.7000 ;
	    RECT 1492.2001 594.3000 1493.4000 599.7000 ;
	    RECT 1465.8000 593.4000 1466.7001 593.7000 ;
	    RECT 1461.3000 592.5000 1466.7001 593.4000 ;
	    RECT 1463.4000 590.4000 1464.6000 591.6000 ;
	    RECT 1434.6000 589.5000 1435.8000 589.8000 ;
	    RECT 1465.8000 589.5000 1466.7001 592.5000 ;
	    RECT 1490.1000 593.4000 1491.0000 593.7000 ;
	    RECT 1494.6000 593.7000 1495.8000 599.7000 ;
	    RECT 1497.0000 593.7000 1498.2001 599.7000 ;
	    RECT 1494.6000 593.4000 1495.5000 593.7000 ;
	    RECT 1490.1000 592.5000 1495.5000 593.4000 ;
	    RECT 1490.1000 589.5000 1491.0000 592.5000 ;
	    RECT 1492.2001 590.4000 1493.4000 591.6000 ;
	    RECT 1463.4000 589.2000 1464.6000 589.5000 ;
	    RECT 1492.2001 589.2000 1493.4000 589.5000 ;
	    RECT 1434.6000 587.4000 1435.8000 588.6000 ;
	    RECT 1449.0000 588.4500 1450.2001 588.6000 ;
	    RECT 1458.6000 588.4500 1459.8000 588.6000 ;
	    RECT 1449.0000 587.5500 1459.8000 588.4500 ;
	    RECT 1449.0000 587.4000 1450.2001 587.5500 ;
	    RECT 1458.6000 587.4000 1459.8000 587.5500 ;
	    RECT 1465.8000 588.4500 1467.0000 588.6000 ;
	    RECT 1487.4000 588.4500 1488.6000 588.6000 ;
	    RECT 1465.8000 587.5500 1488.6000 588.4500 ;
	    RECT 1465.8000 587.4000 1467.0000 587.5500 ;
	    RECT 1487.4000 587.4000 1488.6000 587.5500 ;
	    RECT 1489.8000 587.4000 1491.0000 588.6000 ;
	    RECT 1497.0000 587.4000 1498.2001 588.6000 ;
	    RECT 1521.0000 587.7000 1522.2001 599.7000 ;
	    RECT 1524.9000 588.6000 1526.1000 599.7000 ;
	    RECT 1527.3000 593.7000 1528.5000 599.7000 ;
	    RECT 1542.6000 593.7000 1543.8000 599.7000 ;
	    RECT 1527.0000 590.4000 1528.2001 591.6000 ;
	    RECT 1527.3000 589.5000 1528.2001 590.4000 ;
	    RECT 1524.9000 587.7000 1526.4000 588.6000 ;
	    RECT 1297.8000 586.2000 1299.0000 586.5000 ;
	    RECT 1259.4000 585.4500 1260.6000 585.6000 ;
	    RECT 1271.4000 585.4500 1272.6000 585.6000 ;
	    RECT 1259.4000 584.5500 1272.6000 585.4500 ;
	    RECT 1259.4000 584.4000 1260.6000 584.5500 ;
	    RECT 1271.4000 584.4000 1272.6000 584.5500 ;
	    RECT 1300.2001 584.4000 1301.4000 585.6000 ;
	    RECT 1302.3000 584.4000 1302.6000 585.6000 ;
	    RECT 1218.6000 581.4000 1219.8000 582.6000 ;
	    RECT 1242.6000 581.4000 1243.8000 582.6000 ;
	    RECT 1244.7001 580.8000 1245.0000 582.3000 ;
	    RECT 1247.1000 581.4000 1248.9000 582.6000 ;
	    RECT 1249.8000 582.4500 1251.0000 582.6000 ;
	    RECT 1261.8000 582.4500 1263.0000 582.6000 ;
	    RECT 1249.8000 581.5500 1263.0000 582.4500 ;
	    RECT 1249.8000 581.4000 1251.0000 581.5500 ;
	    RECT 1261.8000 581.4000 1263.0000 581.5500 ;
	    RECT 1264.2001 582.4500 1265.4000 582.6000 ;
	    RECT 1269.0000 582.4500 1270.2001 582.6000 ;
	    RECT 1264.2001 581.5500 1270.2001 582.4500 ;
	    RECT 1264.2001 581.4000 1265.4000 581.5500 ;
	    RECT 1269.0000 581.4000 1270.2001 581.5500 ;
	    RECT 1218.6000 580.2000 1219.8000 580.5000 ;
	    RECT 1242.9000 579.3000 1248.3000 579.9000 ;
	    RECT 1249.8000 579.3000 1250.7001 580.5000 ;
	    RECT 1269.0000 580.2000 1270.2001 580.5000 ;
	    RECT 1271.4000 579.3000 1272.6000 583.5000 ;
	    RECT 1305.0000 582.6000 1305.9000 586.5000 ;
	    RECT 1331.4000 586.2000 1332.6000 586.5000 ;
	    RECT 1333.8000 584.4000 1335.0000 585.6000 ;
	    RECT 1335.9000 584.4000 1336.2001 585.6000 ;
	    RECT 1338.6000 582.6000 1339.5000 586.5000 ;
	    RECT 1372.2001 586.2000 1373.4000 586.5000 ;
	    RECT 1374.6000 584.4000 1375.8000 585.6000 ;
	    RECT 1376.7001 584.4000 1377.0000 585.6000 ;
	    RECT 1379.4000 582.6000 1380.3000 586.5000 ;
	    RECT 1403.4000 586.2000 1404.6000 586.5000 ;
	    RECT 1405.8000 584.4000 1407.0000 585.6000 ;
	    RECT 1407.9000 584.4000 1408.2001 585.6000 ;
	    RECT 1410.6000 582.6000 1411.5000 586.5000 ;
	    RECT 1458.6000 586.2000 1459.8000 586.5000 ;
	    RECT 1432.2001 584.4000 1433.4000 585.6000 ;
	    RECT 1461.0000 584.4000 1462.2001 585.6000 ;
	    RECT 1463.1000 584.4000 1463.4000 585.6000 ;
	    RECT 1303.5000 582.3000 1305.9000 582.6000 ;
	    RECT 1337.1000 582.3000 1339.5000 582.6000 ;
	    RECT 1377.9000 582.3000 1380.3000 582.6000 ;
	    RECT 1409.1000 582.3000 1411.5000 582.6000 ;
	    RECT 1168.2001 573.3000 1169.4000 579.0000 ;
	    RECT 1170.6000 573.3000 1171.8000 576.3000 ;
	    RECT 1189.8000 573.3000 1191.0000 579.3000 ;
	    RECT 1192.2001 578.4000 1194.9000 579.3000 ;
	    RECT 1193.7001 573.3000 1194.9000 578.4000 ;
	    RECT 1214.7001 578.4000 1217.4000 579.3000 ;
	    RECT 1214.7001 573.3000 1215.9000 578.4000 ;
	    RECT 1218.6000 573.3000 1219.8000 579.3000 ;
	    RECT 1242.6000 579.0000 1248.6000 579.3000 ;
	    RECT 1242.6000 573.3000 1243.8000 579.0000 ;
	    RECT 1245.0000 573.3000 1246.2001 578.1000 ;
	    RECT 1247.4000 573.3000 1248.6000 579.0000 ;
	    RECT 1249.8000 573.3000 1251.0000 579.3000 ;
	    RECT 1269.0000 573.3000 1270.2001 579.3000 ;
	    RECT 1271.4000 578.4000 1274.1000 579.3000 ;
	    RECT 1272.9000 573.3000 1274.1000 578.4000 ;
	    RECT 1297.8000 573.3000 1299.0000 582.3000 ;
	    RECT 1303.2001 581.7000 1305.9000 582.3000 ;
	    RECT 1303.2001 573.3000 1304.4000 581.7000 ;
	    RECT 1331.4000 573.3000 1332.6000 582.3000 ;
	    RECT 1336.8000 581.7000 1339.5000 582.3000 ;
	    RECT 1336.8000 573.3000 1338.0000 581.7000 ;
	    RECT 1372.2001 573.3000 1373.4000 582.3000 ;
	    RECT 1377.6000 581.7000 1380.3000 582.3000 ;
	    RECT 1377.6000 573.3000 1378.8000 581.7000 ;
	    RECT 1403.4000 573.3000 1404.6000 582.3000 ;
	    RECT 1408.8000 581.7000 1411.5000 582.3000 ;
	    RECT 1417.8000 582.4500 1419.0000 582.6000 ;
	    RECT 1429.8000 582.4500 1431.0000 582.6000 ;
	    RECT 1408.8000 573.3000 1410.0000 581.7000 ;
	    RECT 1417.8000 581.5500 1431.0000 582.4500 ;
	    RECT 1417.8000 581.4000 1419.0000 581.5500 ;
	    RECT 1429.8000 581.4000 1431.0000 581.5500 ;
	    RECT 1429.8000 580.2000 1431.0000 580.5000 ;
	    RECT 1432.2001 579.3000 1433.4000 583.5000 ;
	    RECT 1465.8000 582.6000 1466.7001 586.5000 ;
	    RECT 1464.3000 582.3000 1466.7001 582.6000 ;
	    RECT 1429.8000 573.3000 1431.0000 579.3000 ;
	    RECT 1432.2001 578.4000 1434.9000 579.3000 ;
	    RECT 1433.7001 573.3000 1434.9000 578.4000 ;
	    RECT 1458.6000 573.3000 1459.8000 582.3000 ;
	    RECT 1464.0000 581.7000 1466.7001 582.3000 ;
	    RECT 1490.1000 582.6000 1491.0000 586.5000 ;
	    RECT 1497.0000 586.2000 1498.2001 586.5000 ;
	    RECT 1493.4000 584.4000 1493.7001 585.6000 ;
	    RECT 1494.6000 584.4000 1495.8000 585.6000 ;
	    RECT 1501.8000 585.4500 1503.0000 585.6000 ;
	    RECT 1523.4000 585.4500 1524.6000 585.6000 ;
	    RECT 1501.8000 584.5500 1524.6000 585.4500 ;
	    RECT 1501.8000 584.4000 1503.0000 584.5500 ;
	    RECT 1523.4000 584.4000 1524.6000 584.5500 ;
	    RECT 1523.4000 583.2000 1524.6000 583.5000 ;
	    RECT 1525.5000 582.6000 1526.4000 587.7000 ;
	    RECT 1528.2001 588.4500 1529.4000 588.6000 ;
	    RECT 1533.0000 588.4500 1534.2001 588.6000 ;
	    RECT 1528.2001 587.5500 1534.2001 588.4500 ;
	    RECT 1528.2001 587.4000 1529.4000 587.5500 ;
	    RECT 1533.0000 587.4000 1534.2001 587.5500 ;
	    RECT 1545.0000 583.5000 1546.2001 599.7000 ;
	    RECT 1490.1000 582.3000 1492.5000 582.6000 ;
	    RECT 1490.1000 581.7000 1492.8000 582.3000 ;
	    RECT 1464.0000 573.3000 1465.2001 581.7000 ;
	    RECT 1491.6000 573.3000 1492.8000 581.7000 ;
	    RECT 1497.0000 573.3000 1498.2001 582.3000 ;
	    RECT 1521.0000 581.4000 1522.2001 582.6000 ;
	    RECT 1523.1000 580.8000 1523.4000 582.3000 ;
	    RECT 1525.5000 581.4000 1527.3000 582.6000 ;
	    RECT 1528.2001 582.4500 1529.4000 582.6000 ;
	    RECT 1537.8000 582.4500 1539.0000 582.6000 ;
	    RECT 1528.2001 581.5500 1539.0000 582.4500 ;
	    RECT 1528.2001 581.4000 1529.4000 581.5500 ;
	    RECT 1537.8000 581.4000 1539.0000 581.5500 ;
	    RECT 1545.0000 581.4000 1546.2001 582.6000 ;
	    RECT 1521.3000 579.3000 1526.7001 579.9000 ;
	    RECT 1528.2001 579.3000 1529.1000 580.5000 ;
	    RECT 1521.0000 579.0000 1527.0000 579.3000 ;
	    RECT 1521.0000 573.3000 1522.2001 579.0000 ;
	    RECT 1523.4000 573.3000 1524.6000 578.1000 ;
	    RECT 1525.8000 573.3000 1527.0000 579.0000 ;
	    RECT 1528.2001 573.3000 1529.4000 579.3000 ;
	    RECT 1542.6000 578.4000 1543.8000 579.6000 ;
	    RECT 1542.6000 577.2000 1543.8000 577.5000 ;
	    RECT 1542.6000 573.3000 1543.8000 576.3000 ;
	    RECT 1545.0000 573.3000 1546.2001 580.5000 ;
	    RECT 1.2000 570.6000 1569.0000 572.4000 ;
	    RECT 18.6000 562.5000 19.8000 569.7000 ;
	    RECT 21.0000 563.7000 22.2000 569.7000 ;
	    RECT 23.4000 562.8000 24.6000 569.7000 ;
	    RECT 49.8000 563.7000 51.0000 569.7000 ;
	    RECT 52.2000 564.0000 53.4000 569.7000 ;
	    RECT 54.6000 564.9000 55.8000 569.7000 ;
	    RECT 57.0000 564.0000 58.2000 569.7000 ;
	    RECT 52.2000 563.7000 58.2000 564.0000 ;
	    RECT 21.3000 561.9000 24.6000 562.8000 ;
	    RECT 50.1000 562.5000 51.0000 563.7000 ;
	    RECT 52.5000 563.1000 57.9000 563.7000 ;
	    RECT 69.0000 562.5000 70.2000 569.7000 ;
	    RECT 71.4000 566.7000 72.6000 569.7000 ;
	    RECT 71.4000 565.5000 72.6000 565.8000 ;
	    RECT 71.4000 564.4500 72.6000 564.6000 ;
	    RECT 93.0000 564.4500 94.2000 564.6000 ;
	    RECT 71.4000 563.5500 94.2000 564.4500 ;
	    RECT 95.4000 563.7000 96.6000 569.7000 ;
	    RECT 97.8000 564.0000 99.0000 569.7000 ;
	    RECT 100.2000 564.9000 101.4000 569.7000 ;
	    RECT 102.6000 564.0000 103.8000 569.7000 ;
	    RECT 117.0000 566.7000 118.2000 569.7000 ;
	    RECT 117.0000 565.5000 118.2000 565.8000 ;
	    RECT 97.8000 563.7000 103.8000 564.0000 ;
	    RECT 71.4000 563.4000 72.6000 563.5500 ;
	    RECT 93.0000 563.4000 94.2000 563.5500 ;
	    RECT 95.7000 562.5000 96.6000 563.7000 ;
	    RECT 98.1000 563.1000 103.5000 563.7000 ;
	    RECT 117.0000 563.4000 118.2000 564.6000 ;
	    RECT 119.4000 562.5000 120.6000 569.7000 ;
	    RECT 131.4000 566.7000 132.6000 569.7000 ;
	    RECT 131.4000 565.5000 132.6000 565.8000 ;
	    RECT 131.4000 563.4000 132.6000 564.6000 ;
	    RECT 133.8000 562.5000 135.0000 569.7000 ;
	    RECT 18.6000 560.4000 19.8000 561.6000 ;
	    RECT 18.6000 558.6000 19.8000 559.5000 ;
	    RECT 18.6000 555.3000 19.5000 558.6000 ;
	    RECT 21.3000 557.4000 22.2000 561.9000 ;
	    RECT 49.8000 560.4000 51.0000 561.6000 ;
	    RECT 51.9000 560.4000 53.7000 561.6000 ;
	    RECT 55.8000 560.7000 56.1000 562.2000 ;
	    RECT 57.0000 560.4000 58.2000 561.6000 ;
	    RECT 69.0000 561.4500 70.2000 561.6000 ;
	    RECT 59.5500 560.5500 70.2000 561.4500 ;
	    RECT 23.4000 559.5000 24.6000 559.8000 ;
	    RECT 23.4000 557.4000 24.6000 558.6000 ;
	    RECT 20.4000 556.2000 22.2000 557.4000 ;
	    RECT 21.3000 555.3000 22.2000 556.2000 ;
	    RECT 47.4000 555.4500 48.6000 555.6000 ;
	    RECT 49.8000 555.4500 51.0000 555.6000 ;
	    RECT 18.6000 543.3000 19.8000 555.3000 ;
	    RECT 21.3000 554.4000 24.6000 555.3000 ;
	    RECT 47.4000 554.5500 51.0000 555.4500 ;
	    RECT 47.4000 554.4000 48.6000 554.5500 ;
	    RECT 49.8000 554.4000 51.0000 554.5500 ;
	    RECT 52.8000 555.3000 53.7000 560.4000 ;
	    RECT 54.6000 559.5000 55.8000 559.8000 ;
	    RECT 54.6000 558.4500 55.8000 558.6000 ;
	    RECT 59.5500 558.4500 60.4500 560.5500 ;
	    RECT 69.0000 560.4000 70.2000 560.5500 ;
	    RECT 95.4000 560.4000 96.6000 561.6000 ;
	    RECT 97.5000 560.4000 99.3000 561.6000 ;
	    RECT 101.4000 560.7000 101.7000 562.2000 ;
	    RECT 102.6000 560.4000 103.8000 561.6000 ;
	    RECT 119.4000 561.4500 120.6000 561.6000 ;
	    RECT 129.0000 561.4500 130.2000 561.6000 ;
	    RECT 119.4000 560.5500 130.2000 561.4500 ;
	    RECT 119.4000 560.4000 120.6000 560.5500 ;
	    RECT 129.0000 560.4000 130.2000 560.5500 ;
	    RECT 133.8000 561.4500 135.0000 561.6000 ;
	    RECT 258.6000 561.4500 259.8000 561.6000 ;
	    RECT 133.8000 560.5500 259.8000 561.4500 ;
	    RECT 133.8000 560.4000 135.0000 560.5500 ;
	    RECT 258.6000 560.4000 259.8000 560.5500 ;
	    RECT 265.8000 560.7000 267.0000 569.7000 ;
	    RECT 270.6000 563.7000 271.8000 569.7000 ;
	    RECT 275.4000 564.9000 276.6000 569.7000 ;
	    RECT 277.8000 565.5000 279.0000 569.7000 ;
	    RECT 280.2000 565.5000 281.4000 569.7000 ;
	    RECT 282.6000 565.5000 283.8000 569.7000 ;
	    RECT 285.0000 566.7000 286.2000 569.7000 ;
	    RECT 287.4000 565.5000 288.6000 569.7000 ;
	    RECT 289.8000 566.7000 291.0000 569.7000 ;
	    RECT 292.2000 565.5000 293.4000 569.7000 ;
	    RECT 294.6000 565.5000 295.8000 569.7000 ;
	    RECT 297.0000 565.5000 298.2000 569.7000 ;
	    RECT 299.4000 565.5000 300.6000 569.7000 ;
	    RECT 272.7000 563.7000 276.6000 564.9000 ;
	    RECT 301.8000 564.9000 303.0000 569.7000 ;
	    RECT 281.7000 563.7000 288.6000 564.6000 ;
	    RECT 272.7000 562.8000 273.9000 563.7000 ;
	    RECT 269.4000 561.6000 273.9000 562.8000 ;
	    RECT 54.6000 557.5500 60.4500 558.4500 ;
	    RECT 54.6000 557.4000 55.8000 557.5500 ;
	    RECT 52.8000 554.4000 54.3000 555.3000 ;
	    RECT 21.0000 543.3000 22.2000 553.5000 ;
	    RECT 23.4000 543.3000 24.6000 554.4000 ;
	    RECT 51.0000 552.6000 51.9000 553.5000 ;
	    RECT 51.0000 551.4000 52.2000 552.6000 ;
	    RECT 50.7000 543.3000 51.9000 549.3000 ;
	    RECT 53.1000 543.3000 54.3000 554.4000 ;
	    RECT 57.0000 543.3000 58.2000 555.3000 ;
	    RECT 69.0000 543.3000 70.2000 559.5000 ;
	    RECT 90.6000 555.4500 91.8000 555.6000 ;
	    RECT 95.4000 555.4500 96.6000 555.6000 ;
	    RECT 90.6000 554.5500 96.6000 555.4500 ;
	    RECT 90.6000 554.4000 91.8000 554.5500 ;
	    RECT 95.4000 554.4000 96.6000 554.5500 ;
	    RECT 98.4000 555.3000 99.3000 560.4000 ;
	    RECT 100.2000 559.5000 101.4000 559.8000 ;
	    RECT 265.8000 559.5000 279.0000 560.7000 ;
	    RECT 281.7000 560.1000 282.9000 563.7000 ;
	    RECT 287.4000 563.4000 288.6000 563.7000 ;
	    RECT 289.8000 563.4000 291.0000 564.6000 ;
	    RECT 291.9000 563.4000 292.2000 564.6000 ;
	    RECT 296.7000 563.4000 298.2000 564.6000 ;
	    RECT 301.8000 563.7000 305.4000 564.9000 ;
	    RECT 306.6000 563.7000 307.8000 569.7000 ;
	    RECT 285.0000 562.5000 286.2000 562.8000 ;
	    RECT 287.4000 562.2000 288.6000 562.5000 ;
	    RECT 285.0000 560.4000 286.2000 561.6000 ;
	    RECT 287.4000 561.3000 294.0000 562.2000 ;
	    RECT 292.8000 561.0000 294.0000 561.3000 ;
	    RECT 100.2000 558.4500 101.4000 558.6000 ;
	    RECT 107.4000 558.4500 108.6000 558.6000 ;
	    RECT 100.2000 557.5500 108.6000 558.4500 ;
	    RECT 100.2000 557.4000 101.4000 557.5500 ;
	    RECT 107.4000 557.4000 108.6000 557.5500 ;
	    RECT 98.4000 554.4000 99.9000 555.3000 ;
	    RECT 96.6000 552.6000 97.5000 553.5000 ;
	    RECT 96.6000 551.4000 97.8000 552.6000 ;
	    RECT 71.4000 543.3000 72.6000 549.3000 ;
	    RECT 96.3000 543.3000 97.5000 549.3000 ;
	    RECT 98.7000 543.3000 99.9000 554.4000 ;
	    RECT 102.6000 543.3000 103.8000 555.3000 ;
	    RECT 117.0000 543.3000 118.2000 549.3000 ;
	    RECT 119.4000 543.3000 120.6000 559.5000 ;
	    RECT 131.4000 543.3000 132.6000 549.3000 ;
	    RECT 133.8000 543.3000 135.0000 559.5000 ;
	    RECT 265.8000 551.1000 267.0000 559.5000 ;
	    RECT 279.9000 558.9000 282.9000 560.1000 ;
	    RECT 288.6000 558.9000 293.4000 560.1000 ;
	    RECT 297.0000 559.2000 298.2000 563.4000 ;
	    RECT 304.2000 562.8000 305.4000 563.7000 ;
	    RECT 304.2000 561.9000 306.9000 562.8000 ;
	    RECT 305.7000 560.1000 306.9000 561.9000 ;
	    RECT 311.4000 561.9000 312.6000 569.7000 ;
	    RECT 313.8000 564.0000 315.0000 569.7000 ;
	    RECT 316.2000 566.7000 317.4000 569.7000 ;
	    RECT 313.8000 562.8000 315.3000 564.0000 ;
	    RECT 311.4000 561.0000 313.2000 561.9000 ;
	    RECT 305.7000 558.9000 311.4000 560.1000 ;
	    RECT 267.9000 558.0000 269.1000 558.3000 ;
	    RECT 267.9000 557.1000 274.5000 558.0000 ;
	    RECT 275.4000 557.4000 276.6000 558.6000 ;
	    RECT 301.8000 558.0000 303.0000 558.9000 ;
	    RECT 312.3000 558.0000 313.2000 561.0000 ;
	    RECT 277.5000 557.1000 303.0000 558.0000 ;
	    RECT 312.0000 557.1000 313.2000 558.0000 ;
	    RECT 309.9000 556.2000 311.1000 556.5000 ;
	    RECT 270.6000 554.4000 271.8000 555.6000 ;
	    RECT 272.7000 555.3000 311.1000 556.2000 ;
	    RECT 275.7000 555.0000 276.9000 555.3000 ;
	    RECT 312.0000 554.4000 312.9000 557.1000 ;
	    RECT 314.1000 556.2000 315.3000 562.8000 ;
	    RECT 328.2000 562.5000 329.4000 569.7000 ;
	    RECT 330.6000 566.7000 331.8000 569.7000 ;
	    RECT 330.6000 565.5000 331.8000 565.8000 ;
	    RECT 330.6000 563.4000 331.8000 564.6000 ;
	    RECT 349.8000 562.8000 351.0000 569.7000 ;
	    RECT 352.2000 563.7000 353.4000 569.7000 ;
	    RECT 349.8000 561.9000 353.1000 562.8000 ;
	    RECT 354.6000 562.5000 355.8000 569.7000 ;
	    RECT 373.8000 563.7000 375.0000 569.7000 ;
	    RECT 377.7000 564.6000 378.9000 569.7000 ;
	    RECT 376.2000 563.7000 378.9000 564.6000 ;
	    RECT 373.8000 562.5000 375.0000 562.8000 ;
	    RECT 328.2000 561.4500 329.4000 561.6000 ;
	    RECT 335.4000 561.4500 336.6000 561.6000 ;
	    RECT 328.2000 560.5500 336.6000 561.4500 ;
	    RECT 328.2000 560.4000 329.4000 560.5500 ;
	    RECT 335.4000 560.4000 336.6000 560.5500 ;
	    RECT 349.8000 559.5000 351.0000 559.8000 ;
	    RECT 280.2000 554.1000 281.4000 554.4000 ;
	    RECT 273.3000 553.5000 281.4000 554.1000 ;
	    RECT 272.1000 553.2000 281.4000 553.5000 ;
	    RECT 282.9000 553.5000 295.8000 554.4000 ;
	    RECT 268.2000 552.0000 270.6000 553.2000 ;
	    RECT 272.1000 552.3000 274.2000 553.2000 ;
	    RECT 282.9000 552.3000 283.8000 553.5000 ;
	    RECT 294.6000 553.2000 295.8000 553.5000 ;
	    RECT 299.4000 553.5000 312.9000 554.4000 ;
	    RECT 313.8000 555.0000 315.3000 556.2000 ;
	    RECT 313.8000 553.5000 315.0000 555.0000 ;
	    RECT 299.4000 553.2000 300.6000 553.5000 ;
	    RECT 269.7000 551.4000 270.6000 552.0000 ;
	    RECT 275.1000 551.4000 283.8000 552.3000 ;
	    RECT 284.7000 551.4000 288.6000 552.6000 ;
	    RECT 265.8000 550.2000 268.8000 551.1000 ;
	    RECT 269.7000 550.2000 276.0000 551.4000 ;
	    RECT 267.9000 549.3000 268.8000 550.2000 ;
	    RECT 265.8000 543.3000 267.0000 549.3000 ;
	    RECT 267.9000 548.4000 269.4000 549.3000 ;
	    RECT 268.2000 543.3000 269.4000 548.4000 ;
	    RECT 270.6000 542.4000 271.8000 549.3000 ;
	    RECT 273.0000 543.3000 274.2000 550.2000 ;
	    RECT 275.4000 543.3000 276.6000 549.3000 ;
	    RECT 277.8000 543.3000 279.0000 547.5000 ;
	    RECT 280.2000 543.3000 281.4000 547.5000 ;
	    RECT 282.6000 543.3000 283.8000 550.5000 ;
	    RECT 285.0000 543.3000 286.2000 549.3000 ;
	    RECT 287.4000 543.3000 288.6000 550.5000 ;
	    RECT 289.8000 543.3000 291.0000 549.3000 ;
	    RECT 292.2000 543.3000 293.4000 552.6000 ;
	    RECT 304.2000 551.4000 308.1000 552.6000 ;
	    RECT 297.0000 550.2000 303.3000 551.4000 ;
	    RECT 294.6000 543.3000 295.8000 547.5000 ;
	    RECT 297.0000 543.3000 298.2000 547.5000 ;
	    RECT 299.4000 543.3000 300.6000 547.5000 ;
	    RECT 301.8000 543.3000 303.0000 549.3000 ;
	    RECT 304.2000 543.3000 305.4000 551.4000 ;
	    RECT 312.0000 551.1000 312.9000 553.5000 ;
	    RECT 313.8000 552.4500 315.0000 552.6000 ;
	    RECT 316.2000 552.4500 317.4000 552.6000 ;
	    RECT 313.8000 551.5500 317.4000 552.4500 ;
	    RECT 313.8000 551.4000 315.0000 551.5500 ;
	    RECT 316.2000 551.4000 317.4000 551.5500 ;
	    RECT 309.0000 550.2000 312.9000 551.1000 ;
	    RECT 306.6000 543.3000 307.8000 549.3000 ;
	    RECT 309.0000 543.3000 310.2000 550.2000 ;
	    RECT 311.4000 543.3000 312.6000 549.3000 ;
	    RECT 313.8000 543.3000 315.0000 550.5000 ;
	    RECT 316.2000 543.3000 317.4000 549.3000 ;
	    RECT 328.2000 543.3000 329.4000 559.5000 ;
	    RECT 340.2000 558.4500 341.4000 558.6000 ;
	    RECT 349.8000 558.4500 351.0000 558.6000 ;
	    RECT 340.2000 557.5500 351.0000 558.4500 ;
	    RECT 340.2000 557.4000 341.4000 557.5500 ;
	    RECT 349.8000 557.4000 351.0000 557.5500 ;
	    RECT 352.2000 557.4000 353.1000 561.9000 ;
	    RECT 354.6000 561.4500 355.8000 561.6000 ;
	    RECT 357.0000 561.4500 358.2000 561.6000 ;
	    RECT 373.8000 561.4500 375.0000 561.6000 ;
	    RECT 354.6000 560.5500 375.0000 561.4500 ;
	    RECT 354.6000 560.4000 355.8000 560.5500 ;
	    RECT 357.0000 560.4000 358.2000 560.5500 ;
	    RECT 373.8000 560.4000 375.0000 560.5500 ;
	    RECT 376.2000 559.5000 377.4000 563.7000 ;
	    RECT 513.0000 560.7000 514.2000 569.7000 ;
	    RECT 517.8000 563.7000 519.0000 569.7000 ;
	    RECT 522.6000 564.9000 523.8000 569.7000 ;
	    RECT 525.0000 565.5000 526.2000 569.7000 ;
	    RECT 527.4000 565.5000 528.6000 569.7000 ;
	    RECT 529.8000 565.5000 531.0000 569.7000 ;
	    RECT 532.2000 566.7000 533.4000 569.7000 ;
	    RECT 534.6000 565.5000 535.8000 569.7000 ;
	    RECT 537.0000 566.7000 538.2000 569.7000 ;
	    RECT 539.4000 565.5000 540.6000 569.7000 ;
	    RECT 541.8000 565.5000 543.0000 569.7000 ;
	    RECT 544.2000 565.5000 545.4000 569.7000 ;
	    RECT 546.6000 565.5000 547.8000 569.7000 ;
	    RECT 519.9000 563.7000 523.8000 564.9000 ;
	    RECT 549.0000 564.9000 550.2000 569.7000 ;
	    RECT 528.9000 563.7000 535.8000 564.6000 ;
	    RECT 519.9000 562.8000 521.1000 563.7000 ;
	    RECT 516.6000 561.6000 521.1000 562.8000 ;
	    RECT 513.0000 559.5000 526.2000 560.7000 ;
	    RECT 528.9000 560.1000 530.1000 563.7000 ;
	    RECT 534.6000 563.4000 535.8000 563.7000 ;
	    RECT 537.0000 563.4000 538.2000 564.6000 ;
	    RECT 539.1000 563.4000 539.4000 564.6000 ;
	    RECT 543.9000 563.4000 545.4000 564.6000 ;
	    RECT 549.0000 563.7000 552.6000 564.9000 ;
	    RECT 553.8000 563.7000 555.0000 569.7000 ;
	    RECT 532.2000 562.5000 533.4000 562.8000 ;
	    RECT 534.6000 562.2000 535.8000 562.5000 ;
	    RECT 532.2000 560.4000 533.4000 561.6000 ;
	    RECT 534.6000 561.3000 541.2000 562.2000 ;
	    RECT 540.0000 561.0000 541.2000 561.3000 ;
	    RECT 354.6000 558.6000 355.8000 559.5000 ;
	    RECT 352.2000 556.2000 354.0000 557.4000 ;
	    RECT 352.2000 555.3000 353.1000 556.2000 ;
	    RECT 354.9000 555.3000 355.8000 558.6000 ;
	    RECT 366.6000 558.4500 367.8000 558.6000 ;
	    RECT 376.2000 558.4500 377.4000 558.6000 ;
	    RECT 366.6000 557.5500 377.4000 558.4500 ;
	    RECT 366.6000 557.4000 367.8000 557.5500 ;
	    RECT 376.2000 557.4000 377.4000 557.5500 ;
	    RECT 349.8000 554.4000 353.1000 555.3000 ;
	    RECT 330.6000 543.3000 331.8000 549.3000 ;
	    RECT 349.8000 543.3000 351.0000 554.4000 ;
	    RECT 352.2000 543.3000 353.4000 553.5000 ;
	    RECT 354.6000 543.3000 355.8000 555.3000 ;
	    RECT 373.8000 543.3000 375.0000 549.3000 ;
	    RECT 376.2000 543.3000 377.4000 556.5000 ;
	    RECT 378.6000 555.4500 379.8000 555.6000 ;
	    RECT 510.6000 555.4500 511.8000 555.6000 ;
	    RECT 378.6000 554.5500 511.8000 555.4500 ;
	    RECT 378.6000 554.4000 379.8000 554.5500 ;
	    RECT 510.6000 554.4000 511.8000 554.5500 ;
	    RECT 378.6000 553.2000 379.8000 553.5000 ;
	    RECT 513.0000 551.1000 514.2000 559.5000 ;
	    RECT 527.1000 558.9000 530.1000 560.1000 ;
	    RECT 535.8000 558.9000 540.6000 560.1000 ;
	    RECT 544.2000 559.2000 545.4000 563.4000 ;
	    RECT 551.4000 562.8000 552.6000 563.7000 ;
	    RECT 551.4000 561.9000 554.1000 562.8000 ;
	    RECT 552.9000 560.1000 554.1000 561.9000 ;
	    RECT 558.6000 561.9000 559.8000 569.7000 ;
	    RECT 561.0000 564.0000 562.2000 569.7000 ;
	    RECT 563.4000 566.7000 564.6000 569.7000 ;
	    RECT 583.5000 564.6000 584.7000 569.7000 ;
	    RECT 561.0000 562.8000 562.5000 564.0000 ;
	    RECT 583.5000 563.7000 586.2000 564.6000 ;
	    RECT 587.4000 563.7000 588.6000 569.7000 ;
	    RECT 601.8000 566.7000 603.0000 569.7000 ;
	    RECT 601.8000 565.5000 603.0000 565.8000 ;
	    RECT 558.6000 561.0000 560.4000 561.9000 ;
	    RECT 552.9000 558.9000 558.6000 560.1000 ;
	    RECT 515.1000 558.0000 516.3000 558.3000 ;
	    RECT 515.1000 557.1000 521.7000 558.0000 ;
	    RECT 522.6000 557.4000 523.8000 558.6000 ;
	    RECT 549.0000 558.0000 550.2000 558.9000 ;
	    RECT 559.5000 558.0000 560.4000 561.0000 ;
	    RECT 524.7000 557.1000 550.2000 558.0000 ;
	    RECT 559.2000 557.1000 560.4000 558.0000 ;
	    RECT 557.1000 556.2000 558.3000 556.5000 ;
	    RECT 515.4000 555.4500 516.6000 555.6000 ;
	    RECT 517.8000 555.4500 519.0000 555.6000 ;
	    RECT 515.4000 554.5500 519.0000 555.4500 ;
	    RECT 519.9000 555.3000 558.3000 556.2000 ;
	    RECT 522.9000 555.0000 524.1000 555.3000 ;
	    RECT 515.4000 554.4000 516.6000 554.5500 ;
	    RECT 517.8000 554.4000 519.0000 554.5500 ;
	    RECT 559.2000 554.4000 560.1000 557.1000 ;
	    RECT 561.3000 556.2000 562.5000 562.8000 ;
	    RECT 585.0000 559.5000 586.2000 563.7000 ;
	    RECT 601.8000 563.4000 603.0000 564.6000 ;
	    RECT 587.4000 562.5000 588.6000 562.8000 ;
	    RECT 604.2000 562.5000 605.4000 569.7000 ;
	    RECT 616.2000 562.5000 617.4000 569.7000 ;
	    RECT 618.6000 566.7000 619.8000 569.7000 ;
	    RECT 618.6000 565.5000 619.8000 565.8000 ;
	    RECT 638.7000 564.6000 639.9000 569.7000 ;
	    RECT 618.6000 563.4000 619.8000 564.6000 ;
	    RECT 638.7000 563.7000 641.4000 564.6000 ;
	    RECT 642.6000 563.7000 643.8000 569.7000 ;
	    RECT 676.2000 563.7000 677.4000 569.7000 ;
	    RECT 678.6000 564.0000 679.8000 569.7000 ;
	    RECT 681.0000 564.9000 682.2000 569.7000 ;
	    RECT 683.4000 564.0000 684.6000 569.7000 ;
	    RECT 678.6000 563.7000 684.6000 564.0000 ;
	    RECT 587.4000 560.4000 588.6000 561.6000 ;
	    RECT 597.0000 561.4500 598.2000 561.6000 ;
	    RECT 601.8000 561.4500 603.0000 561.6000 ;
	    RECT 604.2000 561.4500 605.4000 561.6000 ;
	    RECT 597.0000 560.5500 605.4000 561.4500 ;
	    RECT 597.0000 560.4000 598.2000 560.5500 ;
	    RECT 601.8000 560.4000 603.0000 560.5500 ;
	    RECT 604.2000 560.4000 605.4000 560.5500 ;
	    RECT 616.2000 561.4500 617.4000 561.6000 ;
	    RECT 633.0000 561.4500 634.2000 561.6000 ;
	    RECT 616.2000 560.5500 634.2000 561.4500 ;
	    RECT 616.2000 560.4000 617.4000 560.5500 ;
	    RECT 633.0000 560.4000 634.2000 560.5500 ;
	    RECT 640.2000 559.5000 641.4000 563.7000 ;
	    RECT 642.6000 562.5000 643.8000 562.8000 ;
	    RECT 676.5000 562.5000 677.4000 563.7000 ;
	    RECT 678.9000 563.1000 684.3000 563.7000 ;
	    RECT 695.4000 562.5000 696.6000 569.7000 ;
	    RECT 697.8000 566.7000 699.0000 569.7000 ;
	    RECT 712.2000 566.7000 713.4000 569.7000 ;
	    RECT 697.8000 565.5000 699.0000 565.8000 ;
	    RECT 712.2000 565.5000 713.4000 565.8000 ;
	    RECT 697.8000 564.4500 699.0000 564.6000 ;
	    RECT 707.4000 564.4500 708.6000 564.6000 ;
	    RECT 697.8000 563.5500 708.6000 564.4500 ;
	    RECT 697.8000 563.4000 699.0000 563.5500 ;
	    RECT 707.4000 563.4000 708.6000 563.5500 ;
	    RECT 712.2000 563.4000 713.4000 564.6000 ;
	    RECT 714.6000 562.5000 715.8000 569.7000 ;
	    RECT 642.6000 560.4000 643.8000 561.6000 ;
	    RECT 676.2000 560.4000 677.4000 561.6000 ;
	    RECT 678.3000 560.4000 680.1000 561.6000 ;
	    RECT 682.2000 560.7000 682.5000 562.2000 ;
	    RECT 683.4000 560.4000 684.6000 561.6000 ;
	    RECT 695.4000 561.4500 696.6000 561.6000 ;
	    RECT 685.9500 560.5500 696.6000 561.4500 ;
	    RECT 570.6000 558.4500 571.8000 558.6000 ;
	    RECT 585.0000 558.4500 586.2000 558.6000 ;
	    RECT 570.6000 557.5500 586.2000 558.4500 ;
	    RECT 570.6000 557.4000 571.8000 557.5500 ;
	    RECT 585.0000 557.4000 586.2000 557.5500 ;
	    RECT 527.4000 554.1000 528.6000 554.4000 ;
	    RECT 520.5000 553.5000 528.6000 554.1000 ;
	    RECT 519.3000 553.2000 528.6000 553.5000 ;
	    RECT 530.1000 553.5000 543.0000 554.4000 ;
	    RECT 515.4000 552.0000 517.8000 553.2000 ;
	    RECT 519.3000 552.3000 521.4000 553.2000 ;
	    RECT 530.1000 552.3000 531.0000 553.5000 ;
	    RECT 541.8000 553.2000 543.0000 553.5000 ;
	    RECT 546.6000 553.5000 560.1000 554.4000 ;
	    RECT 561.0000 555.0000 562.5000 556.2000 ;
	    RECT 561.0000 553.5000 562.2000 555.0000 ;
	    RECT 582.6000 554.4000 583.8000 555.6000 ;
	    RECT 546.6000 553.2000 547.8000 553.5000 ;
	    RECT 516.9000 551.4000 517.8000 552.0000 ;
	    RECT 522.3000 551.4000 531.0000 552.3000 ;
	    RECT 531.9000 551.4000 535.8000 552.6000 ;
	    RECT 513.0000 550.2000 516.0000 551.1000 ;
	    RECT 516.9000 550.2000 523.2000 551.4000 ;
	    RECT 515.1000 549.3000 516.0000 550.2000 ;
	    RECT 378.6000 543.3000 379.8000 549.3000 ;
	    RECT 513.0000 543.3000 514.2000 549.3000 ;
	    RECT 515.1000 548.4000 516.6000 549.3000 ;
	    RECT 515.4000 543.3000 516.6000 548.4000 ;
	    RECT 517.8000 542.4000 519.0000 549.3000 ;
	    RECT 520.2000 543.3000 521.4000 550.2000 ;
	    RECT 522.6000 543.3000 523.8000 549.3000 ;
	    RECT 525.0000 543.3000 526.2000 547.5000 ;
	    RECT 527.4000 543.3000 528.6000 547.5000 ;
	    RECT 529.8000 543.3000 531.0000 550.5000 ;
	    RECT 532.2000 543.3000 533.4000 549.3000 ;
	    RECT 534.6000 543.3000 535.8000 550.5000 ;
	    RECT 537.0000 543.3000 538.2000 549.3000 ;
	    RECT 539.4000 543.3000 540.6000 552.6000 ;
	    RECT 551.4000 551.4000 555.3000 552.6000 ;
	    RECT 544.2000 550.2000 550.5000 551.4000 ;
	    RECT 541.8000 543.3000 543.0000 547.5000 ;
	    RECT 544.2000 543.3000 545.4000 547.5000 ;
	    RECT 546.6000 543.3000 547.8000 547.5000 ;
	    RECT 549.0000 543.3000 550.2000 549.3000 ;
	    RECT 551.4000 543.3000 552.6000 551.4000 ;
	    RECT 559.2000 551.1000 560.1000 553.5000 ;
	    RECT 582.6000 553.2000 583.8000 553.5000 ;
	    RECT 561.0000 551.4000 562.2000 552.6000 ;
	    RECT 556.2000 550.2000 560.1000 551.1000 ;
	    RECT 553.8000 543.3000 555.0000 549.3000 ;
	    RECT 556.2000 543.3000 557.4000 550.2000 ;
	    RECT 558.6000 543.3000 559.8000 549.3000 ;
	    RECT 561.0000 543.3000 562.2000 550.5000 ;
	    RECT 563.4000 543.3000 564.6000 549.3000 ;
	    RECT 582.6000 543.3000 583.8000 549.3000 ;
	    RECT 585.0000 543.3000 586.2000 556.5000 ;
	    RECT 587.4000 543.3000 588.6000 549.3000 ;
	    RECT 601.8000 543.3000 603.0000 549.3000 ;
	    RECT 604.2000 543.3000 605.4000 559.5000 ;
	    RECT 616.2000 543.3000 617.4000 559.5000 ;
	    RECT 640.2000 558.4500 641.4000 558.6000 ;
	    RECT 640.2000 557.5500 677.2500 558.4500 ;
	    RECT 640.2000 557.4000 641.4000 557.5500 ;
	    RECT 637.8000 554.4000 639.0000 555.6000 ;
	    RECT 637.8000 553.2000 639.0000 553.5000 ;
	    RECT 618.6000 543.3000 619.8000 549.3000 ;
	    RECT 637.8000 543.3000 639.0000 549.3000 ;
	    RECT 640.2000 543.3000 641.4000 556.5000 ;
	    RECT 676.3500 555.6000 677.2500 557.5500 ;
	    RECT 676.2000 554.4000 677.4000 555.6000 ;
	    RECT 679.2000 555.3000 680.1000 560.4000 ;
	    RECT 681.0000 559.5000 682.2000 559.8000 ;
	    RECT 681.0000 558.4500 682.2000 558.6000 ;
	    RECT 685.9500 558.4500 686.8500 560.5500 ;
	    RECT 695.4000 560.4000 696.6000 560.5500 ;
	    RECT 714.6000 561.4500 715.8000 561.6000 ;
	    RECT 724.2000 561.4500 725.4000 561.6000 ;
	    RECT 714.6000 560.5500 725.4000 561.4500 ;
	    RECT 714.6000 560.4000 715.8000 560.5500 ;
	    RECT 724.2000 560.4000 725.4000 560.5500 ;
	    RECT 839.4000 560.7000 840.6000 569.7000 ;
	    RECT 844.2000 563.7000 845.4000 569.7000 ;
	    RECT 849.0000 564.9000 850.2000 569.7000 ;
	    RECT 851.4000 565.5000 852.6000 569.7000 ;
	    RECT 853.8000 565.5000 855.0000 569.7000 ;
	    RECT 856.2000 565.5000 857.4000 569.7000 ;
	    RECT 858.6000 566.7000 859.8000 569.7000 ;
	    RECT 861.0000 565.5000 862.2000 569.7000 ;
	    RECT 863.4000 566.7000 864.6000 569.7000 ;
	    RECT 865.8000 565.5000 867.0000 569.7000 ;
	    RECT 868.2000 565.5000 869.4000 569.7000 ;
	    RECT 870.6000 565.5000 871.8000 569.7000 ;
	    RECT 873.0000 565.5000 874.2000 569.7000 ;
	    RECT 846.3000 563.7000 850.2000 564.9000 ;
	    RECT 875.4000 564.9000 876.6000 569.7000 ;
	    RECT 855.3000 563.7000 862.2000 564.6000 ;
	    RECT 846.3000 562.8000 847.5000 563.7000 ;
	    RECT 843.0000 561.6000 847.5000 562.8000 ;
	    RECT 839.4000 559.5000 852.6000 560.7000 ;
	    RECT 855.3000 560.1000 856.5000 563.7000 ;
	    RECT 861.0000 563.4000 862.2000 563.7000 ;
	    RECT 863.4000 563.4000 864.6000 564.6000 ;
	    RECT 865.5000 563.4000 865.8000 564.6000 ;
	    RECT 870.3000 563.4000 871.8000 564.6000 ;
	    RECT 875.4000 563.7000 879.0000 564.9000 ;
	    RECT 880.2000 563.7000 881.4000 569.7000 ;
	    RECT 858.6000 562.5000 859.8000 562.8000 ;
	    RECT 861.0000 562.2000 862.2000 562.5000 ;
	    RECT 858.6000 560.4000 859.8000 561.6000 ;
	    RECT 861.0000 561.3000 867.6000 562.2000 ;
	    RECT 866.4000 561.0000 867.6000 561.3000 ;
	    RECT 681.0000 557.5500 686.8500 558.4500 ;
	    RECT 681.0000 557.4000 682.2000 557.5500 ;
	    RECT 679.2000 554.4000 680.7000 555.3000 ;
	    RECT 677.4000 552.6000 678.3000 553.5000 ;
	    RECT 677.4000 551.4000 678.6000 552.6000 ;
	    RECT 642.6000 543.3000 643.8000 549.3000 ;
	    RECT 677.1000 543.3000 678.3000 549.3000 ;
	    RECT 679.5000 543.3000 680.7000 554.4000 ;
	    RECT 683.4000 543.3000 684.6000 555.3000 ;
	    RECT 695.4000 543.3000 696.6000 559.5000 ;
	    RECT 697.8000 543.3000 699.0000 549.3000 ;
	    RECT 712.2000 543.3000 713.4000 549.3000 ;
	    RECT 714.6000 543.3000 715.8000 559.5000 ;
	    RECT 839.4000 551.1000 840.6000 559.5000 ;
	    RECT 853.5000 558.9000 856.5000 560.1000 ;
	    RECT 862.2000 558.9000 867.0000 560.1000 ;
	    RECT 870.6000 559.2000 871.8000 563.4000 ;
	    RECT 877.8000 562.8000 879.0000 563.7000 ;
	    RECT 877.8000 561.9000 880.5000 562.8000 ;
	    RECT 879.3000 560.1000 880.5000 561.9000 ;
	    RECT 885.0000 561.9000 886.2000 569.7000 ;
	    RECT 887.4000 564.0000 888.6000 569.7000 ;
	    RECT 889.8000 566.7000 891.0000 569.7000 ;
	    RECT 887.4000 562.8000 888.9000 564.0000 ;
	    RECT 885.0000 561.0000 886.8000 561.9000 ;
	    RECT 879.3000 558.9000 885.0000 560.1000 ;
	    RECT 841.5000 558.0000 842.7000 558.3000 ;
	    RECT 841.5000 557.1000 848.1000 558.0000 ;
	    RECT 849.0000 557.4000 850.2000 558.6000 ;
	    RECT 875.4000 558.0000 876.6000 558.9000 ;
	    RECT 885.9000 558.0000 886.8000 561.0000 ;
	    RECT 851.1000 557.1000 876.6000 558.0000 ;
	    RECT 885.6000 557.1000 886.8000 558.0000 ;
	    RECT 883.5000 556.2000 884.7000 556.5000 ;
	    RECT 844.2000 554.4000 845.4000 555.6000 ;
	    RECT 846.3000 555.3000 884.7000 556.2000 ;
	    RECT 849.3000 555.0000 850.5000 555.3000 ;
	    RECT 885.6000 554.4000 886.5000 557.1000 ;
	    RECT 887.7000 556.2000 888.9000 562.8000 ;
	    RECT 966.6000 562.5000 967.8000 569.7000 ;
	    RECT 969.0000 563.7000 970.2000 569.7000 ;
	    RECT 973.2000 567.6000 974.4000 569.7000 ;
	    RECT 971.4000 566.7000 974.4000 567.6000 ;
	    RECT 977.1000 566.7000 978.6000 569.7000 ;
	    RECT 979.8000 566.7000 981.0000 569.7000 ;
	    RECT 982.2000 566.7000 983.4000 569.7000 ;
	    RECT 986.1000 567.6000 987.9000 569.7000 ;
	    RECT 985.8000 566.7000 987.9000 567.6000 ;
	    RECT 971.4000 565.5000 972.6000 566.7000 ;
	    RECT 979.8000 565.8000 980.7000 566.7000 ;
	    RECT 973.8000 564.6000 975.0000 565.8000 ;
	    RECT 976.5000 564.9000 980.7000 565.8000 ;
	    RECT 985.8000 565.5000 987.0000 566.7000 ;
	    RECT 976.5000 564.6000 977.7000 564.9000 ;
	    RECT 967.8000 560.4000 968.1000 561.6000 ;
	    RECT 969.0000 560.4000 970.2000 561.6000 ;
	    RECT 974.1000 561.3000 975.0000 564.6000 ;
	    RECT 990.6000 564.0000 991.8000 569.7000 ;
	    RECT 988.5000 563.1000 989.7000 563.4000 ;
	    RECT 993.0000 563.1000 994.2000 569.7000 ;
	    RECT 1013.1000 564.6000 1014.3000 569.7000 ;
	    RECT 1013.1000 563.7000 1015.8000 564.6000 ;
	    RECT 1017.0000 563.7000 1018.2000 569.7000 ;
	    RECT 1043.4000 563.7000 1044.6000 569.7000 ;
	    RECT 1045.8000 564.0000 1047.0000 569.7000 ;
	    RECT 1048.2001 564.9000 1049.4000 569.7000 ;
	    RECT 1050.6000 564.0000 1051.8000 569.7000 ;
	    RECT 1045.8000 563.7000 1051.8000 564.0000 ;
	    RECT 988.5000 562.2000 994.2000 563.1000 ;
	    RECT 982.5000 561.3000 983.7000 561.6000 ;
	    RECT 971.1000 560.4000 984.3000 561.3000 ;
	    RECT 972.3000 560.1000 973.5000 560.4000 ;
	    RECT 969.9000 558.6000 971.1000 558.9000 ;
	    RECT 969.9000 557.7000 975.3000 558.6000 ;
	    RECT 976.2000 557.4000 977.4000 558.6000 ;
	    RECT 853.8000 554.1000 855.0000 554.4000 ;
	    RECT 846.9000 553.5000 855.0000 554.1000 ;
	    RECT 845.7000 553.2000 855.0000 553.5000 ;
	    RECT 856.5000 553.5000 869.4000 554.4000 ;
	    RECT 841.8000 552.0000 844.2000 553.2000 ;
	    RECT 845.7000 552.3000 847.8000 553.2000 ;
	    RECT 856.5000 552.3000 857.4000 553.5000 ;
	    RECT 868.2000 553.2000 869.4000 553.5000 ;
	    RECT 873.0000 553.5000 886.5000 554.4000 ;
	    RECT 887.4000 555.0000 888.9000 556.2000 ;
	    RECT 966.6000 556.5000 975.0000 556.8000 ;
	    RECT 966.6000 556.2000 975.3000 556.5000 ;
	    RECT 966.6000 555.9000 981.3000 556.2000 ;
	    RECT 887.4000 553.5000 888.6000 555.0000 ;
	    RECT 873.0000 553.2000 874.2000 553.5000 ;
	    RECT 843.3000 551.4000 844.2000 552.0000 ;
	    RECT 848.7000 551.4000 857.4000 552.3000 ;
	    RECT 858.3000 551.4000 862.2000 552.6000 ;
	    RECT 839.4000 550.2000 842.4000 551.1000 ;
	    RECT 843.3000 550.2000 849.6000 551.4000 ;
	    RECT 841.5000 549.3000 842.4000 550.2000 ;
	    RECT 839.4000 543.3000 840.6000 549.3000 ;
	    RECT 841.5000 548.4000 843.0000 549.3000 ;
	    RECT 841.8000 543.3000 843.0000 548.4000 ;
	    RECT 844.2000 542.4000 845.4000 549.3000 ;
	    RECT 846.6000 543.3000 847.8000 550.2000 ;
	    RECT 849.0000 543.3000 850.2000 549.3000 ;
	    RECT 851.4000 543.3000 852.6000 547.5000 ;
	    RECT 853.8000 543.3000 855.0000 547.5000 ;
	    RECT 856.2000 543.3000 857.4000 550.5000 ;
	    RECT 858.6000 543.3000 859.8000 549.3000 ;
	    RECT 861.0000 543.3000 862.2000 550.5000 ;
	    RECT 863.4000 543.3000 864.6000 549.3000 ;
	    RECT 865.8000 543.3000 867.0000 552.6000 ;
	    RECT 877.8000 551.4000 881.7000 552.6000 ;
	    RECT 870.6000 550.2000 876.9000 551.4000 ;
	    RECT 868.2000 543.3000 869.4000 547.5000 ;
	    RECT 870.6000 543.3000 871.8000 547.5000 ;
	    RECT 873.0000 543.3000 874.2000 547.5000 ;
	    RECT 875.4000 543.3000 876.6000 549.3000 ;
	    RECT 877.8000 543.3000 879.0000 551.4000 ;
	    RECT 885.6000 551.1000 886.5000 553.5000 ;
	    RECT 887.4000 551.4000 888.6000 552.6000 ;
	    RECT 882.6000 550.2000 886.5000 551.1000 ;
	    RECT 880.2000 543.3000 881.4000 549.3000 ;
	    RECT 882.6000 543.3000 883.8000 550.2000 ;
	    RECT 885.0000 543.3000 886.2000 549.3000 ;
	    RECT 887.4000 543.3000 888.6000 550.5000 ;
	    RECT 889.8000 543.3000 891.0000 549.3000 ;
	    RECT 966.6000 543.3000 967.8000 555.9000 ;
	    RECT 974.1000 555.3000 981.3000 555.9000 ;
	    RECT 969.0000 543.3000 970.2000 555.0000 ;
	    RECT 971.4000 553.5000 979.5000 554.4000 ;
	    RECT 971.4000 553.2000 972.6000 553.5000 ;
	    RECT 978.3000 553.2000 979.5000 553.5000 ;
	    RECT 980.4000 553.5000 981.3000 555.3000 ;
	    RECT 983.4000 555.6000 984.3000 560.4000 ;
	    RECT 993.0000 559.5000 994.2000 562.2000 ;
	    RECT 1014.6000 559.5000 1015.8000 563.7000 ;
	    RECT 1017.0000 562.5000 1018.2000 562.8000 ;
	    RECT 1043.7001 562.5000 1044.6000 563.7000 ;
	    RECT 1046.1000 563.1000 1051.5000 563.7000 ;
	    RECT 1062.6000 562.5000 1063.8000 569.7000 ;
	    RECT 1065.0000 566.7000 1066.2001 569.7000 ;
	    RECT 1065.0000 565.5000 1066.2001 565.8000 ;
	    RECT 1065.0000 564.4500 1066.2001 564.6000 ;
	    RECT 1093.8000 564.4500 1095.0000 564.6000 ;
	    RECT 1065.0000 563.5500 1095.0000 564.4500 ;
	    RECT 1096.8000 563.7000 1098.0000 569.7000 ;
	    RECT 1100.7001 563.7000 1103.1000 569.7000 ;
	    RECT 1105.8000 563.7000 1107.0000 569.7000 ;
	    RECT 1127.4000 567.4500 1128.6000 567.6000 ;
	    RECT 1134.6000 567.4500 1135.8000 567.6000 ;
	    RECT 1127.4000 566.5500 1135.8000 567.4500 ;
	    RECT 1127.4000 566.4000 1128.6000 566.5500 ;
	    RECT 1134.6000 566.4000 1135.8000 566.5500 ;
	    RECT 1137.9000 565.2000 1139.1000 569.7000 ;
	    RECT 1137.0000 563.7000 1139.1000 565.2000 ;
	    RECT 1140.3000 564.0000 1141.5000 569.7000 ;
	    RECT 1144.2001 563.7000 1145.4000 569.7000 ;
	    RECT 1065.0000 563.4000 1066.2001 563.5500 ;
	    RECT 1093.8000 563.4000 1095.0000 563.5500 ;
	    RECT 1017.0000 560.4000 1018.2000 561.6000 ;
	    RECT 1043.4000 560.4000 1044.6000 561.6000 ;
	    RECT 1045.5000 560.4000 1047.3000 561.6000 ;
	    RECT 1049.4000 560.7000 1049.7001 562.2000 ;
	    RECT 1050.6000 560.4000 1051.8000 561.6000 ;
	    RECT 1062.6000 561.4500 1063.8000 561.6000 ;
	    RECT 1053.1500 560.5500 1063.8000 561.4500 ;
	    RECT 985.8000 559.2000 987.0000 559.5000 ;
	    RECT 985.8000 558.3000 991.5000 559.2000 ;
	    RECT 990.3000 558.0000 991.5000 558.3000 ;
	    RECT 993.0000 557.4000 994.2000 558.6000 ;
	    RECT 1014.6000 558.4500 1015.8000 558.6000 ;
	    RECT 1014.6000 557.5500 1044.4501 558.4500 ;
	    RECT 1014.6000 557.4000 1015.8000 557.5500 ;
	    RECT 987.9000 557.1000 989.1000 557.4000 ;
	    RECT 987.9000 556.5000 992.1000 557.1000 ;
	    RECT 987.9000 556.2000 994.2000 556.5000 ;
	    RECT 983.4000 554.7000 987.0000 555.6000 ;
	    RECT 982.5000 553.5000 983.7000 553.8000 ;
	    RECT 980.4000 552.6000 983.7000 553.5000 ;
	    RECT 986.1000 553.2000 987.0000 554.7000 ;
	    RECT 986.1000 552.0000 988.2000 553.2000 ;
	    RECT 976.5000 551.1000 977.7000 551.4000 ;
	    RECT 980.7000 551.1000 981.9000 551.4000 ;
	    RECT 971.4000 549.3000 972.6000 550.5000 ;
	    RECT 976.5000 550.2000 981.9000 551.1000 ;
	    RECT 979.8000 549.3000 980.7000 550.2000 ;
	    RECT 985.8000 549.3000 987.0000 550.5000 ;
	    RECT 971.4000 548.4000 974.4000 549.3000 ;
	    RECT 973.2000 543.3000 974.4000 548.4000 ;
	    RECT 977.4000 543.3000 978.6000 549.3000 ;
	    RECT 979.8000 543.3000 981.0000 549.3000 ;
	    RECT 982.2000 543.3000 983.4000 549.3000 ;
	    RECT 986.1000 543.3000 987.9000 549.3000 ;
	    RECT 990.6000 543.3000 991.8000 555.3000 ;
	    RECT 993.0000 543.3000 994.2000 556.2000 ;
	    RECT 1002.6000 555.4500 1003.8000 555.6000 ;
	    RECT 1012.2000 555.4500 1013.4000 555.6000 ;
	    RECT 1002.6000 554.5500 1013.4000 555.4500 ;
	    RECT 1002.6000 554.4000 1003.8000 554.5500 ;
	    RECT 1012.2000 554.4000 1013.4000 554.5500 ;
	    RECT 1012.2000 553.2000 1013.4000 553.5000 ;
	    RECT 1012.2000 543.3000 1013.4000 549.3000 ;
	    RECT 1014.6000 543.3000 1015.8000 556.5000 ;
	    RECT 1043.5500 555.6000 1044.4501 557.5500 ;
	    RECT 1043.4000 554.4000 1044.6000 555.6000 ;
	    RECT 1046.4000 555.3000 1047.3000 560.4000 ;
	    RECT 1048.2001 559.5000 1049.4000 559.8000 ;
	    RECT 1048.2001 558.4500 1049.4000 558.6000 ;
	    RECT 1053.1500 558.4500 1054.0500 560.5500 ;
	    RECT 1062.6000 560.4000 1063.8000 560.5500 ;
	    RECT 1079.4000 561.4500 1080.6000 561.6000 ;
	    RECT 1098.6000 561.4500 1099.8000 561.6000 ;
	    RECT 1079.4000 560.5500 1099.8000 561.4500 ;
	    RECT 1079.4000 560.4000 1080.6000 560.5500 ;
	    RECT 1098.6000 560.4000 1099.8000 560.5500 ;
	    RECT 1101.3000 559.5000 1102.2001 563.7000 ;
	    RECT 1103.4000 560.4000 1104.6000 561.6000 ;
	    RECT 1137.0000 559.5000 1137.9000 563.7000 ;
	    RECT 1144.2001 563.4000 1145.1000 563.7000 ;
	    RECT 1142.4000 562.8000 1145.1000 563.4000 ;
	    RECT 1138.8000 562.5000 1145.1000 562.8000 ;
	    RECT 1138.8000 561.9000 1143.3000 562.5000 ;
	    RECT 1138.8000 561.6000 1140.0000 561.9000 ;
	    RECT 1048.2001 557.5500 1054.0500 558.4500 ;
	    RECT 1048.2001 557.4000 1049.4000 557.5500 ;
	    RECT 1046.4000 554.4000 1047.9000 555.3000 ;
	    RECT 1044.6000 552.6000 1045.5000 553.5000 ;
	    RECT 1044.6000 551.4000 1045.8000 552.6000 ;
	    RECT 1017.0000 543.3000 1018.2000 549.3000 ;
	    RECT 1044.3000 543.3000 1045.5000 549.3000 ;
	    RECT 1046.7001 543.3000 1047.9000 554.4000 ;
	    RECT 1050.6000 543.3000 1051.8000 555.3000 ;
	    RECT 1062.6000 543.3000 1063.8000 559.5000 ;
	    RECT 1098.6000 559.2000 1099.8000 559.5000 ;
	    RECT 1103.1000 558.6000 1104.3000 559.5000 ;
	    RECT 1084.2001 558.4500 1085.4000 558.6000 ;
	    RECT 1096.2001 558.4500 1097.4000 558.6000 ;
	    RECT 1084.2001 557.5500 1097.4000 558.4500 ;
	    RECT 1084.2001 557.4000 1085.4000 557.5500 ;
	    RECT 1096.2001 557.4000 1097.4000 557.5500 ;
	    RECT 1098.3000 556.8000 1098.6000 558.3000 ;
	    RECT 1101.0000 557.4000 1102.2001 558.6000 ;
	    RECT 1105.8000 558.4500 1107.0000 558.6000 ;
	    RECT 1134.6000 558.4500 1135.8000 558.6000 ;
	    RECT 1105.8000 557.5500 1135.8000 558.4500 ;
	    RECT 1105.8000 557.4000 1107.0000 557.5500 ;
	    RECT 1134.6000 557.4000 1135.8000 557.5500 ;
	    RECT 1137.0000 557.4000 1138.2001 558.6000 ;
	    RECT 1103.1000 556.5000 1104.3000 557.1000 ;
	    RECT 1139.1000 556.5000 1140.0000 561.6000 ;
	    RECT 1141.2001 560.7000 1142.4000 561.0000 ;
	    RECT 1141.2001 559.8000 1142.7001 560.7000 ;
	    RECT 1144.2001 560.4000 1145.4000 561.6000 ;
	    RECT 1168.2001 560.7000 1169.4000 569.7000 ;
	    RECT 1173.6000 561.3000 1174.8000 569.7000 ;
	    RECT 1203.6000 561.3000 1204.8000 569.7000 ;
	    RECT 1173.6000 560.7000 1176.3000 561.3000 ;
	    RECT 1173.9000 560.4000 1176.3000 560.7000 ;
	    RECT 1141.8000 559.5000 1142.7001 559.8000 ;
	    RECT 1144.2001 559.2000 1145.4000 559.5000 ;
	    RECT 1141.8000 557.4000 1143.0000 558.6000 ;
	    RECT 1170.6000 557.4000 1171.8000 558.6000 ;
	    RECT 1172.7001 557.4000 1173.0000 558.6000 ;
	    RECT 1168.2001 556.5000 1169.4000 556.8000 ;
	    RECT 1175.4000 556.5000 1176.3000 560.4000 ;
	    RECT 1202.1000 560.7000 1204.8000 561.3000 ;
	    RECT 1209.0000 560.7000 1210.2001 569.7000 ;
	    RECT 1223.4000 562.5000 1224.6000 569.7000 ;
	    RECT 1225.8000 566.7000 1227.0000 569.7000 ;
	    RECT 1225.8000 565.5000 1227.0000 565.8000 ;
	    RECT 1225.8000 564.4500 1227.0000 564.6000 ;
	    RECT 1245.0000 564.4500 1246.2001 564.6000 ;
	    RECT 1225.8000 563.5500 1246.2001 564.4500 ;
	    RECT 1225.8000 563.4000 1227.0000 563.5500 ;
	    RECT 1245.0000 563.4000 1246.2001 563.5500 ;
	    RECT 1211.4000 561.4500 1212.6000 561.6000 ;
	    RECT 1223.4000 561.4500 1224.6000 561.6000 ;
	    RECT 1240.2001 561.4500 1241.4000 561.6000 ;
	    RECT 1202.1000 560.4000 1204.5000 560.7000 ;
	    RECT 1211.4000 560.5500 1241.4000 561.4500 ;
	    RECT 1251.6000 561.3000 1252.8000 569.7000 ;
	    RECT 1211.4000 560.4000 1212.6000 560.5500 ;
	    RECT 1223.4000 560.4000 1224.6000 560.5500 ;
	    RECT 1240.2001 560.4000 1241.4000 560.5500 ;
	    RECT 1250.1000 560.7000 1252.8000 561.3000 ;
	    RECT 1257.0000 560.7000 1258.2001 569.7000 ;
	    RECT 1281.9000 563.7000 1283.1000 569.7000 ;
	    RECT 1285.8000 563.7000 1287.0000 569.7000 ;
	    RECT 1288.2001 566.7000 1289.4000 569.7000 ;
	    RECT 1287.9000 565.5000 1289.1000 565.8000 ;
	    RECT 1261.8000 561.4500 1263.0000 561.6000 ;
	    RECT 1283.4000 561.4500 1284.6000 561.6000 ;
	    RECT 1250.1000 560.4000 1252.5000 560.7000 ;
	    RECT 1261.8000 560.5500 1284.6000 561.4500 ;
	    RECT 1261.8000 560.4000 1263.0000 560.5500 ;
	    RECT 1283.4000 560.4000 1284.6000 560.5500 ;
	    RECT 1202.1000 556.5000 1203.0000 560.4000 ;
	    RECT 1205.4000 557.4000 1205.7001 558.6000 ;
	    RECT 1206.6000 557.4000 1207.8000 558.6000 ;
	    RECT 1209.0000 556.5000 1210.2001 556.8000 ;
	    RECT 1101.3000 556.2000 1104.3000 556.5000 ;
	    RECT 1105.8000 556.2000 1107.0000 556.5000 ;
	    RECT 1103.4000 555.3000 1104.3000 556.2000 ;
	    RECT 1137.0000 555.3000 1137.9000 556.5000 ;
	    RECT 1139.1000 555.6000 1142.7001 556.5000 ;
	    RECT 1096.2001 554.4000 1102.2001 555.3000 ;
	    RECT 1065.0000 543.3000 1066.2001 549.3000 ;
	    RECT 1096.2001 543.3000 1097.4000 554.4000 ;
	    RECT 1098.6000 543.3000 1099.8000 553.5000 ;
	    RECT 1101.0000 544.2000 1102.2001 554.4000 ;
	    RECT 1103.4000 545.1000 1104.6000 555.3000 ;
	    RECT 1105.8000 544.2000 1107.0000 555.3000 ;
	    RECT 1101.0000 543.3000 1107.0000 544.2000 ;
	    RECT 1137.0000 543.3000 1138.2001 555.3000 ;
	    RECT 1139.4000 543.3000 1140.6000 554.7000 ;
	    RECT 1141.8000 549.3000 1142.7001 555.6000 ;
	    RECT 1168.2001 554.4000 1169.4000 555.6000 ;
	    RECT 1175.4000 555.4500 1176.6000 555.6000 ;
	    RECT 1177.8000 555.4500 1179.0000 555.6000 ;
	    RECT 1175.4000 554.5500 1179.0000 555.4500 ;
	    RECT 1175.4000 554.4000 1176.6000 554.5500 ;
	    RECT 1177.8000 554.4000 1179.0000 554.5500 ;
	    RECT 1201.8000 554.4000 1203.0000 555.6000 ;
	    RECT 1206.6000 555.4500 1207.8000 555.6000 ;
	    RECT 1209.0000 555.4500 1210.2001 555.6000 ;
	    RECT 1211.4000 555.4500 1212.6000 555.6000 ;
	    RECT 1206.6000 554.5500 1212.6000 555.4500 ;
	    RECT 1206.6000 554.4000 1207.8000 554.5500 ;
	    RECT 1209.0000 554.4000 1210.2001 554.5500 ;
	    RECT 1211.4000 554.4000 1212.6000 554.5500 ;
	    RECT 1173.0000 553.5000 1174.2001 553.8000 ;
	    RECT 1204.2001 553.5000 1205.4000 553.8000 ;
	    RECT 1173.0000 551.4000 1174.2001 552.6000 ;
	    RECT 1175.4000 550.5000 1176.3000 553.5000 ;
	    RECT 1170.9000 549.6000 1176.3000 550.5000 ;
	    RECT 1170.9000 549.3000 1171.8000 549.6000 ;
	    RECT 1141.8000 543.3000 1143.0000 549.3000 ;
	    RECT 1144.2001 543.3000 1145.4000 549.3000 ;
	    RECT 1168.2001 543.3000 1169.4000 549.3000 ;
	    RECT 1170.6000 543.3000 1171.8000 549.3000 ;
	    RECT 1175.4000 549.3000 1176.3000 549.6000 ;
	    RECT 1202.1000 550.5000 1203.0000 553.5000 ;
	    RECT 1204.2001 552.4500 1205.4000 552.6000 ;
	    RECT 1213.8000 552.4500 1215.0000 552.6000 ;
	    RECT 1204.2001 551.5500 1215.0000 552.4500 ;
	    RECT 1204.2001 551.4000 1205.4000 551.5500 ;
	    RECT 1213.8000 551.4000 1215.0000 551.5500 ;
	    RECT 1202.1000 549.6000 1207.5000 550.5000 ;
	    RECT 1202.1000 549.3000 1203.0000 549.6000 ;
	    RECT 1173.0000 543.3000 1174.2001 548.7000 ;
	    RECT 1175.4000 543.3000 1176.6000 549.3000 ;
	    RECT 1201.8000 543.3000 1203.0000 549.3000 ;
	    RECT 1206.6000 549.3000 1207.5000 549.6000 ;
	    RECT 1204.2001 543.3000 1205.4000 548.7000 ;
	    RECT 1206.6000 543.3000 1207.8000 549.3000 ;
	    RECT 1209.0000 543.3000 1210.2001 549.3000 ;
	    RECT 1223.4000 543.3000 1224.6000 559.5000 ;
	    RECT 1250.1000 556.5000 1251.0000 560.4000 ;
	    RECT 1283.4000 559.2000 1284.6000 559.5000 ;
	    RECT 1253.4000 557.4000 1253.7001 558.6000 ;
	    RECT 1254.6000 557.4000 1255.8000 558.6000 ;
	    RECT 1281.0000 557.4000 1282.2001 558.6000 ;
	    RECT 1285.8000 558.3000 1286.7001 563.7000 ;
	    RECT 1288.2001 563.4000 1289.4000 564.6000 ;
	    RECT 1314.6000 564.0000 1315.8000 569.7000 ;
	    RECT 1317.0000 564.9000 1318.2001 569.7000 ;
	    RECT 1319.4000 564.0000 1320.6000 569.7000 ;
	    RECT 1314.6000 563.7000 1320.6000 564.0000 ;
	    RECT 1321.8000 563.7000 1323.0000 569.7000 ;
	    RECT 1349.1000 563.7000 1350.3000 569.7000 ;
	    RECT 1353.0000 563.7000 1354.2001 569.7000 ;
	    RECT 1355.4000 566.7000 1356.6000 569.7000 ;
	    RECT 1355.1000 565.5000 1356.3000 565.8000 ;
	    RECT 1355.4000 564.4500 1356.6000 564.6000 ;
	    RECT 1362.6000 564.4500 1363.8000 564.6000 ;
	    RECT 1314.9000 563.1000 1320.3000 563.7000 ;
	    RECT 1321.8000 562.5000 1322.7001 563.7000 ;
	    RECT 1314.6000 560.4000 1315.8000 561.6000 ;
	    RECT 1316.7001 560.7000 1317.0000 562.2000 ;
	    RECT 1319.1000 560.4000 1320.9000 561.6000 ;
	    RECT 1321.8000 561.4500 1323.0000 561.6000 ;
	    RECT 1348.2001 561.4500 1349.4000 561.6000 ;
	    RECT 1321.8000 560.5500 1349.4000 561.4500 ;
	    RECT 1321.8000 560.4000 1323.0000 560.5500 ;
	    RECT 1348.2001 560.4000 1349.4000 560.5500 ;
	    RECT 1350.6000 560.4000 1351.8000 561.6000 ;
	    RECT 1317.0000 559.5000 1318.2001 559.8000 ;
	    RECT 1288.2001 558.4500 1289.4000 558.6000 ;
	    RECT 1317.0000 558.4500 1318.2001 558.6000 ;
	    RECT 1283.1000 556.8000 1283.4000 558.3000 ;
	    RECT 1285.8000 557.4000 1287.3000 558.3000 ;
	    RECT 1288.2001 557.5500 1318.2001 558.4500 ;
	    RECT 1288.2001 557.4000 1289.4000 557.5500 ;
	    RECT 1317.0000 557.4000 1318.2001 557.5500 ;
	    RECT 1257.0000 556.5000 1258.2001 556.8000 ;
	    RECT 1249.8000 554.4000 1251.0000 555.6000 ;
	    RECT 1257.0000 555.4500 1258.2001 555.6000 ;
	    RECT 1259.4000 555.4500 1260.6000 555.6000 ;
	    RECT 1257.0000 554.5500 1260.6000 555.4500 ;
	    RECT 1288.2001 555.3000 1289.1000 556.5000 ;
	    RECT 1319.1000 555.3000 1320.0000 560.4000 ;
	    RECT 1350.6000 559.2000 1351.8000 559.5000 ;
	    RECT 1345.8000 558.4500 1347.0000 558.6000 ;
	    RECT 1348.2001 558.4500 1349.4000 558.6000 ;
	    RECT 1345.8000 557.5500 1349.4000 558.4500 ;
	    RECT 1353.0000 558.3000 1353.9000 563.7000 ;
	    RECT 1355.4000 563.5500 1363.8000 564.4500 ;
	    RECT 1355.4000 563.4000 1356.6000 563.5500 ;
	    RECT 1362.6000 563.4000 1363.8000 563.5500 ;
	    RECT 1389.0000 560.7000 1390.2001 569.7000 ;
	    RECT 1394.4000 561.3000 1395.6000 569.7000 ;
	    RECT 1422.0000 561.3000 1423.2001 569.7000 ;
	    RECT 1394.4000 560.7000 1397.1000 561.3000 ;
	    RECT 1394.7001 560.4000 1397.1000 560.7000 ;
	    RECT 1355.4000 558.4500 1356.6000 558.6000 ;
	    RECT 1386.6000 558.4500 1387.8000 558.6000 ;
	    RECT 1345.8000 557.4000 1347.0000 557.5500 ;
	    RECT 1348.2001 557.4000 1349.4000 557.5500 ;
	    RECT 1350.3000 556.8000 1350.6000 558.3000 ;
	    RECT 1353.0000 557.4000 1354.5000 558.3000 ;
	    RECT 1355.4000 557.5500 1387.8000 558.4500 ;
	    RECT 1355.4000 557.4000 1356.6000 557.5500 ;
	    RECT 1386.6000 557.4000 1387.8000 557.5500 ;
	    RECT 1391.4000 557.4000 1392.6000 558.6000 ;
	    RECT 1393.5000 557.4000 1393.8000 558.6000 ;
	    RECT 1389.0000 556.5000 1390.2001 556.8000 ;
	    RECT 1396.2001 556.5000 1397.1000 560.4000 ;
	    RECT 1420.5000 560.7000 1423.2001 561.3000 ;
	    RECT 1427.4000 560.7000 1428.6000 569.7000 ;
	    RECT 1453.2001 561.3000 1454.4000 569.7000 ;
	    RECT 1451.7001 560.7000 1454.4000 561.3000 ;
	    RECT 1458.6000 560.7000 1459.8000 569.7000 ;
	    RECT 1485.0000 566.7000 1486.2001 569.7000 ;
	    RECT 1485.3000 565.5000 1486.5000 565.8000 ;
	    RECT 1482.6000 564.4500 1483.8000 564.6000 ;
	    RECT 1485.0000 564.4500 1486.2001 564.6000 ;
	    RECT 1482.6000 563.5500 1486.2001 564.4500 ;
	    RECT 1487.4000 563.7000 1488.6000 569.7000 ;
	    RECT 1491.3000 563.7000 1492.5000 569.7000 ;
	    RECT 1511.4000 563.7000 1512.6000 569.7000 ;
	    RECT 1515.3000 564.6000 1516.5000 569.7000 ;
	    RECT 1513.8000 563.7000 1516.5000 564.6000 ;
	    RECT 1540.2001 563.7000 1541.4000 569.7000 ;
	    RECT 1544.1000 564.0000 1545.3000 569.7000 ;
	    RECT 1546.5000 565.2000 1547.7001 569.7000 ;
	    RECT 1546.5000 563.7000 1548.6000 565.2000 ;
	    RECT 1482.6000 563.4000 1483.8000 563.5500 ;
	    RECT 1485.0000 563.4000 1486.2001 563.5500 ;
	    RECT 1420.5000 560.4000 1422.9000 560.7000 ;
	    RECT 1451.7001 560.4000 1454.1000 560.7000 ;
	    RECT 1420.5000 556.5000 1421.4000 560.4000 ;
	    RECT 1423.8000 557.4000 1424.1000 558.6000 ;
	    RECT 1425.0000 557.4000 1426.2001 558.6000 ;
	    RECT 1427.4000 556.5000 1428.6000 556.8000 ;
	    RECT 1451.7001 556.5000 1452.6000 560.4000 ;
	    RECT 1455.0000 557.4000 1455.3000 558.6000 ;
	    RECT 1456.2001 557.4000 1457.4000 558.6000 ;
	    RECT 1485.0000 557.4000 1486.2001 558.6000 ;
	    RECT 1487.7001 558.3000 1488.6000 563.7000 ;
	    RECT 1511.4000 562.5000 1512.6000 562.8000 ;
	    RECT 1489.8000 560.4000 1491.0000 561.6000 ;
	    RECT 1494.6000 561.4500 1495.8000 561.6000 ;
	    RECT 1506.6000 561.4500 1507.8000 561.6000 ;
	    RECT 1511.4000 561.4500 1512.6000 561.6000 ;
	    RECT 1494.6000 560.5500 1512.6000 561.4500 ;
	    RECT 1494.6000 560.4000 1495.8000 560.5500 ;
	    RECT 1506.6000 560.4000 1507.8000 560.5500 ;
	    RECT 1511.4000 560.4000 1512.6000 560.5500 ;
	    RECT 1513.8000 559.5000 1515.0000 563.7000 ;
	    RECT 1540.5000 563.4000 1541.4000 563.7000 ;
	    RECT 1540.5000 562.8000 1543.2001 563.4000 ;
	    RECT 1540.5000 562.5000 1546.8000 562.8000 ;
	    RECT 1542.3000 561.9000 1546.8000 562.5000 ;
	    RECT 1545.6000 561.6000 1546.8000 561.9000 ;
	    RECT 1523.4000 561.4500 1524.6000 561.6000 ;
	    RECT 1540.2001 561.4500 1541.4000 561.6000 ;
	    RECT 1523.4000 560.5500 1541.4000 561.4500 ;
	    RECT 1543.2001 560.7000 1544.4000 561.0000 ;
	    RECT 1523.4000 560.4000 1524.6000 560.5500 ;
	    RECT 1540.2001 560.4000 1541.4000 560.5500 ;
	    RECT 1542.9000 559.8000 1544.4000 560.7000 ;
	    RECT 1542.9000 559.5000 1543.8000 559.8000 ;
	    RECT 1489.8000 559.2000 1491.0000 559.5000 ;
	    RECT 1540.2001 559.2000 1541.4000 559.5000 ;
	    RECT 1487.1000 557.4000 1488.6000 558.3000 ;
	    RECT 1491.0000 556.8000 1491.3000 558.3000 ;
	    RECT 1492.2001 557.4000 1493.4000 558.6000 ;
	    RECT 1513.8000 558.4500 1515.0000 558.6000 ;
	    RECT 1535.4000 558.4500 1536.6000 558.6000 ;
	    RECT 1513.8000 557.5500 1536.6000 558.4500 ;
	    RECT 1513.8000 557.4000 1515.0000 557.5500 ;
	    RECT 1535.4000 557.4000 1536.6000 557.5500 ;
	    RECT 1542.6000 557.4000 1543.8000 558.6000 ;
	    RECT 1458.6000 556.5000 1459.8000 556.8000 ;
	    RECT 1545.6000 556.5000 1546.5000 561.6000 ;
	    RECT 1547.7001 559.5000 1548.6000 563.7000 ;
	    RECT 1547.4000 558.4500 1548.6000 558.6000 ;
	    RECT 1559.4000 558.4500 1560.6000 558.6000 ;
	    RECT 1547.4000 557.5500 1560.6000 558.4500 ;
	    RECT 1547.4000 557.4000 1548.6000 557.5500 ;
	    RECT 1559.4000 557.4000 1560.6000 557.5500 ;
	    RECT 1257.0000 554.4000 1258.2001 554.5500 ;
	    RECT 1259.4000 554.4000 1260.6000 554.5500 ;
	    RECT 1281.0000 554.4000 1287.0000 555.3000 ;
	    RECT 1252.2001 553.5000 1253.4000 553.8000 ;
	    RECT 1250.1000 550.5000 1251.0000 553.5000 ;
	    RECT 1252.2001 551.4000 1253.4000 552.6000 ;
	    RECT 1250.1000 549.6000 1255.5000 550.5000 ;
	    RECT 1250.1000 549.3000 1251.0000 549.6000 ;
	    RECT 1225.8000 543.3000 1227.0000 549.3000 ;
	    RECT 1249.8000 543.3000 1251.0000 549.3000 ;
	    RECT 1254.6000 549.3000 1255.5000 549.6000 ;
	    RECT 1252.2001 543.3000 1253.4000 548.7000 ;
	    RECT 1254.6000 543.3000 1255.8000 549.3000 ;
	    RECT 1257.0000 543.3000 1258.2001 549.3000 ;
	    RECT 1281.0000 543.3000 1282.2001 554.4000 ;
	    RECT 1283.4000 543.3000 1284.6000 553.5000 ;
	    RECT 1285.8000 543.3000 1287.0000 554.4000 ;
	    RECT 1288.2001 543.3000 1289.4000 555.3000 ;
	    RECT 1314.6000 543.3000 1315.8000 555.3000 ;
	    RECT 1318.5000 554.4000 1320.0000 555.3000 ;
	    RECT 1321.8000 555.4500 1323.0000 555.6000 ;
	    RECT 1343.4000 555.4500 1344.6000 555.6000 ;
	    RECT 1321.8000 554.5500 1344.6000 555.4500 ;
	    RECT 1355.4000 555.3000 1356.3000 556.5000 ;
	    RECT 1321.8000 554.4000 1323.0000 554.5500 ;
	    RECT 1343.4000 554.4000 1344.6000 554.5500 ;
	    RECT 1348.2001 554.4000 1354.2001 555.3000 ;
	    RECT 1318.5000 543.3000 1319.7001 554.4000 ;
	    RECT 1320.9000 552.6000 1321.8000 553.5000 ;
	    RECT 1320.6000 551.4000 1321.8000 552.6000 ;
	    RECT 1320.9000 543.3000 1322.1000 549.3000 ;
	    RECT 1348.2001 543.3000 1349.4000 554.4000 ;
	    RECT 1350.6000 543.3000 1351.8000 553.5000 ;
	    RECT 1353.0000 543.3000 1354.2001 554.4000 ;
	    RECT 1355.4000 543.3000 1356.6000 555.3000 ;
	    RECT 1389.0000 554.4000 1390.2001 555.6000 ;
	    RECT 1396.2001 555.4500 1397.4000 555.6000 ;
	    RECT 1417.8000 555.4500 1419.0000 555.6000 ;
	    RECT 1396.2001 554.5500 1419.0000 555.4500 ;
	    RECT 1396.2001 554.4000 1397.4000 554.5500 ;
	    RECT 1417.8000 554.4000 1419.0000 554.5500 ;
	    RECT 1420.2001 554.4000 1421.4000 555.6000 ;
	    RECT 1427.4000 554.4000 1428.6000 555.6000 ;
	    RECT 1446.6000 555.4500 1447.8000 555.6000 ;
	    RECT 1451.4000 555.4500 1452.6000 555.6000 ;
	    RECT 1446.6000 554.5500 1452.6000 555.4500 ;
	    RECT 1446.6000 554.4000 1447.8000 554.5500 ;
	    RECT 1451.4000 554.4000 1452.6000 554.5500 ;
	    RECT 1458.6000 555.4500 1459.8000 555.6000 ;
	    RECT 1475.4000 555.4500 1476.6000 555.6000 ;
	    RECT 1458.6000 554.5500 1476.6000 555.4500 ;
	    RECT 1485.3000 555.3000 1486.2001 556.5000 ;
	    RECT 1458.6000 554.4000 1459.8000 554.5500 ;
	    RECT 1475.4000 554.4000 1476.6000 554.5500 ;
	    RECT 1393.8000 553.5000 1395.0000 553.8000 ;
	    RECT 1422.6000 553.5000 1423.8000 553.8000 ;
	    RECT 1453.8000 553.5000 1455.0000 553.8000 ;
	    RECT 1386.6000 552.4500 1387.8000 552.6000 ;
	    RECT 1393.8000 552.4500 1395.0000 552.6000 ;
	    RECT 1386.6000 551.5500 1395.0000 552.4500 ;
	    RECT 1386.6000 551.4000 1387.8000 551.5500 ;
	    RECT 1393.8000 551.4000 1395.0000 551.5500 ;
	    RECT 1396.2001 550.5000 1397.1000 553.5000 ;
	    RECT 1391.7001 549.6000 1397.1000 550.5000 ;
	    RECT 1391.7001 549.3000 1392.6000 549.6000 ;
	    RECT 1362.6000 546.4500 1363.8000 546.6000 ;
	    RECT 1369.8000 546.4500 1371.0000 546.6000 ;
	    RECT 1362.6000 545.5500 1371.0000 546.4500 ;
	    RECT 1362.6000 545.4000 1363.8000 545.5500 ;
	    RECT 1369.8000 545.4000 1371.0000 545.5500 ;
	    RECT 1389.0000 543.3000 1390.2001 549.3000 ;
	    RECT 1391.4000 543.3000 1392.6000 549.3000 ;
	    RECT 1396.2001 549.3000 1397.1000 549.6000 ;
	    RECT 1420.5000 550.5000 1421.4000 553.5000 ;
	    RECT 1422.6000 551.4000 1423.8000 552.6000 ;
	    RECT 1451.7001 550.5000 1452.6000 553.5000 ;
	    RECT 1453.8000 551.4000 1455.0000 552.6000 ;
	    RECT 1420.5000 549.6000 1425.9000 550.5000 ;
	    RECT 1420.5000 549.3000 1421.4000 549.6000 ;
	    RECT 1393.8000 543.3000 1395.0000 548.7000 ;
	    RECT 1396.2001 543.3000 1397.4000 549.3000 ;
	    RECT 1420.2001 543.3000 1421.4000 549.3000 ;
	    RECT 1425.0000 549.3000 1425.9000 549.6000 ;
	    RECT 1451.7001 549.6000 1457.1000 550.5000 ;
	    RECT 1451.7001 549.3000 1452.6000 549.6000 ;
	    RECT 1422.6000 543.3000 1423.8000 548.7000 ;
	    RECT 1425.0000 543.3000 1426.2001 549.3000 ;
	    RECT 1427.4000 543.3000 1428.6000 549.3000 ;
	    RECT 1451.4000 543.3000 1452.6000 549.3000 ;
	    RECT 1456.2001 549.3000 1457.1000 549.6000 ;
	    RECT 1453.8000 543.3000 1455.0000 548.7000 ;
	    RECT 1456.2001 543.3000 1457.4000 549.3000 ;
	    RECT 1458.6000 543.3000 1459.8000 549.3000 ;
	    RECT 1463.4000 546.4500 1464.6000 546.6000 ;
	    RECT 1473.0000 546.4500 1474.2001 546.6000 ;
	    RECT 1463.4000 545.5500 1474.2001 546.4500 ;
	    RECT 1463.4000 545.4000 1464.6000 545.5500 ;
	    RECT 1473.0000 545.4000 1474.2001 545.5500 ;
	    RECT 1485.0000 543.3000 1486.2001 555.3000 ;
	    RECT 1487.4000 554.4000 1493.4000 555.3000 ;
	    RECT 1487.4000 543.3000 1488.6000 554.4000 ;
	    RECT 1489.8000 543.3000 1491.0000 553.5000 ;
	    RECT 1492.2001 543.3000 1493.4000 554.4000 ;
	    RECT 1511.4000 543.3000 1512.6000 549.3000 ;
	    RECT 1513.8000 543.3000 1515.0000 556.5000 ;
	    RECT 1542.9000 555.6000 1546.5000 556.5000 ;
	    RECT 1516.2001 554.4000 1517.4000 555.6000 ;
	    RECT 1516.2001 553.2000 1517.4000 553.5000 ;
	    RECT 1542.9000 549.3000 1543.8000 555.6000 ;
	    RECT 1547.7001 555.3000 1548.6000 556.5000 ;
	    RECT 1516.2001 543.3000 1517.4000 549.3000 ;
	    RECT 1540.2001 543.3000 1541.4000 549.3000 ;
	    RECT 1542.6000 543.3000 1543.8000 549.3000 ;
	    RECT 1545.0000 543.3000 1546.2001 554.7000 ;
	    RECT 1547.4000 543.3000 1548.6000 555.3000 ;
	    RECT 1.2000 540.6000 1569.0000 542.4000 ;
	    RECT 124.2000 533.7000 125.4000 539.7000 ;
	    RECT 126.6000 534.6000 127.8000 539.7000 ;
	    RECT 126.3000 533.7000 127.8000 534.6000 ;
	    RECT 129.0000 533.7000 130.2000 540.6000 ;
	    RECT 126.3000 532.8000 127.2000 533.7000 ;
	    RECT 131.4000 532.8000 132.6000 539.7000 ;
	    RECT 133.8000 533.7000 135.0000 539.7000 ;
	    RECT 136.2000 535.5000 137.4000 539.7000 ;
	    RECT 138.6000 535.5000 139.8000 539.7000 ;
	    RECT 124.2000 531.9000 127.2000 532.8000 ;
	    RECT 124.2000 523.5000 125.4000 531.9000 ;
	    RECT 128.1000 531.6000 134.4000 532.8000 ;
	    RECT 141.0000 532.5000 142.2000 539.7000 ;
	    RECT 143.4000 533.7000 144.6000 539.7000 ;
	    RECT 145.8000 532.5000 147.0000 539.7000 ;
	    RECT 148.2000 533.7000 149.4000 539.7000 ;
	    RECT 128.1000 531.0000 129.0000 531.6000 ;
	    RECT 126.6000 529.8000 129.0000 531.0000 ;
	    RECT 133.5000 530.7000 142.2000 531.6000 ;
	    RECT 130.5000 529.8000 132.6000 530.7000 ;
	    RECT 130.5000 529.5000 139.8000 529.8000 ;
	    RECT 131.7000 528.9000 139.8000 529.5000 ;
	    RECT 138.6000 528.6000 139.8000 528.9000 ;
	    RECT 141.3000 529.5000 142.2000 530.7000 ;
	    RECT 143.1000 530.4000 147.0000 531.6000 ;
	    RECT 150.6000 530.4000 151.8000 539.7000 ;
	    RECT 153.0000 535.5000 154.2000 539.7000 ;
	    RECT 155.4000 535.5000 156.6000 539.7000 ;
	    RECT 157.8000 535.5000 159.0000 539.7000 ;
	    RECT 160.2000 533.7000 161.4000 539.7000 ;
	    RECT 155.4000 531.6000 161.7000 532.8000 ;
	    RECT 162.6000 531.6000 163.8000 539.7000 ;
	    RECT 165.0000 533.7000 166.2000 539.7000 ;
	    RECT 167.4000 532.8000 168.6000 539.7000 ;
	    RECT 169.8000 533.7000 171.0000 539.7000 ;
	    RECT 167.4000 531.9000 171.3000 532.8000 ;
	    RECT 172.2000 532.5000 173.4000 539.7000 ;
	    RECT 174.6000 533.7000 175.8000 539.7000 ;
	    RECT 193.8000 533.7000 195.0000 539.7000 ;
	    RECT 162.6000 530.4000 166.5000 531.6000 ;
	    RECT 153.0000 529.5000 154.2000 529.8000 ;
	    RECT 141.3000 528.6000 154.2000 529.5000 ;
	    RECT 157.8000 529.5000 159.0000 529.8000 ;
	    RECT 170.4000 529.5000 171.3000 531.9000 ;
	    RECT 172.2000 531.4500 173.4000 531.6000 ;
	    RECT 191.4000 531.4500 192.6000 531.6000 ;
	    RECT 172.2000 530.5500 192.6000 531.4500 ;
	    RECT 172.2000 530.4000 173.4000 530.5500 ;
	    RECT 191.4000 530.4000 192.6000 530.5500 ;
	    RECT 193.8000 529.5000 195.0000 529.8000 ;
	    RECT 157.8000 528.6000 171.3000 529.5000 ;
	    RECT 129.0000 527.4000 130.2000 528.6000 ;
	    RECT 134.1000 527.7000 135.3000 528.0000 ;
	    RECT 131.1000 526.8000 169.5000 527.7000 ;
	    RECT 168.3000 526.5000 169.5000 526.8000 ;
	    RECT 170.4000 525.9000 171.3000 528.6000 ;
	    RECT 172.2000 528.0000 173.4000 529.5000 ;
	    RECT 172.2000 526.8000 173.7000 528.0000 ;
	    RECT 193.8000 527.4000 195.0000 528.6000 ;
	    RECT 126.3000 525.0000 132.9000 525.9000 ;
	    RECT 126.3000 524.7000 127.5000 525.0000 ;
	    RECT 133.8000 524.4000 135.0000 525.6000 ;
	    RECT 135.9000 525.0000 161.4000 525.9000 ;
	    RECT 170.4000 525.0000 171.6000 525.9000 ;
	    RECT 160.2000 524.1000 161.4000 525.0000 ;
	    RECT 124.2000 522.3000 137.4000 523.5000 ;
	    RECT 138.3000 522.9000 141.3000 524.1000 ;
	    RECT 147.0000 522.9000 151.8000 524.1000 ;
	    RECT 124.2000 513.3000 125.4000 522.3000 ;
	    RECT 127.8000 520.2000 132.3000 521.4000 ;
	    RECT 131.1000 519.3000 132.3000 520.2000 ;
	    RECT 140.1000 519.3000 141.3000 522.9000 ;
	    RECT 143.4000 521.4000 144.6000 522.6000 ;
	    RECT 151.2000 521.7000 152.4000 522.0000 ;
	    RECT 145.8000 520.8000 152.4000 521.7000 ;
	    RECT 145.8000 520.5000 147.0000 520.8000 ;
	    RECT 143.4000 520.2000 144.6000 520.5000 ;
	    RECT 155.4000 519.6000 156.6000 523.8000 ;
	    RECT 164.1000 522.9000 169.8000 524.1000 ;
	    RECT 164.1000 521.1000 165.3000 522.9000 ;
	    RECT 170.7000 522.0000 171.6000 525.0000 ;
	    RECT 145.8000 519.3000 147.0000 519.6000 ;
	    RECT 129.0000 513.3000 130.2000 519.3000 ;
	    RECT 131.1000 518.1000 135.0000 519.3000 ;
	    RECT 140.1000 518.4000 147.0000 519.3000 ;
	    RECT 148.2000 518.4000 149.4000 519.6000 ;
	    RECT 150.3000 518.4000 150.6000 519.6000 ;
	    RECT 155.1000 518.4000 156.6000 519.6000 ;
	    RECT 162.6000 520.2000 165.3000 521.1000 ;
	    RECT 169.8000 521.1000 171.6000 522.0000 ;
	    RECT 162.6000 519.3000 163.8000 520.2000 ;
	    RECT 133.8000 513.3000 135.0000 518.1000 ;
	    RECT 160.2000 518.1000 163.8000 519.3000 ;
	    RECT 136.2000 513.3000 137.4000 517.5000 ;
	    RECT 138.6000 513.3000 139.8000 517.5000 ;
	    RECT 141.0000 513.3000 142.2000 517.5000 ;
	    RECT 143.4000 513.3000 144.6000 516.3000 ;
	    RECT 145.8000 513.3000 147.0000 517.5000 ;
	    RECT 148.2000 513.3000 149.4000 516.3000 ;
	    RECT 150.6000 513.3000 151.8000 517.5000 ;
	    RECT 153.0000 513.3000 154.2000 517.5000 ;
	    RECT 155.4000 513.3000 156.6000 517.5000 ;
	    RECT 157.8000 513.3000 159.0000 517.5000 ;
	    RECT 160.2000 513.3000 161.4000 518.1000 ;
	    RECT 165.0000 513.3000 166.2000 519.3000 ;
	    RECT 169.8000 513.3000 171.0000 521.1000 ;
	    RECT 172.5000 520.2000 173.7000 526.8000 ;
	    RECT 196.2000 526.5000 197.4000 539.7000 ;
	    RECT 198.6000 533.7000 199.8000 539.7000 ;
	    RECT 330.6000 533.7000 331.8000 539.7000 ;
	    RECT 333.0000 534.6000 334.2000 539.7000 ;
	    RECT 332.7000 533.7000 334.2000 534.6000 ;
	    RECT 335.4000 533.7000 336.6000 540.6000 ;
	    RECT 332.7000 532.8000 333.6000 533.7000 ;
	    RECT 337.8000 532.8000 339.0000 539.7000 ;
	    RECT 340.2000 533.7000 341.4000 539.7000 ;
	    RECT 342.6000 535.5000 343.8000 539.7000 ;
	    RECT 345.0000 535.5000 346.2000 539.7000 ;
	    RECT 330.6000 531.9000 333.6000 532.8000 ;
	    RECT 196.2000 525.4500 197.4000 525.6000 ;
	    RECT 246.6000 525.4500 247.8000 525.6000 ;
	    RECT 196.2000 524.5500 247.8000 525.4500 ;
	    RECT 196.2000 524.4000 197.4000 524.5500 ;
	    RECT 246.6000 524.4000 247.8000 524.5500 ;
	    RECT 301.8000 525.4500 303.0000 525.6000 ;
	    RECT 306.6000 525.4500 307.8000 525.6000 ;
	    RECT 301.8000 524.5500 307.8000 525.4500 ;
	    RECT 301.8000 524.4000 303.0000 524.5500 ;
	    RECT 306.6000 524.4000 307.8000 524.5500 ;
	    RECT 330.6000 523.5000 331.8000 531.9000 ;
	    RECT 334.5000 531.6000 340.8000 532.8000 ;
	    RECT 347.4000 532.5000 348.6000 539.7000 ;
	    RECT 349.8000 533.7000 351.0000 539.7000 ;
	    RECT 352.2000 532.5000 353.4000 539.7000 ;
	    RECT 354.6000 533.7000 355.8000 539.7000 ;
	    RECT 334.5000 531.0000 335.4000 531.6000 ;
	    RECT 333.0000 529.8000 335.4000 531.0000 ;
	    RECT 339.9000 530.7000 348.6000 531.6000 ;
	    RECT 336.9000 529.8000 339.0000 530.7000 ;
	    RECT 336.9000 529.5000 346.2000 529.8000 ;
	    RECT 338.1000 528.9000 346.2000 529.5000 ;
	    RECT 345.0000 528.6000 346.2000 528.9000 ;
	    RECT 347.7000 529.5000 348.6000 530.7000 ;
	    RECT 349.5000 530.4000 353.4000 531.6000 ;
	    RECT 357.0000 530.4000 358.2000 539.7000 ;
	    RECT 359.4000 535.5000 360.6000 539.7000 ;
	    RECT 361.8000 535.5000 363.0000 539.7000 ;
	    RECT 364.2000 535.5000 365.4000 539.7000 ;
	    RECT 366.6000 533.7000 367.8000 539.7000 ;
	    RECT 361.8000 531.6000 368.1000 532.8000 ;
	    RECT 369.0000 531.6000 370.2000 539.7000 ;
	    RECT 371.4000 533.7000 372.6000 539.7000 ;
	    RECT 373.8000 532.8000 375.0000 539.7000 ;
	    RECT 376.2000 533.7000 377.4000 539.7000 ;
	    RECT 373.8000 531.9000 377.7000 532.8000 ;
	    RECT 378.6000 532.5000 379.8000 539.7000 ;
	    RECT 381.0000 533.7000 382.2000 539.7000 ;
	    RECT 513.0000 533.7000 514.2000 539.7000 ;
	    RECT 515.4000 534.6000 516.6000 539.7000 ;
	    RECT 515.1000 533.7000 516.6000 534.6000 ;
	    RECT 517.8000 533.7000 519.0000 540.6000 ;
	    RECT 515.1000 532.8000 516.0000 533.7000 ;
	    RECT 520.2000 532.8000 521.4000 539.7000 ;
	    RECT 522.6000 533.7000 523.8000 539.7000 ;
	    RECT 525.0000 535.5000 526.2000 539.7000 ;
	    RECT 527.4000 535.5000 528.6000 539.7000 ;
	    RECT 369.0000 530.4000 372.9000 531.6000 ;
	    RECT 359.4000 529.5000 360.6000 529.8000 ;
	    RECT 347.7000 528.6000 360.6000 529.5000 ;
	    RECT 364.2000 529.5000 365.4000 529.8000 ;
	    RECT 376.8000 529.5000 377.7000 531.9000 ;
	    RECT 513.0000 531.9000 516.0000 532.8000 ;
	    RECT 378.6000 530.4000 379.8000 531.6000 ;
	    RECT 364.2000 528.6000 377.7000 529.5000 ;
	    RECT 335.4000 527.4000 336.6000 528.6000 ;
	    RECT 340.5000 527.7000 341.7000 528.0000 ;
	    RECT 337.5000 526.8000 375.9000 527.7000 ;
	    RECT 374.7000 526.5000 375.9000 526.8000 ;
	    RECT 376.8000 525.9000 377.7000 528.6000 ;
	    RECT 378.6000 528.0000 379.8000 529.5000 ;
	    RECT 378.6000 526.8000 380.1000 528.0000 ;
	    RECT 332.7000 525.0000 339.3000 525.9000 ;
	    RECT 332.7000 524.7000 333.9000 525.0000 ;
	    RECT 340.2000 524.4000 341.4000 525.6000 ;
	    RECT 342.3000 525.0000 367.8000 525.9000 ;
	    RECT 376.8000 525.0000 378.0000 525.9000 ;
	    RECT 366.6000 524.1000 367.8000 525.0000 ;
	    RECT 172.2000 519.0000 173.7000 520.2000 ;
	    RECT 196.2000 519.3000 197.4000 523.5000 ;
	    RECT 198.6000 522.4500 199.8000 522.6000 ;
	    RECT 328.2000 522.4500 329.4000 522.6000 ;
	    RECT 198.6000 521.5500 329.4000 522.4500 ;
	    RECT 198.6000 521.4000 199.8000 521.5500 ;
	    RECT 328.2000 521.4000 329.4000 521.5500 ;
	    RECT 330.6000 522.3000 343.8000 523.5000 ;
	    RECT 344.7000 522.9000 347.7000 524.1000 ;
	    RECT 353.4000 522.9000 358.2000 524.1000 ;
	    RECT 198.6000 520.2000 199.8000 520.5000 ;
	    RECT 172.2000 513.3000 173.4000 519.0000 ;
	    RECT 194.7000 518.4000 197.4000 519.3000 ;
	    RECT 174.6000 513.3000 175.8000 516.3000 ;
	    RECT 194.7000 513.3000 195.9000 518.4000 ;
	    RECT 198.6000 513.3000 199.8000 519.3000 ;
	    RECT 330.6000 513.3000 331.8000 522.3000 ;
	    RECT 334.2000 520.2000 338.7000 521.4000 ;
	    RECT 337.5000 519.3000 338.7000 520.2000 ;
	    RECT 346.5000 519.3000 347.7000 522.9000 ;
	    RECT 349.8000 521.4000 351.0000 522.6000 ;
	    RECT 357.6000 521.7000 358.8000 522.0000 ;
	    RECT 352.2000 520.8000 358.8000 521.7000 ;
	    RECT 352.2000 520.5000 353.4000 520.8000 ;
	    RECT 349.8000 520.2000 351.0000 520.5000 ;
	    RECT 361.8000 519.6000 363.0000 523.8000 ;
	    RECT 370.5000 522.9000 376.2000 524.1000 ;
	    RECT 370.5000 521.1000 371.7000 522.9000 ;
	    RECT 377.1000 522.0000 378.0000 525.0000 ;
	    RECT 352.2000 519.3000 353.4000 519.6000 ;
	    RECT 335.4000 513.3000 336.6000 519.3000 ;
	    RECT 337.5000 518.1000 341.4000 519.3000 ;
	    RECT 346.5000 518.4000 353.4000 519.3000 ;
	    RECT 354.6000 518.4000 355.8000 519.6000 ;
	    RECT 356.7000 518.4000 357.0000 519.6000 ;
	    RECT 361.5000 518.4000 363.0000 519.6000 ;
	    RECT 369.0000 520.2000 371.7000 521.1000 ;
	    RECT 376.2000 521.1000 378.0000 522.0000 ;
	    RECT 369.0000 519.3000 370.2000 520.2000 ;
	    RECT 340.2000 513.3000 341.4000 518.1000 ;
	    RECT 366.6000 518.1000 370.2000 519.3000 ;
	    RECT 342.6000 513.3000 343.8000 517.5000 ;
	    RECT 345.0000 513.3000 346.2000 517.5000 ;
	    RECT 347.4000 513.3000 348.6000 517.5000 ;
	    RECT 349.8000 513.3000 351.0000 516.3000 ;
	    RECT 352.2000 513.3000 353.4000 517.5000 ;
	    RECT 354.6000 513.3000 355.8000 516.3000 ;
	    RECT 357.0000 513.3000 358.2000 517.5000 ;
	    RECT 359.4000 513.3000 360.6000 517.5000 ;
	    RECT 361.8000 513.3000 363.0000 517.5000 ;
	    RECT 364.2000 513.3000 365.4000 517.5000 ;
	    RECT 366.6000 513.3000 367.8000 518.1000 ;
	    RECT 371.4000 513.3000 372.6000 519.3000 ;
	    RECT 376.2000 513.3000 377.4000 521.1000 ;
	    RECT 378.9000 520.2000 380.1000 526.8000 ;
	    RECT 378.6000 519.0000 380.1000 520.2000 ;
	    RECT 513.0000 523.5000 514.2000 531.9000 ;
	    RECT 516.9000 531.6000 523.2000 532.8000 ;
	    RECT 529.8000 532.5000 531.0000 539.7000 ;
	    RECT 532.2000 533.7000 533.4000 539.7000 ;
	    RECT 534.6000 532.5000 535.8000 539.7000 ;
	    RECT 537.0000 533.7000 538.2000 539.7000 ;
	    RECT 516.9000 531.0000 517.8000 531.6000 ;
	    RECT 515.4000 529.8000 517.8000 531.0000 ;
	    RECT 522.3000 530.7000 531.0000 531.6000 ;
	    RECT 519.3000 529.8000 521.4000 530.7000 ;
	    RECT 519.3000 529.5000 528.6000 529.8000 ;
	    RECT 520.5000 528.9000 528.6000 529.5000 ;
	    RECT 527.4000 528.6000 528.6000 528.9000 ;
	    RECT 530.1000 529.5000 531.0000 530.7000 ;
	    RECT 531.9000 530.4000 535.8000 531.6000 ;
	    RECT 539.4000 530.4000 540.6000 539.7000 ;
	    RECT 541.8000 535.5000 543.0000 539.7000 ;
	    RECT 544.2000 535.5000 545.4000 539.7000 ;
	    RECT 546.6000 535.5000 547.8000 539.7000 ;
	    RECT 549.0000 533.7000 550.2000 539.7000 ;
	    RECT 544.2000 531.6000 550.5000 532.8000 ;
	    RECT 551.4000 531.6000 552.6000 539.7000 ;
	    RECT 553.8000 533.7000 555.0000 539.7000 ;
	    RECT 556.2000 532.8000 557.4000 539.7000 ;
	    RECT 558.6000 533.7000 559.8000 539.7000 ;
	    RECT 556.2000 531.9000 560.1000 532.8000 ;
	    RECT 561.0000 532.5000 562.2000 539.7000 ;
	    RECT 563.4000 533.7000 564.6000 539.7000 ;
	    RECT 551.4000 530.4000 555.3000 531.6000 ;
	    RECT 541.8000 529.5000 543.0000 529.8000 ;
	    RECT 530.1000 528.6000 543.0000 529.5000 ;
	    RECT 546.6000 529.5000 547.8000 529.8000 ;
	    RECT 559.2000 529.5000 560.1000 531.9000 ;
	    RECT 561.0000 531.4500 562.2000 531.6000 ;
	    RECT 563.4000 531.4500 564.6000 531.6000 ;
	    RECT 561.0000 530.5500 564.6000 531.4500 ;
	    RECT 561.0000 530.4000 562.2000 530.5500 ;
	    RECT 563.4000 530.4000 564.6000 530.5500 ;
	    RECT 546.6000 528.6000 560.1000 529.5000 ;
	    RECT 517.8000 527.4000 519.0000 528.6000 ;
	    RECT 522.9000 527.7000 524.1000 528.0000 ;
	    RECT 519.9000 526.8000 558.3000 527.7000 ;
	    RECT 557.1000 526.5000 558.3000 526.8000 ;
	    RECT 559.2000 525.9000 560.1000 528.6000 ;
	    RECT 561.0000 528.0000 562.2000 529.5000 ;
	    RECT 561.0000 526.8000 562.5000 528.0000 ;
	    RECT 515.1000 525.0000 521.7000 525.9000 ;
	    RECT 515.1000 524.7000 516.3000 525.0000 ;
	    RECT 522.6000 524.4000 523.8000 525.6000 ;
	    RECT 524.7000 525.0000 550.2000 525.9000 ;
	    RECT 559.2000 525.0000 560.4000 525.9000 ;
	    RECT 549.0000 524.1000 550.2000 525.0000 ;
	    RECT 513.0000 522.3000 526.2000 523.5000 ;
	    RECT 527.1000 522.9000 530.1000 524.1000 ;
	    RECT 535.8000 522.9000 540.6000 524.1000 ;
	    RECT 378.6000 513.3000 379.8000 519.0000 ;
	    RECT 381.0000 513.3000 382.2000 516.3000 ;
	    RECT 513.0000 513.3000 514.2000 522.3000 ;
	    RECT 516.6000 520.2000 521.1000 521.4000 ;
	    RECT 519.9000 519.3000 521.1000 520.2000 ;
	    RECT 528.9000 519.3000 530.1000 522.9000 ;
	    RECT 532.2000 521.4000 533.4000 522.6000 ;
	    RECT 540.0000 521.7000 541.2000 522.0000 ;
	    RECT 534.6000 520.8000 541.2000 521.7000 ;
	    RECT 534.6000 520.5000 535.8000 520.8000 ;
	    RECT 532.2000 520.2000 533.4000 520.5000 ;
	    RECT 544.2000 519.6000 545.4000 523.8000 ;
	    RECT 552.9000 522.9000 558.6000 524.1000 ;
	    RECT 552.9000 521.1000 554.1000 522.9000 ;
	    RECT 559.5000 522.0000 560.4000 525.0000 ;
	    RECT 534.6000 519.3000 535.8000 519.6000 ;
	    RECT 517.8000 513.3000 519.0000 519.3000 ;
	    RECT 519.9000 518.1000 523.8000 519.3000 ;
	    RECT 528.9000 518.4000 535.8000 519.3000 ;
	    RECT 537.0000 518.4000 538.2000 519.6000 ;
	    RECT 539.1000 518.4000 539.4000 519.6000 ;
	    RECT 543.9000 518.4000 545.4000 519.6000 ;
	    RECT 551.4000 520.2000 554.1000 521.1000 ;
	    RECT 558.6000 521.1000 560.4000 522.0000 ;
	    RECT 551.4000 519.3000 552.6000 520.2000 ;
	    RECT 522.6000 513.3000 523.8000 518.1000 ;
	    RECT 549.0000 518.1000 552.6000 519.3000 ;
	    RECT 525.0000 513.3000 526.2000 517.5000 ;
	    RECT 527.4000 513.3000 528.6000 517.5000 ;
	    RECT 529.8000 513.3000 531.0000 517.5000 ;
	    RECT 532.2000 513.3000 533.4000 516.3000 ;
	    RECT 534.6000 513.3000 535.8000 517.5000 ;
	    RECT 537.0000 513.3000 538.2000 516.3000 ;
	    RECT 539.4000 513.3000 540.6000 517.5000 ;
	    RECT 541.8000 513.3000 543.0000 517.5000 ;
	    RECT 544.2000 513.3000 545.4000 517.5000 ;
	    RECT 546.6000 513.3000 547.8000 517.5000 ;
	    RECT 549.0000 513.3000 550.2000 518.1000 ;
	    RECT 553.8000 513.3000 555.0000 519.3000 ;
	    RECT 558.6000 513.3000 559.8000 521.1000 ;
	    RECT 561.3000 520.2000 562.5000 526.8000 ;
	    RECT 575.4000 523.5000 576.6000 539.7000 ;
	    RECT 577.8000 533.7000 579.0000 539.7000 ;
	    RECT 630.6000 527.7000 631.8000 539.7000 ;
	    RECT 633.0000 526.8000 634.2000 539.7000 ;
	    RECT 635.4000 527.7000 636.6000 539.7000 ;
	    RECT 637.8000 526.8000 639.0000 539.7000 ;
	    RECT 640.2000 527.7000 641.4000 539.7000 ;
	    RECT 642.6000 526.8000 643.8000 539.7000 ;
	    RECT 645.0000 527.7000 646.2000 539.7000 ;
	    RECT 647.4000 526.8000 648.6000 539.7000 ;
	    RECT 649.8000 527.7000 651.0000 539.7000 ;
	    RECT 671.4000 533.7000 672.6000 539.7000 ;
	    RECT 633.0000 525.6000 635.7000 526.8000 ;
	    RECT 637.8000 525.6000 641.1000 526.8000 ;
	    RECT 642.6000 525.6000 645.9000 526.8000 ;
	    RECT 647.4000 526.5000 651.0000 526.8000 ;
	    RECT 647.4000 525.6000 648.9000 526.5000 ;
	    RECT 634.5000 523.5000 635.7000 525.6000 ;
	    RECT 639.9000 523.5000 641.1000 525.6000 ;
	    RECT 644.7000 523.5000 645.9000 525.6000 ;
	    RECT 649.8000 524.4000 651.0000 525.6000 ;
	    RECT 673.8000 523.5000 675.0000 539.7000 ;
	    RECT 695.4000 539.4000 696.6000 540.6000 ;
	    RECT 697.8000 527.7000 699.0000 539.7000 ;
	    RECT 701.7000 528.6000 702.9000 539.7000 ;
	    RECT 704.1000 533.7000 705.3000 539.7000 ;
	    RECT 724.2000 533.7000 725.4000 539.7000 ;
	    RECT 703.8000 530.4000 705.0000 531.6000 ;
	    RECT 704.1000 529.5000 705.0000 530.4000 ;
	    RECT 701.7000 527.7000 703.2000 528.6000 ;
	    RECT 700.2000 525.4500 701.4000 525.6000 ;
	    RECT 693.1500 524.5500 701.4000 525.4500 ;
	    RECT 575.4000 521.4000 576.6000 522.6000 ;
	    RECT 632.7000 522.3000 633.3000 523.5000 ;
	    RECT 634.5000 522.3000 638.4000 523.5000 ;
	    RECT 639.9000 522.3000 643.5000 523.5000 ;
	    RECT 644.7000 522.3000 648.6000 523.5000 ;
	    RECT 634.5000 521.4000 635.7000 522.3000 ;
	    RECT 639.9000 521.4000 641.1000 522.3000 ;
	    RECT 644.7000 521.4000 645.9000 522.3000 ;
	    RECT 649.8000 521.4000 651.0000 523.5000 ;
	    RECT 673.8000 522.4500 675.0000 522.6000 ;
	    RECT 693.1500 522.4500 694.0500 524.5500 ;
	    RECT 700.2000 524.4000 701.4000 524.5500 ;
	    RECT 700.2000 523.2000 701.4000 523.5000 ;
	    RECT 702.3000 522.6000 703.2000 527.7000 ;
	    RECT 705.0000 527.4000 706.2000 528.6000 ;
	    RECT 705.1500 525.4500 706.0500 527.4000 ;
	    RECT 726.6000 526.5000 727.8000 539.7000 ;
	    RECT 729.0000 533.7000 730.2000 539.7000 ;
	    RECT 743.4000 533.7000 744.6000 539.7000 ;
	    RECT 729.0000 529.5000 730.2000 529.8000 ;
	    RECT 729.0000 528.4500 730.2000 528.6000 ;
	    RECT 743.4000 528.4500 744.6000 528.6000 ;
	    RECT 729.0000 527.5500 744.6000 528.4500 ;
	    RECT 729.0000 527.4000 730.2000 527.5500 ;
	    RECT 743.4000 527.4000 744.6000 527.5500 ;
	    RECT 726.6000 525.4500 727.8000 525.6000 ;
	    RECT 705.1500 524.5500 727.8000 525.4500 ;
	    RECT 726.6000 524.4000 727.8000 524.5500 ;
	    RECT 745.8000 523.5000 747.0000 539.7000 ;
	    RECT 760.2000 533.7000 761.4000 539.7000 ;
	    RECT 762.6000 523.5000 763.8000 539.7000 ;
	    RECT 781.8000 533.7000 783.0000 539.7000 ;
	    RECT 784.2000 526.5000 785.4000 539.7000 ;
	    RECT 786.6000 533.7000 787.8000 539.7000 ;
	    RECT 805.8000 533.7000 807.0000 539.7000 ;
	    RECT 786.6000 529.5000 787.8000 529.8000 ;
	    RECT 805.8000 529.5000 807.0000 529.8000 ;
	    RECT 786.6000 527.4000 787.8000 528.6000 ;
	    RECT 805.8000 527.4000 807.0000 528.6000 ;
	    RECT 784.2000 525.4500 785.4000 525.6000 ;
	    RECT 805.9500 525.4500 806.8500 527.4000 ;
	    RECT 808.2000 526.5000 809.4000 539.7000 ;
	    RECT 810.6000 533.7000 811.8000 539.7000 ;
	    RECT 837.0000 533.7000 838.2000 539.7000 ;
	    RECT 839.4000 533.7000 840.6000 539.7000 ;
	    RECT 841.8000 534.3000 843.0000 539.7000 ;
	    RECT 839.7000 533.4000 840.6000 533.7000 ;
	    RECT 844.2000 533.7000 845.4000 539.7000 ;
	    RECT 858.6000 533.7000 859.8000 539.7000 ;
	    RECT 844.2000 533.4000 845.1000 533.7000 ;
	    RECT 839.7000 532.5000 845.1000 533.4000 ;
	    RECT 810.6000 531.4500 811.8000 531.6000 ;
	    RECT 841.8000 531.4500 843.0000 531.6000 ;
	    RECT 810.6000 530.5500 843.0000 531.4500 ;
	    RECT 810.6000 530.4000 811.8000 530.5500 ;
	    RECT 841.8000 530.4000 843.0000 530.5500 ;
	    RECT 844.2000 529.5000 845.1000 532.5000 ;
	    RECT 841.8000 529.2000 843.0000 529.5000 ;
	    RECT 817.8000 528.4500 819.0000 528.6000 ;
	    RECT 837.0000 528.4500 838.2000 528.6000 ;
	    RECT 817.8000 527.5500 838.2000 528.4500 ;
	    RECT 817.8000 527.4000 819.0000 527.5500 ;
	    RECT 837.0000 527.4000 838.2000 527.5500 ;
	    RECT 844.2000 528.4500 845.4000 528.6000 ;
	    RECT 856.2000 528.4500 857.4000 528.6000 ;
	    RECT 844.2000 527.5500 857.4000 528.4500 ;
	    RECT 844.2000 527.4000 845.4000 527.5500 ;
	    RECT 856.2000 527.4000 857.4000 527.5500 ;
	    RECT 837.0000 526.2000 838.2000 526.5000 ;
	    RECT 784.2000 524.5500 806.8500 525.4500 ;
	    RECT 808.2000 525.4500 809.4000 525.6000 ;
	    RECT 834.6000 525.4500 835.8000 525.6000 ;
	    RECT 808.2000 524.5500 835.8000 525.4500 ;
	    RECT 784.2000 524.4000 785.4000 524.5500 ;
	    RECT 808.2000 524.4000 809.4000 524.5500 ;
	    RECT 834.6000 524.4000 835.8000 524.5500 ;
	    RECT 839.4000 524.4000 840.6000 525.6000 ;
	    RECT 841.5000 524.4000 841.8000 525.6000 ;
	    RECT 673.8000 521.5500 694.0500 522.4500 ;
	    RECT 695.4000 522.4500 696.6000 522.6000 ;
	    RECT 697.8000 522.4500 699.0000 522.6000 ;
	    RECT 695.4000 521.5500 699.0000 522.4500 ;
	    RECT 673.8000 521.4000 675.0000 521.5500 ;
	    RECT 695.4000 521.4000 696.6000 521.5500 ;
	    RECT 697.8000 521.4000 699.0000 521.5500 ;
	    RECT 561.0000 519.0000 562.5000 520.2000 ;
	    RECT 561.0000 513.3000 562.2000 519.0000 ;
	    RECT 563.4000 513.3000 564.6000 516.3000 ;
	    RECT 575.4000 513.3000 576.6000 520.5000 ;
	    RECT 633.0000 520.2000 635.7000 521.4000 ;
	    RECT 637.8000 520.2000 641.1000 521.4000 ;
	    RECT 642.6000 520.2000 645.9000 521.4000 ;
	    RECT 647.4000 520.2000 651.0000 521.4000 ;
	    RECT 699.9000 520.8000 700.2000 522.3000 ;
	    RECT 702.3000 521.4000 704.1000 522.6000 ;
	    RECT 705.0000 522.4500 706.2000 522.6000 ;
	    RECT 721.8000 522.4500 723.0000 522.6000 ;
	    RECT 705.0000 521.5500 723.0000 522.4500 ;
	    RECT 705.0000 521.4000 706.2000 521.5500 ;
	    RECT 721.8000 521.4000 723.0000 521.5500 ;
	    RECT 724.2000 521.4000 725.4000 522.6000 ;
	    RECT 577.8000 519.4500 579.0000 519.6000 ;
	    RECT 594.6000 519.4500 595.8000 519.6000 ;
	    RECT 604.2000 519.4500 605.4000 519.6000 ;
	    RECT 577.8000 518.5500 605.4000 519.4500 ;
	    RECT 577.8000 518.4000 579.0000 518.5500 ;
	    RECT 594.6000 518.4000 595.8000 518.5500 ;
	    RECT 604.2000 518.4000 605.4000 518.5500 ;
	    RECT 577.8000 517.2000 579.0000 517.5000 ;
	    RECT 577.8000 513.3000 579.0000 516.3000 ;
	    RECT 630.6000 513.3000 631.8000 519.3000 ;
	    RECT 633.0000 513.3000 634.2000 520.2000 ;
	    RECT 635.4000 513.3000 636.6000 519.3000 ;
	    RECT 637.8000 513.3000 639.0000 520.2000 ;
	    RECT 640.2000 513.3000 641.4000 519.3000 ;
	    RECT 642.6000 513.3000 643.8000 520.2000 ;
	    RECT 645.0000 513.3000 646.2000 519.3000 ;
	    RECT 647.4000 513.3000 648.6000 520.2000 ;
	    RECT 652.2000 519.4500 653.4000 519.6000 ;
	    RECT 671.4000 519.4500 672.6000 519.6000 ;
	    RECT 649.8000 513.3000 651.0000 519.3000 ;
	    RECT 652.2000 518.5500 672.6000 519.4500 ;
	    RECT 652.2000 518.4000 653.4000 518.5500 ;
	    RECT 671.4000 518.4000 672.6000 518.5500 ;
	    RECT 671.4000 517.2000 672.6000 517.5000 ;
	    RECT 671.4000 513.3000 672.6000 516.3000 ;
	    RECT 673.8000 513.3000 675.0000 520.5000 ;
	    RECT 698.1000 519.3000 703.5000 519.9000 ;
	    RECT 705.0000 519.3000 705.9000 520.5000 ;
	    RECT 724.2000 520.2000 725.4000 520.5000 ;
	    RECT 726.6000 519.3000 727.8000 523.5000 ;
	    RECT 731.4000 522.4500 732.6000 522.6000 ;
	    RECT 745.8000 522.4500 747.0000 522.6000 ;
	    RECT 731.4000 521.5500 747.0000 522.4500 ;
	    RECT 731.4000 521.4000 732.6000 521.5500 ;
	    RECT 745.8000 521.4000 747.0000 521.5500 ;
	    RECT 762.6000 522.4500 763.8000 522.6000 ;
	    RECT 777.0000 522.4500 778.2000 522.6000 ;
	    RECT 762.6000 521.5500 778.2000 522.4500 ;
	    RECT 762.6000 521.4000 763.8000 521.5500 ;
	    RECT 777.0000 521.4000 778.2000 521.5500 ;
	    RECT 781.8000 521.4000 783.0000 522.6000 ;
	    RECT 697.8000 519.0000 703.8000 519.3000 ;
	    RECT 697.8000 513.3000 699.0000 519.0000 ;
	    RECT 700.2000 513.3000 701.4000 518.1000 ;
	    RECT 702.6000 513.3000 703.8000 519.0000 ;
	    RECT 705.0000 513.3000 706.2000 519.3000 ;
	    RECT 724.2000 513.3000 725.4000 519.3000 ;
	    RECT 726.6000 518.4000 729.3000 519.3000 ;
	    RECT 743.4000 518.4000 744.6000 519.6000 ;
	    RECT 728.1000 513.3000 729.3000 518.4000 ;
	    RECT 743.4000 517.2000 744.6000 517.5000 ;
	    RECT 743.4000 513.3000 744.6000 516.3000 ;
	    RECT 745.8000 513.3000 747.0000 520.5000 ;
	    RECT 753.0000 519.4500 754.2000 519.6000 ;
	    RECT 760.2000 519.4500 761.4000 519.6000 ;
	    RECT 753.0000 518.5500 761.4000 519.4500 ;
	    RECT 753.0000 518.4000 754.2000 518.5500 ;
	    RECT 760.2000 518.4000 761.4000 518.5500 ;
	    RECT 760.2000 517.2000 761.4000 517.5000 ;
	    RECT 760.2000 513.3000 761.4000 516.3000 ;
	    RECT 762.6000 513.3000 763.8000 520.5000 ;
	    RECT 781.8000 520.2000 783.0000 520.5000 ;
	    RECT 784.2000 519.3000 785.4000 523.5000 ;
	    RECT 808.2000 519.3000 809.4000 523.5000 ;
	    RECT 844.2000 522.6000 845.1000 526.5000 ;
	    RECT 861.0000 523.5000 862.2000 539.7000 ;
	    RECT 880.2000 533.7000 881.4000 539.7000 ;
	    RECT 882.6000 526.5000 883.8000 539.7000 ;
	    RECT 885.0000 533.7000 886.2000 539.7000 ;
	    RECT 904.2000 533.7000 905.4000 539.7000 ;
	    RECT 885.0000 529.5000 886.2000 529.8000 ;
	    RECT 885.0000 527.4000 886.2000 528.6000 ;
	    RECT 873.0000 525.4500 874.2000 525.6000 ;
	    RECT 882.6000 525.4500 883.8000 525.6000 ;
	    RECT 873.0000 524.5500 883.8000 525.4500 ;
	    RECT 873.0000 524.4000 874.2000 524.5500 ;
	    RECT 882.6000 524.4000 883.8000 524.5500 ;
	    RECT 906.6000 523.5000 907.8000 539.7000 ;
	    RECT 976.2000 527.1000 977.4000 539.7000 ;
	    RECT 978.6000 528.0000 979.8000 539.7000 ;
	    RECT 982.8000 534.6000 984.0000 539.7000 ;
	    RECT 981.0000 533.7000 984.0000 534.6000 ;
	    RECT 987.0000 533.7000 988.2000 539.7000 ;
	    RECT 989.4000 533.7000 990.6000 539.7000 ;
	    RECT 991.8000 533.7000 993.0000 539.7000 ;
	    RECT 995.7000 533.7000 997.5000 539.7000 ;
	    RECT 981.0000 532.5000 982.2000 533.7000 ;
	    RECT 989.4000 532.8000 990.3000 533.7000 ;
	    RECT 986.1000 531.9000 991.5000 532.8000 ;
	    RECT 995.4000 532.5000 996.6000 533.7000 ;
	    RECT 986.1000 531.6000 987.3000 531.9000 ;
	    RECT 990.3000 531.6000 991.5000 531.9000 ;
	    RECT 981.0000 529.5000 982.2000 529.8000 ;
	    RECT 987.9000 529.5000 989.1000 529.8000 ;
	    RECT 981.0000 528.6000 989.1000 529.5000 ;
	    RECT 990.0000 529.5000 993.3000 530.4000 ;
	    RECT 990.0000 527.7000 990.9000 529.5000 ;
	    RECT 992.1000 529.2000 993.3000 529.5000 ;
	    RECT 995.7000 529.8000 997.8000 531.0000 ;
	    RECT 995.7000 528.3000 996.6000 529.8000 ;
	    RECT 983.7000 527.1000 990.9000 527.7000 ;
	    RECT 976.2000 526.8000 990.9000 527.1000 ;
	    RECT 993.0000 527.4000 996.6000 528.3000 ;
	    RECT 1000.2000 527.7000 1001.4000 539.7000 ;
	    RECT 976.2000 526.5000 984.9000 526.8000 ;
	    RECT 976.2000 526.2000 984.6000 526.5000 ;
	    RECT 979.5000 524.4000 984.9000 525.3000 ;
	    RECT 985.8000 524.4000 987.0000 525.6000 ;
	    RECT 979.5000 524.1000 980.7000 524.4000 ;
	    RECT 810.6000 521.4000 811.8000 522.6000 ;
	    RECT 842.7000 522.3000 845.1000 522.6000 ;
	    RECT 810.6000 520.2000 811.8000 520.5000 ;
	    RECT 781.8000 513.3000 783.0000 519.3000 ;
	    RECT 784.2000 518.4000 786.9000 519.3000 ;
	    RECT 785.7000 513.3000 786.9000 518.4000 ;
	    RECT 806.7000 518.4000 809.4000 519.3000 ;
	    RECT 806.7000 513.3000 807.9000 518.4000 ;
	    RECT 810.6000 513.3000 811.8000 519.3000 ;
	    RECT 837.0000 513.3000 838.2000 522.3000 ;
	    RECT 842.4000 521.7000 845.1000 522.3000 ;
	    RECT 861.0000 522.4500 862.2000 522.6000 ;
	    RECT 868.2000 522.4500 869.4000 522.6000 ;
	    RECT 842.4000 513.3000 843.6000 521.7000 ;
	    RECT 861.0000 521.5500 869.4000 522.4500 ;
	    RECT 861.0000 521.4000 862.2000 521.5500 ;
	    RECT 868.2000 521.4000 869.4000 521.5500 ;
	    RECT 870.6000 522.4500 871.8000 522.6000 ;
	    RECT 880.2000 522.4500 881.4000 522.6000 ;
	    RECT 870.6000 521.5500 881.4000 522.4500 ;
	    RECT 870.6000 521.4000 871.8000 521.5500 ;
	    RECT 880.2000 521.4000 881.4000 521.5500 ;
	    RECT 858.6000 518.4000 859.8000 519.6000 ;
	    RECT 858.6000 517.2000 859.8000 517.5000 ;
	    RECT 858.6000 513.3000 859.8000 516.3000 ;
	    RECT 861.0000 513.3000 862.2000 520.5000 ;
	    RECT 880.2000 520.2000 881.4000 520.5000 ;
	    RECT 882.6000 519.3000 883.8000 523.5000 ;
	    RECT 981.9000 522.6000 983.1000 522.9000 ;
	    RECT 993.0000 522.6000 993.9000 527.4000 ;
	    RECT 1002.6000 526.8000 1003.8000 539.7000 ;
	    RECT 1021.8000 528.6000 1023.0000 539.7000 ;
	    RECT 1024.2001 529.5000 1025.4000 539.7000 ;
	    RECT 1021.8000 527.7000 1025.1000 528.6000 ;
	    RECT 1026.6000 527.7000 1027.8000 539.7000 ;
	    RECT 1043.4000 539.4000 1044.6000 540.6000 ;
	    RECT 1045.8000 528.6000 1047.0000 539.7000 ;
	    RECT 1048.2001 529.5000 1049.4000 539.7000 ;
	    RECT 1045.8000 527.7000 1049.1000 528.6000 ;
	    RECT 1050.6000 527.7000 1051.8000 539.7000 ;
	    RECT 1077.0000 533.7000 1078.2001 539.7000 ;
	    RECT 1079.4000 533.7000 1080.6000 539.7000 ;
	    RECT 997.5000 526.5000 1003.8000 526.8000 ;
	    RECT 1024.2001 526.8000 1025.1000 527.7000 ;
	    RECT 997.5000 525.9000 1001.7000 526.5000 ;
	    RECT 997.5000 525.6000 998.7000 525.9000 ;
	    RECT 1024.2001 525.6000 1026.0000 526.8000 ;
	    RECT 999.9000 524.7000 1001.1000 525.0000 ;
	    RECT 995.4000 523.8000 1001.1000 524.7000 ;
	    RECT 1002.6000 524.4000 1003.8000 525.6000 ;
	    RECT 1021.8000 524.4000 1023.0000 525.6000 ;
	    RECT 995.4000 523.5000 996.6000 523.8000 ;
	    RECT 906.6000 522.4500 907.8000 522.6000 ;
	    RECT 973.8000 522.4500 975.0000 522.6000 ;
	    RECT 906.6000 521.5500 975.0000 522.4500 ;
	    RECT 906.6000 521.4000 907.8000 521.5500 ;
	    RECT 973.8000 521.4000 975.0000 521.5500 ;
	    RECT 977.4000 521.4000 977.7000 522.6000 ;
	    RECT 978.6000 521.4000 979.8000 522.6000 ;
	    RECT 980.7000 521.7000 993.9000 522.6000 ;
	    RECT 880.2000 513.3000 881.4000 519.3000 ;
	    RECT 882.6000 518.4000 885.3000 519.3000 ;
	    RECT 904.2000 518.4000 905.4000 519.6000 ;
	    RECT 884.1000 513.3000 885.3000 518.4000 ;
	    RECT 904.2000 517.2000 905.4000 517.5000 ;
	    RECT 904.2000 513.3000 905.4000 516.3000 ;
	    RECT 906.6000 513.3000 907.8000 520.5000 ;
	    RECT 976.2000 513.3000 977.4000 520.5000 ;
	    RECT 978.6000 513.3000 979.8000 519.3000 ;
	    RECT 983.7000 518.4000 984.6000 521.7000 ;
	    RECT 992.1000 521.4000 993.3000 521.7000 ;
	    RECT 1002.6000 520.8000 1003.8000 523.5000 ;
	    RECT 1021.8000 523.2000 1023.0000 523.5000 ;
	    RECT 1024.2001 521.1000 1025.1000 525.6000 ;
	    RECT 1026.9000 524.4000 1027.8000 527.7000 ;
	    RECT 1048.2001 526.8000 1049.1000 527.7000 ;
	    RECT 1048.2001 525.6000 1050.0000 526.8000 ;
	    RECT 1045.8000 524.4000 1047.0000 525.6000 ;
	    RECT 1026.6000 523.5000 1027.8000 524.4000 ;
	    RECT 1045.8000 523.2000 1047.0000 523.5000 ;
	    RECT 1026.6000 522.4500 1027.8000 522.6000 ;
	    RECT 1043.4000 522.4500 1044.6000 522.6000 ;
	    RECT 1026.6000 521.5500 1044.6000 522.4500 ;
	    RECT 1026.6000 521.4000 1027.8000 521.5500 ;
	    RECT 1043.4000 521.4000 1044.6000 521.5500 ;
	    RECT 1048.2001 521.1000 1049.1000 525.6000 ;
	    RECT 1050.9000 524.4000 1051.8000 527.7000 ;
	    RECT 1079.7001 527.4000 1080.6000 533.7000 ;
	    RECT 1081.8000 528.3000 1083.0000 539.7000 ;
	    RECT 1084.2001 527.7000 1085.4000 539.7000 ;
	    RECT 1108.2001 533.7000 1109.4000 539.7000 ;
	    RECT 1110.6000 533.7000 1111.8000 539.7000 ;
	    RECT 1079.7001 526.5000 1083.3000 527.4000 ;
	    RECT 1084.5000 526.5000 1085.4000 527.7000 ;
	    RECT 1110.9000 527.4000 1111.8000 533.7000 ;
	    RECT 1113.0000 528.3000 1114.2001 539.7000 ;
	    RECT 1115.4000 527.7000 1116.6000 539.7000 ;
	    RECT 1141.8000 533.7000 1143.0000 539.7000 ;
	    RECT 1110.9000 526.5000 1114.5000 527.4000 ;
	    RECT 1115.7001 526.5000 1116.6000 527.7000 ;
	    RECT 1144.2001 526.5000 1145.4000 539.7000 ;
	    RECT 1146.6000 533.7000 1147.8000 539.7000 ;
	    RECT 1165.8000 533.7000 1167.0000 539.7000 ;
	    RECT 1146.6000 529.5000 1147.8000 529.8000 ;
	    RECT 1146.6000 527.4000 1147.8000 528.6000 ;
	    RECT 1168.2001 526.5000 1169.4000 539.7000 ;
	    RECT 1170.6000 533.7000 1171.8000 539.7000 ;
	    RECT 1170.6000 529.5000 1171.8000 529.8000 ;
	    RECT 1199.4000 528.6000 1200.6000 539.7000 ;
	    RECT 1201.8000 529.5000 1203.0000 539.7000 ;
	    RECT 1204.2001 538.8000 1210.2001 539.7000 ;
	    RECT 1204.2001 528.6000 1205.4000 538.8000 ;
	    RECT 1170.6000 527.4000 1171.8000 528.6000 ;
	    RECT 1199.4000 527.7000 1205.4000 528.6000 ;
	    RECT 1206.6000 527.7000 1207.8000 537.9000 ;
	    RECT 1209.0000 527.7000 1210.2001 538.8000 ;
	    RECT 1235.4000 533.7000 1236.6000 539.7000 ;
	    RECT 1237.8000 534.3000 1239.0000 539.7000 ;
	    RECT 1235.7001 533.4000 1236.6000 533.7000 ;
	    RECT 1240.2001 533.7000 1241.4000 539.7000 ;
	    RECT 1242.6000 533.7000 1243.8000 539.7000 ;
	    RECT 1266.6000 533.7000 1267.8000 539.7000 ;
	    RECT 1269.0000 533.7000 1270.2001 539.7000 ;
	    RECT 1271.4000 534.3000 1272.6000 539.7000 ;
	    RECT 1240.2001 533.4000 1241.1000 533.7000 ;
	    RECT 1235.7001 532.5000 1241.1000 533.4000 ;
	    RECT 1269.3000 533.4000 1270.2001 533.7000 ;
	    RECT 1273.8000 533.7000 1275.0000 539.7000 ;
	    RECT 1285.8000 533.7000 1287.0000 539.7000 ;
	    RECT 1273.8000 533.4000 1274.7001 533.7000 ;
	    RECT 1269.3000 532.5000 1274.7001 533.4000 ;
	    RECT 1235.7001 529.5000 1236.6000 532.5000 ;
	    RECT 1237.8000 531.4500 1239.0000 531.6000 ;
	    RECT 1271.4000 531.4500 1272.6000 531.6000 ;
	    RECT 1237.8000 530.5500 1272.6000 531.4500 ;
	    RECT 1237.8000 530.4000 1239.0000 530.5500 ;
	    RECT 1271.4000 530.4000 1272.6000 530.5500 ;
	    RECT 1273.8000 529.5000 1274.7001 532.5000 ;
	    RECT 1237.8000 529.2000 1239.0000 529.5000 ;
	    RECT 1271.4000 529.2000 1272.6000 529.5000 ;
	    RECT 1206.6000 526.8000 1207.5000 527.7000 ;
	    RECT 1235.4000 527.4000 1236.6000 528.6000 ;
	    RECT 1242.6000 527.4000 1243.8000 528.6000 ;
	    RECT 1259.4000 528.4500 1260.6000 528.6000 ;
	    RECT 1266.6000 528.4500 1267.8000 528.6000 ;
	    RECT 1259.4000 527.5500 1267.8000 528.4500 ;
	    RECT 1259.4000 527.4000 1260.6000 527.5500 ;
	    RECT 1266.6000 527.4000 1267.8000 527.5500 ;
	    RECT 1273.8000 528.4500 1275.0000 528.6000 ;
	    RECT 1285.8000 528.4500 1287.0000 528.6000 ;
	    RECT 1273.8000 527.5500 1287.0000 528.4500 ;
	    RECT 1273.8000 527.4000 1275.0000 527.5500 ;
	    RECT 1285.8000 527.4000 1287.0000 527.5500 ;
	    RECT 1204.5000 526.5000 1207.5000 526.8000 ;
	    RECT 1209.0000 526.5000 1210.2001 526.8000 ;
	    RECT 1079.4000 524.4000 1080.6000 525.6000 ;
	    RECT 1050.6000 523.5000 1051.8000 524.4000 ;
	    RECT 1077.0000 523.5000 1078.2001 523.8000 ;
	    RECT 1079.7001 523.2000 1080.6000 523.5000 ;
	    RECT 1050.6000 522.4500 1051.8000 522.6000 ;
	    RECT 1060.2001 522.4500 1061.4000 522.6000 ;
	    RECT 1050.6000 521.5500 1061.4000 522.4500 ;
	    RECT 1050.6000 521.4000 1051.8000 521.5500 ;
	    RECT 1060.2001 521.4000 1061.4000 521.5500 ;
	    RECT 1062.6000 522.4500 1063.8000 522.6000 ;
	    RECT 1077.0000 522.4500 1078.2001 522.6000 ;
	    RECT 1062.6000 521.5500 1078.2001 522.4500 ;
	    RECT 1079.7001 522.3000 1081.2001 523.2000 ;
	    RECT 1080.0000 522.0000 1081.2001 522.3000 ;
	    RECT 1062.6000 521.4000 1063.8000 521.5500 ;
	    RECT 1077.0000 521.4000 1078.2001 521.5500 ;
	    RECT 1082.4000 521.4000 1083.3000 526.5000 ;
	    RECT 1084.2001 525.4500 1085.4000 525.6000 ;
	    RECT 1105.8000 525.4500 1107.0000 525.6000 ;
	    RECT 1084.2001 524.5500 1107.0000 525.4500 ;
	    RECT 1084.2001 524.4000 1085.4000 524.5500 ;
	    RECT 1105.8000 524.4000 1107.0000 524.5500 ;
	    RECT 1110.6000 524.4000 1111.8000 525.6000 ;
	    RECT 1108.2001 523.5000 1109.4000 523.8000 ;
	    RECT 1082.4000 521.1000 1083.6000 521.4000 ;
	    RECT 998.1000 519.9000 1003.8000 520.8000 ;
	    RECT 998.1000 519.6000 999.3000 519.9000 ;
	    RECT 981.0000 516.3000 982.2000 517.5000 ;
	    RECT 983.4000 517.2000 984.6000 518.4000 ;
	    RECT 986.1000 518.1000 987.3000 518.4000 ;
	    RECT 986.1000 517.2000 990.3000 518.1000 ;
	    RECT 989.4000 516.3000 990.3000 517.2000 ;
	    RECT 995.4000 516.3000 996.6000 517.5000 ;
	    RECT 981.0000 515.4000 984.0000 516.3000 ;
	    RECT 982.8000 513.3000 984.0000 515.4000 ;
	    RECT 986.7000 513.3000 988.2000 516.3000 ;
	    RECT 989.4000 513.3000 990.6000 516.3000 ;
	    RECT 991.8000 513.3000 993.0000 516.3000 ;
	    RECT 995.4000 515.4000 997.5000 516.3000 ;
	    RECT 995.7000 513.3000 997.5000 515.4000 ;
	    RECT 1000.2000 513.3000 1001.4000 519.0000 ;
	    RECT 1002.6000 513.3000 1003.8000 519.9000 ;
	    RECT 1021.8000 520.2000 1025.1000 521.1000 ;
	    RECT 1021.8000 513.3000 1023.0000 520.2000 ;
	    RECT 1024.2001 513.3000 1025.4000 519.3000 ;
	    RECT 1026.6000 513.3000 1027.8000 520.5000 ;
	    RECT 1045.8000 520.2000 1049.1000 521.1000 ;
	    RECT 1079.1000 520.5000 1083.6000 521.1000 ;
	    RECT 1045.8000 513.3000 1047.0000 520.2000 ;
	    RECT 1048.2001 513.3000 1049.4000 519.3000 ;
	    RECT 1050.6000 513.3000 1051.8000 520.5000 ;
	    RECT 1077.3000 520.2000 1083.6000 520.5000 ;
	    RECT 1077.3000 519.6000 1080.0000 520.2000 ;
	    RECT 1077.3000 519.3000 1078.2001 519.6000 ;
	    RECT 1084.5000 519.3000 1085.4000 523.5000 ;
	    RECT 1110.9000 523.2000 1111.8000 523.5000 ;
	    RECT 1091.4000 522.4500 1092.6000 522.6000 ;
	    RECT 1103.4000 522.4500 1104.6000 522.6000 ;
	    RECT 1108.2001 522.4500 1109.4000 522.6000 ;
	    RECT 1091.4000 521.5500 1109.4000 522.4500 ;
	    RECT 1110.9000 522.3000 1112.4000 523.2000 ;
	    RECT 1111.2001 522.0000 1112.4000 522.3000 ;
	    RECT 1091.4000 521.4000 1092.6000 521.5500 ;
	    RECT 1103.4000 521.4000 1104.6000 521.5500 ;
	    RECT 1108.2001 521.4000 1109.4000 521.5500 ;
	    RECT 1113.6000 521.4000 1114.5000 526.5000 ;
	    RECT 1115.4000 525.4500 1116.6000 525.6000 ;
	    RECT 1141.8000 525.4500 1143.0000 525.6000 ;
	    RECT 1115.4000 524.5500 1143.0000 525.4500 ;
	    RECT 1115.4000 524.4000 1116.6000 524.5500 ;
	    RECT 1141.8000 524.4000 1143.0000 524.5500 ;
	    RECT 1144.2001 525.4500 1145.4000 525.6000 ;
	    RECT 1168.2001 525.4500 1169.4000 525.6000 ;
	    RECT 1192.2001 525.4500 1193.4000 525.6000 ;
	    RECT 1144.2001 524.5500 1166.8500 525.4500 ;
	    RECT 1144.2001 524.4000 1145.4000 524.5500 ;
	    RECT 1113.6000 521.1000 1114.8000 521.4000 ;
	    RECT 1110.3000 520.5000 1114.8000 521.1000 ;
	    RECT 1108.5000 520.2000 1114.8000 520.5000 ;
	    RECT 1108.5000 519.6000 1111.2001 520.2000 ;
	    RECT 1108.5000 519.3000 1109.4000 519.6000 ;
	    RECT 1115.7001 519.3000 1116.6000 523.5000 ;
	    RECT 1117.8000 522.4500 1119.0000 522.6000 ;
	    RECT 1139.4000 522.4500 1140.6000 522.6000 ;
	    RECT 1141.8000 522.4500 1143.0000 522.6000 ;
	    RECT 1117.8000 521.5500 1143.0000 522.4500 ;
	    RECT 1117.8000 521.4000 1119.0000 521.5500 ;
	    RECT 1139.4000 521.4000 1140.6000 521.5500 ;
	    RECT 1141.8000 521.4000 1143.0000 521.5500 ;
	    RECT 1141.8000 520.2000 1143.0000 520.5000 ;
	    RECT 1144.2001 519.3000 1145.4000 523.5000 ;
	    RECT 1165.9501 522.6000 1166.8500 524.5500 ;
	    RECT 1168.2001 524.5500 1193.4000 525.4500 ;
	    RECT 1168.2001 524.4000 1169.4000 524.5500 ;
	    RECT 1192.2001 524.4000 1193.4000 524.5500 ;
	    RECT 1199.4000 524.4000 1200.6000 525.6000 ;
	    RECT 1201.5000 524.7000 1201.8000 526.2000 ;
	    RECT 1206.3000 525.9000 1207.5000 526.5000 ;
	    RECT 1204.2001 524.4000 1205.4000 525.6000 ;
	    RECT 1209.0000 525.4500 1210.2001 525.6000 ;
	    RECT 1228.2001 525.4500 1229.4000 525.6000 ;
	    RECT 1209.0000 524.5500 1229.4000 525.4500 ;
	    RECT 1209.0000 524.4000 1210.2001 524.5500 ;
	    RECT 1228.2001 524.4000 1229.4000 524.5500 ;
	    RECT 1201.8000 523.5000 1203.0000 523.8000 ;
	    RECT 1206.3000 523.5000 1207.5000 524.4000 ;
	    RECT 1165.8000 521.4000 1167.0000 522.6000 ;
	    RECT 1165.8000 520.2000 1167.0000 520.5000 ;
	    RECT 1168.2001 519.3000 1169.4000 523.5000 ;
	    RECT 1170.6000 522.4500 1171.8000 522.6000 ;
	    RECT 1201.8000 522.4500 1203.0000 522.6000 ;
	    RECT 1170.6000 521.5500 1203.0000 522.4500 ;
	    RECT 1170.6000 521.4000 1171.8000 521.5500 ;
	    RECT 1201.8000 521.4000 1203.0000 521.5500 ;
	    RECT 1204.5000 519.3000 1205.4000 523.5000 ;
	    RECT 1235.7001 522.6000 1236.6000 526.5000 ;
	    RECT 1242.6000 526.2000 1243.8000 526.5000 ;
	    RECT 1266.6000 526.2000 1267.8000 526.5000 ;
	    RECT 1239.0000 524.4000 1239.3000 525.6000 ;
	    RECT 1240.2001 524.4000 1241.4000 525.6000 ;
	    RECT 1269.0000 524.4000 1270.2001 525.6000 ;
	    RECT 1271.1000 524.4000 1271.4000 525.6000 ;
	    RECT 1273.8000 522.6000 1274.7001 526.5000 ;
	    RECT 1288.2001 523.5000 1289.4000 539.7000 ;
	    RECT 1312.2001 527.7000 1313.4000 539.7000 ;
	    RECT 1316.1000 528.6000 1317.3000 539.7000 ;
	    RECT 1318.5000 533.7000 1319.7001 539.7000 ;
	    RECT 1333.8000 533.7000 1335.0000 539.7000 ;
	    RECT 1318.2001 530.4000 1319.4000 531.6000 ;
	    RECT 1318.5000 529.5000 1319.4000 530.4000 ;
	    RECT 1316.1000 527.7000 1317.6000 528.6000 ;
	    RECT 1290.6000 525.4500 1291.8000 525.6000 ;
	    RECT 1314.6000 525.4500 1315.8000 525.6000 ;
	    RECT 1290.6000 524.5500 1315.8000 525.4500 ;
	    RECT 1290.6000 524.4000 1291.8000 524.5500 ;
	    RECT 1314.6000 524.4000 1315.8000 524.5500 ;
	    RECT 1314.6000 523.2000 1315.8000 523.5000 ;
	    RECT 1316.7001 522.6000 1317.6000 527.7000 ;
	    RECT 1319.4000 527.4000 1320.6000 528.6000 ;
	    RECT 1336.2001 523.5000 1337.4000 539.7000 ;
	    RECT 1367.4000 533.7000 1368.6000 539.7000 ;
	    RECT 1369.8000 534.3000 1371.0000 539.7000 ;
	    RECT 1367.7001 533.4000 1368.6000 533.7000 ;
	    RECT 1372.2001 533.7000 1373.4000 539.7000 ;
	    RECT 1374.6000 533.7000 1375.8000 539.7000 ;
	    RECT 1401.0000 533.7000 1402.2001 539.7000 ;
	    RECT 1403.4000 533.7000 1404.6000 539.7000 ;
	    RECT 1405.8000 534.3000 1407.0000 539.7000 ;
	    RECT 1372.2001 533.4000 1373.1000 533.7000 ;
	    RECT 1367.7001 532.5000 1373.1000 533.4000 ;
	    RECT 1403.7001 533.4000 1404.6000 533.7000 ;
	    RECT 1408.2001 533.7000 1409.4000 539.7000 ;
	    RECT 1432.2001 533.7000 1433.4000 539.7000 ;
	    RECT 1434.6000 533.7000 1435.8000 539.7000 ;
	    RECT 1437.0000 534.3000 1438.2001 539.7000 ;
	    RECT 1408.2001 533.4000 1409.1000 533.7000 ;
	    RECT 1403.7001 532.5000 1409.1000 533.4000 ;
	    RECT 1434.9000 533.4000 1435.8000 533.7000 ;
	    RECT 1439.4000 533.7000 1440.6000 539.7000 ;
	    RECT 1463.4000 533.7000 1464.6000 539.7000 ;
	    RECT 1465.8000 533.7000 1467.0000 539.7000 ;
	    RECT 1468.2001 534.3000 1469.4000 539.7000 ;
	    RECT 1439.4000 533.4000 1440.3000 533.7000 ;
	    RECT 1434.9000 532.5000 1440.3000 533.4000 ;
	    RECT 1466.1000 533.4000 1467.0000 533.7000 ;
	    RECT 1470.6000 533.7000 1471.8000 539.7000 ;
	    RECT 1494.6000 533.7000 1495.8000 539.7000 ;
	    RECT 1497.0000 534.3000 1498.2001 539.7000 ;
	    RECT 1470.6000 533.4000 1471.5000 533.7000 ;
	    RECT 1466.1000 532.5000 1471.5000 533.4000 ;
	    RECT 1367.7001 529.5000 1368.6000 532.5000 ;
	    RECT 1369.8000 530.4000 1371.0000 531.6000 ;
	    RECT 1386.6000 531.4500 1387.8000 531.6000 ;
	    RECT 1405.8000 531.4500 1407.0000 531.6000 ;
	    RECT 1386.6000 530.5500 1407.0000 531.4500 ;
	    RECT 1386.6000 530.4000 1387.8000 530.5500 ;
	    RECT 1405.8000 530.4000 1407.0000 530.5500 ;
	    RECT 1408.2001 529.5000 1409.1000 532.5000 ;
	    RECT 1437.0000 531.4500 1438.2001 531.6000 ;
	    RECT 1429.9501 530.5500 1438.2001 531.4500 ;
	    RECT 1369.8000 529.2000 1371.0000 529.5000 ;
	    RECT 1405.8000 529.2000 1407.0000 529.5000 ;
	    RECT 1367.4000 527.4000 1368.6000 528.6000 ;
	    RECT 1374.6000 527.4000 1375.8000 528.6000 ;
	    RECT 1379.4000 528.4500 1380.6000 528.6000 ;
	    RECT 1393.8000 528.4500 1395.0000 528.6000 ;
	    RECT 1401.0000 528.4500 1402.2001 528.6000 ;
	    RECT 1379.4000 527.5500 1402.2001 528.4500 ;
	    RECT 1379.4000 527.4000 1380.6000 527.5500 ;
	    RECT 1393.8000 527.4000 1395.0000 527.5500 ;
	    RECT 1401.0000 527.4000 1402.2001 527.5500 ;
	    RECT 1408.2001 528.4500 1409.4000 528.6000 ;
	    RECT 1429.9501 528.4500 1430.8500 530.5500 ;
	    RECT 1437.0000 530.4000 1438.2001 530.5500 ;
	    RECT 1439.4000 529.5000 1440.3000 532.5000 ;
	    RECT 1446.6000 531.4500 1447.8000 531.6000 ;
	    RECT 1465.8000 531.4500 1467.0000 531.6000 ;
	    RECT 1446.6000 530.5500 1467.0000 531.4500 ;
	    RECT 1446.6000 530.4000 1447.8000 530.5500 ;
	    RECT 1465.8000 530.4000 1467.0000 530.5500 ;
	    RECT 1468.2001 530.4000 1469.4000 531.6000 ;
	    RECT 1470.6000 529.5000 1471.5000 532.5000 ;
	    RECT 1494.9000 533.4000 1495.8000 533.7000 ;
	    RECT 1499.4000 533.7000 1500.6000 539.7000 ;
	    RECT 1501.8000 533.7000 1503.0000 539.7000 ;
	    RECT 1521.0000 533.7000 1522.2001 539.7000 ;
	    RECT 1499.4000 533.4000 1500.3000 533.7000 ;
	    RECT 1494.9000 532.5000 1500.3000 533.4000 ;
	    RECT 1494.9000 529.5000 1495.8000 532.5000 ;
	    RECT 1497.0000 530.4000 1498.2001 531.6000 ;
	    RECT 1521.0000 529.5000 1522.2001 529.8000 ;
	    RECT 1437.0000 529.2000 1438.2001 529.5000 ;
	    RECT 1468.2001 529.2000 1469.4000 529.5000 ;
	    RECT 1497.0000 529.2000 1498.2001 529.5000 ;
	    RECT 1408.2001 527.5500 1430.8500 528.4500 ;
	    RECT 1432.2001 528.4500 1433.4000 528.6000 ;
	    RECT 1434.6000 528.4500 1435.8000 528.6000 ;
	    RECT 1432.2001 527.5500 1435.8000 528.4500 ;
	    RECT 1408.2001 527.4000 1409.4000 527.5500 ;
	    RECT 1432.2001 527.4000 1433.4000 527.5500 ;
	    RECT 1434.6000 527.4000 1435.8000 527.5500 ;
	    RECT 1439.4000 528.4500 1440.6000 528.6000 ;
	    RECT 1449.0000 528.4500 1450.2001 528.6000 ;
	    RECT 1439.4000 527.5500 1450.2001 528.4500 ;
	    RECT 1439.4000 527.4000 1440.6000 527.5500 ;
	    RECT 1449.0000 527.4000 1450.2001 527.5500 ;
	    RECT 1461.0000 528.4500 1462.2001 528.6000 ;
	    RECT 1463.4000 528.4500 1464.6000 528.6000 ;
	    RECT 1461.0000 527.5500 1464.6000 528.4500 ;
	    RECT 1461.0000 527.4000 1462.2001 527.5500 ;
	    RECT 1463.4000 527.4000 1464.6000 527.5500 ;
	    RECT 1470.6000 528.4500 1471.8000 528.6000 ;
	    RECT 1473.0000 528.4500 1474.2001 528.6000 ;
	    RECT 1470.6000 527.5500 1474.2001 528.4500 ;
	    RECT 1470.6000 527.4000 1471.8000 527.5500 ;
	    RECT 1473.0000 527.4000 1474.2001 527.5500 ;
	    RECT 1494.6000 527.4000 1495.8000 528.6000 ;
	    RECT 1501.8000 527.4000 1503.0000 528.6000 ;
	    RECT 1521.0000 527.4000 1522.2001 528.6000 ;
	    RECT 1523.4000 526.5000 1524.6000 539.7000 ;
	    RECT 1525.8000 533.7000 1527.0000 539.7000 ;
	    RECT 1557.0000 527.7000 1558.2001 539.7000 ;
	    RECT 1560.9000 527.7000 1563.9000 539.7000 ;
	    RECT 1566.6000 527.7000 1567.8000 539.7000 ;
	    RECT 1367.7001 522.6000 1368.6000 526.5000 ;
	    RECT 1374.6000 526.2000 1375.8000 526.5000 ;
	    RECT 1401.0000 526.2000 1402.2001 526.5000 ;
	    RECT 1371.0000 524.4000 1371.3000 525.6000 ;
	    RECT 1372.2001 524.4000 1373.4000 525.6000 ;
	    RECT 1403.4000 524.4000 1404.6000 525.6000 ;
	    RECT 1405.5000 524.4000 1405.8000 525.6000 ;
	    RECT 1408.2001 522.6000 1409.1000 526.5000 ;
	    RECT 1432.2001 526.2000 1433.4000 526.5000 ;
	    RECT 1434.6000 524.4000 1435.8000 525.6000 ;
	    RECT 1436.7001 524.4000 1437.0000 525.6000 ;
	    RECT 1439.4000 522.6000 1440.3000 526.5000 ;
	    RECT 1463.4000 526.2000 1464.6000 526.5000 ;
	    RECT 1465.8000 524.4000 1467.0000 525.6000 ;
	    RECT 1467.9000 524.4000 1468.2001 525.6000 ;
	    RECT 1470.6000 522.6000 1471.5000 526.5000 ;
	    RECT 1206.6000 521.4000 1207.8000 522.6000 ;
	    RECT 1235.7001 522.3000 1238.1000 522.6000 ;
	    RECT 1272.3000 522.3000 1274.7001 522.6000 ;
	    RECT 1235.7001 521.7000 1238.4000 522.3000 ;
	    RECT 1077.0000 513.3000 1078.2001 519.3000 ;
	    RECT 1080.9000 513.3000 1082.1000 519.0000 ;
	    RECT 1083.3000 517.8000 1085.4000 519.3000 ;
	    RECT 1083.3000 513.3000 1084.5000 517.8000 ;
	    RECT 1108.2001 513.3000 1109.4000 519.3000 ;
	    RECT 1112.1000 513.3000 1113.3000 519.0000 ;
	    RECT 1114.5000 517.8000 1116.6000 519.3000 ;
	    RECT 1114.5000 513.3000 1115.7001 517.8000 ;
	    RECT 1141.8000 513.3000 1143.0000 519.3000 ;
	    RECT 1144.2001 518.4000 1146.9000 519.3000 ;
	    RECT 1145.7001 513.3000 1146.9000 518.4000 ;
	    RECT 1165.8000 513.3000 1167.0000 519.3000 ;
	    RECT 1168.2001 518.4000 1170.9000 519.3000 ;
	    RECT 1169.7001 513.3000 1170.9000 518.4000 ;
	    RECT 1200.0000 513.3000 1201.2001 519.3000 ;
	    RECT 1203.9000 513.3000 1206.3000 519.3000 ;
	    RECT 1209.0000 513.3000 1210.2001 519.3000 ;
	    RECT 1237.2001 513.3000 1238.4000 521.7000 ;
	    RECT 1242.6000 513.3000 1243.8000 522.3000 ;
	    RECT 1266.6000 513.3000 1267.8000 522.3000 ;
	    RECT 1272.0000 521.7000 1274.7001 522.3000 ;
	    RECT 1288.2001 522.4500 1289.4000 522.6000 ;
	    RECT 1302.6000 522.4500 1303.8000 522.6000 ;
	    RECT 1272.0000 513.3000 1273.2001 521.7000 ;
	    RECT 1288.2001 521.5500 1303.8000 522.4500 ;
	    RECT 1288.2001 521.4000 1289.4000 521.5500 ;
	    RECT 1302.6000 521.4000 1303.8000 521.5500 ;
	    RECT 1312.2001 521.4000 1313.4000 522.6000 ;
	    RECT 1314.3000 520.8000 1314.6000 522.3000 ;
	    RECT 1316.7001 521.4000 1318.5000 522.6000 ;
	    RECT 1319.4000 522.4500 1320.6000 522.6000 ;
	    RECT 1333.8000 522.4500 1335.0000 522.6000 ;
	    RECT 1319.4000 521.5500 1335.0000 522.4500 ;
	    RECT 1319.4000 521.4000 1320.6000 521.5500 ;
	    RECT 1333.8000 521.4000 1335.0000 521.5500 ;
	    RECT 1336.2001 522.4500 1337.4000 522.6000 ;
	    RECT 1341.0000 522.4500 1342.2001 522.6000 ;
	    RECT 1336.2001 521.5500 1342.2001 522.4500 ;
	    RECT 1367.7001 522.3000 1370.1000 522.6000 ;
	    RECT 1406.7001 522.3000 1409.1000 522.6000 ;
	    RECT 1437.9000 522.3000 1440.3000 522.6000 ;
	    RECT 1469.1000 522.3000 1471.5000 522.6000 ;
	    RECT 1367.7001 521.7000 1370.4000 522.3000 ;
	    RECT 1336.2001 521.4000 1337.4000 521.5500 ;
	    RECT 1341.0000 521.4000 1342.2001 521.5500 ;
	    RECT 1283.4000 519.4500 1284.6000 519.6000 ;
	    RECT 1285.8000 519.4500 1287.0000 519.6000 ;
	    RECT 1283.4000 518.5500 1287.0000 519.4500 ;
	    RECT 1283.4000 518.4000 1284.6000 518.5500 ;
	    RECT 1285.8000 518.4000 1287.0000 518.5500 ;
	    RECT 1285.8000 517.2000 1287.0000 517.5000 ;
	    RECT 1285.8000 513.3000 1287.0000 516.3000 ;
	    RECT 1288.2001 513.3000 1289.4000 520.5000 ;
	    RECT 1312.5000 519.3000 1317.9000 519.9000 ;
	    RECT 1319.4000 519.3000 1320.3000 520.5000 ;
	    RECT 1331.4000 519.4500 1332.6000 519.6000 ;
	    RECT 1333.8000 519.4500 1335.0000 519.6000 ;
	    RECT 1312.2001 519.0000 1318.2001 519.3000 ;
	    RECT 1312.2001 513.3000 1313.4000 519.0000 ;
	    RECT 1314.6000 513.3000 1315.8000 518.1000 ;
	    RECT 1317.0000 513.3000 1318.2001 519.0000 ;
	    RECT 1319.4000 513.3000 1320.6000 519.3000 ;
	    RECT 1331.4000 518.5500 1335.0000 519.4500 ;
	    RECT 1331.4000 518.4000 1332.6000 518.5500 ;
	    RECT 1333.8000 518.4000 1335.0000 518.5500 ;
	    RECT 1333.8000 517.2000 1335.0000 517.5000 ;
	    RECT 1333.8000 513.3000 1335.0000 516.3000 ;
	    RECT 1336.2001 513.3000 1337.4000 520.5000 ;
	    RECT 1369.2001 513.3000 1370.4000 521.7000 ;
	    RECT 1374.6000 513.3000 1375.8000 522.3000 ;
	    RECT 1401.0000 513.3000 1402.2001 522.3000 ;
	    RECT 1406.4000 521.7000 1409.1000 522.3000 ;
	    RECT 1406.4000 513.3000 1407.6000 521.7000 ;
	    RECT 1432.2001 513.3000 1433.4000 522.3000 ;
	    RECT 1437.6000 521.7000 1440.3000 522.3000 ;
	    RECT 1437.6000 513.3000 1438.8000 521.7000 ;
	    RECT 1463.4000 513.3000 1464.6000 522.3000 ;
	    RECT 1468.8000 521.7000 1471.5000 522.3000 ;
	    RECT 1494.9000 522.6000 1495.8000 526.5000 ;
	    RECT 1501.8000 526.2000 1503.0000 526.5000 ;
	    RECT 1498.2001 524.4000 1498.5000 525.6000 ;
	    RECT 1499.4000 524.4000 1500.6000 525.6000 ;
	    RECT 1504.2001 525.4500 1505.4000 525.6000 ;
	    RECT 1523.4000 525.4500 1524.6000 525.6000 ;
	    RECT 1504.2001 524.5500 1524.6000 525.4500 ;
	    RECT 1504.2001 524.4000 1505.4000 524.5500 ;
	    RECT 1523.4000 524.4000 1524.6000 524.5500 ;
	    RECT 1537.8000 525.4500 1539.0000 525.6000 ;
	    RECT 1537.8000 524.5500 1555.6500 525.4500 ;
	    RECT 1537.8000 524.4000 1539.0000 524.5500 ;
	    RECT 1494.9000 522.3000 1497.3000 522.6000 ;
	    RECT 1494.9000 521.7000 1497.6000 522.3000 ;
	    RECT 1468.8000 513.3000 1470.0000 521.7000 ;
	    RECT 1496.4000 513.3000 1497.6000 521.7000 ;
	    RECT 1501.8000 513.3000 1503.0000 522.3000 ;
	    RECT 1523.4000 519.3000 1524.6000 523.5000 ;
	    RECT 1525.8000 522.4500 1527.0000 522.6000 ;
	    RECT 1545.0000 522.4500 1546.2001 522.6000 ;
	    RECT 1525.8000 521.5500 1546.2001 522.4500 ;
	    RECT 1554.7500 522.4500 1555.6500 524.5500 ;
	    RECT 1559.4000 524.4000 1560.6000 525.6000 ;
	    RECT 1557.0000 523.5000 1558.2001 523.8000 ;
	    RECT 1562.1000 523.5000 1563.0000 527.7000 ;
	    RECT 1564.2001 524.4000 1565.4000 525.6000 ;
	    RECT 1559.4000 523.2000 1560.6000 523.5000 ;
	    RECT 1564.2001 523.2000 1565.4000 523.5000 ;
	    RECT 1557.0000 522.4500 1558.2001 522.6000 ;
	    RECT 1554.7500 521.5500 1558.2001 522.4500 ;
	    RECT 1525.8000 521.4000 1527.0000 521.5500 ;
	    RECT 1545.0000 521.4000 1546.2001 521.5500 ;
	    RECT 1557.0000 521.4000 1558.2001 521.5500 ;
	    RECT 1559.4000 521.4000 1560.9000 522.3000 ;
	    RECT 1561.8000 521.4000 1563.0000 522.6000 ;
	    RECT 1525.8000 520.2000 1527.0000 520.5000 ;
	    RECT 1559.4000 519.3000 1560.3000 521.4000 ;
	    RECT 1565.4000 520.8000 1565.7001 522.3000 ;
	    RECT 1566.6000 521.4000 1567.8000 522.6000 ;
	    RECT 1562.1000 519.3000 1567.5000 519.9000 ;
	    RECT 1521.9000 518.4000 1524.6000 519.3000 ;
	    RECT 1521.9000 513.3000 1523.1000 518.4000 ;
	    RECT 1525.8000 513.3000 1527.0000 519.3000 ;
	    RECT 1557.0000 514.2000 1558.2001 519.3000 ;
	    RECT 1559.4000 515.1000 1560.6000 519.3000 ;
	    RECT 1561.8000 519.0000 1567.8000 519.3000 ;
	    RECT 1561.8000 514.2000 1563.0000 519.0000 ;
	    RECT 1557.0000 513.3000 1563.0000 514.2000 ;
	    RECT 1564.2001 513.3000 1565.4000 518.1000 ;
	    RECT 1566.6000 513.3000 1567.8000 519.0000 ;
	    RECT 1.2000 510.6000 1569.0000 512.4000 ;
	    RECT 126.6000 500.7000 127.8000 509.7000 ;
	    RECT 131.4000 503.7000 132.6000 509.7000 ;
	    RECT 136.2000 504.9000 137.4000 509.7000 ;
	    RECT 138.6000 505.5000 139.8000 509.7000 ;
	    RECT 141.0000 505.5000 142.2000 509.7000 ;
	    RECT 143.4000 505.5000 144.6000 509.7000 ;
	    RECT 145.8000 506.7000 147.0000 509.7000 ;
	    RECT 148.2000 505.5000 149.4000 509.7000 ;
	    RECT 150.6000 506.7000 151.8000 509.7000 ;
	    RECT 153.0000 505.5000 154.2000 509.7000 ;
	    RECT 155.4000 505.5000 156.6000 509.7000 ;
	    RECT 157.8000 505.5000 159.0000 509.7000 ;
	    RECT 160.2000 505.5000 161.4000 509.7000 ;
	    RECT 133.5000 503.7000 137.4000 504.9000 ;
	    RECT 162.6000 504.9000 163.8000 509.7000 ;
	    RECT 142.5000 503.7000 149.4000 504.6000 ;
	    RECT 133.5000 502.8000 134.7000 503.7000 ;
	    RECT 130.2000 501.6000 134.7000 502.8000 ;
	    RECT 126.6000 499.5000 139.8000 500.7000 ;
	    RECT 142.5000 500.1000 143.7000 503.7000 ;
	    RECT 148.2000 503.4000 149.4000 503.7000 ;
	    RECT 150.6000 503.4000 151.8000 504.6000 ;
	    RECT 152.7000 503.4000 153.0000 504.6000 ;
	    RECT 157.5000 503.4000 159.0000 504.6000 ;
	    RECT 162.6000 503.7000 166.2000 504.9000 ;
	    RECT 167.4000 503.7000 168.6000 509.7000 ;
	    RECT 145.8000 502.5000 147.0000 502.8000 ;
	    RECT 148.2000 502.2000 149.4000 502.5000 ;
	    RECT 145.8000 500.4000 147.0000 501.6000 ;
	    RECT 148.2000 501.3000 154.8000 502.2000 ;
	    RECT 153.6000 501.0000 154.8000 501.3000 ;
	    RECT 13.8000 492.4500 15.0000 492.6000 ;
	    RECT 117.0000 492.4500 118.2000 492.6000 ;
	    RECT 13.8000 491.5500 118.2000 492.4500 ;
	    RECT 13.8000 491.4000 15.0000 491.5500 ;
	    RECT 117.0000 491.4000 118.2000 491.5500 ;
	    RECT 126.6000 491.1000 127.8000 499.5000 ;
	    RECT 140.7000 498.9000 143.7000 500.1000 ;
	    RECT 149.4000 498.9000 154.2000 500.1000 ;
	    RECT 157.8000 499.2000 159.0000 503.4000 ;
	    RECT 165.0000 502.8000 166.2000 503.7000 ;
	    RECT 165.0000 501.9000 167.7000 502.8000 ;
	    RECT 166.5000 500.1000 167.7000 501.9000 ;
	    RECT 172.2000 501.9000 173.4000 509.7000 ;
	    RECT 174.6000 504.0000 175.8000 509.7000 ;
	    RECT 177.0000 506.7000 178.2000 509.7000 ;
	    RECT 191.4000 506.7000 192.6000 509.7000 ;
	    RECT 191.4000 505.5000 192.6000 505.8000 ;
	    RECT 184.2000 504.4500 185.4000 504.6000 ;
	    RECT 191.4000 504.4500 192.6000 504.6000 ;
	    RECT 174.6000 502.8000 176.1000 504.0000 ;
	    RECT 184.2000 503.5500 192.6000 504.4500 ;
	    RECT 184.2000 503.4000 185.4000 503.5500 ;
	    RECT 191.4000 503.4000 192.6000 503.5500 ;
	    RECT 172.2000 501.0000 174.0000 501.9000 ;
	    RECT 166.5000 498.9000 172.2000 500.1000 ;
	    RECT 128.7000 498.0000 129.9000 498.3000 ;
	    RECT 128.7000 497.1000 135.3000 498.0000 ;
	    RECT 136.2000 497.4000 137.4000 498.6000 ;
	    RECT 162.6000 498.0000 163.8000 498.9000 ;
	    RECT 173.1000 498.0000 174.0000 501.0000 ;
	    RECT 138.3000 497.1000 163.8000 498.0000 ;
	    RECT 172.8000 497.1000 174.0000 498.0000 ;
	    RECT 170.7000 496.2000 171.9000 496.5000 ;
	    RECT 131.4000 494.4000 132.6000 495.6000 ;
	    RECT 133.5000 495.3000 171.9000 496.2000 ;
	    RECT 136.5000 495.0000 137.7000 495.3000 ;
	    RECT 172.8000 494.4000 173.7000 497.1000 ;
	    RECT 174.9000 496.2000 176.1000 502.8000 ;
	    RECT 193.8000 502.5000 195.0000 509.7000 ;
	    RECT 215.4000 506.7000 216.6000 509.7000 ;
	    RECT 215.4000 505.5000 216.6000 505.8000 ;
	    RECT 215.4000 503.4000 216.6000 504.6000 ;
	    RECT 217.8000 502.5000 219.0000 509.7000 ;
	    RECT 229.8000 506.7000 231.0000 509.7000 ;
	    RECT 229.8000 505.5000 231.0000 505.8000 ;
	    RECT 227.4000 504.4500 228.6000 504.6000 ;
	    RECT 229.8000 504.4500 231.0000 504.6000 ;
	    RECT 227.4000 503.5500 231.0000 504.4500 ;
	    RECT 227.4000 503.4000 228.6000 503.5500 ;
	    RECT 229.8000 503.4000 231.0000 503.5500 ;
	    RECT 232.2000 502.5000 233.4000 509.7000 ;
	    RECT 263.4000 504.0000 264.6000 509.7000 ;
	    RECT 265.8000 504.9000 267.0000 509.7000 ;
	    RECT 268.2000 508.8000 274.2000 509.7000 ;
	    RECT 268.2000 504.0000 269.4000 508.8000 ;
	    RECT 263.4000 503.7000 269.4000 504.0000 ;
	    RECT 270.6000 503.7000 271.8000 507.9000 ;
	    RECT 273.0000 503.7000 274.2000 508.8000 ;
	    RECT 297.0000 504.0000 298.2000 509.7000 ;
	    RECT 299.4000 504.9000 300.6000 509.7000 ;
	    RECT 301.8000 504.0000 303.0000 509.7000 ;
	    RECT 297.0000 503.7000 303.0000 504.0000 ;
	    RECT 304.2000 503.7000 305.4000 509.7000 ;
	    RECT 263.7000 503.1000 269.1000 503.7000 ;
	    RECT 193.8000 501.4500 195.0000 501.6000 ;
	    RECT 213.0000 501.4500 214.2000 501.6000 ;
	    RECT 193.8000 500.5500 214.2000 501.4500 ;
	    RECT 193.8000 500.4000 195.0000 500.5500 ;
	    RECT 213.0000 500.4000 214.2000 500.5500 ;
	    RECT 217.8000 501.4500 219.0000 501.6000 ;
	    RECT 229.8000 501.4500 231.0000 501.6000 ;
	    RECT 217.8000 500.5500 231.0000 501.4500 ;
	    RECT 217.8000 500.4000 219.0000 500.5500 ;
	    RECT 229.8000 500.4000 231.0000 500.5500 ;
	    RECT 232.2000 501.4500 233.4000 501.6000 ;
	    RECT 263.4000 501.4500 264.6000 501.6000 ;
	    RECT 232.2000 500.5500 264.6000 501.4500 ;
	    RECT 265.5000 500.7000 265.8000 502.2000 ;
	    RECT 270.9000 501.6000 271.8000 503.7000 ;
	    RECT 297.3000 503.1000 302.7000 503.7000 ;
	    RECT 304.2000 502.5000 305.1000 503.7000 ;
	    RECT 318.6000 502.5000 319.8000 509.7000 ;
	    RECT 321.0000 506.7000 322.2000 509.7000 ;
	    RECT 321.0000 505.5000 322.2000 505.8000 ;
	    RECT 321.0000 504.4500 322.2000 504.6000 ;
	    RECT 333.0000 504.4500 334.2000 504.6000 ;
	    RECT 321.0000 503.5500 334.2000 504.4500 ;
	    RECT 321.0000 503.4000 322.2000 503.5500 ;
	    RECT 333.0000 503.4000 334.2000 503.5500 ;
	    RECT 335.4000 502.5000 336.6000 509.7000 ;
	    RECT 337.8000 506.7000 339.0000 509.7000 ;
	    RECT 354.6000 507.4500 355.8000 507.6000 ;
	    RECT 445.8000 507.4500 447.0000 507.6000 ;
	    RECT 354.6000 506.5500 447.0000 507.4500 ;
	    RECT 469.8000 506.7000 471.0000 509.7000 ;
	    RECT 354.6000 506.4000 355.8000 506.5500 ;
	    RECT 445.8000 506.4000 447.0000 506.5500 ;
	    RECT 337.8000 505.5000 339.0000 505.8000 ;
	    RECT 337.8000 503.4000 339.0000 504.6000 ;
	    RECT 472.2000 504.0000 473.4000 509.7000 ;
	    RECT 471.9000 502.8000 473.4000 504.0000 ;
	    RECT 232.2000 500.4000 233.4000 500.5500 ;
	    RECT 263.4000 500.4000 264.6000 500.5500 ;
	    RECT 268.2000 500.4000 269.4000 501.6000 ;
	    RECT 270.3000 500.7000 271.8000 501.6000 ;
	    RECT 273.0000 500.4000 274.2000 501.6000 ;
	    RECT 297.0000 500.4000 298.2000 501.6000 ;
	    RECT 299.1000 500.7000 299.4000 502.2000 ;
	    RECT 301.5000 500.4000 303.3000 501.6000 ;
	    RECT 304.2000 501.4500 305.4000 501.6000 ;
	    RECT 306.6000 501.4500 307.8000 501.6000 ;
	    RECT 304.2000 500.5500 307.8000 501.4500 ;
	    RECT 304.2000 500.4000 305.4000 500.5500 ;
	    RECT 306.6000 500.4000 307.8000 500.5500 ;
	    RECT 309.0000 501.4500 310.2000 501.6000 ;
	    RECT 318.6000 501.4500 319.8000 501.6000 ;
	    RECT 309.0000 500.5500 319.8000 501.4500 ;
	    RECT 309.0000 500.4000 310.2000 500.5500 ;
	    RECT 318.6000 500.4000 319.8000 500.5500 ;
	    RECT 330.6000 501.4500 331.8000 501.6000 ;
	    RECT 335.4000 501.4500 336.6000 501.6000 ;
	    RECT 330.6000 500.5500 336.6000 501.4500 ;
	    RECT 330.6000 500.4000 331.8000 500.5500 ;
	    RECT 335.4000 500.4000 336.6000 500.5500 ;
	    RECT 345.0000 501.4500 346.2000 501.6000 ;
	    RECT 455.4000 501.4500 456.6000 501.6000 ;
	    RECT 345.0000 500.5500 456.6000 501.4500 ;
	    RECT 345.0000 500.4000 346.2000 500.5500 ;
	    RECT 455.4000 500.4000 456.6000 500.5500 ;
	    RECT 265.8000 499.5000 267.0000 499.8000 ;
	    RECT 270.6000 499.5000 271.8000 499.8000 ;
	    RECT 299.4000 499.5000 300.6000 499.8000 ;
	    RECT 141.0000 494.1000 142.2000 494.4000 ;
	    RECT 134.1000 493.5000 142.2000 494.1000 ;
	    RECT 132.9000 493.2000 142.2000 493.5000 ;
	    RECT 143.7000 493.5000 156.6000 494.4000 ;
	    RECT 129.0000 492.0000 131.4000 493.2000 ;
	    RECT 132.9000 492.3000 135.0000 493.2000 ;
	    RECT 143.7000 492.3000 144.6000 493.5000 ;
	    RECT 155.4000 493.2000 156.6000 493.5000 ;
	    RECT 160.2000 493.5000 173.7000 494.4000 ;
	    RECT 174.6000 495.0000 176.1000 496.2000 ;
	    RECT 174.6000 493.5000 175.8000 495.0000 ;
	    RECT 160.2000 493.2000 161.4000 493.5000 ;
	    RECT 130.5000 491.4000 131.4000 492.0000 ;
	    RECT 135.9000 491.4000 144.6000 492.3000 ;
	    RECT 145.5000 491.4000 149.4000 492.6000 ;
	    RECT 126.6000 490.2000 129.6000 491.1000 ;
	    RECT 130.5000 490.2000 136.8000 491.4000 ;
	    RECT 128.7000 489.3000 129.6000 490.2000 ;
	    RECT 126.6000 483.3000 127.8000 489.3000 ;
	    RECT 128.7000 488.4000 130.2000 489.3000 ;
	    RECT 129.0000 483.3000 130.2000 488.4000 ;
	    RECT 131.4000 482.4000 132.6000 489.3000 ;
	    RECT 133.8000 483.3000 135.0000 490.2000 ;
	    RECT 136.2000 483.3000 137.4000 489.3000 ;
	    RECT 138.6000 483.3000 139.8000 487.5000 ;
	    RECT 141.0000 483.3000 142.2000 487.5000 ;
	    RECT 143.4000 483.3000 144.6000 490.5000 ;
	    RECT 145.8000 483.3000 147.0000 489.3000 ;
	    RECT 148.2000 483.3000 149.4000 490.5000 ;
	    RECT 150.6000 483.3000 151.8000 489.3000 ;
	    RECT 153.0000 483.3000 154.2000 492.6000 ;
	    RECT 165.0000 491.4000 168.9000 492.6000 ;
	    RECT 157.8000 490.2000 164.1000 491.4000 ;
	    RECT 155.4000 483.3000 156.6000 487.5000 ;
	    RECT 157.8000 483.3000 159.0000 487.5000 ;
	    RECT 160.2000 483.3000 161.4000 487.5000 ;
	    RECT 162.6000 483.3000 163.8000 489.3000 ;
	    RECT 165.0000 483.3000 166.2000 491.4000 ;
	    RECT 172.8000 491.1000 173.7000 493.5000 ;
	    RECT 174.6000 491.4000 175.8000 492.6000 ;
	    RECT 169.8000 490.2000 173.7000 491.1000 ;
	    RECT 167.4000 483.3000 168.6000 489.3000 ;
	    RECT 169.8000 483.3000 171.0000 490.2000 ;
	    RECT 172.2000 483.3000 173.4000 489.3000 ;
	    RECT 174.6000 483.3000 175.8000 490.5000 ;
	    RECT 177.0000 483.3000 178.2000 489.3000 ;
	    RECT 191.4000 483.3000 192.6000 489.3000 ;
	    RECT 193.8000 483.3000 195.0000 499.5000 ;
	    RECT 215.4000 483.3000 216.6000 489.3000 ;
	    RECT 217.8000 483.3000 219.0000 499.5000 ;
	    RECT 229.8000 483.3000 231.0000 489.3000 ;
	    RECT 232.2000 483.3000 233.4000 499.5000 ;
	    RECT 251.4000 498.4500 252.6000 498.6000 ;
	    RECT 265.8000 498.4500 267.0000 498.6000 ;
	    RECT 251.4000 497.5500 267.0000 498.4500 ;
	    RECT 251.4000 497.4000 252.6000 497.5500 ;
	    RECT 265.8000 497.4000 267.0000 497.5500 ;
	    RECT 268.2000 495.3000 269.1000 499.5000 ;
	    RECT 273.0000 499.2000 274.2000 499.5000 ;
	    RECT 270.6000 497.4000 271.8000 498.6000 ;
	    RECT 299.4000 497.4000 300.6000 498.6000 ;
	    RECT 301.5000 495.3000 302.4000 500.4000 ;
	    RECT 263.4000 483.3000 264.6000 495.3000 ;
	    RECT 267.3000 483.3000 270.3000 495.3000 ;
	    RECT 273.0000 483.3000 274.2000 495.3000 ;
	    RECT 297.0000 483.3000 298.2000 495.3000 ;
	    RECT 300.9000 494.4000 302.4000 495.3000 ;
	    RECT 304.2000 494.4000 305.4000 495.6000 ;
	    RECT 300.9000 483.3000 302.1000 494.4000 ;
	    RECT 303.3000 492.6000 304.2000 493.5000 ;
	    RECT 303.0000 491.4000 304.2000 492.6000 ;
	    RECT 303.3000 483.3000 304.5000 489.3000 ;
	    RECT 318.6000 483.3000 319.8000 499.5000 ;
	    RECT 321.0000 483.3000 322.2000 489.3000 ;
	    RECT 335.4000 483.3000 336.6000 499.5000 ;
	    RECT 471.9000 496.2000 473.1000 502.8000 ;
	    RECT 474.6000 501.9000 475.8000 509.7000 ;
	    RECT 479.4000 503.7000 480.6000 509.7000 ;
	    RECT 484.2000 504.9000 485.4000 509.7000 ;
	    RECT 486.6000 505.5000 487.8000 509.7000 ;
	    RECT 489.0000 505.5000 490.2000 509.7000 ;
	    RECT 491.4000 505.5000 492.6000 509.7000 ;
	    RECT 493.8000 505.5000 495.0000 509.7000 ;
	    RECT 496.2000 506.7000 497.4000 509.7000 ;
	    RECT 498.6000 505.5000 499.8000 509.7000 ;
	    RECT 501.0000 506.7000 502.2000 509.7000 ;
	    RECT 503.4000 505.5000 504.6000 509.7000 ;
	    RECT 505.8000 505.5000 507.0000 509.7000 ;
	    RECT 508.2000 505.5000 509.4000 509.7000 ;
	    RECT 481.8000 503.7000 485.4000 504.9000 ;
	    RECT 510.6000 504.9000 511.8000 509.7000 ;
	    RECT 481.8000 502.8000 483.0000 503.7000 ;
	    RECT 474.0000 501.0000 475.8000 501.9000 ;
	    RECT 480.3000 501.9000 483.0000 502.8000 ;
	    RECT 489.0000 503.4000 490.5000 504.6000 ;
	    RECT 495.0000 503.4000 495.3000 504.6000 ;
	    RECT 496.2000 503.4000 497.4000 504.6000 ;
	    RECT 498.6000 503.7000 505.5000 504.6000 ;
	    RECT 510.6000 503.7000 514.5000 504.9000 ;
	    RECT 515.4000 503.7000 516.6000 509.7000 ;
	    RECT 498.6000 503.4000 499.8000 503.7000 ;
	    RECT 474.0000 498.0000 474.9000 501.0000 ;
	    RECT 480.3000 500.1000 481.5000 501.9000 ;
	    RECT 475.8000 498.9000 481.5000 500.1000 ;
	    RECT 489.0000 499.2000 490.2000 503.4000 ;
	    RECT 501.0000 502.5000 502.2000 502.8000 ;
	    RECT 498.6000 502.2000 499.8000 502.5000 ;
	    RECT 493.2000 501.3000 499.8000 502.2000 ;
	    RECT 493.2000 501.0000 494.4000 501.3000 ;
	    RECT 501.0000 500.4000 502.2000 501.6000 ;
	    RECT 504.3000 500.1000 505.5000 503.7000 ;
	    RECT 513.3000 502.8000 514.5000 503.7000 ;
	    RECT 513.3000 501.6000 517.8000 502.8000 ;
	    RECT 520.2000 500.7000 521.4000 509.7000 ;
	    RECT 539.4000 502.5000 540.6000 509.7000 ;
	    RECT 541.8000 503.7000 543.0000 509.7000 ;
	    RECT 544.2000 502.8000 545.4000 509.7000 ;
	    RECT 570.6000 503.7000 571.8000 509.7000 ;
	    RECT 573.0000 504.0000 574.2000 509.7000 ;
	    RECT 575.4000 504.9000 576.6000 509.7000 ;
	    RECT 577.8000 504.0000 579.0000 509.7000 ;
	    RECT 573.0000 503.7000 579.0000 504.0000 ;
	    RECT 542.1000 501.9000 545.4000 502.8000 ;
	    RECT 570.9000 502.5000 571.8000 503.7000 ;
	    RECT 573.3000 503.1000 578.7000 503.7000 ;
	    RECT 597.0000 502.8000 598.2000 509.7000 ;
	    RECT 599.4000 503.7000 600.6000 509.7000 ;
	    RECT 493.8000 498.9000 498.6000 500.1000 ;
	    RECT 504.3000 498.9000 507.3000 500.1000 ;
	    RECT 508.2000 499.5000 521.4000 500.7000 ;
	    RECT 539.4000 500.4000 540.6000 501.6000 ;
	    RECT 484.2000 498.0000 485.4000 498.9000 ;
	    RECT 474.0000 497.1000 475.2000 498.0000 ;
	    RECT 484.2000 497.1000 509.7000 498.0000 ;
	    RECT 510.6000 497.4000 511.8000 498.6000 ;
	    RECT 518.1000 498.0000 519.3000 498.3000 ;
	    RECT 512.7000 497.1000 519.3000 498.0000 ;
	    RECT 347.4000 495.4500 348.6000 495.6000 ;
	    RECT 359.4000 495.4500 360.6000 495.6000 ;
	    RECT 347.4000 494.5500 360.6000 495.4500 ;
	    RECT 471.9000 495.0000 473.4000 496.2000 ;
	    RECT 347.4000 494.4000 348.6000 494.5500 ;
	    RECT 359.4000 494.4000 360.6000 494.5500 ;
	    RECT 472.2000 493.5000 473.4000 495.0000 ;
	    RECT 474.3000 494.4000 475.2000 497.1000 ;
	    RECT 476.1000 496.2000 477.3000 496.5000 ;
	    RECT 476.1000 495.3000 514.5000 496.2000 ;
	    RECT 510.3000 495.0000 511.5000 495.3000 ;
	    RECT 515.4000 494.4000 516.6000 495.6000 ;
	    RECT 474.3000 493.5000 487.8000 494.4000 ;
	    RECT 373.8000 492.4500 375.0000 492.6000 ;
	    RECT 409.8000 492.4500 411.0000 492.6000 ;
	    RECT 472.2000 492.4500 473.4000 492.6000 ;
	    RECT 373.8000 491.5500 473.4000 492.4500 ;
	    RECT 373.8000 491.4000 375.0000 491.5500 ;
	    RECT 409.8000 491.4000 411.0000 491.5500 ;
	    RECT 472.2000 491.4000 473.4000 491.5500 ;
	    RECT 474.3000 491.1000 475.2000 493.5000 ;
	    RECT 486.6000 493.2000 487.8000 493.5000 ;
	    RECT 491.4000 493.5000 504.3000 494.4000 ;
	    RECT 491.4000 493.2000 492.6000 493.5000 ;
	    RECT 479.1000 491.4000 483.0000 492.6000 ;
	    RECT 337.8000 483.3000 339.0000 489.3000 ;
	    RECT 469.8000 483.3000 471.0000 489.3000 ;
	    RECT 472.2000 483.3000 473.4000 490.5000 ;
	    RECT 474.3000 490.2000 478.2000 491.1000 ;
	    RECT 474.6000 483.3000 475.8000 489.3000 ;
	    RECT 477.0000 483.3000 478.2000 490.2000 ;
	    RECT 479.4000 483.3000 480.6000 489.3000 ;
	    RECT 481.8000 483.3000 483.0000 491.4000 ;
	    RECT 483.9000 490.2000 490.2000 491.4000 ;
	    RECT 484.2000 483.3000 485.4000 489.3000 ;
	    RECT 486.6000 483.3000 487.8000 487.5000 ;
	    RECT 489.0000 483.3000 490.2000 487.5000 ;
	    RECT 491.4000 483.3000 492.6000 487.5000 ;
	    RECT 493.8000 483.3000 495.0000 492.6000 ;
	    RECT 498.6000 491.4000 502.5000 492.6000 ;
	    RECT 503.4000 492.3000 504.3000 493.5000 ;
	    RECT 505.8000 494.1000 507.0000 494.4000 ;
	    RECT 505.8000 493.5000 513.9000 494.1000 ;
	    RECT 505.8000 493.2000 515.1000 493.5000 ;
	    RECT 513.0000 492.3000 515.1000 493.2000 ;
	    RECT 503.4000 491.4000 512.1000 492.3000 ;
	    RECT 516.6000 492.0000 519.0000 493.2000 ;
	    RECT 516.6000 491.4000 517.5000 492.0000 ;
	    RECT 496.2000 483.3000 497.4000 489.3000 ;
	    RECT 498.6000 483.3000 499.8000 490.5000 ;
	    RECT 501.0000 483.3000 502.2000 489.3000 ;
	    RECT 503.4000 483.3000 504.6000 490.5000 ;
	    RECT 511.2000 490.2000 517.5000 491.4000 ;
	    RECT 520.2000 491.1000 521.4000 499.5000 ;
	    RECT 518.4000 490.2000 521.4000 491.1000 ;
	    RECT 539.4000 498.6000 540.6000 499.5000 ;
	    RECT 539.4000 495.3000 540.3000 498.6000 ;
	    RECT 542.1000 497.4000 543.0000 501.9000 ;
	    RECT 568.2000 501.4500 569.4000 501.6000 ;
	    RECT 570.6000 501.4500 571.8000 501.6000 ;
	    RECT 568.2000 500.5500 571.8000 501.4500 ;
	    RECT 568.2000 500.4000 569.4000 500.5500 ;
	    RECT 570.6000 500.4000 571.8000 500.5500 ;
	    RECT 572.7000 500.4000 574.5000 501.6000 ;
	    RECT 576.6000 500.7000 576.9000 502.2000 ;
	    RECT 597.0000 501.9000 600.3000 502.8000 ;
	    RECT 601.8000 502.5000 603.0000 509.7000 ;
	    RECT 613.8000 502.5000 615.0000 509.7000 ;
	    RECT 616.2000 506.7000 617.4000 509.7000 ;
	    RECT 635.4000 506.7000 636.6000 509.7000 ;
	    RECT 637.8000 506.7000 639.0000 509.7000 ;
	    RECT 640.2000 506.7000 641.4000 509.7000 ;
	    RECT 772.2000 506.7000 773.4000 509.7000 ;
	    RECT 616.2000 505.5000 617.4000 505.8000 ;
	    RECT 616.2000 503.4000 617.4000 504.6000 ;
	    RECT 637.8000 502.5000 638.7000 506.7000 ;
	    RECT 640.2000 505.5000 641.4000 505.8000 ;
	    RECT 640.2000 504.4500 641.4000 504.6000 ;
	    RECT 647.4000 504.4500 648.6000 504.6000 ;
	    RECT 640.2000 503.5500 648.6000 504.4500 ;
	    RECT 774.6000 504.0000 775.8000 509.7000 ;
	    RECT 640.2000 503.4000 641.4000 503.5500 ;
	    RECT 647.4000 503.4000 648.6000 503.5500 ;
	    RECT 774.3000 502.8000 775.8000 504.0000 ;
	    RECT 577.8000 500.4000 579.0000 501.6000 ;
	    RECT 544.2000 499.5000 545.4000 499.8000 ;
	    RECT 541.2000 496.2000 543.0000 497.4000 ;
	    RECT 542.1000 495.3000 543.0000 496.2000 ;
	    RECT 505.8000 483.3000 507.0000 487.5000 ;
	    RECT 508.2000 483.3000 509.4000 487.5000 ;
	    RECT 510.6000 483.3000 511.8000 489.3000 ;
	    RECT 513.0000 483.3000 514.2000 490.2000 ;
	    RECT 518.4000 489.3000 519.3000 490.2000 ;
	    RECT 515.4000 482.4000 516.6000 489.3000 ;
	    RECT 517.8000 488.4000 519.3000 489.3000 ;
	    RECT 517.8000 483.3000 519.0000 488.4000 ;
	    RECT 520.2000 483.3000 521.4000 489.3000 ;
	    RECT 539.4000 483.3000 540.6000 495.3000 ;
	    RECT 542.1000 494.4000 545.4000 495.3000 ;
	    RECT 570.6000 494.4000 571.8000 495.6000 ;
	    RECT 573.6000 495.3000 574.5000 500.4000 ;
	    RECT 575.4000 499.5000 576.6000 499.8000 ;
	    RECT 597.0000 499.5000 598.2000 499.8000 ;
	    RECT 575.4000 497.4000 576.6000 498.6000 ;
	    RECT 599.4000 497.4000 600.3000 501.9000 ;
	    RECT 601.8000 501.4500 603.0000 501.6000 ;
	    RECT 611.4000 501.4500 612.6000 501.6000 ;
	    RECT 601.8000 500.5500 612.6000 501.4500 ;
	    RECT 601.8000 500.4000 603.0000 500.5500 ;
	    RECT 611.4000 500.4000 612.6000 500.5500 ;
	    RECT 613.8000 501.4500 615.0000 501.6000 ;
	    RECT 635.4000 501.4500 636.6000 501.6000 ;
	    RECT 613.8000 500.5500 636.6000 501.4500 ;
	    RECT 613.8000 500.4000 615.0000 500.5500 ;
	    RECT 635.4000 500.4000 636.6000 500.5500 ;
	    RECT 637.8000 500.4000 639.0000 501.6000 ;
	    RECT 676.2000 501.4500 677.4000 501.6000 ;
	    RECT 681.0000 501.4500 682.2000 501.6000 ;
	    RECT 676.2000 500.5500 682.2000 501.4500 ;
	    RECT 676.2000 500.4000 677.4000 500.5500 ;
	    RECT 681.0000 500.4000 682.2000 500.5500 ;
	    RECT 601.8000 498.6000 603.0000 499.5000 ;
	    RECT 599.4000 496.2000 601.2000 497.4000 ;
	    RECT 599.4000 495.3000 600.3000 496.2000 ;
	    RECT 602.1000 495.3000 603.0000 498.6000 ;
	    RECT 573.6000 494.4000 575.1000 495.3000 ;
	    RECT 541.8000 483.3000 543.0000 493.5000 ;
	    RECT 544.2000 483.3000 545.4000 494.4000 ;
	    RECT 571.8000 492.6000 572.7000 493.5000 ;
	    RECT 571.8000 491.4000 573.0000 492.6000 ;
	    RECT 571.5000 483.3000 572.7000 489.3000 ;
	    RECT 573.9000 483.3000 575.1000 494.4000 ;
	    RECT 577.8000 483.3000 579.0000 495.3000 ;
	    RECT 597.0000 494.4000 600.3000 495.3000 ;
	    RECT 597.0000 483.3000 598.2000 494.4000 ;
	    RECT 599.4000 483.3000 600.6000 493.5000 ;
	    RECT 601.8000 483.3000 603.0000 495.3000 ;
	    RECT 613.8000 483.3000 615.0000 499.5000 ;
	    RECT 635.4000 497.4000 636.6000 498.6000 ;
	    RECT 635.4000 496.2000 636.6000 496.5000 ;
	    RECT 637.8000 495.3000 638.7000 499.5000 ;
	    RECT 774.3000 496.2000 775.5000 502.8000 ;
	    RECT 777.0000 501.9000 778.2000 509.7000 ;
	    RECT 781.8000 503.7000 783.0000 509.7000 ;
	    RECT 786.6000 504.9000 787.8000 509.7000 ;
	    RECT 789.0000 505.5000 790.2000 509.7000 ;
	    RECT 791.4000 505.5000 792.6000 509.7000 ;
	    RECT 793.8000 505.5000 795.0000 509.7000 ;
	    RECT 796.2000 505.5000 797.4000 509.7000 ;
	    RECT 798.6000 506.7000 799.8000 509.7000 ;
	    RECT 801.0000 505.5000 802.2000 509.7000 ;
	    RECT 803.4000 506.7000 804.6000 509.7000 ;
	    RECT 805.8000 505.5000 807.0000 509.7000 ;
	    RECT 808.2000 505.5000 809.4000 509.7000 ;
	    RECT 810.6000 505.5000 811.8000 509.7000 ;
	    RECT 784.2000 503.7000 787.8000 504.9000 ;
	    RECT 813.0000 504.9000 814.2000 509.7000 ;
	    RECT 784.2000 502.8000 785.4000 503.7000 ;
	    RECT 776.4000 501.0000 778.2000 501.9000 ;
	    RECT 782.7000 501.9000 785.4000 502.8000 ;
	    RECT 791.4000 503.4000 792.9000 504.6000 ;
	    RECT 797.4000 503.4000 797.7000 504.6000 ;
	    RECT 798.6000 503.4000 799.8000 504.6000 ;
	    RECT 801.0000 503.7000 807.9000 504.6000 ;
	    RECT 813.0000 503.7000 816.9000 504.9000 ;
	    RECT 817.8000 503.7000 819.0000 509.7000 ;
	    RECT 801.0000 503.4000 802.2000 503.7000 ;
	    RECT 776.4000 498.0000 777.3000 501.0000 ;
	    RECT 782.7000 500.1000 783.9000 501.9000 ;
	    RECT 778.2000 498.9000 783.9000 500.1000 ;
	    RECT 791.4000 499.2000 792.6000 503.4000 ;
	    RECT 803.4000 502.5000 804.6000 502.8000 ;
	    RECT 801.0000 502.2000 802.2000 502.5000 ;
	    RECT 795.6000 501.3000 802.2000 502.2000 ;
	    RECT 795.6000 501.0000 796.8000 501.3000 ;
	    RECT 803.4000 500.4000 804.6000 501.6000 ;
	    RECT 806.7000 500.1000 807.9000 503.7000 ;
	    RECT 815.7000 502.8000 816.9000 503.7000 ;
	    RECT 815.7000 501.6000 820.2000 502.8000 ;
	    RECT 822.6000 500.7000 823.8000 509.7000 ;
	    RECT 837.0000 502.5000 838.2000 509.7000 ;
	    RECT 839.4000 506.7000 840.6000 509.7000 ;
	    RECT 839.4000 505.5000 840.6000 505.8000 ;
	    RECT 839.4000 504.4500 840.6000 504.6000 ;
	    RECT 841.8000 504.4500 843.0000 504.6000 ;
	    RECT 839.4000 503.5500 843.0000 504.4500 ;
	    RECT 863.4000 503.7000 864.6000 509.7000 ;
	    RECT 865.8000 504.0000 867.0000 509.7000 ;
	    RECT 868.2000 504.9000 869.4000 509.7000 ;
	    RECT 870.6000 504.0000 871.8000 509.7000 ;
	    RECT 865.8000 503.7000 871.8000 504.0000 ;
	    RECT 889.8000 503.7000 891.0000 509.7000 ;
	    RECT 893.7000 504.6000 894.9000 509.7000 ;
	    RECT 892.2000 503.7000 894.9000 504.6000 ;
	    RECT 839.4000 503.4000 840.6000 503.5500 ;
	    RECT 841.8000 503.4000 843.0000 503.5500 ;
	    RECT 863.7000 502.5000 864.6000 503.7000 ;
	    RECT 866.1000 503.1000 871.5000 503.7000 ;
	    RECT 889.8000 502.5000 891.0000 502.8000 ;
	    RECT 796.2000 498.9000 801.0000 500.1000 ;
	    RECT 806.7000 498.9000 809.7000 500.1000 ;
	    RECT 810.6000 499.5000 823.8000 500.7000 ;
	    RECT 825.0000 501.4500 826.2000 501.6000 ;
	    RECT 837.0000 501.4500 838.2000 501.6000 ;
	    RECT 861.0000 501.4500 862.2000 501.6000 ;
	    RECT 825.0000 500.5500 862.2000 501.4500 ;
	    RECT 825.0000 500.4000 826.2000 500.5500 ;
	    RECT 837.0000 500.4000 838.2000 500.5500 ;
	    RECT 861.0000 500.4000 862.2000 500.5500 ;
	    RECT 863.4000 500.4000 864.6000 501.6000 ;
	    RECT 865.5000 500.4000 867.3000 501.6000 ;
	    RECT 869.4000 500.7000 869.7000 502.2000 ;
	    RECT 870.6000 500.4000 871.8000 501.6000 ;
	    RECT 889.8000 500.4000 891.0000 501.6000 ;
	    RECT 786.6000 498.0000 787.8000 498.9000 ;
	    RECT 776.4000 497.1000 777.6000 498.0000 ;
	    RECT 786.6000 497.1000 812.1000 498.0000 ;
	    RECT 813.0000 497.4000 814.2000 498.6000 ;
	    RECT 820.5000 498.0000 821.7000 498.3000 ;
	    RECT 815.1000 497.1000 821.7000 498.0000 ;
	    RECT 636.3000 494.1000 639.0000 495.3000 ;
	    RECT 616.2000 483.3000 617.4000 489.3000 ;
	    RECT 636.3000 483.3000 637.5000 494.1000 ;
	    RECT 640.2000 483.3000 641.4000 495.3000 ;
	    RECT 774.3000 495.0000 775.8000 496.2000 ;
	    RECT 774.6000 493.5000 775.8000 495.0000 ;
	    RECT 776.7000 494.4000 777.6000 497.1000 ;
	    RECT 778.5000 496.2000 779.7000 496.5000 ;
	    RECT 778.5000 495.3000 816.9000 496.2000 ;
	    RECT 812.7000 495.0000 813.9000 495.3000 ;
	    RECT 817.8000 494.4000 819.0000 495.6000 ;
	    RECT 776.7000 493.5000 790.2000 494.4000 ;
	    RECT 712.2000 492.4500 713.4000 492.6000 ;
	    RECT 774.6000 492.4500 775.8000 492.6000 ;
	    RECT 712.2000 491.5500 775.8000 492.4500 ;
	    RECT 712.2000 491.4000 713.4000 491.5500 ;
	    RECT 774.6000 491.4000 775.8000 491.5500 ;
	    RECT 776.7000 491.1000 777.6000 493.5000 ;
	    RECT 789.0000 493.2000 790.2000 493.5000 ;
	    RECT 793.8000 493.5000 806.7000 494.4000 ;
	    RECT 793.8000 493.2000 795.0000 493.5000 ;
	    RECT 781.5000 491.4000 785.4000 492.6000 ;
	    RECT 772.2000 483.3000 773.4000 489.3000 ;
	    RECT 774.6000 483.3000 775.8000 490.5000 ;
	    RECT 776.7000 490.2000 780.6000 491.1000 ;
	    RECT 777.0000 483.3000 778.2000 489.3000 ;
	    RECT 779.4000 483.3000 780.6000 490.2000 ;
	    RECT 781.8000 483.3000 783.0000 489.3000 ;
	    RECT 784.2000 483.3000 785.4000 491.4000 ;
	    RECT 786.3000 490.2000 792.6000 491.4000 ;
	    RECT 786.6000 483.3000 787.8000 489.3000 ;
	    RECT 789.0000 483.3000 790.2000 487.5000 ;
	    RECT 791.4000 483.3000 792.6000 487.5000 ;
	    RECT 793.8000 483.3000 795.0000 487.5000 ;
	    RECT 796.2000 483.3000 797.4000 492.6000 ;
	    RECT 801.0000 491.4000 804.9000 492.6000 ;
	    RECT 805.8000 492.3000 806.7000 493.5000 ;
	    RECT 808.2000 494.1000 809.4000 494.4000 ;
	    RECT 808.2000 493.5000 816.3000 494.1000 ;
	    RECT 808.2000 493.2000 817.5000 493.5000 ;
	    RECT 815.4000 492.3000 817.5000 493.2000 ;
	    RECT 805.8000 491.4000 814.5000 492.3000 ;
	    RECT 819.0000 492.0000 821.4000 493.2000 ;
	    RECT 819.0000 491.4000 819.9000 492.0000 ;
	    RECT 798.6000 483.3000 799.8000 489.3000 ;
	    RECT 801.0000 483.3000 802.2000 490.5000 ;
	    RECT 803.4000 483.3000 804.6000 489.3000 ;
	    RECT 805.8000 483.3000 807.0000 490.5000 ;
	    RECT 813.6000 490.2000 819.9000 491.4000 ;
	    RECT 822.6000 491.1000 823.8000 499.5000 ;
	    RECT 820.8000 490.2000 823.8000 491.1000 ;
	    RECT 808.2000 483.3000 809.4000 487.5000 ;
	    RECT 810.6000 483.3000 811.8000 487.5000 ;
	    RECT 813.0000 483.3000 814.2000 489.3000 ;
	    RECT 815.4000 483.3000 816.6000 490.2000 ;
	    RECT 820.8000 489.3000 821.7000 490.2000 ;
	    RECT 817.8000 482.4000 819.0000 489.3000 ;
	    RECT 820.2000 488.4000 821.7000 489.3000 ;
	    RECT 820.2000 483.3000 821.4000 488.4000 ;
	    RECT 822.6000 483.3000 823.8000 489.3000 ;
	    RECT 837.0000 483.3000 838.2000 499.5000 ;
	    RECT 863.4000 494.4000 864.6000 495.6000 ;
	    RECT 866.4000 495.3000 867.3000 500.4000 ;
	    RECT 868.2000 499.5000 869.4000 499.8000 ;
	    RECT 892.2000 499.5000 893.4000 503.7000 ;
	    RECT 1026.6000 500.7000 1027.8000 509.7000 ;
	    RECT 1031.4000 503.7000 1032.6000 509.7000 ;
	    RECT 1036.2001 504.9000 1037.4000 509.7000 ;
	    RECT 1038.6000 505.5000 1039.8000 509.7000 ;
	    RECT 1041.0000 505.5000 1042.2001 509.7000 ;
	    RECT 1043.4000 505.5000 1044.6000 509.7000 ;
	    RECT 1045.8000 506.7000 1047.0000 509.7000 ;
	    RECT 1048.2001 505.5000 1049.4000 509.7000 ;
	    RECT 1050.6000 506.7000 1051.8000 509.7000 ;
	    RECT 1053.0000 505.5000 1054.2001 509.7000 ;
	    RECT 1055.4000 505.5000 1056.6000 509.7000 ;
	    RECT 1057.8000 505.5000 1059.0000 509.7000 ;
	    RECT 1060.2001 505.5000 1061.4000 509.7000 ;
	    RECT 1033.5000 503.7000 1037.4000 504.9000 ;
	    RECT 1062.6000 504.9000 1063.8000 509.7000 ;
	    RECT 1042.5000 503.7000 1049.4000 504.6000 ;
	    RECT 1033.5000 502.8000 1034.7001 503.7000 ;
	    RECT 1030.2001 501.6000 1034.7001 502.8000 ;
	    RECT 1026.6000 499.5000 1039.8000 500.7000 ;
	    RECT 1042.5000 500.1000 1043.7001 503.7000 ;
	    RECT 1048.2001 503.4000 1049.4000 503.7000 ;
	    RECT 1050.6000 503.4000 1051.8000 504.6000 ;
	    RECT 1052.7001 503.4000 1053.0000 504.6000 ;
	    RECT 1057.5000 503.4000 1059.0000 504.6000 ;
	    RECT 1062.6000 503.7000 1066.2001 504.9000 ;
	    RECT 1067.4000 503.7000 1068.6000 509.7000 ;
	    RECT 1045.8000 502.5000 1047.0000 502.8000 ;
	    RECT 1048.2001 502.2000 1049.4000 502.5000 ;
	    RECT 1045.8000 500.4000 1047.0000 501.6000 ;
	    RECT 1048.2001 501.3000 1054.8000 502.2000 ;
	    RECT 1053.6000 501.0000 1054.8000 501.3000 ;
	    RECT 868.2000 497.4000 869.4000 498.6000 ;
	    RECT 870.6000 498.4500 871.8000 498.6000 ;
	    RECT 892.2000 498.4500 893.4000 498.6000 ;
	    RECT 870.6000 497.5500 893.4000 498.4500 ;
	    RECT 870.6000 497.4000 871.8000 497.5500 ;
	    RECT 892.2000 497.4000 893.4000 497.5500 ;
	    RECT 866.4000 494.4000 867.9000 495.3000 ;
	    RECT 864.6000 492.6000 865.5000 493.5000 ;
	    RECT 864.6000 491.4000 865.8000 492.6000 ;
	    RECT 839.4000 483.3000 840.6000 489.3000 ;
	    RECT 864.3000 483.3000 865.5000 489.3000 ;
	    RECT 866.7000 483.3000 867.9000 494.4000 ;
	    RECT 870.6000 483.3000 871.8000 495.3000 ;
	    RECT 889.8000 483.3000 891.0000 489.3000 ;
	    RECT 892.2000 483.3000 893.4000 496.5000 ;
	    RECT 894.6000 495.4500 895.8000 495.6000 ;
	    RECT 906.6000 495.4500 907.8000 495.6000 ;
	    RECT 928.2000 495.4500 929.4000 495.6000 ;
	    RECT 894.6000 494.5500 929.4000 495.4500 ;
	    RECT 894.6000 494.4000 895.8000 494.5500 ;
	    RECT 906.6000 494.4000 907.8000 494.5500 ;
	    RECT 928.2000 494.4000 929.4000 494.5500 ;
	    RECT 894.6000 493.2000 895.8000 493.5000 ;
	    RECT 1026.6000 491.1000 1027.8000 499.5000 ;
	    RECT 1040.7001 498.9000 1043.7001 500.1000 ;
	    RECT 1049.4000 498.9000 1054.2001 500.1000 ;
	    RECT 1057.8000 499.2000 1059.0000 503.4000 ;
	    RECT 1065.0000 502.8000 1066.2001 503.7000 ;
	    RECT 1065.0000 501.9000 1067.7001 502.8000 ;
	    RECT 1066.5000 500.1000 1067.7001 501.9000 ;
	    RECT 1072.2001 501.9000 1073.4000 509.7000 ;
	    RECT 1074.6000 504.0000 1075.8000 509.7000 ;
	    RECT 1077.0000 506.7000 1078.2001 509.7000 ;
	    RECT 1074.6000 502.8000 1076.1000 504.0000 ;
	    RECT 1096.2001 503.7000 1097.4000 509.7000 ;
	    RECT 1100.1000 504.6000 1101.3000 509.7000 ;
	    RECT 1098.6000 503.7000 1101.3000 504.6000 ;
	    RECT 1072.2001 501.0000 1074.0000 501.9000 ;
	    RECT 1066.5000 498.9000 1072.2001 500.1000 ;
	    RECT 1028.7001 498.0000 1029.9000 498.3000 ;
	    RECT 1028.7001 497.1000 1035.3000 498.0000 ;
	    RECT 1036.2001 497.4000 1037.4000 498.6000 ;
	    RECT 1062.6000 498.0000 1063.8000 498.9000 ;
	    RECT 1073.1000 498.0000 1074.0000 501.0000 ;
	    RECT 1038.3000 497.1000 1063.8000 498.0000 ;
	    RECT 1072.8000 497.1000 1074.0000 498.0000 ;
	    RECT 1070.7001 496.2000 1071.9000 496.5000 ;
	    RECT 1031.4000 494.4000 1032.6000 495.6000 ;
	    RECT 1033.5000 495.3000 1071.9000 496.2000 ;
	    RECT 1036.5000 495.0000 1037.7001 495.3000 ;
	    RECT 1072.8000 494.4000 1073.7001 497.1000 ;
	    RECT 1074.9000 496.2000 1076.1000 502.8000 ;
	    RECT 1096.2001 502.5000 1097.4000 502.8000 ;
	    RECT 1091.4000 501.4500 1092.6000 501.6000 ;
	    RECT 1096.2001 501.4500 1097.4000 501.6000 ;
	    RECT 1091.4000 500.5500 1097.4000 501.4500 ;
	    RECT 1091.4000 500.4000 1092.6000 500.5500 ;
	    RECT 1096.2001 500.4000 1097.4000 500.5500 ;
	    RECT 1098.6000 499.5000 1099.8000 503.7000 ;
	    RECT 1134.6000 500.7000 1135.8000 509.7000 ;
	    RECT 1140.0000 501.3000 1141.2001 509.7000 ;
	    RECT 1161.0000 503.7000 1162.2001 509.7000 ;
	    RECT 1164.9000 504.6000 1166.1000 509.7000 ;
	    RECT 1163.4000 503.7000 1166.1000 504.6000 ;
	    RECT 1161.0000 502.5000 1162.2001 502.8000 ;
	    RECT 1140.0000 500.7000 1142.7001 501.3000 ;
	    RECT 1140.3000 500.4000 1142.7001 500.7000 ;
	    RECT 1161.0000 500.4000 1162.2001 501.6000 ;
	    RECT 1098.6000 498.4500 1099.8000 498.6000 ;
	    RECT 1132.2001 498.4500 1133.4000 498.6000 ;
	    RECT 1098.6000 497.5500 1133.4000 498.4500 ;
	    RECT 1098.6000 497.4000 1099.8000 497.5500 ;
	    RECT 1132.2001 497.4000 1133.4000 497.5500 ;
	    RECT 1137.0000 497.4000 1138.2001 498.6000 ;
	    RECT 1139.1000 497.4000 1139.4000 498.6000 ;
	    RECT 1134.6000 496.5000 1135.8000 496.8000 ;
	    RECT 1141.8000 496.5000 1142.7001 500.4000 ;
	    RECT 1163.4000 499.5000 1164.6000 503.7000 ;
	    RECT 1191.6000 501.3000 1192.8000 509.7000 ;
	    RECT 1190.1000 500.7000 1192.8000 501.3000 ;
	    RECT 1197.0000 500.7000 1198.2001 509.7000 ;
	    RECT 1221.0000 500.7000 1222.2001 509.7000 ;
	    RECT 1226.4000 501.3000 1227.6000 509.7000 ;
	    RECT 1255.5000 503.7000 1256.7001 509.7000 ;
	    RECT 1259.4000 503.7000 1260.6000 509.7000 ;
	    RECT 1261.8000 506.7000 1263.0000 509.7000 ;
	    RECT 1261.5000 505.5000 1262.7001 505.8000 ;
	    RECT 1226.4000 500.7000 1229.1000 501.3000 ;
	    RECT 1190.1000 500.4000 1192.5000 500.7000 ;
	    RECT 1226.7001 500.4000 1229.1000 500.7000 ;
	    RECT 1257.0000 500.4000 1258.2001 501.6000 ;
	    RECT 1163.4000 498.4500 1164.6000 498.6000 ;
	    RECT 1187.4000 498.4500 1188.6000 498.6000 ;
	    RECT 1163.4000 497.5500 1188.6000 498.4500 ;
	    RECT 1163.4000 497.4000 1164.6000 497.5500 ;
	    RECT 1187.4000 497.4000 1188.6000 497.5500 ;
	    RECT 1190.1000 496.5000 1191.0000 500.4000 ;
	    RECT 1193.4000 497.4000 1193.7001 498.6000 ;
	    RECT 1194.6000 497.4000 1195.8000 498.6000 ;
	    RECT 1223.4000 497.4000 1224.6000 498.6000 ;
	    RECT 1225.5000 497.4000 1225.8000 498.6000 ;
	    RECT 1197.0000 496.5000 1198.2001 496.8000 ;
	    RECT 1221.0000 496.5000 1222.2001 496.8000 ;
	    RECT 1228.2001 496.5000 1229.1000 500.4000 ;
	    RECT 1257.0000 499.2000 1258.2001 499.5000 ;
	    RECT 1254.6000 497.4000 1255.8000 498.6000 ;
	    RECT 1259.4000 498.3000 1260.3000 503.7000 ;
	    RECT 1261.8000 503.4000 1263.0000 504.6000 ;
	    RECT 1285.8000 504.0000 1287.0000 509.7000 ;
	    RECT 1288.2001 504.9000 1289.4000 509.7000 ;
	    RECT 1290.6000 504.0000 1291.8000 509.7000 ;
	    RECT 1285.8000 503.7000 1291.8000 504.0000 ;
	    RECT 1293.0000 503.7000 1294.2001 509.7000 ;
	    RECT 1317.9000 503.7000 1319.1000 509.7000 ;
	    RECT 1321.8000 503.7000 1323.0000 509.7000 ;
	    RECT 1324.2001 506.7000 1325.4000 509.7000 ;
	    RECT 1323.9000 505.5000 1325.1000 505.8000 ;
	    RECT 1286.1000 503.1000 1291.5000 503.7000 ;
	    RECT 1293.0000 502.5000 1293.9000 503.7000 ;
	    RECT 1285.8000 500.4000 1287.0000 501.6000 ;
	    RECT 1287.9000 500.7000 1288.2001 502.2000 ;
	    RECT 1290.3000 500.4000 1292.1000 501.6000 ;
	    RECT 1293.0000 501.4500 1294.2001 501.6000 ;
	    RECT 1317.0000 501.4500 1318.2001 501.6000 ;
	    RECT 1293.0000 500.5500 1318.2001 501.4500 ;
	    RECT 1293.0000 500.4000 1294.2001 500.5500 ;
	    RECT 1317.0000 500.4000 1318.2001 500.5500 ;
	    RECT 1319.4000 500.4000 1320.6000 501.6000 ;
	    RECT 1288.2001 499.5000 1289.4000 499.8000 ;
	    RECT 1261.8000 498.4500 1263.0000 498.6000 ;
	    RECT 1288.2001 498.4500 1289.4000 498.6000 ;
	    RECT 1256.7001 496.8000 1257.0000 498.3000 ;
	    RECT 1259.4000 497.4000 1260.9000 498.3000 ;
	    RECT 1261.8000 497.5500 1289.4000 498.4500 ;
	    RECT 1261.8000 497.4000 1263.0000 497.5500 ;
	    RECT 1288.2001 497.4000 1289.4000 497.5500 ;
	    RECT 1041.0000 494.1000 1042.2001 494.4000 ;
	    RECT 1034.1000 493.5000 1042.2001 494.1000 ;
	    RECT 1032.9000 493.2000 1042.2001 493.5000 ;
	    RECT 1043.7001 493.5000 1056.6000 494.4000 ;
	    RECT 1029.0000 492.0000 1031.4000 493.2000 ;
	    RECT 1032.9000 492.3000 1035.0000 493.2000 ;
	    RECT 1043.7001 492.3000 1044.6000 493.5000 ;
	    RECT 1055.4000 493.2000 1056.6000 493.5000 ;
	    RECT 1060.2001 493.5000 1073.7001 494.4000 ;
	    RECT 1074.6000 495.0000 1076.1000 496.2000 ;
	    RECT 1074.6000 493.5000 1075.8000 495.0000 ;
	    RECT 1060.2001 493.2000 1061.4000 493.5000 ;
	    RECT 1030.5000 491.4000 1031.4000 492.0000 ;
	    RECT 1035.9000 491.4000 1044.6000 492.3000 ;
	    RECT 1045.5000 491.4000 1049.4000 492.6000 ;
	    RECT 1026.6000 490.2000 1029.6000 491.1000 ;
	    RECT 1030.5000 490.2000 1036.8000 491.4000 ;
	    RECT 1028.7001 489.3000 1029.6000 490.2000 ;
	    RECT 894.6000 483.3000 895.8000 489.3000 ;
	    RECT 1026.6000 483.3000 1027.8000 489.3000 ;
	    RECT 1028.7001 488.4000 1030.2001 489.3000 ;
	    RECT 1029.0000 483.3000 1030.2001 488.4000 ;
	    RECT 1031.4000 482.4000 1032.6000 489.3000 ;
	    RECT 1033.8000 483.3000 1035.0000 490.2000 ;
	    RECT 1036.2001 483.3000 1037.4000 489.3000 ;
	    RECT 1038.6000 483.3000 1039.8000 487.5000 ;
	    RECT 1041.0000 483.3000 1042.2001 487.5000 ;
	    RECT 1043.4000 483.3000 1044.6000 490.5000 ;
	    RECT 1045.8000 483.3000 1047.0000 489.3000 ;
	    RECT 1048.2001 483.3000 1049.4000 490.5000 ;
	    RECT 1050.6000 483.3000 1051.8000 489.3000 ;
	    RECT 1053.0000 483.3000 1054.2001 492.6000 ;
	    RECT 1065.0000 491.4000 1068.9000 492.6000 ;
	    RECT 1057.8000 490.2000 1064.1000 491.4000 ;
	    RECT 1055.4000 483.3000 1056.6000 487.5000 ;
	    RECT 1057.8000 483.3000 1059.0000 487.5000 ;
	    RECT 1060.2001 483.3000 1061.4000 487.5000 ;
	    RECT 1062.6000 483.3000 1063.8000 489.3000 ;
	    RECT 1065.0000 483.3000 1066.2001 491.4000 ;
	    RECT 1072.8000 491.1000 1073.7001 493.5000 ;
	    RECT 1074.6000 491.4000 1075.8000 492.6000 ;
	    RECT 1069.8000 490.2000 1073.7001 491.1000 ;
	    RECT 1067.4000 483.3000 1068.6000 489.3000 ;
	    RECT 1069.8000 483.3000 1071.0000 490.2000 ;
	    RECT 1072.2001 483.3000 1073.4000 489.3000 ;
	    RECT 1074.6000 483.3000 1075.8000 490.5000 ;
	    RECT 1077.0000 483.3000 1078.2001 489.3000 ;
	    RECT 1096.2001 483.3000 1097.4000 489.3000 ;
	    RECT 1098.6000 483.3000 1099.8000 496.5000 ;
	    RECT 1101.0000 495.4500 1102.2001 495.6000 ;
	    RECT 1103.4000 495.4500 1104.6000 495.6000 ;
	    RECT 1110.6000 495.4500 1111.8000 495.6000 ;
	    RECT 1101.0000 494.5500 1111.8000 495.4500 ;
	    RECT 1101.0000 494.4000 1102.2001 494.5500 ;
	    RECT 1103.4000 494.4000 1104.6000 494.5500 ;
	    RECT 1110.6000 494.4000 1111.8000 494.5500 ;
	    RECT 1127.4000 495.4500 1128.6000 495.6000 ;
	    RECT 1134.6000 495.4500 1135.8000 495.6000 ;
	    RECT 1127.4000 494.5500 1135.8000 495.4500 ;
	    RECT 1127.4000 494.4000 1128.6000 494.5500 ;
	    RECT 1134.6000 494.4000 1135.8000 494.5500 ;
	    RECT 1141.8000 495.4500 1143.0000 495.6000 ;
	    RECT 1161.0000 495.4500 1162.2001 495.6000 ;
	    RECT 1141.8000 494.5500 1162.2001 495.4500 ;
	    RECT 1141.8000 494.4000 1143.0000 494.5500 ;
	    RECT 1161.0000 494.4000 1162.2001 494.5500 ;
	    RECT 1139.4000 493.5000 1140.6000 493.8000 ;
	    RECT 1101.0000 493.2000 1102.2001 493.5000 ;
	    RECT 1132.2001 492.4500 1133.4000 492.6000 ;
	    RECT 1139.4000 492.4500 1140.6000 492.6000 ;
	    RECT 1132.2001 491.5500 1140.6000 492.4500 ;
	    RECT 1132.2001 491.4000 1133.4000 491.5500 ;
	    RECT 1139.4000 491.4000 1140.6000 491.5500 ;
	    RECT 1141.8000 490.5000 1142.7001 493.5000 ;
	    RECT 1137.3000 489.6000 1142.7001 490.5000 ;
	    RECT 1137.3000 489.3000 1138.2001 489.6000 ;
	    RECT 1101.0000 483.3000 1102.2001 489.3000 ;
	    RECT 1134.6000 483.3000 1135.8000 489.3000 ;
	    RECT 1137.0000 483.3000 1138.2001 489.3000 ;
	    RECT 1141.8000 489.3000 1142.7001 489.6000 ;
	    RECT 1139.4000 483.3000 1140.6000 488.7000 ;
	    RECT 1141.8000 483.3000 1143.0000 489.3000 ;
	    RECT 1161.0000 483.3000 1162.2001 489.3000 ;
	    RECT 1163.4000 483.3000 1164.6000 496.5000 ;
	    RECT 1165.8000 494.4000 1167.0000 495.6000 ;
	    RECT 1189.8000 494.4000 1191.0000 495.6000 ;
	    RECT 1197.0000 494.4000 1198.2001 495.6000 ;
	    RECT 1199.4000 495.4500 1200.6000 495.6000 ;
	    RECT 1221.0000 495.4500 1222.2001 495.6000 ;
	    RECT 1199.4000 494.5500 1222.2001 495.4500 ;
	    RECT 1199.4000 494.4000 1200.6000 494.5500 ;
	    RECT 1221.0000 494.4000 1222.2001 494.5500 ;
	    RECT 1228.2001 495.4500 1229.4000 495.6000 ;
	    RECT 1252.2001 495.4500 1253.4000 495.6000 ;
	    RECT 1228.2001 494.5500 1253.4000 495.4500 ;
	    RECT 1261.8000 495.3000 1262.7001 496.5000 ;
	    RECT 1290.3000 495.3000 1291.2001 500.4000 ;
	    RECT 1319.4000 499.2000 1320.6000 499.5000 ;
	    RECT 1302.6000 498.4500 1303.8000 498.6000 ;
	    RECT 1317.0000 498.4500 1318.2001 498.6000 ;
	    RECT 1302.6000 497.5500 1318.2001 498.4500 ;
	    RECT 1321.8000 498.3000 1322.7001 503.7000 ;
	    RECT 1324.2001 503.4000 1325.4000 504.6000 ;
	    RECT 1350.0000 501.3000 1351.2001 509.7000 ;
	    RECT 1348.5000 500.7000 1351.2001 501.3000 ;
	    RECT 1355.4000 500.7000 1356.6000 509.7000 ;
	    RECT 1387.5000 503.7000 1388.7001 509.7000 ;
	    RECT 1391.4000 503.7000 1392.6000 509.7000 ;
	    RECT 1393.8000 506.7000 1395.0000 509.7000 ;
	    RECT 1393.5000 505.5000 1394.7001 505.8000 ;
	    RECT 1393.8000 504.4500 1395.0000 504.6000 ;
	    RECT 1415.4000 504.4500 1416.6000 504.6000 ;
	    RECT 1348.5000 500.4000 1350.9000 500.7000 ;
	    RECT 1389.0000 500.4000 1390.2001 501.6000 ;
	    RECT 1324.2001 498.4500 1325.4000 498.6000 ;
	    RECT 1326.6000 498.4500 1327.8000 498.6000 ;
	    RECT 1302.6000 497.4000 1303.8000 497.5500 ;
	    RECT 1317.0000 497.4000 1318.2001 497.5500 ;
	    RECT 1319.1000 496.8000 1319.4000 498.3000 ;
	    RECT 1321.8000 497.4000 1323.3000 498.3000 ;
	    RECT 1324.2001 497.5500 1327.8000 498.4500 ;
	    RECT 1324.2001 497.4000 1325.4000 497.5500 ;
	    RECT 1326.6000 497.4000 1327.8000 497.5500 ;
	    RECT 1348.5000 496.5000 1349.4000 500.4000 ;
	    RECT 1389.0000 499.2000 1390.2001 499.5000 ;
	    RECT 1351.8000 497.4000 1352.1000 498.6000 ;
	    RECT 1353.0000 497.4000 1354.2001 498.6000 ;
	    RECT 1386.6000 497.4000 1387.8000 498.6000 ;
	    RECT 1391.4000 498.3000 1392.3000 503.7000 ;
	    RECT 1393.8000 503.5500 1416.6000 504.4500 ;
	    RECT 1393.8000 503.4000 1395.0000 503.5500 ;
	    RECT 1415.4000 503.4000 1416.6000 503.5500 ;
	    RECT 1417.8000 500.7000 1419.0000 509.7000 ;
	    RECT 1423.2001 501.3000 1424.4000 509.7000 ;
	    RECT 1423.2001 500.7000 1425.9000 501.3000 ;
	    RECT 1451.4000 500.7000 1452.6000 509.7000 ;
	    RECT 1456.8000 501.3000 1458.0000 509.7000 ;
	    RECT 1456.8000 500.7000 1459.5000 501.3000 ;
	    RECT 1485.0000 500.7000 1486.2001 509.7000 ;
	    RECT 1490.4000 501.3000 1491.6000 509.7000 ;
	    RECT 1512.3000 504.6000 1513.5000 509.7000 ;
	    RECT 1512.3000 503.7000 1515.0000 504.6000 ;
	    RECT 1516.2001 503.7000 1517.4000 509.7000 ;
	    RECT 1542.6000 506.7000 1543.8000 509.7000 ;
	    RECT 1542.9000 505.5000 1544.1000 505.8000 ;
	    RECT 1518.6000 504.4500 1519.8000 504.6000 ;
	    RECT 1535.4000 504.4500 1536.6000 504.6000 ;
	    RECT 1542.6000 504.4500 1543.8000 504.6000 ;
	    RECT 1490.4000 500.7000 1493.1000 501.3000 ;
	    RECT 1423.5000 500.4000 1425.9000 500.7000 ;
	    RECT 1457.1000 500.4000 1459.5000 500.7000 ;
	    RECT 1490.7001 500.4000 1493.1000 500.7000 ;
	    RECT 1393.8000 498.4500 1395.0000 498.6000 ;
	    RECT 1410.6000 498.4500 1411.8000 498.6000 ;
	    RECT 1388.7001 496.8000 1389.0000 498.3000 ;
	    RECT 1391.4000 497.4000 1392.9000 498.3000 ;
	    RECT 1393.8000 497.5500 1411.8000 498.4500 ;
	    RECT 1393.8000 497.4000 1395.0000 497.5500 ;
	    RECT 1410.6000 497.4000 1411.8000 497.5500 ;
	    RECT 1420.2001 497.4000 1421.4000 498.6000 ;
	    RECT 1422.3000 497.4000 1422.6000 498.6000 ;
	    RECT 1355.4000 496.5000 1356.6000 496.8000 ;
	    RECT 1417.8000 496.5000 1419.0000 496.8000 ;
	    RECT 1425.0000 496.5000 1425.9000 500.4000 ;
	    RECT 1453.8000 497.4000 1455.0000 498.6000 ;
	    RECT 1455.9000 497.4000 1456.2001 498.6000 ;
	    RECT 1451.4000 496.5000 1452.6000 496.8000 ;
	    RECT 1458.6000 496.5000 1459.5000 500.4000 ;
	    RECT 1487.4000 497.4000 1488.6000 498.6000 ;
	    RECT 1489.5000 497.4000 1489.8000 498.6000 ;
	    RECT 1485.0000 496.5000 1486.2001 496.8000 ;
	    RECT 1492.2001 496.5000 1493.1000 500.4000 ;
	    RECT 1513.8000 499.5000 1515.0000 503.7000 ;
	    RECT 1518.6000 503.5500 1543.8000 504.4500 ;
	    RECT 1545.0000 503.7000 1546.2001 509.7000 ;
	    RECT 1548.9000 503.7000 1550.1000 509.7000 ;
	    RECT 1518.6000 503.4000 1519.8000 503.5500 ;
	    RECT 1535.4000 503.4000 1536.6000 503.5500 ;
	    RECT 1542.6000 503.4000 1543.8000 503.5500 ;
	    RECT 1516.2001 502.5000 1517.4000 502.8000 ;
	    RECT 1516.2001 500.4000 1517.4000 501.6000 ;
	    RECT 1513.8000 498.4500 1515.0000 498.6000 ;
	    RECT 1530.6000 498.4500 1531.8000 498.6000 ;
	    RECT 1513.8000 497.5500 1531.8000 498.4500 ;
	    RECT 1513.8000 497.4000 1515.0000 497.5500 ;
	    RECT 1530.6000 497.4000 1531.8000 497.5500 ;
	    RECT 1542.6000 497.4000 1543.8000 498.6000 ;
	    RECT 1545.3000 498.3000 1546.2001 503.7000 ;
	    RECT 1547.4000 500.4000 1548.6000 501.6000 ;
	    RECT 1547.4000 499.2000 1548.6000 499.5000 ;
	    RECT 1544.7001 497.4000 1546.2001 498.3000 ;
	    RECT 1548.6000 496.8000 1548.9000 498.3000 ;
	    RECT 1549.8000 497.4000 1551.0000 498.6000 ;
	    RECT 1228.2001 494.4000 1229.4000 494.5500 ;
	    RECT 1252.2001 494.4000 1253.4000 494.5500 ;
	    RECT 1254.6000 494.4000 1260.6000 495.3000 ;
	    RECT 1192.2001 493.5000 1193.4000 493.8000 ;
	    RECT 1165.8000 493.2000 1167.0000 493.5000 ;
	    RECT 1190.1000 490.5000 1191.0000 493.5000 ;
	    RECT 1192.2001 491.4000 1193.4000 492.6000 ;
	    RECT 1197.1500 492.4500 1198.0500 494.4000 ;
	    RECT 1225.8000 493.5000 1227.0000 493.8000 ;
	    RECT 1221.0000 492.4500 1222.2001 492.6000 ;
	    RECT 1197.1500 491.5500 1222.2001 492.4500 ;
	    RECT 1221.0000 491.4000 1222.2001 491.5500 ;
	    RECT 1225.8000 491.4000 1227.0000 492.6000 ;
	    RECT 1228.2001 490.5000 1229.1000 493.5000 ;
	    RECT 1190.1000 489.6000 1195.5000 490.5000 ;
	    RECT 1190.1000 489.3000 1191.0000 489.6000 ;
	    RECT 1165.8000 483.3000 1167.0000 489.3000 ;
	    RECT 1189.8000 483.3000 1191.0000 489.3000 ;
	    RECT 1194.6000 489.3000 1195.5000 489.6000 ;
	    RECT 1223.7001 489.6000 1229.1000 490.5000 ;
	    RECT 1223.7001 489.3000 1224.6000 489.6000 ;
	    RECT 1192.2001 483.3000 1193.4000 488.7000 ;
	    RECT 1194.6000 483.3000 1195.8000 489.3000 ;
	    RECT 1197.0000 483.3000 1198.2001 489.3000 ;
	    RECT 1221.0000 483.3000 1222.2001 489.3000 ;
	    RECT 1223.4000 483.3000 1224.6000 489.3000 ;
	    RECT 1228.2001 489.3000 1229.1000 489.6000 ;
	    RECT 1225.8000 483.3000 1227.0000 488.7000 ;
	    RECT 1228.2001 483.3000 1229.4000 489.3000 ;
	    RECT 1254.6000 483.3000 1255.8000 494.4000 ;
	    RECT 1257.0000 483.3000 1258.2001 493.5000 ;
	    RECT 1259.4000 483.3000 1260.6000 494.4000 ;
	    RECT 1261.8000 483.3000 1263.0000 495.3000 ;
	    RECT 1285.8000 483.3000 1287.0000 495.3000 ;
	    RECT 1289.7001 494.4000 1291.2001 495.3000 ;
	    RECT 1293.0000 495.4500 1294.2001 495.6000 ;
	    RECT 1314.6000 495.4500 1315.8000 495.6000 ;
	    RECT 1293.0000 494.5500 1315.8000 495.4500 ;
	    RECT 1324.2001 495.3000 1325.1000 496.5000 ;
	    RECT 1345.8000 495.4500 1347.0000 495.6000 ;
	    RECT 1348.2001 495.4500 1349.4000 495.6000 ;
	    RECT 1293.0000 494.4000 1294.2001 494.5500 ;
	    RECT 1314.6000 494.4000 1315.8000 494.5500 ;
	    RECT 1317.0000 494.4000 1323.0000 495.3000 ;
	    RECT 1289.7001 483.3000 1290.9000 494.4000 ;
	    RECT 1292.1000 492.6000 1293.0000 493.5000 ;
	    RECT 1291.8000 491.4000 1293.0000 492.6000 ;
	    RECT 1292.1000 483.3000 1293.3000 489.3000 ;
	    RECT 1317.0000 483.3000 1318.2001 494.4000 ;
	    RECT 1319.4000 483.3000 1320.6000 493.5000 ;
	    RECT 1321.8000 483.3000 1323.0000 494.4000 ;
	    RECT 1324.2001 483.3000 1325.4000 495.3000 ;
	    RECT 1345.8000 494.5500 1349.4000 495.4500 ;
	    RECT 1345.8000 494.4000 1347.0000 494.5500 ;
	    RECT 1348.2001 494.4000 1349.4000 494.5500 ;
	    RECT 1355.4000 494.4000 1356.6000 495.6000 ;
	    RECT 1393.8000 495.3000 1394.7001 496.5000 ;
	    RECT 1415.4000 495.4500 1416.6000 495.6000 ;
	    RECT 1417.8000 495.4500 1419.0000 495.6000 ;
	    RECT 1386.6000 494.4000 1392.6000 495.3000 ;
	    RECT 1350.6000 493.5000 1351.8000 493.8000 ;
	    RECT 1348.5000 490.5000 1349.4000 493.5000 ;
	    RECT 1350.6000 491.4000 1351.8000 492.6000 ;
	    RECT 1348.5000 489.6000 1353.9000 490.5000 ;
	    RECT 1348.5000 489.3000 1349.4000 489.6000 ;
	    RECT 1348.2001 483.3000 1349.4000 489.3000 ;
	    RECT 1353.0000 489.3000 1353.9000 489.6000 ;
	    RECT 1350.6000 483.3000 1351.8000 488.7000 ;
	    RECT 1353.0000 483.3000 1354.2001 489.3000 ;
	    RECT 1355.4000 483.3000 1356.6000 489.3000 ;
	    RECT 1386.6000 483.3000 1387.8000 494.4000 ;
	    RECT 1389.0000 483.3000 1390.2001 493.5000 ;
	    RECT 1391.4000 483.3000 1392.6000 494.4000 ;
	    RECT 1393.8000 483.3000 1395.0000 495.3000 ;
	    RECT 1415.4000 494.5500 1419.0000 495.4500 ;
	    RECT 1415.4000 494.4000 1416.6000 494.5500 ;
	    RECT 1417.8000 494.4000 1419.0000 494.5500 ;
	    RECT 1425.0000 494.4000 1426.2001 495.6000 ;
	    RECT 1441.8000 495.4500 1443.0000 495.6000 ;
	    RECT 1451.4000 495.4500 1452.6000 495.6000 ;
	    RECT 1441.8000 494.5500 1452.6000 495.4500 ;
	    RECT 1441.8000 494.4000 1443.0000 494.5500 ;
	    RECT 1451.4000 494.4000 1452.6000 494.5500 ;
	    RECT 1458.6000 495.4500 1459.8000 495.6000 ;
	    RECT 1461.0000 495.4500 1462.2001 495.6000 ;
	    RECT 1485.0000 495.4500 1486.2001 495.6000 ;
	    RECT 1458.6000 494.5500 1486.2001 495.4500 ;
	    RECT 1458.6000 494.4000 1459.8000 494.5500 ;
	    RECT 1461.0000 494.4000 1462.2001 494.5500 ;
	    RECT 1485.0000 494.4000 1486.2001 494.5500 ;
	    RECT 1492.2001 494.4000 1493.4000 495.6000 ;
	    RECT 1494.6000 495.4500 1495.8000 495.6000 ;
	    RECT 1511.4000 495.4500 1512.6000 495.6000 ;
	    RECT 1494.6000 494.5500 1512.6000 495.4500 ;
	    RECT 1494.6000 494.4000 1495.8000 494.5500 ;
	    RECT 1511.4000 494.4000 1512.6000 494.5500 ;
	    RECT 1422.6000 493.5000 1423.8000 493.8000 ;
	    RECT 1456.2001 493.5000 1457.4000 493.8000 ;
	    RECT 1489.8000 493.5000 1491.0000 493.8000 ;
	    RECT 1422.6000 491.4000 1423.8000 492.6000 ;
	    RECT 1425.0000 490.5000 1425.9000 493.5000 ;
	    RECT 1427.4000 492.4500 1428.6000 492.6000 ;
	    RECT 1456.2001 492.4500 1457.4000 492.6000 ;
	    RECT 1427.4000 491.5500 1457.4000 492.4500 ;
	    RECT 1427.4000 491.4000 1428.6000 491.5500 ;
	    RECT 1456.2001 491.4000 1457.4000 491.5500 ;
	    RECT 1458.6000 490.5000 1459.5000 493.5000 ;
	    RECT 1489.8000 491.4000 1491.0000 492.6000 ;
	    RECT 1492.2001 490.5000 1493.1000 493.5000 ;
	    RECT 1511.4000 493.2000 1512.6000 493.5000 ;
	    RECT 1420.5000 489.6000 1425.9000 490.5000 ;
	    RECT 1420.5000 489.3000 1421.4000 489.6000 ;
	    RECT 1417.8000 483.3000 1419.0000 489.3000 ;
	    RECT 1420.2001 483.3000 1421.4000 489.3000 ;
	    RECT 1425.0000 489.3000 1425.9000 489.6000 ;
	    RECT 1454.1000 489.6000 1459.5000 490.5000 ;
	    RECT 1454.1000 489.3000 1455.0000 489.6000 ;
	    RECT 1422.6000 483.3000 1423.8000 488.7000 ;
	    RECT 1425.0000 483.3000 1426.2001 489.3000 ;
	    RECT 1451.4000 483.3000 1452.6000 489.3000 ;
	    RECT 1453.8000 483.3000 1455.0000 489.3000 ;
	    RECT 1458.6000 489.3000 1459.5000 489.6000 ;
	    RECT 1487.7001 489.6000 1493.1000 490.5000 ;
	    RECT 1487.7001 489.3000 1488.6000 489.6000 ;
	    RECT 1456.2001 483.3000 1457.4000 488.7000 ;
	    RECT 1458.6000 483.3000 1459.8000 489.3000 ;
	    RECT 1485.0000 483.3000 1486.2001 489.3000 ;
	    RECT 1487.4000 483.3000 1488.6000 489.3000 ;
	    RECT 1492.2001 489.3000 1493.1000 489.6000 ;
	    RECT 1489.8000 483.3000 1491.0000 488.7000 ;
	    RECT 1492.2001 483.3000 1493.4000 489.3000 ;
	    RECT 1511.4000 483.3000 1512.6000 489.3000 ;
	    RECT 1513.8000 483.3000 1515.0000 496.5000 ;
	    RECT 1542.9000 495.3000 1543.8000 496.5000 ;
	    RECT 1516.2001 483.3000 1517.4000 489.3000 ;
	    RECT 1542.6000 483.3000 1543.8000 495.3000 ;
	    RECT 1545.0000 494.4000 1551.0000 495.3000 ;
	    RECT 1545.0000 483.3000 1546.2001 494.4000 ;
	    RECT 1547.4000 483.3000 1548.6000 493.5000 ;
	    RECT 1549.8000 483.3000 1551.0000 494.4000 ;
	    RECT 1.2000 480.6000 1569.0000 482.4000 ;
	    RECT 124.2000 473.7000 125.4000 479.7000 ;
	    RECT 126.6000 474.6000 127.8000 479.7000 ;
	    RECT 126.3000 473.7000 127.8000 474.6000 ;
	    RECT 129.0000 473.7000 130.2000 480.6000 ;
	    RECT 126.3000 472.8000 127.2000 473.7000 ;
	    RECT 131.4000 472.8000 132.6000 479.7000 ;
	    RECT 133.8000 473.7000 135.0000 479.7000 ;
	    RECT 136.2000 475.5000 137.4000 479.7000 ;
	    RECT 138.6000 475.5000 139.8000 479.7000 ;
	    RECT 124.2000 471.9000 127.2000 472.8000 ;
	    RECT 124.2000 463.5000 125.4000 471.9000 ;
	    RECT 128.1000 471.6000 134.4000 472.8000 ;
	    RECT 141.0000 472.5000 142.2000 479.7000 ;
	    RECT 143.4000 473.7000 144.6000 479.7000 ;
	    RECT 145.8000 472.5000 147.0000 479.7000 ;
	    RECT 148.2000 473.7000 149.4000 479.7000 ;
	    RECT 128.1000 471.0000 129.0000 471.6000 ;
	    RECT 126.6000 469.8000 129.0000 471.0000 ;
	    RECT 133.5000 470.7000 142.2000 471.6000 ;
	    RECT 130.5000 469.8000 132.6000 470.7000 ;
	    RECT 130.5000 469.5000 139.8000 469.8000 ;
	    RECT 131.7000 468.9000 139.8000 469.5000 ;
	    RECT 138.6000 468.6000 139.8000 468.9000 ;
	    RECT 141.3000 469.5000 142.2000 470.7000 ;
	    RECT 143.1000 470.4000 147.0000 471.6000 ;
	    RECT 150.6000 470.4000 151.8000 479.7000 ;
	    RECT 153.0000 475.5000 154.2000 479.7000 ;
	    RECT 155.4000 475.5000 156.6000 479.7000 ;
	    RECT 157.8000 475.5000 159.0000 479.7000 ;
	    RECT 160.2000 473.7000 161.4000 479.7000 ;
	    RECT 155.4000 471.6000 161.7000 472.8000 ;
	    RECT 162.6000 471.6000 163.8000 479.7000 ;
	    RECT 165.0000 473.7000 166.2000 479.7000 ;
	    RECT 167.4000 472.8000 168.6000 479.7000 ;
	    RECT 169.8000 473.7000 171.0000 479.7000 ;
	    RECT 167.4000 471.9000 171.3000 472.8000 ;
	    RECT 172.2000 472.5000 173.4000 479.7000 ;
	    RECT 174.6000 473.7000 175.8000 479.7000 ;
	    RECT 162.6000 470.4000 166.5000 471.6000 ;
	    RECT 153.0000 469.5000 154.2000 469.8000 ;
	    RECT 141.3000 468.6000 154.2000 469.5000 ;
	    RECT 157.8000 469.5000 159.0000 469.8000 ;
	    RECT 170.4000 469.5000 171.3000 471.9000 ;
	    RECT 172.2000 470.4000 173.4000 471.6000 ;
	    RECT 157.8000 468.6000 171.3000 469.5000 ;
	    RECT 129.0000 467.4000 130.2000 468.6000 ;
	    RECT 134.1000 467.7000 135.3000 468.0000 ;
	    RECT 131.1000 466.8000 169.5000 467.7000 ;
	    RECT 168.3000 466.5000 169.5000 466.8000 ;
	    RECT 170.4000 465.9000 171.3000 468.6000 ;
	    RECT 172.2000 468.0000 173.4000 469.5000 ;
	    RECT 194.7000 468.9000 195.9000 479.7000 ;
	    RECT 172.2000 466.8000 173.7000 468.0000 ;
	    RECT 194.7000 467.7000 197.4000 468.9000 ;
	    RECT 198.6000 467.7000 199.8000 479.7000 ;
	    RECT 220.2000 473.7000 221.4000 479.7000 ;
	    RECT 126.3000 465.0000 132.9000 465.9000 ;
	    RECT 126.3000 464.7000 127.5000 465.0000 ;
	    RECT 133.8000 464.4000 135.0000 465.6000 ;
	    RECT 135.9000 465.0000 161.4000 465.9000 ;
	    RECT 170.4000 465.0000 171.6000 465.9000 ;
	    RECT 160.2000 464.1000 161.4000 465.0000 ;
	    RECT 124.2000 462.3000 137.4000 463.5000 ;
	    RECT 138.3000 462.9000 141.3000 464.1000 ;
	    RECT 147.0000 462.9000 151.8000 464.1000 ;
	    RECT 124.2000 453.3000 125.4000 462.3000 ;
	    RECT 127.8000 460.2000 132.3000 461.4000 ;
	    RECT 131.1000 459.3000 132.3000 460.2000 ;
	    RECT 140.1000 459.3000 141.3000 462.9000 ;
	    RECT 143.4000 461.4000 144.6000 462.6000 ;
	    RECT 151.2000 461.7000 152.4000 462.0000 ;
	    RECT 145.8000 460.8000 152.4000 461.7000 ;
	    RECT 145.8000 460.5000 147.0000 460.8000 ;
	    RECT 143.4000 460.2000 144.6000 460.5000 ;
	    RECT 155.4000 459.6000 156.6000 463.8000 ;
	    RECT 164.1000 462.9000 169.8000 464.1000 ;
	    RECT 164.1000 461.1000 165.3000 462.9000 ;
	    RECT 170.7000 462.0000 171.6000 465.0000 ;
	    RECT 145.8000 459.3000 147.0000 459.6000 ;
	    RECT 129.0000 453.3000 130.2000 459.3000 ;
	    RECT 131.1000 458.1000 135.0000 459.3000 ;
	    RECT 140.1000 458.4000 147.0000 459.3000 ;
	    RECT 148.2000 458.4000 149.4000 459.6000 ;
	    RECT 150.3000 458.4000 150.6000 459.6000 ;
	    RECT 155.1000 458.4000 156.6000 459.6000 ;
	    RECT 162.6000 460.2000 165.3000 461.1000 ;
	    RECT 169.8000 461.1000 171.6000 462.0000 ;
	    RECT 162.6000 459.3000 163.8000 460.2000 ;
	    RECT 133.8000 453.3000 135.0000 458.1000 ;
	    RECT 160.2000 458.1000 163.8000 459.3000 ;
	    RECT 136.2000 453.3000 137.4000 457.5000 ;
	    RECT 138.6000 453.3000 139.8000 457.5000 ;
	    RECT 141.0000 453.3000 142.2000 457.5000 ;
	    RECT 143.4000 453.3000 144.6000 456.3000 ;
	    RECT 145.8000 453.3000 147.0000 457.5000 ;
	    RECT 148.2000 453.3000 149.4000 456.3000 ;
	    RECT 150.6000 453.3000 151.8000 457.5000 ;
	    RECT 153.0000 453.3000 154.2000 457.5000 ;
	    RECT 155.4000 453.3000 156.6000 457.5000 ;
	    RECT 157.8000 453.3000 159.0000 457.5000 ;
	    RECT 160.2000 453.3000 161.4000 458.1000 ;
	    RECT 165.0000 453.3000 166.2000 459.3000 ;
	    RECT 169.8000 453.3000 171.0000 461.1000 ;
	    RECT 172.5000 460.2000 173.7000 466.8000 ;
	    RECT 193.8000 466.5000 195.0000 466.8000 ;
	    RECT 193.8000 464.4000 195.0000 465.6000 ;
	    RECT 196.2000 463.5000 197.1000 467.7000 ;
	    RECT 222.6000 463.5000 223.8000 479.7000 ;
	    RECT 253.8000 467.7000 255.0000 479.7000 ;
	    RECT 257.7000 467.7000 260.7000 479.7000 ;
	    RECT 263.4000 467.7000 264.6000 479.7000 ;
	    RECT 283.5000 468.9000 284.7000 479.7000 ;
	    RECT 265.8000 468.4500 267.0000 468.6000 ;
	    RECT 275.4000 468.4500 276.6000 468.6000 ;
	    RECT 256.2000 464.4000 257.4000 465.6000 ;
	    RECT 258.6000 463.5000 259.5000 467.7000 ;
	    RECT 265.8000 467.5500 276.6000 468.4500 ;
	    RECT 283.5000 467.7000 286.2000 468.9000 ;
	    RECT 287.4000 467.7000 288.6000 479.7000 ;
	    RECT 297.0000 479.4000 298.2000 480.6000 ;
	    RECT 301.8000 473.7000 303.0000 479.7000 ;
	    RECT 265.8000 467.4000 267.0000 467.5500 ;
	    RECT 275.4000 467.4000 276.6000 467.5500 ;
	    RECT 282.6000 466.5000 283.8000 466.8000 ;
	    RECT 261.0000 464.4000 262.2000 465.6000 ;
	    RECT 273.0000 465.4500 274.2000 465.6000 ;
	    RECT 282.6000 465.4500 283.8000 465.6000 ;
	    RECT 273.0000 464.5500 283.8000 465.4500 ;
	    RECT 273.0000 464.4000 274.2000 464.5500 ;
	    RECT 282.6000 464.4000 283.8000 464.5500 ;
	    RECT 263.4000 463.5000 264.6000 463.8000 ;
	    RECT 285.0000 463.5000 285.9000 467.7000 ;
	    RECT 304.2000 463.5000 305.4000 479.7000 ;
	    RECT 318.6000 479.4000 319.8000 480.6000 ;
	    RECT 328.2000 467.7000 329.4000 479.7000 ;
	    RECT 332.1000 468.6000 333.3000 479.7000 ;
	    RECT 334.5000 473.7000 335.7000 479.7000 ;
	    RECT 354.6000 473.7000 355.8000 479.7000 ;
	    RECT 334.2000 470.4000 335.4000 471.6000 ;
	    RECT 334.5000 469.5000 335.4000 470.4000 ;
	    RECT 332.1000 467.7000 333.6000 468.6000 ;
	    RECT 330.6000 465.4500 331.8000 465.6000 ;
	    RECT 325.9500 464.5500 331.8000 465.4500 ;
	    RECT 256.2000 463.2000 257.4000 463.5000 ;
	    RECT 261.0000 463.2000 262.2000 463.5000 ;
	    RECT 196.2000 462.4500 197.4000 462.6000 ;
	    RECT 198.6000 462.4500 199.8000 462.6000 ;
	    RECT 196.2000 461.5500 199.8000 462.4500 ;
	    RECT 196.2000 461.4000 197.4000 461.5500 ;
	    RECT 198.6000 461.4000 199.8000 461.5500 ;
	    RECT 222.6000 462.4500 223.8000 462.6000 ;
	    RECT 241.8000 462.4500 243.0000 462.6000 ;
	    RECT 222.6000 461.5500 243.0000 462.4500 ;
	    RECT 222.6000 461.4000 223.8000 461.5500 ;
	    RECT 241.8000 461.4000 243.0000 461.5500 ;
	    RECT 244.2000 462.4500 245.4000 462.6000 ;
	    RECT 253.8000 462.4500 255.0000 462.6000 ;
	    RECT 244.2000 461.5500 255.0000 462.4500 ;
	    RECT 244.2000 461.4000 245.4000 461.5500 ;
	    RECT 253.8000 461.4000 255.0000 461.5500 ;
	    RECT 255.9000 460.8000 256.2000 462.3000 ;
	    RECT 258.6000 461.4000 259.8000 462.6000 ;
	    RECT 260.7000 461.4000 262.2000 462.3000 ;
	    RECT 263.4000 461.4000 264.6000 462.6000 ;
	    RECT 285.0000 462.4500 286.2000 462.6000 ;
	    RECT 294.6000 462.4500 295.8000 462.6000 ;
	    RECT 285.0000 461.5500 295.8000 462.4500 ;
	    RECT 285.0000 461.4000 286.2000 461.5500 ;
	    RECT 294.6000 461.4000 295.8000 461.5500 ;
	    RECT 304.2000 462.4500 305.4000 462.6000 ;
	    RECT 325.9500 462.4500 326.8500 464.5500 ;
	    RECT 330.6000 464.4000 331.8000 464.5500 ;
	    RECT 330.6000 463.2000 331.8000 463.5000 ;
	    RECT 332.7000 462.6000 333.6000 467.7000 ;
	    RECT 335.4000 467.4000 336.6000 468.6000 ;
	    RECT 357.0000 466.5000 358.2000 479.7000 ;
	    RECT 359.4000 473.7000 360.6000 479.7000 ;
	    RECT 373.8000 473.7000 375.0000 479.7000 ;
	    RECT 359.4000 469.5000 360.6000 469.8000 ;
	    RECT 359.4000 467.4000 360.6000 468.6000 ;
	    RECT 342.6000 465.4500 343.8000 465.6000 ;
	    RECT 357.0000 465.4500 358.2000 465.6000 ;
	    RECT 342.6000 464.5500 358.2000 465.4500 ;
	    RECT 342.6000 464.4000 343.8000 464.5500 ;
	    RECT 357.0000 464.4000 358.2000 464.5500 ;
	    RECT 376.2000 463.5000 377.4000 479.7000 ;
	    RECT 395.4000 473.7000 396.6000 479.7000 ;
	    RECT 397.8000 466.5000 399.0000 479.7000 ;
	    RECT 400.2000 473.7000 401.4000 479.7000 ;
	    RECT 400.2000 469.5000 401.4000 469.8000 ;
	    RECT 400.2000 467.4000 401.4000 468.6000 ;
	    RECT 424.2000 467.7000 425.4000 479.7000 ;
	    RECT 428.1000 468.6000 429.3000 479.7000 ;
	    RECT 430.5000 473.7000 431.7000 479.7000 ;
	    RECT 453.0000 473.7000 454.2000 479.7000 ;
	    RECT 430.2000 470.4000 431.4000 471.6000 ;
	    RECT 430.5000 469.5000 431.4000 470.4000 ;
	    RECT 428.1000 467.7000 429.6000 468.6000 ;
	    RECT 383.4000 465.4500 384.6000 465.6000 ;
	    RECT 397.8000 465.4500 399.0000 465.6000 ;
	    RECT 383.4000 464.5500 399.0000 465.4500 ;
	    RECT 383.4000 464.4000 384.6000 464.5500 ;
	    RECT 397.8000 464.4000 399.0000 464.5500 ;
	    RECT 426.6000 464.4000 427.8000 465.6000 ;
	    RECT 304.2000 461.5500 326.8500 462.4500 ;
	    RECT 304.2000 461.4000 305.4000 461.5500 ;
	    RECT 328.2000 461.4000 329.4000 462.6000 ;
	    RECT 172.2000 459.0000 173.7000 460.2000 ;
	    RECT 172.2000 453.3000 173.4000 459.0000 ;
	    RECT 196.2000 456.3000 197.1000 460.5000 ;
	    RECT 198.6000 458.4000 199.8000 459.6000 ;
	    RECT 213.0000 459.4500 214.2000 459.6000 ;
	    RECT 220.2000 459.4500 221.4000 459.6000 ;
	    RECT 213.0000 458.5500 221.4000 459.4500 ;
	    RECT 213.0000 458.4000 214.2000 458.5500 ;
	    RECT 220.2000 458.4000 221.4000 458.5500 ;
	    RECT 198.6000 457.2000 199.8000 457.5000 ;
	    RECT 220.2000 457.2000 221.4000 457.5000 ;
	    RECT 174.6000 453.3000 175.8000 456.3000 ;
	    RECT 193.8000 453.3000 195.0000 456.3000 ;
	    RECT 196.2000 453.3000 197.4000 456.3000 ;
	    RECT 198.6000 453.3000 199.8000 456.3000 ;
	    RECT 220.2000 453.3000 221.4000 456.3000 ;
	    RECT 222.6000 453.3000 223.8000 460.5000 ;
	    RECT 254.1000 459.3000 259.5000 459.9000 ;
	    RECT 261.3000 459.3000 262.2000 461.4000 ;
	    RECT 330.3000 460.8000 330.6000 462.3000 ;
	    RECT 332.7000 461.4000 334.5000 462.6000 ;
	    RECT 335.4000 461.4000 336.6000 462.6000 ;
	    RECT 352.2000 462.4500 353.4000 462.6000 ;
	    RECT 354.6000 462.4500 355.8000 462.6000 ;
	    RECT 352.2000 461.5500 355.8000 462.4500 ;
	    RECT 352.2000 461.4000 353.4000 461.5500 ;
	    RECT 354.6000 461.4000 355.8000 461.5500 ;
	    RECT 253.8000 459.0000 259.8000 459.3000 ;
	    RECT 253.8000 453.3000 255.0000 459.0000 ;
	    RECT 256.2000 453.3000 257.4000 458.1000 ;
	    RECT 258.6000 454.2000 259.8000 459.0000 ;
	    RECT 261.0000 455.1000 262.2000 459.3000 ;
	    RECT 263.4000 454.2000 264.6000 459.3000 ;
	    RECT 285.0000 456.3000 285.9000 460.5000 ;
	    RECT 287.4000 458.4000 288.6000 459.6000 ;
	    RECT 301.8000 458.4000 303.0000 459.6000 ;
	    RECT 287.4000 457.2000 288.6000 457.5000 ;
	    RECT 301.8000 457.2000 303.0000 457.5000 ;
	    RECT 258.6000 453.3000 264.6000 454.2000 ;
	    RECT 282.6000 453.3000 283.8000 456.3000 ;
	    RECT 285.0000 453.3000 286.2000 456.3000 ;
	    RECT 287.4000 453.3000 288.6000 456.3000 ;
	    RECT 301.8000 453.3000 303.0000 456.3000 ;
	    RECT 304.2000 453.3000 305.4000 460.5000 ;
	    RECT 328.5000 459.3000 333.9000 459.9000 ;
	    RECT 335.4000 459.3000 336.3000 460.5000 ;
	    RECT 354.6000 460.2000 355.8000 460.5000 ;
	    RECT 357.0000 459.3000 358.2000 463.5000 ;
	    RECT 376.2000 462.4500 377.4000 462.6000 ;
	    RECT 393.0000 462.4500 394.2000 462.6000 ;
	    RECT 376.2000 461.5500 394.2000 462.4500 ;
	    RECT 376.2000 461.4000 377.4000 461.5500 ;
	    RECT 393.0000 461.4000 394.2000 461.5500 ;
	    RECT 395.4000 461.4000 396.6000 462.6000 ;
	    RECT 328.2000 459.0000 334.2000 459.3000 ;
	    RECT 328.2000 453.3000 329.4000 459.0000 ;
	    RECT 330.6000 453.3000 331.8000 458.1000 ;
	    RECT 333.0000 453.3000 334.2000 459.0000 ;
	    RECT 335.4000 453.3000 336.6000 459.3000 ;
	    RECT 354.6000 453.3000 355.8000 459.3000 ;
	    RECT 357.0000 458.4000 359.7000 459.3000 ;
	    RECT 373.8000 458.4000 375.0000 459.6000 ;
	    RECT 358.5000 453.3000 359.7000 458.4000 ;
	    RECT 373.8000 457.2000 375.0000 457.5000 ;
	    RECT 373.8000 453.3000 375.0000 456.3000 ;
	    RECT 376.2000 453.3000 377.4000 460.5000 ;
	    RECT 395.4000 460.2000 396.6000 460.5000 ;
	    RECT 397.8000 459.3000 399.0000 463.5000 ;
	    RECT 426.6000 463.2000 427.8000 463.5000 ;
	    RECT 428.7000 462.6000 429.6000 467.7000 ;
	    RECT 431.4000 467.4000 432.6000 468.6000 ;
	    RECT 455.4000 463.5000 456.6000 479.7000 ;
	    RECT 467.4000 473.7000 468.6000 479.7000 ;
	    RECT 469.8000 463.5000 471.0000 479.7000 ;
	    RECT 594.6000 473.7000 595.8000 479.7000 ;
	    RECT 597.0000 474.6000 598.2000 479.7000 ;
	    RECT 596.7000 473.7000 598.2000 474.6000 ;
	    RECT 599.4000 473.7000 600.6000 480.6000 ;
	    RECT 596.7000 472.8000 597.6000 473.7000 ;
	    RECT 601.8000 472.8000 603.0000 479.7000 ;
	    RECT 604.2000 473.7000 605.4000 479.7000 ;
	    RECT 606.6000 475.5000 607.8000 479.7000 ;
	    RECT 609.0000 475.5000 610.2000 479.7000 ;
	    RECT 594.6000 471.9000 597.6000 472.8000 ;
	    RECT 594.6000 463.5000 595.8000 471.9000 ;
	    RECT 598.5000 471.6000 604.8000 472.8000 ;
	    RECT 611.4000 472.5000 612.6000 479.7000 ;
	    RECT 613.8000 473.7000 615.0000 479.7000 ;
	    RECT 616.2000 472.5000 617.4000 479.7000 ;
	    RECT 618.6000 473.7000 619.8000 479.7000 ;
	    RECT 598.5000 471.0000 599.4000 471.6000 ;
	    RECT 597.0000 469.8000 599.4000 471.0000 ;
	    RECT 603.9000 470.7000 612.6000 471.6000 ;
	    RECT 600.9000 469.8000 603.0000 470.7000 ;
	    RECT 600.9000 469.5000 610.2000 469.8000 ;
	    RECT 602.1000 468.9000 610.2000 469.5000 ;
	    RECT 609.0000 468.6000 610.2000 468.9000 ;
	    RECT 611.7000 469.5000 612.6000 470.7000 ;
	    RECT 613.5000 470.4000 617.4000 471.6000 ;
	    RECT 621.0000 470.4000 622.2000 479.7000 ;
	    RECT 623.4000 475.5000 624.6000 479.7000 ;
	    RECT 625.8000 475.5000 627.0000 479.7000 ;
	    RECT 628.2000 475.5000 629.4000 479.7000 ;
	    RECT 630.6000 473.7000 631.8000 479.7000 ;
	    RECT 625.8000 471.6000 632.1000 472.8000 ;
	    RECT 633.0000 471.6000 634.2000 479.7000 ;
	    RECT 635.4000 473.7000 636.6000 479.7000 ;
	    RECT 637.8000 472.8000 639.0000 479.7000 ;
	    RECT 640.2000 473.7000 641.4000 479.7000 ;
	    RECT 637.8000 471.9000 641.7000 472.8000 ;
	    RECT 642.6000 472.5000 643.8000 479.7000 ;
	    RECT 645.0000 473.7000 646.2000 479.7000 ;
	    RECT 657.0000 473.7000 658.2000 479.7000 ;
	    RECT 633.0000 470.4000 636.9000 471.6000 ;
	    RECT 623.4000 469.5000 624.6000 469.8000 ;
	    RECT 611.7000 468.6000 624.6000 469.5000 ;
	    RECT 628.2000 469.5000 629.4000 469.8000 ;
	    RECT 640.8000 469.5000 641.7000 471.9000 ;
	    RECT 642.6000 470.4000 643.8000 471.6000 ;
	    RECT 628.2000 468.6000 641.7000 469.5000 ;
	    RECT 599.4000 467.4000 600.6000 468.6000 ;
	    RECT 604.5000 467.7000 605.7000 468.0000 ;
	    RECT 601.5000 466.8000 639.9000 467.7000 ;
	    RECT 638.7000 466.5000 639.9000 466.8000 ;
	    RECT 640.8000 465.9000 641.7000 468.6000 ;
	    RECT 642.6000 468.0000 643.8000 469.5000 ;
	    RECT 642.6000 466.8000 644.1000 468.0000 ;
	    RECT 596.7000 465.0000 603.3000 465.9000 ;
	    RECT 596.7000 464.7000 597.9000 465.0000 ;
	    RECT 604.2000 464.4000 605.4000 465.6000 ;
	    RECT 606.3000 465.0000 631.8000 465.9000 ;
	    RECT 640.8000 465.0000 642.0000 465.9000 ;
	    RECT 630.6000 464.1000 631.8000 465.0000 ;
	    RECT 421.8000 462.4500 423.0000 462.6000 ;
	    RECT 424.2000 462.4500 425.4000 462.6000 ;
	    RECT 421.8000 461.5500 425.4000 462.4500 ;
	    RECT 421.8000 461.4000 423.0000 461.5500 ;
	    RECT 424.2000 461.4000 425.4000 461.5500 ;
	    RECT 426.3000 460.8000 426.6000 462.3000 ;
	    RECT 428.7000 461.4000 430.5000 462.6000 ;
	    RECT 431.4000 462.4500 432.6000 462.6000 ;
	    RECT 450.6000 462.4500 451.8000 462.6000 ;
	    RECT 431.4000 461.5500 451.8000 462.4500 ;
	    RECT 431.4000 461.4000 432.6000 461.5500 ;
	    RECT 450.6000 461.4000 451.8000 461.5500 ;
	    RECT 455.4000 462.4500 456.6000 462.6000 ;
	    RECT 467.4000 462.4500 468.6000 462.6000 ;
	    RECT 455.4000 461.5500 468.6000 462.4500 ;
	    RECT 455.4000 461.4000 456.6000 461.5500 ;
	    RECT 467.4000 461.4000 468.6000 461.5500 ;
	    RECT 469.8000 461.4000 471.0000 462.6000 ;
	    RECT 594.6000 462.3000 607.8000 463.5000 ;
	    RECT 608.7000 462.9000 611.7000 464.1000 ;
	    RECT 617.4000 462.9000 622.2000 464.1000 ;
	    RECT 424.5000 459.3000 429.9000 459.9000 ;
	    RECT 431.4000 459.3000 432.3000 460.5000 ;
	    RECT 395.4000 453.3000 396.6000 459.3000 ;
	    RECT 397.8000 458.4000 400.5000 459.3000 ;
	    RECT 399.3000 453.3000 400.5000 458.4000 ;
	    RECT 424.2000 459.0000 430.2000 459.3000 ;
	    RECT 424.2000 453.3000 425.4000 459.0000 ;
	    RECT 426.6000 453.3000 427.8000 458.1000 ;
	    RECT 429.0000 453.3000 430.2000 459.0000 ;
	    RECT 431.4000 453.3000 432.6000 459.3000 ;
	    RECT 453.0000 458.4000 454.2000 459.6000 ;
	    RECT 453.0000 457.2000 454.2000 457.5000 ;
	    RECT 453.0000 453.3000 454.2000 456.3000 ;
	    RECT 455.4000 453.3000 456.6000 460.5000 ;
	    RECT 467.4000 458.4000 468.6000 459.6000 ;
	    RECT 467.4000 457.2000 468.6000 457.5000 ;
	    RECT 467.4000 453.3000 468.6000 456.3000 ;
	    RECT 469.8000 453.3000 471.0000 460.5000 ;
	    RECT 594.6000 453.3000 595.8000 462.3000 ;
	    RECT 598.2000 460.2000 602.7000 461.4000 ;
	    RECT 601.5000 459.3000 602.7000 460.2000 ;
	    RECT 610.5000 459.3000 611.7000 462.9000 ;
	    RECT 613.8000 461.4000 615.0000 462.6000 ;
	    RECT 621.6000 461.7000 622.8000 462.0000 ;
	    RECT 616.2000 460.8000 622.8000 461.7000 ;
	    RECT 616.2000 460.5000 617.4000 460.8000 ;
	    RECT 613.8000 460.2000 615.0000 460.5000 ;
	    RECT 625.8000 459.6000 627.0000 463.8000 ;
	    RECT 634.5000 462.9000 640.2000 464.1000 ;
	    RECT 634.5000 461.1000 635.7000 462.9000 ;
	    RECT 641.1000 462.0000 642.0000 465.0000 ;
	    RECT 616.2000 459.3000 617.4000 459.6000 ;
	    RECT 599.4000 453.3000 600.6000 459.3000 ;
	    RECT 601.5000 458.1000 605.4000 459.3000 ;
	    RECT 610.5000 458.4000 617.4000 459.3000 ;
	    RECT 618.6000 458.4000 619.8000 459.6000 ;
	    RECT 620.7000 458.4000 621.0000 459.6000 ;
	    RECT 625.5000 458.4000 627.0000 459.6000 ;
	    RECT 633.0000 460.2000 635.7000 461.1000 ;
	    RECT 640.2000 461.1000 642.0000 462.0000 ;
	    RECT 633.0000 459.3000 634.2000 460.2000 ;
	    RECT 604.2000 453.3000 605.4000 458.1000 ;
	    RECT 630.6000 458.1000 634.2000 459.3000 ;
	    RECT 606.6000 453.3000 607.8000 457.5000 ;
	    RECT 609.0000 453.3000 610.2000 457.5000 ;
	    RECT 611.4000 453.3000 612.6000 457.5000 ;
	    RECT 613.8000 453.3000 615.0000 456.3000 ;
	    RECT 616.2000 453.3000 617.4000 457.5000 ;
	    RECT 618.6000 453.3000 619.8000 456.3000 ;
	    RECT 621.0000 453.3000 622.2000 457.5000 ;
	    RECT 623.4000 453.3000 624.6000 457.5000 ;
	    RECT 625.8000 453.3000 627.0000 457.5000 ;
	    RECT 628.2000 453.3000 629.4000 457.5000 ;
	    RECT 630.6000 453.3000 631.8000 458.1000 ;
	    RECT 635.4000 453.3000 636.6000 459.3000 ;
	    RECT 640.2000 453.3000 641.4000 461.1000 ;
	    RECT 642.9000 460.2000 644.1000 466.8000 ;
	    RECT 659.4000 463.5000 660.6000 479.7000 ;
	    RECT 693.0000 467.7000 694.2000 479.7000 ;
	    RECT 696.9000 468.6000 698.1000 479.7000 ;
	    RECT 699.3000 473.7000 700.5000 479.7000 ;
	    RECT 699.0000 470.4000 700.2000 471.6000 ;
	    RECT 699.3000 469.5000 700.2000 470.4000 ;
	    RECT 719.4000 468.6000 720.6000 479.7000 ;
	    RECT 721.8000 469.5000 723.0000 479.7000 ;
	    RECT 696.9000 467.7000 698.4000 468.6000 ;
	    RECT 695.4000 465.4500 696.6000 465.6000 ;
	    RECT 690.7500 464.5500 696.6000 465.4500 ;
	    RECT 659.4000 462.4500 660.6000 462.6000 ;
	    RECT 690.7500 462.4500 691.6500 464.5500 ;
	    RECT 695.4000 464.4000 696.6000 464.5500 ;
	    RECT 695.4000 463.2000 696.6000 463.5000 ;
	    RECT 697.5000 462.6000 698.4000 467.7000 ;
	    RECT 700.2000 467.4000 701.4000 468.6000 ;
	    RECT 719.4000 467.7000 722.7000 468.6000 ;
	    RECT 724.2000 467.7000 725.4000 479.7000 ;
	    RECT 743.4000 468.6000 744.6000 479.7000 ;
	    RECT 745.8000 469.5000 747.0000 479.7000 ;
	    RECT 743.4000 467.7000 746.7000 468.6000 ;
	    RECT 748.2000 467.7000 749.4000 479.7000 ;
	    RECT 762.6000 473.7000 763.8000 479.7000 ;
	    RECT 721.8000 466.8000 722.7000 467.7000 ;
	    RECT 721.8000 465.6000 723.6000 466.8000 ;
	    RECT 719.4000 464.4000 720.6000 465.6000 ;
	    RECT 719.4000 463.2000 720.6000 463.5000 ;
	    RECT 659.4000 461.5500 691.6500 462.4500 ;
	    RECT 659.4000 461.4000 660.6000 461.5500 ;
	    RECT 693.0000 461.4000 694.2000 462.6000 ;
	    RECT 695.1000 460.8000 695.4000 462.3000 ;
	    RECT 697.5000 461.4000 699.3000 462.6000 ;
	    RECT 700.2000 461.4000 701.4000 462.6000 ;
	    RECT 721.8000 461.1000 722.7000 465.6000 ;
	    RECT 724.5000 464.4000 725.4000 467.7000 ;
	    RECT 745.8000 466.8000 746.7000 467.7000 ;
	    RECT 745.8000 465.6000 747.6000 466.8000 ;
	    RECT 741.0000 465.4500 742.2000 465.6000 ;
	    RECT 743.4000 465.4500 744.6000 465.6000 ;
	    RECT 741.0000 464.5500 744.6000 465.4500 ;
	    RECT 741.0000 464.4000 742.2000 464.5500 ;
	    RECT 743.4000 464.4000 744.6000 464.5500 ;
	    RECT 724.2000 463.5000 725.4000 464.4000 ;
	    RECT 743.4000 463.2000 744.6000 463.5000 ;
	    RECT 724.2000 461.4000 725.4000 462.6000 ;
	    RECT 745.8000 461.1000 746.7000 465.6000 ;
	    RECT 748.5000 464.4000 749.4000 467.7000 ;
	    RECT 748.2000 463.5000 749.4000 464.4000 ;
	    RECT 765.0000 463.5000 766.2000 479.7000 ;
	    RECT 789.9000 473.7000 791.1000 479.7000 ;
	    RECT 790.2000 470.4000 791.4000 471.6000 ;
	    RECT 790.2000 469.5000 791.1000 470.4000 ;
	    RECT 792.3000 468.6000 793.5000 479.7000 ;
	    RECT 786.6000 468.4500 787.8000 468.6000 ;
	    RECT 789.0000 468.4500 790.2000 468.6000 ;
	    RECT 786.6000 467.5500 790.2000 468.4500 ;
	    RECT 786.6000 467.4000 787.8000 467.5500 ;
	    RECT 789.0000 467.4000 790.2000 467.5500 ;
	    RECT 792.0000 467.7000 793.5000 468.6000 ;
	    RECT 796.2000 467.7000 797.4000 479.7000 ;
	    RECT 801.0000 479.4000 802.2000 480.6000 ;
	    RECT 815.4000 468.6000 816.6000 479.7000 ;
	    RECT 817.8000 469.5000 819.0000 479.7000 ;
	    RECT 815.4000 467.7000 818.7000 468.6000 ;
	    RECT 820.2000 467.7000 821.4000 479.7000 ;
	    RECT 839.4000 473.7000 840.6000 479.7000 ;
	    RECT 792.0000 462.6000 792.9000 467.7000 ;
	    RECT 817.8000 466.8000 818.7000 467.7000 ;
	    RECT 817.8000 465.6000 819.6000 466.8000 ;
	    RECT 793.8000 464.4000 795.0000 465.6000 ;
	    RECT 815.4000 464.4000 816.6000 465.6000 ;
	    RECT 793.8000 463.2000 795.0000 463.5000 ;
	    RECT 815.4000 463.2000 816.6000 463.5000 ;
	    RECT 748.2000 461.4000 749.4000 462.6000 ;
	    RECT 765.0000 462.4500 766.2000 462.6000 ;
	    RECT 786.6000 462.4500 787.8000 462.6000 ;
	    RECT 765.0000 461.5500 787.8000 462.4500 ;
	    RECT 765.0000 461.4000 766.2000 461.5500 ;
	    RECT 786.6000 461.4000 787.8000 461.5500 ;
	    RECT 789.0000 461.4000 790.2000 462.6000 ;
	    RECT 791.1000 461.4000 792.9000 462.6000 ;
	    RECT 796.2000 462.4500 797.4000 462.6000 ;
	    RECT 801.0000 462.4500 802.2000 462.6000 ;
	    RECT 642.6000 459.0000 644.1000 460.2000 ;
	    RECT 642.6000 453.3000 643.8000 459.0000 ;
	    RECT 657.0000 458.4000 658.2000 459.6000 ;
	    RECT 657.0000 457.2000 658.2000 457.5000 ;
	    RECT 645.0000 453.3000 646.2000 456.3000 ;
	    RECT 657.0000 453.3000 658.2000 456.3000 ;
	    RECT 659.4000 453.3000 660.6000 460.5000 ;
	    RECT 693.3000 459.3000 698.7000 459.9000 ;
	    RECT 700.2000 459.3000 701.1000 460.5000 ;
	    RECT 719.4000 460.2000 722.7000 461.1000 ;
	    RECT 693.0000 459.0000 699.0000 459.3000 ;
	    RECT 693.0000 453.3000 694.2000 459.0000 ;
	    RECT 695.4000 453.3000 696.6000 458.1000 ;
	    RECT 697.8000 453.3000 699.0000 459.0000 ;
	    RECT 700.2000 453.3000 701.4000 459.3000 ;
	    RECT 719.4000 453.3000 720.6000 460.2000 ;
	    RECT 721.8000 453.3000 723.0000 459.3000 ;
	    RECT 724.2000 453.3000 725.4000 460.5000 ;
	    RECT 743.4000 460.2000 746.7000 461.1000 ;
	    RECT 795.0000 460.8000 795.3000 462.3000 ;
	    RECT 796.2000 461.5500 802.2000 462.4500 ;
	    RECT 796.2000 461.4000 797.4000 461.5500 ;
	    RECT 801.0000 461.4000 802.2000 461.5500 ;
	    RECT 817.8000 461.1000 818.7000 465.6000 ;
	    RECT 820.5000 464.4000 821.4000 467.7000 ;
	    RECT 841.8000 466.5000 843.0000 479.7000 ;
	    RECT 844.2000 473.7000 845.4000 479.7000 ;
	    RECT 844.2000 469.5000 845.4000 469.8000 ;
	    RECT 863.4000 468.6000 864.6000 479.7000 ;
	    RECT 865.8000 469.5000 867.0000 479.7000 ;
	    RECT 844.2000 467.4000 845.4000 468.6000 ;
	    RECT 863.4000 467.7000 866.7000 468.6000 ;
	    RECT 868.2000 467.7000 869.4000 479.7000 ;
	    RECT 889.8000 479.4000 891.0000 480.6000 ;
	    RECT 865.8000 466.8000 866.7000 467.7000 ;
	    RECT 865.8000 465.6000 867.6000 466.8000 ;
	    RECT 825.0000 465.4500 826.2000 465.6000 ;
	    RECT 841.8000 465.4500 843.0000 465.6000 ;
	    RECT 825.0000 464.5500 843.0000 465.4500 ;
	    RECT 825.0000 464.4000 826.2000 464.5500 ;
	    RECT 841.8000 464.4000 843.0000 464.5500 ;
	    RECT 863.4000 464.4000 864.6000 465.6000 ;
	    RECT 820.2000 463.5000 821.4000 464.4000 ;
	    RECT 820.2000 461.4000 821.4000 462.6000 ;
	    RECT 839.4000 461.4000 840.6000 462.6000 ;
	    RECT 743.4000 453.3000 744.6000 460.2000 ;
	    RECT 745.8000 453.3000 747.0000 459.3000 ;
	    RECT 748.2000 453.3000 749.4000 460.5000 ;
	    RECT 750.6000 459.4500 751.8000 459.6000 ;
	    RECT 762.6000 459.4500 763.8000 459.6000 ;
	    RECT 750.6000 458.5500 763.8000 459.4500 ;
	    RECT 750.6000 458.4000 751.8000 458.5500 ;
	    RECT 762.6000 458.4000 763.8000 458.5500 ;
	    RECT 762.6000 457.2000 763.8000 457.5000 ;
	    RECT 762.6000 453.3000 763.8000 456.3000 ;
	    RECT 765.0000 453.3000 766.2000 460.5000 ;
	    RECT 789.3000 459.3000 790.2000 460.5000 ;
	    RECT 815.4000 460.2000 818.7000 461.1000 ;
	    RECT 791.7000 459.3000 797.1000 459.9000 ;
	    RECT 789.0000 453.3000 790.2000 459.3000 ;
	    RECT 791.4000 459.0000 797.4000 459.3000 ;
	    RECT 791.4000 453.3000 792.6000 459.0000 ;
	    RECT 793.8000 453.3000 795.0000 458.1000 ;
	    RECT 796.2000 453.3000 797.4000 459.0000 ;
	    RECT 815.4000 453.3000 816.6000 460.2000 ;
	    RECT 817.8000 453.3000 819.0000 459.3000 ;
	    RECT 820.2000 453.3000 821.4000 460.5000 ;
	    RECT 839.4000 460.2000 840.6000 460.5000 ;
	    RECT 841.8000 459.3000 843.0000 463.5000 ;
	    RECT 863.4000 463.2000 864.6000 463.5000 ;
	    RECT 865.8000 461.1000 866.7000 465.6000 ;
	    RECT 868.5000 464.4000 869.4000 467.7000 ;
	    RECT 945.0000 467.1000 946.2000 479.7000 ;
	    RECT 947.4000 468.0000 948.6000 479.7000 ;
	    RECT 951.6000 474.6000 952.8000 479.7000 ;
	    RECT 949.8000 473.7000 952.8000 474.6000 ;
	    RECT 955.8000 473.7000 957.0000 479.7000 ;
	    RECT 958.2000 473.7000 959.4000 479.7000 ;
	    RECT 960.6000 473.7000 961.8000 479.7000 ;
	    RECT 964.5000 473.7000 966.3000 479.7000 ;
	    RECT 949.8000 472.5000 951.0000 473.7000 ;
	    RECT 958.2000 472.8000 959.1000 473.7000 ;
	    RECT 954.9000 471.9000 960.3000 472.8000 ;
	    RECT 964.2000 472.5000 965.4000 473.7000 ;
	    RECT 954.9000 471.6000 956.1000 471.9000 ;
	    RECT 959.1000 471.6000 960.3000 471.9000 ;
	    RECT 949.8000 469.5000 951.0000 469.8000 ;
	    RECT 956.7000 469.5000 957.9000 469.8000 ;
	    RECT 949.8000 468.6000 957.9000 469.5000 ;
	    RECT 958.8000 469.5000 962.1000 470.4000 ;
	    RECT 958.8000 467.7000 959.7000 469.5000 ;
	    RECT 960.9000 469.2000 962.1000 469.5000 ;
	    RECT 964.5000 469.8000 966.6000 471.0000 ;
	    RECT 964.5000 468.3000 965.4000 469.8000 ;
	    RECT 952.5000 467.1000 959.7000 467.7000 ;
	    RECT 945.0000 466.8000 959.7000 467.1000 ;
	    RECT 961.8000 467.4000 965.4000 468.3000 ;
	    RECT 969.0000 467.7000 970.2000 479.7000 ;
	    RECT 945.0000 466.5000 953.7000 466.8000 ;
	    RECT 945.0000 466.2000 953.4000 466.5000 ;
	    RECT 868.2000 463.5000 869.4000 464.4000 ;
	    RECT 948.3000 464.4000 953.7000 465.3000 ;
	    RECT 954.6000 464.4000 955.8000 465.6000 ;
	    RECT 948.3000 464.1000 949.5000 464.4000 ;
	    RECT 950.7000 462.6000 951.9000 462.9000 ;
	    RECT 961.8000 462.6000 962.7000 467.4000 ;
	    RECT 971.4000 466.8000 972.6000 479.7000 ;
	    RECT 990.6000 468.6000 991.8000 479.7000 ;
	    RECT 993.0000 469.5000 994.2000 479.7000 ;
	    RECT 990.6000 467.7000 993.9000 468.6000 ;
	    RECT 995.4000 467.7000 996.6000 479.7000 ;
	    RECT 1026.6000 478.8000 1032.6000 479.7000 ;
	    RECT 1026.6000 467.7000 1027.8000 478.8000 ;
	    RECT 1029.0000 467.7000 1030.2001 477.9000 ;
	    RECT 1031.4000 468.6000 1032.6000 478.8000 ;
	    RECT 1033.8000 469.5000 1035.0000 479.7000 ;
	    RECT 1036.2001 468.6000 1037.4000 479.7000 ;
	    RECT 1031.4000 467.7000 1037.4000 468.6000 ;
	    RECT 1055.4000 468.6000 1056.6000 479.7000 ;
	    RECT 1057.8000 469.5000 1059.0000 479.7000 ;
	    RECT 1055.4000 467.7000 1058.7001 468.6000 ;
	    RECT 1060.2001 467.7000 1061.4000 479.7000 ;
	    RECT 1091.4000 478.8000 1097.4000 479.7000 ;
	    RECT 1091.4000 467.7000 1092.6000 478.8000 ;
	    RECT 1093.8000 467.7000 1095.0000 477.9000 ;
	    RECT 1096.2001 468.6000 1097.4000 478.8000 ;
	    RECT 1098.6000 469.5000 1099.8000 479.7000 ;
	    RECT 1101.0000 468.6000 1102.2001 479.7000 ;
	    RECT 1132.2001 473.7000 1133.4000 479.7000 ;
	    RECT 1134.6000 473.7000 1135.8000 479.7000 ;
	    RECT 1096.2001 467.7000 1102.2001 468.6000 ;
	    RECT 966.3000 466.5000 972.6000 466.8000 ;
	    RECT 993.0000 466.8000 993.9000 467.7000 ;
	    RECT 966.3000 465.9000 970.5000 466.5000 ;
	    RECT 966.3000 465.6000 967.5000 465.9000 ;
	    RECT 993.0000 465.6000 994.8000 466.8000 ;
	    RECT 968.7000 464.7000 969.9000 465.0000 ;
	    RECT 964.2000 463.8000 969.9000 464.7000 ;
	    RECT 971.4000 464.4000 972.6000 465.6000 ;
	    RECT 990.6000 464.4000 991.8000 465.6000 ;
	    RECT 964.2000 463.5000 965.4000 463.8000 ;
	    RECT 868.2000 461.4000 869.4000 462.6000 ;
	    RECT 946.2000 461.4000 946.5000 462.6000 ;
	    RECT 947.4000 461.4000 948.6000 462.6000 ;
	    RECT 949.5000 461.7000 962.7000 462.6000 ;
	    RECT 863.4000 460.2000 866.7000 461.1000 ;
	    RECT 839.4000 453.3000 840.6000 459.3000 ;
	    RECT 841.8000 458.4000 844.5000 459.3000 ;
	    RECT 843.3000 453.3000 844.5000 458.4000 ;
	    RECT 863.4000 453.3000 864.6000 460.2000 ;
	    RECT 865.8000 453.3000 867.0000 459.3000 ;
	    RECT 868.2000 453.3000 869.4000 460.5000 ;
	    RECT 945.0000 453.3000 946.2000 460.5000 ;
	    RECT 947.4000 453.3000 948.6000 459.3000 ;
	    RECT 952.5000 458.4000 953.4000 461.7000 ;
	    RECT 960.9000 461.4000 962.1000 461.7000 ;
	    RECT 971.4000 460.8000 972.6000 463.5000 ;
	    RECT 990.6000 463.2000 991.8000 463.5000 ;
	    RECT 993.0000 461.1000 993.9000 465.6000 ;
	    RECT 995.7000 464.4000 996.6000 467.7000 ;
	    RECT 1029.3000 466.8000 1030.2001 467.7000 ;
	    RECT 1057.8000 466.8000 1058.7001 467.7000 ;
	    RECT 1026.6000 466.5000 1027.8000 466.8000 ;
	    RECT 1029.3000 466.5000 1032.3000 466.8000 ;
	    RECT 1029.3000 465.9000 1030.5000 466.5000 ;
	    RECT 1026.6000 464.4000 1027.8000 465.6000 ;
	    RECT 1031.4000 464.4000 1032.6000 465.6000 ;
	    RECT 1035.0000 464.7000 1035.3000 466.2000 ;
	    RECT 1057.8000 465.6000 1059.6000 466.8000 ;
	    RECT 1036.2001 464.4000 1037.4000 465.6000 ;
	    RECT 1048.2001 465.4500 1049.4000 465.6000 ;
	    RECT 1055.4000 465.4500 1056.6000 465.6000 ;
	    RECT 1048.2001 464.5500 1056.6000 465.4500 ;
	    RECT 1048.2001 464.4000 1049.4000 464.5500 ;
	    RECT 1055.4000 464.4000 1056.6000 464.5500 ;
	    RECT 995.4000 463.5000 996.6000 464.4000 ;
	    RECT 1029.3000 463.5000 1030.5000 464.4000 ;
	    RECT 1033.8000 463.5000 1035.0000 463.8000 ;
	    RECT 995.4000 462.4500 996.6000 462.6000 ;
	    RECT 1019.4000 462.4500 1020.6000 462.6000 ;
	    RECT 995.4000 461.5500 1020.6000 462.4500 ;
	    RECT 995.4000 461.4000 996.6000 461.5500 ;
	    RECT 1019.4000 461.4000 1020.6000 461.5500 ;
	    RECT 1029.0000 461.4000 1030.2001 462.6000 ;
	    RECT 966.9000 459.9000 972.6000 460.8000 ;
	    RECT 966.9000 459.6000 968.1000 459.9000 ;
	    RECT 949.8000 456.3000 951.0000 457.5000 ;
	    RECT 952.2000 457.2000 953.4000 458.4000 ;
	    RECT 954.9000 458.1000 956.1000 458.4000 ;
	    RECT 954.9000 457.2000 959.1000 458.1000 ;
	    RECT 958.2000 456.3000 959.1000 457.2000 ;
	    RECT 964.2000 456.3000 965.4000 457.5000 ;
	    RECT 949.8000 455.4000 952.8000 456.3000 ;
	    RECT 951.6000 453.3000 952.8000 455.4000 ;
	    RECT 955.5000 453.3000 957.0000 456.3000 ;
	    RECT 958.2000 453.3000 959.4000 456.3000 ;
	    RECT 960.6000 453.3000 961.8000 456.3000 ;
	    RECT 964.2000 455.4000 966.3000 456.3000 ;
	    RECT 964.5000 453.3000 966.3000 455.4000 ;
	    RECT 969.0000 453.3000 970.2000 459.0000 ;
	    RECT 971.4000 453.3000 972.6000 459.9000 ;
	    RECT 990.6000 460.2000 993.9000 461.1000 ;
	    RECT 990.6000 453.3000 991.8000 460.2000 ;
	    RECT 993.0000 453.3000 994.2000 459.3000 ;
	    RECT 995.4000 453.3000 996.6000 460.5000 ;
	    RECT 1031.4000 459.3000 1032.3000 463.5000 ;
	    RECT 1055.4000 463.2000 1056.6000 463.5000 ;
	    RECT 1033.8000 461.4000 1035.0000 462.6000 ;
	    RECT 1057.8000 461.1000 1058.7001 465.6000 ;
	    RECT 1060.5000 464.4000 1061.4000 467.7000 ;
	    RECT 1094.1000 466.8000 1095.0000 467.7000 ;
	    RECT 1134.9000 467.4000 1135.8000 473.7000 ;
	    RECT 1137.0000 468.3000 1138.2001 479.7000 ;
	    RECT 1139.4000 467.7000 1140.6000 479.7000 ;
	    RECT 1153.8000 473.7000 1155.0000 479.7000 ;
	    RECT 1091.4000 466.5000 1092.6000 466.8000 ;
	    RECT 1094.1000 466.5000 1097.1000 466.8000 ;
	    RECT 1134.9000 466.5000 1138.5000 467.4000 ;
	    RECT 1139.7001 466.5000 1140.6000 467.7000 ;
	    RECT 1094.1000 465.9000 1095.3000 466.5000 ;
	    RECT 1079.4000 465.4500 1080.6000 465.6000 ;
	    RECT 1079.4000 464.5500 1090.0500 465.4500 ;
	    RECT 1079.4000 464.4000 1080.6000 464.5500 ;
	    RECT 1060.2001 463.5000 1061.4000 464.4000 ;
	    RECT 1060.2001 462.4500 1061.4000 462.6000 ;
	    RECT 1084.2001 462.4500 1085.4000 462.6000 ;
	    RECT 1060.2001 461.5500 1085.4000 462.4500 ;
	    RECT 1089.1500 462.4500 1090.0500 464.5500 ;
	    RECT 1091.4000 464.4000 1092.6000 465.6000 ;
	    RECT 1096.2001 464.4000 1097.4000 465.6000 ;
	    RECT 1099.8000 464.7000 1100.1000 466.2000 ;
	    RECT 1101.0000 464.4000 1102.2001 465.6000 ;
	    RECT 1134.6000 464.4000 1135.8000 465.6000 ;
	    RECT 1094.1000 463.5000 1095.3000 464.4000 ;
	    RECT 1098.6000 463.5000 1099.8000 463.8000 ;
	    RECT 1132.2001 463.5000 1133.4000 463.8000 ;
	    RECT 1093.8000 462.4500 1095.0000 462.6000 ;
	    RECT 1089.1500 461.5500 1095.0000 462.4500 ;
	    RECT 1060.2001 461.4000 1061.4000 461.5500 ;
	    RECT 1084.2001 461.4000 1085.4000 461.5500 ;
	    RECT 1093.8000 461.4000 1095.0000 461.5500 ;
	    RECT 1055.4000 460.2000 1058.7001 461.1000 ;
	    RECT 1026.6000 453.3000 1027.8000 459.3000 ;
	    RECT 1030.5000 453.3000 1032.9000 459.3000 ;
	    RECT 1035.6000 453.3000 1036.8000 459.3000 ;
	    RECT 1055.4000 453.3000 1056.6000 460.2000 ;
	    RECT 1057.8000 453.3000 1059.0000 459.3000 ;
	    RECT 1060.2001 453.3000 1061.4000 460.5000 ;
	    RECT 1096.2001 459.3000 1097.1000 463.5000 ;
	    RECT 1134.9000 463.2000 1135.8000 463.5000 ;
	    RECT 1098.6000 461.4000 1099.8000 462.6000 ;
	    RECT 1132.2001 461.4000 1133.4000 462.6000 ;
	    RECT 1134.9000 462.3000 1136.4000 463.2000 ;
	    RECT 1135.2001 462.0000 1136.4000 462.3000 ;
	    RECT 1137.6000 461.4000 1138.5000 466.5000 ;
	    RECT 1139.4000 465.4500 1140.6000 465.6000 ;
	    RECT 1153.8000 465.4500 1155.0000 465.6000 ;
	    RECT 1139.4000 464.5500 1155.0000 465.4500 ;
	    RECT 1139.4000 464.4000 1140.6000 464.5500 ;
	    RECT 1153.8000 464.4000 1155.0000 464.5500 ;
	    RECT 1156.2001 463.5000 1157.4000 479.7000 ;
	    RECT 1180.2001 473.7000 1181.4000 479.7000 ;
	    RECT 1182.6000 473.7000 1183.8000 479.7000 ;
	    RECT 1185.0000 474.3000 1186.2001 479.7000 ;
	    RECT 1182.9000 473.4000 1183.8000 473.7000 ;
	    RECT 1187.4000 473.7000 1188.6000 479.7000 ;
	    RECT 1206.6000 473.7000 1207.8000 479.7000 ;
	    RECT 1187.4000 473.4000 1188.3000 473.7000 ;
	    RECT 1182.9000 472.5000 1188.3000 473.4000 ;
	    RECT 1161.0000 471.4500 1162.2001 471.6000 ;
	    RECT 1182.6000 471.4500 1183.8000 471.6000 ;
	    RECT 1161.0000 470.5500 1183.8000 471.4500 ;
	    RECT 1161.0000 470.4000 1162.2001 470.5500 ;
	    RECT 1182.6000 470.4000 1183.8000 470.5500 ;
	    RECT 1185.0000 470.4000 1186.2001 471.6000 ;
	    RECT 1187.4000 469.5000 1188.3000 472.5000 ;
	    RECT 1206.6000 469.5000 1207.8000 469.8000 ;
	    RECT 1185.0000 469.2000 1186.2001 469.5000 ;
	    RECT 1165.8000 468.4500 1167.0000 468.6000 ;
	    RECT 1180.2001 468.4500 1181.4000 468.6000 ;
	    RECT 1165.8000 467.5500 1181.4000 468.4500 ;
	    RECT 1165.8000 467.4000 1167.0000 467.5500 ;
	    RECT 1180.2001 467.4000 1181.4000 467.5500 ;
	    RECT 1187.4000 468.4500 1188.6000 468.6000 ;
	    RECT 1197.0000 468.4500 1198.2001 468.6000 ;
	    RECT 1187.4000 467.5500 1198.2001 468.4500 ;
	    RECT 1187.4000 467.4000 1188.6000 467.5500 ;
	    RECT 1197.0000 467.4000 1198.2001 467.5500 ;
	    RECT 1199.4000 468.4500 1200.6000 468.6000 ;
	    RECT 1206.6000 468.4500 1207.8000 468.6000 ;
	    RECT 1199.4000 467.5500 1207.8000 468.4500 ;
	    RECT 1199.4000 467.4000 1200.6000 467.5500 ;
	    RECT 1206.6000 467.4000 1207.8000 467.5500 ;
	    RECT 1209.0000 466.5000 1210.2001 479.7000 ;
	    RECT 1211.4000 473.7000 1212.6000 479.7000 ;
	    RECT 1236.3000 473.7000 1237.5000 479.7000 ;
	    RECT 1236.6000 470.4000 1237.8000 471.6000 ;
	    RECT 1236.6000 469.5000 1237.5000 470.4000 ;
	    RECT 1238.7001 468.6000 1239.9000 479.7000 ;
	    RECT 1235.4000 467.4000 1236.6000 468.6000 ;
	    RECT 1238.4000 467.7000 1239.9000 468.6000 ;
	    RECT 1242.6000 467.7000 1243.8000 479.7000 ;
	    RECT 1266.6000 468.6000 1267.8000 479.7000 ;
	    RECT 1269.0000 469.5000 1270.2001 479.7000 ;
	    RECT 1271.4000 468.6000 1272.6000 479.7000 ;
	    RECT 1266.6000 467.7000 1272.6000 468.6000 ;
	    RECT 1273.8000 467.7000 1275.0000 479.7000 ;
	    RECT 1300.2001 473.7000 1301.4000 479.7000 ;
	    RECT 1302.6000 473.7000 1303.8000 479.7000 ;
	    RECT 1305.0000 474.3000 1306.2001 479.7000 ;
	    RECT 1302.9000 473.4000 1303.8000 473.7000 ;
	    RECT 1307.4000 473.7000 1308.6000 479.7000 ;
	    RECT 1333.8000 473.7000 1335.0000 479.7000 ;
	    RECT 1336.2001 473.7000 1337.4000 479.7000 ;
	    RECT 1338.6000 474.3000 1339.8000 479.7000 ;
	    RECT 1307.4000 473.4000 1308.3000 473.7000 ;
	    RECT 1302.9000 472.5000 1308.3000 473.4000 ;
	    RECT 1336.5000 473.4000 1337.4000 473.7000 ;
	    RECT 1341.0000 473.7000 1342.2001 479.7000 ;
	    RECT 1341.0000 473.4000 1341.9000 473.7000 ;
	    RECT 1336.5000 472.5000 1341.9000 473.4000 ;
	    RECT 1305.0000 470.4000 1306.2001 471.6000 ;
	    RECT 1307.4000 469.5000 1308.3000 472.5000 ;
	    RECT 1319.4000 471.4500 1320.6000 471.6000 ;
	    RECT 1338.6000 471.4500 1339.8000 471.6000 ;
	    RECT 1319.4000 470.5500 1339.8000 471.4500 ;
	    RECT 1319.4000 470.4000 1320.6000 470.5500 ;
	    RECT 1338.6000 470.4000 1339.8000 470.5500 ;
	    RECT 1341.0000 469.5000 1341.9000 472.5000 ;
	    RECT 1305.0000 469.2000 1306.2001 469.5000 ;
	    RECT 1338.6000 469.2000 1339.8000 469.5000 ;
	    RECT 1288.2001 468.4500 1289.4000 468.6000 ;
	    RECT 1300.2001 468.4500 1301.4000 468.6000 ;
	    RECT 1180.2001 466.2000 1181.4000 466.5000 ;
	    RECT 1182.6000 464.4000 1183.8000 465.6000 ;
	    RECT 1184.7001 464.4000 1185.0000 465.6000 ;
	    RECT 1137.6000 461.1000 1138.8000 461.4000 ;
	    RECT 1134.3000 460.5000 1138.8000 461.1000 ;
	    RECT 1132.5000 460.2000 1138.8000 460.5000 ;
	    RECT 1132.5000 459.6000 1135.2001 460.2000 ;
	    RECT 1132.5000 459.3000 1133.4000 459.6000 ;
	    RECT 1139.7001 459.3000 1140.6000 463.5000 ;
	    RECT 1187.4000 462.6000 1188.3000 466.5000 ;
	    RECT 1209.0000 465.4500 1210.2001 465.6000 ;
	    RECT 1235.5500 465.4500 1236.4501 467.4000 ;
	    RECT 1209.0000 464.5500 1236.4501 465.4500 ;
	    RECT 1209.0000 464.4000 1210.2001 464.5500 ;
	    RECT 1156.2001 462.4500 1157.4000 462.6000 ;
	    RECT 1177.8000 462.4500 1179.0000 462.6000 ;
	    RECT 1156.2001 461.5500 1179.0000 462.4500 ;
	    RECT 1185.9000 462.3000 1188.3000 462.6000 ;
	    RECT 1156.2001 461.4000 1157.4000 461.5500 ;
	    RECT 1177.8000 461.4000 1179.0000 461.5500 ;
	    RECT 1091.4000 453.3000 1092.6000 459.3000 ;
	    RECT 1095.3000 453.3000 1097.7001 459.3000 ;
	    RECT 1100.4000 453.3000 1101.6000 459.3000 ;
	    RECT 1132.2001 453.3000 1133.4000 459.3000 ;
	    RECT 1136.1000 453.3000 1137.3000 459.0000 ;
	    RECT 1138.5000 457.8000 1140.6000 459.3000 ;
	    RECT 1141.8000 459.4500 1143.0000 459.6000 ;
	    RECT 1153.8000 459.4500 1155.0000 459.6000 ;
	    RECT 1141.8000 458.5500 1155.0000 459.4500 ;
	    RECT 1141.8000 458.4000 1143.0000 458.5500 ;
	    RECT 1153.8000 458.4000 1155.0000 458.5500 ;
	    RECT 1138.5000 453.3000 1139.7001 457.8000 ;
	    RECT 1153.8000 457.2000 1155.0000 457.5000 ;
	    RECT 1153.8000 453.3000 1155.0000 456.3000 ;
	    RECT 1156.2001 453.3000 1157.4000 460.5000 ;
	    RECT 1180.2001 453.3000 1181.4000 462.3000 ;
	    RECT 1185.6000 461.7000 1188.3000 462.3000 ;
	    RECT 1185.6000 453.3000 1186.8000 461.7000 ;
	    RECT 1209.0000 459.3000 1210.2001 463.5000 ;
	    RECT 1238.4000 462.6000 1239.3000 467.7000 ;
	    RECT 1273.8000 466.5000 1274.7001 467.7000 ;
	    RECT 1288.2001 467.5500 1301.4000 468.4500 ;
	    RECT 1288.2001 467.4000 1289.4000 467.5500 ;
	    RECT 1300.2001 467.4000 1301.4000 467.5500 ;
	    RECT 1307.4000 468.4500 1308.6000 468.6000 ;
	    RECT 1312.2001 468.4500 1313.4000 468.6000 ;
	    RECT 1307.4000 467.5500 1313.4000 468.4500 ;
	    RECT 1307.4000 467.4000 1308.6000 467.5500 ;
	    RECT 1312.2001 467.4000 1313.4000 467.5500 ;
	    RECT 1314.6000 468.4500 1315.8000 468.6000 ;
	    RECT 1329.0000 468.4500 1330.2001 468.6000 ;
	    RECT 1333.8000 468.4500 1335.0000 468.6000 ;
	    RECT 1314.6000 467.5500 1335.0000 468.4500 ;
	    RECT 1314.6000 467.4000 1315.8000 467.5500 ;
	    RECT 1329.0000 467.4000 1330.2001 467.5500 ;
	    RECT 1333.8000 467.4000 1335.0000 467.5500 ;
	    RECT 1341.0000 468.4500 1342.2001 468.6000 ;
	    RECT 1348.2001 468.4500 1349.4000 468.6000 ;
	    RECT 1341.0000 467.5500 1349.4000 468.4500 ;
	    RECT 1341.0000 467.4000 1342.2001 467.5500 ;
	    RECT 1348.2001 467.4000 1349.4000 467.5500 ;
	    RECT 1300.2001 466.2000 1301.4000 466.5000 ;
	    RECT 1240.2001 464.4000 1241.4000 465.6000 ;
	    RECT 1266.6000 464.4000 1267.8000 465.6000 ;
	    RECT 1268.7001 464.7000 1269.0000 466.2000 ;
	    RECT 1271.4000 464.7000 1272.9000 465.6000 ;
	    RECT 1273.8000 465.4500 1275.0000 465.6000 ;
	    RECT 1285.8000 465.4500 1287.0000 465.6000 ;
	    RECT 1269.0000 463.5000 1270.2001 463.8000 ;
	    RECT 1240.2001 463.2000 1241.4000 463.5000 ;
	    RECT 1211.4000 461.4000 1212.6000 462.6000 ;
	    RECT 1235.4000 461.4000 1236.6000 462.6000 ;
	    RECT 1237.5000 461.4000 1239.3000 462.6000 ;
	    RECT 1242.6000 462.4500 1243.8000 462.6000 ;
	    RECT 1259.4000 462.4500 1260.6000 462.6000 ;
	    RECT 1241.4000 460.8000 1241.7001 462.3000 ;
	    RECT 1242.6000 461.5500 1260.6000 462.4500 ;
	    RECT 1242.6000 461.4000 1243.8000 461.5500 ;
	    RECT 1259.4000 461.4000 1260.6000 461.5500 ;
	    RECT 1269.0000 461.4000 1270.2001 462.6000 ;
	    RECT 1211.4000 460.2000 1212.6000 460.5000 ;
	    RECT 1235.7001 459.3000 1236.6000 460.5000 ;
	    RECT 1238.1000 459.3000 1243.5000 459.9000 ;
	    RECT 1271.4000 459.3000 1272.3000 464.7000 ;
	    RECT 1273.8000 464.5500 1287.0000 465.4500 ;
	    RECT 1273.8000 464.4000 1275.0000 464.5500 ;
	    RECT 1285.8000 464.4000 1287.0000 464.5500 ;
	    RECT 1302.6000 464.4000 1303.8000 465.6000 ;
	    RECT 1304.7001 464.4000 1305.0000 465.6000 ;
	    RECT 1307.4000 462.6000 1308.3000 466.5000 ;
	    RECT 1333.8000 466.2000 1335.0000 466.5000 ;
	    RECT 1336.2001 464.4000 1337.4000 465.6000 ;
	    RECT 1338.3000 464.4000 1338.6000 465.6000 ;
	    RECT 1341.0000 462.6000 1341.9000 466.5000 ;
	    RECT 1353.0000 463.5000 1354.2001 479.7000 ;
	    RECT 1355.4000 473.7000 1356.6000 479.7000 ;
	    RECT 1386.6000 473.7000 1387.8000 479.7000 ;
	    RECT 1389.0000 474.3000 1390.2001 479.7000 ;
	    RECT 1386.9000 473.4000 1387.8000 473.7000 ;
	    RECT 1391.4000 473.7000 1392.6000 479.7000 ;
	    RECT 1393.8000 473.7000 1395.0000 479.7000 ;
	    RECT 1417.8000 473.7000 1419.0000 479.7000 ;
	    RECT 1420.2001 473.7000 1421.4000 479.7000 ;
	    RECT 1422.6000 474.3000 1423.8000 479.7000 ;
	    RECT 1391.4000 473.4000 1392.3000 473.7000 ;
	    RECT 1386.9000 472.5000 1392.3000 473.4000 ;
	    RECT 1420.5000 473.4000 1421.4000 473.7000 ;
	    RECT 1425.0000 473.7000 1426.2001 479.7000 ;
	    RECT 1449.0000 473.7000 1450.2001 479.7000 ;
	    RECT 1451.4000 473.7000 1452.6000 479.7000 ;
	    RECT 1453.8000 474.3000 1455.0000 479.7000 ;
	    RECT 1425.0000 473.4000 1425.9000 473.7000 ;
	    RECT 1420.5000 472.5000 1425.9000 473.4000 ;
	    RECT 1451.7001 473.4000 1452.6000 473.7000 ;
	    RECT 1456.2001 473.7000 1457.4000 479.7000 ;
	    RECT 1480.2001 473.7000 1481.4000 479.7000 ;
	    RECT 1482.6000 473.7000 1483.8000 479.7000 ;
	    RECT 1485.0000 474.3000 1486.2001 479.7000 ;
	    RECT 1456.2001 473.4000 1457.1000 473.7000 ;
	    RECT 1451.7001 472.5000 1457.1000 473.4000 ;
	    RECT 1482.9000 473.4000 1483.8000 473.7000 ;
	    RECT 1487.4000 473.7000 1488.6000 479.7000 ;
	    RECT 1506.6000 473.7000 1507.8000 479.7000 ;
	    RECT 1487.4000 473.4000 1488.3000 473.7000 ;
	    RECT 1482.9000 472.5000 1488.3000 473.4000 ;
	    RECT 1386.9000 469.5000 1387.8000 472.5000 ;
	    RECT 1389.0000 471.4500 1390.2001 471.6000 ;
	    RECT 1422.6000 471.4500 1423.8000 471.6000 ;
	    RECT 1389.0000 470.5500 1423.8000 471.4500 ;
	    RECT 1389.0000 470.4000 1390.2001 470.5500 ;
	    RECT 1422.6000 470.4000 1423.8000 470.5500 ;
	    RECT 1425.0000 469.5000 1425.9000 472.5000 ;
	    RECT 1446.6000 471.4500 1447.8000 471.6000 ;
	    RECT 1446.6000 470.5500 1452.4501 471.4500 ;
	    RECT 1446.6000 470.4000 1447.8000 470.5500 ;
	    RECT 1389.0000 469.2000 1390.2001 469.5000 ;
	    RECT 1422.6000 469.2000 1423.8000 469.5000 ;
	    RECT 1386.6000 467.4000 1387.8000 468.6000 ;
	    RECT 1393.8000 468.4500 1395.0000 468.6000 ;
	    RECT 1415.4000 468.4500 1416.6000 468.6000 ;
	    RECT 1393.8000 467.5500 1416.6000 468.4500 ;
	    RECT 1393.8000 467.4000 1395.0000 467.5500 ;
	    RECT 1415.4000 467.4000 1416.6000 467.5500 ;
	    RECT 1417.8000 467.4000 1419.0000 468.6000 ;
	    RECT 1425.0000 467.4000 1426.2001 468.6000 ;
	    RECT 1449.0000 467.4000 1450.2001 468.6000 ;
	    RECT 1386.9000 462.6000 1387.8000 466.5000 ;
	    RECT 1393.8000 466.2000 1395.0000 466.5000 ;
	    RECT 1417.8000 466.2000 1419.0000 466.5000 ;
	    RECT 1390.2001 464.4000 1390.5000 465.6000 ;
	    RECT 1391.4000 464.4000 1392.6000 465.6000 ;
	    RECT 1420.2001 464.4000 1421.4000 465.6000 ;
	    RECT 1422.3000 464.4000 1422.6000 465.6000 ;
	    RECT 1425.0000 462.6000 1425.9000 466.5000 ;
	    RECT 1449.0000 466.2000 1450.2001 466.5000 ;
	    RECT 1451.5500 465.6000 1452.4501 470.5500 ;
	    RECT 1453.8000 470.4000 1455.0000 471.6000 ;
	    RECT 1456.2001 469.5000 1457.1000 472.5000 ;
	    RECT 1485.0000 470.4000 1486.2001 471.6000 ;
	    RECT 1487.4000 469.5000 1488.3000 472.5000 ;
	    RECT 1453.8000 469.2000 1455.0000 469.5000 ;
	    RECT 1485.0000 469.2000 1486.2001 469.5000 ;
	    RECT 1456.2001 468.4500 1457.4000 468.6000 ;
	    RECT 1477.8000 468.4500 1479.0000 468.6000 ;
	    RECT 1456.2001 467.5500 1479.0000 468.4500 ;
	    RECT 1456.2001 467.4000 1457.4000 467.5500 ;
	    RECT 1477.8000 467.4000 1479.0000 467.5500 ;
	    RECT 1480.2001 467.4000 1481.4000 468.6000 ;
	    RECT 1487.4000 468.4500 1488.6000 468.6000 ;
	    RECT 1506.6000 468.4500 1507.8000 468.6000 ;
	    RECT 1487.4000 467.5500 1507.8000 468.4500 ;
	    RECT 1487.4000 467.4000 1488.6000 467.5500 ;
	    RECT 1506.6000 467.4000 1507.8000 467.5500 ;
	    RECT 1509.0000 466.5000 1510.2001 479.7000 ;
	    RECT 1511.4000 473.7000 1512.6000 479.7000 ;
	    RECT 1535.4000 473.7000 1536.6000 479.7000 ;
	    RECT 1537.8000 474.3000 1539.0000 479.7000 ;
	    RECT 1535.7001 473.4000 1536.6000 473.7000 ;
	    RECT 1540.2001 473.7000 1541.4000 479.7000 ;
	    RECT 1542.6000 473.7000 1543.8000 479.7000 ;
	    RECT 1554.6000 473.7000 1555.8000 479.7000 ;
	    RECT 1540.2001 473.4000 1541.1000 473.7000 ;
	    RECT 1535.7001 472.5000 1541.1000 473.4000 ;
	    RECT 1511.4000 469.5000 1512.6000 469.8000 ;
	    RECT 1535.7001 469.5000 1536.6000 472.5000 ;
	    RECT 1537.8000 471.4500 1539.0000 471.6000 ;
	    RECT 1545.0000 471.4500 1546.2001 471.6000 ;
	    RECT 1549.8000 471.4500 1551.0000 471.6000 ;
	    RECT 1537.8000 470.5500 1551.0000 471.4500 ;
	    RECT 1537.8000 470.4000 1539.0000 470.5500 ;
	    RECT 1545.0000 470.4000 1546.2001 470.5500 ;
	    RECT 1549.8000 470.4000 1551.0000 470.5500 ;
	    RECT 1537.8000 469.2000 1539.0000 469.5000 ;
	    RECT 1511.4000 468.4500 1512.6000 468.6000 ;
	    RECT 1535.4000 468.4500 1536.6000 468.6000 ;
	    RECT 1511.4000 467.5500 1536.6000 468.4500 ;
	    RECT 1511.4000 467.4000 1512.6000 467.5500 ;
	    RECT 1535.4000 467.4000 1536.6000 467.5500 ;
	    RECT 1542.6000 467.4000 1543.8000 468.6000 ;
	    RECT 1451.4000 464.4000 1452.6000 465.6000 ;
	    RECT 1453.5000 464.4000 1453.8000 465.6000 ;
	    RECT 1456.2001 462.6000 1457.1000 466.5000 ;
	    RECT 1480.2001 466.2000 1481.4000 466.5000 ;
	    RECT 1482.6000 464.4000 1483.8000 465.6000 ;
	    RECT 1484.7001 464.4000 1485.0000 465.6000 ;
	    RECT 1487.4000 462.6000 1488.3000 466.5000 ;
	    RECT 1501.8000 465.4500 1503.0000 465.6000 ;
	    RECT 1509.0000 465.4500 1510.2001 465.6000 ;
	    RECT 1501.8000 464.5500 1510.2001 465.4500 ;
	    RECT 1501.8000 464.4000 1503.0000 464.5500 ;
	    RECT 1509.0000 464.4000 1510.2001 464.5500 ;
	    RECT 1305.9000 462.3000 1308.3000 462.6000 ;
	    RECT 1339.5000 462.3000 1341.9000 462.6000 ;
	    RECT 1207.5000 458.4000 1210.2001 459.3000 ;
	    RECT 1207.5000 453.3000 1208.7001 458.4000 ;
	    RECT 1211.4000 453.3000 1212.6000 459.3000 ;
	    RECT 1235.4000 453.3000 1236.6000 459.3000 ;
	    RECT 1237.8000 459.0000 1243.8000 459.3000 ;
	    RECT 1237.8000 453.3000 1239.0000 459.0000 ;
	    RECT 1240.2001 453.3000 1241.4000 458.1000 ;
	    RECT 1242.6000 453.3000 1243.8000 459.0000 ;
	    RECT 1267.5000 453.3000 1268.7001 459.3000 ;
	    RECT 1271.4000 453.3000 1272.6000 459.3000 ;
	    RECT 1273.8000 458.4000 1275.0000 459.6000 ;
	    RECT 1273.5000 457.2000 1274.7001 457.5000 ;
	    RECT 1273.8000 453.3000 1275.0000 456.3000 ;
	    RECT 1300.2001 453.3000 1301.4000 462.3000 ;
	    RECT 1305.6000 461.7000 1308.3000 462.3000 ;
	    RECT 1305.6000 453.3000 1306.8000 461.7000 ;
	    RECT 1333.8000 453.3000 1335.0000 462.3000 ;
	    RECT 1339.2001 461.7000 1341.9000 462.3000 ;
	    RECT 1353.0000 462.4500 1354.2001 462.6000 ;
	    RECT 1384.2001 462.4500 1385.4000 462.6000 ;
	    RECT 1339.2001 453.3000 1340.4000 461.7000 ;
	    RECT 1353.0000 461.5500 1385.4000 462.4500 ;
	    RECT 1386.9000 462.3000 1389.3000 462.6000 ;
	    RECT 1423.5000 462.3000 1425.9000 462.6000 ;
	    RECT 1454.7001 462.3000 1457.1000 462.6000 ;
	    RECT 1485.9000 462.3000 1488.3000 462.6000 ;
	    RECT 1386.9000 461.7000 1389.6000 462.3000 ;
	    RECT 1353.0000 461.4000 1354.2001 461.5500 ;
	    RECT 1384.2001 461.4000 1385.4000 461.5500 ;
	    RECT 1353.0000 453.3000 1354.2001 460.5000 ;
	    RECT 1355.4000 459.4500 1356.6000 459.6000 ;
	    RECT 1367.4000 459.4500 1368.6000 459.6000 ;
	    RECT 1355.4000 458.5500 1368.6000 459.4500 ;
	    RECT 1355.4000 458.4000 1356.6000 458.5500 ;
	    RECT 1367.4000 458.4000 1368.6000 458.5500 ;
	    RECT 1355.4000 457.2000 1356.6000 457.5000 ;
	    RECT 1355.4000 453.3000 1356.6000 456.3000 ;
	    RECT 1388.4000 453.3000 1389.6000 461.7000 ;
	    RECT 1393.8000 453.3000 1395.0000 462.3000 ;
	    RECT 1417.8000 453.3000 1419.0000 462.3000 ;
	    RECT 1423.2001 461.7000 1425.9000 462.3000 ;
	    RECT 1423.2001 453.3000 1424.4000 461.7000 ;
	    RECT 1449.0000 453.3000 1450.2001 462.3000 ;
	    RECT 1454.4000 461.7000 1457.1000 462.3000 ;
	    RECT 1454.4000 453.3000 1455.6000 461.7000 ;
	    RECT 1480.2001 453.3000 1481.4000 462.3000 ;
	    RECT 1485.6000 461.7000 1488.3000 462.3000 ;
	    RECT 1485.6000 453.3000 1486.8000 461.7000 ;
	    RECT 1506.6000 461.4000 1507.8000 462.6000 ;
	    RECT 1506.6000 460.2000 1507.8000 460.5000 ;
	    RECT 1509.0000 459.3000 1510.2001 463.5000 ;
	    RECT 1535.7001 462.6000 1536.6000 466.5000 ;
	    RECT 1542.6000 466.2000 1543.8000 466.5000 ;
	    RECT 1539.0000 464.4000 1539.3000 465.6000 ;
	    RECT 1540.2001 464.4000 1541.4000 465.6000 ;
	    RECT 1557.0000 463.5000 1558.2001 479.7000 ;
	    RECT 1535.7001 462.3000 1538.1000 462.6000 ;
	    RECT 1535.7001 461.7000 1538.4000 462.3000 ;
	    RECT 1506.6000 453.3000 1507.8000 459.3000 ;
	    RECT 1509.0000 458.4000 1511.7001 459.3000 ;
	    RECT 1510.5000 453.3000 1511.7001 458.4000 ;
	    RECT 1537.2001 453.3000 1538.4000 461.7000 ;
	    RECT 1542.6000 453.3000 1543.8000 462.3000 ;
	    RECT 1557.0000 461.4000 1558.2001 462.6000 ;
	    RECT 1554.6000 458.4000 1555.8000 459.6000 ;
	    RECT 1554.6000 457.2000 1555.8000 457.5000 ;
	    RECT 1554.6000 453.3000 1555.8000 456.3000 ;
	    RECT 1557.0000 453.3000 1558.2001 460.5000 ;
	    RECT 1.2000 450.6000 1569.0000 452.4000 ;
	    RECT 13.8000 446.7000 15.0000 449.7000 ;
	    RECT 13.8000 445.5000 15.0000 445.8000 ;
	    RECT 13.8000 443.4000 15.0000 444.6000 ;
	    RECT 16.2000 442.5000 17.4000 449.7000 ;
	    RECT 36.3000 444.6000 37.5000 449.7000 ;
	    RECT 36.3000 443.7000 39.0000 444.6000 ;
	    RECT 40.2000 443.7000 41.4000 449.7000 ;
	    RECT 64.2000 444.0000 65.4000 449.7000 ;
	    RECT 66.6000 444.9000 67.8000 449.7000 ;
	    RECT 69.0000 444.0000 70.2000 449.7000 ;
	    RECT 64.2000 443.7000 70.2000 444.0000 ;
	    RECT 71.4000 443.7000 72.6000 449.7000 ;
	    RECT 90.6000 443.7000 91.8000 449.7000 ;
	    RECT 94.5000 444.6000 95.7000 449.7000 ;
	    RECT 93.0000 443.7000 95.7000 444.6000 ;
	    RECT 126.6000 448.8000 132.6000 449.7000 ;
	    RECT 126.6000 443.7000 127.8000 448.8000 ;
	    RECT 129.0000 443.7000 130.2000 447.9000 ;
	    RECT 131.4000 444.0000 132.6000 448.8000 ;
	    RECT 133.8000 444.9000 135.0000 449.7000 ;
	    RECT 136.2000 444.0000 137.4000 449.7000 ;
	    RECT 131.4000 443.7000 137.4000 444.0000 ;
	    RECT 165.0000 448.8000 171.0000 449.7000 ;
	    RECT 165.0000 443.7000 166.2000 448.8000 ;
	    RECT 167.4000 443.7000 168.6000 447.9000 ;
	    RECT 169.8000 444.0000 171.0000 448.8000 ;
	    RECT 172.2000 444.9000 173.4000 449.7000 ;
	    RECT 174.6000 444.0000 175.8000 449.7000 ;
	    RECT 169.8000 443.7000 175.8000 444.0000 ;
	    RECT 213.0000 444.0000 214.2000 449.7000 ;
	    RECT 215.4000 444.9000 216.6000 449.7000 ;
	    RECT 217.8000 448.8000 223.8000 449.7000 ;
	    RECT 217.8000 444.0000 219.0000 448.8000 ;
	    RECT 213.0000 443.7000 219.0000 444.0000 ;
	    RECT 220.2000 443.7000 221.4000 447.9000 ;
	    RECT 222.6000 443.7000 223.8000 448.8000 ;
	    RECT 234.6000 446.7000 235.8000 449.7000 ;
	    RECT 234.6000 445.5000 235.8000 445.8000 ;
	    RECT 232.2000 444.4500 233.4000 444.6000 ;
	    RECT 234.6000 444.4500 235.8000 444.6000 ;
	    RECT 16.2000 441.4500 17.4000 441.6000 ;
	    RECT 35.4000 441.4500 36.6000 441.6000 ;
	    RECT 16.2000 440.5500 36.6000 441.4500 ;
	    RECT 16.2000 440.4000 17.4000 440.5500 ;
	    RECT 35.4000 440.4000 36.6000 440.5500 ;
	    RECT 37.8000 439.5000 39.0000 443.7000 ;
	    RECT 64.5000 443.1000 69.9000 443.7000 ;
	    RECT 40.2000 442.5000 41.4000 442.8000 ;
	    RECT 71.4000 442.5000 72.3000 443.7000 ;
	    RECT 90.6000 442.5000 91.8000 442.8000 ;
	    RECT 40.2000 440.4000 41.4000 441.6000 ;
	    RECT 64.2000 440.4000 65.4000 441.6000 ;
	    RECT 66.3000 440.7000 66.6000 442.2000 ;
	    RECT 68.7000 440.4000 70.5000 441.6000 ;
	    RECT 71.4000 441.4500 72.6000 441.6000 ;
	    RECT 85.8000 441.4500 87.0000 441.6000 ;
	    RECT 71.4000 440.5500 87.0000 441.4500 ;
	    RECT 71.4000 440.4000 72.6000 440.5500 ;
	    RECT 85.8000 440.4000 87.0000 440.5500 ;
	    RECT 88.2000 441.4500 89.4000 441.6000 ;
	    RECT 90.6000 441.4500 91.8000 441.6000 ;
	    RECT 88.2000 440.5500 91.8000 441.4500 ;
	    RECT 88.2000 440.4000 89.4000 440.5500 ;
	    RECT 90.6000 440.4000 91.8000 440.5500 ;
	    RECT 66.6000 439.5000 67.8000 439.8000 ;
	    RECT 13.8000 423.3000 15.0000 429.3000 ;
	    RECT 16.2000 423.3000 17.4000 439.5000 ;
	    RECT 37.8000 438.4500 39.0000 438.6000 ;
	    RECT 45.0000 438.4500 46.2000 438.6000 ;
	    RECT 37.8000 437.5500 46.2000 438.4500 ;
	    RECT 37.8000 437.4000 39.0000 437.5500 ;
	    RECT 45.0000 437.4000 46.2000 437.5500 ;
	    RECT 66.6000 437.4000 67.8000 438.6000 ;
	    RECT 35.4000 434.4000 36.6000 435.6000 ;
	    RECT 35.4000 433.2000 36.6000 433.5000 ;
	    RECT 35.4000 423.3000 36.6000 429.3000 ;
	    RECT 37.8000 423.3000 39.0000 436.5000 ;
	    RECT 68.7000 435.3000 69.6000 440.4000 ;
	    RECT 93.0000 439.5000 94.2000 443.7000 ;
	    RECT 129.0000 441.6000 129.9000 443.7000 ;
	    RECT 131.7000 443.1000 137.1000 443.7000 ;
	    RECT 126.6000 440.4000 127.8000 441.6000 ;
	    RECT 129.0000 440.7000 130.5000 441.6000 ;
	    RECT 131.4000 440.4000 132.6000 441.6000 ;
	    RECT 135.0000 440.7000 135.3000 442.2000 ;
	    RECT 167.4000 441.6000 168.3000 443.7000 ;
	    RECT 170.1000 443.1000 175.5000 443.7000 ;
	    RECT 213.3000 443.1000 218.7000 443.7000 ;
	    RECT 136.2000 440.4000 137.4000 441.6000 ;
	    RECT 160.2000 441.4500 161.4000 441.6000 ;
	    RECT 165.0000 441.4500 166.2000 441.6000 ;
	    RECT 160.2000 440.5500 166.2000 441.4500 ;
	    RECT 167.4000 440.7000 168.9000 441.6000 ;
	    RECT 160.2000 440.4000 161.4000 440.5500 ;
	    RECT 165.0000 440.4000 166.2000 440.5500 ;
	    RECT 169.8000 440.4000 171.0000 441.6000 ;
	    RECT 173.4000 440.7000 173.7000 442.2000 ;
	    RECT 174.6000 440.4000 175.8000 441.6000 ;
	    RECT 198.6000 441.4500 199.8000 441.6000 ;
	    RECT 213.0000 441.4500 214.2000 441.6000 ;
	    RECT 198.6000 440.5500 214.2000 441.4500 ;
	    RECT 215.1000 440.7000 215.4000 442.2000 ;
	    RECT 220.5000 441.6000 221.4000 443.7000 ;
	    RECT 232.2000 443.5500 235.8000 444.4500 ;
	    RECT 232.2000 443.4000 233.4000 443.5500 ;
	    RECT 234.6000 443.4000 235.8000 443.5500 ;
	    RECT 237.0000 442.5000 238.2000 449.7000 ;
	    RECT 268.2000 448.8000 274.2000 449.7000 ;
	    RECT 268.2000 443.7000 269.4000 448.8000 ;
	    RECT 270.6000 443.7000 271.8000 447.9000 ;
	    RECT 273.0000 444.0000 274.2000 448.8000 ;
	    RECT 275.4000 444.9000 276.6000 449.7000 ;
	    RECT 277.8000 444.0000 279.0000 449.7000 ;
	    RECT 273.0000 443.7000 279.0000 444.0000 ;
	    RECT 270.6000 441.6000 271.5000 443.7000 ;
	    RECT 273.3000 443.1000 278.7000 443.7000 ;
	    RECT 289.8000 442.5000 291.0000 449.7000 ;
	    RECT 292.2000 446.7000 293.4000 449.7000 ;
	    RECT 292.2000 445.5000 293.4000 445.8000 ;
	    RECT 292.2000 444.4500 293.4000 444.6000 ;
	    RECT 313.8000 444.4500 315.0000 444.6000 ;
	    RECT 292.2000 443.5500 315.0000 444.4500 ;
	    RECT 316.2000 443.7000 317.4000 449.7000 ;
	    RECT 318.6000 444.0000 319.8000 449.7000 ;
	    RECT 321.0000 444.9000 322.2000 449.7000 ;
	    RECT 323.4000 444.0000 324.6000 449.7000 ;
	    RECT 318.6000 443.7000 324.6000 444.0000 ;
	    RECT 292.2000 443.4000 293.4000 443.5500 ;
	    RECT 313.8000 443.4000 315.0000 443.5500 ;
	    RECT 316.5000 442.5000 317.4000 443.7000 ;
	    RECT 318.9000 443.1000 324.3000 443.7000 ;
	    RECT 335.4000 442.5000 336.6000 449.7000 ;
	    RECT 337.8000 446.7000 339.0000 449.7000 ;
	    RECT 352.2000 446.7000 353.4000 449.7000 ;
	    RECT 337.8000 445.5000 339.0000 445.8000 ;
	    RECT 352.2000 445.5000 353.4000 445.8000 ;
	    RECT 337.8000 444.4500 339.0000 444.6000 ;
	    RECT 349.8000 444.4500 351.0000 444.6000 ;
	    RECT 337.8000 443.5500 351.0000 444.4500 ;
	    RECT 337.8000 443.4000 339.0000 443.5500 ;
	    RECT 349.8000 443.4000 351.0000 443.5500 ;
	    RECT 352.2000 443.4000 353.4000 444.6000 ;
	    RECT 354.6000 442.5000 355.8000 449.7000 ;
	    RECT 378.6000 444.0000 379.8000 449.7000 ;
	    RECT 381.0000 444.9000 382.2000 449.7000 ;
	    RECT 383.4000 444.0000 384.6000 449.7000 ;
	    RECT 378.6000 443.7000 384.6000 444.0000 ;
	    RECT 385.8000 443.7000 387.0000 449.7000 ;
	    RECT 405.9000 444.6000 407.1000 449.7000 ;
	    RECT 405.9000 443.7000 408.6000 444.6000 ;
	    RECT 409.8000 443.7000 411.0000 449.7000 ;
	    RECT 424.2000 446.7000 425.4000 449.7000 ;
	    RECT 424.2000 445.5000 425.4000 445.8000 ;
	    RECT 424.2000 444.4500 425.4000 444.6000 ;
	    RECT 378.9000 443.1000 384.3000 443.7000 ;
	    RECT 385.8000 442.5000 386.7000 443.7000 ;
	    RECT 198.6000 440.4000 199.8000 440.5500 ;
	    RECT 213.0000 440.4000 214.2000 440.5500 ;
	    RECT 217.8000 440.4000 219.0000 441.6000 ;
	    RECT 219.9000 440.7000 221.4000 441.6000 ;
	    RECT 222.6000 441.4500 223.8000 441.6000 ;
	    RECT 225.0000 441.4500 226.2000 441.6000 ;
	    RECT 222.6000 440.5500 226.2000 441.4500 ;
	    RECT 222.6000 440.4000 223.8000 440.5500 ;
	    RECT 225.0000 440.4000 226.2000 440.5500 ;
	    RECT 237.0000 441.4500 238.2000 441.6000 ;
	    RECT 263.4000 441.4500 264.6000 441.6000 ;
	    RECT 237.0000 440.5500 264.6000 441.4500 ;
	    RECT 237.0000 440.4000 238.2000 440.5500 ;
	    RECT 263.4000 440.4000 264.6000 440.5500 ;
	    RECT 268.2000 440.4000 269.4000 441.6000 ;
	    RECT 270.6000 440.7000 272.1000 441.6000 ;
	    RECT 273.0000 440.4000 274.2000 441.6000 ;
	    RECT 276.6000 440.7000 276.9000 442.2000 ;
	    RECT 277.8000 441.4500 279.0000 441.6000 ;
	    RECT 289.8000 441.4500 291.0000 441.6000 ;
	    RECT 277.8000 440.5500 291.0000 441.4500 ;
	    RECT 277.8000 440.4000 279.0000 440.5500 ;
	    RECT 289.8000 440.4000 291.0000 440.5500 ;
	    RECT 309.0000 441.4500 310.2000 441.6000 ;
	    RECT 316.2000 441.4500 317.4000 441.6000 ;
	    RECT 309.0000 440.5500 317.4000 441.4500 ;
	    RECT 309.0000 440.4000 310.2000 440.5500 ;
	    RECT 316.2000 440.4000 317.4000 440.5500 ;
	    RECT 318.3000 440.4000 320.1000 441.6000 ;
	    RECT 322.2000 440.7000 322.5000 442.2000 ;
	    RECT 323.4000 441.4500 324.6000 441.6000 ;
	    RECT 328.2000 441.4500 329.4000 441.6000 ;
	    RECT 323.4000 440.5500 329.4000 441.4500 ;
	    RECT 323.4000 440.4000 324.6000 440.5500 ;
	    RECT 328.2000 440.4000 329.4000 440.5500 ;
	    RECT 335.4000 441.4500 336.6000 441.6000 ;
	    RECT 345.0000 441.4500 346.2000 441.6000 ;
	    RECT 335.4000 440.5500 346.2000 441.4500 ;
	    RECT 335.4000 440.4000 336.6000 440.5500 ;
	    RECT 345.0000 440.4000 346.2000 440.5500 ;
	    RECT 354.6000 441.4500 355.8000 441.6000 ;
	    RECT 354.6000 440.5500 377.2500 441.4500 ;
	    RECT 354.6000 440.4000 355.8000 440.5500 ;
	    RECT 129.0000 439.5000 130.2000 439.8000 ;
	    RECT 133.8000 439.5000 135.0000 439.8000 ;
	    RECT 167.4000 439.5000 168.6000 439.8000 ;
	    RECT 172.2000 439.5000 173.4000 439.8000 ;
	    RECT 215.4000 439.5000 216.6000 439.8000 ;
	    RECT 220.2000 439.5000 221.4000 439.8000 ;
	    RECT 270.6000 439.5000 271.8000 439.8000 ;
	    RECT 275.4000 439.5000 276.6000 439.8000 ;
	    RECT 126.6000 439.2000 127.8000 439.5000 ;
	    RECT 93.0000 438.4500 94.2000 438.6000 ;
	    RECT 71.5500 437.5500 94.2000 438.4500 ;
	    RECT 71.5500 435.6000 72.4500 437.5500 ;
	    RECT 93.0000 437.4000 94.2000 437.5500 ;
	    RECT 129.0000 437.4000 130.2000 438.6000 ;
	    RECT 40.2000 423.3000 41.4000 429.3000 ;
	    RECT 64.2000 423.3000 65.4000 435.3000 ;
	    RECT 68.1000 434.4000 69.6000 435.3000 ;
	    RECT 71.4000 434.4000 72.6000 435.6000 ;
	    RECT 68.1000 423.3000 69.3000 434.4000 ;
	    RECT 70.5000 432.6000 71.4000 433.5000 ;
	    RECT 70.2000 431.4000 71.4000 432.6000 ;
	    RECT 70.5000 423.3000 71.7000 429.3000 ;
	    RECT 90.6000 423.3000 91.8000 429.3000 ;
	    RECT 93.0000 423.3000 94.2000 436.5000 ;
	    RECT 95.4000 435.4500 96.6000 435.6000 ;
	    RECT 124.2000 435.4500 125.4000 435.6000 ;
	    RECT 95.4000 434.5500 125.4000 435.4500 ;
	    RECT 131.7000 435.3000 132.6000 439.5000 ;
	    RECT 165.0000 439.2000 166.2000 439.5000 ;
	    RECT 133.8000 438.4500 135.0000 438.6000 ;
	    RECT 162.6000 438.4500 163.8000 438.6000 ;
	    RECT 133.8000 437.5500 163.8000 438.4500 ;
	    RECT 133.8000 437.4000 135.0000 437.5500 ;
	    RECT 162.6000 437.4000 163.8000 437.5500 ;
	    RECT 167.4000 437.4000 168.6000 438.6000 ;
	    RECT 170.1000 435.3000 171.0000 439.5000 ;
	    RECT 172.2000 438.4500 173.4000 438.6000 ;
	    RECT 186.6000 438.4500 187.8000 438.6000 ;
	    RECT 172.2000 437.5500 187.8000 438.4500 ;
	    RECT 172.2000 437.4000 173.4000 437.5500 ;
	    RECT 186.6000 437.4000 187.8000 437.5500 ;
	    RECT 193.8000 438.4500 195.0000 438.6000 ;
	    RECT 215.4000 438.4500 216.6000 438.6000 ;
	    RECT 193.8000 437.5500 216.6000 438.4500 ;
	    RECT 193.8000 437.4000 195.0000 437.5500 ;
	    RECT 215.4000 437.4000 216.6000 437.5500 ;
	    RECT 217.8000 435.3000 218.7000 439.5000 ;
	    RECT 222.6000 439.2000 223.8000 439.5000 ;
	    RECT 220.2000 437.4000 221.4000 438.6000 ;
	    RECT 95.4000 434.4000 96.6000 434.5500 ;
	    RECT 124.2000 434.4000 125.4000 434.5500 ;
	    RECT 95.4000 433.2000 96.6000 433.5000 ;
	    RECT 95.4000 423.3000 96.6000 429.3000 ;
	    RECT 126.6000 423.3000 127.8000 435.3000 ;
	    RECT 130.5000 423.3000 133.5000 435.3000 ;
	    RECT 136.2000 423.3000 137.4000 435.3000 ;
	    RECT 165.0000 423.3000 166.2000 435.3000 ;
	    RECT 168.9000 423.3000 171.9000 435.3000 ;
	    RECT 174.6000 423.3000 175.8000 435.3000 ;
	    RECT 213.0000 423.3000 214.2000 435.3000 ;
	    RECT 216.9000 423.3000 219.9000 435.3000 ;
	    RECT 222.6000 423.3000 223.8000 435.3000 ;
	    RECT 234.6000 423.3000 235.8000 429.3000 ;
	    RECT 237.0000 423.3000 238.2000 439.5000 ;
	    RECT 268.2000 439.2000 269.4000 439.5000 ;
	    RECT 270.6000 437.4000 271.8000 438.6000 ;
	    RECT 273.3000 435.3000 274.2000 439.5000 ;
	    RECT 275.4000 437.4000 276.6000 438.6000 ;
	    RECT 268.2000 423.3000 269.4000 435.3000 ;
	    RECT 272.1000 423.3000 275.1000 435.3000 ;
	    RECT 277.8000 423.3000 279.0000 435.3000 ;
	    RECT 289.8000 423.3000 291.0000 439.5000 ;
	    RECT 316.2000 434.4000 317.4000 435.6000 ;
	    RECT 319.2000 435.3000 320.1000 440.4000 ;
	    RECT 321.0000 439.5000 322.2000 439.8000 ;
	    RECT 321.0000 438.4500 322.2000 438.6000 ;
	    RECT 328.2000 438.4500 329.4000 438.6000 ;
	    RECT 321.0000 437.5500 329.4000 438.4500 ;
	    RECT 321.0000 437.4000 322.2000 437.5500 ;
	    RECT 328.2000 437.4000 329.4000 437.5500 ;
	    RECT 319.2000 434.4000 320.7000 435.3000 ;
	    RECT 317.4000 432.6000 318.3000 433.5000 ;
	    RECT 317.4000 431.4000 318.6000 432.6000 ;
	    RECT 292.2000 423.3000 293.4000 429.3000 ;
	    RECT 317.1000 423.3000 318.3000 429.3000 ;
	    RECT 319.5000 423.3000 320.7000 434.4000 ;
	    RECT 323.4000 423.3000 324.6000 435.3000 ;
	    RECT 335.4000 423.3000 336.6000 439.5000 ;
	    RECT 337.8000 423.3000 339.0000 429.3000 ;
	    RECT 352.2000 423.3000 353.4000 429.3000 ;
	    RECT 354.6000 423.3000 355.8000 439.5000 ;
	    RECT 376.3500 438.4500 377.2500 440.5500 ;
	    RECT 378.6000 440.4000 379.8000 441.6000 ;
	    RECT 380.7000 440.7000 381.0000 442.2000 ;
	    RECT 383.1000 440.4000 384.9000 441.6000 ;
	    RECT 385.8000 441.4500 387.0000 441.6000 ;
	    RECT 402.6000 441.4500 403.8000 441.6000 ;
	    RECT 385.8000 440.5500 403.8000 441.4500 ;
	    RECT 385.8000 440.4000 387.0000 440.5500 ;
	    RECT 402.6000 440.4000 403.8000 440.5500 ;
	    RECT 381.0000 439.5000 382.2000 439.8000 ;
	    RECT 381.0000 438.4500 382.2000 438.6000 ;
	    RECT 376.3500 437.5500 382.2000 438.4500 ;
	    RECT 381.0000 437.4000 382.2000 437.5500 ;
	    RECT 383.1000 435.3000 384.0000 440.4000 ;
	    RECT 407.4000 439.5000 408.6000 443.7000 ;
	    RECT 412.3500 443.5500 425.4000 444.4500 ;
	    RECT 409.8000 442.5000 411.0000 442.8000 ;
	    RECT 409.8000 441.4500 411.0000 441.6000 ;
	    RECT 412.3500 441.4500 413.2500 443.5500 ;
	    RECT 424.2000 443.4000 425.4000 443.5500 ;
	    RECT 426.6000 442.5000 427.8000 449.7000 ;
	    RECT 448.2000 442.5000 449.4000 449.7000 ;
	    RECT 450.6000 446.7000 451.8000 449.7000 ;
	    RECT 450.6000 445.5000 451.8000 445.8000 ;
	    RECT 450.6000 444.4500 451.8000 444.6000 ;
	    RECT 453.0000 444.4500 454.2000 444.6000 ;
	    RECT 450.6000 443.5500 454.2000 444.4500 ;
	    RECT 450.6000 443.4000 451.8000 443.5500 ;
	    RECT 453.0000 443.4000 454.2000 443.5500 ;
	    RECT 469.8000 442.8000 471.0000 449.7000 ;
	    RECT 472.2000 443.7000 473.4000 449.7000 ;
	    RECT 469.8000 441.9000 473.1000 442.8000 ;
	    RECT 474.6000 442.5000 475.8000 449.7000 ;
	    RECT 489.0000 442.5000 490.2000 449.7000 ;
	    RECT 491.4000 446.7000 492.6000 449.7000 ;
	    RECT 491.4000 445.5000 492.6000 445.8000 ;
	    RECT 491.4000 443.4000 492.6000 444.6000 ;
	    RECT 409.8000 440.5500 413.2500 441.4500 ;
	    RECT 426.6000 441.4500 427.8000 441.6000 ;
	    RECT 429.0000 441.4500 430.2000 441.6000 ;
	    RECT 426.6000 440.5500 430.2000 441.4500 ;
	    RECT 409.8000 440.4000 411.0000 440.5500 ;
	    RECT 426.6000 440.4000 427.8000 440.5500 ;
	    RECT 429.0000 440.4000 430.2000 440.5500 ;
	    RECT 448.2000 441.4500 449.4000 441.6000 ;
	    RECT 462.6000 441.4500 463.8000 441.6000 ;
	    RECT 448.2000 440.5500 463.8000 441.4500 ;
	    RECT 448.2000 440.4000 449.4000 440.5500 ;
	    RECT 462.6000 440.4000 463.8000 440.5500 ;
	    RECT 469.8000 439.5000 471.0000 439.8000 ;
	    RECT 407.4000 438.4500 408.6000 438.6000 ;
	    RECT 385.9500 437.5500 408.6000 438.4500 ;
	    RECT 385.9500 435.6000 386.8500 437.5500 ;
	    RECT 407.4000 437.4000 408.6000 437.5500 ;
	    RECT 378.6000 423.3000 379.8000 435.3000 ;
	    RECT 382.5000 434.4000 384.0000 435.3000 ;
	    RECT 385.8000 434.4000 387.0000 435.6000 ;
	    RECT 405.0000 434.4000 406.2000 435.6000 ;
	    RECT 382.5000 423.3000 383.7000 434.4000 ;
	    RECT 384.9000 432.6000 385.8000 433.5000 ;
	    RECT 405.0000 433.2000 406.2000 433.5000 ;
	    RECT 384.6000 431.4000 385.8000 432.6000 ;
	    RECT 384.9000 423.3000 386.1000 429.3000 ;
	    RECT 405.0000 423.3000 406.2000 429.3000 ;
	    RECT 407.4000 423.3000 408.6000 436.5000 ;
	    RECT 409.8000 423.3000 411.0000 429.3000 ;
	    RECT 424.2000 423.3000 425.4000 429.3000 ;
	    RECT 426.6000 423.3000 427.8000 439.5000 ;
	    RECT 448.2000 423.3000 449.4000 439.5000 ;
	    RECT 472.2000 437.4000 473.1000 441.9000 ;
	    RECT 474.6000 441.4500 475.8000 441.6000 ;
	    RECT 486.6000 441.4500 487.8000 441.6000 ;
	    RECT 474.6000 440.5500 487.8000 441.4500 ;
	    RECT 474.6000 440.4000 475.8000 440.5500 ;
	    RECT 486.6000 440.4000 487.8000 440.5500 ;
	    RECT 489.0000 441.4500 490.2000 441.6000 ;
	    RECT 522.6000 441.4500 523.8000 441.6000 ;
	    RECT 489.0000 440.5500 523.8000 441.4500 ;
	    RECT 489.0000 440.4000 490.2000 440.5500 ;
	    RECT 522.6000 440.4000 523.8000 440.5500 ;
	    RECT 618.6000 440.7000 619.8000 449.7000 ;
	    RECT 623.4000 443.7000 624.6000 449.7000 ;
	    RECT 628.2000 444.9000 629.4000 449.7000 ;
	    RECT 630.6000 445.5000 631.8000 449.7000 ;
	    RECT 633.0000 445.5000 634.2000 449.7000 ;
	    RECT 635.4000 445.5000 636.6000 449.7000 ;
	    RECT 637.8000 446.7000 639.0000 449.7000 ;
	    RECT 640.2000 445.5000 641.4000 449.7000 ;
	    RECT 642.6000 446.7000 643.8000 449.7000 ;
	    RECT 645.0000 445.5000 646.2000 449.7000 ;
	    RECT 647.4000 445.5000 648.6000 449.7000 ;
	    RECT 649.8000 445.5000 651.0000 449.7000 ;
	    RECT 652.2000 445.5000 653.4000 449.7000 ;
	    RECT 625.5000 443.7000 629.4000 444.9000 ;
	    RECT 654.6000 444.9000 655.8000 449.7000 ;
	    RECT 634.5000 443.7000 641.4000 444.6000 ;
	    RECT 625.5000 442.8000 626.7000 443.7000 ;
	    RECT 622.2000 441.6000 626.7000 442.8000 ;
	    RECT 618.6000 439.5000 631.8000 440.7000 ;
	    RECT 634.5000 440.1000 635.7000 443.7000 ;
	    RECT 640.2000 443.4000 641.4000 443.7000 ;
	    RECT 642.6000 443.4000 643.8000 444.6000 ;
	    RECT 644.7000 443.4000 645.0000 444.6000 ;
	    RECT 649.5000 443.4000 651.0000 444.6000 ;
	    RECT 654.6000 443.7000 658.2000 444.9000 ;
	    RECT 659.4000 443.7000 660.6000 449.7000 ;
	    RECT 637.8000 442.5000 639.0000 442.8000 ;
	    RECT 640.2000 442.2000 641.4000 442.5000 ;
	    RECT 637.8000 440.4000 639.0000 441.6000 ;
	    RECT 640.2000 441.3000 646.8000 442.2000 ;
	    RECT 645.6000 441.0000 646.8000 441.3000 ;
	    RECT 474.6000 438.6000 475.8000 439.5000 ;
	    RECT 472.2000 436.2000 474.0000 437.4000 ;
	    RECT 472.2000 435.3000 473.1000 436.2000 ;
	    RECT 474.9000 435.3000 475.8000 438.6000 ;
	    RECT 469.8000 434.4000 473.1000 435.3000 ;
	    RECT 450.6000 423.3000 451.8000 429.3000 ;
	    RECT 469.8000 423.3000 471.0000 434.4000 ;
	    RECT 472.2000 423.3000 473.4000 433.5000 ;
	    RECT 474.6000 423.3000 475.8000 435.3000 ;
	    RECT 489.0000 423.3000 490.2000 439.5000 ;
	    RECT 618.6000 431.1000 619.8000 439.5000 ;
	    RECT 632.7000 438.9000 635.7000 440.1000 ;
	    RECT 641.4000 438.9000 646.2000 440.1000 ;
	    RECT 649.8000 439.2000 651.0000 443.4000 ;
	    RECT 657.0000 442.8000 658.2000 443.7000 ;
	    RECT 657.0000 441.9000 659.7000 442.8000 ;
	    RECT 658.5000 440.1000 659.7000 441.9000 ;
	    RECT 664.2000 441.9000 665.4000 449.7000 ;
	    RECT 666.6000 444.0000 667.8000 449.7000 ;
	    RECT 669.0000 446.7000 670.2000 449.7000 ;
	    RECT 719.4000 449.4000 720.6000 450.6000 ;
	    RECT 666.6000 442.8000 668.1000 444.0000 ;
	    RECT 664.2000 441.0000 666.0000 441.9000 ;
	    RECT 658.5000 438.9000 664.2000 440.1000 ;
	    RECT 620.7000 438.0000 621.9000 438.3000 ;
	    RECT 620.7000 437.1000 627.3000 438.0000 ;
	    RECT 628.2000 437.4000 629.4000 438.6000 ;
	    RECT 654.6000 438.0000 655.8000 438.9000 ;
	    RECT 665.1000 438.0000 666.0000 441.0000 ;
	    RECT 630.3000 437.1000 655.8000 438.0000 ;
	    RECT 664.8000 437.1000 666.0000 438.0000 ;
	    RECT 662.7000 436.2000 663.9000 436.5000 ;
	    RECT 623.4000 434.4000 624.6000 435.6000 ;
	    RECT 625.5000 435.3000 663.9000 436.2000 ;
	    RECT 628.5000 435.0000 629.7000 435.3000 ;
	    RECT 664.8000 434.4000 665.7000 437.1000 ;
	    RECT 666.9000 436.2000 668.1000 442.8000 ;
	    RECT 745.8000 443.1000 747.0000 449.7000 ;
	    RECT 748.2000 444.0000 749.4000 449.7000 ;
	    RECT 752.1000 447.6000 753.9000 449.7000 ;
	    RECT 752.1000 446.7000 754.2000 447.6000 ;
	    RECT 756.6000 446.7000 757.8000 449.7000 ;
	    RECT 759.0000 446.7000 760.2000 449.7000 ;
	    RECT 761.4000 446.7000 762.9000 449.7000 ;
	    RECT 765.6000 447.6000 766.8000 449.7000 ;
	    RECT 765.6000 446.7000 768.6000 447.6000 ;
	    RECT 753.0000 445.5000 754.2000 446.7000 ;
	    RECT 759.3000 445.8000 760.2000 446.7000 ;
	    RECT 759.3000 444.9000 763.5000 445.8000 ;
	    RECT 762.3000 444.6000 763.5000 444.9000 ;
	    RECT 765.0000 444.6000 766.2000 445.8000 ;
	    RECT 767.4000 445.5000 768.6000 446.7000 ;
	    RECT 750.3000 443.1000 751.5000 443.4000 ;
	    RECT 745.8000 442.2000 751.5000 443.1000 ;
	    RECT 745.8000 439.5000 747.0000 442.2000 ;
	    RECT 756.3000 441.3000 757.5000 441.6000 ;
	    RECT 765.0000 441.3000 765.9000 444.6000 ;
	    RECT 769.8000 443.7000 771.0000 449.7000 ;
	    RECT 772.2000 442.5000 773.4000 449.7000 ;
	    RECT 786.6000 446.7000 787.8000 449.7000 ;
	    RECT 786.6000 445.5000 787.8000 445.8000 ;
	    RECT 786.6000 443.4000 787.8000 444.6000 ;
	    RECT 789.0000 442.5000 790.2000 449.7000 ;
	    RECT 801.0000 446.7000 802.2000 449.7000 ;
	    RECT 801.0000 445.5000 802.2000 445.8000 ;
	    RECT 796.2000 444.4500 797.4000 444.6000 ;
	    RECT 801.0000 444.4500 802.2000 444.6000 ;
	    RECT 796.2000 443.5500 802.2000 444.4500 ;
	    RECT 796.2000 443.4000 797.4000 443.5500 ;
	    RECT 801.0000 443.4000 802.2000 443.5500 ;
	    RECT 803.4000 442.5000 804.6000 449.7000 ;
	    RECT 815.4000 449.4000 816.6000 450.6000 ;
	    RECT 863.4000 449.4000 864.6000 450.6000 ;
	    RECT 873.0000 442.5000 874.2000 449.7000 ;
	    RECT 875.4000 443.7000 876.6000 449.7000 ;
	    RECT 879.6000 447.6000 880.8000 449.7000 ;
	    RECT 877.8000 446.7000 880.8000 447.6000 ;
	    RECT 883.5000 446.7000 885.0000 449.7000 ;
	    RECT 886.2000 446.7000 887.4000 449.7000 ;
	    RECT 888.6000 446.7000 889.8000 449.7000 ;
	    RECT 892.5000 447.6000 894.3000 449.7000 ;
	    RECT 892.2000 446.7000 894.3000 447.6000 ;
	    RECT 877.8000 445.5000 879.0000 446.7000 ;
	    RECT 886.2000 445.8000 887.1000 446.7000 ;
	    RECT 880.2000 444.6000 881.4000 445.8000 ;
	    RECT 882.9000 444.9000 887.1000 445.8000 ;
	    RECT 892.2000 445.5000 893.4000 446.7000 ;
	    RECT 882.9000 444.6000 884.1000 444.9000 ;
	    RECT 755.7000 440.4000 768.9000 441.3000 ;
	    RECT 769.8000 440.4000 771.0000 441.6000 ;
	    RECT 771.9000 440.4000 772.2000 441.6000 ;
	    RECT 784.2000 441.4500 785.4000 441.6000 ;
	    RECT 789.0000 441.4500 790.2000 441.6000 ;
	    RECT 784.2000 440.5500 790.2000 441.4500 ;
	    RECT 784.2000 440.4000 785.4000 440.5500 ;
	    RECT 789.0000 440.4000 790.2000 440.5500 ;
	    RECT 803.4000 441.4500 804.6000 441.6000 ;
	    RECT 870.6000 441.4500 871.8000 441.6000 ;
	    RECT 803.4000 440.5500 871.8000 441.4500 ;
	    RECT 803.4000 440.4000 804.6000 440.5500 ;
	    RECT 870.6000 440.4000 871.8000 440.5500 ;
	    RECT 874.2000 440.4000 874.5000 441.6000 ;
	    RECT 875.4000 440.4000 876.6000 441.6000 ;
	    RECT 880.5000 441.3000 881.4000 444.6000 ;
	    RECT 897.0000 444.0000 898.2000 449.7000 ;
	    RECT 894.9000 443.1000 896.1000 443.4000 ;
	    RECT 899.4000 443.1000 900.6000 449.7000 ;
	    RECT 918.6000 446.7000 919.8000 449.7000 ;
	    RECT 918.6000 445.5000 919.8000 445.8000 ;
	    RECT 904.2000 444.4500 905.4000 444.6000 ;
	    RECT 918.6000 444.4500 919.8000 444.6000 ;
	    RECT 904.2000 443.5500 919.8000 444.4500 ;
	    RECT 904.2000 443.4000 905.4000 443.5500 ;
	    RECT 918.6000 443.4000 919.8000 443.5500 ;
	    RECT 894.9000 442.2000 900.6000 443.1000 ;
	    RECT 921.0000 442.5000 922.2000 449.7000 ;
	    RECT 993.0000 444.4500 994.2000 444.6000 ;
	    RECT 1033.8000 444.4500 1035.0000 444.6000 ;
	    RECT 993.0000 443.5500 1035.0000 444.4500 ;
	    RECT 993.0000 443.4000 994.2000 443.5500 ;
	    RECT 1033.8000 443.4000 1035.0000 443.5500 ;
	    RECT 888.9000 441.3000 890.1000 441.6000 ;
	    RECT 877.5000 440.4000 890.7000 441.3000 ;
	    RECT 753.0000 439.2000 754.2000 439.5000 ;
	    RECT 745.8000 437.4000 747.0000 438.6000 ;
	    RECT 748.5000 438.3000 754.2000 439.2000 ;
	    RECT 748.5000 438.0000 749.7000 438.3000 ;
	    RECT 750.9000 437.1000 752.1000 437.4000 ;
	    RECT 747.9000 436.5000 752.1000 437.1000 ;
	    RECT 633.0000 434.1000 634.2000 434.4000 ;
	    RECT 626.1000 433.5000 634.2000 434.1000 ;
	    RECT 624.9000 433.2000 634.2000 433.5000 ;
	    RECT 635.7000 433.5000 648.6000 434.4000 ;
	    RECT 621.0000 432.0000 623.4000 433.2000 ;
	    RECT 624.9000 432.3000 627.0000 433.2000 ;
	    RECT 635.7000 432.3000 636.6000 433.5000 ;
	    RECT 647.4000 433.2000 648.6000 433.5000 ;
	    RECT 652.2000 433.5000 665.7000 434.4000 ;
	    RECT 666.6000 435.0000 668.1000 436.2000 ;
	    RECT 745.8000 436.2000 752.1000 436.5000 ;
	    RECT 666.6000 433.5000 667.8000 435.0000 ;
	    RECT 652.2000 433.2000 653.4000 433.5000 ;
	    RECT 622.5000 431.4000 623.4000 432.0000 ;
	    RECT 627.9000 431.4000 636.6000 432.3000 ;
	    RECT 637.5000 431.4000 641.4000 432.6000 ;
	    RECT 618.6000 430.2000 621.6000 431.1000 ;
	    RECT 622.5000 430.2000 628.8000 431.4000 ;
	    RECT 620.7000 429.3000 621.6000 430.2000 ;
	    RECT 491.4000 423.3000 492.6000 429.3000 ;
	    RECT 618.6000 423.3000 619.8000 429.3000 ;
	    RECT 620.7000 428.4000 622.2000 429.3000 ;
	    RECT 621.0000 423.3000 622.2000 428.4000 ;
	    RECT 623.4000 422.4000 624.6000 429.3000 ;
	    RECT 625.8000 423.3000 627.0000 430.2000 ;
	    RECT 628.2000 423.3000 629.4000 429.3000 ;
	    RECT 630.6000 423.3000 631.8000 427.5000 ;
	    RECT 633.0000 423.3000 634.2000 427.5000 ;
	    RECT 635.4000 423.3000 636.6000 430.5000 ;
	    RECT 637.8000 423.3000 639.0000 429.3000 ;
	    RECT 640.2000 423.3000 641.4000 430.5000 ;
	    RECT 642.6000 423.3000 643.8000 429.3000 ;
	    RECT 645.0000 423.3000 646.2000 432.6000 ;
	    RECT 657.0000 431.4000 660.9000 432.6000 ;
	    RECT 649.8000 430.2000 656.1000 431.4000 ;
	    RECT 647.4000 423.3000 648.6000 427.5000 ;
	    RECT 649.8000 423.3000 651.0000 427.5000 ;
	    RECT 652.2000 423.3000 653.4000 427.5000 ;
	    RECT 654.6000 423.3000 655.8000 429.3000 ;
	    RECT 657.0000 423.3000 658.2000 431.4000 ;
	    RECT 664.8000 431.1000 665.7000 433.5000 ;
	    RECT 666.6000 431.4000 667.8000 432.6000 ;
	    RECT 661.8000 430.2000 665.7000 431.1000 ;
	    RECT 659.4000 423.3000 660.6000 429.3000 ;
	    RECT 661.8000 423.3000 663.0000 430.2000 ;
	    RECT 664.2000 423.3000 665.4000 429.3000 ;
	    RECT 666.6000 423.3000 667.8000 430.5000 ;
	    RECT 669.0000 423.3000 670.2000 429.3000 ;
	    RECT 693.0000 426.4500 694.2000 426.6000 ;
	    RECT 719.4000 426.4500 720.6000 426.6000 ;
	    RECT 693.0000 425.5500 720.6000 426.4500 ;
	    RECT 693.0000 425.4000 694.2000 425.5500 ;
	    RECT 719.4000 425.4000 720.6000 425.5500 ;
	    RECT 745.8000 423.3000 747.0000 436.2000 ;
	    RECT 755.7000 435.6000 756.6000 440.4000 ;
	    RECT 766.5000 440.1000 767.7000 440.4000 ;
	    RECT 878.7000 440.1000 879.9000 440.4000 ;
	    RECT 768.9000 438.6000 770.1000 438.9000 ;
	    RECT 762.6000 437.4000 763.8000 438.6000 ;
	    RECT 764.7000 437.7000 770.1000 438.6000 ;
	    RECT 765.0000 436.5000 773.4000 436.8000 ;
	    RECT 764.7000 436.2000 773.4000 436.5000 ;
	    RECT 748.2000 423.3000 749.4000 435.3000 ;
	    RECT 753.0000 434.7000 756.6000 435.6000 ;
	    RECT 758.7000 435.9000 773.4000 436.2000 ;
	    RECT 758.7000 435.3000 765.9000 435.9000 ;
	    RECT 753.0000 433.2000 753.9000 434.7000 ;
	    RECT 751.8000 432.0000 753.9000 433.2000 ;
	    RECT 756.3000 433.5000 757.5000 433.8000 ;
	    RECT 758.7000 433.5000 759.6000 435.3000 ;
	    RECT 756.3000 432.6000 759.6000 433.5000 ;
	    RECT 760.5000 433.5000 768.6000 434.4000 ;
	    RECT 760.5000 433.2000 761.7000 433.5000 ;
	    RECT 767.4000 433.2000 768.6000 433.5000 ;
	    RECT 758.1000 431.1000 759.3000 431.4000 ;
	    RECT 762.3000 431.1000 763.5000 431.4000 ;
	    RECT 753.0000 429.3000 754.2000 430.5000 ;
	    RECT 758.1000 430.2000 763.5000 431.1000 ;
	    RECT 759.3000 429.3000 760.2000 430.2000 ;
	    RECT 767.4000 429.3000 768.6000 430.5000 ;
	    RECT 752.1000 423.3000 753.9000 429.3000 ;
	    RECT 756.6000 423.3000 757.8000 429.3000 ;
	    RECT 759.0000 423.3000 760.2000 429.3000 ;
	    RECT 761.4000 423.3000 762.6000 429.3000 ;
	    RECT 765.6000 428.4000 768.6000 429.3000 ;
	    RECT 765.6000 423.3000 766.8000 428.4000 ;
	    RECT 769.8000 423.3000 771.0000 435.0000 ;
	    RECT 772.2000 423.3000 773.4000 435.9000 ;
	    RECT 786.6000 423.3000 787.8000 429.3000 ;
	    RECT 789.0000 423.3000 790.2000 439.5000 ;
	    RECT 801.0000 423.3000 802.2000 429.3000 ;
	    RECT 803.4000 423.3000 804.6000 439.5000 ;
	    RECT 876.3000 438.6000 877.5000 438.9000 ;
	    RECT 876.3000 437.7000 881.7000 438.6000 ;
	    RECT 882.6000 437.4000 883.8000 438.6000 ;
	    RECT 873.0000 436.5000 881.4000 436.8000 ;
	    RECT 873.0000 436.2000 881.7000 436.5000 ;
	    RECT 873.0000 435.9000 887.7000 436.2000 ;
	    RECT 873.0000 423.3000 874.2000 435.9000 ;
	    RECT 880.5000 435.3000 887.7000 435.9000 ;
	    RECT 875.4000 423.3000 876.6000 435.0000 ;
	    RECT 877.8000 433.5000 885.9000 434.4000 ;
	    RECT 877.8000 433.2000 879.0000 433.5000 ;
	    RECT 884.7000 433.2000 885.9000 433.5000 ;
	    RECT 886.8000 433.5000 887.7000 435.3000 ;
	    RECT 889.8000 435.6000 890.7000 440.4000 ;
	    RECT 899.4000 439.5000 900.6000 442.2000 ;
	    RECT 921.0000 441.4500 922.2000 441.6000 ;
	    RECT 957.0000 441.4500 958.2000 441.6000 ;
	    RECT 921.0000 440.5500 958.2000 441.4500 ;
	    RECT 921.0000 440.4000 922.2000 440.5500 ;
	    RECT 957.0000 440.4000 958.2000 440.5500 ;
	    RECT 971.4000 441.4500 972.6000 441.6000 ;
	    RECT 1005.0000 441.4500 1006.2000 441.6000 ;
	    RECT 971.4000 440.5500 1006.2000 441.4500 ;
	    RECT 971.4000 440.4000 972.6000 440.5500 ;
	    RECT 1005.0000 440.4000 1006.2000 440.5500 ;
	    RECT 1045.8000 440.7000 1047.0000 449.7000 ;
	    RECT 1050.6000 443.7000 1051.8000 449.7000 ;
	    RECT 1055.4000 444.9000 1056.6000 449.7000 ;
	    RECT 1057.8000 445.5000 1059.0000 449.7000 ;
	    RECT 1060.2001 445.5000 1061.4000 449.7000 ;
	    RECT 1062.6000 445.5000 1063.8000 449.7000 ;
	    RECT 1065.0000 446.7000 1066.2001 449.7000 ;
	    RECT 1067.4000 445.5000 1068.6000 449.7000 ;
	    RECT 1069.8000 446.7000 1071.0000 449.7000 ;
	    RECT 1072.2001 445.5000 1073.4000 449.7000 ;
	    RECT 1074.6000 445.5000 1075.8000 449.7000 ;
	    RECT 1077.0000 445.5000 1078.2001 449.7000 ;
	    RECT 1079.4000 445.5000 1080.6000 449.7000 ;
	    RECT 1052.7001 443.7000 1056.6000 444.9000 ;
	    RECT 1081.8000 444.9000 1083.0000 449.7000 ;
	    RECT 1061.7001 443.7000 1068.6000 444.6000 ;
	    RECT 1052.7001 442.8000 1053.9000 443.7000 ;
	    RECT 1049.4000 441.6000 1053.9000 442.8000 ;
	    RECT 1045.8000 439.5000 1059.0000 440.7000 ;
	    RECT 1061.7001 440.1000 1062.9000 443.7000 ;
	    RECT 1067.4000 443.4000 1068.6000 443.7000 ;
	    RECT 1069.8000 443.4000 1071.0000 444.6000 ;
	    RECT 1071.9000 443.4000 1072.2001 444.6000 ;
	    RECT 1076.7001 443.4000 1078.2001 444.6000 ;
	    RECT 1081.8000 443.7000 1085.4000 444.9000 ;
	    RECT 1086.6000 443.7000 1087.8000 449.7000 ;
	    RECT 1065.0000 442.5000 1066.2001 442.8000 ;
	    RECT 1067.4000 442.2000 1068.6000 442.5000 ;
	    RECT 1065.0000 440.4000 1066.2001 441.6000 ;
	    RECT 1067.4000 441.3000 1074.0000 442.2000 ;
	    RECT 1072.8000 441.0000 1074.0000 441.3000 ;
	    RECT 892.2000 439.2000 893.4000 439.5000 ;
	    RECT 892.2000 438.3000 897.9000 439.2000 ;
	    RECT 896.7000 438.0000 897.9000 438.3000 ;
	    RECT 899.4000 437.4000 900.6000 438.6000 ;
	    RECT 894.3000 437.1000 895.5000 437.4000 ;
	    RECT 894.3000 436.5000 898.5000 437.1000 ;
	    RECT 894.3000 436.2000 900.6000 436.5000 ;
	    RECT 889.8000 434.7000 893.4000 435.6000 ;
	    RECT 888.9000 433.5000 890.1000 433.8000 ;
	    RECT 886.8000 432.6000 890.1000 433.5000 ;
	    RECT 892.5000 433.2000 893.4000 434.7000 ;
	    RECT 892.5000 432.0000 894.6000 433.2000 ;
	    RECT 882.9000 431.1000 884.1000 431.4000 ;
	    RECT 887.1000 431.1000 888.3000 431.4000 ;
	    RECT 877.8000 429.3000 879.0000 430.5000 ;
	    RECT 882.9000 430.2000 888.3000 431.1000 ;
	    RECT 886.2000 429.3000 887.1000 430.2000 ;
	    RECT 892.2000 429.3000 893.4000 430.5000 ;
	    RECT 877.8000 428.4000 880.8000 429.3000 ;
	    RECT 879.6000 423.3000 880.8000 428.4000 ;
	    RECT 883.8000 423.3000 885.0000 429.3000 ;
	    RECT 886.2000 423.3000 887.4000 429.3000 ;
	    RECT 888.6000 423.3000 889.8000 429.3000 ;
	    RECT 892.5000 423.3000 894.3000 429.3000 ;
	    RECT 897.0000 423.3000 898.2000 435.3000 ;
	    RECT 899.4000 423.3000 900.6000 436.2000 ;
	    RECT 918.6000 423.3000 919.8000 429.3000 ;
	    RECT 921.0000 423.3000 922.2000 439.5000 ;
	    RECT 1045.8000 431.1000 1047.0000 439.5000 ;
	    RECT 1059.9000 438.9000 1062.9000 440.1000 ;
	    RECT 1068.6000 438.9000 1073.4000 440.1000 ;
	    RECT 1077.0000 439.2000 1078.2001 443.4000 ;
	    RECT 1084.2001 442.8000 1085.4000 443.7000 ;
	    RECT 1084.2001 441.9000 1086.9000 442.8000 ;
	    RECT 1085.7001 440.1000 1086.9000 441.9000 ;
	    RECT 1091.4000 441.9000 1092.6000 449.7000 ;
	    RECT 1093.8000 444.0000 1095.0000 449.7000 ;
	    RECT 1096.2001 446.7000 1097.4000 449.7000 ;
	    RECT 1116.3000 444.6000 1117.5000 449.7000 ;
	    RECT 1093.8000 442.8000 1095.3000 444.0000 ;
	    RECT 1116.3000 443.7000 1119.0000 444.6000 ;
	    RECT 1120.2001 443.7000 1121.4000 449.7000 ;
	    RECT 1141.8000 446.7000 1143.0000 449.7000 ;
	    RECT 1141.8000 445.5000 1143.0000 445.8000 ;
	    RECT 1122.6000 444.4500 1123.8000 444.6000 ;
	    RECT 1141.8000 444.4500 1143.0000 444.6000 ;
	    RECT 1091.4000 441.0000 1093.2001 441.9000 ;
	    RECT 1085.7001 438.9000 1091.4000 440.1000 ;
	    RECT 1047.9000 438.0000 1049.1000 438.3000 ;
	    RECT 1047.9000 437.1000 1054.5000 438.0000 ;
	    RECT 1055.4000 437.4000 1056.6000 438.6000 ;
	    RECT 1081.8000 438.0000 1083.0000 438.9000 ;
	    RECT 1092.3000 438.0000 1093.2001 441.0000 ;
	    RECT 1057.5000 437.1000 1083.0000 438.0000 ;
	    RECT 1092.0000 437.1000 1093.2001 438.0000 ;
	    RECT 1089.9000 436.2000 1091.1000 436.5000 ;
	    RECT 1050.6000 434.4000 1051.8000 435.6000 ;
	    RECT 1052.7001 435.3000 1091.1000 436.2000 ;
	    RECT 1055.7001 435.0000 1056.9000 435.3000 ;
	    RECT 1092.0000 434.4000 1092.9000 437.1000 ;
	    RECT 1094.1000 436.2000 1095.3000 442.8000 ;
	    RECT 1117.8000 439.5000 1119.0000 443.7000 ;
	    RECT 1122.6000 443.5500 1143.0000 444.4500 ;
	    RECT 1122.6000 443.4000 1123.8000 443.5500 ;
	    RECT 1141.8000 443.4000 1143.0000 443.5500 ;
	    RECT 1120.2001 442.5000 1121.4000 442.8000 ;
	    RECT 1144.2001 442.5000 1145.4000 449.7000 ;
	    RECT 1164.3000 444.6000 1165.5000 449.7000 ;
	    RECT 1164.3000 443.7000 1167.0000 444.6000 ;
	    RECT 1168.2001 443.7000 1169.4000 449.7000 ;
	    RECT 1192.2001 444.0000 1193.4000 449.7000 ;
	    RECT 1194.6000 444.9000 1195.8000 449.7000 ;
	    RECT 1197.0000 444.0000 1198.2001 449.7000 ;
	    RECT 1192.2001 443.7000 1198.2001 444.0000 ;
	    RECT 1199.4000 443.7000 1200.6000 449.7000 ;
	    RECT 1213.8000 446.7000 1215.0000 449.7000 ;
	    RECT 1213.8000 445.5000 1215.0000 445.8000 ;
	    RECT 1201.8000 444.4500 1203.0000 444.6000 ;
	    RECT 1213.8000 444.4500 1215.0000 444.6000 ;
	    RECT 1120.2001 440.4000 1121.4000 441.6000 ;
	    RECT 1144.2001 441.4500 1145.4000 441.6000 ;
	    RECT 1163.4000 441.4500 1164.6000 441.6000 ;
	    RECT 1144.2001 440.5500 1164.6000 441.4500 ;
	    RECT 1144.2001 440.4000 1145.4000 440.5500 ;
	    RECT 1163.4000 440.4000 1164.6000 440.5500 ;
	    RECT 1165.8000 439.5000 1167.0000 443.7000 ;
	    RECT 1192.5000 443.1000 1197.9000 443.7000 ;
	    RECT 1168.2001 442.5000 1169.4000 442.8000 ;
	    RECT 1199.4000 442.5000 1200.3000 443.7000 ;
	    RECT 1201.8000 443.5500 1215.0000 444.4500 ;
	    RECT 1201.8000 443.4000 1203.0000 443.5500 ;
	    RECT 1213.8000 443.4000 1215.0000 443.5500 ;
	    RECT 1216.2001 442.5000 1217.4000 449.7000 ;
	    RECT 1168.2001 441.4500 1169.4000 441.6000 ;
	    RECT 1175.4000 441.4500 1176.6000 441.6000 ;
	    RECT 1168.2001 440.5500 1176.6000 441.4500 ;
	    RECT 1168.2001 440.4000 1169.4000 440.5500 ;
	    RECT 1175.4000 440.4000 1176.6000 440.5500 ;
	    RECT 1192.2001 440.4000 1193.4000 441.6000 ;
	    RECT 1194.3000 440.7000 1194.6000 442.2000 ;
	    RECT 1196.7001 440.4000 1198.5000 441.6000 ;
	    RECT 1199.4000 441.4500 1200.6000 441.6000 ;
	    RECT 1213.8000 441.4500 1215.0000 441.6000 ;
	    RECT 1199.4000 440.5500 1215.0000 441.4500 ;
	    RECT 1199.4000 440.4000 1200.6000 440.5500 ;
	    RECT 1213.8000 440.4000 1215.0000 440.5500 ;
	    RECT 1216.2001 441.4500 1217.4000 441.6000 ;
	    RECT 1221.0000 441.4500 1222.2001 441.6000 ;
	    RECT 1216.2001 440.5500 1222.2001 441.4500 ;
	    RECT 1242.6000 440.7000 1243.8000 449.7000 ;
	    RECT 1248.0000 441.3000 1249.2001 449.7000 ;
	    RECT 1248.0000 440.7000 1250.7001 441.3000 ;
	    RECT 1273.8000 440.7000 1275.0000 449.7000 ;
	    RECT 1279.2001 441.3000 1280.4000 449.7000 ;
	    RECT 1300.2001 443.7000 1301.4000 449.7000 ;
	    RECT 1304.1000 444.6000 1305.3000 449.7000 ;
	    RECT 1302.6000 443.7000 1305.3000 444.6000 ;
	    RECT 1329.0000 443.7000 1330.2001 449.7000 ;
	    RECT 1331.4000 444.0000 1332.6000 449.7000 ;
	    RECT 1333.8000 444.9000 1335.0000 449.7000 ;
	    RECT 1336.2001 444.0000 1337.4000 449.7000 ;
	    RECT 1331.4000 443.7000 1337.4000 444.0000 ;
	    RECT 1369.8000 444.0000 1371.0000 449.7000 ;
	    RECT 1372.2001 444.9000 1373.4000 449.7000 ;
	    RECT 1374.6000 444.0000 1375.8000 449.7000 ;
	    RECT 1369.8000 443.7000 1375.8000 444.0000 ;
	    RECT 1377.0000 443.7000 1378.2001 449.7000 ;
	    RECT 1403.4000 444.0000 1404.6000 449.7000 ;
	    RECT 1405.8000 444.9000 1407.0000 449.7000 ;
	    RECT 1408.2001 444.0000 1409.4000 449.7000 ;
	    RECT 1403.4000 443.7000 1409.4000 444.0000 ;
	    RECT 1410.6000 443.7000 1411.8000 449.7000 ;
	    RECT 1300.2001 442.5000 1301.4000 442.8000 ;
	    RECT 1295.4000 441.4500 1296.6000 441.6000 ;
	    RECT 1300.2001 441.4500 1301.4000 441.6000 ;
	    RECT 1279.2001 440.7000 1281.9000 441.3000 ;
	    RECT 1216.2001 440.4000 1217.4000 440.5500 ;
	    RECT 1221.0000 440.4000 1222.2001 440.5500 ;
	    RECT 1248.3000 440.4000 1250.7001 440.7000 ;
	    RECT 1279.5000 440.4000 1281.9000 440.7000 ;
	    RECT 1295.4000 440.5500 1301.4000 441.4500 ;
	    RECT 1295.4000 440.4000 1296.6000 440.5500 ;
	    RECT 1300.2001 440.4000 1301.4000 440.5500 ;
	    RECT 1194.6000 439.5000 1195.8000 439.8000 ;
	    RECT 1117.8000 438.4500 1119.0000 438.6000 ;
	    RECT 1141.8000 438.4500 1143.0000 438.6000 ;
	    RECT 1117.8000 437.5500 1143.0000 438.4500 ;
	    RECT 1117.8000 437.4000 1119.0000 437.5500 ;
	    RECT 1141.8000 437.4000 1143.0000 437.5500 ;
	    RECT 1060.2001 434.1000 1061.4000 434.4000 ;
	    RECT 1053.3000 433.5000 1061.4000 434.1000 ;
	    RECT 1052.1000 433.2000 1061.4000 433.5000 ;
	    RECT 1062.9000 433.5000 1075.8000 434.4000 ;
	    RECT 1048.2001 432.0000 1050.6000 433.2000 ;
	    RECT 1052.1000 432.3000 1054.2001 433.2000 ;
	    RECT 1062.9000 432.3000 1063.8000 433.5000 ;
	    RECT 1074.6000 433.2000 1075.8000 433.5000 ;
	    RECT 1079.4000 433.5000 1092.9000 434.4000 ;
	    RECT 1093.8000 435.0000 1095.3000 436.2000 ;
	    RECT 1093.8000 433.5000 1095.0000 435.0000 ;
	    RECT 1115.4000 434.4000 1116.6000 435.6000 ;
	    RECT 1079.4000 433.2000 1080.6000 433.5000 ;
	    RECT 1049.7001 431.4000 1050.6000 432.0000 ;
	    RECT 1055.1000 431.4000 1063.8000 432.3000 ;
	    RECT 1064.7001 431.4000 1068.6000 432.6000 ;
	    RECT 1045.8000 430.2000 1048.8000 431.1000 ;
	    RECT 1049.7001 430.2000 1056.0000 431.4000 ;
	    RECT 1047.9000 429.3000 1048.8000 430.2000 ;
	    RECT 947.4000 426.4500 948.6000 426.6000 ;
	    RECT 971.4000 426.4500 972.6000 426.6000 ;
	    RECT 978.6000 426.4500 979.8000 426.6000 ;
	    RECT 947.4000 425.5500 979.8000 426.4500 ;
	    RECT 947.4000 425.4000 948.6000 425.5500 ;
	    RECT 971.4000 425.4000 972.6000 425.5500 ;
	    RECT 978.6000 425.4000 979.8000 425.5500 ;
	    RECT 1045.8000 423.3000 1047.0000 429.3000 ;
	    RECT 1047.9000 428.4000 1049.4000 429.3000 ;
	    RECT 1048.2001 423.3000 1049.4000 428.4000 ;
	    RECT 1050.6000 422.4000 1051.8000 429.3000 ;
	    RECT 1053.0000 423.3000 1054.2001 430.2000 ;
	    RECT 1055.4000 423.3000 1056.6000 429.3000 ;
	    RECT 1057.8000 423.3000 1059.0000 427.5000 ;
	    RECT 1060.2001 423.3000 1061.4000 427.5000 ;
	    RECT 1062.6000 423.3000 1063.8000 430.5000 ;
	    RECT 1065.0000 423.3000 1066.2001 429.3000 ;
	    RECT 1067.4000 423.3000 1068.6000 430.5000 ;
	    RECT 1069.8000 423.3000 1071.0000 429.3000 ;
	    RECT 1072.2001 423.3000 1073.4000 432.6000 ;
	    RECT 1084.2001 431.4000 1088.1000 432.6000 ;
	    RECT 1077.0000 430.2000 1083.3000 431.4000 ;
	    RECT 1074.6000 423.3000 1075.8000 427.5000 ;
	    RECT 1077.0000 423.3000 1078.2001 427.5000 ;
	    RECT 1079.4000 423.3000 1080.6000 427.5000 ;
	    RECT 1081.8000 423.3000 1083.0000 429.3000 ;
	    RECT 1084.2001 423.3000 1085.4000 431.4000 ;
	    RECT 1092.0000 431.1000 1092.9000 433.5000 ;
	    RECT 1115.4000 433.2000 1116.6000 433.5000 ;
	    RECT 1093.8000 431.4000 1095.0000 432.6000 ;
	    RECT 1089.0000 430.2000 1092.9000 431.1000 ;
	    RECT 1086.6000 423.3000 1087.8000 429.3000 ;
	    RECT 1089.0000 423.3000 1090.2001 430.2000 ;
	    RECT 1091.4000 423.3000 1092.6000 429.3000 ;
	    RECT 1093.8000 423.3000 1095.0000 430.5000 ;
	    RECT 1096.2001 423.3000 1097.4000 429.3000 ;
	    RECT 1115.4000 423.3000 1116.6000 429.3000 ;
	    RECT 1117.8000 423.3000 1119.0000 436.5000 ;
	    RECT 1120.2001 423.3000 1121.4000 429.3000 ;
	    RECT 1141.8000 423.3000 1143.0000 429.3000 ;
	    RECT 1144.2001 423.3000 1145.4000 439.5000 ;
	    RECT 1165.8000 437.4000 1167.0000 438.6000 ;
	    RECT 1194.6000 437.4000 1195.8000 438.6000 ;
	    RECT 1146.6000 435.4500 1147.8000 435.6000 ;
	    RECT 1163.4000 435.4500 1164.6000 435.6000 ;
	    RECT 1146.6000 434.5500 1164.6000 435.4500 ;
	    RECT 1146.6000 434.4000 1147.8000 434.5500 ;
	    RECT 1163.4000 434.4000 1164.6000 434.5500 ;
	    RECT 1163.4000 433.2000 1164.6000 433.5000 ;
	    RECT 1163.4000 423.3000 1164.6000 429.3000 ;
	    RECT 1165.8000 423.3000 1167.0000 436.5000 ;
	    RECT 1196.7001 435.3000 1197.6000 440.4000 ;
	    RECT 1168.2001 423.3000 1169.4000 429.3000 ;
	    RECT 1192.2001 423.3000 1193.4000 435.3000 ;
	    RECT 1196.1000 434.4000 1197.6000 435.3000 ;
	    RECT 1199.4000 435.4500 1200.6000 435.6000 ;
	    RECT 1211.4000 435.4500 1212.6000 435.6000 ;
	    RECT 1199.4000 434.5500 1212.6000 435.4500 ;
	    RECT 1199.4000 434.4000 1200.6000 434.5500 ;
	    RECT 1211.4000 434.4000 1212.6000 434.5500 ;
	    RECT 1196.1000 423.3000 1197.3000 434.4000 ;
	    RECT 1198.5000 432.6000 1199.4000 433.5000 ;
	    RECT 1198.2001 431.4000 1199.4000 432.6000 ;
	    RECT 1198.5000 423.3000 1199.7001 429.3000 ;
	    RECT 1213.8000 423.3000 1215.0000 429.3000 ;
	    RECT 1216.2001 423.3000 1217.4000 439.5000 ;
	    RECT 1245.0000 437.4000 1246.2001 438.6000 ;
	    RECT 1247.1000 437.4000 1247.4000 438.6000 ;
	    RECT 1242.6000 436.5000 1243.8000 436.8000 ;
	    RECT 1249.8000 436.5000 1250.7001 440.4000 ;
	    RECT 1276.2001 437.4000 1277.4000 438.6000 ;
	    RECT 1278.3000 437.4000 1278.6000 438.6000 ;
	    RECT 1273.8000 436.5000 1275.0000 436.8000 ;
	    RECT 1281.0000 436.5000 1281.9000 440.4000 ;
	    RECT 1302.6000 439.5000 1303.8000 443.7000 ;
	    RECT 1329.3000 442.5000 1330.2001 443.7000 ;
	    RECT 1331.7001 443.1000 1337.1000 443.7000 ;
	    RECT 1370.1000 443.1000 1375.5000 443.7000 ;
	    RECT 1377.0000 442.5000 1377.9000 443.7000 ;
	    RECT 1403.7001 443.1000 1409.1000 443.7000 ;
	    RECT 1410.6000 442.5000 1411.5000 443.7000 ;
	    RECT 1329.0000 440.4000 1330.2001 441.6000 ;
	    RECT 1331.1000 440.4000 1332.9000 441.6000 ;
	    RECT 1335.0000 440.7000 1335.3000 442.2000 ;
	    RECT 1336.2001 440.4000 1337.4000 441.6000 ;
	    RECT 1345.8000 441.4500 1347.0000 441.6000 ;
	    RECT 1369.8000 441.4500 1371.0000 441.6000 ;
	    RECT 1345.8000 440.5500 1371.0000 441.4500 ;
	    RECT 1371.9000 440.7000 1372.2001 442.2000 ;
	    RECT 1345.8000 440.4000 1347.0000 440.5500 ;
	    RECT 1369.8000 440.4000 1371.0000 440.5500 ;
	    RECT 1374.3000 440.4000 1376.1000 441.6000 ;
	    RECT 1377.0000 440.4000 1378.2001 441.6000 ;
	    RECT 1384.2001 441.4500 1385.4000 441.6000 ;
	    RECT 1403.4000 441.4500 1404.6000 441.6000 ;
	    RECT 1384.2001 440.5500 1404.6000 441.4500 ;
	    RECT 1405.5000 440.7000 1405.8000 442.2000 ;
	    RECT 1384.2001 440.4000 1385.4000 440.5500 ;
	    RECT 1403.4000 440.4000 1404.6000 440.5500 ;
	    RECT 1407.9000 440.4000 1409.7001 441.6000 ;
	    RECT 1410.6000 441.4500 1411.8000 441.6000 ;
	    RECT 1420.2001 441.4500 1421.4000 441.6000 ;
	    RECT 1410.6000 440.5500 1421.4000 441.4500 ;
	    RECT 1434.6000 440.7000 1435.8000 449.7000 ;
	    RECT 1440.0000 441.3000 1441.2001 449.7000 ;
	    RECT 1461.0000 443.7000 1462.2001 449.7000 ;
	    RECT 1464.9000 444.6000 1466.1000 449.7000 ;
	    RECT 1468.2001 447.4500 1469.4000 447.6000 ;
	    RECT 1482.6000 447.4500 1483.8000 447.6000 ;
	    RECT 1468.2001 446.5500 1483.8000 447.4500 ;
	    RECT 1468.2001 446.4000 1469.4000 446.5500 ;
	    RECT 1482.6000 446.4000 1483.8000 446.5500 ;
	    RECT 1463.4000 443.7000 1466.1000 444.6000 ;
	    RECT 1461.0000 442.5000 1462.2001 442.8000 ;
	    RECT 1440.0000 440.7000 1442.7001 441.3000 ;
	    RECT 1410.6000 440.4000 1411.8000 440.5500 ;
	    RECT 1420.2001 440.4000 1421.4000 440.5500 ;
	    RECT 1440.3000 440.4000 1442.7001 440.7000 ;
	    RECT 1461.0000 440.4000 1462.2001 441.6000 ;
	    RECT 1302.6000 438.4500 1303.8000 438.6000 ;
	    RECT 1329.0000 438.4500 1330.2001 438.6000 ;
	    RECT 1302.6000 437.5500 1330.2001 438.4500 ;
	    RECT 1302.6000 437.4000 1303.8000 437.5500 ;
	    RECT 1329.0000 437.4000 1330.2001 437.5500 ;
	    RECT 1237.8000 435.4500 1239.0000 435.6000 ;
	    RECT 1242.6000 435.4500 1243.8000 435.6000 ;
	    RECT 1237.8000 434.5500 1243.8000 435.4500 ;
	    RECT 1237.8000 434.4000 1239.0000 434.5500 ;
	    RECT 1242.6000 434.4000 1243.8000 434.5500 ;
	    RECT 1249.8000 435.4500 1251.0000 435.6000 ;
	    RECT 1254.6000 435.4500 1255.8000 435.6000 ;
	    RECT 1249.8000 434.5500 1255.8000 435.4500 ;
	    RECT 1249.8000 434.4000 1251.0000 434.5500 ;
	    RECT 1254.6000 434.4000 1255.8000 434.5500 ;
	    RECT 1261.8000 435.4500 1263.0000 435.6000 ;
	    RECT 1273.8000 435.4500 1275.0000 435.6000 ;
	    RECT 1261.8000 434.5500 1275.0000 435.4500 ;
	    RECT 1261.8000 434.4000 1263.0000 434.5500 ;
	    RECT 1273.8000 434.4000 1275.0000 434.5500 ;
	    RECT 1281.0000 434.4000 1282.2001 435.6000 ;
	    RECT 1247.4000 433.5000 1248.6000 433.8000 ;
	    RECT 1278.6000 433.5000 1279.8000 433.8000 ;
	    RECT 1247.4000 431.4000 1248.6000 432.6000 ;
	    RECT 1249.8000 430.5000 1250.7001 433.5000 ;
	    RECT 1273.8000 432.4500 1275.0000 432.6000 ;
	    RECT 1278.6000 432.4500 1279.8000 432.6000 ;
	    RECT 1273.8000 431.5500 1279.8000 432.4500 ;
	    RECT 1273.8000 431.4000 1275.0000 431.5500 ;
	    RECT 1278.6000 431.4000 1279.8000 431.5500 ;
	    RECT 1281.0000 430.5000 1281.9000 433.5000 ;
	    RECT 1245.3000 429.6000 1250.7001 430.5000 ;
	    RECT 1245.3000 429.3000 1246.2001 429.6000 ;
	    RECT 1242.6000 423.3000 1243.8000 429.3000 ;
	    RECT 1245.0000 423.3000 1246.2001 429.3000 ;
	    RECT 1249.8000 429.3000 1250.7001 429.6000 ;
	    RECT 1276.5000 429.6000 1281.9000 430.5000 ;
	    RECT 1276.5000 429.3000 1277.4000 429.6000 ;
	    RECT 1247.4000 423.3000 1248.6000 428.7000 ;
	    RECT 1249.8000 423.3000 1251.0000 429.3000 ;
	    RECT 1273.8000 423.3000 1275.0000 429.3000 ;
	    RECT 1276.2001 423.3000 1277.4000 429.3000 ;
	    RECT 1281.0000 429.3000 1281.9000 429.6000 ;
	    RECT 1278.6000 423.3000 1279.8000 428.7000 ;
	    RECT 1281.0000 423.3000 1282.2001 429.3000 ;
	    RECT 1300.2001 423.3000 1301.4000 429.3000 ;
	    RECT 1302.6000 423.3000 1303.8000 436.5000 ;
	    RECT 1305.0000 434.4000 1306.2001 435.6000 ;
	    RECT 1321.8000 435.4500 1323.0000 435.6000 ;
	    RECT 1329.0000 435.4500 1330.2001 435.6000 ;
	    RECT 1321.8000 434.5500 1330.2001 435.4500 ;
	    RECT 1321.8000 434.4000 1323.0000 434.5500 ;
	    RECT 1329.0000 434.4000 1330.2001 434.5500 ;
	    RECT 1332.0000 435.3000 1332.9000 440.4000 ;
	    RECT 1333.8000 439.5000 1335.0000 439.8000 ;
	    RECT 1372.2001 439.5000 1373.4000 439.8000 ;
	    RECT 1333.8000 437.4000 1335.0000 438.6000 ;
	    RECT 1338.6000 438.4500 1339.8000 438.6000 ;
	    RECT 1372.2001 438.4500 1373.4000 438.6000 ;
	    RECT 1338.6000 437.5500 1373.4000 438.4500 ;
	    RECT 1338.6000 437.4000 1339.8000 437.5500 ;
	    RECT 1372.2001 437.4000 1373.4000 437.5500 ;
	    RECT 1374.3000 435.3000 1375.2001 440.4000 ;
	    RECT 1405.8000 439.5000 1407.0000 439.8000 ;
	    RECT 1405.8000 437.4000 1407.0000 438.6000 ;
	    RECT 1332.0000 434.4000 1333.5000 435.3000 ;
	    RECT 1305.0000 433.2000 1306.2001 433.5000 ;
	    RECT 1330.2001 432.6000 1331.1000 433.5000 ;
	    RECT 1330.2001 431.4000 1331.4000 432.6000 ;
	    RECT 1305.0000 423.3000 1306.2001 429.3000 ;
	    RECT 1329.9000 423.3000 1331.1000 429.3000 ;
	    RECT 1332.3000 423.3000 1333.5000 434.4000 ;
	    RECT 1336.2001 423.3000 1337.4000 435.3000 ;
	    RECT 1369.8000 423.3000 1371.0000 435.3000 ;
	    RECT 1373.7001 434.4000 1375.2001 435.3000 ;
	    RECT 1377.0000 435.4500 1378.2001 435.6000 ;
	    RECT 1379.4000 435.4500 1380.6000 435.6000 ;
	    RECT 1377.0000 434.5500 1380.6000 435.4500 ;
	    RECT 1407.9000 435.3000 1408.8000 440.4000 ;
	    RECT 1437.0000 437.4000 1438.2001 438.6000 ;
	    RECT 1439.1000 437.4000 1439.4000 438.6000 ;
	    RECT 1434.6000 436.5000 1435.8000 436.8000 ;
	    RECT 1441.8000 436.5000 1442.7001 440.4000 ;
	    RECT 1463.4000 439.5000 1464.6000 443.7000 ;
	    RECT 1535.4000 442.5000 1536.6000 449.7000 ;
	    RECT 1537.8000 443.7000 1539.0000 449.7000 ;
	    RECT 1542.0000 447.6000 1543.2001 449.7000 ;
	    RECT 1540.2001 446.7000 1543.2001 447.6000 ;
	    RECT 1545.9000 446.7000 1547.4000 449.7000 ;
	    RECT 1548.6000 446.7000 1549.8000 449.7000 ;
	    RECT 1551.0000 446.7000 1552.2001 449.7000 ;
	    RECT 1554.9000 447.6000 1556.7001 449.7000 ;
	    RECT 1554.6000 446.7000 1556.7001 447.6000 ;
	    RECT 1540.2001 445.5000 1541.4000 446.7000 ;
	    RECT 1548.6000 445.8000 1549.5000 446.7000 ;
	    RECT 1542.6000 444.6000 1543.8000 445.8000 ;
	    RECT 1545.3000 444.9000 1549.5000 445.8000 ;
	    RECT 1554.6000 445.5000 1555.8000 446.7000 ;
	    RECT 1545.3000 444.6000 1546.5000 444.9000 ;
	    RECT 1536.6000 440.4000 1536.9000 441.6000 ;
	    RECT 1537.8000 440.4000 1539.0000 441.6000 ;
	    RECT 1542.9000 441.3000 1543.8000 444.6000 ;
	    RECT 1559.4000 444.0000 1560.6000 449.7000 ;
	    RECT 1557.3000 443.1000 1558.5000 443.4000 ;
	    RECT 1561.8000 443.1000 1563.0000 449.7000 ;
	    RECT 1557.3000 442.2000 1563.0000 443.1000 ;
	    RECT 1551.3000 441.3000 1552.5000 441.6000 ;
	    RECT 1539.9000 440.4000 1553.1000 441.3000 ;
	    RECT 1541.1000 440.1000 1542.3000 440.4000 ;
	    RECT 1538.7001 438.6000 1539.9000 438.9000 ;
	    RECT 1463.4000 438.4500 1464.6000 438.6000 ;
	    RECT 1470.6000 438.4500 1471.8000 438.6000 ;
	    RECT 1463.4000 437.5500 1471.8000 438.4500 ;
	    RECT 1538.7001 437.7000 1544.1000 438.6000 ;
	    RECT 1463.4000 437.4000 1464.6000 437.5500 ;
	    RECT 1470.6000 437.4000 1471.8000 437.5500 ;
	    RECT 1545.0000 437.4000 1546.2001 438.6000 ;
	    RECT 1535.4000 436.5000 1543.8000 436.8000 ;
	    RECT 1377.0000 434.4000 1378.2001 434.5500 ;
	    RECT 1379.4000 434.4000 1380.6000 434.5500 ;
	    RECT 1373.7001 423.3000 1374.9000 434.4000 ;
	    RECT 1376.1000 432.6000 1377.0000 433.5000 ;
	    RECT 1375.8000 431.4000 1377.0000 432.6000 ;
	    RECT 1376.1000 423.3000 1377.3000 429.3000 ;
	    RECT 1403.4000 423.3000 1404.6000 435.3000 ;
	    RECT 1407.3000 434.4000 1408.8000 435.3000 ;
	    RECT 1410.6000 434.4000 1411.8000 435.6000 ;
	    RECT 1415.4000 435.4500 1416.6000 435.6000 ;
	    RECT 1427.4000 435.4500 1428.6000 435.6000 ;
	    RECT 1434.6000 435.4500 1435.8000 435.6000 ;
	    RECT 1415.4000 434.5500 1435.8000 435.4500 ;
	    RECT 1415.4000 434.4000 1416.6000 434.5500 ;
	    RECT 1427.4000 434.4000 1428.6000 434.5500 ;
	    RECT 1434.6000 434.4000 1435.8000 434.5500 ;
	    RECT 1441.8000 435.4500 1443.0000 435.6000 ;
	    RECT 1444.2001 435.4500 1445.4000 435.6000 ;
	    RECT 1441.8000 434.5500 1445.4000 435.4500 ;
	    RECT 1441.8000 434.4000 1443.0000 434.5500 ;
	    RECT 1444.2001 434.4000 1445.4000 434.5500 ;
	    RECT 1407.3000 423.3000 1408.5000 434.4000 ;
	    RECT 1439.4000 433.5000 1440.6000 433.8000 ;
	    RECT 1409.7001 432.6000 1410.6000 433.5000 ;
	    RECT 1409.4000 431.4000 1410.6000 432.6000 ;
	    RECT 1420.2001 432.4500 1421.4000 432.6000 ;
	    RECT 1439.4000 432.4500 1440.6000 432.6000 ;
	    RECT 1420.2001 431.5500 1440.6000 432.4500 ;
	    RECT 1420.2001 431.4000 1421.4000 431.5500 ;
	    RECT 1439.4000 431.4000 1440.6000 431.5500 ;
	    RECT 1441.8000 430.5000 1442.7001 433.5000 ;
	    RECT 1437.3000 429.6000 1442.7001 430.5000 ;
	    RECT 1437.3000 429.3000 1438.2001 429.6000 ;
	    RECT 1409.7001 423.3000 1410.9000 429.3000 ;
	    RECT 1434.6000 423.3000 1435.8000 429.3000 ;
	    RECT 1437.0000 423.3000 1438.2001 429.3000 ;
	    RECT 1441.8000 429.3000 1442.7001 429.6000 ;
	    RECT 1439.4000 423.3000 1440.6000 428.7000 ;
	    RECT 1441.8000 423.3000 1443.0000 429.3000 ;
	    RECT 1461.0000 423.3000 1462.2001 429.3000 ;
	    RECT 1463.4000 423.3000 1464.6000 436.5000 ;
	    RECT 1535.4000 436.2000 1544.1000 436.5000 ;
	    RECT 1535.4000 435.9000 1550.1000 436.2000 ;
	    RECT 1465.8000 434.4000 1467.0000 435.6000 ;
	    RECT 1465.8000 433.2000 1467.0000 433.5000 ;
	    RECT 1465.8000 423.3000 1467.0000 429.3000 ;
	    RECT 1504.2001 426.4500 1505.4000 426.6000 ;
	    RECT 1523.4000 426.4500 1524.6000 426.6000 ;
	    RECT 1504.2001 425.5500 1524.6000 426.4500 ;
	    RECT 1504.2001 425.4000 1505.4000 425.5500 ;
	    RECT 1523.4000 425.4000 1524.6000 425.5500 ;
	    RECT 1535.4000 423.3000 1536.6000 435.9000 ;
	    RECT 1542.9000 435.3000 1550.1000 435.9000 ;
	    RECT 1537.8000 423.3000 1539.0000 435.0000 ;
	    RECT 1540.2001 433.5000 1548.3000 434.4000 ;
	    RECT 1540.2001 433.2000 1541.4000 433.5000 ;
	    RECT 1547.1000 433.2000 1548.3000 433.5000 ;
	    RECT 1549.2001 433.5000 1550.1000 435.3000 ;
	    RECT 1552.2001 435.6000 1553.1000 440.4000 ;
	    RECT 1561.8000 439.5000 1563.0000 442.2000 ;
	    RECT 1554.6000 439.2000 1555.8000 439.5000 ;
	    RECT 1554.6000 438.3000 1560.3000 439.2000 ;
	    RECT 1559.1000 438.0000 1560.3000 438.3000 ;
	    RECT 1561.8000 437.4000 1563.0000 438.6000 ;
	    RECT 1556.7001 437.1000 1557.9000 437.4000 ;
	    RECT 1556.7001 436.5000 1560.9000 437.1000 ;
	    RECT 1556.7001 436.2000 1563.0000 436.5000 ;
	    RECT 1552.2001 434.7000 1555.8000 435.6000 ;
	    RECT 1551.3000 433.5000 1552.5000 433.8000 ;
	    RECT 1549.2001 432.6000 1552.5000 433.5000 ;
	    RECT 1554.9000 433.2000 1555.8000 434.7000 ;
	    RECT 1554.9000 432.0000 1557.0000 433.2000 ;
	    RECT 1545.3000 431.1000 1546.5000 431.4000 ;
	    RECT 1549.5000 431.1000 1550.7001 431.4000 ;
	    RECT 1540.2001 429.3000 1541.4000 430.5000 ;
	    RECT 1545.3000 430.2000 1550.7001 431.1000 ;
	    RECT 1548.6000 429.3000 1549.5000 430.2000 ;
	    RECT 1554.6000 429.3000 1555.8000 430.5000 ;
	    RECT 1540.2001 428.4000 1543.2001 429.3000 ;
	    RECT 1542.0000 423.3000 1543.2001 428.4000 ;
	    RECT 1546.2001 423.3000 1547.4000 429.3000 ;
	    RECT 1548.6000 423.3000 1549.8000 429.3000 ;
	    RECT 1551.0000 423.3000 1552.2001 429.3000 ;
	    RECT 1554.9000 423.3000 1556.7001 429.3000 ;
	    RECT 1559.4000 423.3000 1560.6000 435.3000 ;
	    RECT 1561.8000 423.3000 1563.0000 436.2000 ;
	    RECT 1.2000 420.6000 1569.0000 422.4000 ;
	    RECT 13.8000 403.5000 15.0000 419.7000 ;
	    RECT 16.2000 413.7000 17.4000 419.7000 ;
	    RECT 35.4000 413.7000 36.6000 419.7000 ;
	    RECT 35.4000 409.5000 36.6000 409.8000 ;
	    RECT 35.4000 407.4000 36.6000 408.6000 ;
	    RECT 37.8000 406.5000 39.0000 419.7000 ;
	    RECT 40.2000 413.7000 41.4000 419.7000 ;
	    RECT 65.1000 413.7000 66.3000 419.7000 ;
	    RECT 65.4000 410.4000 66.6000 411.6000 ;
	    RECT 65.4000 409.5000 66.3000 410.4000 ;
	    RECT 67.5000 408.6000 68.7000 419.7000 ;
	    RECT 64.2000 407.4000 65.4000 408.6000 ;
	    RECT 67.2000 407.7000 68.7000 408.6000 ;
	    RECT 71.4000 407.7000 72.6000 419.7000 ;
	    RECT 37.8000 405.4500 39.0000 405.6000 ;
	    RECT 64.3500 405.4500 65.2500 407.4000 ;
	    RECT 37.8000 404.5500 65.2500 405.4500 ;
	    RECT 37.8000 404.4000 39.0000 404.5500 ;
	    RECT 13.8000 402.4500 15.0000 402.6000 ;
	    RECT 33.0000 402.4500 34.2000 402.6000 ;
	    RECT 13.8000 401.5500 34.2000 402.4500 ;
	    RECT 13.8000 401.4000 15.0000 401.5500 ;
	    RECT 33.0000 401.4000 34.2000 401.5500 ;
	    RECT 13.8000 393.3000 15.0000 400.5000 ;
	    RECT 16.2000 398.4000 17.4000 399.6000 ;
	    RECT 37.8000 399.3000 39.0000 403.5000 ;
	    RECT 67.2000 402.6000 68.1000 407.7000 ;
	    RECT 69.0000 405.4500 70.2000 405.6000 ;
	    RECT 69.0000 404.5500 74.8500 405.4500 ;
	    RECT 69.0000 404.4000 70.2000 404.5500 ;
	    RECT 69.0000 403.2000 70.2000 403.5000 ;
	    RECT 40.2000 402.4500 41.4000 402.6000 ;
	    RECT 42.6000 402.4500 43.8000 402.6000 ;
	    RECT 40.2000 401.5500 43.8000 402.4500 ;
	    RECT 40.2000 401.4000 41.4000 401.5500 ;
	    RECT 42.6000 401.4000 43.8000 401.5500 ;
	    RECT 64.2000 401.4000 65.4000 402.6000 ;
	    RECT 66.3000 401.4000 68.1000 402.6000 ;
	    RECT 70.2000 400.8000 70.5000 402.3000 ;
	    RECT 71.4000 401.4000 72.6000 402.6000 ;
	    RECT 73.9500 402.4500 74.8500 404.5500 ;
	    RECT 85.8000 403.5000 87.0000 419.7000 ;
	    RECT 88.2000 413.7000 89.4000 419.7000 ;
	    RECT 102.6000 413.7000 103.8000 419.7000 ;
	    RECT 105.0000 403.5000 106.2000 419.7000 ;
	    RECT 119.4000 413.7000 120.6000 419.7000 ;
	    RECT 121.8000 403.5000 123.0000 419.7000 ;
	    RECT 136.2000 413.7000 137.4000 419.7000 ;
	    RECT 138.6000 403.5000 139.8000 419.7000 ;
	    RECT 167.4000 417.4500 168.6000 417.6000 ;
	    RECT 270.6000 417.4500 271.8000 417.6000 ;
	    RECT 167.4000 416.5500 271.8000 417.4500 ;
	    RECT 167.4000 416.4000 168.6000 416.5500 ;
	    RECT 270.6000 416.4000 271.8000 416.5500 ;
	    RECT 273.0000 413.7000 274.2000 419.7000 ;
	    RECT 275.4000 412.5000 276.6000 419.7000 ;
	    RECT 277.8000 413.7000 279.0000 419.7000 ;
	    RECT 280.2000 412.8000 281.4000 419.7000 ;
	    RECT 282.6000 413.7000 283.8000 419.7000 ;
	    RECT 277.5000 411.9000 281.4000 412.8000 ;
	    RECT 220.2000 411.4500 221.4000 411.6000 ;
	    RECT 232.2000 411.4500 233.4000 411.6000 ;
	    RECT 275.4000 411.4500 276.6000 411.6000 ;
	    RECT 220.2000 410.5500 276.6000 411.4500 ;
	    RECT 220.2000 410.4000 221.4000 410.5500 ;
	    RECT 232.2000 410.4000 233.4000 410.5500 ;
	    RECT 275.4000 410.4000 276.6000 410.5500 ;
	    RECT 277.5000 409.5000 278.4000 411.9000 ;
	    RECT 285.0000 411.6000 286.2000 419.7000 ;
	    RECT 287.4000 413.7000 288.6000 419.7000 ;
	    RECT 289.8000 415.5000 291.0000 419.7000 ;
	    RECT 292.2000 415.5000 293.4000 419.7000 ;
	    RECT 294.6000 415.5000 295.8000 419.7000 ;
	    RECT 287.1000 411.6000 293.4000 412.8000 ;
	    RECT 282.3000 410.4000 286.2000 411.6000 ;
	    RECT 297.0000 410.4000 298.2000 419.7000 ;
	    RECT 299.4000 413.7000 300.6000 419.7000 ;
	    RECT 301.8000 412.5000 303.0000 419.7000 ;
	    RECT 304.2000 413.7000 305.4000 419.7000 ;
	    RECT 306.6000 412.5000 307.8000 419.7000 ;
	    RECT 309.0000 415.5000 310.2000 419.7000 ;
	    RECT 311.4000 415.5000 312.6000 419.7000 ;
	    RECT 313.8000 413.7000 315.0000 419.7000 ;
	    RECT 316.2000 412.8000 317.4000 419.7000 ;
	    RECT 318.6000 413.7000 319.8000 420.6000 ;
	    RECT 321.0000 414.6000 322.2000 419.7000 ;
	    RECT 321.0000 413.7000 322.5000 414.6000 ;
	    RECT 323.4000 413.7000 324.6000 419.7000 ;
	    RECT 321.6000 412.8000 322.5000 413.7000 ;
	    RECT 314.4000 411.6000 320.7000 412.8000 ;
	    RECT 321.6000 411.9000 324.6000 412.8000 ;
	    RECT 301.8000 410.4000 305.7000 411.6000 ;
	    RECT 306.6000 410.7000 315.3000 411.6000 ;
	    RECT 319.8000 411.0000 320.7000 411.6000 ;
	    RECT 289.8000 409.5000 291.0000 409.8000 ;
	    RECT 275.4000 408.0000 276.6000 409.5000 ;
	    RECT 275.1000 406.8000 276.6000 408.0000 ;
	    RECT 277.5000 408.6000 291.0000 409.5000 ;
	    RECT 294.6000 409.5000 295.8000 409.8000 ;
	    RECT 306.6000 409.5000 307.5000 410.7000 ;
	    RECT 316.2000 409.8000 318.3000 410.7000 ;
	    RECT 319.8000 409.8000 322.2000 411.0000 ;
	    RECT 294.6000 408.6000 307.5000 409.5000 ;
	    RECT 309.0000 409.5000 318.3000 409.8000 ;
	    RECT 309.0000 408.9000 317.1000 409.5000 ;
	    RECT 309.0000 408.6000 310.2000 408.9000 ;
	    RECT 85.8000 402.4500 87.0000 402.6000 ;
	    RECT 73.9500 401.5500 87.0000 402.4500 ;
	    RECT 85.8000 401.4000 87.0000 401.5500 ;
	    RECT 105.0000 402.4500 106.2000 402.6000 ;
	    RECT 119.4000 402.4500 120.6000 402.6000 ;
	    RECT 105.0000 401.5500 120.6000 402.4500 ;
	    RECT 105.0000 401.4000 106.2000 401.5500 ;
	    RECT 119.4000 401.4000 120.6000 401.5500 ;
	    RECT 121.8000 402.4500 123.0000 402.6000 ;
	    RECT 136.2000 402.4500 137.4000 402.6000 ;
	    RECT 121.8000 401.5500 137.4000 402.4500 ;
	    RECT 121.8000 401.4000 123.0000 401.5500 ;
	    RECT 136.2000 401.4000 137.4000 401.5500 ;
	    RECT 138.6000 402.4500 139.8000 402.6000 ;
	    RECT 198.6000 402.4500 199.8000 402.6000 ;
	    RECT 138.6000 401.5500 199.8000 402.4500 ;
	    RECT 138.6000 401.4000 139.8000 401.5500 ;
	    RECT 198.6000 401.4000 199.8000 401.5500 ;
	    RECT 40.2000 400.2000 41.4000 400.5000 ;
	    RECT 64.5000 399.3000 65.4000 400.5000 ;
	    RECT 66.9000 399.3000 72.3000 399.9000 ;
	    RECT 36.3000 398.4000 39.0000 399.3000 ;
	    RECT 16.2000 397.2000 17.4000 397.5000 ;
	    RECT 16.2000 393.3000 17.4000 396.3000 ;
	    RECT 36.3000 393.3000 37.5000 398.4000 ;
	    RECT 40.2000 393.3000 41.4000 399.3000 ;
	    RECT 64.2000 393.3000 65.4000 399.3000 ;
	    RECT 66.6000 399.0000 72.6000 399.3000 ;
	    RECT 66.6000 393.3000 67.8000 399.0000 ;
	    RECT 69.0000 393.3000 70.2000 398.1000 ;
	    RECT 71.4000 393.3000 72.6000 399.0000 ;
	    RECT 85.8000 393.3000 87.0000 400.5000 ;
	    RECT 88.2000 398.4000 89.4000 399.6000 ;
	    RECT 90.6000 399.4500 91.8000 399.6000 ;
	    RECT 102.6000 399.4500 103.8000 399.6000 ;
	    RECT 90.6000 398.5500 103.8000 399.4500 ;
	    RECT 90.6000 398.4000 91.8000 398.5500 ;
	    RECT 102.6000 398.4000 103.8000 398.5500 ;
	    RECT 88.2000 397.2000 89.4000 397.5000 ;
	    RECT 102.6000 397.2000 103.8000 397.5000 ;
	    RECT 88.2000 393.3000 89.4000 396.3000 ;
	    RECT 102.6000 393.3000 103.8000 396.3000 ;
	    RECT 105.0000 393.3000 106.2000 400.5000 ;
	    RECT 119.4000 398.4000 120.6000 399.6000 ;
	    RECT 119.4000 397.2000 120.6000 397.5000 ;
	    RECT 119.4000 393.3000 120.6000 396.3000 ;
	    RECT 121.8000 393.3000 123.0000 400.5000 ;
	    RECT 131.4000 399.4500 132.6000 399.6000 ;
	    RECT 136.2000 399.4500 137.4000 399.6000 ;
	    RECT 131.4000 398.5500 137.4000 399.4500 ;
	    RECT 131.4000 398.4000 132.6000 398.5500 ;
	    RECT 136.2000 398.4000 137.4000 398.5500 ;
	    RECT 136.2000 397.2000 137.4000 397.5000 ;
	    RECT 136.2000 393.3000 137.4000 396.3000 ;
	    RECT 138.6000 393.3000 139.8000 400.5000 ;
	    RECT 275.1000 400.2000 276.3000 406.8000 ;
	    RECT 277.5000 405.9000 278.4000 408.6000 ;
	    RECT 313.5000 407.7000 314.7000 408.0000 ;
	    RECT 279.3000 406.8000 317.7000 407.7000 ;
	    RECT 318.6000 407.4000 319.8000 408.6000 ;
	    RECT 279.3000 406.5000 280.5000 406.8000 ;
	    RECT 277.2000 405.0000 278.4000 405.9000 ;
	    RECT 287.4000 405.0000 312.9000 405.9000 ;
	    RECT 277.2000 402.0000 278.1000 405.0000 ;
	    RECT 287.4000 404.1000 288.6000 405.0000 ;
	    RECT 313.8000 404.4000 315.0000 405.6000 ;
	    RECT 315.9000 405.0000 322.5000 405.9000 ;
	    RECT 321.3000 404.7000 322.5000 405.0000 ;
	    RECT 279.0000 402.9000 284.7000 404.1000 ;
	    RECT 277.2000 401.1000 279.0000 402.0000 ;
	    RECT 275.1000 399.0000 276.6000 400.2000 ;
	    RECT 273.0000 393.3000 274.2000 396.3000 ;
	    RECT 275.4000 393.3000 276.6000 399.0000 ;
	    RECT 277.8000 393.3000 279.0000 401.1000 ;
	    RECT 283.5000 401.1000 284.7000 402.9000 ;
	    RECT 283.5000 400.2000 286.2000 401.1000 ;
	    RECT 285.0000 399.3000 286.2000 400.2000 ;
	    RECT 292.2000 399.6000 293.4000 403.8000 ;
	    RECT 297.0000 402.9000 301.8000 404.1000 ;
	    RECT 307.5000 402.9000 310.5000 404.1000 ;
	    RECT 323.4000 403.5000 324.6000 411.9000 ;
	    RECT 337.8000 403.5000 339.0000 419.7000 ;
	    RECT 340.2000 413.7000 341.4000 419.7000 ;
	    RECT 378.6000 419.4000 379.8000 420.6000 ;
	    RECT 405.0000 419.4000 406.2000 420.6000 ;
	    RECT 421.8000 417.4500 423.0000 417.6000 ;
	    RECT 424.3500 417.4500 425.2500 420.6000 ;
	    RECT 448.2000 419.4000 449.4000 420.6000 ;
	    RECT 421.8000 416.5500 425.2500 417.4500 ;
	    RECT 421.8000 416.4000 423.0000 416.5500 ;
	    RECT 472.2000 413.7000 473.4000 419.7000 ;
	    RECT 474.6000 412.5000 475.8000 419.7000 ;
	    RECT 477.0000 413.7000 478.2000 419.7000 ;
	    RECT 479.4000 412.8000 480.6000 419.7000 ;
	    RECT 481.8000 413.7000 483.0000 419.7000 ;
	    RECT 476.7000 411.9000 480.6000 412.8000 ;
	    RECT 424.2000 411.4500 425.4000 411.6000 ;
	    RECT 474.6000 411.4500 475.8000 411.6000 ;
	    RECT 424.2000 410.5500 475.8000 411.4500 ;
	    RECT 424.2000 410.4000 425.4000 410.5500 ;
	    RECT 474.6000 410.4000 475.8000 410.5500 ;
	    RECT 476.7000 409.5000 477.6000 411.9000 ;
	    RECT 484.2000 411.6000 485.4000 419.7000 ;
	    RECT 486.6000 413.7000 487.8000 419.7000 ;
	    RECT 489.0000 415.5000 490.2000 419.7000 ;
	    RECT 491.4000 415.5000 492.6000 419.7000 ;
	    RECT 493.8000 415.5000 495.0000 419.7000 ;
	    RECT 486.3000 411.6000 492.6000 412.8000 ;
	    RECT 481.5000 410.4000 485.4000 411.6000 ;
	    RECT 496.2000 410.4000 497.4000 419.7000 ;
	    RECT 498.6000 413.7000 499.8000 419.7000 ;
	    RECT 501.0000 412.5000 502.2000 419.7000 ;
	    RECT 503.4000 413.7000 504.6000 419.7000 ;
	    RECT 505.8000 412.5000 507.0000 419.7000 ;
	    RECT 508.2000 415.5000 509.4000 419.7000 ;
	    RECT 510.6000 415.5000 511.8000 419.7000 ;
	    RECT 513.0000 413.7000 514.2000 419.7000 ;
	    RECT 515.4000 412.8000 516.6000 419.7000 ;
	    RECT 517.8000 413.7000 519.0000 420.6000 ;
	    RECT 520.2000 414.6000 521.4000 419.7000 ;
	    RECT 520.2000 413.7000 521.7000 414.6000 ;
	    RECT 522.6000 413.7000 523.8000 419.7000 ;
	    RECT 537.0000 413.7000 538.2000 419.7000 ;
	    RECT 520.8000 412.8000 521.7000 413.7000 ;
	    RECT 513.6000 411.6000 519.9000 412.8000 ;
	    RECT 520.8000 411.9000 523.8000 412.8000 ;
	    RECT 501.0000 410.4000 504.9000 411.6000 ;
	    RECT 505.8000 410.7000 514.5000 411.6000 ;
	    RECT 519.0000 411.0000 519.9000 411.6000 ;
	    RECT 489.0000 409.5000 490.2000 409.8000 ;
	    RECT 474.6000 408.0000 475.8000 409.5000 ;
	    RECT 474.3000 406.8000 475.8000 408.0000 ;
	    RECT 476.7000 408.6000 490.2000 409.5000 ;
	    RECT 493.8000 409.5000 495.0000 409.8000 ;
	    RECT 505.8000 409.5000 506.7000 410.7000 ;
	    RECT 515.4000 409.8000 517.5000 410.7000 ;
	    RECT 519.0000 409.8000 521.4000 411.0000 ;
	    RECT 493.8000 408.6000 506.7000 409.5000 ;
	    RECT 508.2000 409.5000 517.5000 409.8000 ;
	    RECT 508.2000 408.9000 516.3000 409.5000 ;
	    RECT 508.2000 408.6000 509.4000 408.9000 ;
	    RECT 296.4000 401.7000 297.6000 402.0000 ;
	    RECT 296.4000 400.8000 303.0000 401.7000 ;
	    RECT 304.2000 401.4000 305.4000 402.6000 ;
	    RECT 301.8000 400.5000 303.0000 400.8000 ;
	    RECT 304.2000 400.2000 305.4000 400.5000 ;
	    RECT 282.6000 393.3000 283.8000 399.3000 ;
	    RECT 285.0000 398.1000 288.6000 399.3000 ;
	    RECT 292.2000 398.4000 293.7000 399.6000 ;
	    RECT 298.2000 398.4000 298.5000 399.6000 ;
	    RECT 299.4000 398.4000 300.6000 399.6000 ;
	    RECT 301.8000 399.3000 303.0000 399.6000 ;
	    RECT 307.5000 399.3000 308.7000 402.9000 ;
	    RECT 311.4000 402.3000 324.6000 403.5000 ;
	    RECT 316.5000 400.2000 321.0000 401.4000 ;
	    RECT 316.5000 399.3000 317.7000 400.2000 ;
	    RECT 301.8000 398.4000 308.7000 399.3000 ;
	    RECT 287.4000 393.3000 288.6000 398.1000 ;
	    RECT 313.8000 398.1000 317.7000 399.3000 ;
	    RECT 289.8000 393.3000 291.0000 397.5000 ;
	    RECT 292.2000 393.3000 293.4000 397.5000 ;
	    RECT 294.6000 393.3000 295.8000 397.5000 ;
	    RECT 297.0000 393.3000 298.2000 397.5000 ;
	    RECT 299.4000 393.3000 300.6000 396.3000 ;
	    RECT 301.8000 393.3000 303.0000 397.5000 ;
	    RECT 304.2000 393.3000 305.4000 396.3000 ;
	    RECT 306.6000 393.3000 307.8000 397.5000 ;
	    RECT 309.0000 393.3000 310.2000 397.5000 ;
	    RECT 311.4000 393.3000 312.6000 397.5000 ;
	    RECT 313.8000 393.3000 315.0000 398.1000 ;
	    RECT 318.6000 393.3000 319.8000 399.3000 ;
	    RECT 323.4000 393.3000 324.6000 402.3000 ;
	    RECT 328.2000 402.4500 329.4000 402.6000 ;
	    RECT 337.8000 402.4500 339.0000 402.6000 ;
	    RECT 328.2000 401.5500 339.0000 402.4500 ;
	    RECT 328.2000 401.4000 329.4000 401.5500 ;
	    RECT 337.8000 401.4000 339.0000 401.5500 ;
	    RECT 337.8000 393.3000 339.0000 400.5000 ;
	    RECT 474.3000 400.2000 475.5000 406.8000 ;
	    RECT 476.7000 405.9000 477.6000 408.6000 ;
	    RECT 512.7000 407.7000 513.9000 408.0000 ;
	    RECT 478.5000 406.8000 516.9000 407.7000 ;
	    RECT 517.8000 407.4000 519.0000 408.6000 ;
	    RECT 478.5000 406.5000 479.7000 406.8000 ;
	    RECT 476.4000 405.0000 477.6000 405.9000 ;
	    RECT 486.6000 405.0000 512.1000 405.9000 ;
	    RECT 476.4000 402.0000 477.3000 405.0000 ;
	    RECT 486.6000 404.1000 487.8000 405.0000 ;
	    RECT 513.0000 404.4000 514.2000 405.6000 ;
	    RECT 515.1000 405.0000 521.7000 405.9000 ;
	    RECT 520.5000 404.7000 521.7000 405.0000 ;
	    RECT 478.2000 402.9000 483.9000 404.1000 ;
	    RECT 476.4000 401.1000 478.2000 402.0000 ;
	    RECT 340.2000 399.4500 341.4000 399.6000 ;
	    RECT 371.4000 399.4500 372.6000 399.6000 ;
	    RECT 393.0000 399.4500 394.2000 399.6000 ;
	    RECT 340.2000 398.5500 394.2000 399.4500 ;
	    RECT 474.3000 399.0000 475.8000 400.2000 ;
	    RECT 340.2000 398.4000 341.4000 398.5500 ;
	    RECT 371.4000 398.4000 372.6000 398.5500 ;
	    RECT 393.0000 398.4000 394.2000 398.5500 ;
	    RECT 340.2000 397.2000 341.4000 397.5000 ;
	    RECT 340.2000 393.3000 341.4000 396.3000 ;
	    RECT 472.2000 393.3000 473.4000 396.3000 ;
	    RECT 474.6000 393.3000 475.8000 399.0000 ;
	    RECT 477.0000 393.3000 478.2000 401.1000 ;
	    RECT 482.7000 401.1000 483.9000 402.9000 ;
	    RECT 482.7000 400.2000 485.4000 401.1000 ;
	    RECT 484.2000 399.3000 485.4000 400.2000 ;
	    RECT 491.4000 399.6000 492.6000 403.8000 ;
	    RECT 496.2000 402.9000 501.0000 404.1000 ;
	    RECT 506.7000 402.9000 509.7000 404.1000 ;
	    RECT 522.6000 403.5000 523.8000 411.9000 ;
	    RECT 539.4000 403.5000 540.6000 419.7000 ;
	    RECT 673.8000 413.7000 675.0000 419.7000 ;
	    RECT 676.2000 412.5000 677.4000 419.7000 ;
	    RECT 678.6000 413.7000 679.8000 419.7000 ;
	    RECT 681.0000 412.8000 682.2000 419.7000 ;
	    RECT 683.4000 413.7000 684.6000 419.7000 ;
	    RECT 678.3000 411.9000 682.2000 412.8000 ;
	    RECT 621.0000 411.4500 622.2000 411.6000 ;
	    RECT 676.2000 411.4500 677.4000 411.6000 ;
	    RECT 621.0000 410.5500 677.4000 411.4500 ;
	    RECT 621.0000 410.4000 622.2000 410.5500 ;
	    RECT 676.2000 410.4000 677.4000 410.5500 ;
	    RECT 678.3000 409.5000 679.2000 411.9000 ;
	    RECT 685.8000 411.6000 687.0000 419.7000 ;
	    RECT 688.2000 413.7000 689.4000 419.7000 ;
	    RECT 690.6000 415.5000 691.8000 419.7000 ;
	    RECT 693.0000 415.5000 694.2000 419.7000 ;
	    RECT 695.4000 415.5000 696.6000 419.7000 ;
	    RECT 687.9000 411.6000 694.2000 412.8000 ;
	    RECT 683.1000 410.4000 687.0000 411.6000 ;
	    RECT 697.8000 410.4000 699.0000 419.7000 ;
	    RECT 700.2000 413.7000 701.4000 419.7000 ;
	    RECT 702.6000 412.5000 703.8000 419.7000 ;
	    RECT 705.0000 413.7000 706.2000 419.7000 ;
	    RECT 707.4000 412.5000 708.6000 419.7000 ;
	    RECT 709.8000 415.5000 711.0000 419.7000 ;
	    RECT 712.2000 415.5000 713.4000 419.7000 ;
	    RECT 714.6000 413.7000 715.8000 419.7000 ;
	    RECT 717.0000 412.8000 718.2000 419.7000 ;
	    RECT 719.4000 413.7000 720.6000 420.6000 ;
	    RECT 721.8000 414.6000 723.0000 419.7000 ;
	    RECT 721.8000 413.7000 723.3000 414.6000 ;
	    RECT 724.2000 413.7000 725.4000 419.7000 ;
	    RECT 738.6000 413.7000 739.8000 419.7000 ;
	    RECT 722.4000 412.8000 723.3000 413.7000 ;
	    RECT 715.2000 411.6000 721.5000 412.8000 ;
	    RECT 722.4000 411.9000 725.4000 412.8000 ;
	    RECT 702.6000 410.4000 706.5000 411.6000 ;
	    RECT 707.4000 410.7000 716.1000 411.6000 ;
	    RECT 720.6000 411.0000 721.5000 411.6000 ;
	    RECT 690.6000 409.5000 691.8000 409.8000 ;
	    RECT 616.2000 408.4500 617.4000 408.6000 ;
	    RECT 659.4000 408.4500 660.6000 408.6000 ;
	    RECT 616.2000 407.5500 660.6000 408.4500 ;
	    RECT 676.2000 408.0000 677.4000 409.5000 ;
	    RECT 616.2000 407.4000 617.4000 407.5500 ;
	    RECT 659.4000 407.4000 660.6000 407.5500 ;
	    RECT 675.9000 406.8000 677.4000 408.0000 ;
	    RECT 678.3000 408.6000 691.8000 409.5000 ;
	    RECT 695.4000 409.5000 696.6000 409.8000 ;
	    RECT 707.4000 409.5000 708.3000 410.7000 ;
	    RECT 717.0000 409.8000 719.1000 410.7000 ;
	    RECT 720.6000 409.8000 723.0000 411.0000 ;
	    RECT 695.4000 408.6000 708.3000 409.5000 ;
	    RECT 709.8000 409.5000 719.1000 409.8000 ;
	    RECT 709.8000 408.9000 717.9000 409.5000 ;
	    RECT 709.8000 408.6000 711.0000 408.9000 ;
	    RECT 495.6000 401.7000 496.8000 402.0000 ;
	    RECT 495.6000 400.8000 502.2000 401.7000 ;
	    RECT 503.4000 401.4000 504.6000 402.6000 ;
	    RECT 501.0000 400.5000 502.2000 400.8000 ;
	    RECT 503.4000 400.2000 504.6000 400.5000 ;
	    RECT 481.8000 393.3000 483.0000 399.3000 ;
	    RECT 484.2000 398.1000 487.8000 399.3000 ;
	    RECT 491.4000 398.4000 492.9000 399.6000 ;
	    RECT 497.4000 398.4000 497.7000 399.6000 ;
	    RECT 498.6000 398.4000 499.8000 399.6000 ;
	    RECT 501.0000 399.3000 502.2000 399.6000 ;
	    RECT 506.7000 399.3000 507.9000 402.9000 ;
	    RECT 510.6000 402.3000 523.8000 403.5000 ;
	    RECT 515.7000 400.2000 520.2000 401.4000 ;
	    RECT 515.7000 399.3000 516.9000 400.2000 ;
	    RECT 501.0000 398.4000 507.9000 399.3000 ;
	    RECT 486.6000 393.3000 487.8000 398.1000 ;
	    RECT 513.0000 398.1000 516.9000 399.3000 ;
	    RECT 489.0000 393.3000 490.2000 397.5000 ;
	    RECT 491.4000 393.3000 492.6000 397.5000 ;
	    RECT 493.8000 393.3000 495.0000 397.5000 ;
	    RECT 496.2000 393.3000 497.4000 397.5000 ;
	    RECT 498.6000 393.3000 499.8000 396.3000 ;
	    RECT 501.0000 393.3000 502.2000 397.5000 ;
	    RECT 503.4000 393.3000 504.6000 396.3000 ;
	    RECT 505.8000 393.3000 507.0000 397.5000 ;
	    RECT 508.2000 393.3000 509.4000 397.5000 ;
	    RECT 510.6000 393.3000 511.8000 397.5000 ;
	    RECT 513.0000 393.3000 514.2000 398.1000 ;
	    RECT 517.8000 393.3000 519.0000 399.3000 ;
	    RECT 522.6000 393.3000 523.8000 402.3000 ;
	    RECT 539.4000 402.4500 540.6000 402.6000 ;
	    RECT 585.0000 402.4500 586.2000 402.6000 ;
	    RECT 539.4000 401.5500 586.2000 402.4500 ;
	    RECT 539.4000 401.4000 540.6000 401.5500 ;
	    RECT 585.0000 401.4000 586.2000 401.5500 ;
	    RECT 599.4000 402.4500 600.6000 402.6000 ;
	    RECT 623.4000 402.4500 624.6000 402.6000 ;
	    RECT 599.4000 401.5500 624.6000 402.4500 ;
	    RECT 599.4000 401.4000 600.6000 401.5500 ;
	    RECT 623.4000 401.4000 624.6000 401.5500 ;
	    RECT 537.0000 398.4000 538.2000 399.6000 ;
	    RECT 537.0000 397.2000 538.2000 397.5000 ;
	    RECT 537.0000 393.3000 538.2000 396.3000 ;
	    RECT 539.4000 393.3000 540.6000 400.5000 ;
	    RECT 675.9000 400.2000 677.1000 406.8000 ;
	    RECT 678.3000 405.9000 679.2000 408.6000 ;
	    RECT 714.3000 407.7000 715.5000 408.0000 ;
	    RECT 680.1000 406.8000 718.5000 407.7000 ;
	    RECT 719.4000 407.4000 720.6000 408.6000 ;
	    RECT 680.1000 406.5000 681.3000 406.8000 ;
	    RECT 678.0000 405.0000 679.2000 405.9000 ;
	    RECT 688.2000 405.0000 713.7000 405.9000 ;
	    RECT 678.0000 402.0000 678.9000 405.0000 ;
	    RECT 688.2000 404.1000 689.4000 405.0000 ;
	    RECT 714.6000 404.4000 715.8000 405.6000 ;
	    RECT 716.7000 405.0000 723.3000 405.9000 ;
	    RECT 722.1000 404.7000 723.3000 405.0000 ;
	    RECT 679.8000 402.9000 685.5000 404.1000 ;
	    RECT 678.0000 401.1000 679.8000 402.0000 ;
	    RECT 675.9000 399.0000 677.4000 400.2000 ;
	    RECT 673.8000 393.3000 675.0000 396.3000 ;
	    RECT 676.2000 393.3000 677.4000 399.0000 ;
	    RECT 678.6000 393.3000 679.8000 401.1000 ;
	    RECT 684.3000 401.1000 685.5000 402.9000 ;
	    RECT 684.3000 400.2000 687.0000 401.1000 ;
	    RECT 685.8000 399.3000 687.0000 400.2000 ;
	    RECT 693.0000 399.6000 694.2000 403.8000 ;
	    RECT 697.8000 402.9000 702.6000 404.1000 ;
	    RECT 708.3000 402.9000 711.3000 404.1000 ;
	    RECT 724.2000 403.5000 725.4000 411.9000 ;
	    RECT 741.0000 403.5000 742.2000 419.7000 ;
	    RECT 767.4000 407.7000 768.6000 419.7000 ;
	    RECT 771.3000 408.6000 772.5000 419.7000 ;
	    RECT 773.7000 413.7000 774.9000 419.7000 ;
	    RECT 773.4000 410.4000 774.6000 411.6000 ;
	    RECT 773.7000 409.5000 774.6000 410.4000 ;
	    RECT 771.3000 407.7000 772.8000 408.6000 ;
	    RECT 769.8000 404.4000 771.0000 405.6000 ;
	    RECT 697.2000 401.7000 698.4000 402.0000 ;
	    RECT 697.2000 400.8000 703.8000 401.7000 ;
	    RECT 705.0000 401.4000 706.2000 402.6000 ;
	    RECT 702.6000 400.5000 703.8000 400.8000 ;
	    RECT 705.0000 400.2000 706.2000 400.5000 ;
	    RECT 683.4000 393.3000 684.6000 399.3000 ;
	    RECT 685.8000 398.1000 689.4000 399.3000 ;
	    RECT 693.0000 398.4000 694.5000 399.6000 ;
	    RECT 699.0000 398.4000 699.3000 399.6000 ;
	    RECT 700.2000 398.4000 701.4000 399.6000 ;
	    RECT 702.6000 399.3000 703.8000 399.6000 ;
	    RECT 708.3000 399.3000 709.5000 402.9000 ;
	    RECT 712.2000 402.3000 725.4000 403.5000 ;
	    RECT 769.8000 403.2000 771.0000 403.5000 ;
	    RECT 771.9000 402.6000 772.8000 407.7000 ;
	    RECT 774.6000 407.4000 775.8000 408.6000 ;
	    RECT 786.6000 403.5000 787.8000 419.7000 ;
	    RECT 789.0000 413.7000 790.2000 419.7000 ;
	    RECT 801.0000 419.4000 802.2000 420.6000 ;
	    RECT 808.2000 413.7000 809.4000 419.7000 ;
	    RECT 810.6000 406.5000 811.8000 419.7000 ;
	    RECT 813.0000 413.7000 814.2000 419.7000 ;
	    RECT 947.4000 413.7000 948.6000 419.7000 ;
	    RECT 949.8000 414.6000 951.0000 419.7000 ;
	    RECT 949.5000 413.7000 951.0000 414.6000 ;
	    RECT 952.2000 413.7000 953.4000 420.6000 ;
	    RECT 949.5000 412.8000 950.4000 413.7000 ;
	    RECT 954.6000 412.8000 955.8000 419.7000 ;
	    RECT 957.0000 413.7000 958.2000 419.7000 ;
	    RECT 959.4000 415.5000 960.6000 419.7000 ;
	    RECT 961.8000 415.5000 963.0000 419.7000 ;
	    RECT 947.4000 411.9000 950.4000 412.8000 ;
	    RECT 813.0000 409.5000 814.2000 409.8000 ;
	    RECT 813.0000 407.4000 814.2000 408.6000 ;
	    RECT 810.6000 405.4500 811.8000 405.6000 ;
	    RECT 945.0000 405.4500 946.2000 405.6000 ;
	    RECT 810.6000 404.5500 946.2000 405.4500 ;
	    RECT 810.6000 404.4000 811.8000 404.5500 ;
	    RECT 945.0000 404.4000 946.2000 404.5500 ;
	    RECT 947.4000 403.5000 948.6000 411.9000 ;
	    RECT 951.3000 411.6000 957.6000 412.8000 ;
	    RECT 964.2000 412.5000 965.4000 419.7000 ;
	    RECT 966.6000 413.7000 967.8000 419.7000 ;
	    RECT 969.0000 412.5000 970.2000 419.7000 ;
	    RECT 971.4000 413.7000 972.6000 419.7000 ;
	    RECT 951.3000 411.0000 952.2000 411.6000 ;
	    RECT 949.8000 409.8000 952.2000 411.0000 ;
	    RECT 956.7000 410.7000 965.4000 411.6000 ;
	    RECT 953.7000 409.8000 955.8000 410.7000 ;
	    RECT 953.7000 409.5000 963.0000 409.8000 ;
	    RECT 954.9000 408.9000 963.0000 409.5000 ;
	    RECT 961.8000 408.6000 963.0000 408.9000 ;
	    RECT 964.5000 409.5000 965.4000 410.7000 ;
	    RECT 966.3000 410.4000 970.2000 411.6000 ;
	    RECT 973.8000 410.4000 975.0000 419.7000 ;
	    RECT 976.2000 415.5000 977.4000 419.7000 ;
	    RECT 978.6000 415.5000 979.8000 419.7000 ;
	    RECT 981.0000 415.5000 982.2000 419.7000 ;
	    RECT 983.4000 413.7000 984.6000 419.7000 ;
	    RECT 978.6000 411.6000 984.9000 412.8000 ;
	    RECT 985.8000 411.6000 987.0000 419.7000 ;
	    RECT 988.2000 413.7000 989.4000 419.7000 ;
	    RECT 990.6000 412.8000 991.8000 419.7000 ;
	    RECT 993.0000 413.7000 994.2000 419.7000 ;
	    RECT 990.6000 411.9000 994.5000 412.8000 ;
	    RECT 995.4000 412.5000 996.6000 419.7000 ;
	    RECT 997.8000 413.7000 999.0000 419.7000 ;
	    RECT 985.8000 410.4000 989.7000 411.6000 ;
	    RECT 976.2000 409.5000 977.4000 409.8000 ;
	    RECT 964.5000 408.6000 977.4000 409.5000 ;
	    RECT 981.0000 409.5000 982.2000 409.8000 ;
	    RECT 993.6000 409.5000 994.5000 411.9000 ;
	    RECT 995.4000 410.4000 996.6000 411.6000 ;
	    RECT 981.0000 408.6000 994.5000 409.5000 ;
	    RECT 952.2000 407.4000 953.4000 408.6000 ;
	    RECT 957.3000 407.7000 958.5000 408.0000 ;
	    RECT 954.3000 406.8000 992.7000 407.7000 ;
	    RECT 991.5000 406.5000 992.7000 406.8000 ;
	    RECT 993.6000 405.9000 994.5000 408.6000 ;
	    RECT 995.4000 408.0000 996.6000 409.5000 ;
	    RECT 995.4000 406.8000 996.9000 408.0000 ;
	    RECT 949.5000 405.0000 956.1000 405.9000 ;
	    RECT 949.5000 404.7000 950.7000 405.0000 ;
	    RECT 957.0000 404.4000 958.2000 405.6000 ;
	    RECT 959.1000 405.0000 984.6000 405.9000 ;
	    RECT 993.6000 405.0000 994.8000 405.9000 ;
	    RECT 983.4000 404.1000 984.6000 405.0000 ;
	    RECT 717.3000 400.2000 721.8000 401.4000 ;
	    RECT 717.3000 399.3000 718.5000 400.2000 ;
	    RECT 702.6000 398.4000 709.5000 399.3000 ;
	    RECT 688.2000 393.3000 689.4000 398.1000 ;
	    RECT 714.6000 398.1000 718.5000 399.3000 ;
	    RECT 690.6000 393.3000 691.8000 397.5000 ;
	    RECT 693.0000 393.3000 694.2000 397.5000 ;
	    RECT 695.4000 393.3000 696.6000 397.5000 ;
	    RECT 697.8000 393.3000 699.0000 397.5000 ;
	    RECT 700.2000 393.3000 701.4000 396.3000 ;
	    RECT 702.6000 393.3000 703.8000 397.5000 ;
	    RECT 705.0000 393.3000 706.2000 396.3000 ;
	    RECT 707.4000 393.3000 708.6000 397.5000 ;
	    RECT 709.8000 393.3000 711.0000 397.5000 ;
	    RECT 712.2000 393.3000 713.4000 397.5000 ;
	    RECT 714.6000 393.3000 715.8000 398.1000 ;
	    RECT 719.4000 393.3000 720.6000 399.3000 ;
	    RECT 724.2000 393.3000 725.4000 402.3000 ;
	    RECT 741.0000 402.4500 742.2000 402.6000 ;
	    RECT 765.0000 402.4500 766.2000 402.6000 ;
	    RECT 741.0000 401.5500 766.2000 402.4500 ;
	    RECT 741.0000 401.4000 742.2000 401.5500 ;
	    RECT 765.0000 401.4000 766.2000 401.5500 ;
	    RECT 767.4000 401.4000 768.6000 402.6000 ;
	    RECT 769.5000 400.8000 769.8000 402.3000 ;
	    RECT 771.9000 401.4000 773.7000 402.6000 ;
	    RECT 774.6000 401.4000 775.8000 402.6000 ;
	    RECT 777.0000 402.4500 778.2000 402.6000 ;
	    RECT 786.6000 402.4500 787.8000 402.6000 ;
	    RECT 777.0000 401.5500 787.8000 402.4500 ;
	    RECT 777.0000 401.4000 778.2000 401.5500 ;
	    RECT 786.6000 401.4000 787.8000 401.5500 ;
	    RECT 801.0000 402.4500 802.2000 402.6000 ;
	    RECT 808.2000 402.4500 809.4000 402.6000 ;
	    RECT 801.0000 401.5500 809.4000 402.4500 ;
	    RECT 801.0000 401.4000 802.2000 401.5500 ;
	    RECT 808.2000 401.4000 809.4000 401.5500 ;
	    RECT 738.6000 398.4000 739.8000 399.6000 ;
	    RECT 738.6000 397.2000 739.8000 397.5000 ;
	    RECT 738.6000 393.3000 739.8000 396.3000 ;
	    RECT 741.0000 393.3000 742.2000 400.5000 ;
	    RECT 767.7000 399.3000 773.1000 399.9000 ;
	    RECT 774.6000 399.3000 775.5000 400.5000 ;
	    RECT 767.4000 399.0000 773.4000 399.3000 ;
	    RECT 767.4000 393.3000 768.6000 399.0000 ;
	    RECT 769.8000 393.3000 771.0000 398.1000 ;
	    RECT 772.2000 393.3000 773.4000 399.0000 ;
	    RECT 774.6000 393.3000 775.8000 399.3000 ;
	    RECT 786.6000 393.3000 787.8000 400.5000 ;
	    RECT 808.2000 400.2000 809.4000 400.5000 ;
	    RECT 789.0000 399.4500 790.2000 399.6000 ;
	    RECT 805.8000 399.4500 807.0000 399.6000 ;
	    RECT 789.0000 398.5500 807.0000 399.4500 ;
	    RECT 810.6000 399.3000 811.8000 403.5000 ;
	    RECT 947.4000 402.3000 960.6000 403.5000 ;
	    RECT 961.5000 402.9000 964.5000 404.1000 ;
	    RECT 970.2000 402.9000 975.0000 404.1000 ;
	    RECT 789.0000 398.4000 790.2000 398.5500 ;
	    RECT 805.8000 398.4000 807.0000 398.5500 ;
	    RECT 789.0000 397.2000 790.2000 397.5000 ;
	    RECT 789.0000 393.3000 790.2000 396.3000 ;
	    RECT 808.2000 393.3000 809.4000 399.3000 ;
	    RECT 810.6000 398.4000 813.3000 399.3000 ;
	    RECT 812.1000 393.3000 813.3000 398.4000 ;
	    RECT 947.4000 393.3000 948.6000 402.3000 ;
	    RECT 951.0000 400.2000 955.5000 401.4000 ;
	    RECT 954.3000 399.3000 955.5000 400.2000 ;
	    RECT 963.3000 399.3000 964.5000 402.9000 ;
	    RECT 966.6000 401.4000 967.8000 402.6000 ;
	    RECT 974.4000 401.7000 975.6000 402.0000 ;
	    RECT 969.0000 400.8000 975.6000 401.7000 ;
	    RECT 969.0000 400.5000 970.2000 400.8000 ;
	    RECT 966.6000 400.2000 967.8000 400.5000 ;
	    RECT 978.6000 399.6000 979.8000 403.8000 ;
	    RECT 987.3000 402.9000 993.0000 404.1000 ;
	    RECT 987.3000 401.1000 988.5000 402.9000 ;
	    RECT 993.9000 402.0000 994.8000 405.0000 ;
	    RECT 969.0000 399.3000 970.2000 399.6000 ;
	    RECT 952.2000 393.3000 953.4000 399.3000 ;
	    RECT 954.3000 398.1000 958.2000 399.3000 ;
	    RECT 963.3000 398.4000 970.2000 399.3000 ;
	    RECT 971.4000 398.4000 972.6000 399.6000 ;
	    RECT 973.5000 398.4000 973.8000 399.6000 ;
	    RECT 978.3000 398.4000 979.8000 399.6000 ;
	    RECT 985.8000 400.2000 988.5000 401.1000 ;
	    RECT 993.0000 401.1000 994.8000 402.0000 ;
	    RECT 985.8000 399.3000 987.0000 400.2000 ;
	    RECT 957.0000 393.3000 958.2000 398.1000 ;
	    RECT 983.4000 398.1000 987.0000 399.3000 ;
	    RECT 959.4000 393.3000 960.6000 397.5000 ;
	    RECT 961.8000 393.3000 963.0000 397.5000 ;
	    RECT 964.2000 393.3000 965.4000 397.5000 ;
	    RECT 966.6000 393.3000 967.8000 396.3000 ;
	    RECT 969.0000 393.3000 970.2000 397.5000 ;
	    RECT 971.4000 393.3000 972.6000 396.3000 ;
	    RECT 973.8000 393.3000 975.0000 397.5000 ;
	    RECT 976.2000 393.3000 977.4000 397.5000 ;
	    RECT 978.6000 393.3000 979.8000 397.5000 ;
	    RECT 981.0000 393.3000 982.2000 397.5000 ;
	    RECT 983.4000 393.3000 984.6000 398.1000 ;
	    RECT 988.2000 393.3000 989.4000 399.3000 ;
	    RECT 993.0000 393.3000 994.2000 401.1000 ;
	    RECT 995.7000 400.2000 996.9000 406.8000 ;
	    RECT 1012.2000 403.5000 1013.4000 419.7000 ;
	    RECT 1014.6000 413.7000 1015.8000 419.7000 ;
	    RECT 1041.9000 413.7000 1043.1000 419.7000 ;
	    RECT 1042.2001 410.4000 1043.4000 411.6000 ;
	    RECT 1042.2001 409.5000 1043.1000 410.4000 ;
	    RECT 1044.3000 408.6000 1045.5000 419.7000 ;
	    RECT 1041.0000 407.4000 1042.2001 408.6000 ;
	    RECT 1044.0000 407.7000 1045.5000 408.6000 ;
	    RECT 1048.2001 407.7000 1049.4000 419.7000 ;
	    RECT 1060.2001 413.7000 1061.4000 419.7000 ;
	    RECT 1044.0000 402.6000 1044.9000 407.7000 ;
	    RECT 1045.8000 405.4500 1047.0000 405.6000 ;
	    RECT 1045.8000 404.5500 1051.6500 405.4500 ;
	    RECT 1045.8000 404.4000 1047.0000 404.5500 ;
	    RECT 1045.8000 403.2000 1047.0000 403.5000 ;
	    RECT 1009.8000 402.4500 1011.0000 402.6000 ;
	    RECT 1012.2000 402.4500 1013.4000 402.6000 ;
	    RECT 1009.8000 401.5500 1013.4000 402.4500 ;
	    RECT 1009.8000 401.4000 1011.0000 401.5500 ;
	    RECT 1012.2000 401.4000 1013.4000 401.5500 ;
	    RECT 1036.2001 402.4500 1037.4000 402.6000 ;
	    RECT 1041.0000 402.4500 1042.2001 402.6000 ;
	    RECT 1036.2001 401.5500 1042.2001 402.4500 ;
	    RECT 1036.2001 401.4000 1037.4000 401.5500 ;
	    RECT 1041.0000 401.4000 1042.2001 401.5500 ;
	    RECT 1043.1000 401.4000 1044.9000 402.6000 ;
	    RECT 1047.0000 400.8000 1047.3000 402.3000 ;
	    RECT 1048.2001 401.4000 1049.4000 402.6000 ;
	    RECT 1050.7500 402.4500 1051.6500 404.5500 ;
	    RECT 1062.6000 403.5000 1063.8000 419.7000 ;
	    RECT 1067.4000 419.4000 1068.6000 420.6000 ;
	    RECT 1103.4000 408.6000 1104.6000 419.7000 ;
	    RECT 1105.8000 409.8000 1107.3000 419.7000 ;
	    RECT 1105.5000 408.6000 1106.7001 408.9000 ;
	    RECT 1103.4000 407.7000 1106.7001 408.6000 ;
	    RECT 1110.0000 408.6000 1112.4000 419.7000 ;
	    RECT 1115.1000 409.8000 1116.6000 419.7000 ;
	    RECT 1115.4000 408.6000 1116.6000 408.9000 ;
	    RECT 1117.8000 408.6000 1119.0000 419.7000 ;
	    RECT 1110.0000 407.7000 1113.0000 408.6000 ;
	    RECT 1115.4000 407.7000 1119.0000 408.6000 ;
	    RECT 1156.2001 407.7000 1157.4000 419.7000 ;
	    RECT 1160.1000 407.7000 1163.1000 419.7000 ;
	    RECT 1165.8000 407.7000 1167.0000 419.7000 ;
	    RECT 1189.8000 407.7000 1191.0000 419.7000 ;
	    RECT 1193.7001 408.6000 1194.9000 419.7000 ;
	    RECT 1196.1000 413.7000 1197.3000 419.7000 ;
	    RECT 1195.8000 410.4000 1197.0000 411.6000 ;
	    RECT 1196.1000 409.5000 1197.0000 410.4000 ;
	    RECT 1193.7001 407.7000 1195.2001 408.6000 ;
	    RECT 1105.8000 406.8000 1106.7001 407.7000 ;
	    RECT 1105.8000 405.9000 1110.9000 406.8000 ;
	    RECT 1112.1000 406.5000 1113.0000 407.7000 ;
	    RECT 1109.7001 405.6000 1110.9000 405.9000 ;
	    RECT 1113.0000 405.4500 1114.2001 405.6000 ;
	    RECT 1146.6000 405.4500 1147.8000 405.6000 ;
	    RECT 1106.4000 404.7000 1107.6000 405.0000 ;
	    RECT 1106.4000 403.8000 1110.3000 404.7000 ;
	    RECT 1109.4000 402.9000 1110.3000 403.8000 ;
	    RECT 1111.5000 403.5000 1112.1000 404.7000 ;
	    RECT 1113.0000 404.5500 1147.8000 405.4500 ;
	    RECT 1113.0000 404.4000 1114.2001 404.5500 ;
	    RECT 1146.6000 404.4000 1147.8000 404.5500 ;
	    RECT 1149.0000 405.4500 1150.2001 405.6000 ;
	    RECT 1158.6000 405.4500 1159.8000 405.6000 ;
	    RECT 1149.0000 404.5500 1159.8000 405.4500 ;
	    RECT 1149.0000 404.4000 1150.2001 404.5500 ;
	    RECT 1158.6000 404.4000 1159.8000 404.5500 ;
	    RECT 1161.0000 403.5000 1161.9000 407.7000 ;
	    RECT 1163.4000 404.4000 1164.6000 405.6000 ;
	    RECT 1192.2001 404.4000 1193.4000 405.6000 ;
	    RECT 1165.8000 403.5000 1167.0000 403.8000 ;
	    RECT 1062.6000 402.4500 1063.8000 402.6000 ;
	    RECT 1050.7500 401.5500 1063.8000 402.4500 ;
	    RECT 1062.6000 401.4000 1063.8000 401.5500 ;
	    RECT 1079.4000 402.4500 1080.6000 402.6000 ;
	    RECT 1103.4000 402.4500 1104.6000 402.6000 ;
	    RECT 1079.4000 401.5500 1104.6000 402.4500 ;
	    RECT 1079.4000 401.4000 1080.6000 401.5500 ;
	    RECT 1103.4000 401.4000 1104.6000 401.5500 ;
	    RECT 1105.5000 402.3000 1105.8000 402.6000 ;
	    RECT 1105.5000 401.4000 1108.5000 402.3000 ;
	    RECT 1109.4000 401.7000 1110.6000 402.9000 ;
	    RECT 1107.6000 400.8000 1108.5000 401.4000 ;
	    RECT 995.4000 399.0000 996.9000 400.2000 ;
	    RECT 995.4000 393.3000 996.6000 399.0000 ;
	    RECT 997.8000 393.3000 999.0000 396.3000 ;
	    RECT 1012.2000 393.3000 1013.4000 400.5000 ;
	    RECT 1014.6000 398.4000 1015.8000 399.6000 ;
	    RECT 1041.3000 399.3000 1042.2001 400.5000 ;
	    RECT 1043.7001 399.3000 1049.1000 399.9000 ;
	    RECT 1014.6000 397.2000 1015.8000 397.5000 ;
	    RECT 1014.6000 393.3000 1015.8000 396.3000 ;
	    RECT 1041.0000 393.3000 1042.2001 399.3000 ;
	    RECT 1043.4000 399.0000 1049.4000 399.3000 ;
	    RECT 1043.4000 393.3000 1044.6000 399.0000 ;
	    RECT 1045.8000 393.3000 1047.0000 398.1000 ;
	    RECT 1048.2001 393.3000 1049.4000 399.0000 ;
	    RECT 1060.2001 398.4000 1061.4000 399.6000 ;
	    RECT 1060.2001 397.2000 1061.4000 397.5000 ;
	    RECT 1060.2001 393.3000 1061.4000 396.3000 ;
	    RECT 1062.6000 393.3000 1063.8000 400.5000 ;
	    RECT 1105.5000 400.2000 1106.7001 400.5000 ;
	    RECT 1103.4000 399.3000 1106.7001 400.2000 ;
	    RECT 1107.6000 399.9000 1110.6000 400.8000 ;
	    RECT 1108.2001 399.6000 1110.6000 399.9000 ;
	    RECT 1103.4000 393.3000 1104.6000 399.3000 ;
	    RECT 1111.5000 398.7000 1112.4000 403.5000 ;
	    RECT 1158.6000 403.2000 1159.8000 403.5000 ;
	    RECT 1163.4000 403.2000 1164.6000 403.5000 ;
	    RECT 1192.2001 403.2000 1193.4000 403.5000 ;
	    RECT 1194.3000 402.6000 1195.2001 407.7000 ;
	    RECT 1197.0000 407.4000 1198.2001 408.6000 ;
	    RECT 1209.0000 405.4500 1210.2001 405.6000 ;
	    RECT 1199.5500 404.5500 1210.2001 405.4500 ;
	    RECT 1113.6000 401.4000 1114.8000 402.6000 ;
	    RECT 1116.6000 401.4000 1116.9000 402.6000 ;
	    RECT 1117.8000 401.4000 1119.0000 402.6000 ;
	    RECT 1141.8000 402.4500 1143.0000 402.6000 ;
	    RECT 1156.2001 402.4500 1157.4000 402.6000 ;
	    RECT 1141.8000 401.5500 1157.4000 402.4500 ;
	    RECT 1141.8000 401.4000 1143.0000 401.5500 ;
	    RECT 1156.2001 401.4000 1157.4000 401.5500 ;
	    RECT 1113.6000 400.8000 1114.5000 401.4000 ;
	    RECT 1158.3000 400.8000 1158.6000 402.3000 ;
	    RECT 1161.0000 401.4000 1162.2001 402.6000 ;
	    RECT 1163.1000 401.4000 1164.6000 402.3000 ;
	    RECT 1165.8000 401.4000 1167.0000 402.6000 ;
	    RECT 1189.8000 401.4000 1191.0000 402.6000 ;
	    RECT 1113.3000 399.6000 1114.5000 400.8000 ;
	    RECT 1115.4000 400.2000 1116.6000 400.5000 ;
	    RECT 1115.4000 399.3000 1119.0000 400.2000 ;
	    RECT 1156.5000 399.3000 1161.9000 399.9000 ;
	    RECT 1163.7001 399.3000 1164.6000 401.4000 ;
	    RECT 1191.9000 400.8000 1192.2001 402.3000 ;
	    RECT 1194.3000 401.4000 1196.1000 402.6000 ;
	    RECT 1197.0000 402.4500 1198.2001 402.6000 ;
	    RECT 1199.5500 402.4500 1200.4501 404.5500 ;
	    RECT 1209.0000 404.4000 1210.2001 404.5500 ;
	    RECT 1211.4000 403.5000 1212.6000 419.7000 ;
	    RECT 1213.8000 413.7000 1215.0000 419.7000 ;
	    RECT 1238.7001 413.7000 1239.9000 419.7000 ;
	    RECT 1239.0000 410.4000 1240.2001 411.6000 ;
	    RECT 1239.0000 409.5000 1239.9000 410.4000 ;
	    RECT 1241.1000 408.6000 1242.3000 419.7000 ;
	    RECT 1237.8000 407.4000 1239.0000 408.6000 ;
	    RECT 1240.8000 407.7000 1242.3000 408.6000 ;
	    RECT 1245.0000 407.7000 1246.2001 419.7000 ;
	    RECT 1273.8000 407.7000 1275.0000 419.7000 ;
	    RECT 1277.7001 407.7000 1280.7001 419.7000 ;
	    RECT 1283.4000 407.7000 1284.6000 419.7000 ;
	    RECT 1297.8000 413.7000 1299.0000 419.7000 ;
	    RECT 1240.8000 402.6000 1241.7001 407.7000 ;
	    RECT 1242.6000 404.4000 1243.8000 405.6000 ;
	    RECT 1276.2001 404.4000 1277.4000 405.6000 ;
	    RECT 1278.6000 403.5000 1279.5000 407.7000 ;
	    RECT 1281.0000 404.4000 1282.2001 405.6000 ;
	    RECT 1283.4000 403.5000 1284.6000 403.8000 ;
	    RECT 1300.2001 403.5000 1301.4000 419.7000 ;
	    RECT 1319.4000 413.7000 1320.6000 419.7000 ;
	    RECT 1321.8000 406.5000 1323.0000 419.7000 ;
	    RECT 1324.2001 413.7000 1325.4000 419.7000 ;
	    RECT 1329.0000 419.4000 1330.2001 420.6000 ;
	    RECT 1351.5000 413.7000 1352.7001 419.7000 ;
	    RECT 1351.8000 410.4000 1353.0000 411.6000 ;
	    RECT 1324.2001 409.5000 1325.4000 409.8000 ;
	    RECT 1351.8000 409.5000 1352.7001 410.4000 ;
	    RECT 1353.9000 408.6000 1355.1000 419.7000 ;
	    RECT 1324.2001 408.4500 1325.4000 408.6000 ;
	    RECT 1341.0000 408.4500 1342.2001 408.6000 ;
	    RECT 1324.2001 407.5500 1342.2001 408.4500 ;
	    RECT 1324.2001 407.4000 1325.4000 407.5500 ;
	    RECT 1341.0000 407.4000 1342.2001 407.5500 ;
	    RECT 1350.6000 407.4000 1351.8000 408.6000 ;
	    RECT 1353.6000 407.7000 1355.1000 408.6000 ;
	    RECT 1357.8000 407.7000 1359.0000 419.7000 ;
	    RECT 1389.0000 413.7000 1390.2001 419.7000 ;
	    RECT 1391.4000 413.7000 1392.6000 419.7000 ;
	    RECT 1393.8000 414.3000 1395.0000 419.7000 ;
	    RECT 1391.7001 413.4000 1392.6000 413.7000 ;
	    RECT 1396.2001 413.7000 1397.4000 419.7000 ;
	    RECT 1396.2001 413.4000 1397.1000 413.7000 ;
	    RECT 1391.7001 412.5000 1397.1000 413.4000 ;
	    RECT 1393.8000 410.4000 1395.0000 411.6000 ;
	    RECT 1396.2001 409.5000 1397.1000 412.5000 ;
	    RECT 1393.8000 409.2000 1395.0000 409.5000 ;
	    RECT 1360.2001 408.4500 1361.4000 408.6000 ;
	    RECT 1386.6000 408.4500 1387.8000 408.6000 ;
	    RECT 1389.0000 408.4500 1390.2001 408.6000 ;
	    RECT 1321.8000 405.4500 1323.0000 405.6000 ;
	    RECT 1345.8000 405.4500 1347.0000 405.6000 ;
	    RECT 1321.8000 404.5500 1347.0000 405.4500 ;
	    RECT 1321.8000 404.4000 1323.0000 404.5500 ;
	    RECT 1345.8000 404.4000 1347.0000 404.5500 ;
	    RECT 1242.6000 403.2000 1243.8000 403.5000 ;
	    RECT 1276.2001 403.2000 1277.4000 403.5000 ;
	    RECT 1281.0000 403.2000 1282.2001 403.5000 ;
	    RECT 1197.0000 401.5500 1200.4501 402.4500 ;
	    RECT 1201.8000 402.4500 1203.0000 402.6000 ;
	    RECT 1211.4000 402.4500 1212.6000 402.6000 ;
	    RECT 1201.8000 401.5500 1212.6000 402.4500 ;
	    RECT 1197.0000 401.4000 1198.2001 401.5500 ;
	    RECT 1201.8000 401.4000 1203.0000 401.5500 ;
	    RECT 1211.4000 401.4000 1212.6000 401.5500 ;
	    RECT 1233.0000 402.4500 1234.2001 402.6000 ;
	    RECT 1237.8000 402.4500 1239.0000 402.6000 ;
	    RECT 1233.0000 401.5500 1239.0000 402.4500 ;
	    RECT 1233.0000 401.4000 1234.2001 401.5500 ;
	    RECT 1237.8000 401.4000 1239.0000 401.5500 ;
	    RECT 1239.9000 401.4000 1241.7001 402.6000 ;
	    RECT 1245.0000 402.4500 1246.2001 402.6000 ;
	    RECT 1271.4000 402.4500 1272.6000 402.6000 ;
	    RECT 1243.8000 400.8000 1244.1000 402.3000 ;
	    RECT 1245.0000 401.5500 1272.6000 402.4500 ;
	    RECT 1245.0000 401.4000 1246.2001 401.5500 ;
	    RECT 1271.4000 401.4000 1272.6000 401.5500 ;
	    RECT 1273.8000 401.4000 1275.0000 402.6000 ;
	    RECT 1275.9000 400.8000 1276.2001 402.3000 ;
	    RECT 1278.6000 401.4000 1279.8000 402.6000 ;
	    RECT 1283.4000 402.4500 1284.6000 402.6000 ;
	    RECT 1285.8000 402.4500 1287.0000 402.6000 ;
	    RECT 1280.7001 401.4000 1282.2001 402.3000 ;
	    RECT 1283.4000 401.5500 1287.0000 402.4500 ;
	    RECT 1283.4000 401.4000 1284.6000 401.5500 ;
	    RECT 1285.8000 401.4000 1287.0000 401.5500 ;
	    RECT 1300.2001 402.4500 1301.4000 402.6000 ;
	    RECT 1314.6000 402.4500 1315.8000 402.6000 ;
	    RECT 1319.4000 402.4500 1320.6000 402.6000 ;
	    RECT 1300.2001 401.5500 1313.2500 402.4500 ;
	    RECT 1300.2001 401.4000 1301.4000 401.5500 ;
	    RECT 1190.1000 399.3000 1195.5000 399.9000 ;
	    RECT 1197.0000 399.3000 1197.9000 400.5000 ;
	    RECT 1105.8000 393.3000 1107.3000 398.4000 ;
	    RECT 1110.0000 393.3000 1112.4000 398.7000 ;
	    RECT 1115.1000 393.3000 1116.6000 398.4000 ;
	    RECT 1117.8000 393.3000 1119.0000 399.3000 ;
	    RECT 1156.2001 399.0000 1162.2001 399.3000 ;
	    RECT 1156.2001 393.3000 1157.4000 399.0000 ;
	    RECT 1158.6000 393.3000 1159.8000 398.1000 ;
	    RECT 1161.0000 394.2000 1162.2001 399.0000 ;
	    RECT 1163.4000 395.1000 1164.6000 399.3000 ;
	    RECT 1165.8000 394.2000 1167.0000 399.3000 ;
	    RECT 1161.0000 393.3000 1167.0000 394.2000 ;
	    RECT 1189.8000 399.0000 1195.8000 399.3000 ;
	    RECT 1189.8000 393.3000 1191.0000 399.0000 ;
	    RECT 1192.2001 393.3000 1193.4000 398.1000 ;
	    RECT 1194.6000 393.3000 1195.8000 399.0000 ;
	    RECT 1197.0000 393.3000 1198.2001 399.3000 ;
	    RECT 1211.4000 393.3000 1212.6000 400.5000 ;
	    RECT 1213.8000 399.4500 1215.0000 399.6000 ;
	    RECT 1218.6000 399.4500 1219.8000 399.6000 ;
	    RECT 1213.8000 398.5500 1219.8000 399.4500 ;
	    RECT 1238.1000 399.3000 1239.0000 400.5000 ;
	    RECT 1240.5000 399.3000 1245.9000 399.9000 ;
	    RECT 1274.1000 399.3000 1279.5000 399.9000 ;
	    RECT 1281.3000 399.3000 1282.2001 401.4000 ;
	    RECT 1293.0000 399.4500 1294.2001 399.6000 ;
	    RECT 1297.8000 399.4500 1299.0000 399.6000 ;
	    RECT 1213.8000 398.4000 1215.0000 398.5500 ;
	    RECT 1218.6000 398.4000 1219.8000 398.5500 ;
	    RECT 1213.8000 397.2000 1215.0000 397.5000 ;
	    RECT 1213.8000 393.3000 1215.0000 396.3000 ;
	    RECT 1237.8000 393.3000 1239.0000 399.3000 ;
	    RECT 1240.2001 399.0000 1246.2001 399.3000 ;
	    RECT 1240.2001 393.3000 1241.4000 399.0000 ;
	    RECT 1242.6000 393.3000 1243.8000 398.1000 ;
	    RECT 1245.0000 393.3000 1246.2001 399.0000 ;
	    RECT 1273.8000 399.0000 1279.8000 399.3000 ;
	    RECT 1273.8000 393.3000 1275.0000 399.0000 ;
	    RECT 1276.2001 393.3000 1277.4000 398.1000 ;
	    RECT 1278.6000 394.2000 1279.8000 399.0000 ;
	    RECT 1281.0000 395.1000 1282.2001 399.3000 ;
	    RECT 1283.4000 394.2000 1284.6000 399.3000 ;
	    RECT 1293.0000 398.5500 1299.0000 399.4500 ;
	    RECT 1293.0000 398.4000 1294.2001 398.5500 ;
	    RECT 1297.8000 398.4000 1299.0000 398.5500 ;
	    RECT 1297.8000 397.2000 1299.0000 397.5000 ;
	    RECT 1278.6000 393.3000 1284.6000 394.2000 ;
	    RECT 1297.8000 393.3000 1299.0000 396.3000 ;
	    RECT 1300.2001 393.3000 1301.4000 400.5000 ;
	    RECT 1312.3500 399.4500 1313.2500 401.5500 ;
	    RECT 1314.6000 401.5500 1320.6000 402.4500 ;
	    RECT 1314.6000 401.4000 1315.8000 401.5500 ;
	    RECT 1319.4000 401.4000 1320.6000 401.5500 ;
	    RECT 1319.4000 400.2000 1320.6000 400.5000 ;
	    RECT 1317.0000 399.4500 1318.2001 399.6000 ;
	    RECT 1312.3500 398.5500 1318.2001 399.4500 ;
	    RECT 1321.8000 399.3000 1323.0000 403.5000 ;
	    RECT 1353.6000 402.6000 1354.5000 407.7000 ;
	    RECT 1360.2001 407.5500 1390.2001 408.4500 ;
	    RECT 1360.2001 407.4000 1361.4000 407.5500 ;
	    RECT 1386.6000 407.4000 1387.8000 407.5500 ;
	    RECT 1389.0000 407.4000 1390.2001 407.5500 ;
	    RECT 1396.2001 408.4500 1397.4000 408.6000 ;
	    RECT 1403.4000 408.4500 1404.6000 408.6000 ;
	    RECT 1396.2001 407.5500 1404.6000 408.4500 ;
	    RECT 1422.6000 407.7000 1423.8000 419.7000 ;
	    RECT 1426.5000 408.6000 1427.7001 419.7000 ;
	    RECT 1428.9000 413.7000 1430.1000 419.7000 ;
	    RECT 1428.6000 410.4000 1429.8000 411.6000 ;
	    RECT 1428.9000 409.5000 1429.8000 410.4000 ;
	    RECT 1426.5000 407.7000 1428.0000 408.6000 ;
	    RECT 1396.2001 407.4000 1397.4000 407.5500 ;
	    RECT 1403.4000 407.4000 1404.6000 407.5500 ;
	    RECT 1389.0000 406.2000 1390.2001 406.5000 ;
	    RECT 1355.4000 405.4500 1356.6000 405.6000 ;
	    RECT 1367.4000 405.4500 1368.6000 405.6000 ;
	    RECT 1355.4000 404.5500 1368.6000 405.4500 ;
	    RECT 1355.4000 404.4000 1356.6000 404.5500 ;
	    RECT 1367.4000 404.4000 1368.6000 404.5500 ;
	    RECT 1391.4000 404.4000 1392.6000 405.6000 ;
	    RECT 1393.5000 404.4000 1393.8000 405.6000 ;
	    RECT 1355.4000 403.2000 1356.6000 403.5000 ;
	    RECT 1396.2001 402.6000 1397.1000 406.5000 ;
	    RECT 1425.0000 404.4000 1426.2001 405.6000 ;
	    RECT 1425.0000 403.2000 1426.2001 403.5000 ;
	    RECT 1427.1000 402.6000 1428.0000 407.7000 ;
	    RECT 1429.8000 408.4500 1431.0000 408.6000 ;
	    RECT 1439.4000 408.4500 1440.6000 408.6000 ;
	    RECT 1429.8000 407.5500 1440.6000 408.4500 ;
	    RECT 1429.8000 407.4000 1431.0000 407.5500 ;
	    RECT 1439.4000 407.4000 1440.6000 407.5500 ;
	    RECT 1444.2001 403.5000 1445.4000 419.7000 ;
	    RECT 1446.6000 413.7000 1447.8000 419.7000 ;
	    RECT 1461.0000 419.4000 1462.2001 420.6000 ;
	    RECT 1465.8000 413.7000 1467.0000 419.7000 ;
	    RECT 1465.8000 409.5000 1467.0000 409.8000 ;
	    RECT 1461.0000 408.4500 1462.2001 408.6000 ;
	    RECT 1465.8000 408.4500 1467.0000 408.6000 ;
	    RECT 1461.0000 407.5500 1467.0000 408.4500 ;
	    RECT 1461.0000 407.4000 1462.2001 407.5500 ;
	    RECT 1465.8000 407.4000 1467.0000 407.5500 ;
	    RECT 1468.2001 406.5000 1469.4000 419.7000 ;
	    RECT 1470.6000 413.7000 1471.8000 419.7000 ;
	    RECT 1465.8000 405.4500 1467.0000 405.6000 ;
	    RECT 1468.2001 405.4500 1469.4000 405.6000 ;
	    RECT 1465.8000 404.5500 1469.4000 405.4500 ;
	    RECT 1465.8000 404.4000 1467.0000 404.5500 ;
	    RECT 1468.2001 404.4000 1469.4000 404.5500 ;
	    RECT 1485.0000 403.5000 1486.2001 419.7000 ;
	    RECT 1487.4000 413.7000 1488.6000 419.7000 ;
	    RECT 1511.4000 413.7000 1512.6000 419.7000 ;
	    RECT 1513.8000 414.3000 1515.0000 419.7000 ;
	    RECT 1511.7001 413.4000 1512.6000 413.7000 ;
	    RECT 1516.2001 413.7000 1517.4000 419.7000 ;
	    RECT 1518.6000 413.7000 1519.8000 419.7000 ;
	    RECT 1516.2001 413.4000 1517.1000 413.7000 ;
	    RECT 1511.7001 412.5000 1517.1000 413.4000 ;
	    RECT 1511.7001 409.5000 1512.6000 412.5000 ;
	    RECT 1513.8000 411.4500 1515.0000 411.6000 ;
	    RECT 1521.0000 411.4500 1522.2001 411.6000 ;
	    RECT 1513.8000 410.5500 1522.2001 411.4500 ;
	    RECT 1513.8000 410.4000 1515.0000 410.5500 ;
	    RECT 1521.0000 410.4000 1522.2001 410.5500 ;
	    RECT 1513.8000 409.2000 1515.0000 409.5000 ;
	    RECT 1506.6000 408.4500 1507.8000 408.6000 ;
	    RECT 1511.4000 408.4500 1512.6000 408.6000 ;
	    RECT 1506.6000 407.5500 1512.6000 408.4500 ;
	    RECT 1506.6000 407.4000 1507.8000 407.5500 ;
	    RECT 1511.4000 407.4000 1512.6000 407.5500 ;
	    RECT 1518.6000 407.4000 1519.8000 408.6000 ;
	    RECT 1542.6000 407.7000 1543.8000 419.7000 ;
	    RECT 1545.0000 408.6000 1546.2001 419.7000 ;
	    RECT 1547.4000 409.5000 1548.6000 419.7000 ;
	    RECT 1549.8000 408.6000 1551.0000 419.7000 ;
	    RECT 1545.0000 407.7000 1551.0000 408.6000 ;
	    RECT 1542.9000 406.5000 1543.8000 407.7000 ;
	    RECT 1350.6000 401.4000 1351.8000 402.6000 ;
	    RECT 1352.7001 401.4000 1354.5000 402.6000 ;
	    RECT 1356.6000 400.8000 1356.9000 402.3000 ;
	    RECT 1357.8000 401.4000 1359.0000 402.6000 ;
	    RECT 1394.7001 402.3000 1397.1000 402.6000 ;
	    RECT 1350.9000 399.3000 1351.8000 400.5000 ;
	    RECT 1353.3000 399.3000 1358.7001 399.9000 ;
	    RECT 1317.0000 398.4000 1318.2001 398.5500 ;
	    RECT 1319.4000 393.3000 1320.6000 399.3000 ;
	    RECT 1321.8000 398.4000 1324.5000 399.3000 ;
	    RECT 1323.3000 393.3000 1324.5000 398.4000 ;
	    RECT 1350.6000 393.3000 1351.8000 399.3000 ;
	    RECT 1353.0000 399.0000 1359.0000 399.3000 ;
	    RECT 1353.0000 393.3000 1354.2001 399.0000 ;
	    RECT 1355.4000 393.3000 1356.6000 398.1000 ;
	    RECT 1357.8000 393.3000 1359.0000 399.0000 ;
	    RECT 1389.0000 393.3000 1390.2001 402.3000 ;
	    RECT 1394.4000 401.7000 1397.1000 402.3000 ;
	    RECT 1394.4000 393.3000 1395.6000 401.7000 ;
	    RECT 1422.6000 401.4000 1423.8000 402.6000 ;
	    RECT 1424.7001 400.8000 1425.0000 402.3000 ;
	    RECT 1427.1000 401.4000 1428.9000 402.6000 ;
	    RECT 1429.8000 402.4500 1431.0000 402.6000 ;
	    RECT 1434.6000 402.4500 1435.8000 402.6000 ;
	    RECT 1429.8000 401.5500 1435.8000 402.4500 ;
	    RECT 1429.8000 401.4000 1431.0000 401.5500 ;
	    RECT 1434.6000 401.4000 1435.8000 401.5500 ;
	    RECT 1439.4000 402.4500 1440.6000 402.6000 ;
	    RECT 1444.2001 402.4500 1445.4000 402.6000 ;
	    RECT 1461.0000 402.4500 1462.2001 402.6000 ;
	    RECT 1439.4000 401.5500 1462.2001 402.4500 ;
	    RECT 1439.4000 401.4000 1440.6000 401.5500 ;
	    RECT 1444.2001 401.4000 1445.4000 401.5500 ;
	    RECT 1461.0000 401.4000 1462.2001 401.5500 ;
	    RECT 1422.9000 399.3000 1428.3000 399.9000 ;
	    RECT 1429.8000 399.3000 1430.7001 400.5000 ;
	    RECT 1422.6000 399.0000 1428.6000 399.3000 ;
	    RECT 1422.6000 393.3000 1423.8000 399.0000 ;
	    RECT 1425.0000 393.3000 1426.2001 398.1000 ;
	    RECT 1427.4000 393.3000 1428.6000 399.0000 ;
	    RECT 1429.8000 393.3000 1431.0000 399.3000 ;
	    RECT 1444.2001 393.3000 1445.4000 400.5000 ;
	    RECT 1446.6000 398.4000 1447.8000 399.6000 ;
	    RECT 1468.2001 399.3000 1469.4000 403.5000 ;
	    RECT 1511.7001 402.6000 1512.6000 406.5000 ;
	    RECT 1518.6000 406.2000 1519.8000 406.5000 ;
	    RECT 1515.0000 404.4000 1515.3000 405.6000 ;
	    RECT 1516.2001 404.4000 1517.4000 405.6000 ;
	    RECT 1540.2001 405.4500 1541.4000 405.6000 ;
	    RECT 1542.6000 405.4500 1543.8000 405.6000 ;
	    RECT 1540.2001 404.5500 1543.8000 405.4500 ;
	    RECT 1544.7001 404.7000 1546.2001 405.6000 ;
	    RECT 1548.6000 404.7000 1548.9000 406.2000 ;
	    RECT 1540.2001 404.4000 1541.4000 404.5500 ;
	    RECT 1542.6000 404.4000 1543.8000 404.5500 ;
	    RECT 1470.6000 401.4000 1471.8000 402.6000 ;
	    RECT 1485.0000 402.4500 1486.2001 402.6000 ;
	    RECT 1504.2001 402.4500 1505.4000 402.6000 ;
	    RECT 1485.0000 401.5500 1505.4000 402.4500 ;
	    RECT 1511.7001 402.3000 1514.1000 402.6000 ;
	    RECT 1511.7001 401.7000 1514.4000 402.3000 ;
	    RECT 1485.0000 401.4000 1486.2001 401.5500 ;
	    RECT 1504.2001 401.4000 1505.4000 401.5500 ;
	    RECT 1470.6000 400.2000 1471.8000 400.5000 ;
	    RECT 1466.7001 398.4000 1469.4000 399.3000 ;
	    RECT 1446.6000 397.2000 1447.8000 397.5000 ;
	    RECT 1446.6000 393.3000 1447.8000 396.3000 ;
	    RECT 1466.7001 393.3000 1467.9000 398.4000 ;
	    RECT 1470.6000 393.3000 1471.8000 399.3000 ;
	    RECT 1485.0000 393.3000 1486.2001 400.5000 ;
	    RECT 1487.4000 398.4000 1488.6000 399.6000 ;
	    RECT 1487.4000 397.2000 1488.6000 397.5000 ;
	    RECT 1487.4000 393.3000 1488.6000 396.3000 ;
	    RECT 1513.2001 393.3000 1514.4000 401.7000 ;
	    RECT 1518.6000 393.3000 1519.8000 402.3000 ;
	    RECT 1523.4000 399.4500 1524.6000 399.6000 ;
	    RECT 1542.6000 399.4500 1543.8000 399.6000 ;
	    RECT 1523.4000 398.5500 1543.8000 399.4500 ;
	    RECT 1545.3000 399.3000 1546.2001 404.7000 ;
	    RECT 1549.8000 404.4000 1551.0000 405.6000 ;
	    RECT 1547.4000 403.5000 1548.6000 403.8000 ;
	    RECT 1547.4000 402.4500 1548.6000 402.6000 ;
	    RECT 1552.2001 402.4500 1553.4000 402.6000 ;
	    RECT 1547.4000 401.5500 1553.4000 402.4500 ;
	    RECT 1547.4000 401.4000 1548.6000 401.5500 ;
	    RECT 1552.2001 401.4000 1553.4000 401.5500 ;
	    RECT 1523.4000 398.4000 1524.6000 398.5500 ;
	    RECT 1542.6000 398.4000 1543.8000 398.5500 ;
	    RECT 1542.9000 397.2000 1544.1000 397.5000 ;
	    RECT 1542.6000 393.3000 1543.8000 396.3000 ;
	    RECT 1545.0000 393.3000 1546.2001 399.3000 ;
	    RECT 1548.9000 393.3000 1550.1000 399.3000 ;
	    RECT 1.2000 390.6000 1569.0000 392.4000 ;
	    RECT 124.2000 380.7000 125.4000 389.7000 ;
	    RECT 129.0000 383.7000 130.2000 389.7000 ;
	    RECT 133.8000 384.9000 135.0000 389.7000 ;
	    RECT 136.2000 385.5000 137.4000 389.7000 ;
	    RECT 138.6000 385.5000 139.8000 389.7000 ;
	    RECT 141.0000 385.5000 142.2000 389.7000 ;
	    RECT 143.4000 386.7000 144.6000 389.7000 ;
	    RECT 145.8000 385.5000 147.0000 389.7000 ;
	    RECT 148.2000 386.7000 149.4000 389.7000 ;
	    RECT 150.6000 385.5000 151.8000 389.7000 ;
	    RECT 153.0000 385.5000 154.2000 389.7000 ;
	    RECT 155.4000 385.5000 156.6000 389.7000 ;
	    RECT 157.8000 385.5000 159.0000 389.7000 ;
	    RECT 131.1000 383.7000 135.0000 384.9000 ;
	    RECT 160.2000 384.9000 161.4000 389.7000 ;
	    RECT 140.1000 383.7000 147.0000 384.6000 ;
	    RECT 131.1000 382.8000 132.3000 383.7000 ;
	    RECT 127.8000 381.6000 132.3000 382.8000 ;
	    RECT 124.2000 379.5000 137.4000 380.7000 ;
	    RECT 140.1000 380.1000 141.3000 383.7000 ;
	    RECT 145.8000 383.4000 147.0000 383.7000 ;
	    RECT 148.2000 383.4000 149.4000 384.6000 ;
	    RECT 150.3000 383.4000 150.6000 384.6000 ;
	    RECT 155.1000 383.4000 156.6000 384.6000 ;
	    RECT 160.2000 383.7000 163.8000 384.9000 ;
	    RECT 165.0000 383.7000 166.2000 389.7000 ;
	    RECT 143.4000 382.5000 144.6000 382.8000 ;
	    RECT 145.8000 382.2000 147.0000 382.5000 ;
	    RECT 143.4000 380.4000 144.6000 381.6000 ;
	    RECT 145.8000 381.3000 152.4000 382.2000 ;
	    RECT 151.2000 381.0000 152.4000 381.3000 ;
	    RECT 124.2000 371.1000 125.4000 379.5000 ;
	    RECT 138.3000 378.9000 141.3000 380.1000 ;
	    RECT 147.0000 378.9000 151.8000 380.1000 ;
	    RECT 155.4000 379.2000 156.6000 383.4000 ;
	    RECT 162.6000 382.8000 163.8000 383.7000 ;
	    RECT 162.6000 381.9000 165.3000 382.8000 ;
	    RECT 164.1000 380.1000 165.3000 381.9000 ;
	    RECT 169.8000 381.9000 171.0000 389.7000 ;
	    RECT 172.2000 384.0000 173.4000 389.7000 ;
	    RECT 174.6000 386.7000 175.8000 389.7000 ;
	    RECT 172.2000 382.8000 173.7000 384.0000 ;
	    RECT 193.8000 383.7000 195.0000 389.7000 ;
	    RECT 197.7000 384.6000 198.9000 389.7000 ;
	    RECT 220.2000 386.7000 221.4000 389.7000 ;
	    RECT 220.2000 385.5000 221.4000 385.8000 ;
	    RECT 196.2000 383.7000 198.9000 384.6000 ;
	    RECT 169.8000 381.0000 171.6000 381.9000 ;
	    RECT 164.1000 378.9000 169.8000 380.1000 ;
	    RECT 126.3000 378.0000 127.5000 378.3000 ;
	    RECT 126.3000 377.1000 132.9000 378.0000 ;
	    RECT 133.8000 377.4000 135.0000 378.6000 ;
	    RECT 160.2000 378.0000 161.4000 378.9000 ;
	    RECT 170.7000 378.0000 171.6000 381.0000 ;
	    RECT 135.9000 377.1000 161.4000 378.0000 ;
	    RECT 170.4000 377.1000 171.6000 378.0000 ;
	    RECT 168.3000 376.2000 169.5000 376.5000 ;
	    RECT 129.0000 374.4000 130.2000 375.6000 ;
	    RECT 131.1000 375.3000 169.5000 376.2000 ;
	    RECT 134.1000 375.0000 135.3000 375.3000 ;
	    RECT 170.4000 374.4000 171.3000 377.1000 ;
	    RECT 172.5000 376.2000 173.7000 382.8000 ;
	    RECT 193.8000 382.5000 195.0000 382.8000 ;
	    RECT 186.6000 381.4500 187.8000 381.6000 ;
	    RECT 193.8000 381.4500 195.0000 381.6000 ;
	    RECT 186.6000 380.5500 195.0000 381.4500 ;
	    RECT 186.6000 380.4000 187.8000 380.5500 ;
	    RECT 193.8000 380.4000 195.0000 380.5500 ;
	    RECT 196.2000 379.5000 197.4000 383.7000 ;
	    RECT 220.2000 383.4000 221.4000 384.6000 ;
	    RECT 222.6000 382.5000 223.8000 389.7000 ;
	    RECT 246.6000 384.0000 247.8000 389.7000 ;
	    RECT 249.0000 384.9000 250.2000 389.7000 ;
	    RECT 251.4000 384.0000 252.6000 389.7000 ;
	    RECT 246.6000 383.7000 252.6000 384.0000 ;
	    RECT 253.8000 383.7000 255.0000 389.7000 ;
	    RECT 273.0000 383.7000 274.2000 389.7000 ;
	    RECT 276.9000 384.6000 278.1000 389.7000 ;
	    RECT 275.4000 383.7000 278.1000 384.6000 ;
	    RECT 297.9000 384.6000 299.1000 389.7000 ;
	    RECT 297.9000 383.7000 300.6000 384.6000 ;
	    RECT 301.8000 383.7000 303.0000 389.7000 ;
	    RECT 316.2000 386.7000 317.4000 389.7000 ;
	    RECT 316.2000 385.5000 317.4000 385.8000 ;
	    RECT 246.9000 383.1000 252.3000 383.7000 ;
	    RECT 253.8000 382.5000 254.7000 383.7000 ;
	    RECT 273.0000 382.5000 274.2000 382.8000 ;
	    RECT 222.6000 381.4500 223.8000 381.6000 ;
	    RECT 222.6000 380.5500 245.2500 381.4500 ;
	    RECT 222.6000 380.4000 223.8000 380.5500 ;
	    RECT 174.6000 378.4500 175.8000 378.6000 ;
	    RECT 196.2000 378.4500 197.4000 378.6000 ;
	    RECT 174.6000 377.5500 197.4000 378.4500 ;
	    RECT 174.6000 377.4000 175.8000 377.5500 ;
	    RECT 196.2000 377.4000 197.4000 377.5500 ;
	    RECT 138.6000 374.1000 139.8000 374.4000 ;
	    RECT 131.7000 373.5000 139.8000 374.1000 ;
	    RECT 130.5000 373.2000 139.8000 373.5000 ;
	    RECT 141.3000 373.5000 154.2000 374.4000 ;
	    RECT 126.6000 372.0000 129.0000 373.2000 ;
	    RECT 130.5000 372.3000 132.6000 373.2000 ;
	    RECT 141.3000 372.3000 142.2000 373.5000 ;
	    RECT 153.0000 373.2000 154.2000 373.5000 ;
	    RECT 157.8000 373.5000 171.3000 374.4000 ;
	    RECT 172.2000 375.0000 173.7000 376.2000 ;
	    RECT 172.2000 373.5000 173.4000 375.0000 ;
	    RECT 157.8000 373.2000 159.0000 373.5000 ;
	    RECT 128.1000 371.4000 129.0000 372.0000 ;
	    RECT 133.5000 371.4000 142.2000 372.3000 ;
	    RECT 143.1000 371.4000 147.0000 372.6000 ;
	    RECT 124.2000 370.2000 127.2000 371.1000 ;
	    RECT 128.1000 370.2000 134.4000 371.4000 ;
	    RECT 126.3000 369.3000 127.2000 370.2000 ;
	    RECT 124.2000 363.3000 125.4000 369.3000 ;
	    RECT 126.3000 368.4000 127.8000 369.3000 ;
	    RECT 126.6000 363.3000 127.8000 368.4000 ;
	    RECT 129.0000 362.4000 130.2000 369.3000 ;
	    RECT 131.4000 363.3000 132.6000 370.2000 ;
	    RECT 133.8000 363.3000 135.0000 369.3000 ;
	    RECT 136.2000 363.3000 137.4000 367.5000 ;
	    RECT 138.6000 363.3000 139.8000 367.5000 ;
	    RECT 141.0000 363.3000 142.2000 370.5000 ;
	    RECT 143.4000 363.3000 144.6000 369.3000 ;
	    RECT 145.8000 363.3000 147.0000 370.5000 ;
	    RECT 148.2000 363.3000 149.4000 369.3000 ;
	    RECT 150.6000 363.3000 151.8000 372.6000 ;
	    RECT 162.6000 371.4000 166.5000 372.6000 ;
	    RECT 155.4000 370.2000 161.7000 371.4000 ;
	    RECT 153.0000 363.3000 154.2000 367.5000 ;
	    RECT 155.4000 363.3000 156.6000 367.5000 ;
	    RECT 157.8000 363.3000 159.0000 367.5000 ;
	    RECT 160.2000 363.3000 161.4000 369.3000 ;
	    RECT 162.6000 363.3000 163.8000 371.4000 ;
	    RECT 170.4000 371.1000 171.3000 373.5000 ;
	    RECT 172.2000 371.4000 173.4000 372.6000 ;
	    RECT 167.4000 370.2000 171.3000 371.1000 ;
	    RECT 165.0000 363.3000 166.2000 369.3000 ;
	    RECT 167.4000 363.3000 168.6000 370.2000 ;
	    RECT 169.8000 363.3000 171.0000 369.3000 ;
	    RECT 172.2000 363.3000 173.4000 370.5000 ;
	    RECT 174.6000 363.3000 175.8000 369.3000 ;
	    RECT 193.8000 363.3000 195.0000 369.3000 ;
	    RECT 196.2000 363.3000 197.4000 376.5000 ;
	    RECT 198.6000 374.4000 199.8000 375.6000 ;
	    RECT 198.6000 373.2000 199.8000 373.5000 ;
	    RECT 198.6000 363.3000 199.8000 369.3000 ;
	    RECT 220.2000 363.3000 221.4000 369.3000 ;
	    RECT 222.6000 363.3000 223.8000 379.5000 ;
	    RECT 244.3500 378.4500 245.2500 380.5500 ;
	    RECT 246.6000 380.4000 247.8000 381.6000 ;
	    RECT 248.7000 380.7000 249.0000 382.2000 ;
	    RECT 251.1000 380.4000 252.9000 381.6000 ;
	    RECT 253.8000 381.4500 255.0000 381.6000 ;
	    RECT 270.6000 381.4500 271.8000 381.6000 ;
	    RECT 253.8000 380.5500 271.8000 381.4500 ;
	    RECT 253.8000 380.4000 255.0000 380.5500 ;
	    RECT 270.6000 380.4000 271.8000 380.5500 ;
	    RECT 273.0000 380.4000 274.2000 381.6000 ;
	    RECT 249.0000 379.5000 250.2000 379.8000 ;
	    RECT 249.0000 378.4500 250.2000 378.6000 ;
	    RECT 244.3500 377.5500 250.2000 378.4500 ;
	    RECT 249.0000 377.4000 250.2000 377.5500 ;
	    RECT 251.1000 375.3000 252.0000 380.4000 ;
	    RECT 275.4000 379.5000 276.6000 383.7000 ;
	    RECT 299.4000 379.5000 300.6000 383.7000 ;
	    RECT 316.2000 383.4000 317.4000 384.6000 ;
	    RECT 301.8000 382.5000 303.0000 382.8000 ;
	    RECT 318.6000 382.5000 319.8000 389.7000 ;
	    RECT 342.6000 384.0000 343.8000 389.7000 ;
	    RECT 345.0000 384.9000 346.2000 389.7000 ;
	    RECT 347.4000 384.0000 348.6000 389.7000 ;
	    RECT 342.6000 383.7000 348.6000 384.0000 ;
	    RECT 349.8000 383.7000 351.0000 389.7000 ;
	    RECT 481.8000 386.7000 483.0000 389.7000 ;
	    RECT 484.2000 384.0000 485.4000 389.7000 ;
	    RECT 342.9000 383.1000 348.3000 383.7000 ;
	    RECT 349.8000 382.5000 350.7000 383.7000 ;
	    RECT 483.9000 382.8000 485.4000 384.0000 ;
	    RECT 301.8000 380.4000 303.0000 381.6000 ;
	    RECT 318.6000 381.4500 319.8000 381.6000 ;
	    RECT 318.6000 380.5500 341.2500 381.4500 ;
	    RECT 318.6000 380.4000 319.8000 380.5500 ;
	    RECT 275.4000 378.4500 276.6000 378.6000 ;
	    RECT 253.9500 377.5500 276.6000 378.4500 ;
	    RECT 253.9500 375.6000 254.8500 377.5500 ;
	    RECT 275.4000 377.4000 276.6000 377.5500 ;
	    RECT 299.4000 378.4500 300.6000 378.6000 ;
	    RECT 316.2000 378.4500 317.4000 378.6000 ;
	    RECT 299.4000 377.5500 317.4000 378.4500 ;
	    RECT 299.4000 377.4000 300.6000 377.5500 ;
	    RECT 316.2000 377.4000 317.4000 377.5500 ;
	    RECT 246.6000 363.3000 247.8000 375.3000 ;
	    RECT 250.5000 374.4000 252.0000 375.3000 ;
	    RECT 253.8000 374.4000 255.0000 375.6000 ;
	    RECT 250.5000 363.3000 251.7000 374.4000 ;
	    RECT 252.9000 372.6000 253.8000 373.5000 ;
	    RECT 252.6000 371.4000 253.8000 372.6000 ;
	    RECT 252.9000 363.3000 254.1000 369.3000 ;
	    RECT 273.0000 363.3000 274.2000 369.3000 ;
	    RECT 275.4000 363.3000 276.6000 376.5000 ;
	    RECT 277.8000 375.4500 279.0000 375.6000 ;
	    RECT 287.4000 375.4500 288.6000 375.6000 ;
	    RECT 297.0000 375.4500 298.2000 375.6000 ;
	    RECT 277.8000 374.5500 281.2500 375.4500 ;
	    RECT 277.8000 374.4000 279.0000 374.5500 ;
	    RECT 277.8000 373.2000 279.0000 373.5000 ;
	    RECT 280.3500 372.4500 281.2500 374.5500 ;
	    RECT 287.4000 374.5500 298.2000 375.4500 ;
	    RECT 287.4000 374.4000 288.6000 374.5500 ;
	    RECT 297.0000 374.4000 298.2000 374.5500 ;
	    RECT 297.0000 373.2000 298.2000 373.5000 ;
	    RECT 294.6000 372.4500 295.8000 372.6000 ;
	    RECT 280.3500 371.5500 295.8000 372.4500 ;
	    RECT 294.6000 371.4000 295.8000 371.5500 ;
	    RECT 277.8000 363.3000 279.0000 369.3000 ;
	    RECT 297.0000 363.3000 298.2000 369.3000 ;
	    RECT 299.4000 363.3000 300.6000 376.5000 ;
	    RECT 301.8000 363.3000 303.0000 369.3000 ;
	    RECT 316.2000 363.3000 317.4000 369.3000 ;
	    RECT 318.6000 363.3000 319.8000 379.5000 ;
	    RECT 340.3500 378.4500 341.2500 380.5500 ;
	    RECT 342.6000 380.4000 343.8000 381.6000 ;
	    RECT 344.7000 380.7000 345.0000 382.2000 ;
	    RECT 347.1000 380.4000 348.9000 381.6000 ;
	    RECT 349.8000 381.4500 351.0000 381.6000 ;
	    RECT 402.6000 381.4500 403.8000 381.6000 ;
	    RECT 349.8000 380.5500 403.8000 381.4500 ;
	    RECT 349.8000 380.4000 351.0000 380.5500 ;
	    RECT 402.6000 380.4000 403.8000 380.5500 ;
	    RECT 345.0000 379.5000 346.2000 379.8000 ;
	    RECT 345.0000 378.4500 346.2000 378.6000 ;
	    RECT 340.3500 377.5500 346.2000 378.4500 ;
	    RECT 345.0000 377.4000 346.2000 377.5500 ;
	    RECT 347.1000 375.3000 348.0000 380.4000 ;
	    RECT 483.9000 376.2000 485.1000 382.8000 ;
	    RECT 486.6000 381.9000 487.8000 389.7000 ;
	    RECT 491.4000 383.7000 492.6000 389.7000 ;
	    RECT 496.2000 384.9000 497.4000 389.7000 ;
	    RECT 498.6000 385.5000 499.8000 389.7000 ;
	    RECT 501.0000 385.5000 502.2000 389.7000 ;
	    RECT 503.4000 385.5000 504.6000 389.7000 ;
	    RECT 505.8000 385.5000 507.0000 389.7000 ;
	    RECT 508.2000 386.7000 509.4000 389.7000 ;
	    RECT 510.6000 385.5000 511.8000 389.7000 ;
	    RECT 513.0000 386.7000 514.2000 389.7000 ;
	    RECT 515.4000 385.5000 516.6000 389.7000 ;
	    RECT 517.8000 385.5000 519.0000 389.7000 ;
	    RECT 520.2000 385.5000 521.4000 389.7000 ;
	    RECT 493.8000 383.7000 497.4000 384.9000 ;
	    RECT 522.6000 384.9000 523.8000 389.7000 ;
	    RECT 493.8000 382.8000 495.0000 383.7000 ;
	    RECT 486.0000 381.0000 487.8000 381.9000 ;
	    RECT 492.3000 381.9000 495.0000 382.8000 ;
	    RECT 501.0000 383.4000 502.5000 384.6000 ;
	    RECT 507.0000 383.4000 507.3000 384.6000 ;
	    RECT 508.2000 383.4000 509.4000 384.6000 ;
	    RECT 510.6000 383.7000 517.5000 384.6000 ;
	    RECT 522.6000 383.7000 526.5000 384.9000 ;
	    RECT 527.4000 383.7000 528.6000 389.7000 ;
	    RECT 510.6000 383.4000 511.8000 383.7000 ;
	    RECT 486.0000 378.0000 486.9000 381.0000 ;
	    RECT 492.3000 380.1000 493.5000 381.9000 ;
	    RECT 487.8000 378.9000 493.5000 380.1000 ;
	    RECT 501.0000 379.2000 502.2000 383.4000 ;
	    RECT 513.0000 382.5000 514.2000 382.8000 ;
	    RECT 510.6000 382.2000 511.8000 382.5000 ;
	    RECT 505.2000 381.3000 511.8000 382.2000 ;
	    RECT 505.2000 381.0000 506.4000 381.3000 ;
	    RECT 513.0000 380.4000 514.2000 381.6000 ;
	    RECT 516.3000 380.1000 517.5000 383.7000 ;
	    RECT 525.3000 382.8000 526.5000 383.7000 ;
	    RECT 525.3000 381.6000 529.8000 382.8000 ;
	    RECT 532.2000 380.7000 533.4000 389.7000 ;
	    RECT 552.3000 384.6000 553.5000 389.7000 ;
	    RECT 552.3000 383.7000 555.0000 384.6000 ;
	    RECT 556.2000 383.7000 557.4000 389.7000 ;
	    RECT 580.2000 383.7000 581.4000 389.7000 ;
	    RECT 582.6000 384.0000 583.8000 389.7000 ;
	    RECT 585.0000 384.9000 586.2000 389.7000 ;
	    RECT 587.4000 384.0000 588.6000 389.7000 ;
	    RECT 606.6000 386.7000 607.8000 389.7000 ;
	    RECT 609.0000 386.7000 610.2000 389.7000 ;
	    RECT 611.4000 386.7000 612.6000 389.7000 ;
	    RECT 623.4000 386.7000 624.6000 389.7000 ;
	    RECT 582.6000 383.7000 588.6000 384.0000 ;
	    RECT 505.8000 378.9000 510.6000 380.1000 ;
	    RECT 516.3000 378.9000 519.3000 380.1000 ;
	    RECT 520.2000 379.5000 533.4000 380.7000 ;
	    RECT 553.8000 379.5000 555.0000 383.7000 ;
	    RECT 556.2000 382.5000 557.4000 382.8000 ;
	    RECT 580.5000 382.5000 581.4000 383.7000 ;
	    RECT 582.9000 383.1000 588.3000 383.7000 ;
	    RECT 609.0000 382.5000 609.9000 386.7000 ;
	    RECT 611.4000 385.5000 612.6000 385.8000 ;
	    RECT 623.4000 385.5000 624.6000 385.8000 ;
	    RECT 611.4000 384.4500 612.6000 384.6000 ;
	    RECT 616.2000 384.4500 617.4000 384.6000 ;
	    RECT 611.4000 383.5500 617.4000 384.4500 ;
	    RECT 611.4000 383.4000 612.6000 383.5500 ;
	    RECT 616.2000 383.4000 617.4000 383.5500 ;
	    RECT 621.0000 384.4500 622.2000 384.6000 ;
	    RECT 623.4000 384.4500 624.6000 384.6000 ;
	    RECT 621.0000 383.5500 624.6000 384.4500 ;
	    RECT 621.0000 383.4000 622.2000 383.5500 ;
	    RECT 623.4000 383.4000 624.6000 383.5500 ;
	    RECT 625.8000 382.5000 627.0000 389.7000 ;
	    RECT 652.2000 384.0000 653.4000 389.7000 ;
	    RECT 654.6000 384.9000 655.8000 389.7000 ;
	    RECT 657.0000 384.0000 658.2000 389.7000 ;
	    RECT 652.2000 383.7000 658.2000 384.0000 ;
	    RECT 659.4000 383.7000 660.6000 389.7000 ;
	    RECT 681.0000 386.7000 682.2000 389.7000 ;
	    RECT 681.0000 385.5000 682.2000 385.8000 ;
	    RECT 671.4000 384.4500 672.6000 384.6000 ;
	    RECT 681.0000 384.4500 682.2000 384.6000 ;
	    RECT 652.5000 383.1000 657.9000 383.7000 ;
	    RECT 659.4000 382.5000 660.3000 383.7000 ;
	    RECT 671.4000 383.5500 682.2000 384.4500 ;
	    RECT 671.4000 383.4000 672.6000 383.5500 ;
	    RECT 681.0000 383.4000 682.2000 383.5500 ;
	    RECT 683.4000 382.5000 684.6000 389.7000 ;
	    RECT 738.6000 389.4000 739.8000 390.6000 ;
	    RECT 700.2000 387.4500 701.4000 387.6000 ;
	    RECT 798.6000 387.4500 799.8000 387.6000 ;
	    RECT 700.2000 386.5500 799.8000 387.4500 ;
	    RECT 808.2000 386.7000 809.4000 389.7000 ;
	    RECT 700.2000 386.4000 701.4000 386.5500 ;
	    RECT 798.6000 386.4000 799.8000 386.5500 ;
	    RECT 810.6000 384.0000 811.8000 389.7000 ;
	    RECT 810.3000 382.8000 811.8000 384.0000 ;
	    RECT 556.2000 381.4500 557.4000 381.6000 ;
	    RECT 563.4000 381.4500 564.6000 381.6000 ;
	    RECT 556.2000 380.5500 564.6000 381.4500 ;
	    RECT 556.2000 380.4000 557.4000 380.5500 ;
	    RECT 563.4000 380.4000 564.6000 380.5500 ;
	    RECT 580.2000 380.4000 581.4000 381.6000 ;
	    RECT 582.3000 380.4000 584.1000 381.6000 ;
	    RECT 586.2000 380.7000 586.5000 382.2000 ;
	    RECT 587.4000 381.4500 588.6000 381.6000 ;
	    RECT 599.4000 381.4500 600.6000 381.6000 ;
	    RECT 587.4000 380.5500 600.6000 381.4500 ;
	    RECT 587.4000 380.4000 588.6000 380.5500 ;
	    RECT 599.4000 380.4000 600.6000 380.5500 ;
	    RECT 609.0000 380.4000 610.2000 381.6000 ;
	    RECT 625.8000 381.4500 627.0000 381.6000 ;
	    RECT 647.4000 381.4500 648.6000 381.6000 ;
	    RECT 652.2000 381.4500 653.4000 381.6000 ;
	    RECT 625.8000 380.5500 646.0500 381.4500 ;
	    RECT 625.8000 380.4000 627.0000 380.5500 ;
	    RECT 496.2000 378.0000 497.4000 378.9000 ;
	    RECT 486.0000 377.1000 487.2000 378.0000 ;
	    RECT 496.2000 377.1000 521.7000 378.0000 ;
	    RECT 522.6000 377.4000 523.8000 378.6000 ;
	    RECT 530.1000 378.0000 531.3000 378.3000 ;
	    RECT 524.7000 377.1000 531.3000 378.0000 ;
	    RECT 342.6000 363.3000 343.8000 375.3000 ;
	    RECT 346.5000 374.4000 348.0000 375.3000 ;
	    RECT 349.8000 374.4000 351.0000 375.6000 ;
	    RECT 483.9000 375.0000 485.4000 376.2000 ;
	    RECT 346.5000 363.3000 347.7000 374.4000 ;
	    RECT 484.2000 373.5000 485.4000 375.0000 ;
	    RECT 486.3000 374.4000 487.2000 377.1000 ;
	    RECT 488.1000 376.2000 489.3000 376.5000 ;
	    RECT 488.1000 375.3000 526.5000 376.2000 ;
	    RECT 522.3000 375.0000 523.5000 375.3000 ;
	    RECT 527.4000 374.4000 528.6000 375.6000 ;
	    RECT 486.3000 373.5000 499.8000 374.4000 ;
	    RECT 348.9000 372.6000 349.8000 373.5000 ;
	    RECT 348.6000 371.4000 349.8000 372.6000 ;
	    RECT 352.2000 372.4500 353.4000 372.6000 ;
	    RECT 484.2000 372.4500 485.4000 372.6000 ;
	    RECT 352.2000 371.5500 485.4000 372.4500 ;
	    RECT 352.2000 371.4000 353.4000 371.5500 ;
	    RECT 484.2000 371.4000 485.4000 371.5500 ;
	    RECT 486.3000 371.1000 487.2000 373.5000 ;
	    RECT 498.6000 373.2000 499.8000 373.5000 ;
	    RECT 503.4000 373.5000 516.3000 374.4000 ;
	    RECT 503.4000 373.2000 504.6000 373.5000 ;
	    RECT 491.1000 371.4000 495.0000 372.6000 ;
	    RECT 348.9000 363.3000 350.1000 369.3000 ;
	    RECT 481.8000 363.3000 483.0000 369.3000 ;
	    RECT 484.2000 363.3000 485.4000 370.5000 ;
	    RECT 486.3000 370.2000 490.2000 371.1000 ;
	    RECT 486.6000 363.3000 487.8000 369.3000 ;
	    RECT 489.0000 363.3000 490.2000 370.2000 ;
	    RECT 491.4000 363.3000 492.6000 369.3000 ;
	    RECT 493.8000 363.3000 495.0000 371.4000 ;
	    RECT 495.9000 370.2000 502.2000 371.4000 ;
	    RECT 496.2000 363.3000 497.4000 369.3000 ;
	    RECT 498.6000 363.3000 499.8000 367.5000 ;
	    RECT 501.0000 363.3000 502.2000 367.5000 ;
	    RECT 503.4000 363.3000 504.6000 367.5000 ;
	    RECT 505.8000 363.3000 507.0000 372.6000 ;
	    RECT 510.6000 371.4000 514.5000 372.6000 ;
	    RECT 515.4000 372.3000 516.3000 373.5000 ;
	    RECT 517.8000 374.1000 519.0000 374.4000 ;
	    RECT 517.8000 373.5000 525.9000 374.1000 ;
	    RECT 517.8000 373.2000 527.1000 373.5000 ;
	    RECT 525.0000 372.3000 527.1000 373.2000 ;
	    RECT 515.4000 371.4000 524.1000 372.3000 ;
	    RECT 528.6000 372.0000 531.0000 373.2000 ;
	    RECT 528.6000 371.4000 529.5000 372.0000 ;
	    RECT 508.2000 363.3000 509.4000 369.3000 ;
	    RECT 510.6000 363.3000 511.8000 370.5000 ;
	    RECT 513.0000 363.3000 514.2000 369.3000 ;
	    RECT 515.4000 363.3000 516.6000 370.5000 ;
	    RECT 523.2000 370.2000 529.5000 371.4000 ;
	    RECT 532.2000 371.1000 533.4000 379.5000 ;
	    RECT 534.6000 378.4500 535.8000 378.6000 ;
	    RECT 553.8000 378.4500 555.0000 378.6000 ;
	    RECT 534.6000 377.5500 555.0000 378.4500 ;
	    RECT 534.6000 377.4000 535.8000 377.5500 ;
	    RECT 553.8000 377.4000 555.0000 377.5500 ;
	    RECT 551.4000 374.4000 552.6000 375.6000 ;
	    RECT 551.4000 373.2000 552.6000 373.5000 ;
	    RECT 530.4000 370.2000 533.4000 371.1000 ;
	    RECT 517.8000 363.3000 519.0000 367.5000 ;
	    RECT 520.2000 363.3000 521.4000 367.5000 ;
	    RECT 522.6000 363.3000 523.8000 369.3000 ;
	    RECT 525.0000 363.3000 526.2000 370.2000 ;
	    RECT 530.4000 369.3000 531.3000 370.2000 ;
	    RECT 527.4000 362.4000 528.6000 369.3000 ;
	    RECT 529.8000 368.4000 531.3000 369.3000 ;
	    RECT 529.8000 363.3000 531.0000 368.4000 ;
	    RECT 532.2000 363.3000 533.4000 369.3000 ;
	    RECT 551.4000 363.3000 552.6000 369.3000 ;
	    RECT 553.8000 363.3000 555.0000 376.5000 ;
	    RECT 577.8000 375.4500 579.0000 375.6000 ;
	    RECT 580.2000 375.4500 581.4000 375.6000 ;
	    RECT 577.8000 374.5500 581.4000 375.4500 ;
	    RECT 577.8000 374.4000 579.0000 374.5500 ;
	    RECT 580.2000 374.4000 581.4000 374.5500 ;
	    RECT 583.2000 375.3000 584.1000 380.4000 ;
	    RECT 585.0000 379.5000 586.2000 379.8000 ;
	    RECT 585.0000 377.4000 586.2000 378.6000 ;
	    RECT 606.6000 377.4000 607.8000 378.6000 ;
	    RECT 606.6000 376.2000 607.8000 376.5000 ;
	    RECT 609.0000 375.3000 609.9000 379.5000 ;
	    RECT 583.2000 374.4000 584.7000 375.3000 ;
	    RECT 581.4000 372.6000 582.3000 373.5000 ;
	    RECT 581.4000 371.4000 582.6000 372.6000 ;
	    RECT 556.2000 363.3000 557.4000 369.3000 ;
	    RECT 581.1000 363.3000 582.3000 369.3000 ;
	    RECT 583.5000 363.3000 584.7000 374.4000 ;
	    RECT 587.4000 363.3000 588.6000 375.3000 ;
	    RECT 607.5000 374.1000 610.2000 375.3000 ;
	    RECT 607.5000 363.3000 608.7000 374.1000 ;
	    RECT 611.4000 363.3000 612.6000 375.3000 ;
	    RECT 623.4000 363.3000 624.6000 369.3000 ;
	    RECT 625.8000 363.3000 627.0000 379.5000 ;
	    RECT 645.1500 378.4500 646.0500 380.5500 ;
	    RECT 647.4000 380.5500 653.4000 381.4500 ;
	    RECT 654.3000 380.7000 654.6000 382.2000 ;
	    RECT 647.4000 380.4000 648.6000 380.5500 ;
	    RECT 652.2000 380.4000 653.4000 380.5500 ;
	    RECT 656.7000 380.4000 658.5000 381.6000 ;
	    RECT 659.4000 381.4500 660.6000 381.6000 ;
	    RECT 681.0000 381.4500 682.2000 381.6000 ;
	    RECT 659.4000 380.5500 682.2000 381.4500 ;
	    RECT 659.4000 380.4000 660.6000 380.5500 ;
	    RECT 681.0000 380.4000 682.2000 380.5500 ;
	    RECT 683.4000 381.4500 684.6000 381.6000 ;
	    RECT 685.8000 381.4500 687.0000 381.6000 ;
	    RECT 683.4000 380.5500 687.0000 381.4500 ;
	    RECT 683.4000 380.4000 684.6000 380.5500 ;
	    RECT 685.8000 380.4000 687.0000 380.5500 ;
	    RECT 654.6000 379.5000 655.8000 379.8000 ;
	    RECT 654.6000 378.4500 655.8000 378.6000 ;
	    RECT 645.1500 377.5500 655.8000 378.4500 ;
	    RECT 654.6000 377.4000 655.8000 377.5500 ;
	    RECT 656.7000 375.3000 657.6000 380.4000 ;
	    RECT 652.2000 363.3000 653.4000 375.3000 ;
	    RECT 656.1000 374.4000 657.6000 375.3000 ;
	    RECT 659.4000 374.4000 660.6000 375.6000 ;
	    RECT 656.1000 363.3000 657.3000 374.4000 ;
	    RECT 658.5000 372.6000 659.4000 373.5000 ;
	    RECT 658.2000 371.4000 659.4000 372.6000 ;
	    RECT 658.5000 363.3000 659.7000 369.3000 ;
	    RECT 681.0000 363.3000 682.2000 369.3000 ;
	    RECT 683.4000 363.3000 684.6000 379.5000 ;
	    RECT 810.3000 376.2000 811.5000 382.8000 ;
	    RECT 813.0000 381.9000 814.2000 389.7000 ;
	    RECT 817.8000 383.7000 819.0000 389.7000 ;
	    RECT 822.6000 384.9000 823.8000 389.7000 ;
	    RECT 825.0000 385.5000 826.2000 389.7000 ;
	    RECT 827.4000 385.5000 828.6000 389.7000 ;
	    RECT 829.8000 385.5000 831.0000 389.7000 ;
	    RECT 832.2000 385.5000 833.4000 389.7000 ;
	    RECT 834.6000 386.7000 835.8000 389.7000 ;
	    RECT 837.0000 385.5000 838.2000 389.7000 ;
	    RECT 839.4000 386.7000 840.6000 389.7000 ;
	    RECT 841.8000 385.5000 843.0000 389.7000 ;
	    RECT 844.2000 385.5000 845.4000 389.7000 ;
	    RECT 846.6000 385.5000 847.8000 389.7000 ;
	    RECT 820.2000 383.7000 823.8000 384.9000 ;
	    RECT 849.0000 384.9000 850.2000 389.7000 ;
	    RECT 820.2000 382.8000 821.4000 383.7000 ;
	    RECT 812.4000 381.0000 814.2000 381.9000 ;
	    RECT 818.7000 381.9000 821.4000 382.8000 ;
	    RECT 827.4000 383.4000 828.9000 384.6000 ;
	    RECT 833.4000 383.4000 833.7000 384.6000 ;
	    RECT 834.6000 383.4000 835.8000 384.6000 ;
	    RECT 837.0000 383.7000 843.9000 384.6000 ;
	    RECT 849.0000 383.7000 852.9000 384.9000 ;
	    RECT 853.8000 383.7000 855.0000 389.7000 ;
	    RECT 837.0000 383.4000 838.2000 383.7000 ;
	    RECT 812.4000 378.0000 813.3000 381.0000 ;
	    RECT 818.7000 380.1000 819.9000 381.9000 ;
	    RECT 814.2000 378.9000 819.9000 380.1000 ;
	    RECT 827.4000 379.2000 828.6000 383.4000 ;
	    RECT 839.4000 382.5000 840.6000 382.8000 ;
	    RECT 837.0000 382.2000 838.2000 382.5000 ;
	    RECT 831.6000 381.3000 838.2000 382.2000 ;
	    RECT 831.6000 381.0000 832.8000 381.3000 ;
	    RECT 839.4000 380.4000 840.6000 381.6000 ;
	    RECT 842.7000 380.1000 843.9000 383.7000 ;
	    RECT 851.7000 382.8000 852.9000 383.7000 ;
	    RECT 851.7000 381.6000 856.2000 382.8000 ;
	    RECT 858.6000 380.7000 859.8000 389.7000 ;
	    RECT 877.8000 383.7000 879.0000 389.7000 ;
	    RECT 881.7000 384.6000 882.9000 389.7000 ;
	    RECT 880.2000 383.7000 882.9000 384.6000 ;
	    RECT 916.2000 383.7000 917.4000 389.7000 ;
	    RECT 918.6000 384.0000 919.8000 389.7000 ;
	    RECT 921.0000 384.9000 922.2000 389.7000 ;
	    RECT 923.4000 384.0000 924.6000 389.7000 ;
	    RECT 918.6000 383.7000 924.6000 384.0000 ;
	    RECT 877.8000 382.5000 879.0000 382.8000 ;
	    RECT 832.2000 378.9000 837.0000 380.1000 ;
	    RECT 842.7000 378.9000 845.7000 380.1000 ;
	    RECT 846.6000 379.5000 859.8000 380.7000 ;
	    RECT 877.8000 380.4000 879.0000 381.6000 ;
	    RECT 880.2000 379.5000 881.4000 383.7000 ;
	    RECT 916.5000 382.5000 917.4000 383.7000 ;
	    RECT 918.9000 383.1000 924.3000 383.7000 ;
	    RECT 935.4000 382.5000 936.6000 389.7000 ;
	    RECT 937.8000 386.7000 939.0000 389.7000 ;
	    RECT 937.8000 385.5000 939.0000 385.8000 ;
	    RECT 937.8000 384.4500 939.0000 384.6000 ;
	    RECT 969.0000 384.4500 970.2000 384.6000 ;
	    RECT 937.8000 383.5500 970.2000 384.4500 ;
	    RECT 990.6000 383.7000 991.8000 389.7000 ;
	    RECT 937.8000 383.4000 939.0000 383.5500 ;
	    RECT 969.0000 383.4000 970.2000 383.5500 ;
	    RECT 993.0000 382.8000 994.2000 389.7000 ;
	    RECT 995.4000 383.7000 996.6000 389.7000 ;
	    RECT 997.8000 382.8000 999.0000 389.7000 ;
	    RECT 1000.2000 383.7000 1001.4000 389.7000 ;
	    RECT 1002.6000 382.8000 1003.8000 389.7000 ;
	    RECT 1005.0000 383.7000 1006.2000 389.7000 ;
	    RECT 1007.4000 382.8000 1008.6000 389.7000 ;
	    RECT 1009.8000 383.7000 1011.0000 389.7000 ;
	    RECT 1012.2000 389.4000 1013.4000 390.6000 ;
	    RECT 1029.9000 384.6000 1031.1000 389.7000 ;
	    RECT 1029.9000 383.7000 1032.6000 384.6000 ;
	    RECT 1033.8000 383.7000 1035.0000 389.7000 ;
	    RECT 1060.2001 383.7000 1061.4000 389.7000 ;
	    RECT 1062.6000 384.0000 1063.8000 389.7000 ;
	    RECT 1065.0000 384.9000 1066.2001 389.7000 ;
	    RECT 1067.4000 384.0000 1068.6000 389.7000 ;
	    RECT 1062.6000 383.7000 1068.6000 384.0000 ;
	    RECT 916.2000 380.4000 917.4000 381.6000 ;
	    RECT 918.3000 380.4000 920.1000 381.6000 ;
	    RECT 922.2000 380.7000 922.5000 382.2000 ;
	    RECT 990.6000 381.6000 994.2000 382.8000 ;
	    RECT 995.7000 381.6000 999.0000 382.8000 ;
	    RECT 1000.5000 381.6000 1003.8000 382.8000 ;
	    RECT 1005.9000 381.6000 1008.6000 382.8000 ;
	    RECT 923.4000 380.4000 924.6000 381.6000 ;
	    RECT 935.4000 381.4500 936.6000 381.6000 ;
	    RECT 925.9500 380.5500 936.6000 381.4500 ;
	    RECT 822.6000 378.0000 823.8000 378.9000 ;
	    RECT 812.4000 377.1000 813.6000 378.0000 ;
	    RECT 822.6000 377.1000 848.1000 378.0000 ;
	    RECT 849.0000 377.4000 850.2000 378.6000 ;
	    RECT 856.5000 378.0000 857.7000 378.3000 ;
	    RECT 851.1000 377.1000 857.7000 378.0000 ;
	    RECT 810.3000 375.0000 811.8000 376.2000 ;
	    RECT 810.6000 373.5000 811.8000 375.0000 ;
	    RECT 812.7000 374.4000 813.6000 377.1000 ;
	    RECT 814.5000 376.2000 815.7000 376.5000 ;
	    RECT 814.5000 375.3000 852.9000 376.2000 ;
	    RECT 848.7000 375.0000 849.9000 375.3000 ;
	    RECT 853.8000 374.4000 855.0000 375.6000 ;
	    RECT 812.7000 373.5000 826.2000 374.4000 ;
	    RECT 750.6000 372.4500 751.8000 372.6000 ;
	    RECT 810.6000 372.4500 811.8000 372.6000 ;
	    RECT 750.6000 371.5500 811.8000 372.4500 ;
	    RECT 750.6000 371.4000 751.8000 371.5500 ;
	    RECT 810.6000 371.4000 811.8000 371.5500 ;
	    RECT 812.7000 371.1000 813.6000 373.5000 ;
	    RECT 825.0000 373.2000 826.2000 373.5000 ;
	    RECT 829.8000 373.5000 842.7000 374.4000 ;
	    RECT 829.8000 373.2000 831.0000 373.5000 ;
	    RECT 817.5000 371.4000 821.4000 372.6000 ;
	    RECT 808.2000 363.3000 809.4000 369.3000 ;
	    RECT 810.6000 363.3000 811.8000 370.5000 ;
	    RECT 812.7000 370.2000 816.6000 371.1000 ;
	    RECT 813.0000 363.3000 814.2000 369.3000 ;
	    RECT 815.4000 363.3000 816.6000 370.2000 ;
	    RECT 817.8000 363.3000 819.0000 369.3000 ;
	    RECT 820.2000 363.3000 821.4000 371.4000 ;
	    RECT 822.3000 370.2000 828.6000 371.4000 ;
	    RECT 822.6000 363.3000 823.8000 369.3000 ;
	    RECT 825.0000 363.3000 826.2000 367.5000 ;
	    RECT 827.4000 363.3000 828.6000 367.5000 ;
	    RECT 829.8000 363.3000 831.0000 367.5000 ;
	    RECT 832.2000 363.3000 833.4000 372.6000 ;
	    RECT 837.0000 371.4000 840.9000 372.6000 ;
	    RECT 841.8000 372.3000 842.7000 373.5000 ;
	    RECT 844.2000 374.1000 845.4000 374.4000 ;
	    RECT 844.2000 373.5000 852.3000 374.1000 ;
	    RECT 844.2000 373.2000 853.5000 373.5000 ;
	    RECT 851.4000 372.3000 853.5000 373.2000 ;
	    RECT 841.8000 371.4000 850.5000 372.3000 ;
	    RECT 855.0000 372.0000 857.4000 373.2000 ;
	    RECT 855.0000 371.4000 855.9000 372.0000 ;
	    RECT 834.6000 363.3000 835.8000 369.3000 ;
	    RECT 837.0000 363.3000 838.2000 370.5000 ;
	    RECT 839.4000 363.3000 840.6000 369.3000 ;
	    RECT 841.8000 363.3000 843.0000 370.5000 ;
	    RECT 849.6000 370.2000 855.9000 371.4000 ;
	    RECT 858.6000 371.1000 859.8000 379.5000 ;
	    RECT 880.2000 378.4500 881.4000 378.6000 ;
	    RECT 880.2000 377.5500 917.2500 378.4500 ;
	    RECT 880.2000 377.4000 881.4000 377.5500 ;
	    RECT 856.8000 370.2000 859.8000 371.1000 ;
	    RECT 844.2000 363.3000 845.4000 367.5000 ;
	    RECT 846.6000 363.3000 847.8000 367.5000 ;
	    RECT 849.0000 363.3000 850.2000 369.3000 ;
	    RECT 851.4000 363.3000 852.6000 370.2000 ;
	    RECT 856.8000 369.3000 857.7000 370.2000 ;
	    RECT 853.8000 362.4000 855.0000 369.3000 ;
	    RECT 856.2000 368.4000 857.7000 369.3000 ;
	    RECT 856.2000 363.3000 857.4000 368.4000 ;
	    RECT 858.6000 363.3000 859.8000 369.3000 ;
	    RECT 877.8000 363.3000 879.0000 369.3000 ;
	    RECT 880.2000 363.3000 881.4000 376.5000 ;
	    RECT 916.3500 375.6000 917.2500 377.5500 ;
	    RECT 882.6000 374.4000 883.8000 375.6000 ;
	    RECT 916.2000 374.4000 917.4000 375.6000 ;
	    RECT 919.2000 375.3000 920.1000 380.4000 ;
	    RECT 921.0000 379.5000 922.2000 379.8000 ;
	    RECT 921.0000 378.4500 922.2000 378.6000 ;
	    RECT 925.9500 378.4500 926.8500 380.5500 ;
	    RECT 935.4000 380.4000 936.6000 380.5500 ;
	    RECT 990.6000 379.5000 991.8000 381.6000 ;
	    RECT 995.7000 380.7000 996.9000 381.6000 ;
	    RECT 1000.5000 380.7000 1001.7000 381.6000 ;
	    RECT 1005.9000 380.7000 1007.1000 381.6000 ;
	    RECT 993.0000 379.5000 996.9000 380.7000 ;
	    RECT 998.1000 379.5000 1001.7000 380.7000 ;
	    RECT 1003.2000 379.5000 1007.1000 380.7000 ;
	    RECT 1008.3000 379.5000 1008.9000 380.7000 ;
	    RECT 1031.4000 379.5000 1032.6000 383.7000 ;
	    RECT 1033.8000 382.5000 1035.0000 382.8000 ;
	    RECT 1060.5000 382.5000 1061.4000 383.7000 ;
	    RECT 1062.9000 383.1000 1068.3000 383.7000 ;
	    RECT 1079.4000 382.5000 1080.6000 389.7000 ;
	    RECT 1081.8000 386.7000 1083.0000 389.7000 ;
	    RECT 1081.8000 385.5000 1083.0000 385.8000 ;
	    RECT 1081.8000 384.4500 1083.0000 384.6000 ;
	    RECT 1093.8000 384.4500 1095.0000 384.6000 ;
	    RECT 1081.8000 383.5500 1095.0000 384.4500 ;
	    RECT 1101.0000 383.7000 1102.2001 389.7000 ;
	    RECT 1104.9000 384.6000 1106.1000 389.7000 ;
	    RECT 1117.8000 386.7000 1119.0000 389.7000 ;
	    RECT 1117.8000 385.5000 1119.0000 385.8000 ;
	    RECT 1103.4000 383.7000 1106.1000 384.6000 ;
	    RECT 1081.8000 383.4000 1083.0000 383.5500 ;
	    RECT 1093.8000 383.4000 1095.0000 383.5500 ;
	    RECT 1101.0000 382.5000 1102.2001 382.8000 ;
	    RECT 1033.8000 380.4000 1035.0000 381.6000 ;
	    RECT 1057.8000 381.4500 1059.0000 381.6000 ;
	    RECT 1060.2001 381.4500 1061.4000 381.6000 ;
	    RECT 1057.8000 380.5500 1061.4000 381.4500 ;
	    RECT 1057.8000 380.4000 1059.0000 380.5500 ;
	    RECT 1060.2001 380.4000 1061.4000 380.5500 ;
	    RECT 1062.3000 380.4000 1064.1000 381.6000 ;
	    RECT 1066.2001 380.7000 1066.5000 382.2000 ;
	    RECT 1067.4000 380.4000 1068.6000 381.6000 ;
	    RECT 1079.4000 381.4500 1080.6000 381.6000 ;
	    RECT 1069.9501 380.5500 1080.6000 381.4500 ;
	    RECT 921.0000 377.5500 926.8500 378.4500 ;
	    RECT 921.0000 377.4000 922.2000 377.5500 ;
	    RECT 919.2000 374.4000 920.7000 375.3000 ;
	    RECT 882.6000 373.2000 883.8000 373.5000 ;
	    RECT 917.4000 372.6000 918.3000 373.5000 ;
	    RECT 917.4000 371.4000 918.6000 372.6000 ;
	    RECT 882.6000 363.3000 883.8000 369.3000 ;
	    RECT 917.1000 363.3000 918.3000 369.3000 ;
	    RECT 919.5000 363.3000 920.7000 374.4000 ;
	    RECT 923.4000 363.3000 924.6000 375.3000 ;
	    RECT 935.4000 363.3000 936.6000 379.5000 ;
	    RECT 971.4000 378.4500 972.6000 378.6000 ;
	    RECT 990.6000 378.4500 991.8000 378.6000 ;
	    RECT 971.4000 377.5500 991.8000 378.4500 ;
	    RECT 971.4000 377.4000 972.6000 377.5500 ;
	    RECT 990.6000 377.4000 991.8000 377.5500 ;
	    RECT 995.7000 377.4000 996.9000 379.5000 ;
	    RECT 1000.5000 377.4000 1001.7000 379.5000 ;
	    RECT 1005.9000 377.4000 1007.1000 379.5000 ;
	    RECT 1031.4000 378.4500 1032.6000 378.6000 ;
	    RECT 1031.4000 377.5500 1061.2500 378.4500 ;
	    RECT 1031.4000 377.4000 1032.6000 377.5500 ;
	    RECT 992.7000 376.5000 994.2000 377.4000 ;
	    RECT 990.6000 376.2000 994.2000 376.5000 ;
	    RECT 995.7000 376.2000 999.0000 377.4000 ;
	    RECT 1000.5000 376.2000 1003.8000 377.4000 ;
	    RECT 1005.9000 376.2000 1008.6000 377.4000 ;
	    RECT 937.8000 363.3000 939.0000 369.3000 ;
	    RECT 990.6000 363.3000 991.8000 375.3000 ;
	    RECT 993.0000 363.3000 994.2000 376.2000 ;
	    RECT 995.4000 363.3000 996.6000 375.3000 ;
	    RECT 997.8000 363.3000 999.0000 376.2000 ;
	    RECT 1000.2000 363.3000 1001.4000 375.3000 ;
	    RECT 1002.6000 363.3000 1003.8000 376.2000 ;
	    RECT 1005.0000 363.3000 1006.2000 375.3000 ;
	    RECT 1007.4000 363.3000 1008.6000 376.2000 ;
	    RECT 1012.2000 375.4500 1013.4000 375.6000 ;
	    RECT 1029.0000 375.4500 1030.2001 375.6000 ;
	    RECT 1009.8000 363.3000 1011.0000 375.3000 ;
	    RECT 1012.2000 374.5500 1030.2001 375.4500 ;
	    RECT 1012.2000 374.4000 1013.4000 374.5500 ;
	    RECT 1029.0000 374.4000 1030.2001 374.5500 ;
	    RECT 1029.0000 373.2000 1030.2001 373.5000 ;
	    RECT 1029.0000 363.3000 1030.2001 369.3000 ;
	    RECT 1031.4000 363.3000 1032.6000 376.5000 ;
	    RECT 1060.3500 375.6000 1061.2500 377.5500 ;
	    RECT 1060.2001 374.4000 1061.4000 375.6000 ;
	    RECT 1063.2001 375.3000 1064.1000 380.4000 ;
	    RECT 1065.0000 379.5000 1066.2001 379.8000 ;
	    RECT 1065.0000 378.4500 1066.2001 378.6000 ;
	    RECT 1069.9501 378.4500 1070.8500 380.5500 ;
	    RECT 1079.4000 380.4000 1080.6000 380.5500 ;
	    RECT 1089.0000 381.4500 1090.2001 381.6000 ;
	    RECT 1101.0000 381.4500 1102.2001 381.6000 ;
	    RECT 1089.0000 380.5500 1102.2001 381.4500 ;
	    RECT 1089.0000 380.4000 1090.2001 380.5500 ;
	    RECT 1101.0000 380.4000 1102.2001 380.5500 ;
	    RECT 1103.4000 379.5000 1104.6000 383.7000 ;
	    RECT 1117.8000 383.4000 1119.0000 384.6000 ;
	    RECT 1120.2001 382.5000 1121.4000 389.7000 ;
	    RECT 1153.8000 383.7000 1155.0000 389.7000 ;
	    RECT 1156.2001 384.0000 1157.4000 389.7000 ;
	    RECT 1158.6000 384.9000 1159.8000 389.7000 ;
	    RECT 1161.0000 384.0000 1162.2001 389.7000 ;
	    RECT 1175.4000 386.7000 1176.6000 389.7000 ;
	    RECT 1175.4000 385.5000 1176.6000 385.8000 ;
	    RECT 1156.2001 383.7000 1162.2001 384.0000 ;
	    RECT 1165.8000 384.4500 1167.0000 384.6000 ;
	    RECT 1175.4000 384.4500 1176.6000 384.6000 ;
	    RECT 1154.1000 382.5000 1155.0000 383.7000 ;
	    RECT 1156.5000 383.1000 1161.9000 383.7000 ;
	    RECT 1165.8000 383.5500 1176.6000 384.4500 ;
	    RECT 1165.8000 383.4000 1167.0000 383.5500 ;
	    RECT 1175.4000 383.4000 1176.6000 383.5500 ;
	    RECT 1177.8000 382.5000 1179.0000 389.7000 ;
	    RECT 1192.2001 386.7000 1193.4000 389.7000 ;
	    RECT 1192.2001 385.5000 1193.4000 385.8000 ;
	    RECT 1180.2001 384.4500 1181.4000 384.6000 ;
	    RECT 1192.2001 384.4500 1193.4000 384.6000 ;
	    RECT 1180.2001 383.5500 1193.4000 384.4500 ;
	    RECT 1180.2001 383.4000 1181.4000 383.5500 ;
	    RECT 1192.2001 383.4000 1193.4000 383.5500 ;
	    RECT 1194.6000 382.5000 1195.8000 389.7000 ;
	    RECT 1249.8000 387.4500 1251.0000 387.6000 ;
	    RECT 1314.6000 387.4500 1315.8000 387.6000 ;
	    RECT 1249.8000 386.5500 1315.8000 387.4500 ;
	    RECT 1249.8000 386.4000 1251.0000 386.5500 ;
	    RECT 1314.6000 386.4000 1315.8000 386.5500 ;
	    RECT 1120.2001 381.4500 1121.4000 381.6000 ;
	    RECT 1151.4000 381.4500 1152.6000 381.6000 ;
	    RECT 1120.2001 380.5500 1152.6000 381.4500 ;
	    RECT 1120.2001 380.4000 1121.4000 380.5500 ;
	    RECT 1151.4000 380.4000 1152.6000 380.5500 ;
	    RECT 1153.8000 380.4000 1155.0000 381.6000 ;
	    RECT 1155.9000 380.4000 1157.7001 381.6000 ;
	    RECT 1159.8000 380.7000 1160.1000 382.2000 ;
	    RECT 1161.0000 381.4500 1162.2001 381.6000 ;
	    RECT 1170.6000 381.4500 1171.8000 381.6000 ;
	    RECT 1161.0000 380.5500 1171.8000 381.4500 ;
	    RECT 1161.0000 380.4000 1162.2001 380.5500 ;
	    RECT 1170.6000 380.4000 1171.8000 380.5500 ;
	    RECT 1177.8000 381.4500 1179.0000 381.6000 ;
	    RECT 1189.8000 381.4500 1191.0000 381.6000 ;
	    RECT 1177.8000 380.5500 1191.0000 381.4500 ;
	    RECT 1177.8000 380.4000 1179.0000 380.5500 ;
	    RECT 1189.8000 380.4000 1191.0000 380.5500 ;
	    RECT 1194.6000 381.4500 1195.8000 381.6000 ;
	    RECT 1317.0000 381.4500 1318.2001 381.6000 ;
	    RECT 1194.6000 380.5500 1318.2001 381.4500 ;
	    RECT 1194.6000 380.4000 1195.8000 380.5500 ;
	    RECT 1317.0000 380.4000 1318.2001 380.5500 ;
	    RECT 1319.4000 380.7000 1320.6000 389.7000 ;
	    RECT 1324.2001 383.7000 1325.4000 389.7000 ;
	    RECT 1329.0000 384.9000 1330.2001 389.7000 ;
	    RECT 1331.4000 385.5000 1332.6000 389.7000 ;
	    RECT 1333.8000 385.5000 1335.0000 389.7000 ;
	    RECT 1336.2001 385.5000 1337.4000 389.7000 ;
	    RECT 1338.6000 386.7000 1339.8000 389.7000 ;
	    RECT 1341.0000 385.5000 1342.2001 389.7000 ;
	    RECT 1343.4000 386.7000 1344.6000 389.7000 ;
	    RECT 1345.8000 385.5000 1347.0000 389.7000 ;
	    RECT 1348.2001 385.5000 1349.4000 389.7000 ;
	    RECT 1350.6000 385.5000 1351.8000 389.7000 ;
	    RECT 1353.0000 385.5000 1354.2001 389.7000 ;
	    RECT 1326.3000 383.7000 1330.2001 384.9000 ;
	    RECT 1355.4000 384.9000 1356.6000 389.7000 ;
	    RECT 1335.3000 383.7000 1342.2001 384.6000 ;
	    RECT 1326.3000 382.8000 1327.5000 383.7000 ;
	    RECT 1323.0000 381.6000 1327.5000 382.8000 ;
	    RECT 1065.0000 377.5500 1070.8500 378.4500 ;
	    RECT 1065.0000 377.4000 1066.2001 377.5500 ;
	    RECT 1063.2001 374.4000 1064.7001 375.3000 ;
	    RECT 1061.4000 372.6000 1062.3000 373.5000 ;
	    RECT 1061.4000 371.4000 1062.6000 372.6000 ;
	    RECT 1033.8000 363.3000 1035.0000 369.3000 ;
	    RECT 1061.1000 363.3000 1062.3000 369.3000 ;
	    RECT 1063.5000 363.3000 1064.7001 374.4000 ;
	    RECT 1067.4000 363.3000 1068.6000 375.3000 ;
	    RECT 1079.4000 363.3000 1080.6000 379.5000 ;
	    RECT 1103.4000 378.4500 1104.6000 378.6000 ;
	    RECT 1108.2001 378.4500 1109.4000 378.6000 ;
	    RECT 1103.4000 377.5500 1109.4000 378.4500 ;
	    RECT 1103.4000 377.4000 1104.6000 377.5500 ;
	    RECT 1108.2001 377.4000 1109.4000 377.5500 ;
	    RECT 1081.8000 363.3000 1083.0000 369.3000 ;
	    RECT 1101.0000 363.3000 1102.2001 369.3000 ;
	    RECT 1103.4000 363.3000 1104.6000 376.5000 ;
	    RECT 1105.8000 375.4500 1107.0000 375.6000 ;
	    RECT 1117.8000 375.4500 1119.0000 375.6000 ;
	    RECT 1105.8000 374.5500 1119.0000 375.4500 ;
	    RECT 1105.8000 374.4000 1107.0000 374.5500 ;
	    RECT 1117.8000 374.4000 1119.0000 374.5500 ;
	    RECT 1105.8000 373.2000 1107.0000 373.5000 ;
	    RECT 1105.8000 363.3000 1107.0000 369.3000 ;
	    RECT 1117.8000 363.3000 1119.0000 369.3000 ;
	    RECT 1120.2001 363.3000 1121.4000 379.5000 ;
	    RECT 1149.0000 375.4500 1150.2001 375.6000 ;
	    RECT 1153.8000 375.4500 1155.0000 375.6000 ;
	    RECT 1149.0000 374.5500 1155.0000 375.4500 ;
	    RECT 1149.0000 374.4000 1150.2001 374.5500 ;
	    RECT 1153.8000 374.4000 1155.0000 374.5500 ;
	    RECT 1156.8000 375.3000 1157.7001 380.4000 ;
	    RECT 1158.6000 379.5000 1159.8000 379.8000 ;
	    RECT 1319.4000 379.5000 1332.6000 380.7000 ;
	    RECT 1335.3000 380.1000 1336.5000 383.7000 ;
	    RECT 1341.0000 383.4000 1342.2001 383.7000 ;
	    RECT 1343.4000 383.4000 1344.6000 384.6000 ;
	    RECT 1345.5000 383.4000 1345.8000 384.6000 ;
	    RECT 1350.3000 383.4000 1351.8000 384.6000 ;
	    RECT 1355.4000 383.7000 1359.0000 384.9000 ;
	    RECT 1360.2001 383.7000 1361.4000 389.7000 ;
	    RECT 1338.6000 382.5000 1339.8000 382.8000 ;
	    RECT 1341.0000 382.2000 1342.2001 382.5000 ;
	    RECT 1338.6000 380.4000 1339.8000 381.6000 ;
	    RECT 1341.0000 381.3000 1347.6000 382.2000 ;
	    RECT 1346.4000 381.0000 1347.6000 381.3000 ;
	    RECT 1158.6000 377.4000 1159.8000 378.6000 ;
	    RECT 1156.8000 374.4000 1158.3000 375.3000 ;
	    RECT 1155.0000 372.6000 1155.9000 373.5000 ;
	    RECT 1155.0000 371.4000 1156.2001 372.6000 ;
	    RECT 1154.7001 363.3000 1155.9000 369.3000 ;
	    RECT 1157.1000 363.3000 1158.3000 374.4000 ;
	    RECT 1161.0000 363.3000 1162.2001 375.3000 ;
	    RECT 1175.4000 363.3000 1176.6000 369.3000 ;
	    RECT 1177.8000 363.3000 1179.0000 379.5000 ;
	    RECT 1192.2001 363.3000 1193.4000 369.3000 ;
	    RECT 1194.6000 363.3000 1195.8000 379.5000 ;
	    RECT 1276.2001 378.4500 1277.4000 378.6000 ;
	    RECT 1283.4000 378.4500 1284.6000 378.6000 ;
	    RECT 1276.2001 377.5500 1284.6000 378.4500 ;
	    RECT 1276.2001 377.4000 1277.4000 377.5500 ;
	    RECT 1283.4000 377.4000 1284.6000 377.5500 ;
	    RECT 1319.4000 371.1000 1320.6000 379.5000 ;
	    RECT 1333.5000 378.9000 1336.5000 380.1000 ;
	    RECT 1342.2001 378.9000 1347.0000 380.1000 ;
	    RECT 1350.6000 379.2000 1351.8000 383.4000 ;
	    RECT 1357.8000 382.8000 1359.0000 383.7000 ;
	    RECT 1357.8000 381.9000 1360.5000 382.8000 ;
	    RECT 1359.3000 380.1000 1360.5000 381.9000 ;
	    RECT 1365.0000 381.9000 1366.2001 389.7000 ;
	    RECT 1367.4000 384.0000 1368.6000 389.7000 ;
	    RECT 1369.8000 386.7000 1371.0000 389.7000 ;
	    RECT 1401.0000 384.0000 1402.2001 389.7000 ;
	    RECT 1403.4000 384.9000 1404.6000 389.7000 ;
	    RECT 1405.8000 384.0000 1407.0000 389.7000 ;
	    RECT 1367.4000 382.8000 1368.9000 384.0000 ;
	    RECT 1401.0000 383.7000 1407.0000 384.0000 ;
	    RECT 1408.2001 383.7000 1409.4000 389.7000 ;
	    RECT 1432.2001 384.0000 1433.4000 389.7000 ;
	    RECT 1434.6000 384.9000 1435.8000 389.7000 ;
	    RECT 1437.0000 384.0000 1438.2001 389.7000 ;
	    RECT 1432.2001 383.7000 1438.2001 384.0000 ;
	    RECT 1439.4000 383.7000 1440.6000 389.7000 ;
	    RECT 1459.5000 384.6000 1460.7001 389.7000 ;
	    RECT 1459.5000 383.7000 1462.2001 384.6000 ;
	    RECT 1463.4000 383.7000 1464.6000 389.7000 ;
	    RECT 1482.6000 386.7000 1483.8000 389.7000 ;
	    RECT 1485.0000 386.7000 1486.2001 389.7000 ;
	    RECT 1487.4000 386.7000 1488.6000 389.7000 ;
	    RECT 1501.8000 386.7000 1503.0000 389.7000 ;
	    RECT 1482.6000 385.5000 1483.8000 385.8000 ;
	    RECT 1401.3000 383.1000 1406.7001 383.7000 ;
	    RECT 1365.0000 381.0000 1366.8000 381.9000 ;
	    RECT 1359.3000 378.9000 1365.0000 380.1000 ;
	    RECT 1321.5000 378.0000 1322.7001 378.3000 ;
	    RECT 1321.5000 377.1000 1328.1000 378.0000 ;
	    RECT 1329.0000 377.4000 1330.2001 378.6000 ;
	    RECT 1355.4000 378.0000 1356.6000 378.9000 ;
	    RECT 1365.9000 378.0000 1366.8000 381.0000 ;
	    RECT 1331.1000 377.1000 1356.6000 378.0000 ;
	    RECT 1365.6000 377.1000 1366.8000 378.0000 ;
	    RECT 1363.5000 376.2000 1364.7001 376.5000 ;
	    RECT 1324.2001 374.4000 1325.4000 375.6000 ;
	    RECT 1326.3000 375.3000 1364.7001 376.2000 ;
	    RECT 1329.3000 375.0000 1330.5000 375.3000 ;
	    RECT 1365.6000 374.4000 1366.5000 377.1000 ;
	    RECT 1367.7001 376.2000 1368.9000 382.8000 ;
	    RECT 1408.2001 382.5000 1409.1000 383.7000 ;
	    RECT 1432.5000 383.1000 1437.9000 383.7000 ;
	    RECT 1439.4000 382.5000 1440.3000 383.7000 ;
	    RECT 1386.6000 381.4500 1387.8000 381.6000 ;
	    RECT 1401.0000 381.4500 1402.2001 381.6000 ;
	    RECT 1386.6000 380.5500 1402.2001 381.4500 ;
	    RECT 1403.1000 380.7000 1403.4000 382.2000 ;
	    RECT 1386.6000 380.4000 1387.8000 380.5500 ;
	    RECT 1401.0000 380.4000 1402.2001 380.5500 ;
	    RECT 1405.5000 380.4000 1407.3000 381.6000 ;
	    RECT 1408.2001 381.4500 1409.4000 381.6000 ;
	    RECT 1417.8000 381.4500 1419.0000 381.6000 ;
	    RECT 1408.2001 380.5500 1419.0000 381.4500 ;
	    RECT 1408.2001 380.4000 1409.4000 380.5500 ;
	    RECT 1417.8000 380.4000 1419.0000 380.5500 ;
	    RECT 1422.6000 381.4500 1423.8000 381.6000 ;
	    RECT 1432.2001 381.4500 1433.4000 381.6000 ;
	    RECT 1422.6000 380.5500 1433.4000 381.4500 ;
	    RECT 1434.3000 380.7000 1434.6000 382.2000 ;
	    RECT 1422.6000 380.4000 1423.8000 380.5500 ;
	    RECT 1432.2001 380.4000 1433.4000 380.5500 ;
	    RECT 1436.7001 380.4000 1438.5000 381.6000 ;
	    RECT 1439.4000 381.4500 1440.6000 381.6000 ;
	    RECT 1449.0000 381.4500 1450.2001 381.6000 ;
	    RECT 1439.4000 380.5500 1450.2001 381.4500 ;
	    RECT 1439.4000 380.4000 1440.6000 380.5500 ;
	    RECT 1449.0000 380.4000 1450.2001 380.5500 ;
	    RECT 1403.4000 379.5000 1404.6000 379.8000 ;
	    RECT 1393.8000 378.4500 1395.0000 378.6000 ;
	    RECT 1403.4000 378.4500 1404.6000 378.6000 ;
	    RECT 1393.8000 377.5500 1404.6000 378.4500 ;
	    RECT 1393.8000 377.4000 1395.0000 377.5500 ;
	    RECT 1403.4000 377.4000 1404.6000 377.5500 ;
	    RECT 1333.8000 374.1000 1335.0000 374.4000 ;
	    RECT 1326.9000 373.5000 1335.0000 374.1000 ;
	    RECT 1325.7001 373.2000 1335.0000 373.5000 ;
	    RECT 1336.5000 373.5000 1349.4000 374.4000 ;
	    RECT 1321.8000 372.0000 1324.2001 373.2000 ;
	    RECT 1325.7001 372.3000 1327.8000 373.2000 ;
	    RECT 1336.5000 372.3000 1337.4000 373.5000 ;
	    RECT 1348.2001 373.2000 1349.4000 373.5000 ;
	    RECT 1353.0000 373.5000 1366.5000 374.4000 ;
	    RECT 1367.4000 375.0000 1368.9000 376.2000 ;
	    RECT 1405.5000 375.3000 1406.4000 380.4000 ;
	    RECT 1434.6000 379.5000 1435.8000 379.8000 ;
	    RECT 1434.6000 377.4000 1435.8000 378.6000 ;
	    RECT 1367.4000 373.5000 1368.6000 375.0000 ;
	    RECT 1353.0000 373.2000 1354.2001 373.5000 ;
	    RECT 1323.3000 371.4000 1324.2001 372.0000 ;
	    RECT 1328.7001 371.4000 1337.4000 372.3000 ;
	    RECT 1338.3000 371.4000 1342.2001 372.6000 ;
	    RECT 1319.4000 370.2000 1322.4000 371.1000 ;
	    RECT 1323.3000 370.2000 1329.6000 371.4000 ;
	    RECT 1257.0000 369.4500 1258.2001 369.6000 ;
	    RECT 1312.2001 369.4500 1313.4000 369.6000 ;
	    RECT 1257.0000 368.5500 1313.4000 369.4500 ;
	    RECT 1321.5000 369.3000 1322.4000 370.2000 ;
	    RECT 1257.0000 368.4000 1258.2001 368.5500 ;
	    RECT 1312.2001 368.4000 1313.4000 368.5500 ;
	    RECT 1319.4000 363.3000 1320.6000 369.3000 ;
	    RECT 1321.5000 368.4000 1323.0000 369.3000 ;
	    RECT 1321.8000 363.3000 1323.0000 368.4000 ;
	    RECT 1324.2001 362.4000 1325.4000 369.3000 ;
	    RECT 1326.6000 363.3000 1327.8000 370.2000 ;
	    RECT 1329.0000 363.3000 1330.2001 369.3000 ;
	    RECT 1331.4000 363.3000 1332.6000 367.5000 ;
	    RECT 1333.8000 363.3000 1335.0000 367.5000 ;
	    RECT 1336.2001 363.3000 1337.4000 370.5000 ;
	    RECT 1338.6000 363.3000 1339.8000 369.3000 ;
	    RECT 1341.0000 363.3000 1342.2001 370.5000 ;
	    RECT 1343.4000 363.3000 1344.6000 369.3000 ;
	    RECT 1345.8000 363.3000 1347.0000 372.6000 ;
	    RECT 1357.8000 371.4000 1361.7001 372.6000 ;
	    RECT 1350.6000 370.2000 1356.9000 371.4000 ;
	    RECT 1348.2001 363.3000 1349.4000 367.5000 ;
	    RECT 1350.6000 363.3000 1351.8000 367.5000 ;
	    RECT 1353.0000 363.3000 1354.2001 367.5000 ;
	    RECT 1355.4000 363.3000 1356.6000 369.3000 ;
	    RECT 1357.8000 363.3000 1359.0000 371.4000 ;
	    RECT 1365.6000 371.1000 1366.5000 373.5000 ;
	    RECT 1367.4000 371.4000 1368.6000 372.6000 ;
	    RECT 1362.6000 370.2000 1366.5000 371.1000 ;
	    RECT 1360.2001 363.3000 1361.4000 369.3000 ;
	    RECT 1362.6000 363.3000 1363.8000 370.2000 ;
	    RECT 1365.0000 363.3000 1366.2001 369.3000 ;
	    RECT 1367.4000 363.3000 1368.6000 370.5000 ;
	    RECT 1369.8000 363.3000 1371.0000 369.3000 ;
	    RECT 1401.0000 363.3000 1402.2001 375.3000 ;
	    RECT 1404.9000 374.4000 1406.4000 375.3000 ;
	    RECT 1408.2001 374.4000 1409.4000 375.6000 ;
	    RECT 1436.7001 375.3000 1437.6000 380.4000 ;
	    RECT 1461.0000 379.5000 1462.2001 383.7000 ;
	    RECT 1482.6000 383.4000 1483.8000 384.6000 ;
	    RECT 1463.4000 382.5000 1464.6000 382.8000 ;
	    RECT 1485.3000 382.5000 1486.2001 386.7000 ;
	    RECT 1501.8000 385.5000 1503.0000 385.8000 ;
	    RECT 1489.8000 384.4500 1491.0000 384.6000 ;
	    RECT 1501.8000 384.4500 1503.0000 384.6000 ;
	    RECT 1489.8000 383.5500 1503.0000 384.4500 ;
	    RECT 1489.8000 383.4000 1491.0000 383.5500 ;
	    RECT 1501.8000 383.4000 1503.0000 383.5500 ;
	    RECT 1504.2001 382.5000 1505.4000 389.7000 ;
	    RECT 1463.4000 381.4500 1464.6000 381.6000 ;
	    RECT 1470.6000 381.4500 1471.8000 381.6000 ;
	    RECT 1485.0000 381.4500 1486.2001 381.6000 ;
	    RECT 1463.4000 380.5500 1486.2001 381.4500 ;
	    RECT 1463.4000 380.4000 1464.6000 380.5500 ;
	    RECT 1470.6000 380.4000 1471.8000 380.5500 ;
	    RECT 1485.0000 380.4000 1486.2001 380.5500 ;
	    RECT 1504.2001 381.4500 1505.4000 381.6000 ;
	    RECT 1518.6000 381.4500 1519.8000 381.6000 ;
	    RECT 1504.2001 380.5500 1519.8000 381.4500 ;
	    RECT 1532.4000 381.3000 1533.6000 389.7000 ;
	    RECT 1504.2001 380.4000 1505.4000 380.5500 ;
	    RECT 1518.6000 380.4000 1519.8000 380.5500 ;
	    RECT 1530.9000 380.7000 1533.6000 381.3000 ;
	    RECT 1537.8000 380.7000 1539.0000 389.7000 ;
	    RECT 1557.9000 384.6000 1559.1000 389.7000 ;
	    RECT 1557.9000 383.7000 1560.6000 384.6000 ;
	    RECT 1561.8000 383.7000 1563.0000 389.7000 ;
	    RECT 1530.9000 380.4000 1533.3000 380.7000 ;
	    RECT 1461.0000 377.4000 1462.2001 378.6000 ;
	    RECT 1404.9000 363.3000 1406.1000 374.4000 ;
	    RECT 1407.3000 372.6000 1408.2001 373.5000 ;
	    RECT 1407.0000 371.4000 1408.2001 372.6000 ;
	    RECT 1407.3000 363.3000 1408.5000 369.3000 ;
	    RECT 1432.2001 363.3000 1433.4000 375.3000 ;
	    RECT 1436.1000 374.4000 1437.6000 375.3000 ;
	    RECT 1439.4000 375.4500 1440.6000 375.6000 ;
	    RECT 1446.6000 375.4500 1447.8000 375.6000 ;
	    RECT 1458.6000 375.4500 1459.8000 375.6000 ;
	    RECT 1439.4000 374.5500 1459.8000 375.4500 ;
	    RECT 1439.4000 374.4000 1440.6000 374.5500 ;
	    RECT 1446.6000 374.4000 1447.8000 374.5500 ;
	    RECT 1458.6000 374.4000 1459.8000 374.5500 ;
	    RECT 1436.1000 363.3000 1437.3000 374.4000 ;
	    RECT 1438.5000 372.6000 1439.4000 373.5000 ;
	    RECT 1458.6000 373.2000 1459.8000 373.5000 ;
	    RECT 1438.2001 371.4000 1439.4000 372.6000 ;
	    RECT 1438.5000 363.3000 1439.7001 369.3000 ;
	    RECT 1458.6000 363.3000 1459.8000 369.3000 ;
	    RECT 1461.0000 363.3000 1462.2001 376.5000 ;
	    RECT 1485.3000 375.3000 1486.2001 379.5000 ;
	    RECT 1487.4000 377.4000 1488.6000 378.6000 ;
	    RECT 1487.4000 376.2000 1488.6000 376.5000 ;
	    RECT 1463.4000 363.3000 1464.6000 369.3000 ;
	    RECT 1482.6000 363.3000 1483.8000 375.3000 ;
	    RECT 1485.0000 374.1000 1487.7001 375.3000 ;
	    RECT 1486.5000 363.3000 1487.7001 374.1000 ;
	    RECT 1501.8000 363.3000 1503.0000 369.3000 ;
	    RECT 1504.2001 363.3000 1505.4000 379.5000 ;
	    RECT 1530.9000 376.5000 1531.8000 380.4000 ;
	    RECT 1559.4000 379.5000 1560.6000 383.7000 ;
	    RECT 1561.8000 382.5000 1563.0000 382.8000 ;
	    RECT 1561.8000 380.4000 1563.0000 381.6000 ;
	    RECT 1534.2001 377.4000 1534.5000 378.6000 ;
	    RECT 1535.4000 377.4000 1536.6000 378.6000 ;
	    RECT 1552.2001 378.4500 1553.4000 378.6000 ;
	    RECT 1559.4000 378.4500 1560.6000 378.6000 ;
	    RECT 1552.2001 377.5500 1560.6000 378.4500 ;
	    RECT 1552.2001 377.4000 1553.4000 377.5500 ;
	    RECT 1559.4000 377.4000 1560.6000 377.5500 ;
	    RECT 1537.8000 376.5000 1539.0000 376.8000 ;
	    RECT 1509.0000 375.4500 1510.2001 375.6000 ;
	    RECT 1530.6000 375.4500 1531.8000 375.6000 ;
	    RECT 1509.0000 374.5500 1531.8000 375.4500 ;
	    RECT 1509.0000 374.4000 1510.2001 374.5500 ;
	    RECT 1530.6000 374.4000 1531.8000 374.5500 ;
	    RECT 1537.8000 374.4000 1539.0000 375.6000 ;
	    RECT 1557.0000 375.4500 1558.2001 375.6000 ;
	    RECT 1545.1500 374.5500 1558.2001 375.4500 ;
	    RECT 1533.0000 373.5000 1534.2001 373.8000 ;
	    RECT 1530.9000 370.5000 1531.8000 373.5000 ;
	    RECT 1533.0000 371.4000 1534.2001 372.6000 ;
	    RECT 1535.4000 372.4500 1536.6000 372.6000 ;
	    RECT 1545.1500 372.4500 1546.0500 374.5500 ;
	    RECT 1557.0000 374.4000 1558.2001 374.5500 ;
	    RECT 1557.0000 373.2000 1558.2001 373.5000 ;
	    RECT 1535.4000 371.5500 1546.0500 372.4500 ;
	    RECT 1535.4000 371.4000 1536.6000 371.5500 ;
	    RECT 1530.9000 369.6000 1536.3000 370.5000 ;
	    RECT 1530.9000 369.3000 1531.8000 369.6000 ;
	    RECT 1530.6000 363.3000 1531.8000 369.3000 ;
	    RECT 1535.4000 369.3000 1536.3000 369.6000 ;
	    RECT 1533.0000 363.3000 1534.2001 368.7000 ;
	    RECT 1535.4000 363.3000 1536.6000 369.3000 ;
	    RECT 1537.8000 363.3000 1539.0000 369.3000 ;
	    RECT 1557.0000 363.3000 1558.2001 369.3000 ;
	    RECT 1559.4000 363.3000 1560.6000 376.5000 ;
	    RECT 1561.8000 363.3000 1563.0000 369.3000 ;
	    RECT 1.2000 360.6000 1569.0000 362.4000 ;
	    RECT 18.6000 347.7000 19.8000 359.7000 ;
	    RECT 21.0000 349.5000 22.2000 359.7000 ;
	    RECT 23.4000 348.6000 24.6000 359.7000 ;
	    RECT 42.6000 353.7000 43.8000 359.7000 ;
	    RECT 42.6000 349.5000 43.8000 349.8000 ;
	    RECT 21.3000 347.7000 24.6000 348.6000 ;
	    RECT 40.2000 348.4500 41.4000 348.6000 ;
	    RECT 42.6000 348.4500 43.8000 348.6000 ;
	    RECT 18.6000 344.4000 19.5000 347.7000 ;
	    RECT 21.3000 346.8000 22.2000 347.7000 ;
	    RECT 40.2000 347.5500 43.8000 348.4500 ;
	    RECT 40.2000 347.4000 41.4000 347.5500 ;
	    RECT 42.6000 347.4000 43.8000 347.5500 ;
	    RECT 20.4000 345.6000 22.2000 346.8000 ;
	    RECT 45.0000 346.5000 46.2000 359.7000 ;
	    RECT 47.4000 353.7000 48.6000 359.7000 ;
	    RECT 66.6000 348.6000 67.8000 359.7000 ;
	    RECT 69.0000 349.5000 70.2000 359.7000 ;
	    RECT 66.6000 347.7000 69.9000 348.6000 ;
	    RECT 71.4000 347.7000 72.6000 359.7000 ;
	    RECT 83.4000 353.7000 84.6000 359.7000 ;
	    RECT 69.0000 346.8000 69.9000 347.7000 ;
	    RECT 69.0000 345.6000 70.8000 346.8000 ;
	    RECT 18.6000 343.5000 19.8000 344.4000 ;
	    RECT 18.6000 341.4000 19.8000 342.6000 ;
	    RECT 21.3000 341.1000 22.2000 345.6000 ;
	    RECT 23.4000 344.4000 24.6000 345.6000 ;
	    RECT 30.6000 345.4500 31.8000 345.6000 ;
	    RECT 45.0000 345.4500 46.2000 345.6000 ;
	    RECT 30.6000 344.5500 46.2000 345.4500 ;
	    RECT 30.6000 344.4000 31.8000 344.5500 ;
	    RECT 45.0000 344.4000 46.2000 344.5500 ;
	    RECT 66.6000 344.4000 67.8000 345.6000 ;
	    RECT 23.4000 343.2000 24.6000 343.5000 ;
	    RECT 18.6000 333.3000 19.8000 340.5000 ;
	    RECT 21.3000 340.2000 24.6000 341.1000 ;
	    RECT 21.0000 333.3000 22.2000 339.3000 ;
	    RECT 23.4000 333.3000 24.6000 340.2000 ;
	    RECT 45.0000 339.3000 46.2000 343.5000 ;
	    RECT 66.6000 343.2000 67.8000 343.5000 ;
	    RECT 47.4000 341.4000 48.6000 342.6000 ;
	    RECT 69.0000 341.1000 69.9000 345.6000 ;
	    RECT 71.7000 344.4000 72.6000 347.7000 ;
	    RECT 71.4000 343.5000 72.6000 344.4000 ;
	    RECT 85.8000 343.5000 87.0000 359.7000 ;
	    RECT 109.8000 347.7000 111.0000 359.7000 ;
	    RECT 113.7000 348.6000 114.9000 359.7000 ;
	    RECT 116.1000 353.7000 117.3000 359.7000 ;
	    RECT 115.8000 350.4000 117.0000 351.6000 ;
	    RECT 116.1000 349.5000 117.0000 350.4000 ;
	    RECT 113.7000 347.7000 115.2000 348.6000 ;
	    RECT 112.2000 344.4000 113.4000 345.6000 ;
	    RECT 112.2000 343.2000 113.4000 343.5000 ;
	    RECT 114.3000 342.6000 115.2000 347.7000 ;
	    RECT 117.0000 348.4500 118.2000 348.6000 ;
	    RECT 121.8000 348.4500 123.0000 348.6000 ;
	    RECT 117.0000 347.5500 123.0000 348.4500 ;
	    RECT 117.0000 347.4000 118.2000 347.5500 ;
	    RECT 121.8000 347.4000 123.0000 347.5500 ;
	    RECT 131.4000 343.5000 132.6000 359.7000 ;
	    RECT 133.8000 353.7000 135.0000 359.7000 ;
	    RECT 161.1000 353.7000 162.3000 359.7000 ;
	    RECT 161.4000 350.4000 162.6000 351.6000 ;
	    RECT 161.4000 349.5000 162.3000 350.4000 ;
	    RECT 163.5000 348.6000 164.7000 359.7000 ;
	    RECT 160.2000 347.4000 161.4000 348.6000 ;
	    RECT 163.2000 347.7000 164.7000 348.6000 ;
	    RECT 167.4000 347.7000 168.6000 359.7000 ;
	    RECT 163.2000 342.6000 164.1000 347.7000 ;
	    RECT 165.0000 345.4500 166.2000 345.6000 ;
	    RECT 165.0000 344.5500 170.8500 345.4500 ;
	    RECT 165.0000 344.4000 166.2000 344.5500 ;
	    RECT 165.0000 343.2000 166.2000 343.5000 ;
	    RECT 71.4000 341.4000 72.6000 342.6000 ;
	    RECT 85.8000 342.4500 87.0000 342.6000 ;
	    RECT 107.4000 342.4500 108.6000 342.6000 ;
	    RECT 85.8000 341.5500 108.6000 342.4500 ;
	    RECT 85.8000 341.4000 87.0000 341.5500 ;
	    RECT 107.4000 341.4000 108.6000 341.5500 ;
	    RECT 109.8000 341.4000 111.0000 342.6000 ;
	    RECT 47.4000 340.2000 48.6000 340.5000 ;
	    RECT 66.6000 340.2000 69.9000 341.1000 ;
	    RECT 111.9000 340.8000 112.2000 342.3000 ;
	    RECT 114.3000 341.4000 116.1000 342.6000 ;
	    RECT 117.0000 341.4000 118.2000 342.6000 ;
	    RECT 119.4000 342.4500 120.6000 342.6000 ;
	    RECT 131.4000 342.4500 132.6000 342.6000 ;
	    RECT 119.4000 341.5500 132.6000 342.4500 ;
	    RECT 119.4000 341.4000 120.6000 341.5500 ;
	    RECT 131.4000 341.4000 132.6000 341.5500 ;
	    RECT 160.2000 341.4000 161.4000 342.6000 ;
	    RECT 162.3000 341.4000 164.1000 342.6000 ;
	    RECT 166.2000 340.8000 166.5000 342.3000 ;
	    RECT 167.4000 341.4000 168.6000 342.6000 ;
	    RECT 169.9500 342.4500 170.8500 344.5500 ;
	    RECT 179.4000 343.5000 180.6000 359.7000 ;
	    RECT 181.8000 353.7000 183.0000 359.7000 ;
	    RECT 196.2000 343.5000 197.4000 359.7000 ;
	    RECT 198.6000 353.7000 199.8000 359.7000 ;
	    RECT 258.6000 347.7000 259.8000 359.7000 ;
	    RECT 261.0000 346.8000 262.2000 359.7000 ;
	    RECT 263.4000 347.7000 264.6000 359.7000 ;
	    RECT 265.8000 346.8000 267.0000 359.7000 ;
	    RECT 268.2000 347.7000 269.4000 359.7000 ;
	    RECT 270.6000 346.8000 271.8000 359.7000 ;
	    RECT 273.0000 347.7000 274.2000 359.7000 ;
	    RECT 275.4000 346.8000 276.6000 359.7000 ;
	    RECT 277.8000 347.7000 279.0000 359.7000 ;
	    RECT 261.0000 345.6000 263.7000 346.8000 ;
	    RECT 265.8000 345.6000 269.1000 346.8000 ;
	    RECT 270.6000 345.6000 273.9000 346.8000 ;
	    RECT 275.4000 346.5000 279.0000 346.8000 ;
	    RECT 275.4000 345.6000 276.9000 346.5000 ;
	    RECT 262.5000 343.5000 263.7000 345.6000 ;
	    RECT 267.9000 343.5000 269.1000 345.6000 ;
	    RECT 272.7000 343.5000 273.9000 345.6000 ;
	    RECT 277.8000 345.4500 279.0000 345.6000 ;
	    RECT 287.4000 345.4500 288.6000 345.6000 ;
	    RECT 277.8000 344.5500 288.6000 345.4500 ;
	    RECT 277.8000 344.4000 279.0000 344.5500 ;
	    RECT 287.4000 344.4000 288.6000 344.5500 ;
	    RECT 292.2000 343.5000 293.4000 359.7000 ;
	    RECT 294.6000 353.7000 295.8000 359.7000 ;
	    RECT 313.8000 347.7000 315.0000 359.7000 ;
	    RECT 316.2000 349.5000 317.4000 359.7000 ;
	    RECT 318.6000 348.6000 319.8000 359.7000 ;
	    RECT 337.8000 353.7000 339.0000 359.7000 ;
	    RECT 316.5000 347.7000 319.8000 348.6000 ;
	    RECT 313.8000 344.4000 314.7000 347.7000 ;
	    RECT 316.5000 346.8000 317.4000 347.7000 ;
	    RECT 315.6000 345.6000 317.4000 346.8000 ;
	    RECT 340.2000 346.5000 341.4000 359.7000 ;
	    RECT 342.6000 353.7000 343.8000 359.7000 ;
	    RECT 347.4000 359.4000 348.6000 360.6000 ;
	    RECT 357.0000 353.7000 358.2000 359.7000 ;
	    RECT 342.6000 349.5000 343.8000 349.8000 ;
	    RECT 342.6000 348.4500 343.8000 348.6000 ;
	    RECT 347.4000 348.4500 348.6000 348.6000 ;
	    RECT 342.6000 347.5500 348.6000 348.4500 ;
	    RECT 342.6000 347.4000 343.8000 347.5500 ;
	    RECT 347.4000 347.4000 348.6000 347.5500 ;
	    RECT 313.8000 343.5000 315.0000 344.4000 ;
	    RECT 179.4000 342.4500 180.6000 342.6000 ;
	    RECT 169.9500 341.5500 180.6000 342.4500 ;
	    RECT 179.4000 341.4000 180.6000 341.5500 ;
	    RECT 189.0000 342.4500 190.2000 342.6000 ;
	    RECT 196.2000 342.4500 197.4000 342.6000 ;
	    RECT 189.0000 341.5500 197.4000 342.4500 ;
	    RECT 189.0000 341.4000 190.2000 341.5500 ;
	    RECT 196.2000 341.4000 197.4000 341.5500 ;
	    RECT 229.8000 342.4500 231.0000 342.6000 ;
	    RECT 258.6000 342.4500 259.8000 342.6000 ;
	    RECT 229.8000 341.5500 259.8000 342.4500 ;
	    RECT 260.7000 342.3000 261.3000 343.5000 ;
	    RECT 262.5000 342.3000 266.4000 343.5000 ;
	    RECT 267.9000 342.3000 271.5000 343.5000 ;
	    RECT 272.7000 342.3000 276.6000 343.5000 ;
	    RECT 229.8000 341.4000 231.0000 341.5500 ;
	    RECT 258.6000 341.4000 259.8000 341.5500 ;
	    RECT 262.5000 341.4000 263.7000 342.3000 ;
	    RECT 267.9000 341.4000 269.1000 342.3000 ;
	    RECT 272.7000 341.4000 273.9000 342.3000 ;
	    RECT 277.8000 341.4000 279.0000 343.5000 ;
	    RECT 280.2000 342.4500 281.4000 342.6000 ;
	    RECT 292.2000 342.4500 293.4000 342.6000 ;
	    RECT 280.2000 341.5500 293.4000 342.4500 ;
	    RECT 280.2000 341.4000 281.4000 341.5500 ;
	    RECT 292.2000 341.4000 293.4000 341.5500 ;
	    RECT 301.8000 342.4500 303.0000 342.6000 ;
	    RECT 313.8000 342.4500 315.0000 342.6000 ;
	    RECT 301.8000 341.5500 315.0000 342.4500 ;
	    RECT 301.8000 341.4000 303.0000 341.5500 ;
	    RECT 313.8000 341.4000 315.0000 341.5500 ;
	    RECT 43.5000 338.4000 46.2000 339.3000 ;
	    RECT 43.5000 333.3000 44.7000 338.4000 ;
	    RECT 47.4000 333.3000 48.6000 339.3000 ;
	    RECT 66.6000 333.3000 67.8000 340.2000 ;
	    RECT 69.0000 333.3000 70.2000 339.3000 ;
	    RECT 71.4000 333.3000 72.6000 340.5000 ;
	    RECT 73.8000 339.4500 75.0000 339.6000 ;
	    RECT 83.4000 339.4500 84.6000 339.6000 ;
	    RECT 73.8000 338.5500 84.6000 339.4500 ;
	    RECT 73.8000 338.4000 75.0000 338.5500 ;
	    RECT 83.4000 338.4000 84.6000 338.5500 ;
	    RECT 83.4000 337.2000 84.6000 337.5000 ;
	    RECT 83.4000 333.3000 84.6000 336.3000 ;
	    RECT 85.8000 333.3000 87.0000 340.5000 ;
	    RECT 110.1000 339.3000 115.5000 339.9000 ;
	    RECT 117.0000 339.3000 117.9000 340.5000 ;
	    RECT 109.8000 339.0000 115.8000 339.3000 ;
	    RECT 109.8000 333.3000 111.0000 339.0000 ;
	    RECT 112.2000 333.3000 113.4000 338.1000 ;
	    RECT 114.6000 333.3000 115.8000 339.0000 ;
	    RECT 117.0000 333.3000 118.2000 339.3000 ;
	    RECT 131.4000 333.3000 132.6000 340.5000 ;
	    RECT 133.8000 339.4500 135.0000 339.6000 ;
	    RECT 157.8000 339.4500 159.0000 339.6000 ;
	    RECT 133.8000 338.5500 159.0000 339.4500 ;
	    RECT 160.5000 339.3000 161.4000 340.5000 ;
	    RECT 162.9000 339.3000 168.3000 339.9000 ;
	    RECT 133.8000 338.4000 135.0000 338.5500 ;
	    RECT 157.8000 338.4000 159.0000 338.5500 ;
	    RECT 133.8000 337.2000 135.0000 337.5000 ;
	    RECT 133.8000 333.3000 135.0000 336.3000 ;
	    RECT 160.2000 333.3000 161.4000 339.3000 ;
	    RECT 162.6000 339.0000 168.6000 339.3000 ;
	    RECT 162.6000 333.3000 163.8000 339.0000 ;
	    RECT 165.0000 333.3000 166.2000 338.1000 ;
	    RECT 167.4000 333.3000 168.6000 339.0000 ;
	    RECT 179.4000 333.3000 180.6000 340.5000 ;
	    RECT 181.8000 339.4500 183.0000 339.6000 ;
	    RECT 193.8000 339.4500 195.0000 339.6000 ;
	    RECT 181.8000 338.5500 195.0000 339.4500 ;
	    RECT 181.8000 338.4000 183.0000 338.5500 ;
	    RECT 193.8000 338.4000 195.0000 338.5500 ;
	    RECT 181.8000 337.2000 183.0000 337.5000 ;
	    RECT 181.8000 333.3000 183.0000 336.3000 ;
	    RECT 196.2000 333.3000 197.4000 340.5000 ;
	    RECT 261.0000 340.2000 263.7000 341.4000 ;
	    RECT 265.8000 340.2000 269.1000 341.4000 ;
	    RECT 270.6000 340.2000 273.9000 341.4000 ;
	    RECT 275.4000 340.2000 279.0000 341.4000 ;
	    RECT 316.5000 341.1000 317.4000 345.6000 ;
	    RECT 318.6000 345.4500 319.8000 345.6000 ;
	    RECT 323.4000 345.4500 324.6000 345.6000 ;
	    RECT 318.6000 344.5500 324.6000 345.4500 ;
	    RECT 318.6000 344.4000 319.8000 344.5500 ;
	    RECT 323.4000 344.4000 324.6000 344.5500 ;
	    RECT 340.2000 345.4500 341.4000 345.6000 ;
	    RECT 342.6000 345.4500 343.8000 345.6000 ;
	    RECT 340.2000 344.5500 343.8000 345.4500 ;
	    RECT 340.2000 344.4000 341.4000 344.5500 ;
	    RECT 342.6000 344.4000 343.8000 344.5500 ;
	    RECT 359.4000 343.5000 360.6000 359.7000 ;
	    RECT 384.3000 353.7000 385.5000 359.7000 ;
	    RECT 384.6000 350.4000 385.8000 351.6000 ;
	    RECT 384.6000 349.5000 385.5000 350.4000 ;
	    RECT 386.7000 348.6000 387.9000 359.7000 ;
	    RECT 383.4000 347.4000 384.6000 348.6000 ;
	    RECT 386.4000 347.7000 387.9000 348.6000 ;
	    RECT 390.6000 347.7000 391.8000 359.7000 ;
	    RECT 409.8000 353.7000 411.0000 359.7000 ;
	    RECT 318.6000 343.2000 319.8000 343.5000 ;
	    RECT 333.0000 342.4500 334.2000 342.6000 ;
	    RECT 337.8000 342.4500 339.0000 342.6000 ;
	    RECT 333.0000 341.5500 339.0000 342.4500 ;
	    RECT 333.0000 341.4000 334.2000 341.5500 ;
	    RECT 337.8000 341.4000 339.0000 341.5500 ;
	    RECT 198.6000 338.4000 199.8000 339.6000 ;
	    RECT 198.6000 337.2000 199.8000 337.5000 ;
	    RECT 198.6000 333.3000 199.8000 336.3000 ;
	    RECT 258.6000 333.3000 259.8000 339.3000 ;
	    RECT 261.0000 333.3000 262.2000 340.2000 ;
	    RECT 263.4000 333.3000 264.6000 339.3000 ;
	    RECT 265.8000 333.3000 267.0000 340.2000 ;
	    RECT 268.2000 333.3000 269.4000 339.3000 ;
	    RECT 270.6000 333.3000 271.8000 340.2000 ;
	    RECT 273.0000 333.3000 274.2000 339.3000 ;
	    RECT 275.4000 333.3000 276.6000 340.2000 ;
	    RECT 277.8000 333.3000 279.0000 339.3000 ;
	    RECT 292.2000 333.3000 293.4000 340.5000 ;
	    RECT 294.6000 339.4500 295.8000 339.6000 ;
	    RECT 306.6000 339.4500 307.8000 339.6000 ;
	    RECT 294.6000 338.5500 307.8000 339.4500 ;
	    RECT 294.6000 338.4000 295.8000 338.5500 ;
	    RECT 306.6000 338.4000 307.8000 338.5500 ;
	    RECT 294.6000 337.2000 295.8000 337.5000 ;
	    RECT 294.6000 333.3000 295.8000 336.3000 ;
	    RECT 313.8000 333.3000 315.0000 340.5000 ;
	    RECT 316.5000 340.2000 319.8000 341.1000 ;
	    RECT 337.8000 340.2000 339.0000 340.5000 ;
	    RECT 316.2000 333.3000 317.4000 339.3000 ;
	    RECT 318.6000 333.3000 319.8000 340.2000 ;
	    RECT 340.2000 339.3000 341.4000 343.5000 ;
	    RECT 386.4000 342.6000 387.3000 347.7000 ;
	    RECT 412.2000 346.5000 413.4000 359.7000 ;
	    RECT 414.6000 353.7000 415.8000 359.7000 ;
	    RECT 441.0000 353.7000 442.2000 359.7000 ;
	    RECT 414.6000 349.5000 415.8000 349.8000 ;
	    RECT 414.6000 348.4500 415.8000 348.6000 ;
	    RECT 417.0000 348.4500 418.2000 348.6000 ;
	    RECT 414.6000 347.5500 418.2000 348.4500 ;
	    RECT 414.6000 347.4000 415.8000 347.5500 ;
	    RECT 417.0000 347.4000 418.2000 347.5500 ;
	    RECT 443.4000 346.5000 444.6000 359.7000 ;
	    RECT 445.8000 353.7000 447.0000 359.7000 ;
	    RECT 470.7000 353.7000 471.9000 359.7000 ;
	    RECT 471.0000 350.4000 472.2000 351.6000 ;
	    RECT 445.8000 349.5000 447.0000 349.8000 ;
	    RECT 471.0000 349.5000 471.9000 350.4000 ;
	    RECT 473.1000 348.6000 474.3000 359.7000 ;
	    RECT 445.8000 348.4500 447.0000 348.6000 ;
	    RECT 448.2000 348.4500 449.4000 348.6000 ;
	    RECT 445.8000 347.5500 449.4000 348.4500 ;
	    RECT 445.8000 347.4000 447.0000 347.5500 ;
	    RECT 448.2000 347.4000 449.4000 347.5500 ;
	    RECT 469.8000 347.4000 471.0000 348.6000 ;
	    RECT 472.8000 347.7000 474.3000 348.6000 ;
	    RECT 477.0000 347.7000 478.2000 359.7000 ;
	    RECT 601.8000 353.7000 603.0000 359.7000 ;
	    RECT 604.2000 352.5000 605.4000 359.7000 ;
	    RECT 606.6000 353.7000 607.8000 359.7000 ;
	    RECT 609.0000 352.8000 610.2000 359.7000 ;
	    RECT 611.4000 353.7000 612.6000 359.7000 ;
	    RECT 606.3000 351.9000 610.2000 352.8000 ;
	    RECT 537.0000 351.4500 538.2000 351.6000 ;
	    RECT 544.2000 351.4500 545.4000 351.6000 ;
	    RECT 604.2000 351.4500 605.4000 351.6000 ;
	    RECT 537.0000 350.5500 605.4000 351.4500 ;
	    RECT 537.0000 350.4000 538.2000 350.5500 ;
	    RECT 544.2000 350.4000 545.4000 350.5500 ;
	    RECT 604.2000 350.4000 605.4000 350.5500 ;
	    RECT 606.3000 349.5000 607.2000 351.9000 ;
	    RECT 613.8000 351.6000 615.0000 359.7000 ;
	    RECT 616.2000 353.7000 617.4000 359.7000 ;
	    RECT 618.6000 355.5000 619.8000 359.7000 ;
	    RECT 621.0000 355.5000 622.2000 359.7000 ;
	    RECT 623.4000 355.5000 624.6000 359.7000 ;
	    RECT 615.9000 351.6000 622.2000 352.8000 ;
	    RECT 611.1000 350.4000 615.0000 351.6000 ;
	    RECT 625.8000 350.4000 627.0000 359.7000 ;
	    RECT 628.2000 353.7000 629.4000 359.7000 ;
	    RECT 630.6000 352.5000 631.8000 359.7000 ;
	    RECT 633.0000 353.7000 634.2000 359.7000 ;
	    RECT 635.4000 352.5000 636.6000 359.7000 ;
	    RECT 637.8000 355.5000 639.0000 359.7000 ;
	    RECT 640.2000 355.5000 641.4000 359.7000 ;
	    RECT 642.6000 353.7000 643.8000 359.7000 ;
	    RECT 645.0000 352.8000 646.2000 359.7000 ;
	    RECT 647.4000 353.7000 648.6000 360.6000 ;
	    RECT 649.8000 354.6000 651.0000 359.7000 ;
	    RECT 649.8000 353.7000 651.3000 354.6000 ;
	    RECT 652.2000 353.7000 653.4000 359.7000 ;
	    RECT 678.6000 353.7000 679.8000 359.7000 ;
	    RECT 650.4000 352.8000 651.3000 353.7000 ;
	    RECT 643.2000 351.6000 649.5000 352.8000 ;
	    RECT 650.4000 351.9000 653.4000 352.8000 ;
	    RECT 630.6000 350.4000 634.5000 351.6000 ;
	    RECT 635.4000 350.7000 644.1000 351.6000 ;
	    RECT 648.6000 351.0000 649.5000 351.6000 ;
	    RECT 618.6000 349.5000 619.8000 349.8000 ;
	    RECT 604.2000 348.0000 605.4000 349.5000 ;
	    RECT 388.2000 344.4000 389.4000 345.6000 ;
	    RECT 390.6000 345.4500 391.8000 345.6000 ;
	    RECT 412.2000 345.4500 413.4000 345.6000 ;
	    RECT 390.6000 344.5500 413.4000 345.4500 ;
	    RECT 390.6000 344.4000 391.8000 344.5500 ;
	    RECT 412.2000 344.4000 413.4000 344.5500 ;
	    RECT 443.4000 345.4500 444.6000 345.6000 ;
	    RECT 469.9500 345.4500 470.8500 347.4000 ;
	    RECT 443.4000 344.5500 470.8500 345.4500 ;
	    RECT 443.4000 344.4000 444.6000 344.5500 ;
	    RECT 388.2000 343.2000 389.4000 343.5000 ;
	    RECT 359.4000 342.4500 360.6000 342.6000 ;
	    RECT 381.0000 342.4500 382.2000 342.6000 ;
	    RECT 359.4000 341.5500 382.2000 342.4500 ;
	    RECT 359.4000 341.4000 360.6000 341.5500 ;
	    RECT 381.0000 341.4000 382.2000 341.5500 ;
	    RECT 383.4000 341.4000 384.6000 342.6000 ;
	    RECT 385.5000 341.4000 387.3000 342.6000 ;
	    RECT 390.6000 342.4500 391.8000 342.6000 ;
	    RECT 405.0000 342.4500 406.2000 342.6000 ;
	    RECT 389.4000 340.8000 389.7000 342.3000 ;
	    RECT 390.6000 341.5500 406.2000 342.4500 ;
	    RECT 390.6000 341.4000 391.8000 341.5500 ;
	    RECT 405.0000 341.4000 406.2000 341.5500 ;
	    RECT 409.8000 341.4000 411.0000 342.6000 ;
	    RECT 337.8000 333.3000 339.0000 339.3000 ;
	    RECT 340.2000 338.4000 342.9000 339.3000 ;
	    RECT 357.0000 338.4000 358.2000 339.6000 ;
	    RECT 341.7000 333.3000 342.9000 338.4000 ;
	    RECT 357.0000 337.2000 358.2000 337.5000 ;
	    RECT 357.0000 333.3000 358.2000 336.3000 ;
	    RECT 359.4000 333.3000 360.6000 340.5000 ;
	    RECT 383.7000 339.3000 384.6000 340.5000 ;
	    RECT 409.8000 340.2000 411.0000 340.5000 ;
	    RECT 386.1000 339.3000 391.5000 339.9000 ;
	    RECT 412.2000 339.3000 413.4000 343.5000 ;
	    RECT 441.0000 341.4000 442.2000 342.6000 ;
	    RECT 441.0000 340.2000 442.2000 340.5000 ;
	    RECT 443.4000 339.3000 444.6000 343.5000 ;
	    RECT 472.8000 342.6000 473.7000 347.7000 ;
	    RECT 603.9000 346.8000 605.4000 348.0000 ;
	    RECT 606.3000 348.6000 619.8000 349.5000 ;
	    RECT 623.4000 349.5000 624.6000 349.8000 ;
	    RECT 635.4000 349.5000 636.3000 350.7000 ;
	    RECT 645.0000 349.8000 647.1000 350.7000 ;
	    RECT 648.6000 349.8000 651.0000 351.0000 ;
	    RECT 623.4000 348.6000 636.3000 349.5000 ;
	    RECT 637.8000 349.5000 647.1000 349.8000 ;
	    RECT 637.8000 348.9000 645.9000 349.5000 ;
	    RECT 637.8000 348.6000 639.0000 348.9000 ;
	    RECT 474.6000 344.4000 475.8000 345.6000 ;
	    RECT 474.6000 343.2000 475.8000 343.5000 ;
	    RECT 469.8000 341.4000 471.0000 342.6000 ;
	    RECT 471.9000 341.4000 473.7000 342.6000 ;
	    RECT 477.0000 342.4500 478.2000 342.6000 ;
	    RECT 501.0000 342.4500 502.2000 342.6000 ;
	    RECT 475.8000 340.8000 476.1000 342.3000 ;
	    RECT 477.0000 341.5500 502.2000 342.4500 ;
	    RECT 477.0000 341.4000 478.2000 341.5500 ;
	    RECT 501.0000 341.4000 502.2000 341.5500 ;
	    RECT 470.1000 339.3000 471.0000 340.5000 ;
	    RECT 603.9000 340.2000 605.1000 346.8000 ;
	    RECT 606.3000 345.9000 607.2000 348.6000 ;
	    RECT 642.3000 347.7000 643.5000 348.0000 ;
	    RECT 608.1000 346.8000 646.5000 347.7000 ;
	    RECT 647.4000 347.4000 648.6000 348.6000 ;
	    RECT 608.1000 346.5000 609.3000 346.8000 ;
	    RECT 606.0000 345.0000 607.2000 345.9000 ;
	    RECT 616.2000 345.0000 641.7000 345.9000 ;
	    RECT 606.0000 342.0000 606.9000 345.0000 ;
	    RECT 616.2000 344.1000 617.4000 345.0000 ;
	    RECT 642.6000 344.4000 643.8000 345.6000 ;
	    RECT 644.7000 345.0000 651.3000 345.9000 ;
	    RECT 650.1000 344.7000 651.3000 345.0000 ;
	    RECT 607.8000 342.9000 613.5000 344.1000 ;
	    RECT 606.0000 341.1000 607.8000 342.0000 ;
	    RECT 472.5000 339.3000 477.9000 339.9000 ;
	    RECT 383.4000 333.3000 384.6000 339.3000 ;
	    RECT 385.8000 339.0000 391.8000 339.3000 ;
	    RECT 385.8000 333.3000 387.0000 339.0000 ;
	    RECT 388.2000 333.3000 389.4000 338.1000 ;
	    RECT 390.6000 333.3000 391.8000 339.0000 ;
	    RECT 409.8000 333.3000 411.0000 339.3000 ;
	    RECT 412.2000 338.4000 414.9000 339.3000 ;
	    RECT 413.7000 333.3000 414.9000 338.4000 ;
	    RECT 441.0000 333.3000 442.2000 339.3000 ;
	    RECT 443.4000 338.4000 446.1000 339.3000 ;
	    RECT 444.9000 333.3000 446.1000 338.4000 ;
	    RECT 469.8000 333.3000 471.0000 339.3000 ;
	    RECT 472.2000 339.0000 478.2000 339.3000 ;
	    RECT 603.9000 339.0000 605.4000 340.2000 ;
	    RECT 472.2000 333.3000 473.4000 339.0000 ;
	    RECT 474.6000 333.3000 475.8000 338.1000 ;
	    RECT 477.0000 333.3000 478.2000 339.0000 ;
	    RECT 601.8000 333.3000 603.0000 336.3000 ;
	    RECT 604.2000 333.3000 605.4000 339.0000 ;
	    RECT 606.6000 333.3000 607.8000 341.1000 ;
	    RECT 612.3000 341.1000 613.5000 342.9000 ;
	    RECT 612.3000 340.2000 615.0000 341.1000 ;
	    RECT 613.8000 339.3000 615.0000 340.2000 ;
	    RECT 621.0000 339.6000 622.2000 343.8000 ;
	    RECT 625.8000 342.9000 630.6000 344.1000 ;
	    RECT 636.3000 342.9000 639.3000 344.1000 ;
	    RECT 652.2000 343.5000 653.4000 351.9000 ;
	    RECT 681.0000 346.5000 682.2000 359.7000 ;
	    RECT 683.4000 353.7000 684.6000 359.7000 ;
	    RECT 774.6000 354.4500 775.8000 354.6000 ;
	    RECT 805.8000 354.4500 807.0000 354.6000 ;
	    RECT 774.6000 353.5500 807.0000 354.4500 ;
	    RECT 808.2000 353.7000 809.4000 359.7000 ;
	    RECT 810.6000 354.6000 811.8000 359.7000 ;
	    RECT 810.3000 353.7000 811.8000 354.6000 ;
	    RECT 813.0000 353.7000 814.2000 360.6000 ;
	    RECT 774.6000 353.4000 775.8000 353.5500 ;
	    RECT 805.8000 353.4000 807.0000 353.5500 ;
	    RECT 810.3000 352.8000 811.2000 353.7000 ;
	    RECT 815.4000 352.8000 816.6000 359.7000 ;
	    RECT 817.8000 353.7000 819.0000 359.7000 ;
	    RECT 820.2000 355.5000 821.4000 359.7000 ;
	    RECT 822.6000 355.5000 823.8000 359.7000 ;
	    RECT 808.2000 351.9000 811.2000 352.8000 ;
	    RECT 683.4000 349.5000 684.6000 349.8000 ;
	    RECT 683.4000 348.4500 684.6000 348.6000 ;
	    RECT 690.6000 348.4500 691.8000 348.6000 ;
	    RECT 683.4000 347.5500 691.8000 348.4500 ;
	    RECT 683.4000 347.4000 684.6000 347.5500 ;
	    RECT 690.6000 347.4000 691.8000 347.5500 ;
	    RECT 659.4000 345.4500 660.6000 345.6000 ;
	    RECT 681.0000 345.4500 682.2000 345.6000 ;
	    RECT 659.4000 344.5500 682.2000 345.4500 ;
	    RECT 659.4000 344.4000 660.6000 344.5500 ;
	    RECT 681.0000 344.4000 682.2000 344.5500 ;
	    RECT 808.2000 343.5000 809.4000 351.9000 ;
	    RECT 812.1000 351.6000 818.4000 352.8000 ;
	    RECT 825.0000 352.5000 826.2000 359.7000 ;
	    RECT 827.4000 353.7000 828.6000 359.7000 ;
	    RECT 829.8000 352.5000 831.0000 359.7000 ;
	    RECT 832.2000 353.7000 833.4000 359.7000 ;
	    RECT 812.1000 351.0000 813.0000 351.6000 ;
	    RECT 810.6000 349.8000 813.0000 351.0000 ;
	    RECT 817.5000 350.7000 826.2000 351.6000 ;
	    RECT 814.5000 349.8000 816.6000 350.7000 ;
	    RECT 814.5000 349.5000 823.8000 349.8000 ;
	    RECT 815.7000 348.9000 823.8000 349.5000 ;
	    RECT 822.6000 348.6000 823.8000 348.9000 ;
	    RECT 825.3000 349.5000 826.2000 350.7000 ;
	    RECT 827.1000 350.4000 831.0000 351.6000 ;
	    RECT 834.6000 350.4000 835.8000 359.7000 ;
	    RECT 837.0000 355.5000 838.2000 359.7000 ;
	    RECT 839.4000 355.5000 840.6000 359.7000 ;
	    RECT 841.8000 355.5000 843.0000 359.7000 ;
	    RECT 844.2000 353.7000 845.4000 359.7000 ;
	    RECT 839.4000 351.6000 845.7000 352.8000 ;
	    RECT 846.6000 351.6000 847.8000 359.7000 ;
	    RECT 849.0000 353.7000 850.2000 359.7000 ;
	    RECT 851.4000 352.8000 852.6000 359.7000 ;
	    RECT 853.8000 353.7000 855.0000 359.7000 ;
	    RECT 851.4000 351.9000 855.3000 352.8000 ;
	    RECT 856.2000 352.5000 857.4000 359.7000 ;
	    RECT 858.6000 353.7000 859.8000 359.7000 ;
	    RECT 877.8000 353.7000 879.0000 359.7000 ;
	    RECT 846.6000 350.4000 850.5000 351.6000 ;
	    RECT 837.0000 349.5000 838.2000 349.8000 ;
	    RECT 825.3000 348.6000 838.2000 349.5000 ;
	    RECT 841.8000 349.5000 843.0000 349.8000 ;
	    RECT 854.4000 349.5000 855.3000 351.9000 ;
	    RECT 856.2000 350.4000 857.4000 351.6000 ;
	    RECT 841.8000 348.6000 855.3000 349.5000 ;
	    RECT 813.0000 347.4000 814.2000 348.6000 ;
	    RECT 818.1000 347.7000 819.3000 348.0000 ;
	    RECT 815.1000 346.8000 853.5000 347.7000 ;
	    RECT 852.3000 346.5000 853.5000 346.8000 ;
	    RECT 854.4000 345.9000 855.3000 348.6000 ;
	    RECT 856.2000 348.0000 857.4000 349.5000 ;
	    RECT 856.2000 346.8000 857.7000 348.0000 ;
	    RECT 810.3000 345.0000 816.9000 345.9000 ;
	    RECT 810.3000 344.7000 811.5000 345.0000 ;
	    RECT 817.8000 344.4000 819.0000 345.6000 ;
	    RECT 819.9000 345.0000 845.4000 345.9000 ;
	    RECT 854.4000 345.0000 855.6000 345.9000 ;
	    RECT 844.2000 344.1000 845.4000 345.0000 ;
	    RECT 625.2000 341.7000 626.4000 342.0000 ;
	    RECT 625.2000 340.8000 631.8000 341.7000 ;
	    RECT 633.0000 341.4000 634.2000 342.6000 ;
	    RECT 630.6000 340.5000 631.8000 340.8000 ;
	    RECT 633.0000 340.2000 634.2000 340.5000 ;
	    RECT 611.4000 333.3000 612.6000 339.3000 ;
	    RECT 613.8000 338.1000 617.4000 339.3000 ;
	    RECT 621.0000 338.4000 622.5000 339.6000 ;
	    RECT 627.0000 338.4000 627.3000 339.6000 ;
	    RECT 628.2000 338.4000 629.4000 339.6000 ;
	    RECT 630.6000 339.3000 631.8000 339.6000 ;
	    RECT 636.3000 339.3000 637.5000 342.9000 ;
	    RECT 640.2000 342.3000 653.4000 343.5000 ;
	    RECT 645.3000 340.2000 649.8000 341.4000 ;
	    RECT 645.3000 339.3000 646.5000 340.2000 ;
	    RECT 630.6000 338.4000 637.5000 339.3000 ;
	    RECT 616.2000 333.3000 617.4000 338.1000 ;
	    RECT 642.6000 338.1000 646.5000 339.3000 ;
	    RECT 618.6000 333.3000 619.8000 337.5000 ;
	    RECT 621.0000 333.3000 622.2000 337.5000 ;
	    RECT 623.4000 333.3000 624.6000 337.5000 ;
	    RECT 625.8000 333.3000 627.0000 337.5000 ;
	    RECT 628.2000 333.3000 629.4000 336.3000 ;
	    RECT 630.6000 333.3000 631.8000 337.5000 ;
	    RECT 633.0000 333.3000 634.2000 336.3000 ;
	    RECT 635.4000 333.3000 636.6000 337.5000 ;
	    RECT 637.8000 333.3000 639.0000 337.5000 ;
	    RECT 640.2000 333.3000 641.4000 337.5000 ;
	    RECT 642.6000 333.3000 643.8000 338.1000 ;
	    RECT 647.4000 333.3000 648.6000 339.3000 ;
	    RECT 652.2000 333.3000 653.4000 342.3000 ;
	    RECT 654.6000 342.4500 655.8000 342.6000 ;
	    RECT 678.6000 342.4500 679.8000 342.6000 ;
	    RECT 654.6000 341.5500 679.8000 342.4500 ;
	    RECT 654.6000 341.4000 655.8000 341.5500 ;
	    RECT 678.6000 341.4000 679.8000 341.5500 ;
	    RECT 678.6000 340.2000 679.8000 340.5000 ;
	    RECT 681.0000 339.3000 682.2000 343.5000 ;
	    RECT 808.2000 342.3000 821.4000 343.5000 ;
	    RECT 822.3000 342.9000 825.3000 344.1000 ;
	    RECT 831.0000 342.9000 835.8000 344.1000 ;
	    RECT 678.6000 333.3000 679.8000 339.3000 ;
	    RECT 681.0000 338.4000 683.7000 339.3000 ;
	    RECT 682.5000 333.3000 683.7000 338.4000 ;
	    RECT 808.2000 333.3000 809.4000 342.3000 ;
	    RECT 811.8000 340.2000 816.3000 341.4000 ;
	    RECT 815.1000 339.3000 816.3000 340.2000 ;
	    RECT 824.1000 339.3000 825.3000 342.9000 ;
	    RECT 827.4000 341.4000 828.6000 342.6000 ;
	    RECT 835.2000 341.7000 836.4000 342.0000 ;
	    RECT 829.8000 340.8000 836.4000 341.7000 ;
	    RECT 829.8000 340.5000 831.0000 340.8000 ;
	    RECT 827.4000 340.2000 828.6000 340.5000 ;
	    RECT 839.4000 339.6000 840.6000 343.8000 ;
	    RECT 848.1000 342.9000 853.8000 344.1000 ;
	    RECT 848.1000 341.1000 849.3000 342.9000 ;
	    RECT 854.7000 342.0000 855.6000 345.0000 ;
	    RECT 829.8000 339.3000 831.0000 339.6000 ;
	    RECT 813.0000 333.3000 814.2000 339.3000 ;
	    RECT 815.1000 338.1000 819.0000 339.3000 ;
	    RECT 824.1000 338.4000 831.0000 339.3000 ;
	    RECT 832.2000 338.4000 833.4000 339.6000 ;
	    RECT 834.3000 338.4000 834.6000 339.6000 ;
	    RECT 839.1000 338.4000 840.6000 339.6000 ;
	    RECT 846.6000 340.2000 849.3000 341.1000 ;
	    RECT 853.8000 341.1000 855.6000 342.0000 ;
	    RECT 846.6000 339.3000 847.8000 340.2000 ;
	    RECT 817.8000 333.3000 819.0000 338.1000 ;
	    RECT 844.2000 338.1000 847.8000 339.3000 ;
	    RECT 820.2000 333.3000 821.4000 337.5000 ;
	    RECT 822.6000 333.3000 823.8000 337.5000 ;
	    RECT 825.0000 333.3000 826.2000 337.5000 ;
	    RECT 827.4000 333.3000 828.6000 336.3000 ;
	    RECT 829.8000 333.3000 831.0000 337.5000 ;
	    RECT 832.2000 333.3000 833.4000 336.3000 ;
	    RECT 834.6000 333.3000 835.8000 337.5000 ;
	    RECT 837.0000 333.3000 838.2000 337.5000 ;
	    RECT 839.4000 333.3000 840.6000 337.5000 ;
	    RECT 841.8000 333.3000 843.0000 337.5000 ;
	    RECT 844.2000 333.3000 845.4000 338.1000 ;
	    RECT 849.0000 333.3000 850.2000 339.3000 ;
	    RECT 853.8000 333.3000 855.0000 341.1000 ;
	    RECT 856.5000 340.2000 857.7000 346.8000 ;
	    RECT 880.2000 346.5000 881.4000 359.7000 ;
	    RECT 882.6000 353.7000 883.8000 359.7000 ;
	    RECT 1014.6000 353.7000 1015.8000 359.7000 ;
	    RECT 1017.0000 354.6000 1018.2000 359.7000 ;
	    RECT 1016.7000 353.7000 1018.2000 354.6000 ;
	    RECT 1019.4000 353.7000 1020.6000 360.6000 ;
	    RECT 1016.7000 352.8000 1017.6000 353.7000 ;
	    RECT 1021.8000 352.8000 1023.0000 359.7000 ;
	    RECT 1024.2001 353.7000 1025.4000 359.7000 ;
	    RECT 1026.6000 355.5000 1027.8000 359.7000 ;
	    RECT 1029.0000 355.5000 1030.2001 359.7000 ;
	    RECT 1014.6000 351.9000 1017.6000 352.8000 ;
	    RECT 882.6000 349.5000 883.8000 349.8000 ;
	    RECT 882.6000 348.4500 883.8000 348.6000 ;
	    RECT 921.0000 348.4500 922.2000 348.6000 ;
	    RECT 882.6000 347.5500 922.2000 348.4500 ;
	    RECT 882.6000 347.4000 883.8000 347.5500 ;
	    RECT 921.0000 347.4000 922.2000 347.5500 ;
	    RECT 861.0000 345.4500 862.2000 345.6000 ;
	    RECT 880.2000 345.4500 881.4000 345.6000 ;
	    RECT 861.0000 344.5500 881.4000 345.4500 ;
	    RECT 861.0000 344.4000 862.2000 344.5500 ;
	    RECT 880.2000 344.4000 881.4000 344.5500 ;
	    RECT 1014.6000 343.5000 1015.8000 351.9000 ;
	    RECT 1018.5000 351.6000 1024.8000 352.8000 ;
	    RECT 1031.4000 352.5000 1032.6000 359.7000 ;
	    RECT 1033.8000 353.7000 1035.0000 359.7000 ;
	    RECT 1036.2001 352.5000 1037.4000 359.7000 ;
	    RECT 1038.6000 353.7000 1039.8000 359.7000 ;
	    RECT 1018.5000 351.0000 1019.4000 351.6000 ;
	    RECT 1017.0000 349.8000 1019.4000 351.0000 ;
	    RECT 1023.9000 350.7000 1032.6000 351.6000 ;
	    RECT 1020.9000 349.8000 1023.0000 350.7000 ;
	    RECT 1020.9000 349.5000 1030.2001 349.8000 ;
	    RECT 1022.1000 348.9000 1030.2001 349.5000 ;
	    RECT 1029.0000 348.6000 1030.2001 348.9000 ;
	    RECT 1031.7001 349.5000 1032.6000 350.7000 ;
	    RECT 1033.5000 350.4000 1037.4000 351.6000 ;
	    RECT 1041.0000 350.4000 1042.2001 359.7000 ;
	    RECT 1043.4000 355.5000 1044.6000 359.7000 ;
	    RECT 1045.8000 355.5000 1047.0000 359.7000 ;
	    RECT 1048.2001 355.5000 1049.4000 359.7000 ;
	    RECT 1050.6000 353.7000 1051.8000 359.7000 ;
	    RECT 1045.8000 351.6000 1052.1000 352.8000 ;
	    RECT 1053.0000 351.6000 1054.2001 359.7000 ;
	    RECT 1055.4000 353.7000 1056.6000 359.7000 ;
	    RECT 1057.8000 352.8000 1059.0000 359.7000 ;
	    RECT 1060.2001 353.7000 1061.4000 359.7000 ;
	    RECT 1057.8000 351.9000 1061.7001 352.8000 ;
	    RECT 1062.6000 352.5000 1063.8000 359.7000 ;
	    RECT 1065.0000 353.7000 1066.2001 359.7000 ;
	    RECT 1089.0000 353.7000 1090.2001 359.7000 ;
	    RECT 1091.4000 354.3000 1092.6000 359.7000 ;
	    RECT 1089.3000 353.4000 1090.2001 353.7000 ;
	    RECT 1093.8000 353.7000 1095.0000 359.7000 ;
	    RECT 1096.2001 353.7000 1097.4000 359.7000 ;
	    RECT 1115.4000 353.7000 1116.6000 359.7000 ;
	    RECT 1093.8000 353.4000 1094.7001 353.7000 ;
	    RECT 1089.3000 352.5000 1094.7001 353.4000 ;
	    RECT 1053.0000 350.4000 1056.9000 351.6000 ;
	    RECT 1043.4000 349.5000 1044.6000 349.8000 ;
	    RECT 1031.7001 348.6000 1044.6000 349.5000 ;
	    RECT 1048.2001 349.5000 1049.4000 349.8000 ;
	    RECT 1060.8000 349.5000 1061.7001 351.9000 ;
	    RECT 1062.6000 350.4000 1063.8000 351.6000 ;
	    RECT 1089.3000 349.5000 1090.2001 352.5000 ;
	    RECT 1091.4000 351.4500 1092.6000 351.6000 ;
	    RECT 1098.6000 351.4500 1099.8000 351.6000 ;
	    RECT 1091.4000 350.5500 1099.8000 351.4500 ;
	    RECT 1091.4000 350.4000 1092.6000 350.5500 ;
	    RECT 1098.6000 350.4000 1099.8000 350.5500 ;
	    RECT 1115.4000 349.5000 1116.6000 349.8000 ;
	    RECT 1048.2001 348.6000 1061.7001 349.5000 ;
	    RECT 1019.4000 347.4000 1020.6000 348.6000 ;
	    RECT 1024.5000 347.7000 1025.7001 348.0000 ;
	    RECT 1021.5000 346.8000 1059.9000 347.7000 ;
	    RECT 1058.7001 346.5000 1059.9000 346.8000 ;
	    RECT 1060.8000 345.9000 1061.7001 348.6000 ;
	    RECT 1062.6000 348.0000 1063.8000 349.5000 ;
	    RECT 1091.4000 349.2000 1092.6000 349.5000 ;
	    RECT 1084.2001 348.4500 1085.4000 348.6000 ;
	    RECT 1089.0000 348.4500 1090.2001 348.6000 ;
	    RECT 1062.6000 346.8000 1064.1000 348.0000 ;
	    RECT 1084.2001 347.5500 1090.2001 348.4500 ;
	    RECT 1084.2001 347.4000 1085.4000 347.5500 ;
	    RECT 1089.0000 347.4000 1090.2001 347.5500 ;
	    RECT 1096.2001 348.4500 1097.4000 348.6000 ;
	    RECT 1101.0000 348.4500 1102.2001 348.6000 ;
	    RECT 1096.2001 347.5500 1102.2001 348.4500 ;
	    RECT 1096.2001 347.4000 1097.4000 347.5500 ;
	    RECT 1101.0000 347.4000 1102.2001 347.5500 ;
	    RECT 1115.4000 347.4000 1116.6000 348.6000 ;
	    RECT 1016.7000 345.0000 1023.3000 345.9000 ;
	    RECT 1016.7000 344.7000 1017.9000 345.0000 ;
	    RECT 1024.2001 344.4000 1025.4000 345.6000 ;
	    RECT 1026.3000 345.0000 1051.8000 345.9000 ;
	    RECT 1060.8000 345.0000 1062.0000 345.9000 ;
	    RECT 1050.6000 344.1000 1051.8000 345.0000 ;
	    RECT 858.6000 342.4500 859.8000 342.6000 ;
	    RECT 875.4000 342.4500 876.6000 342.6000 ;
	    RECT 877.8000 342.4500 879.0000 342.6000 ;
	    RECT 858.6000 341.5500 879.0000 342.4500 ;
	    RECT 858.6000 341.4000 859.8000 341.5500 ;
	    RECT 875.4000 341.4000 876.6000 341.5500 ;
	    RECT 877.8000 341.4000 879.0000 341.5500 ;
	    RECT 877.8000 340.2000 879.0000 340.5000 ;
	    RECT 856.2000 339.0000 857.7000 340.2000 ;
	    RECT 880.2000 339.3000 881.4000 343.5000 ;
	    RECT 1014.6000 342.3000 1027.8000 343.5000 ;
	    RECT 1028.7001 342.9000 1031.7001 344.1000 ;
	    RECT 1037.4000 342.9000 1042.2001 344.1000 ;
	    RECT 856.2000 333.3000 857.4000 339.0000 ;
	    RECT 858.6000 333.3000 859.8000 336.3000 ;
	    RECT 877.8000 333.3000 879.0000 339.3000 ;
	    RECT 880.2000 338.4000 882.9000 339.3000 ;
	    RECT 881.7000 333.3000 882.9000 338.4000 ;
	    RECT 1014.6000 333.3000 1015.8000 342.3000 ;
	    RECT 1018.2000 340.2000 1022.7000 341.4000 ;
	    RECT 1021.5000 339.3000 1022.7000 340.2000 ;
	    RECT 1030.5000 339.3000 1031.7001 342.9000 ;
	    RECT 1033.8000 341.4000 1035.0000 342.6000 ;
	    RECT 1041.6000 341.7000 1042.8000 342.0000 ;
	    RECT 1036.2001 340.8000 1042.8000 341.7000 ;
	    RECT 1036.2001 340.5000 1037.4000 340.8000 ;
	    RECT 1033.8000 340.2000 1035.0000 340.5000 ;
	    RECT 1045.8000 339.6000 1047.0000 343.8000 ;
	    RECT 1054.5000 342.9000 1060.2001 344.1000 ;
	    RECT 1054.5000 341.1000 1055.7001 342.9000 ;
	    RECT 1061.1000 342.0000 1062.0000 345.0000 ;
	    RECT 1036.2001 339.3000 1037.4000 339.6000 ;
	    RECT 1019.4000 333.3000 1020.6000 339.3000 ;
	    RECT 1021.5000 338.1000 1025.4000 339.3000 ;
	    RECT 1030.5000 338.4000 1037.4000 339.3000 ;
	    RECT 1038.6000 338.4000 1039.8000 339.6000 ;
	    RECT 1040.7001 338.4000 1041.0000 339.6000 ;
	    RECT 1045.5000 338.4000 1047.0000 339.6000 ;
	    RECT 1053.0000 340.2000 1055.7001 341.1000 ;
	    RECT 1060.2001 341.1000 1062.0000 342.0000 ;
	    RECT 1053.0000 339.3000 1054.2001 340.2000 ;
	    RECT 1024.2001 333.3000 1025.4000 338.1000 ;
	    RECT 1050.6000 338.1000 1054.2001 339.3000 ;
	    RECT 1026.6000 333.3000 1027.8000 337.5000 ;
	    RECT 1029.0000 333.3000 1030.2001 337.5000 ;
	    RECT 1031.4000 333.3000 1032.6000 337.5000 ;
	    RECT 1033.8000 333.3000 1035.0000 336.3000 ;
	    RECT 1036.2001 333.3000 1037.4000 337.5000 ;
	    RECT 1038.6000 333.3000 1039.8000 336.3000 ;
	    RECT 1041.0000 333.3000 1042.2001 337.5000 ;
	    RECT 1043.4000 333.3000 1044.6000 337.5000 ;
	    RECT 1045.8000 333.3000 1047.0000 337.5000 ;
	    RECT 1048.2001 333.3000 1049.4000 337.5000 ;
	    RECT 1050.6000 333.3000 1051.8000 338.1000 ;
	    RECT 1055.4000 333.3000 1056.6000 339.3000 ;
	    RECT 1060.2001 333.3000 1061.4000 341.1000 ;
	    RECT 1062.9000 340.2000 1064.1000 346.8000 ;
	    RECT 1117.8000 346.5000 1119.0000 359.7000 ;
	    RECT 1120.2001 353.7000 1121.4000 359.7000 ;
	    RECT 1151.4000 353.7000 1152.6000 359.7000 ;
	    RECT 1153.8000 353.7000 1155.0000 359.7000 ;
	    RECT 1154.1000 347.4000 1155.0000 353.7000 ;
	    RECT 1156.2001 348.3000 1157.4000 359.7000 ;
	    RECT 1158.6000 347.7000 1159.8000 359.7000 ;
	    RECT 1154.1000 346.5000 1157.7001 347.4000 ;
	    RECT 1158.9000 346.5000 1159.8000 347.7000 ;
	    RECT 1089.3000 342.6000 1090.2001 346.5000 ;
	    RECT 1096.2001 346.2000 1097.4000 346.5000 ;
	    RECT 1092.6000 344.4000 1092.9000 345.6000 ;
	    RECT 1093.8000 344.4000 1095.0000 345.6000 ;
	    RECT 1098.6000 345.4500 1099.8000 345.6000 ;
	    RECT 1110.6000 345.4500 1111.8000 345.6000 ;
	    RECT 1117.8000 345.4500 1119.0000 345.6000 ;
	    RECT 1149.0000 345.4500 1150.2001 345.6000 ;
	    RECT 1098.6000 344.5500 1150.2001 345.4500 ;
	    RECT 1098.6000 344.4000 1099.8000 344.5500 ;
	    RECT 1110.6000 344.4000 1111.8000 344.5500 ;
	    RECT 1117.8000 344.4000 1119.0000 344.5500 ;
	    RECT 1149.0000 344.4000 1150.2001 344.5500 ;
	    RECT 1153.8000 344.4000 1155.0000 345.6000 ;
	    RECT 1151.4000 343.5000 1152.6000 343.8000 ;
	    RECT 1089.3000 342.3000 1091.7001 342.6000 ;
	    RECT 1089.3000 341.7000 1092.0000 342.3000 ;
	    RECT 1062.6000 339.0000 1064.1000 340.2000 ;
	    RECT 1062.6000 333.3000 1063.8000 339.0000 ;
	    RECT 1065.0000 333.3000 1066.2001 336.3000 ;
	    RECT 1090.8000 333.3000 1092.0000 341.7000 ;
	    RECT 1096.2001 333.3000 1097.4000 342.3000 ;
	    RECT 1117.8000 339.3000 1119.0000 343.5000 ;
	    RECT 1154.1000 343.2000 1155.0000 343.5000 ;
	    RECT 1120.2001 342.4500 1121.4000 342.6000 ;
	    RECT 1151.4000 342.4500 1152.6000 342.6000 ;
	    RECT 1120.2001 341.5500 1152.6000 342.4500 ;
	    RECT 1154.1000 342.3000 1155.6000 343.2000 ;
	    RECT 1154.4000 342.0000 1155.6000 342.3000 ;
	    RECT 1120.2001 341.4000 1121.4000 341.5500 ;
	    RECT 1151.4000 341.4000 1152.6000 341.5500 ;
	    RECT 1156.8000 341.4000 1157.7001 346.5000 ;
	    RECT 1158.6000 344.4000 1159.8000 345.6000 ;
	    RECT 1173.0000 343.5000 1174.2001 359.7000 ;
	    RECT 1175.4000 353.7000 1176.6000 359.7000 ;
	    RECT 1206.6000 358.8000 1212.6000 359.7000 ;
	    RECT 1206.6000 347.7000 1207.8000 358.8000 ;
	    RECT 1209.0000 347.7000 1210.2001 357.9000 ;
	    RECT 1211.4000 348.6000 1212.6000 358.8000 ;
	    RECT 1213.8000 349.5000 1215.0000 359.7000 ;
	    RECT 1216.2001 348.6000 1217.4000 359.7000 ;
	    RECT 1235.4000 353.7000 1236.6000 359.7000 ;
	    RECT 1211.4000 347.7000 1217.4000 348.6000 ;
	    RECT 1209.3000 346.8000 1210.2001 347.7000 ;
	    RECT 1206.6000 346.5000 1207.8000 346.8000 ;
	    RECT 1209.3000 346.5000 1212.3000 346.8000 ;
	    RECT 1237.8000 346.5000 1239.0000 359.7000 ;
	    RECT 1240.2001 353.7000 1241.4000 359.7000 ;
	    RECT 1259.4000 353.7000 1260.6000 359.7000 ;
	    RECT 1240.2001 349.5000 1241.4000 349.8000 ;
	    RECT 1259.4000 349.5000 1260.6000 349.8000 ;
	    RECT 1240.2001 347.4000 1241.4000 348.6000 ;
	    RECT 1247.4000 348.4500 1248.6000 348.6000 ;
	    RECT 1242.7500 347.5500 1248.6000 348.4500 ;
	    RECT 1209.3000 345.9000 1210.5000 346.5000 ;
	    RECT 1204.2001 345.4500 1205.4000 345.6000 ;
	    RECT 1206.6000 345.4500 1207.8000 345.6000 ;
	    RECT 1204.2001 344.5500 1207.8000 345.4500 ;
	    RECT 1204.2001 344.4000 1205.4000 344.5500 ;
	    RECT 1206.6000 344.4000 1207.8000 344.5500 ;
	    RECT 1211.4000 344.4000 1212.6000 345.6000 ;
	    RECT 1215.0000 344.7000 1215.3000 346.2000 ;
	    RECT 1216.2001 344.4000 1217.4000 345.6000 ;
	    RECT 1237.8000 345.4500 1239.0000 345.6000 ;
	    RECT 1242.7500 345.4500 1243.6500 347.5500 ;
	    RECT 1247.4000 347.4000 1248.6000 347.5500 ;
	    RECT 1259.4000 347.4000 1260.6000 348.6000 ;
	    RECT 1261.8000 346.5000 1263.0000 359.7000 ;
	    RECT 1264.2001 353.7000 1265.4000 359.7000 ;
	    RECT 1237.8000 344.5500 1243.6500 345.4500 ;
	    RECT 1245.0000 345.4500 1246.2001 345.6000 ;
	    RECT 1261.8000 345.4500 1263.0000 345.6000 ;
	    RECT 1273.8000 345.4500 1275.0000 345.6000 ;
	    RECT 1245.0000 344.5500 1275.0000 345.4500 ;
	    RECT 1237.8000 344.4000 1239.0000 344.5500 ;
	    RECT 1245.0000 344.4000 1246.2001 344.5500 ;
	    RECT 1261.8000 344.4000 1263.0000 344.5500 ;
	    RECT 1273.8000 344.4000 1275.0000 344.5500 ;
	    RECT 1209.3000 343.5000 1210.5000 344.4000 ;
	    RECT 1213.8000 343.5000 1215.0000 343.8000 ;
	    RECT 1156.8000 341.1000 1158.0000 341.4000 ;
	    RECT 1153.5000 340.5000 1158.0000 341.1000 ;
	    RECT 1120.2001 340.2000 1121.4000 340.5000 ;
	    RECT 1151.7001 340.2000 1158.0000 340.5000 ;
	    RECT 1151.7001 339.6000 1154.4000 340.2000 ;
	    RECT 1151.7001 339.3000 1152.6000 339.6000 ;
	    RECT 1158.9000 339.3000 1159.8000 343.5000 ;
	    RECT 1173.0000 342.4500 1174.2001 342.6000 ;
	    RECT 1182.6000 342.4500 1183.8000 342.6000 ;
	    RECT 1194.6000 342.4500 1195.8000 342.6000 ;
	    RECT 1173.0000 341.5500 1195.8000 342.4500 ;
	    RECT 1173.0000 341.4000 1174.2001 341.5500 ;
	    RECT 1182.6000 341.4000 1183.8000 341.5500 ;
	    RECT 1194.6000 341.4000 1195.8000 341.5500 ;
	    RECT 1209.0000 341.4000 1210.2001 342.6000 ;
	    RECT 1116.3000 338.4000 1119.0000 339.3000 ;
	    RECT 1116.3000 333.3000 1117.5000 338.4000 ;
	    RECT 1120.2001 333.3000 1121.4000 339.3000 ;
	    RECT 1151.4000 333.3000 1152.6000 339.3000 ;
	    RECT 1155.3000 333.3000 1156.5000 339.0000 ;
	    RECT 1157.7001 337.8000 1159.8000 339.3000 ;
	    RECT 1157.7001 333.3000 1158.9000 337.8000 ;
	    RECT 1173.0000 333.3000 1174.2001 340.5000 ;
	    RECT 1175.4000 338.4000 1176.6000 339.6000 ;
	    RECT 1211.4000 339.3000 1212.3000 343.5000 ;
	    RECT 1213.8000 341.4000 1215.0000 342.6000 ;
	    RECT 1216.3500 342.4500 1217.2500 344.4000 ;
	    RECT 1276.2001 343.5000 1277.4000 359.7000 ;
	    RECT 1278.6000 353.7000 1279.8000 359.7000 ;
	    RECT 1297.8000 353.7000 1299.0000 359.7000 ;
	    RECT 1297.8000 349.5000 1299.0000 349.8000 ;
	    RECT 1297.8000 347.4000 1299.0000 348.6000 ;
	    RECT 1300.2001 346.5000 1301.4000 359.7000 ;
	    RECT 1302.6000 353.7000 1303.8000 359.7000 ;
	    RECT 1329.9000 353.7000 1331.1000 359.7000 ;
	    RECT 1330.2001 350.4000 1331.4000 351.6000 ;
	    RECT 1330.2001 349.5000 1331.1000 350.4000 ;
	    RECT 1332.3000 348.6000 1333.5000 359.7000 ;
	    RECT 1321.8000 348.4500 1323.0000 348.6000 ;
	    RECT 1329.0000 348.4500 1330.2001 348.6000 ;
	    RECT 1321.8000 347.5500 1330.2001 348.4500 ;
	    RECT 1321.8000 347.4000 1323.0000 347.5500 ;
	    RECT 1329.0000 347.4000 1330.2001 347.5500 ;
	    RECT 1332.0000 347.7000 1333.5000 348.6000 ;
	    RECT 1336.2001 347.7000 1337.4000 359.7000 ;
	    RECT 1369.8000 348.6000 1371.0000 359.7000 ;
	    RECT 1372.2001 349.5000 1373.4000 359.7000 ;
	    RECT 1374.6000 348.6000 1375.8000 359.7000 ;
	    RECT 1369.8000 347.7000 1375.8000 348.6000 ;
	    RECT 1377.0000 347.7000 1378.2001 359.7000 ;
	    RECT 1401.9000 353.7000 1403.1000 359.7000 ;
	    RECT 1402.2001 350.4000 1403.4000 351.6000 ;
	    RECT 1402.2001 349.5000 1403.1000 350.4000 ;
	    RECT 1404.3000 348.6000 1405.5000 359.7000 ;
	    RECT 1391.4000 348.4500 1392.6000 348.6000 ;
	    RECT 1401.0000 348.4500 1402.2001 348.6000 ;
	    RECT 1281.0000 345.4500 1282.2001 345.6000 ;
	    RECT 1300.2001 345.4500 1301.4000 345.6000 ;
	    RECT 1281.0000 344.5500 1301.4000 345.4500 ;
	    RECT 1281.0000 344.4000 1282.2001 344.5500 ;
	    RECT 1300.2001 344.4000 1301.4000 344.5500 ;
	    RECT 1235.4000 342.4500 1236.6000 342.6000 ;
	    RECT 1216.3500 341.5500 1236.6000 342.4500 ;
	    RECT 1235.4000 341.4000 1236.6000 341.5500 ;
	    RECT 1235.4000 340.2000 1236.6000 340.5000 ;
	    RECT 1237.8000 339.3000 1239.0000 343.5000 ;
	    RECT 1261.8000 339.3000 1263.0000 343.5000 ;
	    RECT 1264.2001 341.4000 1265.4000 342.6000 ;
	    RECT 1276.2001 342.4500 1277.4000 342.6000 ;
	    RECT 1285.8000 342.4500 1287.0000 342.6000 ;
	    RECT 1276.2001 341.5500 1287.0000 342.4500 ;
	    RECT 1276.2001 341.4000 1277.4000 341.5500 ;
	    RECT 1285.8000 341.4000 1287.0000 341.5500 ;
	    RECT 1264.2001 340.2000 1265.4000 340.5000 ;
	    RECT 1175.4000 337.2000 1176.6000 337.5000 ;
	    RECT 1175.4000 333.3000 1176.6000 336.3000 ;
	    RECT 1206.6000 333.3000 1207.8000 339.3000 ;
	    RECT 1210.5000 333.3000 1212.9000 339.3000 ;
	    RECT 1215.6000 333.3000 1216.8000 339.3000 ;
	    RECT 1235.4000 333.3000 1236.6000 339.3000 ;
	    RECT 1237.8000 338.4000 1240.5000 339.3000 ;
	    RECT 1239.3000 333.3000 1240.5000 338.4000 ;
	    RECT 1260.3000 338.4000 1263.0000 339.3000 ;
	    RECT 1260.3000 333.3000 1261.5000 338.4000 ;
	    RECT 1264.2001 333.3000 1265.4000 339.3000 ;
	    RECT 1276.2001 333.3000 1277.4000 340.5000 ;
	    RECT 1278.6000 339.4500 1279.8000 339.6000 ;
	    RECT 1295.4000 339.4500 1296.6000 339.6000 ;
	    RECT 1278.6000 338.5500 1296.6000 339.4500 ;
	    RECT 1300.2001 339.3000 1301.4000 343.5000 ;
	    RECT 1332.0000 342.6000 1332.9000 347.7000 ;
	    RECT 1377.0000 346.5000 1377.9000 347.7000 ;
	    RECT 1391.4000 347.5500 1402.2001 348.4500 ;
	    RECT 1391.4000 347.4000 1392.6000 347.5500 ;
	    RECT 1401.0000 347.4000 1402.2001 347.5500 ;
	    RECT 1404.0000 347.7000 1405.5000 348.6000 ;
	    RECT 1408.2001 347.7000 1409.4000 359.7000 ;
	    RECT 1434.6000 348.6000 1435.8000 359.7000 ;
	    RECT 1437.0000 349.5000 1438.2001 359.7000 ;
	    RECT 1439.4000 348.6000 1440.6000 359.7000 ;
	    RECT 1434.6000 347.7000 1440.6000 348.6000 ;
	    RECT 1441.8000 347.7000 1443.0000 359.7000 ;
	    RECT 1468.2001 353.7000 1469.4000 359.7000 ;
	    RECT 1470.6000 354.3000 1471.8000 359.7000 ;
	    RECT 1468.5000 353.4000 1469.4000 353.7000 ;
	    RECT 1473.0000 353.7000 1474.2001 359.7000 ;
	    RECT 1475.4000 353.7000 1476.6000 359.7000 ;
	    RECT 1473.0000 353.4000 1473.9000 353.7000 ;
	    RECT 1468.5000 352.5000 1473.9000 353.4000 ;
	    RECT 1468.5000 349.5000 1469.4000 352.5000 ;
	    RECT 1470.6000 350.4000 1471.8000 351.6000 ;
	    RECT 1470.6000 349.2000 1471.8000 349.5000 ;
	    RECT 1518.6000 348.6000 1519.8000 359.7000 ;
	    RECT 1521.0000 349.8000 1522.5000 359.7000 ;
	    RECT 1521.3000 348.6000 1522.5000 348.9000 ;
	    RECT 1333.8000 344.4000 1335.0000 345.6000 ;
	    RECT 1348.2001 345.4500 1349.4000 345.6000 ;
	    RECT 1369.8000 345.4500 1371.0000 345.6000 ;
	    RECT 1348.2001 344.5500 1371.0000 345.4500 ;
	    RECT 1371.9000 344.7000 1372.2001 346.2000 ;
	    RECT 1374.6000 344.7000 1376.1000 345.6000 ;
	    RECT 1377.0000 345.4500 1378.2001 345.6000 ;
	    RECT 1393.8000 345.4500 1395.0000 345.6000 ;
	    RECT 1348.2001 344.4000 1349.4000 344.5500 ;
	    RECT 1369.8000 344.4000 1371.0000 344.5500 ;
	    RECT 1372.2001 343.5000 1373.4000 343.8000 ;
	    RECT 1333.8000 343.2000 1335.0000 343.5000 ;
	    RECT 1302.6000 342.4500 1303.8000 342.6000 ;
	    RECT 1314.6000 342.4500 1315.8000 342.6000 ;
	    RECT 1302.6000 341.5500 1315.8000 342.4500 ;
	    RECT 1302.6000 341.4000 1303.8000 341.5500 ;
	    RECT 1314.6000 341.4000 1315.8000 341.5500 ;
	    RECT 1324.2001 342.4500 1325.4000 342.6000 ;
	    RECT 1329.0000 342.4500 1330.2001 342.6000 ;
	    RECT 1324.2001 341.5500 1330.2001 342.4500 ;
	    RECT 1324.2001 341.4000 1325.4000 341.5500 ;
	    RECT 1329.0000 341.4000 1330.2001 341.5500 ;
	    RECT 1331.1000 341.4000 1332.9000 342.6000 ;
	    RECT 1335.0000 340.8000 1335.3000 342.3000 ;
	    RECT 1336.2001 341.4000 1337.4000 342.6000 ;
	    RECT 1343.4000 342.4500 1344.6000 342.6000 ;
	    RECT 1372.2001 342.4500 1373.4000 342.6000 ;
	    RECT 1343.4000 341.5500 1373.4000 342.4500 ;
	    RECT 1343.4000 341.4000 1344.6000 341.5500 ;
	    RECT 1372.2001 341.4000 1373.4000 341.5500 ;
	    RECT 1302.6000 340.2000 1303.8000 340.5000 ;
	    RECT 1329.3000 339.3000 1330.2001 340.5000 ;
	    RECT 1331.7001 339.3000 1337.1000 339.9000 ;
	    RECT 1374.6000 339.3000 1375.5000 344.7000 ;
	    RECT 1377.0000 344.5500 1395.0000 345.4500 ;
	    RECT 1377.0000 344.4000 1378.2001 344.5500 ;
	    RECT 1393.8000 344.4000 1395.0000 344.5500 ;
	    RECT 1404.0000 342.6000 1404.9000 347.7000 ;
	    RECT 1441.8000 346.5000 1442.7001 347.7000 ;
	    RECT 1468.2001 347.4000 1469.4000 348.6000 ;
	    RECT 1475.4000 348.4500 1476.6000 348.6000 ;
	    RECT 1485.0000 348.4500 1486.2001 348.6000 ;
	    RECT 1513.8000 348.4500 1515.0000 348.6000 ;
	    RECT 1475.4000 347.5500 1515.0000 348.4500 ;
	    RECT 1518.6000 347.7000 1522.5000 348.6000 ;
	    RECT 1525.2001 347.7000 1527.6000 359.7000 ;
	    RECT 1530.3000 349.8000 1531.8000 359.7000 ;
	    RECT 1530.6000 348.6000 1531.8000 348.9000 ;
	    RECT 1533.0000 348.6000 1534.2001 359.7000 ;
	    RECT 1559.4000 353.7000 1560.6000 359.7000 ;
	    RECT 1561.8000 353.7000 1563.0000 359.7000 ;
	    RECT 1564.2001 354.3000 1565.4000 359.7000 ;
	    RECT 1562.1000 353.4000 1563.0000 353.7000 ;
	    RECT 1566.6000 353.7000 1567.8000 359.7000 ;
	    RECT 1566.6000 353.4000 1567.5000 353.7000 ;
	    RECT 1562.1000 352.5000 1567.5000 353.4000 ;
	    RECT 1564.2001 350.4000 1565.4000 351.6000 ;
	    RECT 1566.6000 349.5000 1567.5000 352.5000 ;
	    RECT 1564.2001 349.2000 1565.4000 349.5000 ;
	    RECT 1530.6000 347.7000 1534.2001 348.6000 ;
	    RECT 1540.2001 348.4500 1541.4000 348.6000 ;
	    RECT 1559.4000 348.4500 1560.6000 348.6000 ;
	    RECT 1475.4000 347.4000 1476.6000 347.5500 ;
	    RECT 1485.0000 347.4000 1486.2001 347.5500 ;
	    RECT 1513.8000 347.4000 1515.0000 347.5500 ;
	    RECT 1526.1000 346.5000 1527.0000 347.7000 ;
	    RECT 1540.2001 347.5500 1560.6000 348.4500 ;
	    RECT 1540.2001 347.4000 1541.4000 347.5500 ;
	    RECT 1559.4000 347.4000 1560.6000 347.5500 ;
	    RECT 1566.6000 347.4000 1567.8000 348.6000 ;
	    RECT 1405.8000 344.4000 1407.0000 345.6000 ;
	    RECT 1427.4000 345.4500 1428.6000 345.6000 ;
	    RECT 1434.6000 345.4500 1435.8000 345.6000 ;
	    RECT 1427.4000 344.5500 1435.8000 345.4500 ;
	    RECT 1436.7001 344.7000 1437.0000 346.2000 ;
	    RECT 1439.4000 344.7000 1440.9000 345.6000 ;
	    RECT 1441.8000 345.4500 1443.0000 345.6000 ;
	    RECT 1451.4000 345.4500 1452.6000 345.6000 ;
	    RECT 1458.6000 345.4500 1459.8000 345.6000 ;
	    RECT 1427.4000 344.4000 1428.6000 344.5500 ;
	    RECT 1434.6000 344.4000 1435.8000 344.5500 ;
	    RECT 1437.0000 343.5000 1438.2001 343.8000 ;
	    RECT 1405.8000 343.2000 1407.0000 343.5000 ;
	    RECT 1389.0000 342.4500 1390.2001 342.6000 ;
	    RECT 1401.0000 342.4500 1402.2001 342.6000 ;
	    RECT 1389.0000 341.5500 1402.2001 342.4500 ;
	    RECT 1389.0000 341.4000 1390.2001 341.5500 ;
	    RECT 1401.0000 341.4000 1402.2001 341.5500 ;
	    RECT 1403.1000 341.4000 1404.9000 342.6000 ;
	    RECT 1407.0000 340.8000 1407.3000 342.3000 ;
	    RECT 1408.2001 341.4000 1409.4000 342.6000 ;
	    RECT 1422.6000 342.4500 1423.8000 342.6000 ;
	    RECT 1437.0000 342.4500 1438.2001 342.6000 ;
	    RECT 1422.6000 341.5500 1438.2001 342.4500 ;
	    RECT 1422.6000 341.4000 1423.8000 341.5500 ;
	    RECT 1437.0000 341.4000 1438.2001 341.5500 ;
	    RECT 1377.0000 339.4500 1378.2001 339.6000 ;
	    RECT 1391.4000 339.4500 1392.6000 339.6000 ;
	    RECT 1278.6000 338.4000 1279.8000 338.5500 ;
	    RECT 1295.4000 338.4000 1296.6000 338.5500 ;
	    RECT 1298.7001 338.4000 1301.4000 339.3000 ;
	    RECT 1278.6000 337.2000 1279.8000 337.5000 ;
	    RECT 1278.6000 333.3000 1279.8000 336.3000 ;
	    RECT 1298.7001 333.3000 1299.9000 338.4000 ;
	    RECT 1302.6000 333.3000 1303.8000 339.3000 ;
	    RECT 1329.0000 333.3000 1330.2001 339.3000 ;
	    RECT 1331.4000 339.0000 1337.4000 339.3000 ;
	    RECT 1331.4000 333.3000 1332.6000 339.0000 ;
	    RECT 1333.8000 333.3000 1335.0000 338.1000 ;
	    RECT 1336.2001 333.3000 1337.4000 339.0000 ;
	    RECT 1370.7001 333.3000 1371.9000 339.3000 ;
	    RECT 1374.6000 333.3000 1375.8000 339.3000 ;
	    RECT 1377.0000 338.5500 1392.6000 339.4500 ;
	    RECT 1401.3000 339.3000 1402.2001 340.5000 ;
	    RECT 1403.7001 339.3000 1409.1000 339.9000 ;
	    RECT 1439.4000 339.3000 1440.3000 344.7000 ;
	    RECT 1441.8000 344.5500 1459.8000 345.4500 ;
	    RECT 1441.8000 344.4000 1443.0000 344.5500 ;
	    RECT 1451.4000 344.4000 1452.6000 344.5500 ;
	    RECT 1458.6000 344.4000 1459.8000 344.5500 ;
	    RECT 1468.5000 342.6000 1469.4000 346.5000 ;
	    RECT 1475.4000 346.2000 1476.6000 346.5000 ;
	    RECT 1559.4000 346.2000 1560.6000 346.5000 ;
	    RECT 1523.1000 345.6000 1524.3000 345.9000 ;
	    RECT 1471.8000 344.4000 1472.1000 345.6000 ;
	    RECT 1473.0000 344.4000 1474.2001 345.6000 ;
	    RECT 1521.9000 344.7000 1524.3000 345.6000 ;
	    RECT 1525.8000 345.4500 1527.0000 345.6000 ;
	    RECT 1537.8000 345.4500 1539.0000 345.6000 ;
	    RECT 1521.9000 344.4000 1523.1000 344.7000 ;
	    RECT 1525.8000 344.5500 1539.0000 345.4500 ;
	    RECT 1525.8000 344.4000 1527.0000 344.5500 ;
	    RECT 1537.8000 344.4000 1539.0000 344.5500 ;
	    RECT 1561.8000 344.4000 1563.0000 345.6000 ;
	    RECT 1563.9000 344.4000 1564.2001 345.6000 ;
	    RECT 1524.0000 342.9000 1525.2001 343.2000 ;
	    RECT 1521.0000 342.6000 1525.2001 342.9000 ;
	    RECT 1468.5000 342.3000 1470.9000 342.6000 ;
	    RECT 1501.8000 342.4500 1503.0000 342.6000 ;
	    RECT 1509.0000 342.4500 1510.2001 342.6000 ;
	    RECT 1518.6000 342.4500 1519.8000 342.6000 ;
	    RECT 1468.5000 341.7000 1471.2001 342.3000 ;
	    RECT 1377.0000 338.4000 1378.2001 338.5500 ;
	    RECT 1391.4000 338.4000 1392.6000 338.5500 ;
	    RECT 1376.7001 337.2000 1377.9000 337.5000 ;
	    RECT 1377.0000 333.3000 1378.2001 336.3000 ;
	    RECT 1401.0000 333.3000 1402.2001 339.3000 ;
	    RECT 1403.4000 339.0000 1409.4000 339.3000 ;
	    RECT 1403.4000 333.3000 1404.6000 339.0000 ;
	    RECT 1405.8000 333.3000 1407.0000 338.1000 ;
	    RECT 1408.2001 333.3000 1409.4000 339.0000 ;
	    RECT 1435.5000 333.3000 1436.7001 339.3000 ;
	    RECT 1439.4000 333.3000 1440.6000 339.3000 ;
	    RECT 1441.8000 338.4000 1443.0000 339.6000 ;
	    RECT 1441.5000 337.2000 1442.7001 337.5000 ;
	    RECT 1446.6000 336.4500 1447.8000 336.6000 ;
	    RECT 1461.0000 336.4500 1462.2001 336.6000 ;
	    RECT 1441.8000 333.3000 1443.0000 336.3000 ;
	    RECT 1446.6000 335.5500 1462.2001 336.4500 ;
	    RECT 1446.6000 335.4000 1447.8000 335.5500 ;
	    RECT 1461.0000 335.4000 1462.2001 335.5500 ;
	    RECT 1470.0000 333.3000 1471.2001 341.7000 ;
	    RECT 1475.4000 333.3000 1476.6000 342.3000 ;
	    RECT 1501.8000 341.5500 1519.8000 342.4500 ;
	    RECT 1501.8000 341.4000 1503.0000 341.5500 ;
	    RECT 1509.0000 341.4000 1510.2001 341.5500 ;
	    RECT 1518.6000 341.4000 1519.8000 341.5500 ;
	    RECT 1520.7001 342.0000 1525.2001 342.6000 ;
	    RECT 1526.1000 342.6000 1527.0000 343.5000 ;
	    RECT 1566.6000 342.6000 1567.5000 346.5000 ;
	    RECT 1520.7001 341.7000 1521.9000 342.0000 ;
	    RECT 1526.1000 341.7000 1527.6000 342.6000 ;
	    RECT 1520.7001 341.4000 1521.0000 341.7000 ;
	    RECT 1521.3000 340.2000 1522.5000 340.5000 ;
	    RECT 1518.6000 339.3000 1522.5000 340.2000 ;
	    RECT 1523.4000 339.6000 1525.8000 340.8000 ;
	    RECT 1518.6000 333.3000 1519.8000 339.3000 ;
	    RECT 1526.7001 338.7000 1527.6000 341.7000 ;
	    RECT 1528.8000 341.4000 1530.0000 342.6000 ;
	    RECT 1531.8000 341.4000 1532.1000 342.6000 ;
	    RECT 1533.0000 342.4500 1534.2001 342.6000 ;
	    RECT 1540.2001 342.4500 1541.4000 342.6000 ;
	    RECT 1533.0000 341.5500 1541.4000 342.4500 ;
	    RECT 1565.1000 342.3000 1567.5000 342.6000 ;
	    RECT 1533.0000 341.4000 1534.2001 341.5500 ;
	    RECT 1540.2001 341.4000 1541.4000 341.5500 ;
	    RECT 1528.8000 340.8000 1529.7001 341.4000 ;
	    RECT 1528.5000 339.6000 1529.7001 340.8000 ;
	    RECT 1530.6000 340.2000 1531.8000 340.5000 ;
	    RECT 1530.6000 339.3000 1534.2001 340.2000 ;
	    RECT 1521.0000 333.3000 1522.5000 338.4000 ;
	    RECT 1525.2001 333.3000 1527.6000 338.7000 ;
	    RECT 1530.3000 333.3000 1531.8000 338.4000 ;
	    RECT 1533.0000 333.3000 1534.2001 339.3000 ;
	    RECT 1559.4000 333.3000 1560.6000 342.3000 ;
	    RECT 1564.8000 341.7000 1567.5000 342.3000 ;
	    RECT 1564.8000 333.3000 1566.0000 341.7000 ;
	    RECT 1.2000 330.6000 1569.0000 332.4000 ;
	    RECT 25.8000 324.0000 27.0000 329.7000 ;
	    RECT 28.2000 324.9000 29.4000 329.7000 ;
	    RECT 30.6000 324.0000 31.8000 329.7000 ;
	    RECT 25.8000 323.7000 31.8000 324.0000 ;
	    RECT 33.0000 323.7000 34.2000 329.7000 ;
	    RECT 26.1000 323.1000 31.5000 323.7000 ;
	    RECT 33.0000 322.5000 33.9000 323.7000 ;
	    RECT 45.0000 322.5000 46.2000 329.7000 ;
	    RECT 47.4000 326.7000 48.6000 329.7000 ;
	    RECT 47.4000 325.5000 48.6000 325.8000 ;
	    RECT 67.5000 324.6000 68.7000 329.7000 ;
	    RECT 47.4000 324.4500 48.6000 324.6000 ;
	    RECT 64.2000 324.4500 65.4000 324.6000 ;
	    RECT 47.4000 323.5500 65.4000 324.4500 ;
	    RECT 67.5000 323.7000 70.2000 324.6000 ;
	    RECT 71.4000 323.7000 72.6000 329.7000 ;
	    RECT 47.4000 323.4000 48.6000 323.5500 ;
	    RECT 64.2000 323.4000 65.4000 323.5500 ;
	    RECT 25.8000 320.4000 27.0000 321.6000 ;
	    RECT 27.9000 320.7000 28.2000 322.2000 ;
	    RECT 30.3000 320.4000 32.1000 321.6000 ;
	    RECT 33.0000 320.4000 34.2000 321.6000 ;
	    RECT 35.4000 321.4500 36.6000 321.6000 ;
	    RECT 45.0000 321.4500 46.2000 321.6000 ;
	    RECT 35.4000 320.5500 46.2000 321.4500 ;
	    RECT 35.4000 320.4000 36.6000 320.5500 ;
	    RECT 45.0000 320.4000 46.2000 320.5500 ;
	    RECT 28.2000 319.5000 29.4000 319.8000 ;
	    RECT 28.2000 317.4000 29.4000 318.6000 ;
	    RECT 30.3000 315.3000 31.2000 320.4000 ;
	    RECT 69.0000 319.5000 70.2000 323.7000 ;
	    RECT 71.4000 322.5000 72.6000 322.8000 ;
	    RECT 85.8000 322.5000 87.0000 329.7000 ;
	    RECT 88.2000 326.7000 89.4000 329.7000 ;
	    RECT 88.2000 325.5000 89.4000 325.8000 ;
	    RECT 88.2000 324.4500 89.4000 324.6000 ;
	    RECT 141.0000 324.4500 142.2000 324.6000 ;
	    RECT 88.2000 323.5500 142.2000 324.4500 ;
	    RECT 143.4000 323.7000 144.6000 329.7000 ;
	    RECT 88.2000 323.4000 89.4000 323.5500 ;
	    RECT 141.0000 323.4000 142.2000 323.5500 ;
	    RECT 145.8000 322.8000 147.0000 329.7000 ;
	    RECT 148.2000 323.7000 149.4000 329.7000 ;
	    RECT 150.6000 322.8000 151.8000 329.7000 ;
	    RECT 153.0000 323.7000 154.2000 329.7000 ;
	    RECT 155.4000 322.8000 156.6000 329.7000 ;
	    RECT 157.8000 323.7000 159.0000 329.7000 ;
	    RECT 160.2000 322.8000 161.4000 329.7000 ;
	    RECT 162.6000 323.7000 163.8000 329.7000 ;
	    RECT 174.6000 326.7000 175.8000 329.7000 ;
	    RECT 174.6000 325.5000 175.8000 325.8000 ;
	    RECT 174.6000 323.4000 175.8000 324.6000 ;
	    RECT 145.8000 321.6000 148.5000 322.8000 ;
	    RECT 150.6000 321.6000 153.9000 322.8000 ;
	    RECT 155.4000 321.6000 158.7000 322.8000 ;
	    RECT 160.2000 321.6000 163.8000 322.8000 ;
	    RECT 177.0000 322.5000 178.2000 329.7000 ;
	    RECT 196.2000 323.7000 197.4000 329.7000 ;
	    RECT 200.1000 324.6000 201.3000 329.7000 ;
	    RECT 198.6000 323.7000 201.3000 324.6000 ;
	    RECT 232.2000 323.7000 233.4000 329.7000 ;
	    RECT 234.6000 324.0000 235.8000 329.7000 ;
	    RECT 237.0000 324.9000 238.2000 329.7000 ;
	    RECT 239.4000 324.0000 240.6000 329.7000 ;
	    RECT 234.6000 323.7000 240.6000 324.0000 ;
	    RECT 196.2000 322.5000 197.4000 322.8000 ;
	    RECT 71.4000 321.4500 72.6000 321.6000 ;
	    RECT 73.8000 321.4500 75.0000 321.6000 ;
	    RECT 71.4000 320.5500 75.0000 321.4500 ;
	    RECT 71.4000 320.4000 72.6000 320.5500 ;
	    RECT 73.8000 320.4000 75.0000 320.5500 ;
	    RECT 76.2000 321.4500 77.4000 321.6000 ;
	    RECT 85.8000 321.4500 87.0000 321.6000 ;
	    RECT 76.2000 320.5500 87.0000 321.4500 ;
	    RECT 76.2000 320.4000 77.4000 320.5500 ;
	    RECT 85.8000 320.4000 87.0000 320.5500 ;
	    RECT 105.0000 321.4500 106.2000 321.6000 ;
	    RECT 143.4000 321.4500 144.6000 321.6000 ;
	    RECT 105.0000 320.5500 144.6000 321.4500 ;
	    RECT 147.3000 320.7000 148.5000 321.6000 ;
	    RECT 152.7000 320.7000 153.9000 321.6000 ;
	    RECT 157.5000 320.7000 158.7000 321.6000 ;
	    RECT 105.0000 320.4000 106.2000 320.5500 ;
	    RECT 143.4000 320.4000 144.6000 320.5500 ;
	    RECT 145.5000 319.5000 146.1000 320.7000 ;
	    RECT 147.3000 319.5000 151.2000 320.7000 ;
	    RECT 152.7000 319.5000 156.3000 320.7000 ;
	    RECT 157.5000 319.5000 161.4000 320.7000 ;
	    RECT 162.6000 319.5000 163.8000 321.6000 ;
	    RECT 177.0000 321.4500 178.2000 321.6000 ;
	    RECT 184.2000 321.4500 185.4000 321.6000 ;
	    RECT 177.0000 320.5500 185.4000 321.4500 ;
	    RECT 177.0000 320.4000 178.2000 320.5500 ;
	    RECT 184.2000 320.4000 185.4000 320.5500 ;
	    RECT 186.6000 321.4500 187.8000 321.6000 ;
	    RECT 196.2000 321.4500 197.4000 321.6000 ;
	    RECT 186.6000 320.5500 197.4000 321.4500 ;
	    RECT 186.6000 320.4000 187.8000 320.5500 ;
	    RECT 196.2000 320.4000 197.4000 320.5500 ;
	    RECT 198.6000 319.5000 199.8000 323.7000 ;
	    RECT 232.5000 322.5000 233.4000 323.7000 ;
	    RECT 234.9000 323.1000 240.3000 323.7000 ;
	    RECT 253.8000 322.5000 255.0000 329.7000 ;
	    RECT 256.2000 326.7000 257.4000 329.7000 ;
	    RECT 256.2000 325.5000 257.4000 325.8000 ;
	    RECT 256.2000 323.4000 257.4000 324.6000 ;
	    RECT 275.4000 323.7000 276.6000 329.7000 ;
	    RECT 279.3000 324.6000 280.5000 329.7000 ;
	    RECT 405.0000 326.7000 406.2000 329.7000 ;
	    RECT 277.8000 323.7000 280.5000 324.6000 ;
	    RECT 407.4000 324.0000 408.6000 329.7000 ;
	    RECT 275.4000 322.5000 276.6000 322.8000 ;
	    RECT 232.2000 320.4000 233.4000 321.6000 ;
	    RECT 234.3000 320.4000 236.1000 321.6000 ;
	    RECT 238.2000 320.7000 238.5000 322.2000 ;
	    RECT 239.4000 320.4000 240.6000 321.6000 ;
	    RECT 253.8000 321.4500 255.0000 321.6000 ;
	    RECT 241.9500 320.5500 255.0000 321.4500 ;
	    RECT 25.8000 303.3000 27.0000 315.3000 ;
	    RECT 29.7000 314.4000 31.2000 315.3000 ;
	    RECT 33.0000 315.4500 34.2000 315.6000 ;
	    RECT 40.2000 315.4500 41.4000 315.6000 ;
	    RECT 33.0000 314.5500 41.4000 315.4500 ;
	    RECT 33.0000 314.4000 34.2000 314.5500 ;
	    RECT 40.2000 314.4000 41.4000 314.5500 ;
	    RECT 29.7000 303.3000 30.9000 314.4000 ;
	    RECT 32.1000 312.6000 33.0000 313.5000 ;
	    RECT 31.8000 311.4000 33.0000 312.6000 ;
	    RECT 32.1000 303.3000 33.3000 309.3000 ;
	    RECT 45.0000 303.3000 46.2000 319.5000 ;
	    RECT 47.4000 318.4500 48.6000 318.6000 ;
	    RECT 69.0000 318.4500 70.2000 318.6000 ;
	    RECT 47.4000 317.5500 70.2000 318.4500 ;
	    RECT 47.4000 317.4000 48.6000 317.5500 ;
	    RECT 69.0000 317.4000 70.2000 317.5500 ;
	    RECT 66.6000 314.4000 67.8000 315.6000 ;
	    RECT 66.6000 313.2000 67.8000 313.5000 ;
	    RECT 47.4000 303.3000 48.6000 309.3000 ;
	    RECT 66.6000 303.3000 67.8000 309.3000 ;
	    RECT 69.0000 303.3000 70.2000 316.5000 ;
	    RECT 71.4000 303.3000 72.6000 309.3000 ;
	    RECT 85.8000 303.3000 87.0000 319.5000 ;
	    RECT 147.3000 317.4000 148.5000 319.5000 ;
	    RECT 152.7000 317.4000 153.9000 319.5000 ;
	    RECT 157.5000 317.4000 158.7000 319.5000 ;
	    RECT 162.6000 318.4500 163.8000 318.6000 ;
	    RECT 167.4000 318.4500 168.6000 318.6000 ;
	    RECT 162.6000 317.5500 168.6000 318.4500 ;
	    RECT 162.6000 317.4000 163.8000 317.5500 ;
	    RECT 167.4000 317.4000 168.6000 317.5500 ;
	    RECT 145.8000 316.2000 148.5000 317.4000 ;
	    RECT 150.6000 316.2000 153.9000 317.4000 ;
	    RECT 155.4000 316.2000 158.7000 317.4000 ;
	    RECT 160.2000 316.5000 161.7000 317.4000 ;
	    RECT 160.2000 316.2000 163.8000 316.5000 ;
	    RECT 88.2000 303.3000 89.4000 309.3000 ;
	    RECT 143.4000 303.3000 144.6000 315.3000 ;
	    RECT 145.8000 303.3000 147.0000 316.2000 ;
	    RECT 148.2000 303.3000 149.4000 315.3000 ;
	    RECT 150.6000 303.3000 151.8000 316.2000 ;
	    RECT 153.0000 303.3000 154.2000 315.3000 ;
	    RECT 155.4000 303.3000 156.6000 316.2000 ;
	    RECT 157.8000 303.3000 159.0000 315.3000 ;
	    RECT 160.2000 303.3000 161.4000 316.2000 ;
	    RECT 162.6000 303.3000 163.8000 315.3000 ;
	    RECT 174.6000 303.3000 175.8000 309.3000 ;
	    RECT 177.0000 303.3000 178.2000 319.5000 ;
	    RECT 198.6000 318.4500 199.8000 318.6000 ;
	    RECT 198.6000 317.5500 233.2500 318.4500 ;
	    RECT 198.6000 317.4000 199.8000 317.5500 ;
	    RECT 196.2000 303.3000 197.4000 309.3000 ;
	    RECT 198.6000 303.3000 199.8000 316.5000 ;
	    RECT 232.3500 315.6000 233.2500 317.5500 ;
	    RECT 201.0000 314.4000 202.2000 315.6000 ;
	    RECT 232.2000 314.4000 233.4000 315.6000 ;
	    RECT 235.2000 315.3000 236.1000 320.4000 ;
	    RECT 237.0000 319.5000 238.2000 319.8000 ;
	    RECT 237.0000 318.4500 238.2000 318.6000 ;
	    RECT 241.9500 318.4500 242.8500 320.5500 ;
	    RECT 253.8000 320.4000 255.0000 320.5500 ;
	    RECT 273.0000 321.4500 274.2000 321.6000 ;
	    RECT 275.4000 321.4500 276.6000 321.6000 ;
	    RECT 273.0000 320.5500 276.6000 321.4500 ;
	    RECT 273.0000 320.4000 274.2000 320.5500 ;
	    RECT 275.4000 320.4000 276.6000 320.5500 ;
	    RECT 277.8000 319.5000 279.0000 323.7000 ;
	    RECT 407.1000 322.8000 408.6000 324.0000 ;
	    RECT 237.0000 317.5500 242.8500 318.4500 ;
	    RECT 237.0000 317.4000 238.2000 317.5500 ;
	    RECT 235.2000 314.4000 236.7000 315.3000 ;
	    RECT 201.0000 313.2000 202.2000 313.5000 ;
	    RECT 233.4000 312.6000 234.3000 313.5000 ;
	    RECT 233.4000 311.4000 234.6000 312.6000 ;
	    RECT 201.0000 303.3000 202.2000 309.3000 ;
	    RECT 233.1000 303.3000 234.3000 309.3000 ;
	    RECT 235.5000 303.3000 236.7000 314.4000 ;
	    RECT 239.4000 303.3000 240.6000 315.3000 ;
	    RECT 253.8000 303.3000 255.0000 319.5000 ;
	    RECT 277.8000 318.4500 279.0000 318.6000 ;
	    RECT 280.2000 318.4500 281.4000 318.6000 ;
	    RECT 277.8000 317.5500 281.4000 318.4500 ;
	    RECT 277.8000 317.4000 279.0000 317.5500 ;
	    RECT 280.2000 317.4000 281.4000 317.5500 ;
	    RECT 256.2000 303.3000 257.4000 309.3000 ;
	    RECT 275.4000 303.3000 276.6000 309.3000 ;
	    RECT 277.8000 303.3000 279.0000 316.5000 ;
	    RECT 407.1000 316.2000 408.3000 322.8000 ;
	    RECT 409.8000 321.9000 411.0000 329.7000 ;
	    RECT 414.6000 323.7000 415.8000 329.7000 ;
	    RECT 419.4000 324.9000 420.6000 329.7000 ;
	    RECT 421.8000 325.5000 423.0000 329.7000 ;
	    RECT 424.2000 325.5000 425.4000 329.7000 ;
	    RECT 426.6000 325.5000 427.8000 329.7000 ;
	    RECT 429.0000 325.5000 430.2000 329.7000 ;
	    RECT 431.4000 326.7000 432.6000 329.7000 ;
	    RECT 433.8000 325.5000 435.0000 329.7000 ;
	    RECT 436.2000 326.7000 437.4000 329.7000 ;
	    RECT 438.6000 325.5000 439.8000 329.7000 ;
	    RECT 441.0000 325.5000 442.2000 329.7000 ;
	    RECT 443.4000 325.5000 444.6000 329.7000 ;
	    RECT 417.0000 323.7000 420.6000 324.9000 ;
	    RECT 445.8000 324.9000 447.0000 329.7000 ;
	    RECT 417.0000 322.8000 418.2000 323.7000 ;
	    RECT 409.2000 321.0000 411.0000 321.9000 ;
	    RECT 415.5000 321.9000 418.2000 322.8000 ;
	    RECT 424.2000 323.4000 425.7000 324.6000 ;
	    RECT 430.2000 323.4000 430.5000 324.6000 ;
	    RECT 431.4000 323.4000 432.6000 324.6000 ;
	    RECT 433.8000 323.7000 440.7000 324.6000 ;
	    RECT 445.8000 323.7000 449.7000 324.9000 ;
	    RECT 450.6000 323.7000 451.8000 329.7000 ;
	    RECT 433.8000 323.4000 435.0000 323.7000 ;
	    RECT 409.2000 318.0000 410.1000 321.0000 ;
	    RECT 415.5000 320.1000 416.7000 321.9000 ;
	    RECT 411.0000 318.9000 416.7000 320.1000 ;
	    RECT 424.2000 319.2000 425.4000 323.4000 ;
	    RECT 436.2000 322.5000 437.4000 322.8000 ;
	    RECT 433.8000 322.2000 435.0000 322.5000 ;
	    RECT 428.4000 321.3000 435.0000 322.2000 ;
	    RECT 428.4000 321.0000 429.6000 321.3000 ;
	    RECT 436.2000 320.4000 437.4000 321.6000 ;
	    RECT 439.5000 320.1000 440.7000 323.7000 ;
	    RECT 448.5000 322.8000 449.7000 323.7000 ;
	    RECT 448.5000 321.6000 453.0000 322.8000 ;
	    RECT 455.4000 320.7000 456.6000 329.7000 ;
	    RECT 477.0000 322.5000 478.2000 329.7000 ;
	    RECT 479.4000 326.7000 480.6000 329.7000 ;
	    RECT 479.4000 325.5000 480.6000 325.8000 ;
	    RECT 479.4000 323.4000 480.6000 324.6000 ;
	    RECT 479.5500 321.6000 480.4500 323.4000 ;
	    RECT 498.6000 322.5000 499.8000 329.7000 ;
	    RECT 501.0000 323.7000 502.2000 329.7000 ;
	    RECT 503.4000 322.8000 504.6000 329.7000 ;
	    RECT 529.8000 323.7000 531.0000 329.7000 ;
	    RECT 532.2000 324.0000 533.4000 329.7000 ;
	    RECT 534.6000 324.9000 535.8000 329.7000 ;
	    RECT 537.0000 324.0000 538.2000 329.7000 ;
	    RECT 532.2000 323.7000 538.2000 324.0000 ;
	    RECT 501.3000 321.9000 504.6000 322.8000 ;
	    RECT 530.1000 322.5000 531.0000 323.7000 ;
	    RECT 532.5000 323.1000 537.9000 323.7000 ;
	    RECT 549.0000 322.5000 550.2000 329.7000 ;
	    RECT 551.4000 326.7000 552.6000 329.7000 ;
	    RECT 551.4000 325.5000 552.6000 325.8000 ;
	    RECT 578.7000 325.2000 579.9000 329.7000 ;
	    RECT 551.4000 324.4500 552.6000 324.6000 ;
	    RECT 565.8000 324.4500 567.0000 324.6000 ;
	    RECT 575.4000 324.4500 576.6000 324.6000 ;
	    RECT 551.4000 323.5500 576.6000 324.4500 ;
	    RECT 551.4000 323.4000 552.6000 323.5500 ;
	    RECT 565.8000 323.4000 567.0000 323.5500 ;
	    RECT 575.4000 323.4000 576.6000 323.5500 ;
	    RECT 577.8000 323.7000 579.9000 325.2000 ;
	    RECT 581.1000 324.0000 582.3000 329.7000 ;
	    RECT 585.0000 323.7000 586.2000 329.7000 ;
	    RECT 429.0000 318.9000 433.8000 320.1000 ;
	    RECT 439.5000 318.9000 442.5000 320.1000 ;
	    RECT 443.4000 319.5000 456.6000 320.7000 ;
	    RECT 457.8000 321.4500 459.0000 321.6000 ;
	    RECT 477.0000 321.4500 478.2000 321.6000 ;
	    RECT 457.8000 320.5500 478.2000 321.4500 ;
	    RECT 457.8000 320.4000 459.0000 320.5500 ;
	    RECT 477.0000 320.4000 478.2000 320.5500 ;
	    RECT 479.4000 321.4500 480.6000 321.6000 ;
	    RECT 498.6000 321.4500 499.8000 321.6000 ;
	    RECT 479.4000 320.5500 499.8000 321.4500 ;
	    RECT 479.4000 320.4000 480.6000 320.5500 ;
	    RECT 498.6000 320.4000 499.8000 320.5500 ;
	    RECT 419.4000 318.0000 420.6000 318.9000 ;
	    RECT 409.2000 317.1000 410.4000 318.0000 ;
	    RECT 419.4000 317.1000 444.9000 318.0000 ;
	    RECT 445.8000 317.4000 447.0000 318.6000 ;
	    RECT 453.3000 318.0000 454.5000 318.3000 ;
	    RECT 447.9000 317.1000 454.5000 318.0000 ;
	    RECT 280.2000 315.4500 281.4000 315.6000 ;
	    RECT 282.6000 315.4500 283.8000 315.6000 ;
	    RECT 280.2000 314.5500 283.8000 315.4500 ;
	    RECT 280.2000 314.4000 281.4000 314.5500 ;
	    RECT 282.6000 314.4000 283.8000 314.5500 ;
	    RECT 306.6000 315.4500 307.8000 315.6000 ;
	    RECT 385.8000 315.4500 387.0000 315.6000 ;
	    RECT 306.6000 314.5500 387.0000 315.4500 ;
	    RECT 407.1000 315.0000 408.6000 316.2000 ;
	    RECT 306.6000 314.4000 307.8000 314.5500 ;
	    RECT 385.8000 314.4000 387.0000 314.5500 ;
	    RECT 407.4000 313.5000 408.6000 315.0000 ;
	    RECT 409.5000 314.4000 410.4000 317.1000 ;
	    RECT 411.3000 316.2000 412.5000 316.5000 ;
	    RECT 411.3000 315.3000 449.7000 316.2000 ;
	    RECT 445.5000 315.0000 446.7000 315.3000 ;
	    RECT 450.6000 314.4000 451.8000 315.6000 ;
	    RECT 409.5000 313.5000 423.0000 314.4000 ;
	    RECT 280.2000 313.2000 281.4000 313.5000 ;
	    RECT 357.0000 312.4500 358.2000 312.6000 ;
	    RECT 407.4000 312.4500 408.6000 312.6000 ;
	    RECT 357.0000 311.5500 408.6000 312.4500 ;
	    RECT 357.0000 311.4000 358.2000 311.5500 ;
	    RECT 407.4000 311.4000 408.6000 311.5500 ;
	    RECT 409.5000 311.1000 410.4000 313.5000 ;
	    RECT 421.8000 313.2000 423.0000 313.5000 ;
	    RECT 426.6000 313.5000 439.5000 314.4000 ;
	    RECT 426.6000 313.2000 427.8000 313.5000 ;
	    RECT 414.3000 311.4000 418.2000 312.6000 ;
	    RECT 280.2000 303.3000 281.4000 309.3000 ;
	    RECT 287.4000 306.4500 288.6000 306.6000 ;
	    RECT 323.4000 306.4500 324.6000 306.6000 ;
	    RECT 364.2000 306.4500 365.4000 306.6000 ;
	    RECT 287.4000 305.5500 365.4000 306.4500 ;
	    RECT 287.4000 305.4000 288.6000 305.5500 ;
	    RECT 323.4000 305.4000 324.6000 305.5500 ;
	    RECT 364.2000 305.4000 365.4000 305.5500 ;
	    RECT 405.0000 303.3000 406.2000 309.3000 ;
	    RECT 407.4000 303.3000 408.6000 310.5000 ;
	    RECT 409.5000 310.2000 413.4000 311.1000 ;
	    RECT 409.8000 303.3000 411.0000 309.3000 ;
	    RECT 412.2000 303.3000 413.4000 310.2000 ;
	    RECT 414.6000 303.3000 415.8000 309.3000 ;
	    RECT 417.0000 303.3000 418.2000 311.4000 ;
	    RECT 419.1000 310.2000 425.4000 311.4000 ;
	    RECT 419.4000 303.3000 420.6000 309.3000 ;
	    RECT 421.8000 303.3000 423.0000 307.5000 ;
	    RECT 424.2000 303.3000 425.4000 307.5000 ;
	    RECT 426.6000 303.3000 427.8000 307.5000 ;
	    RECT 429.0000 303.3000 430.2000 312.6000 ;
	    RECT 433.8000 311.4000 437.7000 312.6000 ;
	    RECT 438.6000 312.3000 439.5000 313.5000 ;
	    RECT 441.0000 314.1000 442.2000 314.4000 ;
	    RECT 441.0000 313.5000 449.1000 314.1000 ;
	    RECT 441.0000 313.2000 450.3000 313.5000 ;
	    RECT 448.2000 312.3000 450.3000 313.2000 ;
	    RECT 438.6000 311.4000 447.3000 312.3000 ;
	    RECT 451.8000 312.0000 454.2000 313.2000 ;
	    RECT 451.8000 311.4000 452.7000 312.0000 ;
	    RECT 431.4000 303.3000 432.6000 309.3000 ;
	    RECT 433.8000 303.3000 435.0000 310.5000 ;
	    RECT 436.2000 303.3000 437.4000 309.3000 ;
	    RECT 438.6000 303.3000 439.8000 310.5000 ;
	    RECT 446.4000 310.2000 452.7000 311.4000 ;
	    RECT 455.4000 311.1000 456.6000 319.5000 ;
	    RECT 453.6000 310.2000 456.6000 311.1000 ;
	    RECT 441.0000 303.3000 442.2000 307.5000 ;
	    RECT 443.4000 303.3000 444.6000 307.5000 ;
	    RECT 445.8000 303.3000 447.0000 309.3000 ;
	    RECT 448.2000 303.3000 449.4000 310.2000 ;
	    RECT 453.6000 309.3000 454.5000 310.2000 ;
	    RECT 450.6000 302.4000 451.8000 309.3000 ;
	    RECT 453.0000 308.4000 454.5000 309.3000 ;
	    RECT 453.0000 303.3000 454.2000 308.4000 ;
	    RECT 455.4000 303.3000 456.6000 309.3000 ;
	    RECT 477.0000 303.3000 478.2000 319.5000 ;
	    RECT 498.6000 318.6000 499.8000 319.5000 ;
	    RECT 498.6000 315.3000 499.5000 318.6000 ;
	    RECT 501.3000 317.4000 502.2000 321.9000 ;
	    RECT 529.8000 320.4000 531.0000 321.6000 ;
	    RECT 531.9000 320.4000 533.7000 321.6000 ;
	    RECT 535.8000 320.7000 536.1000 322.2000 ;
	    RECT 537.0000 320.4000 538.2000 321.6000 ;
	    RECT 549.0000 321.4500 550.2000 321.6000 ;
	    RECT 539.5500 320.5500 550.2000 321.4500 ;
	    RECT 503.4000 319.5000 504.6000 319.8000 ;
	    RECT 500.4000 316.2000 502.2000 317.4000 ;
	    RECT 501.3000 315.3000 502.2000 316.2000 ;
	    RECT 527.4000 315.4500 528.6000 315.6000 ;
	    RECT 529.8000 315.4500 531.0000 315.6000 ;
	    RECT 479.4000 303.3000 480.6000 309.3000 ;
	    RECT 498.6000 303.3000 499.8000 315.3000 ;
	    RECT 501.3000 314.4000 504.6000 315.3000 ;
	    RECT 527.4000 314.5500 531.0000 315.4500 ;
	    RECT 527.4000 314.4000 528.6000 314.5500 ;
	    RECT 529.8000 314.4000 531.0000 314.5500 ;
	    RECT 532.8000 315.3000 533.7000 320.4000 ;
	    RECT 534.6000 319.5000 535.8000 319.8000 ;
	    RECT 534.6000 318.4500 535.8000 318.6000 ;
	    RECT 539.5500 318.4500 540.4500 320.5500 ;
	    RECT 549.0000 320.4000 550.2000 320.5500 ;
	    RECT 577.8000 319.5000 578.7000 323.7000 ;
	    RECT 585.0000 323.4000 585.9000 323.7000 ;
	    RECT 583.2000 322.8000 585.9000 323.4000 ;
	    RECT 579.6000 322.5000 585.9000 322.8000 ;
	    RECT 661.8000 322.5000 663.0000 329.7000 ;
	    RECT 664.2000 323.7000 665.4000 329.7000 ;
	    RECT 668.4000 327.6000 669.6000 329.7000 ;
	    RECT 666.6000 326.7000 669.6000 327.6000 ;
	    RECT 672.3000 326.7000 673.8000 329.7000 ;
	    RECT 675.0000 326.7000 676.2000 329.7000 ;
	    RECT 677.4000 326.7000 678.6000 329.7000 ;
	    RECT 681.3000 327.6000 683.1000 329.7000 ;
	    RECT 681.0000 326.7000 683.1000 327.6000 ;
	    RECT 666.6000 325.5000 667.8000 326.7000 ;
	    RECT 675.0000 325.8000 675.9000 326.7000 ;
	    RECT 669.0000 324.6000 670.2000 325.8000 ;
	    RECT 671.7000 324.9000 675.9000 325.8000 ;
	    RECT 681.0000 325.5000 682.2000 326.7000 ;
	    RECT 671.7000 324.6000 672.9000 324.9000 ;
	    RECT 579.6000 321.9000 584.1000 322.5000 ;
	    RECT 579.6000 321.6000 580.8000 321.9000 ;
	    RECT 534.6000 317.5500 540.4500 318.4500 ;
	    RECT 534.6000 317.4000 535.8000 317.5500 ;
	    RECT 532.8000 314.4000 534.3000 315.3000 ;
	    RECT 501.0000 303.3000 502.2000 313.5000 ;
	    RECT 503.4000 303.3000 504.6000 314.4000 ;
	    RECT 531.0000 312.6000 531.9000 313.5000 ;
	    RECT 531.0000 311.4000 532.2000 312.6000 ;
	    RECT 530.7000 303.3000 531.9000 309.3000 ;
	    RECT 533.1000 303.3000 534.3000 314.4000 ;
	    RECT 537.0000 303.3000 538.2000 315.3000 ;
	    RECT 549.0000 303.3000 550.2000 319.5000 ;
	    RECT 577.8000 317.4000 579.0000 318.6000 ;
	    RECT 579.9000 316.5000 580.8000 321.6000 ;
	    RECT 585.0000 321.4500 586.2000 321.6000 ;
	    RECT 609.0000 321.4500 610.2000 321.6000 ;
	    RECT 582.0000 320.7000 583.2000 321.0000 ;
	    RECT 582.0000 319.8000 583.5000 320.7000 ;
	    RECT 585.0000 320.5500 610.2000 321.4500 ;
	    RECT 585.0000 320.4000 586.2000 320.5500 ;
	    RECT 609.0000 320.4000 610.2000 320.5500 ;
	    RECT 663.0000 320.4000 663.3000 321.6000 ;
	    RECT 664.2000 320.4000 665.4000 321.6000 ;
	    RECT 669.3000 321.3000 670.2000 324.6000 ;
	    RECT 685.8000 324.0000 687.0000 329.7000 ;
	    RECT 683.7000 323.1000 684.9000 323.4000 ;
	    RECT 688.2000 323.1000 689.4000 329.7000 ;
	    RECT 683.7000 322.2000 689.4000 323.1000 ;
	    RECT 702.6000 322.5000 703.8000 329.7000 ;
	    RECT 705.0000 326.7000 706.2000 329.7000 ;
	    RECT 705.0000 325.5000 706.2000 325.8000 ;
	    RECT 705.0000 324.4500 706.2000 324.6000 ;
	    RECT 717.0000 324.4500 718.2000 324.6000 ;
	    RECT 705.0000 323.5500 718.2000 324.4500 ;
	    RECT 705.0000 323.4000 706.2000 323.5500 ;
	    RECT 717.0000 323.4000 718.2000 323.5500 ;
	    RECT 724.2000 322.5000 725.4000 329.7000 ;
	    RECT 726.6000 323.7000 727.8000 329.7000 ;
	    RECT 729.0000 322.8000 730.2000 329.7000 ;
	    RECT 677.7000 321.3000 678.9000 321.6000 ;
	    RECT 666.3000 320.4000 679.5000 321.3000 ;
	    RECT 667.5000 320.1000 668.7000 320.4000 ;
	    RECT 582.6000 319.5000 583.5000 319.8000 ;
	    RECT 585.0000 319.2000 586.2000 319.5000 ;
	    RECT 665.1000 318.6000 666.3000 318.9000 ;
	    RECT 582.6000 317.4000 583.8000 318.6000 ;
	    RECT 665.1000 317.7000 670.5000 318.6000 ;
	    RECT 671.4000 317.4000 672.6000 318.6000 ;
	    RECT 661.8000 316.5000 670.2000 316.8000 ;
	    RECT 577.8000 315.3000 578.7000 316.5000 ;
	    RECT 579.9000 315.6000 583.5000 316.5000 ;
	    RECT 551.4000 303.3000 552.6000 309.3000 ;
	    RECT 577.8000 303.3000 579.0000 315.3000 ;
	    RECT 580.2000 303.3000 581.4000 314.7000 ;
	    RECT 582.6000 309.3000 583.5000 315.6000 ;
	    RECT 661.8000 316.2000 670.5000 316.5000 ;
	    RECT 661.8000 315.9000 676.5000 316.2000 ;
	    RECT 582.6000 303.3000 583.8000 309.3000 ;
	    RECT 585.0000 303.3000 586.2000 309.3000 ;
	    RECT 661.8000 303.3000 663.0000 315.9000 ;
	    RECT 669.3000 315.3000 676.5000 315.9000 ;
	    RECT 664.2000 303.3000 665.4000 315.0000 ;
	    RECT 666.6000 313.5000 674.7000 314.4000 ;
	    RECT 666.6000 313.2000 667.8000 313.5000 ;
	    RECT 673.5000 313.2000 674.7000 313.5000 ;
	    RECT 675.6000 313.5000 676.5000 315.3000 ;
	    RECT 678.6000 315.6000 679.5000 320.4000 ;
	    RECT 688.2000 319.5000 689.4000 322.2000 ;
	    RECT 726.9000 321.9000 730.2000 322.8000 ;
	    RECT 748.2000 322.5000 749.4000 329.7000 ;
	    RECT 750.6000 323.7000 751.8000 329.7000 ;
	    RECT 753.0000 322.8000 754.2000 329.7000 ;
	    RECT 777.0000 324.0000 778.2000 329.7000 ;
	    RECT 779.4000 324.9000 780.6000 329.7000 ;
	    RECT 781.8000 324.0000 783.0000 329.7000 ;
	    RECT 777.0000 323.7000 783.0000 324.0000 ;
	    RECT 784.2000 323.7000 785.4000 329.7000 ;
	    RECT 916.2000 326.7000 917.4000 329.7000 ;
	    RECT 918.6000 324.0000 919.8000 329.7000 ;
	    RECT 777.3000 323.1000 782.7000 323.7000 ;
	    RECT 750.9000 321.9000 754.2000 322.8000 ;
	    RECT 784.2000 322.5000 785.1000 323.7000 ;
	    RECT 918.3000 322.8000 919.8000 324.0000 ;
	    RECT 702.6000 321.4500 703.8000 321.6000 ;
	    RECT 721.8000 321.4500 723.0000 321.6000 ;
	    RECT 702.6000 320.5500 723.0000 321.4500 ;
	    RECT 702.6000 320.4000 703.8000 320.5500 ;
	    RECT 721.8000 320.4000 723.0000 320.5500 ;
	    RECT 724.2000 320.4000 725.4000 321.6000 ;
	    RECT 681.0000 319.2000 682.2000 319.5000 ;
	    RECT 681.0000 318.3000 686.7000 319.2000 ;
	    RECT 685.5000 318.0000 686.7000 318.3000 ;
	    RECT 688.2000 317.4000 689.4000 318.6000 ;
	    RECT 683.1000 317.1000 684.3000 317.4000 ;
	    RECT 683.1000 316.5000 687.3000 317.1000 ;
	    RECT 683.1000 316.2000 689.4000 316.5000 ;
	    RECT 678.6000 314.7000 682.2000 315.6000 ;
	    RECT 677.7000 313.5000 678.9000 313.8000 ;
	    RECT 675.6000 312.6000 678.9000 313.5000 ;
	    RECT 681.3000 313.2000 682.2000 314.7000 ;
	    RECT 681.3000 312.0000 683.4000 313.2000 ;
	    RECT 671.7000 311.1000 672.9000 311.4000 ;
	    RECT 675.9000 311.1000 677.1000 311.4000 ;
	    RECT 666.6000 309.3000 667.8000 310.5000 ;
	    RECT 671.7000 310.2000 677.1000 311.1000 ;
	    RECT 675.0000 309.3000 675.9000 310.2000 ;
	    RECT 681.0000 309.3000 682.2000 310.5000 ;
	    RECT 666.6000 308.4000 669.6000 309.3000 ;
	    RECT 668.4000 303.3000 669.6000 308.4000 ;
	    RECT 672.6000 303.3000 673.8000 309.3000 ;
	    RECT 675.0000 303.3000 676.2000 309.3000 ;
	    RECT 677.4000 303.3000 678.6000 309.3000 ;
	    RECT 681.3000 303.3000 683.1000 309.3000 ;
	    RECT 685.8000 303.3000 687.0000 315.3000 ;
	    RECT 688.2000 303.3000 689.4000 316.2000 ;
	    RECT 702.6000 303.3000 703.8000 319.5000 ;
	    RECT 724.2000 318.6000 725.4000 319.5000 ;
	    RECT 724.2000 315.3000 725.1000 318.6000 ;
	    RECT 726.9000 317.4000 727.8000 321.9000 ;
	    RECT 748.2000 320.4000 749.4000 321.6000 ;
	    RECT 729.0000 319.5000 730.2000 319.8000 ;
	    RECT 748.2000 318.6000 749.4000 319.5000 ;
	    RECT 729.0000 318.4500 730.2000 318.6000 ;
	    RECT 738.6000 318.4500 739.8000 318.6000 ;
	    RECT 729.0000 317.5500 739.8000 318.4500 ;
	    RECT 729.0000 317.4000 730.2000 317.5500 ;
	    RECT 738.6000 317.4000 739.8000 317.5500 ;
	    RECT 726.0000 316.2000 727.8000 317.4000 ;
	    RECT 726.9000 315.3000 727.8000 316.2000 ;
	    RECT 748.2000 315.3000 749.1000 318.6000 ;
	    RECT 750.9000 317.4000 751.8000 321.9000 ;
	    RECT 755.4000 321.4500 756.6000 321.6000 ;
	    RECT 767.4000 321.4500 768.6000 321.6000 ;
	    RECT 777.0000 321.4500 778.2000 321.6000 ;
	    RECT 755.4000 320.5500 778.2000 321.4500 ;
	    RECT 779.1000 320.7000 779.4000 322.2000 ;
	    RECT 755.4000 320.4000 756.6000 320.5500 ;
	    RECT 767.4000 320.4000 768.6000 320.5500 ;
	    RECT 777.0000 320.4000 778.2000 320.5500 ;
	    RECT 781.5000 320.4000 783.3000 321.6000 ;
	    RECT 784.2000 321.4500 785.4000 321.6000 ;
	    RECT 916.2000 321.4500 917.4000 321.6000 ;
	    RECT 784.2000 320.5500 917.4000 321.4500 ;
	    RECT 784.2000 320.4000 785.4000 320.5500 ;
	    RECT 916.2000 320.4000 917.4000 320.5500 ;
	    RECT 753.0000 319.5000 754.2000 319.8000 ;
	    RECT 779.4000 319.5000 780.6000 319.8000 ;
	    RECT 753.0000 317.4000 754.2000 318.6000 ;
	    RECT 779.4000 317.4000 780.6000 318.6000 ;
	    RECT 750.0000 316.2000 751.8000 317.4000 ;
	    RECT 750.9000 315.3000 751.8000 316.2000 ;
	    RECT 781.5000 315.3000 782.4000 320.4000 ;
	    RECT 918.3000 316.2000 919.5000 322.8000 ;
	    RECT 921.0000 321.9000 922.2000 329.7000 ;
	    RECT 925.8000 323.7000 927.0000 329.7000 ;
	    RECT 930.6000 324.9000 931.8000 329.7000 ;
	    RECT 933.0000 325.5000 934.2000 329.7000 ;
	    RECT 935.4000 325.5000 936.6000 329.7000 ;
	    RECT 937.8000 325.5000 939.0000 329.7000 ;
	    RECT 940.2000 325.5000 941.4000 329.7000 ;
	    RECT 942.6000 326.7000 943.8000 329.7000 ;
	    RECT 945.0000 325.5000 946.2000 329.7000 ;
	    RECT 947.4000 326.7000 948.6000 329.7000 ;
	    RECT 949.8000 325.5000 951.0000 329.7000 ;
	    RECT 952.2000 325.5000 953.4000 329.7000 ;
	    RECT 954.6000 325.5000 955.8000 329.7000 ;
	    RECT 928.2000 323.7000 931.8000 324.9000 ;
	    RECT 957.0000 324.9000 958.2000 329.7000 ;
	    RECT 928.2000 322.8000 929.4000 323.7000 ;
	    RECT 920.4000 321.0000 922.2000 321.9000 ;
	    RECT 926.7000 321.9000 929.4000 322.8000 ;
	    RECT 935.4000 323.4000 936.9000 324.6000 ;
	    RECT 941.4000 323.4000 941.7000 324.6000 ;
	    RECT 942.6000 323.4000 943.8000 324.6000 ;
	    RECT 945.0000 323.7000 951.9000 324.6000 ;
	    RECT 957.0000 323.7000 960.9000 324.9000 ;
	    RECT 961.8000 323.7000 963.0000 329.7000 ;
	    RECT 945.0000 323.4000 946.2000 323.7000 ;
	    RECT 920.4000 318.0000 921.3000 321.0000 ;
	    RECT 926.7000 320.1000 927.9000 321.9000 ;
	    RECT 922.2000 318.9000 927.9000 320.1000 ;
	    RECT 935.4000 319.2000 936.6000 323.4000 ;
	    RECT 947.4000 322.5000 948.6000 322.8000 ;
	    RECT 945.0000 322.2000 946.2000 322.5000 ;
	    RECT 939.6000 321.3000 946.2000 322.2000 ;
	    RECT 939.6000 321.0000 940.8000 321.3000 ;
	    RECT 947.4000 320.4000 948.6000 321.6000 ;
	    RECT 950.7000 320.1000 951.9000 323.7000 ;
	    RECT 959.7000 322.8000 960.9000 323.7000 ;
	    RECT 959.7000 321.6000 964.2000 322.8000 ;
	    RECT 966.6000 320.7000 967.8000 329.7000 ;
	    RECT 998.4000 323.7000 999.6000 329.7000 ;
	    RECT 1002.3000 323.7000 1004.7000 329.7000 ;
	    RECT 1007.4000 323.7000 1008.6000 329.7000 ;
	    RECT 1034.7001 325.2000 1035.9000 329.7000 ;
	    RECT 1033.8000 323.7000 1035.9000 325.2000 ;
	    RECT 1037.1000 324.0000 1038.3000 329.7000 ;
	    RECT 1041.0000 323.7000 1042.2001 329.7000 ;
	    RECT 940.2000 318.9000 945.0000 320.1000 ;
	    RECT 950.7000 318.9000 953.7000 320.1000 ;
	    RECT 954.6000 319.5000 967.8000 320.7000 ;
	    RECT 1000.2000 320.4000 1001.4000 321.6000 ;
	    RECT 1002.9000 319.5000 1003.8000 323.7000 ;
	    RECT 1005.0000 320.4000 1006.2000 321.6000 ;
	    RECT 1033.8000 319.5000 1034.7001 323.7000 ;
	    RECT 1041.0000 323.4000 1041.9000 323.7000 ;
	    RECT 1039.2001 322.8000 1041.9000 323.4000 ;
	    RECT 1035.6000 322.5000 1041.9000 322.8000 ;
	    RECT 1035.6000 321.9000 1040.1000 322.5000 ;
	    RECT 1035.6000 321.6000 1036.8000 321.9000 ;
	    RECT 930.6000 318.0000 931.8000 318.9000 ;
	    RECT 920.4000 317.1000 921.6000 318.0000 ;
	    RECT 930.6000 317.1000 956.1000 318.0000 ;
	    RECT 957.0000 317.4000 958.2000 318.6000 ;
	    RECT 964.5000 318.0000 965.7000 318.3000 ;
	    RECT 959.1000 317.1000 965.7000 318.0000 ;
	    RECT 705.0000 303.3000 706.2000 309.3000 ;
	    RECT 724.2000 303.3000 725.4000 315.3000 ;
	    RECT 726.9000 314.4000 730.2000 315.3000 ;
	    RECT 726.6000 303.3000 727.8000 313.5000 ;
	    RECT 729.0000 303.3000 730.2000 314.4000 ;
	    RECT 748.2000 303.3000 749.4000 315.3000 ;
	    RECT 750.9000 314.4000 754.2000 315.3000 ;
	    RECT 750.6000 303.3000 751.8000 313.5000 ;
	    RECT 753.0000 303.3000 754.2000 314.4000 ;
	    RECT 777.0000 303.3000 778.2000 315.3000 ;
	    RECT 780.9000 314.4000 782.4000 315.3000 ;
	    RECT 784.2000 315.4500 785.4000 315.6000 ;
	    RECT 861.0000 315.4500 862.2000 315.6000 ;
	    RECT 784.2000 314.5500 862.2000 315.4500 ;
	    RECT 918.3000 315.0000 919.8000 316.2000 ;
	    RECT 784.2000 314.4000 785.4000 314.5500 ;
	    RECT 861.0000 314.4000 862.2000 314.5500 ;
	    RECT 780.9000 303.3000 782.1000 314.4000 ;
	    RECT 918.6000 313.5000 919.8000 315.0000 ;
	    RECT 920.7000 314.4000 921.6000 317.1000 ;
	    RECT 922.5000 316.2000 923.7000 316.5000 ;
	    RECT 922.5000 315.3000 960.9000 316.2000 ;
	    RECT 956.7000 315.0000 957.9000 315.3000 ;
	    RECT 961.8000 314.4000 963.0000 315.6000 ;
	    RECT 920.7000 313.5000 934.2000 314.4000 ;
	    RECT 783.3000 312.6000 784.2000 313.5000 ;
	    RECT 783.0000 311.4000 784.2000 312.6000 ;
	    RECT 786.6000 312.4500 787.8000 312.6000 ;
	    RECT 918.6000 312.4500 919.8000 312.6000 ;
	    RECT 786.6000 311.5500 919.8000 312.4500 ;
	    RECT 786.6000 311.4000 787.8000 311.5500 ;
	    RECT 918.6000 311.4000 919.8000 311.5500 ;
	    RECT 920.7000 311.1000 921.6000 313.5000 ;
	    RECT 933.0000 313.2000 934.2000 313.5000 ;
	    RECT 937.8000 313.5000 950.7000 314.4000 ;
	    RECT 937.8000 313.2000 939.0000 313.5000 ;
	    RECT 925.5000 311.4000 929.4000 312.6000 ;
	    RECT 783.3000 303.3000 784.5000 309.3000 ;
	    RECT 916.2000 303.3000 917.4000 309.3000 ;
	    RECT 918.6000 303.3000 919.8000 310.5000 ;
	    RECT 920.7000 310.2000 924.6000 311.1000 ;
	    RECT 921.0000 303.3000 922.2000 309.3000 ;
	    RECT 923.4000 303.3000 924.6000 310.2000 ;
	    RECT 925.8000 303.3000 927.0000 309.3000 ;
	    RECT 928.2000 303.3000 929.4000 311.4000 ;
	    RECT 930.3000 310.2000 936.6000 311.4000 ;
	    RECT 930.6000 303.3000 931.8000 309.3000 ;
	    RECT 933.0000 303.3000 934.2000 307.5000 ;
	    RECT 935.4000 303.3000 936.6000 307.5000 ;
	    RECT 937.8000 303.3000 939.0000 307.5000 ;
	    RECT 940.2000 303.3000 941.4000 312.6000 ;
	    RECT 945.0000 311.4000 948.9000 312.6000 ;
	    RECT 949.8000 312.3000 950.7000 313.5000 ;
	    RECT 952.2000 314.1000 953.4000 314.4000 ;
	    RECT 952.2000 313.5000 960.3000 314.1000 ;
	    RECT 952.2000 313.2000 961.5000 313.5000 ;
	    RECT 959.4000 312.3000 961.5000 313.2000 ;
	    RECT 949.8000 311.4000 958.5000 312.3000 ;
	    RECT 963.0000 312.0000 965.4000 313.2000 ;
	    RECT 963.0000 311.4000 963.9000 312.0000 ;
	    RECT 942.6000 303.3000 943.8000 309.3000 ;
	    RECT 945.0000 303.3000 946.2000 310.5000 ;
	    RECT 947.4000 303.3000 948.6000 309.3000 ;
	    RECT 949.8000 303.3000 951.0000 310.5000 ;
	    RECT 957.6000 310.2000 963.9000 311.4000 ;
	    RECT 966.6000 311.1000 967.8000 319.5000 ;
	    RECT 1000.2000 319.2000 1001.4000 319.5000 ;
	    RECT 1004.7000 318.6000 1005.9000 319.5000 ;
	    RECT 969.0000 318.4500 970.2000 318.6000 ;
	    RECT 997.8000 318.4500 999.0000 318.6000 ;
	    RECT 969.0000 317.5500 999.0000 318.4500 ;
	    RECT 969.0000 317.4000 970.2000 317.5500 ;
	    RECT 997.8000 317.4000 999.0000 317.5500 ;
	    RECT 999.9000 316.8000 1000.2000 318.3000 ;
	    RECT 1002.6000 317.4000 1003.8000 318.6000 ;
	    RECT 1007.4000 318.4500 1008.6000 318.6000 ;
	    RECT 1014.6000 318.4500 1015.8000 318.6000 ;
	    RECT 1007.4000 317.5500 1015.8000 318.4500 ;
	    RECT 1007.4000 317.4000 1008.6000 317.5500 ;
	    RECT 1014.6000 317.4000 1015.8000 317.5500 ;
	    RECT 1033.8000 317.4000 1035.0000 318.6000 ;
	    RECT 1004.7000 316.5000 1005.9000 317.1000 ;
	    RECT 1035.9000 316.5000 1036.8000 321.6000 ;
	    RECT 1041.0000 321.4500 1042.2001 321.6000 ;
	    RECT 1050.6000 321.4500 1051.8000 321.6000 ;
	    RECT 1038.0000 320.7000 1039.2001 321.0000 ;
	    RECT 1038.0000 319.8000 1039.5000 320.7000 ;
	    RECT 1041.0000 320.5500 1051.8000 321.4500 ;
	    RECT 1067.4000 320.7000 1068.6000 329.7000 ;
	    RECT 1072.8000 321.3000 1074.0000 329.7000 ;
	    RECT 1077.0000 327.4500 1078.2001 327.6000 ;
	    RECT 1093.8000 327.4500 1095.0000 327.6000 ;
	    RECT 1077.0000 326.5500 1095.0000 327.4500 ;
	    RECT 1077.0000 326.4000 1078.2001 326.5500 ;
	    RECT 1093.8000 326.4000 1095.0000 326.5500 ;
	    RECT 1072.8000 320.7000 1075.5000 321.3000 ;
	    RECT 1098.6000 320.7000 1099.8000 329.7000 ;
	    RECT 1104.0000 321.3000 1105.2001 329.7000 ;
	    RECT 1133.1000 324.6000 1134.3000 329.7000 ;
	    RECT 1133.1000 323.7000 1135.8000 324.6000 ;
	    RECT 1137.0000 323.7000 1138.2001 329.7000 ;
	    RECT 1104.0000 320.7000 1106.7001 321.3000 ;
	    RECT 1041.0000 320.4000 1042.2001 320.5500 ;
	    RECT 1050.6000 320.4000 1051.8000 320.5500 ;
	    RECT 1073.1000 320.4000 1075.5000 320.7000 ;
	    RECT 1104.3000 320.4000 1106.7001 320.7000 ;
	    RECT 1038.6000 319.5000 1039.5000 319.8000 ;
	    RECT 1041.0000 319.2000 1042.2001 319.5000 ;
	    RECT 1038.6000 317.4000 1039.8000 318.6000 ;
	    RECT 1069.8000 317.4000 1071.0000 318.6000 ;
	    RECT 1071.9000 317.4000 1072.2001 318.6000 ;
	    RECT 1067.4000 316.5000 1068.6000 316.8000 ;
	    RECT 1074.6000 316.5000 1075.5000 320.4000 ;
	    RECT 1101.0000 317.4000 1102.2001 318.6000 ;
	    RECT 1103.1000 317.4000 1103.4000 318.6000 ;
	    RECT 1098.6000 316.5000 1099.8000 316.8000 ;
	    RECT 1105.8000 316.5000 1106.7001 320.4000 ;
	    RECT 1134.6000 319.5000 1135.8000 323.7000 ;
	    RECT 1137.0000 322.5000 1138.2001 322.8000 ;
	    RECT 1137.0000 321.4500 1138.2001 321.6000 ;
	    RECT 1158.6000 321.4500 1159.8000 321.6000 ;
	    RECT 1137.0000 320.5500 1159.8000 321.4500 ;
	    RECT 1165.2001 321.3000 1166.4000 329.7000 ;
	    RECT 1137.0000 320.4000 1138.2001 320.5500 ;
	    RECT 1158.6000 320.4000 1159.8000 320.5500 ;
	    RECT 1163.7001 320.7000 1166.4000 321.3000 ;
	    RECT 1170.6000 320.7000 1171.8000 329.7000 ;
	    RECT 1197.9000 323.7000 1199.1000 329.7000 ;
	    RECT 1201.8000 323.7000 1203.0000 329.7000 ;
	    RECT 1204.2001 326.7000 1205.4000 329.7000 ;
	    RECT 1203.9000 325.5000 1205.1000 325.8000 ;
	    RECT 1204.2001 324.4500 1205.4000 324.6000 ;
	    RECT 1211.4000 324.4500 1212.6000 324.6000 ;
	    RECT 1194.6000 321.4500 1195.8000 321.6000 ;
	    RECT 1199.4000 321.4500 1200.6000 321.6000 ;
	    RECT 1163.7001 320.4000 1166.1000 320.7000 ;
	    RECT 1194.6000 320.5500 1200.6000 321.4500 ;
	    RECT 1194.6000 320.4000 1195.8000 320.5500 ;
	    RECT 1199.4000 320.4000 1200.6000 320.5500 ;
	    RECT 1134.6000 318.4500 1135.8000 318.6000 ;
	    RECT 1149.0000 318.4500 1150.2001 318.6000 ;
	    RECT 1134.6000 317.5500 1150.2001 318.4500 ;
	    RECT 1134.6000 317.4000 1135.8000 317.5500 ;
	    RECT 1149.0000 317.4000 1150.2001 317.5500 ;
	    RECT 1163.7001 316.5000 1164.6000 320.4000 ;
	    RECT 1199.4000 319.2000 1200.6000 319.5000 ;
	    RECT 1167.0000 317.4000 1167.3000 318.6000 ;
	    RECT 1168.2001 317.4000 1169.4000 318.6000 ;
	    RECT 1189.8000 318.4500 1191.0000 318.6000 ;
	    RECT 1197.0000 318.4500 1198.2001 318.6000 ;
	    RECT 1189.8000 317.5500 1198.2001 318.4500 ;
	    RECT 1201.8000 318.3000 1202.7001 323.7000 ;
	    RECT 1204.2001 323.5500 1212.6000 324.4500 ;
	    RECT 1230.6000 323.7000 1231.8000 329.7000 ;
	    RECT 1234.5000 324.0000 1235.7001 329.7000 ;
	    RECT 1236.9000 325.2000 1238.1000 329.7000 ;
	    RECT 1236.9000 323.7000 1239.0000 325.2000 ;
	    RECT 1262.7001 323.7000 1263.9000 329.7000 ;
	    RECT 1266.6000 323.7000 1267.8000 329.7000 ;
	    RECT 1269.0000 326.7000 1270.2001 329.7000 ;
	    RECT 1268.7001 325.5000 1269.9000 325.8000 ;
	    RECT 1269.0000 324.4500 1270.2001 324.6000 ;
	    RECT 1285.8000 324.4500 1287.0000 324.6000 ;
	    RECT 1204.2001 323.4000 1205.4000 323.5500 ;
	    RECT 1211.4000 323.4000 1212.6000 323.5500 ;
	    RECT 1230.9000 323.4000 1231.8000 323.7000 ;
	    RECT 1230.9000 322.8000 1233.6000 323.4000 ;
	    RECT 1230.9000 322.5000 1237.2001 322.8000 ;
	    RECT 1232.7001 321.9000 1237.2001 322.5000 ;
	    RECT 1236.0000 321.6000 1237.2001 321.9000 ;
	    RECT 1225.8000 321.4500 1227.0000 321.6000 ;
	    RECT 1230.6000 321.4500 1231.8000 321.6000 ;
	    RECT 1225.8000 320.5500 1231.8000 321.4500 ;
	    RECT 1233.6000 320.7000 1234.8000 321.0000 ;
	    RECT 1225.8000 320.4000 1227.0000 320.5500 ;
	    RECT 1230.6000 320.4000 1231.8000 320.5500 ;
	    RECT 1233.3000 319.8000 1234.8000 320.7000 ;
	    RECT 1233.3000 319.5000 1234.2001 319.8000 ;
	    RECT 1230.6000 319.2000 1231.8000 319.5000 ;
	    RECT 1204.2001 318.4500 1205.4000 318.6000 ;
	    RECT 1221.0000 318.4500 1222.2001 318.6000 ;
	    RECT 1189.8000 317.4000 1191.0000 317.5500 ;
	    RECT 1197.0000 317.4000 1198.2001 317.5500 ;
	    RECT 1199.1000 316.8000 1199.4000 318.3000 ;
	    RECT 1201.8000 317.4000 1203.3000 318.3000 ;
	    RECT 1204.2001 317.5500 1222.2001 318.4500 ;
	    RECT 1204.2001 317.4000 1205.4000 317.5500 ;
	    RECT 1221.0000 317.4000 1222.2001 317.5500 ;
	    RECT 1233.0000 317.4000 1234.2001 318.6000 ;
	    RECT 1170.6000 316.5000 1171.8000 316.8000 ;
	    RECT 1236.0000 316.5000 1236.9000 321.6000 ;
	    RECT 1238.1000 319.5000 1239.0000 323.7000 ;
	    RECT 1254.6000 321.4500 1255.8000 321.6000 ;
	    RECT 1264.2001 321.4500 1265.4000 321.6000 ;
	    RECT 1254.6000 320.5500 1265.4000 321.4500 ;
	    RECT 1254.6000 320.4000 1255.8000 320.5500 ;
	    RECT 1264.2001 320.4000 1265.4000 320.5500 ;
	    RECT 1264.2001 319.2000 1265.4000 319.5000 ;
	    RECT 1237.8000 318.4500 1239.0000 318.6000 ;
	    RECT 1249.8000 318.4500 1251.0000 318.6000 ;
	    RECT 1237.8000 317.5500 1251.0000 318.4500 ;
	    RECT 1237.8000 317.4000 1239.0000 317.5500 ;
	    RECT 1249.8000 317.4000 1251.0000 317.5500 ;
	    RECT 1252.2001 318.4500 1253.4000 318.6000 ;
	    RECT 1261.8000 318.4500 1263.0000 318.6000 ;
	    RECT 1252.2001 317.5500 1263.0000 318.4500 ;
	    RECT 1266.6000 318.3000 1267.5000 323.7000 ;
	    RECT 1269.0000 323.5500 1287.0000 324.4500 ;
	    RECT 1293.0000 324.0000 1294.2001 329.7000 ;
	    RECT 1295.4000 324.9000 1296.6000 329.7000 ;
	    RECT 1297.8000 324.0000 1299.0000 329.7000 ;
	    RECT 1293.0000 323.7000 1299.0000 324.0000 ;
	    RECT 1300.2001 323.7000 1301.4000 329.7000 ;
	    RECT 1324.2001 324.0000 1325.4000 329.7000 ;
	    RECT 1326.6000 324.9000 1327.8000 329.7000 ;
	    RECT 1329.0000 324.0000 1330.2001 329.7000 ;
	    RECT 1324.2001 323.7000 1330.2001 324.0000 ;
	    RECT 1331.4000 323.7000 1332.6000 329.7000 ;
	    RECT 1363.5000 323.7000 1364.7001 329.7000 ;
	    RECT 1367.4000 323.7000 1368.6000 329.7000 ;
	    RECT 1369.8000 326.7000 1371.0000 329.7000 ;
	    RECT 1369.5000 325.5000 1370.7001 325.8000 ;
	    RECT 1369.8000 324.4500 1371.0000 324.6000 ;
	    RECT 1389.0000 324.4500 1390.2001 324.6000 ;
	    RECT 1269.0000 323.4000 1270.2001 323.5500 ;
	    RECT 1285.8000 323.4000 1287.0000 323.5500 ;
	    RECT 1293.3000 323.1000 1298.7001 323.7000 ;
	    RECT 1300.2001 322.5000 1301.1000 323.7000 ;
	    RECT 1324.5000 323.1000 1329.9000 323.7000 ;
	    RECT 1331.4000 322.5000 1332.3000 323.7000 ;
	    RECT 1293.0000 320.4000 1294.2001 321.6000 ;
	    RECT 1295.1000 320.7000 1295.4000 322.2000 ;
	    RECT 1297.5000 320.4000 1299.3000 321.6000 ;
	    RECT 1300.2001 321.4500 1301.4000 321.6000 ;
	    RECT 1319.4000 321.4500 1320.6000 321.6000 ;
	    RECT 1300.2001 320.5500 1320.6000 321.4500 ;
	    RECT 1300.2001 320.4000 1301.4000 320.5500 ;
	    RECT 1319.4000 320.4000 1320.6000 320.5500 ;
	    RECT 1324.2001 320.4000 1325.4000 321.6000 ;
	    RECT 1326.3000 320.7000 1326.6000 322.2000 ;
	    RECT 1328.7001 320.4000 1330.5000 321.6000 ;
	    RECT 1331.4000 321.4500 1332.6000 321.6000 ;
	    RECT 1362.6000 321.4500 1363.8000 321.6000 ;
	    RECT 1365.0000 321.4500 1366.2001 321.6000 ;
	    RECT 1331.4000 320.5500 1361.2500 321.4500 ;
	    RECT 1331.4000 320.4000 1332.6000 320.5500 ;
	    RECT 1295.4000 319.5000 1296.6000 319.8000 ;
	    RECT 1269.0000 318.4500 1270.2001 318.6000 ;
	    RECT 1271.4000 318.4500 1272.6000 318.6000 ;
	    RECT 1252.2001 317.4000 1253.4000 317.5500 ;
	    RECT 1261.8000 317.4000 1263.0000 317.5500 ;
	    RECT 1263.9000 316.8000 1264.2001 318.3000 ;
	    RECT 1266.6000 317.4000 1268.1000 318.3000 ;
	    RECT 1269.0000 317.5500 1272.6000 318.4500 ;
	    RECT 1269.0000 317.4000 1270.2001 317.5500 ;
	    RECT 1271.4000 317.4000 1272.6000 317.5500 ;
	    RECT 1273.8000 318.4500 1275.0000 318.6000 ;
	    RECT 1295.4000 318.4500 1296.6000 318.6000 ;
	    RECT 1273.8000 317.5500 1296.6000 318.4500 ;
	    RECT 1273.8000 317.4000 1275.0000 317.5500 ;
	    RECT 1295.4000 317.4000 1296.6000 317.5500 ;
	    RECT 1002.9000 316.2000 1005.9000 316.5000 ;
	    RECT 1007.4000 316.2000 1008.6000 316.5000 ;
	    RECT 1005.0000 315.3000 1005.9000 316.2000 ;
	    RECT 1033.8000 315.3000 1034.7001 316.5000 ;
	    RECT 1035.9000 315.6000 1039.5000 316.5000 ;
	    RECT 964.8000 310.2000 967.8000 311.1000 ;
	    RECT 997.8000 314.4000 1003.8000 315.3000 ;
	    RECT 952.2000 303.3000 953.4000 307.5000 ;
	    RECT 954.6000 303.3000 955.8000 307.5000 ;
	    RECT 957.0000 303.3000 958.2000 309.3000 ;
	    RECT 959.4000 303.3000 960.6000 310.2000 ;
	    RECT 964.8000 309.3000 965.7000 310.2000 ;
	    RECT 961.8000 302.4000 963.0000 309.3000 ;
	    RECT 964.2000 308.4000 965.7000 309.3000 ;
	    RECT 964.2000 303.3000 965.4000 308.4000 ;
	    RECT 966.6000 303.3000 967.8000 309.3000 ;
	    RECT 997.8000 303.3000 999.0000 314.4000 ;
	    RECT 1000.2000 303.3000 1001.4000 313.5000 ;
	    RECT 1002.6000 304.2000 1003.8000 314.4000 ;
	    RECT 1005.0000 305.1000 1006.2000 315.3000 ;
	    RECT 1007.4000 304.2000 1008.6000 315.3000 ;
	    RECT 1002.6000 303.3000 1008.6000 304.2000 ;
	    RECT 1033.8000 303.3000 1035.0000 315.3000 ;
	    RECT 1036.2001 303.3000 1037.4000 314.7000 ;
	    RECT 1038.6000 309.3000 1039.5000 315.6000 ;
	    RECT 1043.4000 315.4500 1044.6000 315.6000 ;
	    RECT 1062.6000 315.4500 1063.8000 315.6000 ;
	    RECT 1067.4000 315.4500 1068.6000 315.6000 ;
	    RECT 1043.4000 314.5500 1068.6000 315.4500 ;
	    RECT 1043.4000 314.4000 1044.6000 314.5500 ;
	    RECT 1062.6000 314.4000 1063.8000 314.5500 ;
	    RECT 1067.4000 314.4000 1068.6000 314.5500 ;
	    RECT 1074.6000 315.4500 1075.8000 315.6000 ;
	    RECT 1096.2001 315.4500 1097.4000 315.6000 ;
	    RECT 1098.6000 315.4500 1099.8000 315.6000 ;
	    RECT 1074.6000 314.5500 1094.8500 315.4500 ;
	    RECT 1074.6000 314.4000 1075.8000 314.5500 ;
	    RECT 1072.2001 313.5000 1073.4000 313.8000 ;
	    RECT 1072.2001 311.4000 1073.4000 312.6000 ;
	    RECT 1074.6000 310.5000 1075.5000 313.5000 ;
	    RECT 1093.9501 312.4500 1094.8500 314.5500 ;
	    RECT 1096.2001 314.5500 1099.8000 315.4500 ;
	    RECT 1096.2001 314.4000 1097.4000 314.5500 ;
	    RECT 1098.6000 314.4000 1099.8000 314.5500 ;
	    RECT 1105.8000 315.4500 1107.0000 315.6000 ;
	    RECT 1129.8000 315.4500 1131.0000 315.6000 ;
	    RECT 1105.8000 314.5500 1131.0000 315.4500 ;
	    RECT 1105.8000 314.4000 1107.0000 314.5500 ;
	    RECT 1129.8000 314.4000 1131.0000 314.5500 ;
	    RECT 1132.2001 314.4000 1133.4000 315.6000 ;
	    RECT 1103.4000 313.5000 1104.6000 313.8000 ;
	    RECT 1101.0000 312.4500 1102.2001 312.6000 ;
	    RECT 1103.4000 312.4500 1104.6000 312.6000 ;
	    RECT 1093.9501 311.5500 1104.6000 312.4500 ;
	    RECT 1101.0000 311.4000 1102.2001 311.5500 ;
	    RECT 1103.4000 311.4000 1104.6000 311.5500 ;
	    RECT 1105.8000 310.5000 1106.7001 313.5000 ;
	    RECT 1132.2001 313.2000 1133.4000 313.5000 ;
	    RECT 1070.1000 309.6000 1075.5000 310.5000 ;
	    RECT 1070.1000 309.3000 1071.0000 309.6000 ;
	    RECT 1038.6000 303.3000 1039.8000 309.3000 ;
	    RECT 1041.0000 303.3000 1042.2001 309.3000 ;
	    RECT 1067.4000 303.3000 1068.6000 309.3000 ;
	    RECT 1069.8000 303.3000 1071.0000 309.3000 ;
	    RECT 1074.6000 309.3000 1075.5000 309.6000 ;
	    RECT 1101.3000 309.6000 1106.7001 310.5000 ;
	    RECT 1101.3000 309.3000 1102.2001 309.6000 ;
	    RECT 1072.2001 303.3000 1073.4000 308.7000 ;
	    RECT 1074.6000 303.3000 1075.8000 309.3000 ;
	    RECT 1098.6000 303.3000 1099.8000 309.3000 ;
	    RECT 1101.0000 303.3000 1102.2001 309.3000 ;
	    RECT 1105.8000 309.3000 1106.7001 309.6000 ;
	    RECT 1103.4000 303.3000 1104.6000 308.7000 ;
	    RECT 1105.8000 303.3000 1107.0000 309.3000 ;
	    RECT 1132.2001 303.3000 1133.4000 309.3000 ;
	    RECT 1134.6000 303.3000 1135.8000 316.5000 ;
	    RECT 1163.4000 314.4000 1164.6000 315.6000 ;
	    RECT 1170.6000 314.4000 1171.8000 315.6000 ;
	    RECT 1204.2001 315.3000 1205.1000 316.5000 ;
	    RECT 1233.3000 315.6000 1236.9000 316.5000 ;
	    RECT 1197.0000 314.4000 1203.0000 315.3000 ;
	    RECT 1165.8000 313.5000 1167.0000 313.8000 ;
	    RECT 1163.7001 310.5000 1164.6000 313.5000 ;
	    RECT 1165.8000 311.4000 1167.0000 312.6000 ;
	    RECT 1168.2001 312.4500 1169.4000 312.6000 ;
	    RECT 1187.4000 312.4500 1188.6000 312.6000 ;
	    RECT 1194.6000 312.4500 1195.8000 312.6000 ;
	    RECT 1168.2001 311.5500 1195.8000 312.4500 ;
	    RECT 1168.2001 311.4000 1169.4000 311.5500 ;
	    RECT 1187.4000 311.4000 1188.6000 311.5500 ;
	    RECT 1194.6000 311.4000 1195.8000 311.5500 ;
	    RECT 1163.7001 309.6000 1169.1000 310.5000 ;
	    RECT 1163.7001 309.3000 1164.6000 309.6000 ;
	    RECT 1137.0000 303.3000 1138.2001 309.3000 ;
	    RECT 1163.4000 303.3000 1164.6000 309.3000 ;
	    RECT 1168.2001 309.3000 1169.1000 309.6000 ;
	    RECT 1165.8000 303.3000 1167.0000 308.7000 ;
	    RECT 1168.2001 303.3000 1169.4000 309.3000 ;
	    RECT 1170.6000 303.3000 1171.8000 309.3000 ;
	    RECT 1197.0000 303.3000 1198.2001 314.4000 ;
	    RECT 1199.4000 303.3000 1200.6000 313.5000 ;
	    RECT 1201.8000 303.3000 1203.0000 314.4000 ;
	    RECT 1204.2001 303.3000 1205.4000 315.3000 ;
	    RECT 1233.3000 309.3000 1234.2001 315.6000 ;
	    RECT 1238.1000 315.3000 1239.0000 316.5000 ;
	    RECT 1269.0000 315.3000 1269.9000 316.5000 ;
	    RECT 1297.5000 315.3000 1298.4000 320.4000 ;
	    RECT 1326.6000 319.5000 1327.8000 319.8000 ;
	    RECT 1305.0000 318.4500 1306.2001 318.6000 ;
	    RECT 1326.6000 318.4500 1327.8000 318.6000 ;
	    RECT 1305.0000 317.5500 1327.8000 318.4500 ;
	    RECT 1305.0000 317.4000 1306.2001 317.5500 ;
	    RECT 1326.6000 317.4000 1327.8000 317.5500 ;
	    RECT 1230.6000 303.3000 1231.8000 309.3000 ;
	    RECT 1233.0000 303.3000 1234.2001 309.3000 ;
	    RECT 1235.4000 303.3000 1236.6000 314.7000 ;
	    RECT 1237.8000 303.3000 1239.0000 315.3000 ;
	    RECT 1261.8000 314.4000 1267.8000 315.3000 ;
	    RECT 1261.8000 303.3000 1263.0000 314.4000 ;
	    RECT 1264.2001 303.3000 1265.4000 313.5000 ;
	    RECT 1266.6000 303.3000 1267.8000 314.4000 ;
	    RECT 1269.0000 303.3000 1270.2001 315.3000 ;
	    RECT 1293.0000 303.3000 1294.2001 315.3000 ;
	    RECT 1296.9000 314.4000 1298.4000 315.3000 ;
	    RECT 1300.2001 315.4500 1301.4000 315.6000 ;
	    RECT 1309.8000 315.4500 1311.0000 315.6000 ;
	    RECT 1300.2001 314.5500 1311.0000 315.4500 ;
	    RECT 1328.7001 315.3000 1329.6000 320.4000 ;
	    RECT 1360.3500 318.4500 1361.2500 320.5500 ;
	    RECT 1362.6000 320.5500 1366.2001 321.4500 ;
	    RECT 1362.6000 320.4000 1363.8000 320.5500 ;
	    RECT 1365.0000 320.4000 1366.2001 320.5500 ;
	    RECT 1365.0000 319.2000 1366.2001 319.5000 ;
	    RECT 1362.6000 318.4500 1363.8000 318.6000 ;
	    RECT 1360.3500 317.5500 1363.8000 318.4500 ;
	    RECT 1367.4000 318.3000 1368.3000 323.7000 ;
	    RECT 1369.8000 323.5500 1390.2001 324.4500 ;
	    RECT 1393.8000 324.0000 1395.0000 329.7000 ;
	    RECT 1396.2001 324.9000 1397.4000 329.7000 ;
	    RECT 1398.6000 324.0000 1399.8000 329.7000 ;
	    RECT 1393.8000 323.7000 1399.8000 324.0000 ;
	    RECT 1401.0000 323.7000 1402.2001 329.7000 ;
	    RECT 1369.8000 323.4000 1371.0000 323.5500 ;
	    RECT 1389.0000 323.4000 1390.2001 323.5500 ;
	    RECT 1394.1000 323.1000 1399.5000 323.7000 ;
	    RECT 1401.0000 322.5000 1401.9000 323.7000 ;
	    RECT 1393.8000 320.4000 1395.0000 321.6000 ;
	    RECT 1395.9000 320.7000 1396.2001 322.2000 ;
	    RECT 1398.3000 320.4000 1400.1000 321.6000 ;
	    RECT 1401.0000 321.4500 1402.2001 321.6000 ;
	    RECT 1422.6000 321.4500 1423.8000 321.6000 ;
	    RECT 1401.0000 320.5500 1423.8000 321.4500 ;
	    RECT 1425.0000 320.7000 1426.2001 329.7000 ;
	    RECT 1430.4000 321.3000 1431.6000 329.7000 ;
	    RECT 1458.0000 321.3000 1459.2001 329.7000 ;
	    RECT 1430.4000 320.7000 1433.1000 321.3000 ;
	    RECT 1401.0000 320.4000 1402.2001 320.5500 ;
	    RECT 1422.6000 320.4000 1423.8000 320.5500 ;
	    RECT 1430.7001 320.4000 1433.1000 320.7000 ;
	    RECT 1396.2001 319.5000 1397.4000 319.8000 ;
	    RECT 1369.8000 318.4500 1371.0000 318.6000 ;
	    RECT 1391.4000 318.4500 1392.6000 318.6000 ;
	    RECT 1362.6000 317.4000 1363.8000 317.5500 ;
	    RECT 1364.7001 316.8000 1365.0000 318.3000 ;
	    RECT 1367.4000 317.4000 1368.9000 318.3000 ;
	    RECT 1369.8000 317.5500 1392.6000 318.4500 ;
	    RECT 1369.8000 317.4000 1371.0000 317.5500 ;
	    RECT 1391.4000 317.4000 1392.6000 317.5500 ;
	    RECT 1396.2001 317.4000 1397.4000 318.6000 ;
	    RECT 1300.2001 314.4000 1301.4000 314.5500 ;
	    RECT 1309.8000 314.4000 1311.0000 314.5500 ;
	    RECT 1296.9000 303.3000 1298.1000 314.4000 ;
	    RECT 1299.3000 312.6000 1300.2001 313.5000 ;
	    RECT 1299.0000 311.4000 1300.2001 312.6000 ;
	    RECT 1299.3000 303.3000 1300.5000 309.3000 ;
	    RECT 1324.2001 303.3000 1325.4000 315.3000 ;
	    RECT 1328.1000 314.4000 1329.6000 315.3000 ;
	    RECT 1331.4000 315.4500 1332.6000 315.6000 ;
	    RECT 1333.8000 315.4500 1335.0000 315.6000 ;
	    RECT 1331.4000 314.5500 1335.0000 315.4500 ;
	    RECT 1369.8000 315.3000 1370.7001 316.5000 ;
	    RECT 1398.3000 315.3000 1399.2001 320.4000 ;
	    RECT 1427.4000 317.4000 1428.6000 318.6000 ;
	    RECT 1429.5000 317.4000 1429.8000 318.6000 ;
	    RECT 1425.0000 316.5000 1426.2001 316.8000 ;
	    RECT 1432.2001 316.5000 1433.1000 320.4000 ;
	    RECT 1456.5000 320.7000 1459.2001 321.3000 ;
	    RECT 1463.4000 320.7000 1464.6000 329.7000 ;
	    RECT 1487.4000 320.7000 1488.6000 329.7000 ;
	    RECT 1492.8000 321.3000 1494.0000 329.7000 ;
	    RECT 1514.7001 324.6000 1515.9000 329.7000 ;
	    RECT 1514.7001 323.7000 1517.4000 324.6000 ;
	    RECT 1518.6000 323.7000 1519.8000 329.7000 ;
	    RECT 1542.6000 323.7000 1543.8000 329.7000 ;
	    RECT 1545.0000 324.0000 1546.2001 329.7000 ;
	    RECT 1547.4000 324.9000 1548.6000 329.7000 ;
	    RECT 1549.8000 324.0000 1551.0000 329.7000 ;
	    RECT 1545.0000 323.7000 1551.0000 324.0000 ;
	    RECT 1492.8000 320.7000 1495.5000 321.3000 ;
	    RECT 1456.5000 320.4000 1458.9000 320.7000 ;
	    RECT 1493.1000 320.4000 1495.5000 320.7000 ;
	    RECT 1456.5000 316.5000 1457.4000 320.4000 ;
	    RECT 1459.8000 317.4000 1460.1000 318.6000 ;
	    RECT 1461.0000 317.4000 1462.2001 318.6000 ;
	    RECT 1489.8000 317.4000 1491.0000 318.6000 ;
	    RECT 1491.9000 317.4000 1492.2001 318.6000 ;
	    RECT 1463.4000 316.5000 1464.6000 316.8000 ;
	    RECT 1487.4000 316.5000 1488.6000 316.8000 ;
	    RECT 1494.6000 316.5000 1495.5000 320.4000 ;
	    RECT 1516.2001 319.5000 1517.4000 323.7000 ;
	    RECT 1518.6000 322.5000 1519.8000 322.8000 ;
	    RECT 1542.9000 322.5000 1543.8000 323.7000 ;
	    RECT 1545.3000 323.1000 1550.7001 323.7000 ;
	    RECT 1518.6000 321.4500 1519.8000 321.6000 ;
	    RECT 1521.0000 321.4500 1522.2001 321.6000 ;
	    RECT 1540.2001 321.4500 1541.4000 321.6000 ;
	    RECT 1518.6000 320.5500 1541.4000 321.4500 ;
	    RECT 1518.6000 320.4000 1519.8000 320.5500 ;
	    RECT 1521.0000 320.4000 1522.2001 320.5500 ;
	    RECT 1540.2001 320.4000 1541.4000 320.5500 ;
	    RECT 1542.6000 320.4000 1543.8000 321.6000 ;
	    RECT 1544.7001 320.4000 1546.5000 321.6000 ;
	    RECT 1548.6000 320.7000 1548.9000 322.2000 ;
	    RECT 1549.8000 321.4500 1551.0000 321.6000 ;
	    RECT 1554.6000 321.4500 1555.8000 321.6000 ;
	    RECT 1549.8000 320.5500 1555.8000 321.4500 ;
	    RECT 1549.8000 320.4000 1551.0000 320.5500 ;
	    RECT 1554.6000 320.4000 1555.8000 320.5500 ;
	    RECT 1516.2001 318.4500 1517.4000 318.6000 ;
	    RECT 1535.4000 318.4500 1536.6000 318.6000 ;
	    RECT 1542.6000 318.4500 1543.8000 318.6000 ;
	    RECT 1516.2001 317.5500 1543.8000 318.4500 ;
	    RECT 1516.2001 317.4000 1517.4000 317.5500 ;
	    RECT 1535.4000 317.4000 1536.6000 317.5500 ;
	    RECT 1542.6000 317.4000 1543.8000 317.5500 ;
	    RECT 1331.4000 314.4000 1332.6000 314.5500 ;
	    RECT 1333.8000 314.4000 1335.0000 314.5500 ;
	    RECT 1362.6000 314.4000 1368.6000 315.3000 ;
	    RECT 1328.1000 303.3000 1329.3000 314.4000 ;
	    RECT 1330.5000 312.6000 1331.4000 313.5000 ;
	    RECT 1330.2001 311.4000 1331.4000 312.6000 ;
	    RECT 1330.5000 303.3000 1331.7001 309.3000 ;
	    RECT 1362.6000 303.3000 1363.8000 314.4000 ;
	    RECT 1365.0000 303.3000 1366.2001 313.5000 ;
	    RECT 1367.4000 303.3000 1368.6000 314.4000 ;
	    RECT 1369.8000 303.3000 1371.0000 315.3000 ;
	    RECT 1393.8000 303.3000 1395.0000 315.3000 ;
	    RECT 1397.7001 314.4000 1399.2001 315.3000 ;
	    RECT 1401.0000 314.4000 1402.2001 315.6000 ;
	    RECT 1420.2001 315.4500 1421.4000 315.6000 ;
	    RECT 1425.0000 315.4500 1426.2001 315.6000 ;
	    RECT 1420.2001 314.5500 1426.2001 315.4500 ;
	    RECT 1420.2001 314.4000 1421.4000 314.5500 ;
	    RECT 1425.0000 314.4000 1426.2001 314.5500 ;
	    RECT 1432.2001 315.4500 1433.4000 315.6000 ;
	    RECT 1439.4000 315.4500 1440.6000 315.6000 ;
	    RECT 1432.2001 314.5500 1440.6000 315.4500 ;
	    RECT 1432.2001 314.4000 1433.4000 314.5500 ;
	    RECT 1439.4000 314.4000 1440.6000 314.5500 ;
	    RECT 1456.2001 314.4000 1457.4000 315.6000 ;
	    RECT 1463.4000 314.4000 1464.6000 315.6000 ;
	    RECT 1477.8000 315.4500 1479.0000 315.6000 ;
	    RECT 1482.6000 315.4500 1483.8000 315.6000 ;
	    RECT 1487.4000 315.4500 1488.6000 315.6000 ;
	    RECT 1477.8000 314.5500 1488.6000 315.4500 ;
	    RECT 1477.8000 314.4000 1479.0000 314.5500 ;
	    RECT 1482.6000 314.4000 1483.8000 314.5500 ;
	    RECT 1487.4000 314.4000 1488.6000 314.5500 ;
	    RECT 1494.6000 315.4500 1495.8000 315.6000 ;
	    RECT 1509.0000 315.4500 1510.2001 315.6000 ;
	    RECT 1494.6000 314.5500 1510.2001 315.4500 ;
	    RECT 1494.6000 314.4000 1495.8000 314.5500 ;
	    RECT 1509.0000 314.4000 1510.2001 314.5500 ;
	    RECT 1511.4000 315.4500 1512.6000 315.6000 ;
	    RECT 1513.8000 315.4500 1515.0000 315.6000 ;
	    RECT 1511.4000 314.5500 1515.0000 315.4500 ;
	    RECT 1511.4000 314.4000 1512.6000 314.5500 ;
	    RECT 1513.8000 314.4000 1515.0000 314.5500 ;
	    RECT 1397.7001 303.3000 1398.9000 314.4000 ;
	    RECT 1429.8000 313.5000 1431.0000 313.8000 ;
	    RECT 1458.6000 313.5000 1459.8000 313.8000 ;
	    RECT 1492.2001 313.5000 1493.4000 313.8000 ;
	    RECT 1400.1000 312.6000 1401.0000 313.5000 ;
	    RECT 1399.8000 311.4000 1401.0000 312.6000 ;
	    RECT 1429.8000 311.4000 1431.0000 312.6000 ;
	    RECT 1432.2001 310.5000 1433.1000 313.5000 ;
	    RECT 1437.0000 312.4500 1438.2001 312.6000 ;
	    RECT 1453.8000 312.4500 1455.0000 312.6000 ;
	    RECT 1437.0000 311.5500 1455.0000 312.4500 ;
	    RECT 1437.0000 311.4000 1438.2001 311.5500 ;
	    RECT 1453.8000 311.4000 1455.0000 311.5500 ;
	    RECT 1427.7001 309.6000 1433.1000 310.5000 ;
	    RECT 1427.7001 309.3000 1428.6000 309.6000 ;
	    RECT 1400.1000 303.3000 1401.3000 309.3000 ;
	    RECT 1425.0000 303.3000 1426.2001 309.3000 ;
	    RECT 1427.4000 303.3000 1428.6000 309.3000 ;
	    RECT 1432.2001 309.3000 1433.1000 309.6000 ;
	    RECT 1456.5000 310.5000 1457.4000 313.5000 ;
	    RECT 1458.6000 311.4000 1459.8000 312.6000 ;
	    RECT 1492.2001 311.4000 1493.4000 312.6000 ;
	    RECT 1494.6000 310.5000 1495.5000 313.5000 ;
	    RECT 1513.8000 313.2000 1515.0000 313.5000 ;
	    RECT 1456.5000 309.6000 1461.9000 310.5000 ;
	    RECT 1456.5000 309.3000 1457.4000 309.6000 ;
	    RECT 1429.8000 303.3000 1431.0000 308.7000 ;
	    RECT 1432.2001 303.3000 1433.4000 309.3000 ;
	    RECT 1449.0000 306.4500 1450.2001 306.6000 ;
	    RECT 1453.8000 306.4500 1455.0000 306.6000 ;
	    RECT 1449.0000 305.5500 1455.0000 306.4500 ;
	    RECT 1449.0000 305.4000 1450.2001 305.5500 ;
	    RECT 1453.8000 305.4000 1455.0000 305.5500 ;
	    RECT 1456.2001 303.3000 1457.4000 309.3000 ;
	    RECT 1461.0000 309.3000 1461.9000 309.6000 ;
	    RECT 1490.1000 309.6000 1495.5000 310.5000 ;
	    RECT 1490.1000 309.3000 1491.0000 309.6000 ;
	    RECT 1458.6000 303.3000 1459.8000 308.7000 ;
	    RECT 1461.0000 303.3000 1462.2001 309.3000 ;
	    RECT 1463.4000 303.3000 1464.6000 309.3000 ;
	    RECT 1487.4000 303.3000 1488.6000 309.3000 ;
	    RECT 1489.8000 303.3000 1491.0000 309.3000 ;
	    RECT 1494.6000 309.3000 1495.5000 309.6000 ;
	    RECT 1492.2001 303.3000 1493.4000 308.7000 ;
	    RECT 1494.6000 303.3000 1495.8000 309.3000 ;
	    RECT 1513.8000 303.3000 1515.0000 309.3000 ;
	    RECT 1516.2001 303.3000 1517.4000 316.5000 ;
	    RECT 1518.6000 315.4500 1519.8000 315.6000 ;
	    RECT 1542.6000 315.4500 1543.8000 315.6000 ;
	    RECT 1518.6000 314.5500 1543.8000 315.4500 ;
	    RECT 1518.6000 314.4000 1519.8000 314.5500 ;
	    RECT 1542.6000 314.4000 1543.8000 314.5500 ;
	    RECT 1545.6000 315.3000 1546.5000 320.4000 ;
	    RECT 1547.4000 319.5000 1548.6000 319.8000 ;
	    RECT 1547.4000 318.4500 1548.6000 318.6000 ;
	    RECT 1552.2001 318.4500 1553.4000 318.6000 ;
	    RECT 1547.4000 317.5500 1553.4000 318.4500 ;
	    RECT 1547.4000 317.4000 1548.6000 317.5500 ;
	    RECT 1552.2001 317.4000 1553.4000 317.5500 ;
	    RECT 1545.6000 314.4000 1547.1000 315.3000 ;
	    RECT 1543.8000 312.6000 1544.7001 313.5000 ;
	    RECT 1543.8000 311.4000 1545.0000 312.6000 ;
	    RECT 1518.6000 303.3000 1519.8000 309.3000 ;
	    RECT 1543.5000 303.3000 1544.7001 309.3000 ;
	    RECT 1545.9000 303.3000 1547.1000 314.4000 ;
	    RECT 1549.8000 303.3000 1551.0000 315.3000 ;
	    RECT 1.2000 300.6000 1569.0000 302.4000 ;
	    RECT 23.4000 287.7000 24.6000 299.7000 ;
	    RECT 27.3000 288.6000 28.5000 299.7000 ;
	    RECT 29.7000 293.7000 30.9000 299.7000 ;
	    RECT 157.8000 293.7000 159.0000 299.7000 ;
	    RECT 160.2000 294.6000 161.4000 299.7000 ;
	    RECT 159.9000 293.7000 161.4000 294.6000 ;
	    RECT 162.6000 293.7000 163.8000 300.6000 ;
	    RECT 159.9000 292.8000 160.8000 293.7000 ;
	    RECT 165.0000 292.8000 166.2000 299.7000 ;
	    RECT 167.4000 293.7000 168.6000 299.7000 ;
	    RECT 169.8000 295.5000 171.0000 299.7000 ;
	    RECT 172.2000 295.5000 173.4000 299.7000 ;
	    RECT 157.8000 291.9000 160.8000 292.8000 ;
	    RECT 29.4000 290.4000 30.6000 291.6000 ;
	    RECT 29.7000 289.5000 30.6000 290.4000 ;
	    RECT 27.3000 287.7000 28.8000 288.6000 ;
	    RECT 25.8000 284.4000 27.0000 285.6000 ;
	    RECT 25.8000 283.2000 27.0000 283.5000 ;
	    RECT 27.9000 282.6000 28.8000 287.7000 ;
	    RECT 30.6000 287.4000 31.8000 288.6000 ;
	    RECT 157.8000 283.5000 159.0000 291.9000 ;
	    RECT 161.7000 291.6000 168.0000 292.8000 ;
	    RECT 174.6000 292.5000 175.8000 299.7000 ;
	    RECT 177.0000 293.7000 178.2000 299.7000 ;
	    RECT 179.4000 292.5000 180.6000 299.7000 ;
	    RECT 181.8000 293.7000 183.0000 299.7000 ;
	    RECT 161.7000 291.0000 162.6000 291.6000 ;
	    RECT 160.2000 289.8000 162.6000 291.0000 ;
	    RECT 167.1000 290.7000 175.8000 291.6000 ;
	    RECT 164.1000 289.8000 166.2000 290.7000 ;
	    RECT 164.1000 289.5000 173.4000 289.8000 ;
	    RECT 165.3000 288.9000 173.4000 289.5000 ;
	    RECT 172.2000 288.6000 173.4000 288.9000 ;
	    RECT 174.9000 289.5000 175.8000 290.7000 ;
	    RECT 176.7000 290.4000 180.6000 291.6000 ;
	    RECT 184.2000 290.4000 185.4000 299.7000 ;
	    RECT 186.6000 295.5000 187.8000 299.7000 ;
	    RECT 189.0000 295.5000 190.2000 299.7000 ;
	    RECT 191.4000 295.5000 192.6000 299.7000 ;
	    RECT 193.8000 293.7000 195.0000 299.7000 ;
	    RECT 189.0000 291.6000 195.3000 292.8000 ;
	    RECT 196.2000 291.6000 197.4000 299.7000 ;
	    RECT 198.6000 293.7000 199.8000 299.7000 ;
	    RECT 201.0000 292.8000 202.2000 299.7000 ;
	    RECT 203.4000 293.7000 204.6000 299.7000 ;
	    RECT 201.0000 291.9000 204.9000 292.8000 ;
	    RECT 205.8000 292.5000 207.0000 299.7000 ;
	    RECT 208.2000 293.7000 209.4000 299.7000 ;
	    RECT 340.2000 293.7000 341.4000 299.7000 ;
	    RECT 342.6000 294.6000 343.8000 299.7000 ;
	    RECT 342.3000 293.7000 343.8000 294.6000 ;
	    RECT 345.0000 293.7000 346.2000 300.6000 ;
	    RECT 342.3000 292.8000 343.2000 293.7000 ;
	    RECT 347.4000 292.8000 348.6000 299.7000 ;
	    RECT 349.8000 293.7000 351.0000 299.7000 ;
	    RECT 352.2000 295.5000 353.4000 299.7000 ;
	    RECT 354.6000 295.5000 355.8000 299.7000 ;
	    RECT 196.2000 290.4000 200.1000 291.6000 ;
	    RECT 186.6000 289.5000 187.8000 289.8000 ;
	    RECT 174.9000 288.6000 187.8000 289.5000 ;
	    RECT 191.4000 289.5000 192.6000 289.8000 ;
	    RECT 204.0000 289.5000 204.9000 291.9000 ;
	    RECT 340.2000 291.9000 343.2000 292.8000 ;
	    RECT 205.8000 290.4000 207.0000 291.6000 ;
	    RECT 191.4000 288.6000 204.9000 289.5000 ;
	    RECT 162.6000 287.4000 163.8000 288.6000 ;
	    RECT 167.7000 287.7000 168.9000 288.0000 ;
	    RECT 164.7000 286.8000 203.1000 287.7000 ;
	    RECT 201.9000 286.5000 203.1000 286.8000 ;
	    RECT 204.0000 285.9000 204.9000 288.6000 ;
	    RECT 205.8000 288.0000 207.0000 289.5000 ;
	    RECT 205.8000 286.8000 207.3000 288.0000 ;
	    RECT 159.9000 285.0000 166.5000 285.9000 ;
	    RECT 159.9000 284.7000 161.1000 285.0000 ;
	    RECT 167.4000 284.4000 168.6000 285.6000 ;
	    RECT 169.5000 285.0000 195.0000 285.9000 ;
	    RECT 204.0000 285.0000 205.2000 285.9000 ;
	    RECT 193.8000 284.1000 195.0000 285.0000 ;
	    RECT 18.6000 282.4500 19.8000 282.6000 ;
	    RECT 23.4000 282.4500 24.6000 282.6000 ;
	    RECT 18.6000 281.5500 24.6000 282.4500 ;
	    RECT 18.6000 281.4000 19.8000 281.5500 ;
	    RECT 23.4000 281.4000 24.6000 281.5500 ;
	    RECT 25.5000 280.8000 25.8000 282.3000 ;
	    RECT 27.9000 281.4000 29.7000 282.6000 ;
	    RECT 30.6000 282.4500 31.8000 282.6000 ;
	    RECT 143.4000 282.4500 144.6000 282.6000 ;
	    RECT 30.6000 281.5500 144.6000 282.4500 ;
	    RECT 30.6000 281.4000 31.8000 281.5500 ;
	    RECT 143.4000 281.4000 144.6000 281.5500 ;
	    RECT 157.8000 282.3000 171.0000 283.5000 ;
	    RECT 171.9000 282.9000 174.9000 284.1000 ;
	    RECT 180.6000 282.9000 185.4000 284.1000 ;
	    RECT 23.7000 279.3000 29.1000 279.9000 ;
	    RECT 30.6000 279.3000 31.5000 280.5000 ;
	    RECT 23.4000 279.0000 29.4000 279.3000 ;
	    RECT 23.4000 273.3000 24.6000 279.0000 ;
	    RECT 25.8000 273.3000 27.0000 278.1000 ;
	    RECT 28.2000 273.3000 29.4000 279.0000 ;
	    RECT 30.6000 273.3000 31.8000 279.3000 ;
	    RECT 157.8000 273.3000 159.0000 282.3000 ;
	    RECT 161.4000 280.2000 165.9000 281.4000 ;
	    RECT 164.7000 279.3000 165.9000 280.2000 ;
	    RECT 173.7000 279.3000 174.9000 282.9000 ;
	    RECT 177.0000 281.4000 178.2000 282.6000 ;
	    RECT 184.8000 281.7000 186.0000 282.0000 ;
	    RECT 179.4000 280.8000 186.0000 281.7000 ;
	    RECT 179.4000 280.5000 180.6000 280.8000 ;
	    RECT 177.0000 280.2000 178.2000 280.5000 ;
	    RECT 189.0000 279.6000 190.2000 283.8000 ;
	    RECT 197.7000 282.9000 203.4000 284.1000 ;
	    RECT 197.7000 281.1000 198.9000 282.9000 ;
	    RECT 204.3000 282.0000 205.2000 285.0000 ;
	    RECT 179.4000 279.3000 180.6000 279.6000 ;
	    RECT 162.6000 273.3000 163.8000 279.3000 ;
	    RECT 164.7000 278.1000 168.6000 279.3000 ;
	    RECT 173.7000 278.4000 180.6000 279.3000 ;
	    RECT 181.8000 278.4000 183.0000 279.6000 ;
	    RECT 183.9000 278.4000 184.2000 279.6000 ;
	    RECT 188.7000 278.4000 190.2000 279.6000 ;
	    RECT 196.2000 280.2000 198.9000 281.1000 ;
	    RECT 203.4000 281.1000 205.2000 282.0000 ;
	    RECT 196.2000 279.3000 197.4000 280.2000 ;
	    RECT 167.4000 273.3000 168.6000 278.1000 ;
	    RECT 193.8000 278.1000 197.4000 279.3000 ;
	    RECT 169.8000 273.3000 171.0000 277.5000 ;
	    RECT 172.2000 273.3000 173.4000 277.5000 ;
	    RECT 174.6000 273.3000 175.8000 277.5000 ;
	    RECT 177.0000 273.3000 178.2000 276.3000 ;
	    RECT 179.4000 273.3000 180.6000 277.5000 ;
	    RECT 181.8000 273.3000 183.0000 276.3000 ;
	    RECT 184.2000 273.3000 185.4000 277.5000 ;
	    RECT 186.6000 273.3000 187.8000 277.5000 ;
	    RECT 189.0000 273.3000 190.2000 277.5000 ;
	    RECT 191.4000 273.3000 192.6000 277.5000 ;
	    RECT 193.8000 273.3000 195.0000 278.1000 ;
	    RECT 198.6000 273.3000 199.8000 279.3000 ;
	    RECT 203.4000 273.3000 204.6000 281.1000 ;
	    RECT 206.1000 280.2000 207.3000 286.8000 ;
	    RECT 205.8000 279.0000 207.3000 280.2000 ;
	    RECT 340.2000 283.5000 341.4000 291.9000 ;
	    RECT 344.1000 291.6000 350.4000 292.8000 ;
	    RECT 357.0000 292.5000 358.2000 299.7000 ;
	    RECT 359.4000 293.7000 360.6000 299.7000 ;
	    RECT 361.8000 292.5000 363.0000 299.7000 ;
	    RECT 364.2000 293.7000 365.4000 299.7000 ;
	    RECT 344.1000 291.0000 345.0000 291.6000 ;
	    RECT 342.6000 289.8000 345.0000 291.0000 ;
	    RECT 349.5000 290.7000 358.2000 291.6000 ;
	    RECT 346.5000 289.8000 348.6000 290.7000 ;
	    RECT 346.5000 289.5000 355.8000 289.8000 ;
	    RECT 347.7000 288.9000 355.8000 289.5000 ;
	    RECT 354.6000 288.6000 355.8000 288.9000 ;
	    RECT 357.3000 289.5000 358.2000 290.7000 ;
	    RECT 359.1000 290.4000 363.0000 291.6000 ;
	    RECT 366.6000 290.4000 367.8000 299.7000 ;
	    RECT 369.0000 295.5000 370.2000 299.7000 ;
	    RECT 371.4000 295.5000 372.6000 299.7000 ;
	    RECT 373.8000 295.5000 375.0000 299.7000 ;
	    RECT 376.2000 293.7000 377.4000 299.7000 ;
	    RECT 371.4000 291.6000 377.7000 292.8000 ;
	    RECT 378.6000 291.6000 379.8000 299.7000 ;
	    RECT 381.0000 293.7000 382.2000 299.7000 ;
	    RECT 383.4000 292.8000 384.6000 299.7000 ;
	    RECT 385.8000 293.7000 387.0000 299.7000 ;
	    RECT 383.4000 291.9000 387.3000 292.8000 ;
	    RECT 388.2000 292.5000 389.4000 299.7000 ;
	    RECT 390.6000 293.7000 391.8000 299.7000 ;
	    RECT 405.0000 299.4000 406.2000 300.6000 ;
	    RECT 378.6000 290.4000 382.5000 291.6000 ;
	    RECT 369.0000 289.5000 370.2000 289.8000 ;
	    RECT 357.3000 288.6000 370.2000 289.5000 ;
	    RECT 373.8000 289.5000 375.0000 289.8000 ;
	    RECT 386.4000 289.5000 387.3000 291.9000 ;
	    RECT 388.2000 291.4500 389.4000 291.6000 ;
	    RECT 393.0000 291.4500 394.2000 291.6000 ;
	    RECT 388.2000 290.5500 394.2000 291.4500 ;
	    RECT 388.2000 290.4000 389.4000 290.5500 ;
	    RECT 393.0000 290.4000 394.2000 290.5500 ;
	    RECT 373.8000 288.6000 387.3000 289.5000 ;
	    RECT 345.0000 287.4000 346.2000 288.6000 ;
	    RECT 350.1000 287.7000 351.3000 288.0000 ;
	    RECT 347.1000 286.8000 385.5000 287.7000 ;
	    RECT 384.3000 286.5000 385.5000 286.8000 ;
	    RECT 386.4000 285.9000 387.3000 288.6000 ;
	    RECT 388.2000 288.0000 389.4000 289.5000 ;
	    RECT 388.2000 286.8000 389.7000 288.0000 ;
	    RECT 453.0000 287.7000 454.2000 299.7000 ;
	    RECT 455.4000 286.8000 456.6000 299.7000 ;
	    RECT 457.8000 287.7000 459.0000 299.7000 ;
	    RECT 460.2000 286.8000 461.4000 299.7000 ;
	    RECT 462.6000 287.7000 463.8000 299.7000 ;
	    RECT 465.0000 286.8000 466.2000 299.7000 ;
	    RECT 467.4000 287.7000 468.6000 299.7000 ;
	    RECT 469.8000 286.8000 471.0000 299.7000 ;
	    RECT 472.2000 287.7000 473.4000 299.7000 ;
	    RECT 484.2000 293.7000 485.4000 299.7000 ;
	    RECT 342.3000 285.0000 348.9000 285.9000 ;
	    RECT 342.3000 284.7000 343.5000 285.0000 ;
	    RECT 349.8000 284.4000 351.0000 285.6000 ;
	    RECT 351.9000 285.0000 377.4000 285.9000 ;
	    RECT 386.4000 285.0000 387.6000 285.9000 ;
	    RECT 376.2000 284.1000 377.4000 285.0000 ;
	    RECT 340.2000 282.3000 353.4000 283.5000 ;
	    RECT 354.3000 282.9000 357.3000 284.1000 ;
	    RECT 363.0000 282.9000 367.8000 284.1000 ;
	    RECT 205.8000 273.3000 207.0000 279.0000 ;
	    RECT 208.2000 273.3000 209.4000 276.3000 ;
	    RECT 340.2000 273.3000 341.4000 282.3000 ;
	    RECT 343.8000 280.2000 348.3000 281.4000 ;
	    RECT 347.1000 279.3000 348.3000 280.2000 ;
	    RECT 356.1000 279.3000 357.3000 282.9000 ;
	    RECT 359.4000 281.4000 360.6000 282.6000 ;
	    RECT 367.2000 281.7000 368.4000 282.0000 ;
	    RECT 361.8000 280.8000 368.4000 281.7000 ;
	    RECT 361.8000 280.5000 363.0000 280.8000 ;
	    RECT 359.4000 280.2000 360.6000 280.5000 ;
	    RECT 371.4000 279.6000 372.6000 283.8000 ;
	    RECT 380.1000 282.9000 385.8000 284.1000 ;
	    RECT 380.1000 281.1000 381.3000 282.9000 ;
	    RECT 386.7000 282.0000 387.6000 285.0000 ;
	    RECT 361.8000 279.3000 363.0000 279.6000 ;
	    RECT 345.0000 273.3000 346.2000 279.3000 ;
	    RECT 347.1000 278.1000 351.0000 279.3000 ;
	    RECT 356.1000 278.4000 363.0000 279.3000 ;
	    RECT 364.2000 278.4000 365.4000 279.6000 ;
	    RECT 366.3000 278.4000 366.6000 279.6000 ;
	    RECT 371.1000 278.4000 372.6000 279.6000 ;
	    RECT 378.6000 280.2000 381.3000 281.1000 ;
	    RECT 385.8000 281.1000 387.6000 282.0000 ;
	    RECT 378.6000 279.3000 379.8000 280.2000 ;
	    RECT 349.8000 273.3000 351.0000 278.1000 ;
	    RECT 376.2000 278.1000 379.8000 279.3000 ;
	    RECT 352.2000 273.3000 353.4000 277.5000 ;
	    RECT 354.6000 273.3000 355.8000 277.5000 ;
	    RECT 357.0000 273.3000 358.2000 277.5000 ;
	    RECT 359.4000 273.3000 360.6000 276.3000 ;
	    RECT 361.8000 273.3000 363.0000 277.5000 ;
	    RECT 364.2000 273.3000 365.4000 276.3000 ;
	    RECT 366.6000 273.3000 367.8000 277.5000 ;
	    RECT 369.0000 273.3000 370.2000 277.5000 ;
	    RECT 371.4000 273.3000 372.6000 277.5000 ;
	    RECT 373.8000 273.3000 375.0000 277.5000 ;
	    RECT 376.2000 273.3000 377.4000 278.1000 ;
	    RECT 381.0000 273.3000 382.2000 279.3000 ;
	    RECT 385.8000 273.3000 387.0000 281.1000 ;
	    RECT 388.5000 280.2000 389.7000 286.8000 ;
	    RECT 453.0000 286.5000 456.6000 286.8000 ;
	    RECT 455.1000 285.6000 456.6000 286.5000 ;
	    RECT 458.1000 285.6000 461.4000 286.8000 ;
	    RECT 462.9000 285.6000 466.2000 286.8000 ;
	    RECT 468.3000 285.6000 471.0000 286.8000 ;
	    RECT 453.0000 284.4000 454.2000 285.6000 ;
	    RECT 458.1000 283.5000 459.3000 285.6000 ;
	    RECT 462.9000 283.5000 464.1000 285.6000 ;
	    RECT 468.3000 283.5000 469.5000 285.6000 ;
	    RECT 486.6000 283.5000 487.8000 299.7000 ;
	    RECT 501.0000 299.4000 502.2000 300.6000 ;
	    RECT 513.0000 287.7000 514.2000 299.7000 ;
	    RECT 516.9000 288.6000 518.1000 299.7000 ;
	    RECT 519.3000 293.7000 520.5000 299.7000 ;
	    RECT 539.4000 293.7000 540.6000 299.7000 ;
	    RECT 519.0000 290.4000 520.2000 291.6000 ;
	    RECT 519.3000 289.5000 520.2000 290.4000 ;
	    RECT 516.9000 287.7000 518.4000 288.6000 ;
	    RECT 515.4000 285.4500 516.6000 285.6000 ;
	    RECT 498.7500 284.5500 516.6000 285.4500 ;
	    RECT 453.0000 281.4000 454.2000 283.5000 ;
	    RECT 455.4000 282.3000 459.3000 283.5000 ;
	    RECT 460.5000 282.3000 464.1000 283.5000 ;
	    RECT 465.6000 282.3000 469.5000 283.5000 ;
	    RECT 470.7000 282.3000 471.3000 283.5000 ;
	    RECT 486.6000 282.4500 487.8000 282.6000 ;
	    RECT 498.7500 282.4500 499.6500 284.5500 ;
	    RECT 515.4000 284.4000 516.6000 284.5500 ;
	    RECT 515.4000 283.2000 516.6000 283.5000 ;
	    RECT 517.5000 282.6000 518.4000 287.7000 ;
	    RECT 520.2000 287.4000 521.4000 288.6000 ;
	    RECT 520.3500 285.4500 521.2500 287.4000 ;
	    RECT 541.8000 286.5000 543.0000 299.7000 ;
	    RECT 544.2000 293.7000 545.4000 299.7000 ;
	    RECT 544.2000 289.5000 545.4000 289.8000 ;
	    RECT 568.2000 288.6000 569.4000 299.7000 ;
	    RECT 570.6000 289.5000 571.8000 299.7000 ;
	    RECT 573.0000 288.6000 574.2000 299.7000 ;
	    RECT 544.2000 287.4000 545.4000 288.6000 ;
	    RECT 568.2000 287.7000 574.2000 288.6000 ;
	    RECT 575.4000 287.7000 576.6000 299.7000 ;
	    RECT 707.4000 293.7000 708.6000 299.7000 ;
	    RECT 709.8000 292.5000 711.0000 299.7000 ;
	    RECT 712.2000 293.7000 713.4000 299.7000 ;
	    RECT 714.6000 292.8000 715.8000 299.7000 ;
	    RECT 717.0000 293.7000 718.2000 299.7000 ;
	    RECT 711.9000 291.9000 715.8000 292.8000 ;
	    RECT 709.8000 290.4000 711.0000 291.6000 ;
	    RECT 711.9000 289.5000 712.8000 291.9000 ;
	    RECT 719.4000 291.6000 720.6000 299.7000 ;
	    RECT 721.8000 293.7000 723.0000 299.7000 ;
	    RECT 724.2000 295.5000 725.4000 299.7000 ;
	    RECT 726.6000 295.5000 727.8000 299.7000 ;
	    RECT 729.0000 295.5000 730.2000 299.7000 ;
	    RECT 721.5000 291.6000 727.8000 292.8000 ;
	    RECT 716.7000 290.4000 720.6000 291.6000 ;
	    RECT 731.4000 290.4000 732.6000 299.7000 ;
	    RECT 733.8000 293.7000 735.0000 299.7000 ;
	    RECT 736.2000 292.5000 737.4000 299.7000 ;
	    RECT 738.6000 293.7000 739.8000 299.7000 ;
	    RECT 741.0000 292.5000 742.2000 299.7000 ;
	    RECT 743.4000 295.5000 744.6000 299.7000 ;
	    RECT 745.8000 295.5000 747.0000 299.7000 ;
	    RECT 748.2000 293.7000 749.4000 299.7000 ;
	    RECT 750.6000 292.8000 751.8000 299.7000 ;
	    RECT 753.0000 293.7000 754.2000 300.6000 ;
	    RECT 755.4000 294.6000 756.6000 299.7000 ;
	    RECT 755.4000 293.7000 756.9000 294.6000 ;
	    RECT 757.8000 293.7000 759.0000 299.7000 ;
	    RECT 756.0000 292.8000 756.9000 293.7000 ;
	    RECT 748.8000 291.6000 755.1000 292.8000 ;
	    RECT 756.0000 291.9000 759.0000 292.8000 ;
	    RECT 736.2000 290.4000 740.1000 291.6000 ;
	    RECT 741.0000 290.7000 749.7000 291.6000 ;
	    RECT 754.2000 291.0000 755.1000 291.6000 ;
	    RECT 724.2000 289.5000 725.4000 289.8000 ;
	    RECT 709.8000 288.0000 711.0000 289.5000 ;
	    RECT 575.4000 286.5000 576.3000 287.7000 ;
	    RECT 709.5000 286.8000 711.0000 288.0000 ;
	    RECT 711.9000 288.6000 725.4000 289.5000 ;
	    RECT 729.0000 289.5000 730.2000 289.8000 ;
	    RECT 741.0000 289.5000 741.9000 290.7000 ;
	    RECT 750.6000 289.8000 752.7000 290.7000 ;
	    RECT 754.2000 289.8000 756.6000 291.0000 ;
	    RECT 729.0000 288.6000 741.9000 289.5000 ;
	    RECT 743.4000 289.5000 752.7000 289.8000 ;
	    RECT 743.4000 288.9000 751.5000 289.5000 ;
	    RECT 743.4000 288.6000 744.6000 288.9000 ;
	    RECT 541.8000 285.4500 543.0000 285.6000 ;
	    RECT 520.3500 284.5500 543.0000 285.4500 ;
	    RECT 541.8000 284.4000 543.0000 284.5500 ;
	    RECT 568.2000 284.4000 569.4000 285.6000 ;
	    RECT 570.3000 284.7000 570.6000 286.2000 ;
	    RECT 573.0000 284.7000 574.5000 285.6000 ;
	    RECT 575.4000 285.4500 576.6000 285.6000 ;
	    RECT 707.4000 285.4500 708.6000 285.6000 ;
	    RECT 570.6000 283.5000 571.8000 283.8000 ;
	    RECT 458.1000 281.4000 459.3000 282.3000 ;
	    RECT 462.9000 281.4000 464.1000 282.3000 ;
	    RECT 468.3000 281.4000 469.5000 282.3000 ;
	    RECT 486.6000 281.5500 499.6500 282.4500 ;
	    RECT 501.0000 282.4500 502.2000 282.6000 ;
	    RECT 513.0000 282.4500 514.2000 282.6000 ;
	    RECT 501.0000 281.5500 514.2000 282.4500 ;
	    RECT 486.6000 281.4000 487.8000 281.5500 ;
	    RECT 501.0000 281.4000 502.2000 281.5500 ;
	    RECT 513.0000 281.4000 514.2000 281.5500 ;
	    RECT 453.0000 280.2000 456.6000 281.4000 ;
	    RECT 458.1000 280.2000 461.4000 281.4000 ;
	    RECT 462.9000 280.2000 466.2000 281.4000 ;
	    RECT 468.3000 280.2000 471.0000 281.4000 ;
	    RECT 515.1000 280.8000 515.4000 282.3000 ;
	    RECT 517.5000 281.4000 519.3000 282.6000 ;
	    RECT 520.2000 282.4500 521.4000 282.6000 ;
	    RECT 527.4000 282.4500 528.6000 282.6000 ;
	    RECT 520.2000 281.5500 528.6000 282.4500 ;
	    RECT 520.2000 281.4000 521.4000 281.5500 ;
	    RECT 527.4000 281.4000 528.6000 281.5500 ;
	    RECT 539.4000 281.4000 540.6000 282.6000 ;
	    RECT 388.2000 279.0000 389.7000 280.2000 ;
	    RECT 388.2000 273.3000 389.4000 279.0000 ;
	    RECT 390.6000 273.3000 391.8000 276.3000 ;
	    RECT 453.0000 273.3000 454.2000 279.3000 ;
	    RECT 455.4000 273.3000 456.6000 280.2000 ;
	    RECT 457.8000 273.3000 459.0000 279.3000 ;
	    RECT 460.2000 273.3000 461.4000 280.2000 ;
	    RECT 462.6000 273.3000 463.8000 279.3000 ;
	    RECT 465.0000 273.3000 466.2000 280.2000 ;
	    RECT 467.4000 273.3000 468.6000 279.3000 ;
	    RECT 469.8000 273.3000 471.0000 280.2000 ;
	    RECT 472.2000 273.3000 473.4000 279.3000 ;
	    RECT 484.2000 278.4000 485.4000 279.6000 ;
	    RECT 484.2000 277.2000 485.4000 277.5000 ;
	    RECT 484.2000 273.3000 485.4000 276.3000 ;
	    RECT 486.6000 273.3000 487.8000 280.5000 ;
	    RECT 513.3000 279.3000 518.7000 279.9000 ;
	    RECT 520.2000 279.3000 521.1000 280.5000 ;
	    RECT 539.4000 280.2000 540.6000 280.5000 ;
	    RECT 541.8000 279.3000 543.0000 283.5000 ;
	    RECT 570.6000 281.4000 571.8000 282.6000 ;
	    RECT 573.0000 279.3000 573.9000 284.7000 ;
	    RECT 575.4000 284.5500 708.6000 285.4500 ;
	    RECT 575.4000 284.4000 576.6000 284.5500 ;
	    RECT 707.4000 284.4000 708.6000 284.5500 ;
	    RECT 709.5000 280.2000 710.7000 286.8000 ;
	    RECT 711.9000 285.9000 712.8000 288.6000 ;
	    RECT 747.9000 287.7000 749.1000 288.0000 ;
	    RECT 713.7000 286.8000 752.1000 287.7000 ;
	    RECT 753.0000 287.4000 754.2000 288.6000 ;
	    RECT 713.7000 286.5000 714.9000 286.8000 ;
	    RECT 711.6000 285.0000 712.8000 285.9000 ;
	    RECT 721.8000 285.0000 747.3000 285.9000 ;
	    RECT 711.6000 282.0000 712.5000 285.0000 ;
	    RECT 721.8000 284.1000 723.0000 285.0000 ;
	    RECT 748.2000 284.4000 749.4000 285.6000 ;
	    RECT 750.3000 285.0000 756.9000 285.9000 ;
	    RECT 755.7000 284.7000 756.9000 285.0000 ;
	    RECT 713.4000 282.9000 719.1000 284.1000 ;
	    RECT 711.6000 281.1000 713.4000 282.0000 ;
	    RECT 575.4000 279.4500 576.6000 279.6000 ;
	    RECT 589.8000 279.4500 591.0000 279.6000 ;
	    RECT 513.0000 279.0000 519.0000 279.3000 ;
	    RECT 513.0000 273.3000 514.2000 279.0000 ;
	    RECT 515.4000 273.3000 516.6000 278.1000 ;
	    RECT 517.8000 273.3000 519.0000 279.0000 ;
	    RECT 520.2000 273.3000 521.4000 279.3000 ;
	    RECT 539.4000 273.3000 540.6000 279.3000 ;
	    RECT 541.8000 278.4000 544.5000 279.3000 ;
	    RECT 543.3000 273.3000 544.5000 278.4000 ;
	    RECT 569.1000 273.3000 570.3000 279.3000 ;
	    RECT 573.0000 273.3000 574.2000 279.3000 ;
	    RECT 575.4000 278.5500 591.0000 279.4500 ;
	    RECT 709.5000 279.0000 711.0000 280.2000 ;
	    RECT 575.4000 278.4000 576.6000 278.5500 ;
	    RECT 589.8000 278.4000 591.0000 278.5500 ;
	    RECT 575.1000 277.2000 576.3000 277.5000 ;
	    RECT 606.6000 276.4500 607.8000 276.6000 ;
	    RECT 621.0000 276.4500 622.2000 276.6000 ;
	    RECT 575.4000 273.3000 576.6000 276.3000 ;
	    RECT 606.6000 275.5500 622.2000 276.4500 ;
	    RECT 606.6000 275.4000 607.8000 275.5500 ;
	    RECT 621.0000 275.4000 622.2000 275.5500 ;
	    RECT 707.4000 273.3000 708.6000 276.3000 ;
	    RECT 709.8000 273.3000 711.0000 279.0000 ;
	    RECT 712.2000 273.3000 713.4000 281.1000 ;
	    RECT 717.9000 281.1000 719.1000 282.9000 ;
	    RECT 717.9000 280.2000 720.6000 281.1000 ;
	    RECT 719.4000 279.3000 720.6000 280.2000 ;
	    RECT 726.6000 279.6000 727.8000 283.8000 ;
	    RECT 731.4000 282.9000 736.2000 284.1000 ;
	    RECT 741.9000 282.9000 744.9000 284.1000 ;
	    RECT 757.8000 283.5000 759.0000 291.9000 ;
	    RECT 772.2000 283.5000 773.4000 299.7000 ;
	    RECT 774.6000 293.7000 775.8000 299.7000 ;
	    RECT 781.8000 299.4000 783.0000 300.6000 ;
	    RECT 825.0000 287.7000 826.2000 299.7000 ;
	    RECT 827.4000 286.8000 828.6000 299.7000 ;
	    RECT 829.8000 287.7000 831.0000 299.7000 ;
	    RECT 832.2000 286.8000 833.4000 299.7000 ;
	    RECT 834.6000 287.7000 835.8000 299.7000 ;
	    RECT 837.0000 286.8000 838.2000 299.7000 ;
	    RECT 839.4000 287.7000 840.6000 299.7000 ;
	    RECT 841.8000 286.8000 843.0000 299.7000 ;
	    RECT 844.2000 287.7000 845.4000 299.7000 ;
	    RECT 870.6000 287.7000 871.8000 299.7000 ;
	    RECT 874.5000 288.6000 875.7000 299.7000 ;
	    RECT 876.9000 293.7000 878.1000 299.7000 ;
	    RECT 876.6000 290.4000 877.8000 291.6000 ;
	    RECT 876.9000 289.5000 877.8000 290.4000 ;
	    RECT 874.5000 287.7000 876.0000 288.6000 ;
	    RECT 827.4000 285.6000 830.1000 286.8000 ;
	    RECT 832.2000 285.6000 835.5000 286.8000 ;
	    RECT 837.0000 285.6000 840.3000 286.8000 ;
	    RECT 841.8000 286.5000 845.4000 286.8000 ;
	    RECT 841.8000 285.6000 843.3000 286.5000 ;
	    RECT 828.9000 283.5000 830.1000 285.6000 ;
	    RECT 834.3000 283.5000 835.5000 285.6000 ;
	    RECT 839.1000 283.5000 840.3000 285.6000 ;
	    RECT 844.2000 284.4000 845.4000 285.6000 ;
	    RECT 873.0000 284.4000 874.2000 285.6000 ;
	    RECT 730.8000 281.7000 732.0000 282.0000 ;
	    RECT 730.8000 280.8000 737.4000 281.7000 ;
	    RECT 738.6000 281.4000 739.8000 282.6000 ;
	    RECT 736.2000 280.5000 737.4000 280.8000 ;
	    RECT 738.6000 280.2000 739.8000 280.5000 ;
	    RECT 717.0000 273.3000 718.2000 279.3000 ;
	    RECT 719.4000 278.1000 723.0000 279.3000 ;
	    RECT 726.6000 278.4000 728.1000 279.6000 ;
	    RECT 732.6000 278.4000 732.9000 279.6000 ;
	    RECT 733.8000 278.4000 735.0000 279.6000 ;
	    RECT 736.2000 279.3000 737.4000 279.6000 ;
	    RECT 741.9000 279.3000 743.1000 282.9000 ;
	    RECT 745.8000 282.3000 759.0000 283.5000 ;
	    RECT 750.9000 280.2000 755.4000 281.4000 ;
	    RECT 750.9000 279.3000 752.1000 280.2000 ;
	    RECT 736.2000 278.4000 743.1000 279.3000 ;
	    RECT 721.8000 273.3000 723.0000 278.1000 ;
	    RECT 748.2000 278.1000 752.1000 279.3000 ;
	    RECT 724.2000 273.3000 725.4000 277.5000 ;
	    RECT 726.6000 273.3000 727.8000 277.5000 ;
	    RECT 729.0000 273.3000 730.2000 277.5000 ;
	    RECT 731.4000 273.3000 732.6000 277.5000 ;
	    RECT 733.8000 273.3000 735.0000 276.3000 ;
	    RECT 736.2000 273.3000 737.4000 277.5000 ;
	    RECT 738.6000 273.3000 739.8000 276.3000 ;
	    RECT 741.0000 273.3000 742.2000 277.5000 ;
	    RECT 743.4000 273.3000 744.6000 277.5000 ;
	    RECT 745.8000 273.3000 747.0000 277.5000 ;
	    RECT 748.2000 273.3000 749.4000 278.1000 ;
	    RECT 750.6000 272.4000 751.8000 273.6000 ;
	    RECT 753.0000 273.3000 754.2000 279.3000 ;
	    RECT 757.8000 273.3000 759.0000 282.3000 ;
	    RECT 772.2000 282.4500 773.4000 282.6000 ;
	    RECT 779.4000 282.4500 780.6000 282.6000 ;
	    RECT 772.2000 281.5500 780.6000 282.4500 ;
	    RECT 827.1000 282.3000 827.7000 283.5000 ;
	    RECT 828.9000 282.3000 832.8000 283.5000 ;
	    RECT 834.3000 282.3000 837.9000 283.5000 ;
	    RECT 839.1000 282.3000 843.0000 283.5000 ;
	    RECT 772.2000 281.4000 773.4000 281.5500 ;
	    RECT 779.4000 281.4000 780.6000 281.5500 ;
	    RECT 828.9000 281.4000 830.1000 282.3000 ;
	    RECT 834.3000 281.4000 835.5000 282.3000 ;
	    RECT 839.1000 281.4000 840.3000 282.3000 ;
	    RECT 844.2000 281.4000 845.4000 283.5000 ;
	    RECT 873.0000 283.2000 874.2000 283.5000 ;
	    RECT 875.1000 282.6000 876.0000 287.7000 ;
	    RECT 877.8000 287.4000 879.0000 288.6000 ;
	    RECT 889.8000 283.5000 891.0000 299.7000 ;
	    RECT 892.2000 293.7000 893.4000 299.7000 ;
	    RECT 969.0000 286.8000 970.2000 299.7000 ;
	    RECT 971.4000 287.7000 972.6000 299.7000 ;
	    RECT 975.3000 293.7000 977.1000 299.7000 ;
	    RECT 979.8000 293.7000 981.0000 299.7000 ;
	    RECT 982.2000 293.7000 983.4000 299.7000 ;
	    RECT 984.6000 293.7000 985.8000 299.7000 ;
	    RECT 988.8000 294.6000 990.0000 299.7000 ;
	    RECT 988.8000 293.7000 991.8000 294.6000 ;
	    RECT 976.2000 292.5000 977.4000 293.7000 ;
	    RECT 982.5000 292.8000 983.4000 293.7000 ;
	    RECT 981.3000 291.9000 986.7000 292.8000 ;
	    RECT 990.6000 292.5000 991.8000 293.7000 ;
	    RECT 981.3000 291.6000 982.5000 291.9000 ;
	    RECT 985.5000 291.6000 986.7000 291.9000 ;
	    RECT 975.0000 289.8000 977.1000 291.0000 ;
	    RECT 976.2000 288.3000 977.1000 289.8000 ;
	    RECT 979.5000 289.5000 982.8000 290.4000 ;
	    RECT 979.5000 289.2000 980.7000 289.5000 ;
	    RECT 976.2000 287.4000 979.8000 288.3000 ;
	    RECT 969.0000 286.5000 975.3000 286.8000 ;
	    RECT 971.1000 285.9000 975.3000 286.5000 ;
	    RECT 974.1000 285.6000 975.3000 285.9000 ;
	    RECT 969.0000 284.4000 970.2000 285.6000 ;
	    RECT 971.7000 284.7000 972.9000 285.0000 ;
	    RECT 971.7000 283.8000 977.4000 284.7000 ;
	    RECT 976.2000 283.5000 977.4000 283.8000 ;
	    RECT 858.6000 282.4500 859.8000 282.6000 ;
	    RECT 870.6000 282.4500 871.8000 282.6000 ;
	    RECT 858.6000 281.5500 871.8000 282.4500 ;
	    RECT 858.6000 281.4000 859.8000 281.5500 ;
	    RECT 870.6000 281.4000 871.8000 281.5500 ;
	    RECT 772.2000 273.3000 773.4000 280.5000 ;
	    RECT 827.4000 280.2000 830.1000 281.4000 ;
	    RECT 832.2000 280.2000 835.5000 281.4000 ;
	    RECT 837.0000 280.2000 840.3000 281.4000 ;
	    RECT 841.8000 280.2000 845.4000 281.4000 ;
	    RECT 872.7000 280.8000 873.0000 282.3000 ;
	    RECT 875.1000 281.4000 876.9000 282.6000 ;
	    RECT 877.8000 281.4000 879.0000 282.6000 ;
	    RECT 880.2000 282.4500 881.4000 282.6000 ;
	    RECT 889.8000 282.4500 891.0000 282.6000 ;
	    RECT 880.2000 281.5500 891.0000 282.4500 ;
	    RECT 880.2000 281.4000 881.4000 281.5500 ;
	    RECT 889.8000 281.4000 891.0000 281.5500 ;
	    RECT 969.0000 280.8000 970.2000 283.5000 ;
	    RECT 978.9000 282.6000 979.8000 287.4000 ;
	    RECT 981.9000 287.7000 982.8000 289.5000 ;
	    RECT 983.7000 289.5000 984.9000 289.8000 ;
	    RECT 990.6000 289.5000 991.8000 289.8000 ;
	    RECT 983.7000 288.6000 991.8000 289.5000 ;
	    RECT 993.0000 288.0000 994.2000 299.7000 ;
	    RECT 981.9000 287.1000 989.1000 287.7000 ;
	    RECT 995.4000 287.1000 996.6000 299.7000 ;
	    RECT 1014.6000 293.7000 1015.8000 299.7000 ;
	    RECT 981.9000 286.8000 996.6000 287.1000 ;
	    RECT 987.9000 286.5000 996.6000 286.8000 ;
	    RECT 1017.0000 286.5000 1018.2000 299.7000 ;
	    RECT 1019.4000 293.7000 1020.6000 299.7000 ;
	    RECT 1043.4000 293.7000 1044.6000 299.7000 ;
	    RECT 1045.8000 293.7000 1047.0000 299.7000 ;
	    RECT 1048.2001 294.3000 1049.4000 299.7000 ;
	    RECT 1046.1000 293.4000 1047.0000 293.7000 ;
	    RECT 1050.6000 293.7000 1051.8000 299.7000 ;
	    RECT 1050.6000 293.4000 1051.5000 293.7000 ;
	    RECT 1046.1000 292.5000 1051.5000 293.4000 ;
	    RECT 1045.8000 291.4500 1047.0000 291.6000 ;
	    RECT 1021.9500 290.5500 1047.0000 291.4500 ;
	    RECT 1019.4000 289.5000 1020.6000 289.8000 ;
	    RECT 1019.4000 288.4500 1020.6000 288.6000 ;
	    RECT 1021.9500 288.4500 1022.8500 290.5500 ;
	    RECT 1045.8000 290.4000 1047.0000 290.5500 ;
	    RECT 1048.2001 290.4000 1049.4000 291.6000 ;
	    RECT 1050.6000 289.5000 1051.5000 292.5000 ;
	    RECT 1048.2001 289.2000 1049.4000 289.5000 ;
	    RECT 1019.4000 287.5500 1022.8500 288.4500 ;
	    RECT 1019.4000 287.4000 1020.6000 287.5500 ;
	    RECT 1043.4000 287.4000 1044.6000 288.6000 ;
	    RECT 1050.6000 288.4500 1051.8000 288.6000 ;
	    RECT 1067.4000 288.4500 1068.6000 288.6000 ;
	    RECT 1050.6000 287.5500 1068.6000 288.4500 ;
	    RECT 1069.8000 287.7000 1071.0000 299.7000 ;
	    RECT 1073.7001 288.9000 1074.9000 299.7000 ;
	    RECT 1098.6000 293.7000 1099.8000 299.7000 ;
	    RECT 1101.0000 294.3000 1102.2001 299.7000 ;
	    RECT 1098.9000 293.4000 1099.8000 293.7000 ;
	    RECT 1103.4000 293.7000 1104.6000 299.7000 ;
	    RECT 1105.8000 293.7000 1107.0000 299.7000 ;
	    RECT 1103.4000 293.4000 1104.3000 293.7000 ;
	    RECT 1098.9000 292.5000 1104.3000 293.4000 ;
	    RECT 1098.9000 289.5000 1099.8000 292.5000 ;
	    RECT 1101.0000 290.4000 1102.2001 291.6000 ;
	    RECT 1101.0000 289.2000 1102.2001 289.5000 ;
	    RECT 1072.2001 287.7000 1074.9000 288.9000 ;
	    RECT 1050.6000 287.4000 1051.8000 287.5500 ;
	    RECT 1067.4000 287.4000 1068.6000 287.5500 ;
	    RECT 988.2000 286.2000 996.6000 286.5000 ;
	    RECT 1043.4000 286.2000 1044.6000 286.5000 ;
	    RECT 985.8000 284.4000 987.0000 285.6000 ;
	    RECT 1017.0000 285.4500 1018.2000 285.6000 ;
	    RECT 1041.0000 285.4500 1042.2001 285.6000 ;
	    RECT 987.9000 284.4000 993.3000 285.3000 ;
	    RECT 1017.0000 284.5500 1042.2001 285.4500 ;
	    RECT 1017.0000 284.4000 1018.2000 284.5500 ;
	    RECT 1041.0000 284.4000 1042.2001 284.5500 ;
	    RECT 1045.8000 284.4000 1047.0000 285.6000 ;
	    RECT 1047.9000 284.4000 1048.2001 285.6000 ;
	    RECT 992.1000 284.1000 993.3000 284.4000 ;
	    RECT 989.7000 282.6000 990.9000 282.9000 ;
	    RECT 978.9000 281.7000 992.1000 282.6000 ;
	    RECT 979.5000 281.4000 980.7000 281.7000 ;
	    RECT 774.6000 279.4500 775.8000 279.6000 ;
	    RECT 786.6000 279.4500 787.8000 279.6000 ;
	    RECT 796.2000 279.4500 797.4000 279.6000 ;
	    RECT 774.6000 278.5500 797.4000 279.4500 ;
	    RECT 774.6000 278.4000 775.8000 278.5500 ;
	    RECT 786.6000 278.4000 787.8000 278.5500 ;
	    RECT 796.2000 278.4000 797.4000 278.5500 ;
	    RECT 774.6000 277.2000 775.8000 277.5000 ;
	    RECT 774.6000 273.3000 775.8000 276.3000 ;
	    RECT 825.0000 273.3000 826.2000 279.3000 ;
	    RECT 827.4000 273.3000 828.6000 280.2000 ;
	    RECT 829.8000 273.3000 831.0000 279.3000 ;
	    RECT 832.2000 273.3000 833.4000 280.2000 ;
	    RECT 834.6000 273.3000 835.8000 279.3000 ;
	    RECT 837.0000 273.3000 838.2000 280.2000 ;
	    RECT 839.4000 273.3000 840.6000 279.3000 ;
	    RECT 841.8000 273.3000 843.0000 280.2000 ;
	    RECT 870.9000 279.3000 876.3000 279.9000 ;
	    RECT 877.8000 279.3000 878.7000 280.5000 ;
	    RECT 844.2000 273.3000 845.4000 279.3000 ;
	    RECT 870.6000 279.0000 876.6000 279.3000 ;
	    RECT 870.6000 273.3000 871.8000 279.0000 ;
	    RECT 873.0000 273.3000 874.2000 278.1000 ;
	    RECT 875.4000 273.3000 876.6000 279.0000 ;
	    RECT 877.8000 273.3000 879.0000 279.3000 ;
	    RECT 889.8000 273.3000 891.0000 280.5000 ;
	    RECT 969.0000 279.9000 974.7000 280.8000 ;
	    RECT 892.2000 279.4500 893.4000 279.6000 ;
	    RECT 916.2000 279.4500 917.4000 279.6000 ;
	    RECT 892.2000 278.5500 917.4000 279.4500 ;
	    RECT 892.2000 278.4000 893.4000 278.5500 ;
	    RECT 916.2000 278.4000 917.4000 278.5500 ;
	    RECT 892.2000 277.2000 893.4000 277.5000 ;
	    RECT 892.2000 273.3000 893.4000 276.3000 ;
	    RECT 969.0000 273.3000 970.2000 279.9000 ;
	    RECT 973.5000 279.6000 974.7000 279.9000 ;
	    RECT 971.4000 273.3000 972.6000 279.0000 ;
	    RECT 988.2000 278.4000 989.1000 281.7000 ;
	    RECT 993.0000 281.4000 994.2000 282.6000 ;
	    RECT 995.1000 281.4000 995.4000 282.6000 ;
	    RECT 1014.6000 281.4000 1015.8000 282.6000 ;
	    RECT 985.5000 278.1000 986.7000 278.4000 ;
	    RECT 976.2000 276.3000 977.4000 277.5000 ;
	    RECT 982.5000 277.2000 986.7000 278.1000 ;
	    RECT 988.2000 277.2000 989.4000 278.4000 ;
	    RECT 982.5000 276.3000 983.4000 277.2000 ;
	    RECT 990.6000 276.3000 991.8000 277.5000 ;
	    RECT 975.3000 275.4000 977.4000 276.3000 ;
	    RECT 975.3000 273.3000 977.1000 275.4000 ;
	    RECT 979.8000 273.3000 981.0000 276.3000 ;
	    RECT 982.2000 273.3000 983.4000 276.3000 ;
	    RECT 984.6000 273.3000 986.1000 276.3000 ;
	    RECT 988.8000 275.4000 991.8000 276.3000 ;
	    RECT 988.8000 273.3000 990.0000 275.4000 ;
	    RECT 993.0000 273.3000 994.2000 279.3000 ;
	    RECT 995.4000 273.3000 996.6000 280.5000 ;
	    RECT 1014.6000 280.2000 1015.8000 280.5000 ;
	    RECT 1017.0000 279.3000 1018.2000 283.5000 ;
	    RECT 1050.6000 282.6000 1051.5000 286.5000 ;
	    RECT 1072.5000 283.5000 1073.4000 287.7000 ;
	    RECT 1098.6000 287.4000 1099.8000 288.6000 ;
	    RECT 1105.8000 287.4000 1107.0000 288.6000 ;
	    RECT 1074.6000 286.5000 1075.8000 286.8000 ;
	    RECT 1074.6000 285.4500 1075.8000 285.6000 ;
	    RECT 1084.2001 285.4500 1085.4000 285.6000 ;
	    RECT 1074.6000 284.5500 1085.4000 285.4500 ;
	    RECT 1074.6000 284.4000 1075.8000 284.5500 ;
	    RECT 1084.2001 284.4000 1085.4000 284.5500 ;
	    RECT 1098.9000 282.6000 1099.8000 286.5000 ;
	    RECT 1105.8000 286.2000 1107.0000 286.5000 ;
	    RECT 1102.2001 284.4000 1102.5000 285.6000 ;
	    RECT 1103.4000 284.4000 1104.6000 285.6000 ;
	    RECT 1117.8000 283.5000 1119.0000 299.7000 ;
	    RECT 1120.2001 293.7000 1121.4000 299.7000 ;
	    RECT 1151.4000 293.7000 1152.6000 299.7000 ;
	    RECT 1153.8000 293.7000 1155.0000 299.7000 ;
	    RECT 1156.2001 294.3000 1157.4000 299.7000 ;
	    RECT 1154.1000 293.4000 1155.0000 293.7000 ;
	    RECT 1158.6000 293.7000 1159.8000 299.7000 ;
	    RECT 1163.4000 297.4500 1164.6000 297.6000 ;
	    RECT 1180.2001 297.4500 1181.4000 297.6000 ;
	    RECT 1163.4000 296.5500 1181.4000 297.4500 ;
	    RECT 1163.4000 296.4000 1164.6000 296.5500 ;
	    RECT 1180.2001 296.4000 1181.4000 296.5500 ;
	    RECT 1185.0000 293.7000 1186.2001 299.7000 ;
	    RECT 1187.4000 293.7000 1188.6000 299.7000 ;
	    RECT 1189.8000 294.3000 1191.0000 299.7000 ;
	    RECT 1158.6000 293.4000 1159.5000 293.7000 ;
	    RECT 1154.1000 292.5000 1159.5000 293.4000 ;
	    RECT 1187.7001 293.4000 1188.6000 293.7000 ;
	    RECT 1192.2001 293.7000 1193.4000 299.7000 ;
	    RECT 1216.2001 293.7000 1217.4000 299.7000 ;
	    RECT 1218.6000 293.7000 1219.8000 299.7000 ;
	    RECT 1221.0000 294.3000 1222.2001 299.7000 ;
	    RECT 1192.2001 293.4000 1193.1000 293.7000 ;
	    RECT 1187.7001 292.5000 1193.1000 293.4000 ;
	    RECT 1218.9000 293.4000 1219.8000 293.7000 ;
	    RECT 1223.4000 293.7000 1224.6000 299.7000 ;
	    RECT 1235.4000 299.4000 1236.6000 300.6000 ;
	    RECT 1252.2001 298.8000 1258.2001 299.7000 ;
	    RECT 1228.2001 294.4500 1229.4000 294.6000 ;
	    RECT 1242.6000 294.4500 1243.8000 294.6000 ;
	    RECT 1223.4000 293.4000 1224.3000 293.7000 ;
	    RECT 1228.2001 293.5500 1243.8000 294.4500 ;
	    RECT 1228.2001 293.4000 1229.4000 293.5500 ;
	    RECT 1242.6000 293.4000 1243.8000 293.5500 ;
	    RECT 1218.9000 292.5000 1224.3000 293.4000 ;
	    RECT 1149.0000 291.4500 1150.2001 291.6000 ;
	    RECT 1156.2001 291.4500 1157.4000 291.6000 ;
	    RECT 1149.0000 290.5500 1157.4000 291.4500 ;
	    RECT 1149.0000 290.4000 1150.2001 290.5500 ;
	    RECT 1156.2001 290.4000 1157.4000 290.5500 ;
	    RECT 1158.6000 289.5000 1159.5000 292.5000 ;
	    RECT 1165.8000 291.4500 1167.0000 291.6000 ;
	    RECT 1189.8000 291.4500 1191.0000 291.6000 ;
	    RECT 1165.8000 290.5500 1191.0000 291.4500 ;
	    RECT 1165.8000 290.4000 1167.0000 290.5500 ;
	    RECT 1189.8000 290.4000 1191.0000 290.5500 ;
	    RECT 1192.2001 289.5000 1193.1000 292.5000 ;
	    RECT 1221.0000 290.4000 1222.2001 291.6000 ;
	    RECT 1223.4000 289.5000 1224.3000 292.5000 ;
	    RECT 1156.2001 289.2000 1157.4000 289.5000 ;
	    RECT 1189.8000 289.2000 1191.0000 289.5000 ;
	    RECT 1221.0000 289.2000 1222.2001 289.5000 ;
	    RECT 1120.2001 288.4500 1121.4000 288.6000 ;
	    RECT 1151.4000 288.4500 1152.6000 288.6000 ;
	    RECT 1120.2001 287.5500 1152.6000 288.4500 ;
	    RECT 1120.2001 287.4000 1121.4000 287.5500 ;
	    RECT 1151.4000 287.4000 1152.6000 287.5500 ;
	    RECT 1158.6000 288.4500 1159.8000 288.6000 ;
	    RECT 1165.8000 288.4500 1167.0000 288.6000 ;
	    RECT 1158.6000 287.5500 1167.0000 288.4500 ;
	    RECT 1158.6000 287.4000 1159.8000 287.5500 ;
	    RECT 1165.8000 287.4000 1167.0000 287.5500 ;
	    RECT 1185.0000 287.4000 1186.2001 288.6000 ;
	    RECT 1192.2001 288.4500 1193.4000 288.6000 ;
	    RECT 1204.2001 288.4500 1205.4000 288.6000 ;
	    RECT 1192.2001 287.5500 1205.4000 288.4500 ;
	    RECT 1192.2001 287.4000 1193.4000 287.5500 ;
	    RECT 1204.2001 287.4000 1205.4000 287.5500 ;
	    RECT 1206.6000 288.4500 1207.8000 288.6000 ;
	    RECT 1211.4000 288.4500 1212.6000 288.6000 ;
	    RECT 1216.2001 288.4500 1217.4000 288.6000 ;
	    RECT 1206.6000 287.5500 1217.4000 288.4500 ;
	    RECT 1206.6000 287.4000 1207.8000 287.5500 ;
	    RECT 1211.4000 287.4000 1212.6000 287.5500 ;
	    RECT 1216.2001 287.4000 1217.4000 287.5500 ;
	    RECT 1223.4000 288.4500 1224.6000 288.6000 ;
	    RECT 1223.4000 287.5500 1250.8500 288.4500 ;
	    RECT 1252.2001 287.7000 1253.4000 298.8000 ;
	    RECT 1254.6000 287.7000 1255.8000 297.9000 ;
	    RECT 1257.0000 288.6000 1258.2001 298.8000 ;
	    RECT 1259.4000 289.5000 1260.6000 299.7000 ;
	    RECT 1261.8000 288.6000 1263.0000 299.7000 ;
	    RECT 1257.0000 287.7000 1263.0000 288.6000 ;
	    RECT 1223.4000 287.4000 1224.6000 287.5500 ;
	    RECT 1151.4000 286.2000 1152.6000 286.5000 ;
	    RECT 1153.8000 284.4000 1155.0000 285.6000 ;
	    RECT 1155.9000 284.4000 1156.2001 285.6000 ;
	    RECT 1158.6000 282.6000 1159.5000 286.5000 ;
	    RECT 1185.0000 286.2000 1186.2001 286.5000 ;
	    RECT 1187.4000 284.4000 1188.6000 285.6000 ;
	    RECT 1189.5000 284.4000 1189.8000 285.6000 ;
	    RECT 1192.2001 282.6000 1193.1000 286.5000 ;
	    RECT 1216.2001 286.2000 1217.4000 286.5000 ;
	    RECT 1218.6000 284.4000 1219.8000 285.6000 ;
	    RECT 1220.7001 284.4000 1221.0000 285.6000 ;
	    RECT 1223.4000 282.6000 1224.3000 286.5000 ;
	    RECT 1249.9501 285.4500 1250.8500 287.5500 ;
	    RECT 1254.9000 286.8000 1255.8000 287.7000 ;
	    RECT 1252.2001 286.5000 1253.4000 286.8000 ;
	    RECT 1254.9000 286.5000 1257.9000 286.8000 ;
	    RECT 1254.9000 285.9000 1256.1000 286.5000 ;
	    RECT 1252.2001 285.4500 1253.4000 285.6000 ;
	    RECT 1249.9501 284.5500 1253.4000 285.4500 ;
	    RECT 1252.2001 284.4000 1253.4000 284.5500 ;
	    RECT 1257.0000 284.4000 1258.2001 285.6000 ;
	    RECT 1260.6000 284.7000 1260.9000 286.2000 ;
	    RECT 1261.8000 284.4000 1263.0000 285.6000 ;
	    RECT 1254.9000 283.5000 1256.1000 284.4000 ;
	    RECT 1259.4000 283.5000 1260.6000 283.8000 ;
	    RECT 1273.8000 283.5000 1275.0000 299.7000 ;
	    RECT 1276.2001 293.7000 1277.4000 299.7000 ;
	    RECT 1295.4000 287.7000 1296.6000 299.7000 ;
	    RECT 1297.8000 289.5000 1299.0000 299.7000 ;
	    RECT 1300.2001 288.6000 1301.4000 299.7000 ;
	    RECT 1324.2001 293.7000 1325.4000 299.7000 ;
	    RECT 1326.6000 294.3000 1327.8000 299.7000 ;
	    RECT 1324.5000 293.4000 1325.4000 293.7000 ;
	    RECT 1329.0000 293.7000 1330.2001 299.7000 ;
	    RECT 1331.4000 293.7000 1332.6000 299.7000 ;
	    RECT 1365.0000 293.7000 1366.2001 299.7000 ;
	    RECT 1367.4000 294.3000 1368.6000 299.7000 ;
	    RECT 1329.0000 293.4000 1329.9000 293.7000 ;
	    RECT 1324.5000 292.5000 1329.9000 293.4000 ;
	    RECT 1365.3000 293.4000 1366.2001 293.7000 ;
	    RECT 1369.8000 293.7000 1371.0000 299.7000 ;
	    RECT 1372.2001 293.7000 1373.4000 299.7000 ;
	    RECT 1369.8000 293.4000 1370.7001 293.7000 ;
	    RECT 1365.3000 292.5000 1370.7001 293.4000 ;
	    RECT 1324.5000 289.5000 1325.4000 292.5000 ;
	    RECT 1326.6000 291.4500 1327.8000 291.6000 ;
	    RECT 1333.8000 291.4500 1335.0000 291.6000 ;
	    RECT 1326.6000 290.5500 1335.0000 291.4500 ;
	    RECT 1326.6000 290.4000 1327.8000 290.5500 ;
	    RECT 1333.8000 290.4000 1335.0000 290.5500 ;
	    RECT 1365.3000 289.5000 1366.2001 292.5000 ;
	    RECT 1367.4000 290.4000 1368.6000 291.6000 ;
	    RECT 1326.6000 289.2000 1327.8000 289.5000 ;
	    RECT 1367.4000 289.2000 1368.6000 289.5000 ;
	    RECT 1298.1000 287.7000 1301.4000 288.6000 ;
	    RECT 1295.4000 284.4000 1296.3000 287.7000 ;
	    RECT 1298.1000 286.8000 1299.0000 287.7000 ;
	    RECT 1324.2001 287.4000 1325.4000 288.6000 ;
	    RECT 1331.4000 287.4000 1332.6000 288.6000 ;
	    RECT 1362.6000 288.4500 1363.8000 288.6000 ;
	    RECT 1365.0000 288.4500 1366.2001 288.6000 ;
	    RECT 1362.6000 287.5500 1366.2001 288.4500 ;
	    RECT 1362.6000 287.4000 1363.8000 287.5500 ;
	    RECT 1365.0000 287.4000 1366.2001 287.5500 ;
	    RECT 1372.2001 287.4000 1373.4000 288.6000 ;
	    RECT 1398.6000 287.7000 1399.8000 299.7000 ;
	    RECT 1401.0000 288.6000 1402.2001 299.7000 ;
	    RECT 1403.4000 289.5000 1404.6000 299.7000 ;
	    RECT 1405.8000 288.6000 1407.0000 299.7000 ;
	    RECT 1420.2001 293.7000 1421.4000 299.7000 ;
	    RECT 1401.0000 287.7000 1407.0000 288.6000 ;
	    RECT 1297.2001 285.6000 1299.0000 286.8000 ;
	    RECT 1398.9000 286.5000 1399.8000 287.7000 ;
	    RECT 1295.4000 283.5000 1296.6000 284.4000 ;
	    RECT 1049.1000 282.3000 1051.5000 282.6000 ;
	    RECT 1014.6000 273.3000 1015.8000 279.3000 ;
	    RECT 1017.0000 278.4000 1019.7000 279.3000 ;
	    RECT 1018.5000 273.3000 1019.7000 278.4000 ;
	    RECT 1043.4000 273.3000 1044.6000 282.3000 ;
	    RECT 1048.8000 281.7000 1051.5000 282.3000 ;
	    RECT 1072.2001 282.4500 1073.4000 282.6000 ;
	    RECT 1093.8000 282.4500 1095.0000 282.6000 ;
	    RECT 1048.8000 273.3000 1050.0000 281.7000 ;
	    RECT 1072.2001 281.5500 1095.0000 282.4500 ;
	    RECT 1098.9000 282.3000 1101.3000 282.6000 ;
	    RECT 1115.4000 282.4500 1116.6000 282.6000 ;
	    RECT 1117.8000 282.4500 1119.0000 282.6000 ;
	    RECT 1098.9000 281.7000 1101.6000 282.3000 ;
	    RECT 1072.2001 281.4000 1073.4000 281.5500 ;
	    RECT 1093.8000 281.4000 1095.0000 281.5500 ;
	    RECT 1069.8000 278.4000 1071.0000 279.6000 ;
	    RECT 1069.8000 277.2000 1071.0000 277.5000 ;
	    RECT 1072.5000 276.3000 1073.4000 280.5000 ;
	    RECT 1069.8000 273.3000 1071.0000 276.3000 ;
	    RECT 1072.2001 273.3000 1073.4000 276.3000 ;
	    RECT 1074.6000 273.3000 1075.8000 276.3000 ;
	    RECT 1100.4000 273.3000 1101.6000 281.7000 ;
	    RECT 1105.8000 273.3000 1107.0000 282.3000 ;
	    RECT 1115.4000 281.5500 1119.0000 282.4500 ;
	    RECT 1157.1000 282.3000 1159.5000 282.6000 ;
	    RECT 1190.7001 282.3000 1193.1000 282.6000 ;
	    RECT 1221.9000 282.3000 1224.3000 282.6000 ;
	    RECT 1115.4000 281.4000 1116.6000 281.5500 ;
	    RECT 1117.8000 281.4000 1119.0000 281.5500 ;
	    RECT 1117.8000 273.3000 1119.0000 280.5000 ;
	    RECT 1120.2001 278.4000 1121.4000 279.6000 ;
	    RECT 1120.2001 277.2000 1121.4000 277.5000 ;
	    RECT 1120.2001 273.3000 1121.4000 276.3000 ;
	    RECT 1151.4000 273.3000 1152.6000 282.3000 ;
	    RECT 1156.8000 281.7000 1159.5000 282.3000 ;
	    RECT 1156.8000 273.3000 1158.0000 281.7000 ;
	    RECT 1185.0000 273.3000 1186.2001 282.3000 ;
	    RECT 1190.4000 281.7000 1193.1000 282.3000 ;
	    RECT 1190.4000 273.3000 1191.6000 281.7000 ;
	    RECT 1194.6000 276.4500 1195.8000 276.6000 ;
	    RECT 1213.8000 276.4500 1215.0000 276.6000 ;
	    RECT 1194.6000 275.5500 1215.0000 276.4500 ;
	    RECT 1194.6000 275.4000 1195.8000 275.5500 ;
	    RECT 1213.8000 275.4000 1215.0000 275.5500 ;
	    RECT 1216.2001 273.3000 1217.4000 282.3000 ;
	    RECT 1221.6000 281.7000 1224.3000 282.3000 ;
	    RECT 1221.6000 273.3000 1222.8000 281.7000 ;
	    RECT 1254.6000 281.4000 1255.8000 282.6000 ;
	    RECT 1257.0000 279.3000 1257.9000 283.5000 ;
	    RECT 1259.4000 281.4000 1260.6000 282.6000 ;
	    RECT 1273.8000 282.4500 1275.0000 282.6000 ;
	    RECT 1290.6000 282.4500 1291.8000 282.6000 ;
	    RECT 1295.4000 282.4500 1296.6000 282.6000 ;
	    RECT 1273.8000 281.5500 1291.8000 282.4500 ;
	    RECT 1273.8000 281.4000 1275.0000 281.5500 ;
	    RECT 1290.6000 281.4000 1291.8000 281.5500 ;
	    RECT 1293.1500 281.5500 1296.6000 282.4500 ;
	    RECT 1252.2001 273.3000 1253.4000 279.3000 ;
	    RECT 1256.1000 273.3000 1258.5000 279.3000 ;
	    RECT 1261.2001 273.3000 1262.4000 279.3000 ;
	    RECT 1273.8000 273.3000 1275.0000 280.5000 ;
	    RECT 1276.2001 278.4000 1277.4000 279.6000 ;
	    RECT 1285.8000 279.4500 1287.0000 279.6000 ;
	    RECT 1293.1500 279.4500 1294.0500 281.5500 ;
	    RECT 1295.4000 281.4000 1296.6000 281.5500 ;
	    RECT 1298.1000 281.1000 1299.0000 285.6000 ;
	    RECT 1300.2001 284.4000 1301.4000 285.6000 ;
	    RECT 1300.2001 283.2000 1301.4000 283.5000 ;
	    RECT 1324.5000 282.6000 1325.4000 286.5000 ;
	    RECT 1331.4000 286.2000 1332.6000 286.5000 ;
	    RECT 1327.8000 284.4000 1328.1000 285.6000 ;
	    RECT 1329.0000 284.4000 1330.2001 285.6000 ;
	    RECT 1365.3000 282.6000 1366.2001 286.5000 ;
	    RECT 1372.2001 286.2000 1373.4000 286.5000 ;
	    RECT 1368.6000 284.4000 1368.9000 285.6000 ;
	    RECT 1369.8000 284.4000 1371.0000 285.6000 ;
	    RECT 1393.8000 285.4500 1395.0000 285.6000 ;
	    RECT 1398.6000 285.4500 1399.8000 285.6000 ;
	    RECT 1393.8000 284.5500 1399.8000 285.4500 ;
	    RECT 1400.7001 284.7000 1402.2001 285.6000 ;
	    RECT 1404.6000 284.7000 1404.9000 286.2000 ;
	    RECT 1393.8000 284.4000 1395.0000 284.5500 ;
	    RECT 1398.6000 284.4000 1399.8000 284.5500 ;
	    RECT 1324.5000 282.3000 1326.9000 282.6000 ;
	    RECT 1365.3000 282.3000 1367.7001 282.6000 ;
	    RECT 1324.5000 281.7000 1327.2001 282.3000 ;
	    RECT 1285.8000 278.5500 1294.0500 279.4500 ;
	    RECT 1285.8000 278.4000 1287.0000 278.5500 ;
	    RECT 1276.2001 277.2000 1277.4000 277.5000 ;
	    RECT 1276.2001 273.3000 1277.4000 276.3000 ;
	    RECT 1295.4000 273.3000 1296.6000 280.5000 ;
	    RECT 1298.1000 280.2000 1301.4000 281.1000 ;
	    RECT 1297.8000 273.3000 1299.0000 279.3000 ;
	    RECT 1300.2001 273.3000 1301.4000 280.2000 ;
	    RECT 1326.0000 273.3000 1327.2001 281.7000 ;
	    RECT 1331.4000 273.3000 1332.6000 282.3000 ;
	    RECT 1365.3000 281.7000 1368.0000 282.3000 ;
	    RECT 1366.8000 273.3000 1368.0000 281.7000 ;
	    RECT 1372.2001 273.3000 1373.4000 282.3000 ;
	    RECT 1398.6000 278.4000 1399.8000 279.6000 ;
	    RECT 1401.3000 279.3000 1402.2001 284.7000 ;
	    RECT 1405.8000 284.4000 1407.0000 285.6000 ;
	    RECT 1403.4000 283.5000 1404.6000 283.8000 ;
	    RECT 1422.6000 283.5000 1423.8000 299.7000 ;
	    RECT 1446.6000 293.7000 1447.8000 299.7000 ;
	    RECT 1449.0000 294.3000 1450.2001 299.7000 ;
	    RECT 1446.9000 293.4000 1447.8000 293.7000 ;
	    RECT 1451.4000 293.7000 1452.6000 299.7000 ;
	    RECT 1453.8000 293.7000 1455.0000 299.7000 ;
	    RECT 1477.8000 293.7000 1479.0000 299.7000 ;
	    RECT 1480.2001 293.7000 1481.4000 299.7000 ;
	    RECT 1482.6000 294.3000 1483.8000 299.7000 ;
	    RECT 1451.4000 293.4000 1452.3000 293.7000 ;
	    RECT 1446.9000 292.5000 1452.3000 293.4000 ;
	    RECT 1480.5000 293.4000 1481.4000 293.7000 ;
	    RECT 1485.0000 293.7000 1486.2001 299.7000 ;
	    RECT 1485.0000 293.4000 1485.9000 293.7000 ;
	    RECT 1480.5000 292.5000 1485.9000 293.4000 ;
	    RECT 1446.9000 289.5000 1447.8000 292.5000 ;
	    RECT 1449.0000 291.4500 1450.2001 291.6000 ;
	    RECT 1465.8000 291.4500 1467.0000 291.6000 ;
	    RECT 1482.6000 291.4500 1483.8000 291.6000 ;
	    RECT 1449.0000 290.5500 1483.8000 291.4500 ;
	    RECT 1449.0000 290.4000 1450.2001 290.5500 ;
	    RECT 1465.8000 290.4000 1467.0000 290.5500 ;
	    RECT 1482.6000 290.4000 1483.8000 290.5500 ;
	    RECT 1485.0000 289.5000 1485.9000 292.5000 ;
	    RECT 1449.0000 289.2000 1450.2001 289.5000 ;
	    RECT 1482.6000 289.2000 1483.8000 289.5000 ;
	    RECT 1511.4000 288.6000 1512.6000 299.7000 ;
	    RECT 1513.8000 289.5000 1515.0000 299.7000 ;
	    RECT 1516.2001 288.6000 1517.4000 299.7000 ;
	    RECT 1446.6000 287.4000 1447.8000 288.6000 ;
	    RECT 1453.8000 288.4500 1455.0000 288.6000 ;
	    RECT 1477.8000 288.4500 1479.0000 288.6000 ;
	    RECT 1453.8000 287.5500 1479.0000 288.4500 ;
	    RECT 1453.8000 287.4000 1455.0000 287.5500 ;
	    RECT 1477.8000 287.4000 1479.0000 287.5500 ;
	    RECT 1485.0000 288.4500 1486.2001 288.6000 ;
	    RECT 1506.6000 288.4500 1507.8000 288.6000 ;
	    RECT 1485.0000 287.5500 1507.8000 288.4500 ;
	    RECT 1511.4000 287.7000 1517.4000 288.6000 ;
	    RECT 1518.6000 287.7000 1519.8000 299.7000 ;
	    RECT 1485.0000 287.4000 1486.2001 287.5500 ;
	    RECT 1506.6000 287.4000 1507.8000 287.5500 ;
	    RECT 1518.6000 286.5000 1519.5000 287.7000 ;
	    RECT 1542.6000 286.8000 1543.8000 299.7000 ;
	    RECT 1546.5000 287.7000 1547.7001 299.7000 ;
	    RECT 1548.9000 288.6000 1550.1000 299.7000 ;
	    RECT 1548.9000 287.7000 1551.0000 288.6000 ;
	    RECT 1446.9000 282.6000 1447.8000 286.5000 ;
	    RECT 1453.8000 286.2000 1455.0000 286.5000 ;
	    RECT 1477.8000 286.2000 1479.0000 286.5000 ;
	    RECT 1450.2001 284.4000 1450.5000 285.6000 ;
	    RECT 1451.4000 284.4000 1452.6000 285.6000 ;
	    RECT 1480.2001 284.4000 1481.4000 285.6000 ;
	    RECT 1482.3000 284.4000 1482.6000 285.6000 ;
	    RECT 1485.0000 282.6000 1485.9000 286.5000 ;
	    RECT 1542.6000 286.2000 1548.6000 286.8000 ;
	    RECT 1550.1000 286.5000 1551.0000 287.7000 ;
	    RECT 1511.4000 284.4000 1512.6000 285.6000 ;
	    RECT 1513.5000 284.7000 1513.8000 286.2000 ;
	    RECT 1542.6000 285.9000 1548.9000 286.2000 ;
	    RECT 1516.2001 284.7000 1517.7001 285.6000 ;
	    RECT 1518.6000 285.4500 1519.8000 285.6000 ;
	    RECT 1540.2001 285.4500 1541.4000 285.6000 ;
	    RECT 1513.8000 283.5000 1515.0000 283.8000 ;
	    RECT 1403.4000 281.4000 1404.6000 282.6000 ;
	    RECT 1422.6000 282.4500 1423.8000 282.6000 ;
	    RECT 1441.8000 282.4500 1443.0000 282.6000 ;
	    RECT 1422.6000 281.5500 1443.0000 282.4500 ;
	    RECT 1446.9000 282.3000 1449.3000 282.6000 ;
	    RECT 1483.5000 282.3000 1485.9000 282.6000 ;
	    RECT 1446.9000 281.7000 1449.6000 282.3000 ;
	    RECT 1422.6000 281.4000 1423.8000 281.5500 ;
	    RECT 1441.8000 281.4000 1443.0000 281.5500 ;
	    RECT 1398.9000 277.2000 1400.1000 277.5000 ;
	    RECT 1398.6000 273.3000 1399.8000 276.3000 ;
	    RECT 1401.0000 273.3000 1402.2001 279.3000 ;
	    RECT 1404.9000 273.3000 1406.1000 279.3000 ;
	    RECT 1420.2001 278.4000 1421.4000 279.6000 ;
	    RECT 1420.2001 277.2000 1421.4000 277.5000 ;
	    RECT 1420.2001 273.3000 1421.4000 276.3000 ;
	    RECT 1422.6000 273.3000 1423.8000 280.5000 ;
	    RECT 1448.4000 273.3000 1449.6000 281.7000 ;
	    RECT 1453.8000 273.3000 1455.0000 282.3000 ;
	    RECT 1477.8000 273.3000 1479.0000 282.3000 ;
	    RECT 1483.2001 281.7000 1485.9000 282.3000 ;
	    RECT 1483.2001 273.3000 1484.4000 281.7000 ;
	    RECT 1513.8000 281.4000 1515.0000 282.6000 ;
	    RECT 1516.2001 279.3000 1517.1000 284.7000 ;
	    RECT 1518.6000 284.5500 1541.4000 285.4500 ;
	    RECT 1547.7001 285.0000 1548.9000 285.9000 ;
	    RECT 1518.6000 284.4000 1519.8000 284.5500 ;
	    RECT 1540.2001 284.4000 1541.4000 284.5500 ;
	    RECT 1545.6000 283.5000 1546.8000 283.8000 ;
	    RECT 1537.8000 282.4500 1539.0000 282.6000 ;
	    RECT 1545.0000 282.4500 1546.2001 282.6000 ;
	    RECT 1537.8000 281.5500 1546.2001 282.4500 ;
	    RECT 1537.8000 281.4000 1539.0000 281.5500 ;
	    RECT 1545.0000 281.4000 1546.2001 281.5500 ;
	    RECT 1548.0000 280.5000 1548.9000 285.0000 ;
	    RECT 1549.8000 284.4000 1551.0000 285.6000 ;
	    RECT 1545.3000 279.6000 1548.9000 280.5000 ;
	    RECT 1518.6000 279.4500 1519.8000 279.6000 ;
	    RECT 1540.2001 279.4500 1541.4000 279.6000 ;
	    RECT 1512.3000 273.3000 1513.5000 279.3000 ;
	    RECT 1516.2001 273.3000 1517.4000 279.3000 ;
	    RECT 1518.6000 278.5500 1541.4000 279.4500 ;
	    RECT 1518.6000 278.4000 1519.8000 278.5500 ;
	    RECT 1540.2001 278.4000 1541.4000 278.5500 ;
	    RECT 1542.6000 278.4000 1543.8000 279.6000 ;
	    RECT 1518.3000 277.2000 1519.5000 277.5000 ;
	    RECT 1542.6000 277.2000 1543.8000 277.5000 ;
	    RECT 1545.3000 276.3000 1546.2001 279.6000 ;
	    RECT 1550.1000 279.3000 1551.0000 283.5000 ;
	    RECT 1518.6000 273.3000 1519.8000 276.3000 ;
	    RECT 1542.6000 273.3000 1543.8000 276.3000 ;
	    RECT 1545.0000 273.3000 1546.2001 276.3000 ;
	    RECT 1547.4000 273.3000 1548.6000 278.7000 ;
	    RECT 1549.8000 273.3000 1551.0000 279.3000 ;
	    RECT 1.2000 270.6000 1569.0000 272.4000 ;
	    RECT 124.2000 260.7000 125.4000 269.7000 ;
	    RECT 129.0000 263.7000 130.2000 269.7000 ;
	    RECT 133.8000 264.9000 135.0000 269.7000 ;
	    RECT 136.2000 265.5000 137.4000 269.7000 ;
	    RECT 138.6000 265.5000 139.8000 269.7000 ;
	    RECT 141.0000 265.5000 142.2000 269.7000 ;
	    RECT 143.4000 266.7000 144.6000 269.7000 ;
	    RECT 145.8000 265.5000 147.0000 269.7000 ;
	    RECT 148.2000 266.7000 149.4000 269.7000 ;
	    RECT 150.6000 265.5000 151.8000 269.7000 ;
	    RECT 153.0000 265.5000 154.2000 269.7000 ;
	    RECT 155.4000 265.5000 156.6000 269.7000 ;
	    RECT 157.8000 265.5000 159.0000 269.7000 ;
	    RECT 131.1000 263.7000 135.0000 264.9000 ;
	    RECT 160.2000 264.9000 161.4000 269.7000 ;
	    RECT 140.1000 263.7000 147.0000 264.6000 ;
	    RECT 131.1000 262.8000 132.3000 263.7000 ;
	    RECT 127.8000 261.6000 132.3000 262.8000 ;
	    RECT 124.2000 259.5000 137.4000 260.7000 ;
	    RECT 140.1000 260.1000 141.3000 263.7000 ;
	    RECT 145.8000 263.4000 147.0000 263.7000 ;
	    RECT 148.2000 263.4000 149.4000 264.6000 ;
	    RECT 150.3000 263.4000 150.6000 264.6000 ;
	    RECT 155.1000 263.4000 156.6000 264.6000 ;
	    RECT 160.2000 263.7000 163.8000 264.9000 ;
	    RECT 165.0000 263.7000 166.2000 269.7000 ;
	    RECT 143.4000 262.5000 144.6000 262.8000 ;
	    RECT 145.8000 262.2000 147.0000 262.5000 ;
	    RECT 143.4000 260.4000 144.6000 261.6000 ;
	    RECT 145.8000 261.3000 152.4000 262.2000 ;
	    RECT 151.2000 261.0000 152.4000 261.3000 ;
	    RECT 124.2000 251.1000 125.4000 259.5000 ;
	    RECT 138.3000 258.9000 141.3000 260.1000 ;
	    RECT 147.0000 258.9000 151.8000 260.1000 ;
	    RECT 155.4000 259.2000 156.6000 263.4000 ;
	    RECT 162.6000 262.8000 163.8000 263.7000 ;
	    RECT 162.6000 261.9000 165.3000 262.8000 ;
	    RECT 164.1000 260.1000 165.3000 261.9000 ;
	    RECT 169.8000 261.9000 171.0000 269.7000 ;
	    RECT 172.2000 264.0000 173.4000 269.7000 ;
	    RECT 174.6000 266.7000 175.8000 269.7000 ;
	    RECT 172.2000 262.8000 173.7000 264.0000 ;
	    RECT 232.2000 263.7000 233.4000 269.7000 ;
	    RECT 169.8000 261.0000 171.6000 261.9000 ;
	    RECT 164.1000 258.9000 169.8000 260.1000 ;
	    RECT 126.3000 258.0000 127.5000 258.3000 ;
	    RECT 126.3000 257.1000 132.9000 258.0000 ;
	    RECT 133.8000 257.4000 135.0000 258.6000 ;
	    RECT 160.2000 258.0000 161.4000 258.9000 ;
	    RECT 170.7000 258.0000 171.6000 261.0000 ;
	    RECT 135.9000 257.1000 161.4000 258.0000 ;
	    RECT 170.4000 257.1000 171.6000 258.0000 ;
	    RECT 168.3000 256.2000 169.5000 256.5000 ;
	    RECT 129.0000 254.4000 130.2000 255.6000 ;
	    RECT 131.1000 255.3000 169.5000 256.2000 ;
	    RECT 134.1000 255.0000 135.3000 255.3000 ;
	    RECT 170.4000 254.4000 171.3000 257.1000 ;
	    RECT 172.5000 256.2000 173.7000 262.8000 ;
	    RECT 234.6000 262.8000 235.8000 269.7000 ;
	    RECT 237.0000 263.7000 238.2000 269.7000 ;
	    RECT 239.4000 262.8000 240.6000 269.7000 ;
	    RECT 241.8000 263.7000 243.0000 269.7000 ;
	    RECT 244.2000 262.8000 245.4000 269.7000 ;
	    RECT 246.6000 263.7000 247.8000 269.7000 ;
	    RECT 249.0000 262.8000 250.2000 269.7000 ;
	    RECT 251.4000 263.7000 252.6000 269.7000 ;
	    RECT 234.6000 261.6000 237.3000 262.8000 ;
	    RECT 239.4000 261.6000 242.7000 262.8000 ;
	    RECT 244.2000 261.6000 247.5000 262.8000 ;
	    RECT 249.0000 261.6000 252.6000 262.8000 ;
	    RECT 265.8000 262.5000 267.0000 269.7000 ;
	    RECT 268.2000 266.7000 269.4000 269.7000 ;
	    RECT 268.2000 265.5000 269.4000 265.8000 ;
	    RECT 268.2000 263.4000 269.4000 264.6000 ;
	    RECT 292.2000 263.7000 293.4000 269.7000 ;
	    RECT 294.6000 264.0000 295.8000 269.7000 ;
	    RECT 297.0000 264.9000 298.2000 269.7000 ;
	    RECT 299.4000 264.0000 300.6000 269.7000 ;
	    RECT 294.6000 263.7000 300.6000 264.0000 ;
	    RECT 292.5000 262.5000 293.4000 263.7000 ;
	    RECT 294.9000 263.1000 300.3000 263.7000 ;
	    RECT 313.8000 262.5000 315.0000 269.7000 ;
	    RECT 316.2000 266.7000 317.4000 269.7000 ;
	    RECT 316.2000 265.5000 317.4000 265.8000 ;
	    RECT 336.3000 264.6000 337.5000 269.7000 ;
	    RECT 316.2000 264.4500 317.4000 264.6000 ;
	    RECT 330.6000 264.4500 331.8000 264.6000 ;
	    RECT 333.0000 264.4500 334.2000 264.6000 ;
	    RECT 316.2000 263.5500 334.2000 264.4500 ;
	    RECT 336.3000 263.7000 339.0000 264.6000 ;
	    RECT 340.2000 263.7000 341.4000 269.7000 ;
	    RECT 366.6000 264.0000 367.8000 269.7000 ;
	    RECT 369.0000 264.9000 370.2000 269.7000 ;
	    RECT 371.4000 264.0000 372.6000 269.7000 ;
	    RECT 366.6000 263.7000 372.6000 264.0000 ;
	    RECT 373.8000 263.7000 375.0000 269.7000 ;
	    RECT 385.8000 266.7000 387.0000 269.7000 ;
	    RECT 385.8000 265.5000 387.0000 265.8000 ;
	    RECT 316.2000 263.4000 317.4000 263.5500 ;
	    RECT 330.6000 263.4000 331.8000 263.5500 ;
	    RECT 333.0000 263.4000 334.2000 263.5500 ;
	    RECT 229.8000 261.4500 231.0000 261.6000 ;
	    RECT 232.2000 261.4500 233.4000 261.6000 ;
	    RECT 229.8000 260.5500 233.4000 261.4500 ;
	    RECT 236.1000 260.7000 237.3000 261.6000 ;
	    RECT 241.5000 260.7000 242.7000 261.6000 ;
	    RECT 246.3000 260.7000 247.5000 261.6000 ;
	    RECT 229.8000 260.4000 231.0000 260.5500 ;
	    RECT 232.2000 260.4000 233.4000 260.5500 ;
	    RECT 234.3000 259.5000 234.9000 260.7000 ;
	    RECT 236.1000 259.5000 240.0000 260.7000 ;
	    RECT 241.5000 259.5000 245.1000 260.7000 ;
	    RECT 246.3000 259.5000 250.2000 260.7000 ;
	    RECT 251.4000 259.5000 252.6000 261.6000 ;
	    RECT 253.8000 261.4500 255.0000 261.6000 ;
	    RECT 265.8000 261.4500 267.0000 261.6000 ;
	    RECT 282.6000 261.4500 283.8000 261.6000 ;
	    RECT 253.8000 260.5500 283.8000 261.4500 ;
	    RECT 253.8000 260.4000 255.0000 260.5500 ;
	    RECT 265.8000 260.4000 267.0000 260.5500 ;
	    RECT 282.6000 260.4000 283.8000 260.5500 ;
	    RECT 292.2000 260.4000 293.4000 261.6000 ;
	    RECT 294.3000 260.4000 296.1000 261.6000 ;
	    RECT 298.2000 260.7000 298.5000 262.2000 ;
	    RECT 299.4000 260.4000 300.6000 261.6000 ;
	    RECT 313.8000 261.4500 315.0000 261.6000 ;
	    RECT 301.9500 260.5500 315.0000 261.4500 ;
	    RECT 236.1000 257.4000 237.3000 259.5000 ;
	    RECT 241.5000 257.4000 242.7000 259.5000 ;
	    RECT 246.3000 257.4000 247.5000 259.5000 ;
	    RECT 251.4000 257.4000 252.6000 258.6000 ;
	    RECT 138.6000 254.1000 139.8000 254.4000 ;
	    RECT 131.7000 253.5000 139.8000 254.1000 ;
	    RECT 130.5000 253.2000 139.8000 253.5000 ;
	    RECT 141.3000 253.5000 154.2000 254.4000 ;
	    RECT 126.6000 252.0000 129.0000 253.2000 ;
	    RECT 130.5000 252.3000 132.6000 253.2000 ;
	    RECT 141.3000 252.3000 142.2000 253.5000 ;
	    RECT 153.0000 253.2000 154.2000 253.5000 ;
	    RECT 157.8000 253.5000 171.3000 254.4000 ;
	    RECT 172.2000 255.0000 173.7000 256.2000 ;
	    RECT 234.6000 256.2000 237.3000 257.4000 ;
	    RECT 239.4000 256.2000 242.7000 257.4000 ;
	    RECT 244.2000 256.2000 247.5000 257.4000 ;
	    RECT 249.0000 256.5000 250.5000 257.4000 ;
	    RECT 249.0000 256.2000 252.6000 256.5000 ;
	    RECT 172.2000 253.5000 173.4000 255.0000 ;
	    RECT 157.8000 253.2000 159.0000 253.5000 ;
	    RECT 128.1000 251.4000 129.0000 252.0000 ;
	    RECT 133.5000 251.4000 142.2000 252.3000 ;
	    RECT 143.1000 251.4000 147.0000 252.6000 ;
	    RECT 124.2000 250.2000 127.2000 251.1000 ;
	    RECT 128.1000 250.2000 134.4000 251.4000 ;
	    RECT 126.3000 249.3000 127.2000 250.2000 ;
	    RECT 124.2000 243.3000 125.4000 249.3000 ;
	    RECT 126.3000 248.4000 127.8000 249.3000 ;
	    RECT 126.6000 243.3000 127.8000 248.4000 ;
	    RECT 129.0000 242.4000 130.2000 249.3000 ;
	    RECT 131.4000 243.3000 132.6000 250.2000 ;
	    RECT 133.8000 243.3000 135.0000 249.3000 ;
	    RECT 136.2000 243.3000 137.4000 247.5000 ;
	    RECT 138.6000 243.3000 139.8000 247.5000 ;
	    RECT 141.0000 243.3000 142.2000 250.5000 ;
	    RECT 143.4000 243.3000 144.6000 249.3000 ;
	    RECT 145.8000 243.3000 147.0000 250.5000 ;
	    RECT 148.2000 243.3000 149.4000 249.3000 ;
	    RECT 150.6000 243.3000 151.8000 252.6000 ;
	    RECT 162.6000 251.4000 166.5000 252.6000 ;
	    RECT 155.4000 250.2000 161.7000 251.4000 ;
	    RECT 153.0000 243.3000 154.2000 247.5000 ;
	    RECT 155.4000 243.3000 156.6000 247.5000 ;
	    RECT 157.8000 243.3000 159.0000 247.5000 ;
	    RECT 160.2000 243.3000 161.4000 249.3000 ;
	    RECT 162.6000 243.3000 163.8000 251.4000 ;
	    RECT 170.4000 251.1000 171.3000 253.5000 ;
	    RECT 172.2000 252.4500 173.4000 252.6000 ;
	    RECT 177.0000 252.4500 178.2000 252.6000 ;
	    RECT 172.2000 251.5500 178.2000 252.4500 ;
	    RECT 172.2000 251.4000 173.4000 251.5500 ;
	    RECT 177.0000 251.4000 178.2000 251.5500 ;
	    RECT 167.4000 250.2000 171.3000 251.1000 ;
	    RECT 165.0000 243.3000 166.2000 249.3000 ;
	    RECT 167.4000 243.3000 168.6000 250.2000 ;
	    RECT 169.8000 243.3000 171.0000 249.3000 ;
	    RECT 172.2000 243.3000 173.4000 250.5000 ;
	    RECT 174.6000 243.3000 175.8000 249.3000 ;
	    RECT 232.2000 243.3000 233.4000 255.3000 ;
	    RECT 234.6000 243.3000 235.8000 256.2000 ;
	    RECT 237.0000 243.3000 238.2000 255.3000 ;
	    RECT 239.4000 243.3000 240.6000 256.2000 ;
	    RECT 241.8000 243.3000 243.0000 255.3000 ;
	    RECT 244.2000 243.3000 245.4000 256.2000 ;
	    RECT 246.6000 243.3000 247.8000 255.3000 ;
	    RECT 249.0000 243.3000 250.2000 256.2000 ;
	    RECT 251.4000 243.3000 252.6000 255.3000 ;
	    RECT 265.8000 243.3000 267.0000 259.5000 ;
	    RECT 280.2000 255.4500 281.4000 255.6000 ;
	    RECT 292.2000 255.4500 293.4000 255.6000 ;
	    RECT 280.2000 254.5500 293.4000 255.4500 ;
	    RECT 280.2000 254.4000 281.4000 254.5500 ;
	    RECT 292.2000 254.4000 293.4000 254.5500 ;
	    RECT 295.2000 255.3000 296.1000 260.4000 ;
	    RECT 297.0000 259.5000 298.2000 259.8000 ;
	    RECT 297.0000 258.4500 298.2000 258.6000 ;
	    RECT 301.9500 258.4500 302.8500 260.5500 ;
	    RECT 313.8000 260.4000 315.0000 260.5500 ;
	    RECT 337.8000 259.5000 339.0000 263.7000 ;
	    RECT 366.9000 263.1000 372.3000 263.7000 ;
	    RECT 340.2000 262.5000 341.4000 262.8000 ;
	    RECT 373.8000 262.5000 374.7000 263.7000 ;
	    RECT 385.8000 263.4000 387.0000 264.6000 ;
	    RECT 388.2000 262.5000 389.4000 269.7000 ;
	    RECT 402.6000 262.5000 403.8000 269.7000 ;
	    RECT 405.0000 266.7000 406.2000 269.7000 ;
	    RECT 405.0000 265.5000 406.2000 265.8000 ;
	    RECT 405.0000 264.4500 406.2000 264.6000 ;
	    RECT 479.4000 264.4500 480.6000 264.6000 ;
	    RECT 405.0000 263.5500 480.6000 264.4500 ;
	    RECT 405.0000 263.4000 406.2000 263.5500 ;
	    RECT 479.4000 263.4000 480.6000 263.5500 ;
	    RECT 340.2000 261.4500 341.4000 261.6000 ;
	    RECT 366.6000 261.4500 367.8000 261.6000 ;
	    RECT 340.2000 260.5500 367.8000 261.4500 ;
	    RECT 368.7000 260.7000 369.0000 262.2000 ;
	    RECT 340.2000 260.4000 341.4000 260.5500 ;
	    RECT 366.6000 260.4000 367.8000 260.5500 ;
	    RECT 371.1000 260.4000 372.9000 261.6000 ;
	    RECT 373.8000 260.4000 375.0000 261.6000 ;
	    RECT 376.2000 261.4500 377.4000 261.6000 ;
	    RECT 388.2000 261.4500 389.4000 261.6000 ;
	    RECT 376.2000 260.5500 389.4000 261.4500 ;
	    RECT 376.2000 260.4000 377.4000 260.5500 ;
	    RECT 388.2000 260.4000 389.4000 260.5500 ;
	    RECT 402.6000 261.4500 403.8000 261.6000 ;
	    RECT 445.8000 261.4500 447.0000 261.6000 ;
	    RECT 402.6000 260.5500 447.0000 261.4500 ;
	    RECT 402.6000 260.4000 403.8000 260.5500 ;
	    RECT 445.8000 260.4000 447.0000 260.5500 ;
	    RECT 539.4000 260.7000 540.6000 269.7000 ;
	    RECT 544.2000 263.7000 545.4000 269.7000 ;
	    RECT 549.0000 264.9000 550.2000 269.7000 ;
	    RECT 551.4000 265.5000 552.6000 269.7000 ;
	    RECT 553.8000 265.5000 555.0000 269.7000 ;
	    RECT 556.2000 265.5000 557.4000 269.7000 ;
	    RECT 558.6000 266.7000 559.8000 269.7000 ;
	    RECT 561.0000 265.5000 562.2000 269.7000 ;
	    RECT 563.4000 266.7000 564.6000 269.7000 ;
	    RECT 565.8000 265.5000 567.0000 269.7000 ;
	    RECT 568.2000 265.5000 569.4000 269.7000 ;
	    RECT 570.6000 265.5000 571.8000 269.7000 ;
	    RECT 573.0000 265.5000 574.2000 269.7000 ;
	    RECT 546.3000 263.7000 550.2000 264.9000 ;
	    RECT 575.4000 264.9000 576.6000 269.7000 ;
	    RECT 555.3000 263.7000 562.2000 264.6000 ;
	    RECT 546.3000 262.8000 547.5000 263.7000 ;
	    RECT 543.0000 261.6000 547.5000 262.8000 ;
	    RECT 369.0000 259.5000 370.2000 259.8000 ;
	    RECT 297.0000 257.5500 302.8500 258.4500 ;
	    RECT 297.0000 257.4000 298.2000 257.5500 ;
	    RECT 295.2000 254.4000 296.7000 255.3000 ;
	    RECT 293.4000 252.6000 294.3000 253.5000 ;
	    RECT 293.4000 251.4000 294.6000 252.6000 ;
	    RECT 268.2000 243.3000 269.4000 249.3000 ;
	    RECT 293.1000 243.3000 294.3000 249.3000 ;
	    RECT 295.5000 243.3000 296.7000 254.4000 ;
	    RECT 299.4000 243.3000 300.6000 255.3000 ;
	    RECT 313.8000 243.3000 315.0000 259.5000 ;
	    RECT 337.8000 258.4500 339.0000 258.6000 ;
	    RECT 366.6000 258.4500 367.8000 258.6000 ;
	    RECT 337.8000 257.5500 367.8000 258.4500 ;
	    RECT 337.8000 257.4000 339.0000 257.5500 ;
	    RECT 366.6000 257.4000 367.8000 257.5500 ;
	    RECT 369.0000 257.4000 370.2000 258.6000 ;
	    RECT 333.0000 255.4500 334.2000 255.6000 ;
	    RECT 335.4000 255.4500 336.6000 255.6000 ;
	    RECT 333.0000 254.5500 336.6000 255.4500 ;
	    RECT 333.0000 254.4000 334.2000 254.5500 ;
	    RECT 335.4000 254.4000 336.6000 254.5500 ;
	    RECT 335.4000 253.2000 336.6000 253.5000 ;
	    RECT 316.2000 243.3000 317.4000 249.3000 ;
	    RECT 335.4000 243.3000 336.6000 249.3000 ;
	    RECT 337.8000 243.3000 339.0000 256.5000 ;
	    RECT 371.1000 255.3000 372.0000 260.4000 ;
	    RECT 373.9500 258.4500 374.8500 260.4000 ;
	    RECT 539.4000 259.5000 552.6000 260.7000 ;
	    RECT 555.3000 260.1000 556.5000 263.7000 ;
	    RECT 561.0000 263.4000 562.2000 263.7000 ;
	    RECT 563.4000 263.4000 564.6000 264.6000 ;
	    RECT 565.5000 263.4000 565.8000 264.6000 ;
	    RECT 570.3000 263.4000 571.8000 264.6000 ;
	    RECT 575.4000 263.7000 579.0000 264.9000 ;
	    RECT 580.2000 263.7000 581.4000 269.7000 ;
	    RECT 558.6000 262.5000 559.8000 262.8000 ;
	    RECT 561.0000 262.2000 562.2000 262.5000 ;
	    RECT 558.6000 260.4000 559.8000 261.6000 ;
	    RECT 561.0000 261.3000 567.6000 262.2000 ;
	    RECT 566.4000 261.0000 567.6000 261.3000 ;
	    RECT 383.4000 258.4500 384.6000 258.6000 ;
	    RECT 373.9500 257.5500 384.6000 258.4500 ;
	    RECT 383.4000 257.4000 384.6000 257.5500 ;
	    RECT 340.2000 243.3000 341.4000 249.3000 ;
	    RECT 366.6000 243.3000 367.8000 255.3000 ;
	    RECT 370.5000 254.4000 372.0000 255.3000 ;
	    RECT 373.8000 254.4000 375.0000 255.6000 ;
	    RECT 370.5000 243.3000 371.7000 254.4000 ;
	    RECT 372.9000 252.6000 373.8000 253.5000 ;
	    RECT 372.6000 251.4000 373.8000 252.6000 ;
	    RECT 372.9000 243.3000 374.1000 249.3000 ;
	    RECT 385.8000 243.3000 387.0000 249.3000 ;
	    RECT 388.2000 243.3000 389.4000 259.5000 ;
	    RECT 402.6000 243.3000 403.8000 259.5000 ;
	    RECT 539.4000 251.1000 540.6000 259.5000 ;
	    RECT 553.5000 258.9000 556.5000 260.1000 ;
	    RECT 562.2000 258.9000 567.0000 260.1000 ;
	    RECT 570.6000 259.2000 571.8000 263.4000 ;
	    RECT 577.8000 262.8000 579.0000 263.7000 ;
	    RECT 577.8000 261.9000 580.5000 262.8000 ;
	    RECT 579.3000 260.1000 580.5000 261.9000 ;
	    RECT 585.0000 261.9000 586.2000 269.7000 ;
	    RECT 587.4000 264.0000 588.6000 269.7000 ;
	    RECT 589.8000 266.7000 591.0000 269.7000 ;
	    RECT 587.4000 262.8000 588.9000 264.0000 ;
	    RECT 613.8000 263.7000 615.0000 269.7000 ;
	    RECT 616.2000 264.0000 617.4000 269.7000 ;
	    RECT 618.6000 264.9000 619.8000 269.7000 ;
	    RECT 621.0000 264.0000 622.2000 269.7000 ;
	    RECT 616.2000 263.7000 622.2000 264.0000 ;
	    RECT 585.0000 261.0000 586.8000 261.9000 ;
	    RECT 579.3000 258.9000 585.0000 260.1000 ;
	    RECT 541.5000 258.0000 542.7000 258.3000 ;
	    RECT 541.5000 257.1000 548.1000 258.0000 ;
	    RECT 549.0000 257.4000 550.2000 258.6000 ;
	    RECT 575.4000 258.0000 576.6000 258.9000 ;
	    RECT 585.9000 258.0000 586.8000 261.0000 ;
	    RECT 551.1000 257.1000 576.6000 258.0000 ;
	    RECT 585.6000 257.1000 586.8000 258.0000 ;
	    RECT 583.5000 256.2000 584.7000 256.5000 ;
	    RECT 544.2000 254.4000 545.4000 255.6000 ;
	    RECT 546.3000 255.3000 584.7000 256.2000 ;
	    RECT 549.3000 255.0000 550.5000 255.3000 ;
	    RECT 585.6000 254.4000 586.5000 257.1000 ;
	    RECT 587.7000 256.2000 588.9000 262.8000 ;
	    RECT 614.1000 262.5000 615.0000 263.7000 ;
	    RECT 616.5000 263.1000 621.9000 263.7000 ;
	    RECT 697.8000 262.5000 699.0000 269.7000 ;
	    RECT 700.2000 263.7000 701.4000 269.7000 ;
	    RECT 704.4000 267.6000 705.6000 269.7000 ;
	    RECT 702.6000 266.7000 705.6000 267.6000 ;
	    RECT 708.3000 266.7000 709.8000 269.7000 ;
	    RECT 711.0000 266.7000 712.2000 269.7000 ;
	    RECT 713.4000 266.7000 714.6000 269.7000 ;
	    RECT 717.3000 267.6000 719.1000 269.7000 ;
	    RECT 717.0000 266.7000 719.1000 267.6000 ;
	    RECT 702.6000 265.5000 703.8000 266.7000 ;
	    RECT 711.0000 265.8000 711.9000 266.7000 ;
	    RECT 705.0000 264.6000 706.2000 265.8000 ;
	    RECT 707.7000 264.9000 711.9000 265.8000 ;
	    RECT 717.0000 265.5000 718.2000 266.7000 ;
	    RECT 707.7000 264.6000 708.9000 264.9000 ;
	    RECT 589.8000 261.4500 591.0000 261.6000 ;
	    RECT 613.8000 261.4500 615.0000 261.6000 ;
	    RECT 589.8000 260.5500 615.0000 261.4500 ;
	    RECT 589.8000 260.4000 591.0000 260.5500 ;
	    RECT 613.8000 260.4000 615.0000 260.5500 ;
	    RECT 615.9000 260.4000 617.7000 261.6000 ;
	    RECT 619.8000 260.7000 620.1000 262.2000 ;
	    RECT 621.0000 260.4000 622.2000 261.6000 ;
	    RECT 699.0000 260.4000 699.3000 261.6000 ;
	    RECT 700.2000 260.4000 701.4000 261.6000 ;
	    RECT 705.3000 261.3000 706.2000 264.6000 ;
	    RECT 721.8000 264.0000 723.0000 269.7000 ;
	    RECT 719.7000 263.1000 720.9000 263.4000 ;
	    RECT 724.2000 263.1000 725.4000 269.7000 ;
	    RECT 748.2000 263.7000 749.4000 269.7000 ;
	    RECT 750.6000 264.0000 751.8000 269.7000 ;
	    RECT 753.0000 264.9000 754.2000 269.7000 ;
	    RECT 755.4000 264.0000 756.6000 269.7000 ;
	    RECT 750.6000 263.7000 756.6000 264.0000 ;
	    RECT 719.7000 262.2000 725.4000 263.1000 ;
	    RECT 748.5000 262.5000 749.4000 263.7000 ;
	    RECT 750.9000 263.1000 756.3000 263.7000 ;
	    RECT 769.8000 262.5000 771.0000 269.7000 ;
	    RECT 772.2000 266.7000 773.4000 269.7000 ;
	    RECT 772.2000 265.5000 773.4000 265.8000 ;
	    RECT 772.2000 264.4500 773.4000 264.6000 ;
	    RECT 789.0000 264.4500 790.2000 264.6000 ;
	    RECT 772.2000 263.5500 790.2000 264.4500 ;
	    RECT 791.4000 263.7000 792.6000 269.7000 ;
	    RECT 795.3000 264.6000 796.5000 269.7000 ;
	    RECT 793.8000 263.7000 796.5000 264.6000 ;
	    RECT 815.4000 263.7000 816.6000 269.7000 ;
	    RECT 819.3000 264.6000 820.5000 269.7000 ;
	    RECT 817.8000 263.7000 820.5000 264.6000 ;
	    RECT 772.2000 263.4000 773.4000 263.5500 ;
	    RECT 789.0000 263.4000 790.2000 263.5500 ;
	    RECT 791.4000 262.5000 792.6000 262.8000 ;
	    RECT 713.7000 261.3000 714.9000 261.6000 ;
	    RECT 702.3000 260.4000 715.5000 261.3000 ;
	    RECT 553.8000 254.1000 555.0000 254.4000 ;
	    RECT 546.9000 253.5000 555.0000 254.1000 ;
	    RECT 545.7000 253.2000 555.0000 253.5000 ;
	    RECT 556.5000 253.5000 569.4000 254.4000 ;
	    RECT 541.8000 252.0000 544.2000 253.2000 ;
	    RECT 545.7000 252.3000 547.8000 253.2000 ;
	    RECT 556.5000 252.3000 557.4000 253.5000 ;
	    RECT 568.2000 253.2000 569.4000 253.5000 ;
	    RECT 573.0000 253.5000 586.5000 254.4000 ;
	    RECT 587.4000 255.0000 588.9000 256.2000 ;
	    RECT 601.8000 255.4500 603.0000 255.6000 ;
	    RECT 613.8000 255.4500 615.0000 255.6000 ;
	    RECT 587.4000 253.5000 588.6000 255.0000 ;
	    RECT 601.8000 254.5500 615.0000 255.4500 ;
	    RECT 601.8000 254.4000 603.0000 254.5500 ;
	    RECT 613.8000 254.4000 615.0000 254.5500 ;
	    RECT 616.8000 255.3000 617.7000 260.4000 ;
	    RECT 703.5000 260.1000 704.7000 260.4000 ;
	    RECT 618.6000 259.5000 619.8000 259.8000 ;
	    RECT 701.1000 258.6000 702.3000 258.9000 ;
	    RECT 618.6000 257.4000 619.8000 258.6000 ;
	    RECT 701.1000 257.7000 706.5000 258.6000 ;
	    RECT 707.4000 257.4000 708.6000 258.6000 ;
	    RECT 697.8000 256.5000 706.2000 256.8000 ;
	    RECT 697.8000 256.2000 706.5000 256.5000 ;
	    RECT 697.8000 255.9000 712.5000 256.2000 ;
	    RECT 616.8000 254.4000 618.3000 255.3000 ;
	    RECT 573.0000 253.2000 574.2000 253.5000 ;
	    RECT 543.3000 251.4000 544.2000 252.0000 ;
	    RECT 548.7000 251.4000 557.4000 252.3000 ;
	    RECT 558.3000 251.4000 562.2000 252.6000 ;
	    RECT 539.4000 250.2000 542.4000 251.1000 ;
	    RECT 543.3000 250.2000 549.6000 251.4000 ;
	    RECT 489.0000 249.4500 490.2000 249.6000 ;
	    RECT 501.0000 249.4500 502.2000 249.6000 ;
	    RECT 405.0000 243.3000 406.2000 249.3000 ;
	    RECT 489.0000 248.5500 502.2000 249.4500 ;
	    RECT 541.5000 249.3000 542.4000 250.2000 ;
	    RECT 489.0000 248.4000 490.2000 248.5500 ;
	    RECT 501.0000 248.4000 502.2000 248.5500 ;
	    RECT 419.4000 246.4500 420.6000 246.6000 ;
	    RECT 431.4000 246.4500 432.6000 246.6000 ;
	    RECT 419.4000 245.5500 432.6000 246.4500 ;
	    RECT 419.4000 245.4000 420.6000 245.5500 ;
	    RECT 431.4000 245.4000 432.6000 245.5500 ;
	    RECT 539.4000 243.3000 540.6000 249.3000 ;
	    RECT 541.5000 248.4000 543.0000 249.3000 ;
	    RECT 541.8000 243.3000 543.0000 248.4000 ;
	    RECT 544.2000 242.4000 545.4000 249.3000 ;
	    RECT 546.6000 243.3000 547.8000 250.2000 ;
	    RECT 549.0000 243.3000 550.2000 249.3000 ;
	    RECT 551.4000 243.3000 552.6000 247.5000 ;
	    RECT 553.8000 243.3000 555.0000 247.5000 ;
	    RECT 556.2000 243.3000 557.4000 250.5000 ;
	    RECT 558.6000 243.3000 559.8000 249.3000 ;
	    RECT 561.0000 243.3000 562.2000 250.5000 ;
	    RECT 563.4000 243.3000 564.6000 249.3000 ;
	    RECT 565.8000 243.3000 567.0000 252.6000 ;
	    RECT 577.8000 251.4000 581.7000 252.6000 ;
	    RECT 570.6000 250.2000 576.9000 251.4000 ;
	    RECT 568.2000 243.3000 569.4000 247.5000 ;
	    RECT 570.6000 243.3000 571.8000 247.5000 ;
	    RECT 573.0000 243.3000 574.2000 247.5000 ;
	    RECT 575.4000 243.3000 576.6000 249.3000 ;
	    RECT 577.8000 243.3000 579.0000 251.4000 ;
	    RECT 585.6000 251.1000 586.5000 253.5000 ;
	    RECT 615.0000 252.6000 615.9000 253.5000 ;
	    RECT 587.4000 251.4000 588.6000 252.6000 ;
	    RECT 615.0000 251.4000 616.2000 252.6000 ;
	    RECT 582.6000 250.2000 586.5000 251.1000 ;
	    RECT 580.2000 243.3000 581.4000 249.3000 ;
	    RECT 582.6000 243.3000 583.8000 250.2000 ;
	    RECT 585.0000 243.3000 586.2000 249.3000 ;
	    RECT 587.4000 243.3000 588.6000 250.5000 ;
	    RECT 589.8000 243.3000 591.0000 249.3000 ;
	    RECT 614.7000 243.3000 615.9000 249.3000 ;
	    RECT 617.1000 243.3000 618.3000 254.4000 ;
	    RECT 621.0000 243.3000 622.2000 255.3000 ;
	    RECT 697.8000 243.3000 699.0000 255.9000 ;
	    RECT 705.3000 255.3000 712.5000 255.9000 ;
	    RECT 700.2000 243.3000 701.4000 255.0000 ;
	    RECT 702.6000 253.5000 710.7000 254.4000 ;
	    RECT 702.6000 253.2000 703.8000 253.5000 ;
	    RECT 709.5000 253.2000 710.7000 253.5000 ;
	    RECT 711.6000 253.5000 712.5000 255.3000 ;
	    RECT 714.6000 255.6000 715.5000 260.4000 ;
	    RECT 724.2000 259.5000 725.4000 262.2000 ;
	    RECT 738.6000 261.4500 739.8000 261.6000 ;
	    RECT 748.2000 261.4500 749.4000 261.6000 ;
	    RECT 738.6000 260.5500 749.4000 261.4500 ;
	    RECT 738.6000 260.4000 739.8000 260.5500 ;
	    RECT 748.2000 260.4000 749.4000 260.5500 ;
	    RECT 750.3000 260.4000 752.1000 261.6000 ;
	    RECT 754.2000 260.7000 754.5000 262.2000 ;
	    RECT 755.4000 260.4000 756.6000 261.6000 ;
	    RECT 769.8000 261.4500 771.0000 261.6000 ;
	    RECT 757.9500 260.5500 771.0000 261.4500 ;
	    RECT 717.0000 259.2000 718.2000 259.5000 ;
	    RECT 717.0000 258.3000 722.7000 259.2000 ;
	    RECT 721.5000 258.0000 722.7000 258.3000 ;
	    RECT 724.2000 257.4000 725.4000 258.6000 ;
	    RECT 719.1000 257.1000 720.3000 257.4000 ;
	    RECT 719.1000 256.5000 723.3000 257.1000 ;
	    RECT 719.1000 256.2000 725.4000 256.5000 ;
	    RECT 714.6000 254.7000 718.2000 255.6000 ;
	    RECT 713.7000 253.5000 714.9000 253.8000 ;
	    RECT 711.6000 252.6000 714.9000 253.5000 ;
	    RECT 717.3000 253.2000 718.2000 254.7000 ;
	    RECT 717.3000 252.0000 719.4000 253.2000 ;
	    RECT 707.7000 251.1000 708.9000 251.4000 ;
	    RECT 711.9000 251.1000 713.1000 251.4000 ;
	    RECT 702.6000 249.3000 703.8000 250.5000 ;
	    RECT 707.7000 250.2000 713.1000 251.1000 ;
	    RECT 711.0000 249.3000 711.9000 250.2000 ;
	    RECT 717.0000 249.3000 718.2000 250.5000 ;
	    RECT 702.6000 248.4000 705.6000 249.3000 ;
	    RECT 704.4000 243.3000 705.6000 248.4000 ;
	    RECT 708.6000 243.3000 709.8000 249.3000 ;
	    RECT 711.0000 243.3000 712.2000 249.3000 ;
	    RECT 713.4000 243.3000 714.6000 249.3000 ;
	    RECT 717.3000 243.3000 719.1000 249.3000 ;
	    RECT 721.8000 243.3000 723.0000 255.3000 ;
	    RECT 724.2000 243.3000 725.4000 256.2000 ;
	    RECT 748.2000 254.4000 749.4000 255.6000 ;
	    RECT 751.2000 255.3000 752.1000 260.4000 ;
	    RECT 753.0000 259.5000 754.2000 259.8000 ;
	    RECT 753.0000 258.4500 754.2000 258.6000 ;
	    RECT 757.9500 258.4500 758.8500 260.5500 ;
	    RECT 769.8000 260.4000 771.0000 260.5500 ;
	    RECT 781.8000 261.4500 783.0000 261.6000 ;
	    RECT 791.4000 261.4500 792.6000 261.6000 ;
	    RECT 781.8000 260.5500 792.6000 261.4500 ;
	    RECT 781.8000 260.4000 783.0000 260.5500 ;
	    RECT 791.4000 260.4000 792.6000 260.5500 ;
	    RECT 793.8000 259.5000 795.0000 263.7000 ;
	    RECT 815.4000 262.5000 816.6000 262.8000 ;
	    RECT 815.4000 260.4000 816.6000 261.6000 ;
	    RECT 817.8000 259.5000 819.0000 263.7000 ;
	    RECT 839.4000 262.8000 840.6000 269.7000 ;
	    RECT 841.8000 263.7000 843.0000 269.7000 ;
	    RECT 839.4000 261.9000 842.7000 262.8000 ;
	    RECT 844.2000 262.5000 845.4000 269.7000 ;
	    RECT 863.4000 263.7000 864.6000 269.7000 ;
	    RECT 867.3000 264.6000 868.5000 269.7000 ;
	    RECT 870.6000 269.4000 871.8000 270.6000 ;
	    RECT 865.8000 263.7000 868.5000 264.6000 ;
	    RECT 863.4000 262.5000 864.6000 262.8000 ;
	    RECT 839.4000 259.5000 840.6000 259.8000 ;
	    RECT 753.0000 257.5500 758.8500 258.4500 ;
	    RECT 753.0000 257.4000 754.2000 257.5500 ;
	    RECT 751.2000 254.4000 752.7000 255.3000 ;
	    RECT 749.4000 252.6000 750.3000 253.5000 ;
	    RECT 749.4000 251.4000 750.6000 252.6000 ;
	    RECT 749.1000 243.3000 750.3000 249.3000 ;
	    RECT 751.5000 243.3000 752.7000 254.4000 ;
	    RECT 755.4000 243.3000 756.6000 255.3000 ;
	    RECT 769.8000 243.3000 771.0000 259.5000 ;
	    RECT 793.8000 257.4000 795.0000 258.6000 ;
	    RECT 817.8000 258.4500 819.0000 258.6000 ;
	    RECT 837.0000 258.4500 838.2000 258.6000 ;
	    RECT 817.8000 257.5500 838.2000 258.4500 ;
	    RECT 817.8000 257.4000 819.0000 257.5500 ;
	    RECT 837.0000 257.4000 838.2000 257.5500 ;
	    RECT 839.4000 257.4000 840.6000 258.6000 ;
	    RECT 841.8000 257.4000 842.7000 261.9000 ;
	    RECT 844.2000 260.4000 845.4000 261.6000 ;
	    RECT 858.6000 261.4500 859.8000 261.6000 ;
	    RECT 863.4000 261.4500 864.6000 261.6000 ;
	    RECT 858.6000 260.5500 864.6000 261.4500 ;
	    RECT 858.6000 260.4000 859.8000 260.5500 ;
	    RECT 863.4000 260.4000 864.6000 260.5500 ;
	    RECT 865.8000 259.5000 867.0000 263.7000 ;
	    RECT 1002.6000 260.7000 1003.8000 269.7000 ;
	    RECT 1007.4000 263.7000 1008.6000 269.7000 ;
	    RECT 1012.2000 264.9000 1013.4000 269.7000 ;
	    RECT 1014.6000 265.5000 1015.8000 269.7000 ;
	    RECT 1017.0000 265.5000 1018.2000 269.7000 ;
	    RECT 1019.4000 265.5000 1020.6000 269.7000 ;
	    RECT 1021.8000 266.7000 1023.0000 269.7000 ;
	    RECT 1024.2001 265.5000 1025.4000 269.7000 ;
	    RECT 1026.6000 266.7000 1027.8000 269.7000 ;
	    RECT 1029.0000 265.5000 1030.2001 269.7000 ;
	    RECT 1031.4000 265.5000 1032.6000 269.7000 ;
	    RECT 1033.8000 265.5000 1035.0000 269.7000 ;
	    RECT 1036.2001 265.5000 1037.4000 269.7000 ;
	    RECT 1009.5000 263.7000 1013.4000 264.9000 ;
	    RECT 1038.6000 264.9000 1039.8000 269.7000 ;
	    RECT 1018.5000 263.7000 1025.4000 264.6000 ;
	    RECT 1009.5000 262.8000 1010.7000 263.7000 ;
	    RECT 1006.2000 261.6000 1010.7000 262.8000 ;
	    RECT 1002.6000 259.5000 1015.8000 260.7000 ;
	    RECT 1018.5000 260.1000 1019.7000 263.7000 ;
	    RECT 1024.2001 263.4000 1025.4000 263.7000 ;
	    RECT 1026.6000 263.4000 1027.8000 264.6000 ;
	    RECT 1028.7001 263.4000 1029.0000 264.6000 ;
	    RECT 1033.5000 263.4000 1035.0000 264.6000 ;
	    RECT 1038.6000 263.7000 1042.2001 264.9000 ;
	    RECT 1043.4000 263.7000 1044.6000 269.7000 ;
	    RECT 1021.8000 262.5000 1023.0000 262.8000 ;
	    RECT 1024.2001 262.2000 1025.4000 262.5000 ;
	    RECT 1021.8000 260.4000 1023.0000 261.6000 ;
	    RECT 1024.2001 261.3000 1030.8000 262.2000 ;
	    RECT 1029.6000 261.0000 1030.8000 261.3000 ;
	    RECT 844.2000 258.6000 845.4000 259.5000 ;
	    RECT 772.2000 243.3000 773.4000 249.3000 ;
	    RECT 791.4000 243.3000 792.6000 249.3000 ;
	    RECT 793.8000 243.3000 795.0000 256.5000 ;
	    RECT 796.2000 254.4000 797.4000 255.6000 ;
	    RECT 796.2000 253.2000 797.4000 253.5000 ;
	    RECT 796.2000 243.3000 797.4000 249.3000 ;
	    RECT 815.4000 243.3000 816.6000 249.3000 ;
	    RECT 817.8000 243.3000 819.0000 256.5000 ;
	    RECT 841.8000 256.2000 843.6000 257.4000 ;
	    RECT 820.2000 254.4000 821.4000 255.6000 ;
	    RECT 841.8000 255.3000 842.7000 256.2000 ;
	    RECT 844.5000 255.3000 845.4000 258.6000 ;
	    RECT 865.8000 258.4500 867.0000 258.6000 ;
	    RECT 875.4000 258.4500 876.6000 258.6000 ;
	    RECT 865.8000 257.5500 876.6000 258.4500 ;
	    RECT 865.8000 257.4000 867.0000 257.5500 ;
	    RECT 875.4000 257.4000 876.6000 257.5500 ;
	    RECT 839.4000 254.4000 842.7000 255.3000 ;
	    RECT 820.2000 253.2000 821.4000 253.5000 ;
	    RECT 820.2000 243.3000 821.4000 249.3000 ;
	    RECT 839.4000 243.3000 840.6000 254.4000 ;
	    RECT 841.8000 243.3000 843.0000 253.5000 ;
	    RECT 844.2000 243.3000 845.4000 255.3000 ;
	    RECT 863.4000 243.3000 864.6000 249.3000 ;
	    RECT 865.8000 243.3000 867.0000 256.5000 ;
	    RECT 868.2000 255.4500 869.4000 255.6000 ;
	    RECT 870.6000 255.4500 871.8000 255.6000 ;
	    RECT 868.2000 254.5500 871.8000 255.4500 ;
	    RECT 868.2000 254.4000 869.4000 254.5500 ;
	    RECT 870.6000 254.4000 871.8000 254.5500 ;
	    RECT 868.2000 253.2000 869.4000 253.5000 ;
	    RECT 1002.6000 251.1000 1003.8000 259.5000 ;
	    RECT 1016.7000 258.9000 1019.7000 260.1000 ;
	    RECT 1025.4000 258.9000 1030.2001 260.1000 ;
	    RECT 1033.8000 259.2000 1035.0000 263.4000 ;
	    RECT 1041.0000 262.8000 1042.2001 263.7000 ;
	    RECT 1041.0000 261.9000 1043.7001 262.8000 ;
	    RECT 1042.5000 260.1000 1043.7001 261.9000 ;
	    RECT 1048.2001 261.9000 1049.4000 269.7000 ;
	    RECT 1050.6000 264.0000 1051.8000 269.7000 ;
	    RECT 1053.0000 266.7000 1054.2001 269.7000 ;
	    RECT 1072.2001 266.7000 1073.4000 269.7000 ;
	    RECT 1074.6000 266.7000 1075.8000 269.7000 ;
	    RECT 1077.0000 266.7000 1078.2001 269.7000 ;
	    RECT 1050.6000 262.8000 1052.1000 264.0000 ;
	    RECT 1048.2001 261.0000 1050.0000 261.9000 ;
	    RECT 1042.5000 258.9000 1048.2001 260.1000 ;
	    RECT 1004.7000 258.0000 1005.9000 258.3000 ;
	    RECT 1004.7000 257.1000 1011.3000 258.0000 ;
	    RECT 1012.2000 257.4000 1013.4000 258.6000 ;
	    RECT 1038.6000 258.0000 1039.8000 258.9000 ;
	    RECT 1049.1000 258.0000 1050.0000 261.0000 ;
	    RECT 1014.3000 257.1000 1039.8000 258.0000 ;
	    RECT 1048.8000 257.1000 1050.0000 258.0000 ;
	    RECT 1046.7001 256.2000 1047.9000 256.5000 ;
	    RECT 1007.4000 254.4000 1008.6000 255.6000 ;
	    RECT 1009.5000 255.3000 1047.9000 256.2000 ;
	    RECT 1012.5000 255.0000 1013.7000 255.3000 ;
	    RECT 1048.8000 254.4000 1049.7001 257.1000 ;
	    RECT 1050.9000 256.2000 1052.1000 262.8000 ;
	    RECT 1074.6000 262.5000 1075.5000 266.7000 ;
	    RECT 1077.0000 265.5000 1078.2001 265.8000 ;
	    RECT 1104.3000 265.2000 1105.5000 269.7000 ;
	    RECT 1077.0000 264.4500 1078.2001 264.6000 ;
	    RECT 1084.2001 264.4500 1085.4000 264.6000 ;
	    RECT 1077.0000 263.5500 1085.4000 264.4500 ;
	    RECT 1077.0000 263.4000 1078.2001 263.5500 ;
	    RECT 1084.2001 263.4000 1085.4000 263.5500 ;
	    RECT 1103.4000 263.7000 1105.5000 265.2000 ;
	    RECT 1106.7001 264.0000 1107.9000 269.7000 ;
	    RECT 1110.6000 263.7000 1111.8000 269.7000 ;
	    RECT 1141.8000 264.0000 1143.0000 269.7000 ;
	    RECT 1144.2001 264.9000 1145.4000 269.7000 ;
	    RECT 1146.6000 264.0000 1147.8000 269.7000 ;
	    RECT 1141.8000 263.7000 1147.8000 264.0000 ;
	    RECT 1149.0000 263.7000 1150.2001 269.7000 ;
	    RECT 1173.0000 266.7000 1174.2001 269.7000 ;
	    RECT 1173.3000 265.5000 1174.5000 265.8000 ;
	    RECT 1158.6000 264.4500 1159.8000 264.6000 ;
	    RECT 1173.0000 264.4500 1174.2001 264.6000 ;
	    RECT 1053.0000 261.4500 1054.2001 261.6000 ;
	    RECT 1074.6000 261.4500 1075.8000 261.6000 ;
	    RECT 1053.0000 260.5500 1075.8000 261.4500 ;
	    RECT 1053.0000 260.4000 1054.2001 260.5500 ;
	    RECT 1074.6000 260.4000 1075.8000 260.5500 ;
	    RECT 1103.4000 259.5000 1104.3000 263.7000 ;
	    RECT 1110.6000 263.4000 1111.5000 263.7000 ;
	    RECT 1108.8000 262.8000 1111.5000 263.4000 ;
	    RECT 1142.1000 263.1000 1147.5000 263.7000 ;
	    RECT 1105.2001 262.5000 1111.5000 262.8000 ;
	    RECT 1149.0000 262.5000 1149.9000 263.7000 ;
	    RECT 1158.6000 263.5500 1174.2001 264.4500 ;
	    RECT 1175.4000 263.7000 1176.6000 269.7000 ;
	    RECT 1179.3000 263.7000 1180.5000 269.7000 ;
	    RECT 1158.6000 263.4000 1159.8000 263.5500 ;
	    RECT 1173.0000 263.4000 1174.2001 263.5500 ;
	    RECT 1105.2001 261.9000 1109.7001 262.5000 ;
	    RECT 1105.2001 261.6000 1106.4000 261.9000 ;
	    RECT 1072.2001 257.4000 1073.4000 258.6000 ;
	    RECT 1072.2001 256.2000 1073.4000 256.5000 ;
	    RECT 1017.0000 254.1000 1018.2000 254.4000 ;
	    RECT 1010.1000 253.5000 1018.2000 254.1000 ;
	    RECT 1008.9000 253.2000 1018.2000 253.5000 ;
	    RECT 1019.7000 253.5000 1032.6000 254.4000 ;
	    RECT 1005.0000 252.0000 1007.4000 253.2000 ;
	    RECT 1008.9000 252.3000 1011.0000 253.2000 ;
	    RECT 1019.7000 252.3000 1020.6000 253.5000 ;
	    RECT 1031.4000 253.2000 1032.6000 253.5000 ;
	    RECT 1036.2001 253.5000 1049.7001 254.4000 ;
	    RECT 1050.6000 255.0000 1052.1000 256.2000 ;
	    RECT 1074.6000 255.3000 1075.5000 259.5000 ;
	    RECT 1103.4000 257.4000 1104.6000 258.6000 ;
	    RECT 1105.5000 256.5000 1106.4000 261.6000 ;
	    RECT 1107.6000 260.7000 1108.8000 261.0000 ;
	    RECT 1107.6000 259.8000 1109.1000 260.7000 ;
	    RECT 1110.6000 260.4000 1111.8000 261.6000 ;
	    RECT 1120.2001 261.4500 1121.4000 261.6000 ;
	    RECT 1141.8000 261.4500 1143.0000 261.6000 ;
	    RECT 1120.2001 260.5500 1143.0000 261.4500 ;
	    RECT 1143.9000 260.7000 1144.2001 262.2000 ;
	    RECT 1120.2001 260.4000 1121.4000 260.5500 ;
	    RECT 1141.8000 260.4000 1143.0000 260.5500 ;
	    RECT 1146.3000 260.4000 1148.1000 261.6000 ;
	    RECT 1149.0000 261.4500 1150.2001 261.6000 ;
	    RECT 1151.4000 261.4500 1152.6000 261.6000 ;
	    RECT 1149.0000 260.5500 1152.6000 261.4500 ;
	    RECT 1149.0000 260.4000 1150.2001 260.5500 ;
	    RECT 1151.4000 260.4000 1152.6000 260.5500 ;
	    RECT 1108.2001 259.5000 1109.1000 259.8000 ;
	    RECT 1144.2001 259.5000 1145.4000 259.8000 ;
	    RECT 1110.6000 259.2000 1111.8000 259.5000 ;
	    RECT 1108.2001 257.4000 1109.4000 258.6000 ;
	    RECT 1144.2001 258.4500 1145.4000 258.6000 ;
	    RECT 1139.5500 257.5500 1145.4000 258.4500 ;
	    RECT 1103.4000 255.3000 1104.3000 256.5000 ;
	    RECT 1105.5000 255.6000 1109.1000 256.5000 ;
	    RECT 1050.6000 253.5000 1051.8000 255.0000 ;
	    RECT 1073.1000 254.1000 1075.8000 255.3000 ;
	    RECT 1036.2001 253.2000 1037.4000 253.5000 ;
	    RECT 1006.5000 251.4000 1007.4000 252.0000 ;
	    RECT 1011.9000 251.4000 1020.6000 252.3000 ;
	    RECT 1021.5000 251.4000 1025.4000 252.6000 ;
	    RECT 1002.6000 250.2000 1005.6000 251.1000 ;
	    RECT 1006.5000 250.2000 1012.8000 251.4000 ;
	    RECT 969.0000 249.4500 970.2000 249.6000 ;
	    RECT 988.2000 249.4500 989.4000 249.6000 ;
	    RECT 868.2000 243.3000 869.4000 249.3000 ;
	    RECT 969.0000 248.5500 989.4000 249.4500 ;
	    RECT 1004.7000 249.3000 1005.6000 250.2000 ;
	    RECT 969.0000 248.4000 970.2000 248.5500 ;
	    RECT 988.2000 248.4000 989.4000 248.5500 ;
	    RECT 957.0000 246.4500 958.2000 246.6000 ;
	    RECT 988.2000 246.4500 989.4000 246.6000 ;
	    RECT 957.0000 245.5500 989.4000 246.4500 ;
	    RECT 957.0000 245.4000 958.2000 245.5500 ;
	    RECT 988.2000 245.4000 989.4000 245.5500 ;
	    RECT 1002.6000 243.3000 1003.8000 249.3000 ;
	    RECT 1004.7000 248.4000 1006.2000 249.3000 ;
	    RECT 1005.0000 243.3000 1006.2000 248.4000 ;
	    RECT 1007.4000 242.4000 1008.6000 249.3000 ;
	    RECT 1009.8000 243.3000 1011.0000 250.2000 ;
	    RECT 1012.2000 243.3000 1013.4000 249.3000 ;
	    RECT 1014.6000 243.3000 1015.8000 247.5000 ;
	    RECT 1017.0000 243.3000 1018.2000 247.5000 ;
	    RECT 1019.4000 243.3000 1020.6000 250.5000 ;
	    RECT 1021.8000 243.3000 1023.0000 249.3000 ;
	    RECT 1024.2001 243.3000 1025.4000 250.5000 ;
	    RECT 1026.6000 243.3000 1027.8000 249.3000 ;
	    RECT 1029.0000 243.3000 1030.2001 252.6000 ;
	    RECT 1041.0000 251.4000 1044.9000 252.6000 ;
	    RECT 1033.8000 250.2000 1040.1000 251.4000 ;
	    RECT 1031.4000 243.3000 1032.6000 247.5000 ;
	    RECT 1033.8000 243.3000 1035.0000 247.5000 ;
	    RECT 1036.2001 243.3000 1037.4000 247.5000 ;
	    RECT 1038.6000 243.3000 1039.8000 249.3000 ;
	    RECT 1041.0000 243.3000 1042.2001 251.4000 ;
	    RECT 1048.8000 251.1000 1049.7001 253.5000 ;
	    RECT 1050.6000 251.4000 1051.8000 252.6000 ;
	    RECT 1045.8000 250.2000 1049.7001 251.1000 ;
	    RECT 1043.4000 243.3000 1044.6000 249.3000 ;
	    RECT 1045.8000 243.3000 1047.0000 250.2000 ;
	    RECT 1048.2001 243.3000 1049.4000 249.3000 ;
	    RECT 1050.6000 243.3000 1051.8000 250.5000 ;
	    RECT 1053.0000 243.3000 1054.2001 249.3000 ;
	    RECT 1073.1000 243.3000 1074.3000 254.1000 ;
	    RECT 1077.0000 243.3000 1078.2001 255.3000 ;
	    RECT 1103.4000 243.3000 1104.6000 255.3000 ;
	    RECT 1105.8000 243.3000 1107.0000 254.7000 ;
	    RECT 1108.2001 249.3000 1109.1000 255.6000 ;
	    RECT 1110.6000 255.4500 1111.8000 255.6000 ;
	    RECT 1139.5500 255.4500 1140.4501 257.5500 ;
	    RECT 1144.2001 257.4000 1145.4000 257.5500 ;
	    RECT 1110.6000 254.5500 1140.4501 255.4500 ;
	    RECT 1146.3000 255.3000 1147.2001 260.4000 ;
	    RECT 1158.6000 258.4500 1159.8000 258.6000 ;
	    RECT 1173.0000 258.4500 1174.2001 258.6000 ;
	    RECT 1158.6000 257.5500 1174.2001 258.4500 ;
	    RECT 1175.7001 258.3000 1176.6000 263.7000 ;
	    RECT 1177.8000 260.4000 1179.0000 261.6000 ;
	    RECT 1206.0000 261.3000 1207.2001 269.7000 ;
	    RECT 1204.5000 260.7000 1207.2001 261.3000 ;
	    RECT 1211.4000 260.7000 1212.6000 269.7000 ;
	    RECT 1235.4000 264.0000 1236.6000 269.7000 ;
	    RECT 1237.8000 264.9000 1239.0000 269.7000 ;
	    RECT 1240.2001 264.0000 1241.4000 269.7000 ;
	    RECT 1235.4000 263.7000 1241.4000 264.0000 ;
	    RECT 1242.6000 263.7000 1243.8000 269.7000 ;
	    RECT 1267.5000 263.7000 1268.7001 269.7000 ;
	    RECT 1271.4000 263.7000 1272.6000 269.7000 ;
	    RECT 1273.8000 266.7000 1275.0000 269.7000 ;
	    RECT 1273.5000 265.5000 1274.7001 265.8000 ;
	    RECT 1273.8000 264.4500 1275.0000 264.6000 ;
	    RECT 1276.2001 264.4500 1277.4000 264.6000 ;
	    RECT 1235.7001 263.1000 1241.1000 263.7000 ;
	    RECT 1242.6000 262.5000 1243.5000 263.7000 ;
	    RECT 1204.5000 260.4000 1206.9000 260.7000 ;
	    RECT 1235.4000 260.4000 1236.6000 261.6000 ;
	    RECT 1237.5000 260.7000 1237.8000 262.2000 ;
	    RECT 1239.9000 260.4000 1241.7001 261.6000 ;
	    RECT 1242.6000 261.4500 1243.8000 261.6000 ;
	    RECT 1266.6000 261.4500 1267.8000 261.6000 ;
	    RECT 1242.6000 260.5500 1267.8000 261.4500 ;
	    RECT 1242.6000 260.4000 1243.8000 260.5500 ;
	    RECT 1266.6000 260.4000 1267.8000 260.5500 ;
	    RECT 1269.0000 260.4000 1270.2001 261.6000 ;
	    RECT 1177.8000 259.2000 1179.0000 259.5000 ;
	    RECT 1158.6000 257.4000 1159.8000 257.5500 ;
	    RECT 1173.0000 257.4000 1174.2001 257.5500 ;
	    RECT 1175.1000 257.4000 1176.6000 258.3000 ;
	    RECT 1179.0000 256.8000 1179.3000 258.3000 ;
	    RECT 1180.2001 257.4000 1181.4000 258.6000 ;
	    RECT 1204.5000 256.5000 1205.4000 260.4000 ;
	    RECT 1237.8000 259.5000 1239.0000 259.8000 ;
	    RECT 1207.8000 257.4000 1208.1000 258.6000 ;
	    RECT 1209.0000 257.4000 1210.2001 258.6000 ;
	    RECT 1237.8000 257.4000 1239.0000 258.6000 ;
	    RECT 1211.4000 256.5000 1212.6000 256.8000 ;
	    RECT 1110.6000 254.4000 1111.8000 254.5500 ;
	    RECT 1108.2001 243.3000 1109.4000 249.3000 ;
	    RECT 1110.6000 243.3000 1111.8000 249.3000 ;
	    RECT 1141.8000 243.3000 1143.0000 255.3000 ;
	    RECT 1145.7001 254.4000 1147.2001 255.3000 ;
	    RECT 1149.0000 254.4000 1150.2001 255.6000 ;
	    RECT 1173.3000 255.3000 1174.2001 256.5000 ;
	    RECT 1145.7001 243.3000 1146.9000 254.4000 ;
	    RECT 1148.1000 252.6000 1149.0000 253.5000 ;
	    RECT 1147.8000 251.4000 1149.0000 252.6000 ;
	    RECT 1148.1000 243.3000 1149.3000 249.3000 ;
	    RECT 1173.0000 243.3000 1174.2001 255.3000 ;
	    RECT 1175.4000 254.4000 1181.4000 255.3000 ;
	    RECT 1204.2001 254.4000 1205.4000 255.6000 ;
	    RECT 1211.4000 254.4000 1212.6000 255.6000 ;
	    RECT 1239.9000 255.3000 1240.8000 260.4000 ;
	    RECT 1269.0000 259.2000 1270.2001 259.5000 ;
	    RECT 1247.4000 258.4500 1248.6000 258.6000 ;
	    RECT 1266.6000 258.4500 1267.8000 258.6000 ;
	    RECT 1247.4000 257.5500 1267.8000 258.4500 ;
	    RECT 1271.4000 258.3000 1272.3000 263.7000 ;
	    RECT 1273.8000 263.5500 1277.4000 264.4500 ;
	    RECT 1273.8000 263.4000 1275.0000 263.5500 ;
	    RECT 1276.2001 263.4000 1277.4000 263.5500 ;
	    RECT 1297.8000 260.7000 1299.0000 269.7000 ;
	    RECT 1303.2001 261.3000 1304.4000 269.7000 ;
	    RECT 1325.1000 264.6000 1326.3000 269.7000 ;
	    RECT 1325.1000 263.7000 1327.8000 264.6000 ;
	    RECT 1329.0000 263.7000 1330.2001 269.7000 ;
	    RECT 1360.2001 263.7000 1361.4000 269.7000 ;
	    RECT 1362.6000 264.0000 1363.8000 269.7000 ;
	    RECT 1365.0000 264.9000 1366.2001 269.7000 ;
	    RECT 1367.4000 264.0000 1368.6000 269.7000 ;
	    RECT 1391.4000 266.7000 1392.6000 269.7000 ;
	    RECT 1391.7001 265.5000 1392.9000 265.8000 ;
	    RECT 1362.6000 263.7000 1368.6000 264.0000 ;
	    RECT 1389.0000 264.4500 1390.2001 264.6000 ;
	    RECT 1391.4000 264.4500 1392.6000 264.6000 ;
	    RECT 1303.2001 260.7000 1305.9000 261.3000 ;
	    RECT 1303.5000 260.4000 1305.9000 260.7000 ;
	    RECT 1247.4000 257.4000 1248.6000 257.5500 ;
	    RECT 1266.6000 257.4000 1267.8000 257.5500 ;
	    RECT 1268.7001 256.8000 1269.0000 258.3000 ;
	    RECT 1271.4000 257.4000 1272.9000 258.3000 ;
	    RECT 1273.8000 257.4000 1275.0000 258.6000 ;
	    RECT 1300.2001 257.4000 1301.4000 258.6000 ;
	    RECT 1302.3000 257.4000 1302.6000 258.6000 ;
	    RECT 1297.8000 256.5000 1299.0000 256.8000 ;
	    RECT 1305.0000 256.5000 1305.9000 260.4000 ;
	    RECT 1326.6000 259.5000 1327.8000 263.7000 ;
	    RECT 1329.0000 262.5000 1330.2001 262.8000 ;
	    RECT 1360.5000 262.5000 1361.4000 263.7000 ;
	    RECT 1362.9000 263.1000 1368.3000 263.7000 ;
	    RECT 1389.0000 263.5500 1392.6000 264.4500 ;
	    RECT 1393.8000 263.7000 1395.0000 269.7000 ;
	    RECT 1397.7001 263.7000 1398.9000 269.7000 ;
	    RECT 1427.4000 263.7000 1428.6000 269.7000 ;
	    RECT 1431.3000 263.7000 1433.7001 269.7000 ;
	    RECT 1436.4000 263.7000 1437.6000 269.7000 ;
	    RECT 1456.2001 263.7000 1457.4000 269.7000 ;
	    RECT 1460.1000 264.6000 1461.3000 269.7000 ;
	    RECT 1473.0000 267.4500 1474.2001 267.6000 ;
	    RECT 1480.2001 267.4500 1481.4000 267.6000 ;
	    RECT 1473.0000 266.5500 1481.4000 267.4500 ;
	    RECT 1473.0000 266.4000 1474.2001 266.5500 ;
	    RECT 1480.2001 266.4000 1481.4000 266.5500 ;
	    RECT 1458.6000 263.7000 1461.3000 264.6000 ;
	    RECT 1389.0000 263.4000 1390.2001 263.5500 ;
	    RECT 1391.4000 263.4000 1392.6000 263.5500 ;
	    RECT 1329.0000 260.4000 1330.2001 261.6000 ;
	    RECT 1333.8000 261.4500 1335.0000 261.6000 ;
	    RECT 1360.2001 261.4500 1361.4000 261.6000 ;
	    RECT 1333.8000 260.5500 1361.4000 261.4500 ;
	    RECT 1333.8000 260.4000 1335.0000 260.5500 ;
	    RECT 1360.2001 260.4000 1361.4000 260.5500 ;
	    RECT 1362.3000 260.4000 1364.1000 261.6000 ;
	    RECT 1366.2001 260.7000 1366.5000 262.2000 ;
	    RECT 1367.4000 261.4500 1368.6000 261.6000 ;
	    RECT 1369.8000 261.4500 1371.0000 261.6000 ;
	    RECT 1367.4000 260.5500 1371.0000 261.4500 ;
	    RECT 1367.4000 260.4000 1368.6000 260.5500 ;
	    RECT 1369.8000 260.4000 1371.0000 260.5500 ;
	    RECT 1309.8000 258.4500 1311.0000 258.6000 ;
	    RECT 1326.6000 258.4500 1327.8000 258.6000 ;
	    RECT 1309.8000 257.5500 1327.8000 258.4500 ;
	    RECT 1309.8000 257.4000 1311.0000 257.5500 ;
	    RECT 1326.6000 257.4000 1327.8000 257.5500 ;
	    RECT 1175.4000 243.3000 1176.6000 254.4000 ;
	    RECT 1177.8000 243.3000 1179.0000 253.5000 ;
	    RECT 1180.2001 243.3000 1181.4000 254.4000 ;
	    RECT 1206.6000 253.5000 1207.8000 253.8000 ;
	    RECT 1204.5000 250.5000 1205.4000 253.5000 ;
	    RECT 1206.6000 251.4000 1207.8000 252.6000 ;
	    RECT 1204.5000 249.6000 1209.9000 250.5000 ;
	    RECT 1204.5000 249.3000 1205.4000 249.6000 ;
	    RECT 1204.2001 243.3000 1205.4000 249.3000 ;
	    RECT 1209.0000 249.3000 1209.9000 249.6000 ;
	    RECT 1206.6000 243.3000 1207.8000 248.7000 ;
	    RECT 1209.0000 243.3000 1210.2001 249.3000 ;
	    RECT 1211.4000 243.3000 1212.6000 249.3000 ;
	    RECT 1235.4000 243.3000 1236.6000 255.3000 ;
	    RECT 1239.3000 254.4000 1240.8000 255.3000 ;
	    RECT 1242.6000 254.4000 1243.8000 255.6000 ;
	    RECT 1273.8000 255.3000 1274.7001 256.5000 ;
	    RECT 1276.2001 255.4500 1277.4000 255.6000 ;
	    RECT 1297.8000 255.4500 1299.0000 255.6000 ;
	    RECT 1266.6000 254.4000 1272.6000 255.3000 ;
	    RECT 1239.3000 243.3000 1240.5000 254.4000 ;
	    RECT 1241.7001 252.6000 1242.6000 253.5000 ;
	    RECT 1241.4000 251.4000 1242.6000 252.6000 ;
	    RECT 1241.7001 243.3000 1242.9000 249.3000 ;
	    RECT 1266.6000 243.3000 1267.8000 254.4000 ;
	    RECT 1269.0000 243.3000 1270.2001 253.5000 ;
	    RECT 1271.4000 243.3000 1272.6000 254.4000 ;
	    RECT 1273.8000 243.3000 1275.0000 255.3000 ;
	    RECT 1276.2001 254.5500 1299.0000 255.4500 ;
	    RECT 1276.2001 254.4000 1277.4000 254.5500 ;
	    RECT 1297.8000 254.4000 1299.0000 254.5500 ;
	    RECT 1305.0000 255.4500 1306.2001 255.6000 ;
	    RECT 1321.8000 255.4500 1323.0000 255.6000 ;
	    RECT 1305.0000 254.5500 1323.0000 255.4500 ;
	    RECT 1305.0000 254.4000 1306.2001 254.5500 ;
	    RECT 1321.8000 254.4000 1323.0000 254.5500 ;
	    RECT 1324.2001 254.4000 1325.4000 255.6000 ;
	    RECT 1302.6000 253.5000 1303.8000 253.8000 ;
	    RECT 1293.0000 252.4500 1294.2001 252.6000 ;
	    RECT 1302.6000 252.4500 1303.8000 252.6000 ;
	    RECT 1293.0000 251.5500 1303.8000 252.4500 ;
	    RECT 1293.0000 251.4000 1294.2001 251.5500 ;
	    RECT 1302.6000 251.4000 1303.8000 251.5500 ;
	    RECT 1305.0000 250.5000 1305.9000 253.5000 ;
	    RECT 1324.2001 253.2000 1325.4000 253.5000 ;
	    RECT 1300.5000 249.6000 1305.9000 250.5000 ;
	    RECT 1300.5000 249.3000 1301.4000 249.6000 ;
	    RECT 1297.8000 243.3000 1299.0000 249.3000 ;
	    RECT 1300.2001 243.3000 1301.4000 249.3000 ;
	    RECT 1305.0000 249.3000 1305.9000 249.6000 ;
	    RECT 1302.6000 243.3000 1303.8000 248.7000 ;
	    RECT 1305.0000 243.3000 1306.2001 249.3000 ;
	    RECT 1324.2001 243.3000 1325.4000 249.3000 ;
	    RECT 1326.6000 243.3000 1327.8000 256.5000 ;
	    RECT 1331.4000 255.4500 1332.6000 255.6000 ;
	    RECT 1360.2001 255.4500 1361.4000 255.6000 ;
	    RECT 1331.4000 254.5500 1361.4000 255.4500 ;
	    RECT 1331.4000 254.4000 1332.6000 254.5500 ;
	    RECT 1360.2001 254.4000 1361.4000 254.5500 ;
	    RECT 1363.2001 255.3000 1364.1000 260.4000 ;
	    RECT 1365.0000 259.5000 1366.2001 259.8000 ;
	    RECT 1365.0000 257.4000 1366.2001 258.6000 ;
	    RECT 1391.4000 257.4000 1392.6000 258.6000 ;
	    RECT 1394.1000 258.3000 1395.0000 263.7000 ;
	    RECT 1396.2001 261.4500 1397.4000 261.6000 ;
	    RECT 1403.4000 261.4500 1404.6000 261.6000 ;
	    RECT 1429.8000 261.4500 1431.0000 261.6000 ;
	    RECT 1396.2001 260.5500 1431.0000 261.4500 ;
	    RECT 1396.2001 260.4000 1397.4000 260.5500 ;
	    RECT 1403.4000 260.4000 1404.6000 260.5500 ;
	    RECT 1429.8000 260.4000 1431.0000 260.5500 ;
	    RECT 1432.2001 259.5000 1433.1000 263.7000 ;
	    RECT 1456.2001 262.5000 1457.4000 262.8000 ;
	    RECT 1434.6000 260.4000 1435.8000 261.6000 ;
	    RECT 1456.2001 261.4500 1457.4000 261.6000 ;
	    RECT 1437.1500 260.5500 1457.4000 261.4500 ;
	    RECT 1396.2001 259.2000 1397.4000 259.5000 ;
	    RECT 1430.1000 258.6000 1431.3000 259.5000 ;
	    RECT 1434.6000 259.2000 1435.8000 259.5000 ;
	    RECT 1437.1500 258.6000 1438.0500 260.5500 ;
	    RECT 1456.2001 260.4000 1457.4000 260.5500 ;
	    RECT 1458.6000 259.5000 1459.8000 263.7000 ;
	    RECT 1485.0000 260.7000 1486.2001 269.7000 ;
	    RECT 1490.4000 261.3000 1491.6000 269.7000 ;
	    RECT 1520.4000 261.3000 1521.6000 269.7000 ;
	    RECT 1490.4000 260.7000 1493.1000 261.3000 ;
	    RECT 1490.7001 260.4000 1493.1000 260.7000 ;
	    RECT 1393.5000 257.4000 1395.0000 258.3000 ;
	    RECT 1397.4000 256.8000 1397.7001 258.3000 ;
	    RECT 1398.6000 257.4000 1399.8000 258.6000 ;
	    RECT 1405.8000 258.4500 1407.0000 258.6000 ;
	    RECT 1427.4000 258.4500 1428.6000 258.6000 ;
	    RECT 1405.8000 257.5500 1428.6000 258.4500 ;
	    RECT 1405.8000 257.4000 1407.0000 257.5500 ;
	    RECT 1427.4000 257.4000 1428.6000 257.5500 ;
	    RECT 1432.2001 257.4000 1433.4000 258.6000 ;
	    RECT 1430.1000 256.5000 1431.3000 257.1000 ;
	    RECT 1435.8000 256.8000 1436.1000 258.3000 ;
	    RECT 1437.0000 257.4000 1438.2001 258.6000 ;
	    RECT 1441.8000 258.4500 1443.0000 258.6000 ;
	    RECT 1458.6000 258.4500 1459.8000 258.6000 ;
	    RECT 1441.8000 257.5500 1459.8000 258.4500 ;
	    RECT 1441.8000 257.4000 1443.0000 257.5500 ;
	    RECT 1458.6000 257.4000 1459.8000 257.5500 ;
	    RECT 1487.4000 257.4000 1488.6000 258.6000 ;
	    RECT 1489.5000 257.4000 1489.8000 258.6000 ;
	    RECT 1485.0000 256.5000 1486.2001 256.8000 ;
	    RECT 1492.2001 256.5000 1493.1000 260.4000 ;
	    RECT 1518.9000 260.7000 1521.6000 261.3000 ;
	    RECT 1525.8000 260.7000 1527.0000 269.7000 ;
	    RECT 1549.8000 260.7000 1551.0000 269.7000 ;
	    RECT 1555.2001 261.3000 1556.4000 269.7000 ;
	    RECT 1555.2001 260.7000 1557.9000 261.3000 ;
	    RECT 1518.9000 260.4000 1521.3000 260.7000 ;
	    RECT 1555.5000 260.4000 1557.9000 260.7000 ;
	    RECT 1518.9000 256.5000 1519.8000 260.4000 ;
	    RECT 1522.2001 257.4000 1522.5000 258.6000 ;
	    RECT 1523.4000 257.4000 1524.6000 258.6000 ;
	    RECT 1552.2001 257.4000 1553.4000 258.6000 ;
	    RECT 1554.3000 257.4000 1554.6000 258.6000 ;
	    RECT 1525.8000 256.5000 1527.0000 256.8000 ;
	    RECT 1549.8000 256.5000 1551.0000 256.8000 ;
	    RECT 1557.0000 256.5000 1557.9000 260.4000 ;
	    RECT 1391.7001 255.3000 1392.6000 256.5000 ;
	    RECT 1427.4000 256.2000 1428.6000 256.5000 ;
	    RECT 1430.1000 256.2000 1433.1000 256.5000 ;
	    RECT 1430.1000 255.3000 1431.0000 256.2000 ;
	    RECT 1363.2001 254.4000 1364.7001 255.3000 ;
	    RECT 1361.4000 252.6000 1362.3000 253.5000 ;
	    RECT 1361.4000 251.4000 1362.6000 252.6000 ;
	    RECT 1329.0000 243.3000 1330.2001 249.3000 ;
	    RECT 1361.1000 243.3000 1362.3000 249.3000 ;
	    RECT 1363.5000 243.3000 1364.7001 254.4000 ;
	    RECT 1367.4000 243.3000 1368.6000 255.3000 ;
	    RECT 1391.4000 243.3000 1392.6000 255.3000 ;
	    RECT 1393.8000 254.4000 1399.8000 255.3000 ;
	    RECT 1393.8000 243.3000 1395.0000 254.4000 ;
	    RECT 1396.2001 243.3000 1397.4000 253.5000 ;
	    RECT 1398.6000 243.3000 1399.8000 254.4000 ;
	    RECT 1427.4000 244.2000 1428.6000 255.3000 ;
	    RECT 1429.8000 245.1000 1431.0000 255.3000 ;
	    RECT 1432.2001 254.4000 1438.2001 255.3000 ;
	    RECT 1432.2001 244.2000 1433.4000 254.4000 ;
	    RECT 1427.4000 243.3000 1433.4000 244.2000 ;
	    RECT 1434.6000 243.3000 1435.8000 253.5000 ;
	    RECT 1437.0000 243.3000 1438.2001 254.4000 ;
	    RECT 1456.2001 243.3000 1457.4000 249.3000 ;
	    RECT 1458.6000 243.3000 1459.8000 256.5000 ;
	    RECT 1461.0000 254.4000 1462.2001 255.6000 ;
	    RECT 1470.6000 255.4500 1471.8000 255.6000 ;
	    RECT 1485.0000 255.4500 1486.2001 255.6000 ;
	    RECT 1470.6000 254.5500 1486.2001 255.4500 ;
	    RECT 1470.6000 254.4000 1471.8000 254.5500 ;
	    RECT 1485.0000 254.4000 1486.2001 254.5500 ;
	    RECT 1492.2001 254.4000 1493.4000 255.6000 ;
	    RECT 1497.0000 255.4500 1498.2001 255.6000 ;
	    RECT 1518.6000 255.4500 1519.8000 255.6000 ;
	    RECT 1497.0000 254.5500 1519.8000 255.4500 ;
	    RECT 1497.0000 254.4000 1498.2001 254.5500 ;
	    RECT 1518.6000 254.4000 1519.8000 254.5500 ;
	    RECT 1525.8000 255.4500 1527.0000 255.6000 ;
	    RECT 1545.0000 255.4500 1546.2001 255.6000 ;
	    RECT 1525.8000 254.5500 1546.2001 255.4500 ;
	    RECT 1525.8000 254.4000 1527.0000 254.5500 ;
	    RECT 1545.0000 254.4000 1546.2001 254.5500 ;
	    RECT 1549.8000 254.4000 1551.0000 255.6000 ;
	    RECT 1557.0000 254.4000 1558.2001 255.6000 ;
	    RECT 1489.8000 253.5000 1491.0000 253.8000 ;
	    RECT 1521.0000 253.5000 1522.2001 253.8000 ;
	    RECT 1554.6000 253.5000 1555.8000 253.8000 ;
	    RECT 1461.0000 253.2000 1462.2001 253.5000 ;
	    RECT 1489.8000 251.4000 1491.0000 252.6000 ;
	    RECT 1492.2001 250.5000 1493.1000 253.5000 ;
	    RECT 1487.7001 249.6000 1493.1000 250.5000 ;
	    RECT 1487.7001 249.3000 1488.6000 249.6000 ;
	    RECT 1461.0000 243.3000 1462.2001 249.3000 ;
	    RECT 1485.0000 243.3000 1486.2001 249.3000 ;
	    RECT 1487.4000 243.3000 1488.6000 249.3000 ;
	    RECT 1492.2001 249.3000 1493.1000 249.6000 ;
	    RECT 1518.9000 250.5000 1519.8000 253.5000 ;
	    RECT 1521.0000 251.4000 1522.2001 252.6000 ;
	    RECT 1554.6000 251.4000 1555.8000 252.6000 ;
	    RECT 1557.0000 250.5000 1557.9000 253.5000 ;
	    RECT 1518.9000 249.6000 1524.3000 250.5000 ;
	    RECT 1518.9000 249.3000 1519.8000 249.6000 ;
	    RECT 1489.8000 243.3000 1491.0000 248.7000 ;
	    RECT 1492.2001 243.3000 1493.4000 249.3000 ;
	    RECT 1518.6000 243.3000 1519.8000 249.3000 ;
	    RECT 1523.4000 249.3000 1524.3000 249.6000 ;
	    RECT 1552.5000 249.6000 1557.9000 250.5000 ;
	    RECT 1552.5000 249.3000 1553.4000 249.6000 ;
	    RECT 1521.0000 243.3000 1522.2001 248.7000 ;
	    RECT 1523.4000 243.3000 1524.6000 249.3000 ;
	    RECT 1525.8000 243.3000 1527.0000 249.3000 ;
	    RECT 1549.8000 243.3000 1551.0000 249.3000 ;
	    RECT 1552.2001 243.3000 1553.4000 249.3000 ;
	    RECT 1557.0000 249.3000 1557.9000 249.6000 ;
	    RECT 1554.6000 243.3000 1555.8000 248.7000 ;
	    RECT 1557.0000 243.3000 1558.2001 249.3000 ;
	    RECT 1.2000 240.6000 1569.0000 242.4000 ;
	    RECT 126.6000 233.7000 127.8000 239.7000 ;
	    RECT 129.0000 232.5000 130.2000 239.7000 ;
	    RECT 131.4000 233.7000 132.6000 239.7000 ;
	    RECT 133.8000 232.8000 135.0000 239.7000 ;
	    RECT 136.2000 233.7000 137.4000 239.7000 ;
	    RECT 131.1000 231.9000 135.0000 232.8000 ;
	    RECT 25.8000 231.4500 27.0000 231.6000 ;
	    RECT 64.2000 231.4500 65.4000 231.6000 ;
	    RECT 129.0000 231.4500 130.2000 231.6000 ;
	    RECT 25.8000 230.5500 130.2000 231.4500 ;
	    RECT 25.8000 230.4000 27.0000 230.5500 ;
	    RECT 64.2000 230.4000 65.4000 230.5500 ;
	    RECT 129.0000 230.4000 130.2000 230.5500 ;
	    RECT 131.1000 229.5000 132.0000 231.9000 ;
	    RECT 138.6000 231.6000 139.8000 239.7000 ;
	    RECT 141.0000 233.7000 142.2000 239.7000 ;
	    RECT 143.4000 235.5000 144.6000 239.7000 ;
	    RECT 145.8000 235.5000 147.0000 239.7000 ;
	    RECT 148.2000 235.5000 149.4000 239.7000 ;
	    RECT 140.7000 231.6000 147.0000 232.8000 ;
	    RECT 135.9000 230.4000 139.8000 231.6000 ;
	    RECT 150.6000 230.4000 151.8000 239.7000 ;
	    RECT 153.0000 233.7000 154.2000 239.7000 ;
	    RECT 155.4000 232.5000 156.6000 239.7000 ;
	    RECT 157.8000 233.7000 159.0000 239.7000 ;
	    RECT 160.2000 232.5000 161.4000 239.7000 ;
	    RECT 162.6000 235.5000 163.8000 239.7000 ;
	    RECT 165.0000 235.5000 166.2000 239.7000 ;
	    RECT 167.4000 233.7000 168.6000 239.7000 ;
	    RECT 169.8000 232.8000 171.0000 239.7000 ;
	    RECT 172.2000 233.7000 173.4000 240.6000 ;
	    RECT 174.6000 234.6000 175.8000 239.7000 ;
	    RECT 174.6000 233.7000 176.1000 234.6000 ;
	    RECT 177.0000 233.7000 178.2000 239.7000 ;
	    RECT 209.1000 233.7000 210.3000 239.7000 ;
	    RECT 175.2000 232.8000 176.1000 233.7000 ;
	    RECT 168.0000 231.6000 174.3000 232.8000 ;
	    RECT 175.2000 231.9000 178.2000 232.8000 ;
	    RECT 155.4000 230.4000 159.3000 231.6000 ;
	    RECT 160.2000 230.7000 168.9000 231.6000 ;
	    RECT 173.4000 231.0000 174.3000 231.6000 ;
	    RECT 143.4000 229.5000 144.6000 229.8000 ;
	    RECT 129.0000 228.0000 130.2000 229.5000 ;
	    RECT 128.7000 226.8000 130.2000 228.0000 ;
	    RECT 131.1000 228.6000 144.6000 229.5000 ;
	    RECT 148.2000 229.5000 149.4000 229.8000 ;
	    RECT 160.2000 229.5000 161.1000 230.7000 ;
	    RECT 169.8000 229.8000 171.9000 230.7000 ;
	    RECT 173.4000 229.8000 175.8000 231.0000 ;
	    RECT 148.2000 228.6000 161.1000 229.5000 ;
	    RECT 162.6000 229.5000 171.9000 229.8000 ;
	    RECT 162.6000 228.9000 170.7000 229.5000 ;
	    RECT 162.6000 228.6000 163.8000 228.9000 ;
	    RECT 128.7000 220.2000 129.9000 226.8000 ;
	    RECT 131.1000 225.9000 132.0000 228.6000 ;
	    RECT 167.1000 227.7000 168.3000 228.0000 ;
	    RECT 132.9000 226.8000 171.3000 227.7000 ;
	    RECT 172.2000 227.4000 173.4000 228.6000 ;
	    RECT 132.9000 226.5000 134.1000 226.8000 ;
	    RECT 130.8000 225.0000 132.0000 225.9000 ;
	    RECT 141.0000 225.0000 166.5000 225.9000 ;
	    RECT 130.8000 222.0000 131.7000 225.0000 ;
	    RECT 141.0000 224.1000 142.2000 225.0000 ;
	    RECT 167.4000 224.4000 168.6000 225.6000 ;
	    RECT 169.5000 225.0000 176.1000 225.9000 ;
	    RECT 174.9000 224.7000 176.1000 225.0000 ;
	    RECT 132.6000 222.9000 138.3000 224.1000 ;
	    RECT 130.8000 221.1000 132.6000 222.0000 ;
	    RECT 128.7000 219.0000 130.2000 220.2000 ;
	    RECT 126.6000 213.3000 127.8000 216.3000 ;
	    RECT 129.0000 213.3000 130.2000 219.0000 ;
	    RECT 131.4000 213.3000 132.6000 221.1000 ;
	    RECT 137.1000 221.1000 138.3000 222.9000 ;
	    RECT 137.1000 220.2000 139.8000 221.1000 ;
	    RECT 138.6000 219.3000 139.8000 220.2000 ;
	    RECT 145.8000 219.6000 147.0000 223.8000 ;
	    RECT 150.6000 222.9000 155.4000 224.1000 ;
	    RECT 161.1000 222.9000 164.1000 224.1000 ;
	    RECT 177.0000 223.5000 178.2000 231.9000 ;
	    RECT 209.4000 230.4000 210.6000 231.6000 ;
	    RECT 209.4000 229.5000 210.3000 230.4000 ;
	    RECT 211.5000 228.6000 212.7000 239.7000 ;
	    RECT 205.8000 228.4500 207.0000 228.6000 ;
	    RECT 208.2000 228.4500 209.4000 228.6000 ;
	    RECT 205.8000 227.5500 209.4000 228.4500 ;
	    RECT 205.8000 227.4000 207.0000 227.5500 ;
	    RECT 208.2000 227.4000 209.4000 227.5500 ;
	    RECT 211.2000 227.7000 212.7000 228.6000 ;
	    RECT 215.4000 227.7000 216.6000 239.7000 ;
	    RECT 150.0000 221.7000 151.2000 222.0000 ;
	    RECT 150.0000 220.8000 156.6000 221.7000 ;
	    RECT 157.8000 221.4000 159.0000 222.6000 ;
	    RECT 155.4000 220.5000 156.6000 220.8000 ;
	    RECT 157.8000 220.2000 159.0000 220.5000 ;
	    RECT 136.2000 213.3000 137.4000 219.3000 ;
	    RECT 138.6000 218.1000 142.2000 219.3000 ;
	    RECT 145.8000 218.4000 147.3000 219.6000 ;
	    RECT 151.8000 218.4000 152.1000 219.6000 ;
	    RECT 153.0000 218.4000 154.2000 219.6000 ;
	    RECT 155.4000 219.3000 156.6000 219.6000 ;
	    RECT 161.1000 219.3000 162.3000 222.9000 ;
	    RECT 165.0000 222.3000 178.2000 223.5000 ;
	    RECT 211.2000 222.6000 212.1000 227.7000 ;
	    RECT 213.0000 225.4500 214.2000 225.6000 ;
	    RECT 213.0000 224.5500 218.8500 225.4500 ;
	    RECT 213.0000 224.4000 214.2000 224.5500 ;
	    RECT 213.0000 223.2000 214.2000 223.5000 ;
	    RECT 170.1000 220.2000 174.6000 221.4000 ;
	    RECT 170.1000 219.3000 171.3000 220.2000 ;
	    RECT 155.4000 218.4000 162.3000 219.3000 ;
	    RECT 141.0000 213.3000 142.2000 218.1000 ;
	    RECT 167.4000 218.1000 171.3000 219.3000 ;
	    RECT 143.4000 213.3000 144.6000 217.5000 ;
	    RECT 145.8000 213.3000 147.0000 217.5000 ;
	    RECT 148.2000 213.3000 149.4000 217.5000 ;
	    RECT 150.6000 213.3000 151.8000 217.5000 ;
	    RECT 153.0000 213.3000 154.2000 216.3000 ;
	    RECT 155.4000 213.3000 156.6000 217.5000 ;
	    RECT 157.8000 213.3000 159.0000 216.3000 ;
	    RECT 160.2000 213.3000 161.4000 217.5000 ;
	    RECT 162.6000 213.3000 163.8000 217.5000 ;
	    RECT 165.0000 213.3000 166.2000 217.5000 ;
	    RECT 167.4000 213.3000 168.6000 218.1000 ;
	    RECT 172.2000 213.3000 173.4000 219.3000 ;
	    RECT 177.0000 213.3000 178.2000 222.3000 ;
	    RECT 208.2000 221.4000 209.4000 222.6000 ;
	    RECT 210.3000 221.4000 212.1000 222.6000 ;
	    RECT 214.2000 220.8000 214.5000 222.3000 ;
	    RECT 215.4000 221.4000 216.6000 222.6000 ;
	    RECT 217.9500 222.4500 218.8500 224.5500 ;
	    RECT 229.8000 223.5000 231.0000 239.7000 ;
	    RECT 232.2000 233.7000 233.4000 239.7000 ;
	    RECT 246.6000 223.5000 247.8000 239.7000 ;
	    RECT 249.0000 233.7000 250.2000 239.7000 ;
	    RECT 263.4000 223.5000 264.6000 239.7000 ;
	    RECT 265.8000 233.7000 267.0000 239.7000 ;
	    RECT 390.6000 233.7000 391.8000 239.7000 ;
	    RECT 393.0000 232.5000 394.2000 239.7000 ;
	    RECT 395.4000 233.7000 396.6000 239.7000 ;
	    RECT 397.8000 232.8000 399.0000 239.7000 ;
	    RECT 400.2000 233.7000 401.4000 239.7000 ;
	    RECT 395.1000 231.9000 399.0000 232.8000 ;
	    RECT 385.8000 231.4500 387.0000 231.6000 ;
	    RECT 393.0000 231.4500 394.2000 231.6000 ;
	    RECT 385.8000 230.5500 394.2000 231.4500 ;
	    RECT 385.8000 230.4000 387.0000 230.5500 ;
	    RECT 393.0000 230.4000 394.2000 230.5500 ;
	    RECT 395.1000 229.5000 396.0000 231.9000 ;
	    RECT 402.6000 231.6000 403.8000 239.7000 ;
	    RECT 405.0000 233.7000 406.2000 239.7000 ;
	    RECT 407.4000 235.5000 408.6000 239.7000 ;
	    RECT 409.8000 235.5000 411.0000 239.7000 ;
	    RECT 412.2000 235.5000 413.4000 239.7000 ;
	    RECT 404.7000 231.6000 411.0000 232.8000 ;
	    RECT 399.9000 230.4000 403.8000 231.6000 ;
	    RECT 414.6000 230.4000 415.8000 239.7000 ;
	    RECT 417.0000 233.7000 418.2000 239.7000 ;
	    RECT 419.4000 232.5000 420.6000 239.7000 ;
	    RECT 421.8000 233.7000 423.0000 239.7000 ;
	    RECT 424.2000 232.5000 425.4000 239.7000 ;
	    RECT 426.6000 235.5000 427.8000 239.7000 ;
	    RECT 429.0000 235.5000 430.2000 239.7000 ;
	    RECT 431.4000 233.7000 432.6000 239.7000 ;
	    RECT 433.8000 232.8000 435.0000 239.7000 ;
	    RECT 436.2000 233.7000 437.4000 240.6000 ;
	    RECT 438.6000 234.6000 439.8000 239.7000 ;
	    RECT 438.6000 233.7000 440.1000 234.6000 ;
	    RECT 441.0000 233.7000 442.2000 239.7000 ;
	    RECT 439.2000 232.8000 440.1000 233.7000 ;
	    RECT 432.0000 231.6000 438.3000 232.8000 ;
	    RECT 439.2000 231.9000 442.2000 232.8000 ;
	    RECT 419.4000 230.4000 423.3000 231.6000 ;
	    RECT 424.2000 230.7000 432.9000 231.6000 ;
	    RECT 437.4000 231.0000 438.3000 231.6000 ;
	    RECT 407.4000 229.5000 408.6000 229.8000 ;
	    RECT 393.0000 228.0000 394.2000 229.5000 ;
	    RECT 392.7000 226.8000 394.2000 228.0000 ;
	    RECT 395.1000 228.6000 408.6000 229.5000 ;
	    RECT 412.2000 229.5000 413.4000 229.8000 ;
	    RECT 424.2000 229.5000 425.1000 230.7000 ;
	    RECT 433.8000 229.8000 435.9000 230.7000 ;
	    RECT 437.4000 229.8000 439.8000 231.0000 ;
	    RECT 412.2000 228.6000 425.1000 229.5000 ;
	    RECT 426.6000 229.5000 435.9000 229.8000 ;
	    RECT 426.6000 228.9000 434.7000 229.5000 ;
	    RECT 426.6000 228.6000 427.8000 228.9000 ;
	    RECT 285.0000 225.4500 286.2000 225.6000 ;
	    RECT 347.4000 225.4500 348.6000 225.6000 ;
	    RECT 285.0000 224.5500 348.6000 225.4500 ;
	    RECT 285.0000 224.4000 286.2000 224.5500 ;
	    RECT 347.4000 224.4000 348.6000 224.5500 ;
	    RECT 229.8000 222.4500 231.0000 222.6000 ;
	    RECT 217.9500 221.5500 231.0000 222.4500 ;
	    RECT 229.8000 221.4000 231.0000 221.5500 ;
	    RECT 244.2000 222.4500 245.4000 222.6000 ;
	    RECT 246.6000 222.4500 247.8000 222.6000 ;
	    RECT 244.2000 221.5500 247.8000 222.4500 ;
	    RECT 244.2000 221.4000 245.4000 221.5500 ;
	    RECT 246.6000 221.4000 247.8000 221.5500 ;
	    RECT 249.0000 222.4500 250.2000 222.6000 ;
	    RECT 263.4000 222.4500 264.6000 222.6000 ;
	    RECT 337.8000 222.4500 339.0000 222.6000 ;
	    RECT 249.0000 221.5500 339.0000 222.4500 ;
	    RECT 249.0000 221.4000 250.2000 221.5500 ;
	    RECT 263.4000 221.4000 264.6000 221.5500 ;
	    RECT 337.8000 221.4000 339.0000 221.5500 ;
	    RECT 208.5000 219.3000 209.4000 220.5000 ;
	    RECT 210.9000 219.3000 216.3000 219.9000 ;
	    RECT 208.2000 213.3000 209.4000 219.3000 ;
	    RECT 210.6000 219.0000 216.6000 219.3000 ;
	    RECT 210.6000 213.3000 211.8000 219.0000 ;
	    RECT 213.0000 213.3000 214.2000 218.1000 ;
	    RECT 215.4000 213.3000 216.6000 219.0000 ;
	    RECT 229.8000 213.3000 231.0000 220.5000 ;
	    RECT 232.2000 218.4000 233.4000 219.6000 ;
	    RECT 232.2000 217.2000 233.4000 217.5000 ;
	    RECT 232.2000 213.3000 233.4000 216.3000 ;
	    RECT 246.6000 213.3000 247.8000 220.5000 ;
	    RECT 249.0000 219.4500 250.2000 219.6000 ;
	    RECT 253.8000 219.4500 255.0000 219.6000 ;
	    RECT 249.0000 218.5500 255.0000 219.4500 ;
	    RECT 249.0000 218.4000 250.2000 218.5500 ;
	    RECT 253.8000 218.4000 255.0000 218.5500 ;
	    RECT 249.0000 217.2000 250.2000 217.5000 ;
	    RECT 249.0000 213.3000 250.2000 216.3000 ;
	    RECT 263.4000 213.3000 264.6000 220.5000 ;
	    RECT 392.7000 220.2000 393.9000 226.8000 ;
	    RECT 395.1000 225.9000 396.0000 228.6000 ;
	    RECT 431.1000 227.7000 432.3000 228.0000 ;
	    RECT 396.9000 226.8000 435.3000 227.7000 ;
	    RECT 436.2000 227.4000 437.4000 228.6000 ;
	    RECT 396.9000 226.5000 398.1000 226.8000 ;
	    RECT 394.8000 225.0000 396.0000 225.9000 ;
	    RECT 405.0000 225.0000 430.5000 225.9000 ;
	    RECT 394.8000 222.0000 395.7000 225.0000 ;
	    RECT 405.0000 224.1000 406.2000 225.0000 ;
	    RECT 431.4000 224.4000 432.6000 225.6000 ;
	    RECT 433.5000 225.0000 440.1000 225.9000 ;
	    RECT 438.9000 224.7000 440.1000 225.0000 ;
	    RECT 396.6000 222.9000 402.3000 224.1000 ;
	    RECT 394.8000 221.1000 396.6000 222.0000 ;
	    RECT 265.8000 219.4500 267.0000 219.6000 ;
	    RECT 268.2000 219.4500 269.4000 219.6000 ;
	    RECT 364.2000 219.4500 365.4000 219.6000 ;
	    RECT 265.8000 218.5500 365.4000 219.4500 ;
	    RECT 392.7000 219.0000 394.2000 220.2000 ;
	    RECT 265.8000 218.4000 267.0000 218.5500 ;
	    RECT 268.2000 218.4000 269.4000 218.5500 ;
	    RECT 364.2000 218.4000 365.4000 218.5500 ;
	    RECT 265.8000 217.2000 267.0000 217.5000 ;
	    RECT 333.0000 216.4500 334.2000 216.6000 ;
	    RECT 376.2000 216.4500 377.4000 216.6000 ;
	    RECT 265.8000 213.3000 267.0000 216.3000 ;
	    RECT 333.0000 215.5500 377.4000 216.4500 ;
	    RECT 333.0000 215.4000 334.2000 215.5500 ;
	    RECT 376.2000 215.4000 377.4000 215.5500 ;
	    RECT 390.6000 213.3000 391.8000 216.3000 ;
	    RECT 393.0000 213.3000 394.2000 219.0000 ;
	    RECT 395.4000 213.3000 396.6000 221.1000 ;
	    RECT 401.1000 221.1000 402.3000 222.9000 ;
	    RECT 401.1000 220.2000 403.8000 221.1000 ;
	    RECT 402.6000 219.3000 403.8000 220.2000 ;
	    RECT 409.8000 219.6000 411.0000 223.8000 ;
	    RECT 414.6000 222.9000 419.4000 224.1000 ;
	    RECT 425.1000 222.9000 428.1000 224.1000 ;
	    RECT 441.0000 223.5000 442.2000 231.9000 ;
	    RECT 462.6000 223.5000 463.8000 239.7000 ;
	    RECT 465.0000 233.7000 466.2000 239.7000 ;
	    RECT 489.0000 227.7000 490.2000 239.7000 ;
	    RECT 492.9000 228.6000 494.1000 239.7000 ;
	    RECT 495.3000 233.7000 496.5000 239.7000 ;
	    RECT 495.0000 230.4000 496.2000 231.6000 ;
	    RECT 495.3000 229.5000 496.2000 230.4000 ;
	    RECT 492.9000 227.7000 494.4000 228.6000 ;
	    RECT 491.4000 224.4000 492.6000 225.6000 ;
	    RECT 414.0000 221.7000 415.2000 222.0000 ;
	    RECT 414.0000 220.8000 420.6000 221.7000 ;
	    RECT 421.8000 221.4000 423.0000 222.6000 ;
	    RECT 419.4000 220.5000 420.6000 220.8000 ;
	    RECT 421.8000 220.2000 423.0000 220.5000 ;
	    RECT 400.2000 213.3000 401.4000 219.3000 ;
	    RECT 402.6000 218.1000 406.2000 219.3000 ;
	    RECT 409.8000 218.4000 411.3000 219.6000 ;
	    RECT 415.8000 218.4000 416.1000 219.6000 ;
	    RECT 417.0000 218.4000 418.2000 219.6000 ;
	    RECT 419.4000 219.3000 420.6000 219.6000 ;
	    RECT 425.1000 219.3000 426.3000 222.9000 ;
	    RECT 429.0000 222.3000 442.2000 223.5000 ;
	    RECT 491.4000 223.2000 492.6000 223.5000 ;
	    RECT 493.5000 222.6000 494.4000 227.7000 ;
	    RECT 496.2000 227.4000 497.4000 228.6000 ;
	    RECT 510.6000 223.5000 511.8000 239.7000 ;
	    RECT 513.0000 233.7000 514.2000 239.7000 ;
	    RECT 532.2000 233.7000 533.4000 239.7000 ;
	    RECT 534.6000 226.5000 535.8000 239.7000 ;
	    RECT 537.0000 233.7000 538.2000 239.7000 ;
	    RECT 556.2000 233.7000 557.4000 239.7000 ;
	    RECT 537.0000 229.5000 538.2000 229.8000 ;
	    RECT 537.0000 228.4500 538.2000 228.6000 ;
	    RECT 539.4000 228.4500 540.6000 228.6000 ;
	    RECT 537.0000 227.5500 540.6000 228.4500 ;
	    RECT 537.0000 227.4000 538.2000 227.5500 ;
	    RECT 539.4000 227.4000 540.6000 227.5500 ;
	    RECT 558.6000 226.5000 559.8000 239.7000 ;
	    RECT 561.0000 233.7000 562.2000 239.7000 ;
	    RECT 565.8000 239.4000 567.0000 240.6000 ;
	    RECT 575.4000 233.7000 576.6000 239.7000 ;
	    RECT 561.0000 229.5000 562.2000 229.8000 ;
	    RECT 561.0000 228.4500 562.2000 228.6000 ;
	    RECT 565.8000 228.4500 567.0000 228.6000 ;
	    RECT 561.0000 227.5500 567.0000 228.4500 ;
	    RECT 561.0000 227.4000 562.2000 227.5500 ;
	    RECT 565.8000 227.4000 567.0000 227.5500 ;
	    RECT 513.0000 225.4500 514.2000 225.6000 ;
	    RECT 534.6000 225.4500 535.8000 225.6000 ;
	    RECT 513.0000 224.5500 535.8000 225.4500 ;
	    RECT 513.0000 224.4000 514.2000 224.5500 ;
	    RECT 534.6000 224.4000 535.8000 224.5500 ;
	    RECT 558.6000 225.4500 559.8000 225.6000 ;
	    RECT 575.4000 225.4500 576.6000 225.6000 ;
	    RECT 558.6000 224.5500 576.6000 225.4500 ;
	    RECT 558.6000 224.4000 559.8000 224.5500 ;
	    RECT 575.4000 224.4000 576.6000 224.5500 ;
	    RECT 577.8000 223.5000 579.0000 239.7000 ;
	    RECT 604.2000 227.7000 605.4000 239.7000 ;
	    RECT 606.6000 228.3000 607.8000 239.7000 ;
	    RECT 609.0000 233.7000 610.2000 239.7000 ;
	    RECT 611.4000 233.7000 612.6000 239.7000 ;
	    RECT 604.2000 226.5000 605.1000 227.7000 ;
	    RECT 609.0000 227.4000 609.9000 233.7000 ;
	    RECT 637.8000 227.7000 639.0000 239.7000 ;
	    RECT 641.7000 228.6000 642.9000 239.7000 ;
	    RECT 644.1000 233.7000 645.3000 239.7000 ;
	    RECT 671.4000 233.7000 672.6000 239.7000 ;
	    RECT 643.8000 230.4000 645.0000 231.6000 ;
	    RECT 644.1000 229.5000 645.0000 230.4000 ;
	    RECT 671.4000 229.5000 672.6000 229.8000 ;
	    RECT 641.7000 227.7000 643.2000 228.6000 ;
	    RECT 606.3000 226.5000 609.9000 227.4000 ;
	    RECT 604.2000 224.4000 605.4000 225.6000 ;
	    RECT 434.1000 220.2000 438.6000 221.4000 ;
	    RECT 434.1000 219.3000 435.3000 220.2000 ;
	    RECT 419.4000 218.4000 426.3000 219.3000 ;
	    RECT 405.0000 213.3000 406.2000 218.1000 ;
	    RECT 431.4000 218.1000 435.3000 219.3000 ;
	    RECT 407.4000 213.3000 408.6000 217.5000 ;
	    RECT 409.8000 213.3000 411.0000 217.5000 ;
	    RECT 412.2000 213.3000 413.4000 217.5000 ;
	    RECT 414.6000 213.3000 415.8000 217.5000 ;
	    RECT 417.0000 213.3000 418.2000 216.3000 ;
	    RECT 419.4000 213.3000 420.6000 217.5000 ;
	    RECT 421.8000 213.3000 423.0000 216.3000 ;
	    RECT 424.2000 213.3000 425.4000 217.5000 ;
	    RECT 426.6000 213.3000 427.8000 217.5000 ;
	    RECT 429.0000 213.3000 430.2000 217.5000 ;
	    RECT 431.4000 213.3000 432.6000 218.1000 ;
	    RECT 436.2000 213.3000 437.4000 219.3000 ;
	    RECT 441.0000 213.3000 442.2000 222.3000 ;
	    RECT 443.4000 222.4500 444.6000 222.6000 ;
	    RECT 462.6000 222.4500 463.8000 222.6000 ;
	    RECT 443.4000 221.5500 463.8000 222.4500 ;
	    RECT 443.4000 221.4000 444.6000 221.5500 ;
	    RECT 462.6000 221.4000 463.8000 221.5500 ;
	    RECT 489.0000 221.4000 490.2000 222.6000 ;
	    RECT 491.1000 220.8000 491.4000 222.3000 ;
	    RECT 493.5000 221.4000 495.3000 222.6000 ;
	    RECT 496.2000 221.4000 497.4000 222.6000 ;
	    RECT 498.6000 222.4500 499.8000 222.6000 ;
	    RECT 510.6000 222.4500 511.8000 222.6000 ;
	    RECT 498.6000 221.5500 511.8000 222.4500 ;
	    RECT 498.6000 221.4000 499.8000 221.5500 ;
	    RECT 510.6000 221.4000 511.8000 221.5500 ;
	    RECT 532.2000 221.4000 533.4000 222.6000 ;
	    RECT 462.6000 213.3000 463.8000 220.5000 ;
	    RECT 465.0000 219.4500 466.2000 219.6000 ;
	    RECT 479.4000 219.4500 480.6000 219.6000 ;
	    RECT 465.0000 218.5500 480.6000 219.4500 ;
	    RECT 489.3000 219.3000 494.7000 219.9000 ;
	    RECT 496.2000 219.3000 497.1000 220.5000 ;
	    RECT 465.0000 218.4000 466.2000 218.5500 ;
	    RECT 479.4000 218.4000 480.6000 218.5500 ;
	    RECT 489.0000 219.0000 495.0000 219.3000 ;
	    RECT 465.0000 217.2000 466.2000 217.5000 ;
	    RECT 465.0000 213.3000 466.2000 216.3000 ;
	    RECT 489.0000 213.3000 490.2000 219.0000 ;
	    RECT 491.4000 213.3000 492.6000 218.1000 ;
	    RECT 493.8000 213.3000 495.0000 219.0000 ;
	    RECT 496.2000 213.3000 497.4000 219.3000 ;
	    RECT 510.6000 213.3000 511.8000 220.5000 ;
	    RECT 532.2000 220.2000 533.4000 220.5000 ;
	    RECT 513.0000 219.4500 514.2000 219.6000 ;
	    RECT 529.8000 219.4500 531.0000 219.6000 ;
	    RECT 513.0000 218.5500 531.0000 219.4500 ;
	    RECT 534.6000 219.3000 535.8000 223.5000 ;
	    RECT 546.6000 222.4500 547.8000 222.6000 ;
	    RECT 556.2000 222.4500 557.4000 222.6000 ;
	    RECT 546.6000 221.5500 557.4000 222.4500 ;
	    RECT 546.6000 221.4000 547.8000 221.5500 ;
	    RECT 556.2000 221.4000 557.4000 221.5500 ;
	    RECT 556.2000 220.2000 557.4000 220.5000 ;
	    RECT 558.6000 219.3000 559.8000 223.5000 ;
	    RECT 577.8000 222.4500 579.0000 222.6000 ;
	    RECT 601.8000 222.4500 603.0000 222.6000 ;
	    RECT 577.8000 221.5500 603.0000 222.4500 ;
	    RECT 577.8000 221.4000 579.0000 221.5500 ;
	    RECT 601.8000 221.4000 603.0000 221.5500 ;
	    RECT 513.0000 218.4000 514.2000 218.5500 ;
	    RECT 529.8000 218.4000 531.0000 218.5500 ;
	    RECT 513.0000 217.2000 514.2000 217.5000 ;
	    RECT 513.0000 213.3000 514.2000 216.3000 ;
	    RECT 532.2000 213.3000 533.4000 219.3000 ;
	    RECT 534.6000 218.4000 537.3000 219.3000 ;
	    RECT 536.1000 213.3000 537.3000 218.4000 ;
	    RECT 556.2000 213.3000 557.4000 219.3000 ;
	    RECT 558.6000 218.4000 561.3000 219.3000 ;
	    RECT 575.4000 218.4000 576.6000 219.6000 ;
	    RECT 560.1000 213.3000 561.3000 218.4000 ;
	    RECT 575.4000 217.2000 576.6000 217.5000 ;
	    RECT 575.4000 213.3000 576.6000 216.3000 ;
	    RECT 577.8000 213.3000 579.0000 220.5000 ;
	    RECT 604.2000 219.3000 605.1000 223.5000 ;
	    RECT 606.3000 221.4000 607.2000 226.5000 ;
	    RECT 609.0000 224.4000 610.2000 225.6000 ;
	    RECT 633.0000 225.4500 634.2000 225.6000 ;
	    RECT 640.2000 225.4500 641.4000 225.6000 ;
	    RECT 633.0000 224.5500 641.4000 225.4500 ;
	    RECT 633.0000 224.4000 634.2000 224.5500 ;
	    RECT 640.2000 224.4000 641.4000 224.5500 ;
	    RECT 611.4000 223.5000 612.6000 223.8000 ;
	    RECT 609.0000 223.2000 609.9000 223.5000 ;
	    RECT 640.2000 223.2000 641.4000 223.5000 ;
	    RECT 608.4000 222.3000 609.9000 223.2000 ;
	    RECT 642.3000 222.6000 643.2000 227.7000 ;
	    RECT 645.0000 227.4000 646.2000 228.6000 ;
	    RECT 654.6000 228.4500 655.8000 228.6000 ;
	    RECT 671.4000 228.4500 672.6000 228.6000 ;
	    RECT 654.6000 227.5500 672.6000 228.4500 ;
	    RECT 654.6000 227.4000 655.8000 227.5500 ;
	    RECT 671.4000 227.4000 672.6000 227.5500 ;
	    RECT 673.8000 226.5000 675.0000 239.7000 ;
	    RECT 676.2000 233.7000 677.4000 239.7000 ;
	    RECT 688.2000 233.7000 689.4000 239.7000 ;
	    RECT 673.8000 225.4500 675.0000 225.6000 ;
	    RECT 685.8000 225.4500 687.0000 225.6000 ;
	    RECT 673.8000 224.5500 687.0000 225.4500 ;
	    RECT 673.8000 224.4000 675.0000 224.5500 ;
	    RECT 685.8000 224.4000 687.0000 224.5500 ;
	    RECT 690.6000 223.5000 691.8000 239.7000 ;
	    RECT 717.9000 233.7000 719.1000 239.7000 ;
	    RECT 718.2000 230.4000 719.4000 231.6000 ;
	    RECT 718.2000 229.5000 719.1000 230.4000 ;
	    RECT 720.3000 228.6000 721.5000 239.7000 ;
	    RECT 693.0000 228.4500 694.2000 228.6000 ;
	    RECT 717.0000 228.4500 718.2000 228.6000 ;
	    RECT 693.0000 227.5500 718.2000 228.4500 ;
	    RECT 693.0000 227.4000 694.2000 227.5500 ;
	    RECT 717.0000 227.4000 718.2000 227.5500 ;
	    RECT 720.0000 227.7000 721.5000 228.6000 ;
	    RECT 724.2000 227.7000 725.4000 239.7000 ;
	    RECT 743.4000 227.7000 744.6000 239.7000 ;
	    RECT 745.8000 229.5000 747.0000 239.7000 ;
	    RECT 748.2000 228.6000 749.4000 239.7000 ;
	    RECT 762.6000 233.7000 763.8000 239.7000 ;
	    RECT 746.1000 227.7000 749.4000 228.6000 ;
	    RECT 611.4000 222.4500 612.6000 222.6000 ;
	    RECT 613.8000 222.4500 615.0000 222.6000 ;
	    RECT 637.8000 222.4500 639.0000 222.6000 ;
	    RECT 608.4000 222.0000 609.6000 222.3000 ;
	    RECT 611.4000 221.5500 639.0000 222.4500 ;
	    RECT 611.4000 221.4000 612.6000 221.5500 ;
	    RECT 613.8000 221.4000 615.0000 221.5500 ;
	    RECT 637.8000 221.4000 639.0000 221.5500 ;
	    RECT 606.0000 221.1000 607.2000 221.4000 ;
	    RECT 606.0000 220.5000 610.5000 221.1000 ;
	    RECT 639.9000 220.8000 640.2000 222.3000 ;
	    RECT 642.3000 221.4000 644.1000 222.6000 ;
	    RECT 645.0000 221.4000 646.2000 222.6000 ;
	    RECT 606.0000 220.2000 612.3000 220.5000 ;
	    RECT 609.6000 219.6000 612.3000 220.2000 ;
	    RECT 611.4000 219.3000 612.3000 219.6000 ;
	    RECT 638.1000 219.3000 643.5000 219.9000 ;
	    RECT 645.0000 219.3000 645.9000 220.5000 ;
	    RECT 673.8000 219.3000 675.0000 223.5000 ;
	    RECT 720.0000 222.6000 720.9000 227.7000 ;
	    RECT 721.8000 224.4000 723.0000 225.6000 ;
	    RECT 743.4000 224.4000 744.3000 227.7000 ;
	    RECT 746.1000 226.8000 747.0000 227.7000 ;
	    RECT 745.2000 225.6000 747.0000 226.8000 ;
	    RECT 743.4000 223.5000 744.6000 224.4000 ;
	    RECT 721.8000 223.2000 723.0000 223.5000 ;
	    RECT 676.2000 221.4000 677.4000 222.6000 ;
	    RECT 690.6000 222.4500 691.8000 222.6000 ;
	    RECT 693.0000 222.4500 694.2000 222.6000 ;
	    RECT 690.6000 221.5500 694.2000 222.4500 ;
	    RECT 690.6000 221.4000 691.8000 221.5500 ;
	    RECT 693.0000 221.4000 694.2000 221.5500 ;
	    RECT 695.4000 222.4500 696.6000 222.6000 ;
	    RECT 717.0000 222.4500 718.2000 222.6000 ;
	    RECT 695.4000 221.5500 718.2000 222.4500 ;
	    RECT 695.4000 221.4000 696.6000 221.5500 ;
	    RECT 717.0000 221.4000 718.2000 221.5500 ;
	    RECT 719.1000 221.4000 720.9000 222.6000 ;
	    RECT 723.0000 220.8000 723.3000 222.3000 ;
	    RECT 724.2000 221.4000 725.4000 222.6000 ;
	    RECT 743.4000 221.4000 744.6000 222.6000 ;
	    RECT 746.1000 221.1000 747.0000 225.6000 ;
	    RECT 748.2000 225.4500 749.4000 225.6000 ;
	    RECT 750.6000 225.4500 751.8000 225.6000 ;
	    RECT 748.2000 224.5500 751.8000 225.4500 ;
	    RECT 748.2000 224.4000 749.4000 224.5500 ;
	    RECT 750.6000 224.4000 751.8000 224.5500 ;
	    RECT 765.0000 223.5000 766.2000 239.7000 ;
	    RECT 769.8000 239.4000 771.0000 240.6000 ;
	    RECT 789.0000 227.7000 790.2000 239.7000 ;
	    RECT 792.9000 228.6000 794.1000 239.7000 ;
	    RECT 795.3000 233.7000 796.5000 239.7000 ;
	    RECT 928.2000 233.7000 929.4000 239.7000 ;
	    RECT 930.6000 232.5000 931.8000 239.7000 ;
	    RECT 933.0000 233.7000 934.2000 239.7000 ;
	    RECT 935.4000 232.8000 936.6000 239.7000 ;
	    RECT 937.8000 233.7000 939.0000 239.7000 ;
	    RECT 932.7000 231.9000 936.6000 232.8000 ;
	    RECT 795.0000 230.4000 796.2000 231.6000 ;
	    RECT 930.6000 230.4000 931.8000 231.6000 ;
	    RECT 795.3000 229.5000 796.2000 230.4000 ;
	    RECT 932.7000 229.5000 933.6000 231.9000 ;
	    RECT 940.2000 231.6000 941.4000 239.7000 ;
	    RECT 942.6000 233.7000 943.8000 239.7000 ;
	    RECT 945.0000 235.5000 946.2000 239.7000 ;
	    RECT 947.4000 235.5000 948.6000 239.7000 ;
	    RECT 949.8000 235.5000 951.0000 239.7000 ;
	    RECT 942.3000 231.6000 948.6000 232.8000 ;
	    RECT 937.5000 230.4000 941.4000 231.6000 ;
	    RECT 952.2000 230.4000 953.4000 239.7000 ;
	    RECT 954.6000 233.7000 955.8000 239.7000 ;
	    RECT 957.0000 232.5000 958.2000 239.7000 ;
	    RECT 959.4000 233.7000 960.6000 239.7000 ;
	    RECT 961.8000 232.5000 963.0000 239.7000 ;
	    RECT 964.2000 235.5000 965.4000 239.7000 ;
	    RECT 966.6000 235.5000 967.8000 239.7000 ;
	    RECT 969.0000 233.7000 970.2000 239.7000 ;
	    RECT 971.4000 232.8000 972.6000 239.7000 ;
	    RECT 973.8000 233.7000 975.0000 240.6000 ;
	    RECT 976.2000 234.6000 977.4000 239.7000 ;
	    RECT 976.2000 233.7000 977.7000 234.6000 ;
	    RECT 978.6000 233.7000 979.8000 239.7000 ;
	    RECT 976.8000 232.8000 977.7000 233.7000 ;
	    RECT 969.6000 231.6000 975.9000 232.8000 ;
	    RECT 976.8000 231.9000 979.8000 232.8000 ;
	    RECT 957.0000 230.4000 960.9000 231.6000 ;
	    RECT 961.8000 230.7000 970.5000 231.6000 ;
	    RECT 975.0000 231.0000 975.9000 231.6000 ;
	    RECT 945.0000 229.5000 946.2000 229.8000 ;
	    RECT 792.9000 227.7000 794.4000 228.6000 ;
	    RECT 791.4000 225.4500 792.6000 225.6000 ;
	    RECT 767.5500 224.5500 792.6000 225.4500 ;
	    RECT 748.2000 223.2000 749.4000 223.5000 ;
	    RECT 765.0000 222.4500 766.2000 222.6000 ;
	    RECT 767.5500 222.4500 768.4500 224.5500 ;
	    RECT 791.4000 224.4000 792.6000 224.5500 ;
	    RECT 791.4000 223.2000 792.6000 223.5000 ;
	    RECT 793.5000 222.6000 794.4000 227.7000 ;
	    RECT 796.2000 227.4000 797.4000 228.6000 ;
	    RECT 930.6000 228.0000 931.8000 229.5000 ;
	    RECT 930.3000 226.8000 931.8000 228.0000 ;
	    RECT 932.7000 228.6000 946.2000 229.5000 ;
	    RECT 949.8000 229.5000 951.0000 229.8000 ;
	    RECT 961.8000 229.5000 962.7000 230.7000 ;
	    RECT 971.4000 229.8000 973.5000 230.7000 ;
	    RECT 975.0000 229.8000 977.4000 231.0000 ;
	    RECT 949.8000 228.6000 962.7000 229.5000 ;
	    RECT 964.2000 229.5000 973.5000 229.8000 ;
	    RECT 964.2000 228.9000 972.3000 229.5000 ;
	    RECT 964.2000 228.6000 965.4000 228.9000 ;
	    RECT 765.0000 221.5500 768.4500 222.4500 ;
	    RECT 769.8000 222.4500 771.0000 222.6000 ;
	    RECT 789.0000 222.4500 790.2000 222.6000 ;
	    RECT 769.8000 221.5500 790.2000 222.4500 ;
	    RECT 765.0000 221.4000 766.2000 221.5500 ;
	    RECT 769.8000 221.4000 771.0000 221.5500 ;
	    RECT 789.0000 221.4000 790.2000 221.5500 ;
	    RECT 676.2000 220.2000 677.4000 220.5000 ;
	    RECT 604.2000 217.8000 606.3000 219.3000 ;
	    RECT 605.1000 213.3000 606.3000 217.8000 ;
	    RECT 607.5000 213.3000 608.7000 219.0000 ;
	    RECT 611.4000 213.3000 612.6000 219.3000 ;
	    RECT 637.8000 219.0000 643.8000 219.3000 ;
	    RECT 637.8000 213.3000 639.0000 219.0000 ;
	    RECT 640.2000 213.3000 641.4000 218.1000 ;
	    RECT 642.6000 213.3000 643.8000 219.0000 ;
	    RECT 645.0000 213.3000 646.2000 219.3000 ;
	    RECT 672.3000 218.4000 675.0000 219.3000 ;
	    RECT 672.3000 213.3000 673.5000 218.4000 ;
	    RECT 676.2000 213.3000 677.4000 219.3000 ;
	    RECT 688.2000 218.4000 689.4000 219.6000 ;
	    RECT 688.2000 217.2000 689.4000 217.5000 ;
	    RECT 688.2000 213.3000 689.4000 216.3000 ;
	    RECT 690.6000 213.3000 691.8000 220.5000 ;
	    RECT 717.3000 219.3000 718.2000 220.5000 ;
	    RECT 719.7000 219.3000 725.1000 219.9000 ;
	    RECT 717.0000 213.3000 718.2000 219.3000 ;
	    RECT 719.4000 219.0000 725.4000 219.3000 ;
	    RECT 719.4000 213.3000 720.6000 219.0000 ;
	    RECT 721.8000 213.3000 723.0000 218.1000 ;
	    RECT 724.2000 213.3000 725.4000 219.0000 ;
	    RECT 743.4000 213.3000 744.6000 220.5000 ;
	    RECT 746.1000 220.2000 749.4000 221.1000 ;
	    RECT 791.1000 220.8000 791.4000 222.3000 ;
	    RECT 793.5000 221.4000 795.3000 222.6000 ;
	    RECT 796.2000 222.4500 797.4000 222.6000 ;
	    RECT 928.2000 222.4500 929.4000 222.6000 ;
	    RECT 796.2000 221.5500 929.4000 222.4500 ;
	    RECT 796.2000 221.4000 797.4000 221.5500 ;
	    RECT 928.2000 221.4000 929.4000 221.5500 ;
	    RECT 745.8000 213.3000 747.0000 219.3000 ;
	    RECT 748.2000 213.3000 749.4000 220.2000 ;
	    RECT 762.6000 218.4000 763.8000 219.6000 ;
	    RECT 762.6000 217.2000 763.8000 217.5000 ;
	    RECT 762.6000 213.3000 763.8000 216.3000 ;
	    RECT 765.0000 213.3000 766.2000 220.5000 ;
	    RECT 789.3000 219.3000 794.7000 219.9000 ;
	    RECT 796.2000 219.3000 797.1000 220.5000 ;
	    RECT 930.3000 220.2000 931.5000 226.8000 ;
	    RECT 932.7000 225.9000 933.6000 228.6000 ;
	    RECT 968.7000 227.7000 969.9000 228.0000 ;
	    RECT 934.5000 226.8000 972.9000 227.7000 ;
	    RECT 973.8000 227.4000 975.0000 228.6000 ;
	    RECT 934.5000 226.5000 935.7000 226.8000 ;
	    RECT 932.4000 225.0000 933.6000 225.9000 ;
	    RECT 942.6000 225.0000 968.1000 225.9000 ;
	    RECT 932.4000 222.0000 933.3000 225.0000 ;
	    RECT 942.6000 224.1000 943.8000 225.0000 ;
	    RECT 969.0000 224.4000 970.2000 225.6000 ;
	    RECT 971.1000 225.0000 977.7000 225.9000 ;
	    RECT 976.5000 224.7000 977.7000 225.0000 ;
	    RECT 934.2000 222.9000 939.9000 224.1000 ;
	    RECT 932.4000 221.1000 934.2000 222.0000 ;
	    RECT 789.0000 219.0000 795.0000 219.3000 ;
	    RECT 789.0000 213.3000 790.2000 219.0000 ;
	    RECT 791.4000 213.3000 792.6000 218.1000 ;
	    RECT 793.8000 213.3000 795.0000 219.0000 ;
	    RECT 796.2000 213.3000 797.4000 219.3000 ;
	    RECT 930.3000 219.0000 931.8000 220.2000 ;
	    RECT 928.2000 213.3000 929.4000 216.3000 ;
	    RECT 930.6000 213.3000 931.8000 219.0000 ;
	    RECT 933.0000 213.3000 934.2000 221.1000 ;
	    RECT 938.7000 221.1000 939.9000 222.9000 ;
	    RECT 938.7000 220.2000 941.4000 221.1000 ;
	    RECT 940.2000 219.3000 941.4000 220.2000 ;
	    RECT 947.4000 219.6000 948.6000 223.8000 ;
	    RECT 952.2000 222.9000 957.0000 224.1000 ;
	    RECT 962.7000 222.9000 965.7000 224.1000 ;
	    RECT 978.6000 223.5000 979.8000 231.9000 ;
	    RECT 1002.6000 227.7000 1003.8000 239.7000 ;
	    RECT 1006.5000 228.6000 1007.7000 239.7000 ;
	    RECT 1008.9000 233.7000 1010.1000 239.7000 ;
	    RECT 1029.0000 233.7000 1030.2001 239.7000 ;
	    RECT 1008.6000 230.4000 1009.8000 231.6000 ;
	    RECT 1008.9000 229.5000 1009.8000 230.4000 ;
	    RECT 1029.0000 229.5000 1030.2001 229.8000 ;
	    RECT 1006.5000 227.7000 1008.0000 228.6000 ;
	    RECT 997.8000 225.4500 999.0000 225.6000 ;
	    RECT 1005.0000 225.4500 1006.2000 225.6000 ;
	    RECT 997.8000 224.5500 1006.2000 225.4500 ;
	    RECT 997.8000 224.4000 999.0000 224.5500 ;
	    RECT 1005.0000 224.4000 1006.2000 224.5500 ;
	    RECT 951.6000 221.7000 952.8000 222.0000 ;
	    RECT 951.6000 220.8000 958.2000 221.7000 ;
	    RECT 959.4000 221.4000 960.6000 222.6000 ;
	    RECT 957.0000 220.5000 958.2000 220.8000 ;
	    RECT 959.4000 220.2000 960.6000 220.5000 ;
	    RECT 937.8000 213.3000 939.0000 219.3000 ;
	    RECT 940.2000 218.1000 943.8000 219.3000 ;
	    RECT 947.4000 218.4000 948.9000 219.6000 ;
	    RECT 953.4000 218.4000 953.7000 219.6000 ;
	    RECT 954.6000 218.4000 955.8000 219.6000 ;
	    RECT 957.0000 219.3000 958.2000 219.6000 ;
	    RECT 962.7000 219.3000 963.9000 222.9000 ;
	    RECT 966.6000 222.3000 979.8000 223.5000 ;
	    RECT 1005.0000 223.2000 1006.2000 223.5000 ;
	    RECT 1007.1000 222.6000 1008.0000 227.7000 ;
	    RECT 1009.8000 227.4000 1011.0000 228.6000 ;
	    RECT 1029.0000 227.4000 1030.2001 228.6000 ;
	    RECT 1009.9500 225.4500 1010.8500 227.4000 ;
	    RECT 1031.4000 226.5000 1032.6000 239.7000 ;
	    RECT 1033.8000 233.7000 1035.0000 239.7000 ;
	    RECT 1057.8000 227.7000 1059.0000 239.7000 ;
	    RECT 1061.7001 228.6000 1062.9000 239.7000 ;
	    RECT 1064.1000 233.7000 1065.3000 239.7000 ;
	    RECT 1084.2001 233.7000 1085.4000 239.7000 ;
	    RECT 1063.8000 230.4000 1065.0000 231.6000 ;
	    RECT 1064.1000 229.5000 1065.0000 230.4000 ;
	    RECT 1061.7001 227.7000 1063.2001 228.6000 ;
	    RECT 1017.0000 225.4500 1018.2000 225.6000 ;
	    RECT 1031.4000 225.4500 1032.6000 225.6000 ;
	    RECT 1009.9500 224.5500 1058.8500 225.4500 ;
	    RECT 1017.0000 224.4000 1018.2000 224.5500 ;
	    RECT 1031.4000 224.4000 1032.6000 224.5500 ;
	    RECT 971.7000 220.2000 976.2000 221.4000 ;
	    RECT 971.7000 219.3000 972.9000 220.2000 ;
	    RECT 957.0000 218.4000 963.9000 219.3000 ;
	    RECT 942.6000 213.3000 943.8000 218.1000 ;
	    RECT 969.0000 218.1000 972.9000 219.3000 ;
	    RECT 945.0000 213.3000 946.2000 217.5000 ;
	    RECT 947.4000 213.3000 948.6000 217.5000 ;
	    RECT 949.8000 213.3000 951.0000 217.5000 ;
	    RECT 952.2000 213.3000 953.4000 217.5000 ;
	    RECT 954.6000 213.3000 955.8000 216.3000 ;
	    RECT 957.0000 213.3000 958.2000 217.5000 ;
	    RECT 959.4000 213.3000 960.6000 216.3000 ;
	    RECT 961.8000 213.3000 963.0000 217.5000 ;
	    RECT 964.2000 213.3000 965.4000 217.5000 ;
	    RECT 966.6000 213.3000 967.8000 217.5000 ;
	    RECT 969.0000 213.3000 970.2000 218.1000 ;
	    RECT 973.8000 213.3000 975.0000 219.3000 ;
	    RECT 978.6000 213.3000 979.8000 222.3000 ;
	    RECT 995.4000 222.4500 996.6000 222.6000 ;
	    RECT 1002.6000 222.4500 1003.8000 222.6000 ;
	    RECT 995.4000 221.5500 1003.8000 222.4500 ;
	    RECT 995.4000 221.4000 996.6000 221.5500 ;
	    RECT 1002.6000 221.4000 1003.8000 221.5500 ;
	    RECT 1004.7000 220.8000 1005.0000 222.3000 ;
	    RECT 1007.1000 221.4000 1008.9000 222.6000 ;
	    RECT 1009.8000 222.4500 1011.0000 222.6000 ;
	    RECT 1024.2001 222.4500 1025.4000 222.6000 ;
	    RECT 1009.8000 221.5500 1025.4000 222.4500 ;
	    RECT 1009.8000 221.4000 1011.0000 221.5500 ;
	    RECT 1024.2001 221.4000 1025.4000 221.5500 ;
	    RECT 1002.9000 219.3000 1008.3000 219.9000 ;
	    RECT 1009.8000 219.3000 1010.7000 220.5000 ;
	    RECT 1031.4000 219.3000 1032.6000 223.5000 ;
	    RECT 1057.9501 222.6000 1058.8500 224.5500 ;
	    RECT 1060.2001 224.4000 1061.4000 225.6000 ;
	    RECT 1060.2001 223.2000 1061.4000 223.5000 ;
	    RECT 1062.3000 222.6000 1063.2001 227.7000 ;
	    RECT 1065.0000 228.4500 1066.2001 228.6000 ;
	    RECT 1067.4000 228.4500 1068.6000 228.6000 ;
	    RECT 1065.0000 227.5500 1068.6000 228.4500 ;
	    RECT 1065.0000 227.4000 1066.2001 227.5500 ;
	    RECT 1067.4000 227.4000 1068.6000 227.5500 ;
	    RECT 1086.6000 226.5000 1087.8000 239.7000 ;
	    RECT 1089.0000 233.7000 1090.2001 239.7000 ;
	    RECT 1108.2001 233.7000 1109.4000 239.7000 ;
	    RECT 1089.0000 229.5000 1090.2001 229.8000 ;
	    RECT 1089.0000 227.4000 1090.2001 228.6000 ;
	    RECT 1110.6000 226.5000 1111.8000 239.7000 ;
	    RECT 1113.0000 233.7000 1114.2001 239.7000 ;
	    RECT 1139.4000 233.7000 1140.6000 239.7000 ;
	    RECT 1113.0000 229.5000 1114.2001 229.8000 ;
	    RECT 1139.4000 229.5000 1140.6000 229.8000 ;
	    RECT 1113.0000 228.4500 1114.2001 228.6000 ;
	    RECT 1139.4000 228.4500 1140.6000 228.6000 ;
	    RECT 1113.0000 227.5500 1140.6000 228.4500 ;
	    RECT 1113.0000 227.4000 1114.2001 227.5500 ;
	    RECT 1139.4000 227.4000 1140.6000 227.5500 ;
	    RECT 1141.8000 226.5000 1143.0000 239.7000 ;
	    RECT 1144.2001 233.7000 1145.4000 239.7000 ;
	    RECT 1163.4000 233.7000 1164.6000 239.7000 ;
	    RECT 1165.8000 226.5000 1167.0000 239.7000 ;
	    RECT 1168.2001 233.7000 1169.4000 239.7000 ;
	    RECT 1170.6000 234.4500 1171.8000 234.6000 ;
	    RECT 1192.2001 234.4500 1193.4000 234.6000 ;
	    RECT 1170.6000 233.5500 1193.4000 234.4500 ;
	    RECT 1170.6000 233.4000 1171.8000 233.5500 ;
	    RECT 1192.2001 233.4000 1193.4000 233.5500 ;
	    RECT 1168.2001 229.5000 1169.4000 229.8000 ;
	    RECT 1168.2001 228.4500 1169.4000 228.6000 ;
	    RECT 1173.0000 228.4500 1174.2001 228.6000 ;
	    RECT 1185.0000 228.4500 1186.2001 228.6000 ;
	    RECT 1168.2001 227.5500 1186.2001 228.4500 ;
	    RECT 1194.6000 227.7000 1195.8000 239.7000 ;
	    RECT 1198.5000 228.6000 1199.7001 239.7000 ;
	    RECT 1200.9000 233.7000 1202.1000 239.7000 ;
	    RECT 1200.6000 230.4000 1201.8000 231.6000 ;
	    RECT 1200.9000 229.5000 1201.8000 230.4000 ;
	    RECT 1198.5000 227.7000 1200.0000 228.6000 ;
	    RECT 1168.2001 227.4000 1169.4000 227.5500 ;
	    RECT 1173.0000 227.4000 1174.2001 227.5500 ;
	    RECT 1185.0000 227.4000 1186.2001 227.5500 ;
	    RECT 1086.6000 225.4500 1087.8000 225.6000 ;
	    RECT 1101.0000 225.4500 1102.2001 225.6000 ;
	    RECT 1086.6000 224.5500 1102.2001 225.4500 ;
	    RECT 1086.6000 224.4000 1087.8000 224.5500 ;
	    RECT 1101.0000 224.4000 1102.2001 224.5500 ;
	    RECT 1110.6000 225.4500 1111.8000 225.6000 ;
	    RECT 1137.0000 225.4500 1138.2001 225.6000 ;
	    RECT 1110.6000 224.5500 1138.2001 225.4500 ;
	    RECT 1110.6000 224.4000 1111.8000 224.5500 ;
	    RECT 1137.0000 224.4000 1138.2001 224.5500 ;
	    RECT 1141.8000 225.4500 1143.0000 225.6000 ;
	    RECT 1156.2001 225.4500 1157.4000 225.6000 ;
	    RECT 1141.8000 224.5500 1157.4000 225.4500 ;
	    RECT 1141.8000 224.4000 1143.0000 224.5500 ;
	    RECT 1156.2001 224.4000 1157.4000 224.5500 ;
	    RECT 1165.8000 225.4500 1167.0000 225.6000 ;
	    RECT 1187.4000 225.4500 1188.6000 225.6000 ;
	    RECT 1197.0000 225.4500 1198.2001 225.6000 ;
	    RECT 1165.8000 224.5500 1186.0500 225.4500 ;
	    RECT 1165.8000 224.4000 1167.0000 224.5500 ;
	    RECT 1033.8000 221.4000 1035.0000 222.6000 ;
	    RECT 1057.8000 221.4000 1059.0000 222.6000 ;
	    RECT 1059.9000 220.8000 1060.2001 222.3000 ;
	    RECT 1062.3000 221.4000 1064.1000 222.6000 ;
	    RECT 1065.0000 222.4500 1066.2001 222.6000 ;
	    RECT 1079.4000 222.4500 1080.6000 222.6000 ;
	    RECT 1065.0000 221.5500 1080.6000 222.4500 ;
	    RECT 1065.0000 221.4000 1066.2001 221.5500 ;
	    RECT 1079.4000 221.4000 1080.6000 221.5500 ;
	    RECT 1084.2001 221.4000 1085.4000 222.6000 ;
	    RECT 1033.8000 220.2000 1035.0000 220.5000 ;
	    RECT 1058.1000 219.3000 1063.5000 219.9000 ;
	    RECT 1065.0000 219.3000 1065.9000 220.5000 ;
	    RECT 1084.2001 220.2000 1085.4000 220.5000 ;
	    RECT 1086.6000 219.3000 1087.8000 223.5000 ;
	    RECT 1089.0000 222.4500 1090.2001 222.6000 ;
	    RECT 1108.2001 222.4500 1109.4000 222.6000 ;
	    RECT 1089.0000 221.5500 1109.4000 222.4500 ;
	    RECT 1089.0000 221.4000 1090.2001 221.5500 ;
	    RECT 1108.2001 221.4000 1109.4000 221.5500 ;
	    RECT 1108.2001 220.2000 1109.4000 220.5000 ;
	    RECT 1110.6000 219.3000 1111.8000 223.5000 ;
	    RECT 1141.8000 219.3000 1143.0000 223.5000 ;
	    RECT 1144.2001 222.4500 1145.4000 222.6000 ;
	    RECT 1146.6000 222.4500 1147.8000 222.6000 ;
	    RECT 1144.2001 221.5500 1147.8000 222.4500 ;
	    RECT 1144.2001 221.4000 1145.4000 221.5500 ;
	    RECT 1146.6000 221.4000 1147.8000 221.5500 ;
	    RECT 1163.4000 221.4000 1164.6000 222.6000 ;
	    RECT 1144.2001 220.2000 1145.4000 220.5000 ;
	    RECT 1163.4000 220.2000 1164.6000 220.5000 ;
	    RECT 1165.8000 219.3000 1167.0000 223.5000 ;
	    RECT 1185.1500 222.4500 1186.0500 224.5500 ;
	    RECT 1187.4000 224.5500 1198.2001 225.4500 ;
	    RECT 1187.4000 224.4000 1188.6000 224.5500 ;
	    RECT 1197.0000 224.4000 1198.2001 224.5500 ;
	    RECT 1197.0000 223.2000 1198.2001 223.5000 ;
	    RECT 1199.1000 222.6000 1200.0000 227.7000 ;
	    RECT 1201.8000 228.4500 1203.0000 228.6000 ;
	    RECT 1206.6000 228.4500 1207.8000 228.6000 ;
	    RECT 1201.8000 227.5500 1207.8000 228.4500 ;
	    RECT 1228.2001 227.7000 1229.4000 239.7000 ;
	    RECT 1232.1000 228.6000 1233.3000 239.7000 ;
	    RECT 1234.5000 233.7000 1235.7001 239.7000 ;
	    RECT 1259.4000 233.7000 1260.6000 239.7000 ;
	    RECT 1261.8000 234.3000 1263.0000 239.7000 ;
	    RECT 1259.7001 233.4000 1260.6000 233.7000 ;
	    RECT 1264.2001 233.7000 1265.4000 239.7000 ;
	    RECT 1266.6000 233.7000 1267.8000 239.7000 ;
	    RECT 1290.6000 233.7000 1291.8000 239.7000 ;
	    RECT 1293.0000 233.7000 1294.2001 239.7000 ;
	    RECT 1295.4000 234.3000 1296.6000 239.7000 ;
	    RECT 1264.2001 233.4000 1265.1000 233.7000 ;
	    RECT 1259.7001 232.5000 1265.1000 233.4000 ;
	    RECT 1293.3000 233.4000 1294.2001 233.7000 ;
	    RECT 1297.8000 233.7000 1299.0000 239.7000 ;
	    RECT 1297.8000 233.4000 1298.7001 233.7000 ;
	    RECT 1293.3000 232.5000 1298.7001 233.4000 ;
	    RECT 1234.2001 230.4000 1235.4000 231.6000 ;
	    RECT 1234.5000 229.5000 1235.4000 230.4000 ;
	    RECT 1259.7001 229.5000 1260.6000 232.5000 ;
	    RECT 1261.8000 231.4500 1263.0000 231.6000 ;
	    RECT 1295.4000 231.4500 1296.6000 231.6000 ;
	    RECT 1261.8000 230.5500 1296.6000 231.4500 ;
	    RECT 1261.8000 230.4000 1263.0000 230.5500 ;
	    RECT 1295.4000 230.4000 1296.6000 230.5500 ;
	    RECT 1297.8000 229.5000 1298.7001 232.5000 ;
	    RECT 1261.8000 229.2000 1263.0000 229.5000 ;
	    RECT 1295.4000 229.2000 1296.6000 229.5000 ;
	    RECT 1232.1000 227.7000 1233.6000 228.6000 ;
	    RECT 1201.8000 227.4000 1203.0000 227.5500 ;
	    RECT 1206.6000 227.4000 1207.8000 227.5500 ;
	    RECT 1201.8000 225.4500 1203.0000 225.6000 ;
	    RECT 1209.0000 225.4500 1210.2001 225.6000 ;
	    RECT 1201.8000 224.5500 1210.2001 225.4500 ;
	    RECT 1201.8000 224.4000 1203.0000 224.5500 ;
	    RECT 1209.0000 224.4000 1210.2001 224.5500 ;
	    RECT 1211.4000 225.4500 1212.6000 225.6000 ;
	    RECT 1230.6000 225.4500 1231.8000 225.6000 ;
	    RECT 1211.4000 224.5500 1231.8000 225.4500 ;
	    RECT 1211.4000 224.4000 1212.6000 224.5500 ;
	    RECT 1230.6000 224.4000 1231.8000 224.5500 ;
	    RECT 1230.6000 223.2000 1231.8000 223.5000 ;
	    RECT 1232.7001 222.6000 1233.6000 227.7000 ;
	    RECT 1235.4000 228.4500 1236.6000 228.6000 ;
	    RECT 1245.0000 228.4500 1246.2001 228.6000 ;
	    RECT 1235.4000 227.5500 1246.2001 228.4500 ;
	    RECT 1235.4000 227.4000 1236.6000 227.5500 ;
	    RECT 1245.0000 227.4000 1246.2001 227.5500 ;
	    RECT 1259.4000 227.4000 1260.6000 228.6000 ;
	    RECT 1266.6000 227.4000 1267.8000 228.6000 ;
	    RECT 1290.6000 227.4000 1291.8000 228.6000 ;
	    RECT 1297.8000 228.4500 1299.0000 228.6000 ;
	    RECT 1305.0000 228.4500 1306.2001 228.6000 ;
	    RECT 1297.8000 227.5500 1306.2001 228.4500 ;
	    RECT 1297.8000 227.4000 1299.0000 227.5500 ;
	    RECT 1305.0000 227.4000 1306.2001 227.5500 ;
	    RECT 1259.7001 222.6000 1260.6000 226.5000 ;
	    RECT 1266.6000 226.2000 1267.8000 226.5000 ;
	    RECT 1290.6000 226.2000 1291.8000 226.5000 ;
	    RECT 1263.0000 224.4000 1263.3000 225.6000 ;
	    RECT 1264.2001 224.4000 1265.4000 225.6000 ;
	    RECT 1293.0000 224.4000 1294.2001 225.6000 ;
	    RECT 1295.1000 224.4000 1295.4000 225.6000 ;
	    RECT 1297.8000 222.6000 1298.7001 226.5000 ;
	    RECT 1309.8000 223.5000 1311.0000 239.7000 ;
	    RECT 1312.2001 233.7000 1313.4000 239.7000 ;
	    RECT 1336.2001 233.7000 1337.4000 239.7000 ;
	    RECT 1338.6000 234.3000 1339.8000 239.7000 ;
	    RECT 1336.5000 233.4000 1337.4000 233.7000 ;
	    RECT 1341.0000 233.7000 1342.2001 239.7000 ;
	    RECT 1343.4000 233.7000 1344.6000 239.7000 ;
	    RECT 1377.0000 233.7000 1378.2001 239.7000 ;
	    RECT 1379.4000 233.7000 1380.6000 239.7000 ;
	    RECT 1381.8000 234.3000 1383.0000 239.7000 ;
	    RECT 1341.0000 233.4000 1341.9000 233.7000 ;
	    RECT 1336.5000 232.5000 1341.9000 233.4000 ;
	    RECT 1379.7001 233.4000 1380.6000 233.7000 ;
	    RECT 1384.2001 233.7000 1385.4000 239.7000 ;
	    RECT 1409.1000 233.7000 1410.3000 239.7000 ;
	    RECT 1384.2001 233.4000 1385.1000 233.7000 ;
	    RECT 1379.7001 232.5000 1385.1000 233.4000 ;
	    RECT 1336.5000 229.5000 1337.4000 232.5000 ;
	    RECT 1338.6000 231.4500 1339.8000 231.6000 ;
	    RECT 1343.4000 231.4500 1344.6000 231.6000 ;
	    RECT 1381.8000 231.4500 1383.0000 231.6000 ;
	    RECT 1338.6000 230.5500 1383.0000 231.4500 ;
	    RECT 1338.6000 230.4000 1339.8000 230.5500 ;
	    RECT 1343.4000 230.4000 1344.6000 230.5500 ;
	    RECT 1381.8000 230.4000 1383.0000 230.5500 ;
	    RECT 1384.2001 229.5000 1385.1000 232.5000 ;
	    RECT 1409.4000 230.4000 1410.6000 231.6000 ;
	    RECT 1409.4000 229.5000 1410.3000 230.4000 ;
	    RECT 1338.6000 229.2000 1339.8000 229.5000 ;
	    RECT 1381.8000 229.2000 1383.0000 229.5000 ;
	    RECT 1411.5000 228.6000 1412.7001 239.7000 ;
	    RECT 1329.0000 228.4500 1330.2001 228.6000 ;
	    RECT 1336.2001 228.4500 1337.4000 228.6000 ;
	    RECT 1329.0000 227.5500 1337.4000 228.4500 ;
	    RECT 1329.0000 227.4000 1330.2001 227.5500 ;
	    RECT 1336.2001 227.4000 1337.4000 227.5500 ;
	    RECT 1341.0000 228.4500 1342.2001 228.6000 ;
	    RECT 1343.4000 228.4500 1344.6000 228.6000 ;
	    RECT 1341.0000 227.5500 1344.6000 228.4500 ;
	    RECT 1341.0000 227.4000 1342.2001 227.5500 ;
	    RECT 1343.4000 227.4000 1344.6000 227.5500 ;
	    RECT 1377.0000 227.4000 1378.2001 228.6000 ;
	    RECT 1384.2001 228.4500 1385.4000 228.6000 ;
	    RECT 1405.8000 228.4500 1407.0000 228.6000 ;
	    RECT 1384.2001 227.5500 1407.0000 228.4500 ;
	    RECT 1384.2001 227.4000 1385.4000 227.5500 ;
	    RECT 1405.8000 227.4000 1407.0000 227.5500 ;
	    RECT 1408.2001 227.4000 1409.4000 228.6000 ;
	    RECT 1411.2001 227.7000 1412.7001 228.6000 ;
	    RECT 1415.4000 227.7000 1416.6000 239.7000 ;
	    RECT 1429.8000 233.7000 1431.0000 239.7000 ;
	    RECT 1336.5000 222.6000 1337.4000 226.5000 ;
	    RECT 1343.4000 226.2000 1344.6000 226.5000 ;
	    RECT 1377.0000 226.2000 1378.2001 226.5000 ;
	    RECT 1339.8000 224.4000 1340.1000 225.6000 ;
	    RECT 1341.0000 224.4000 1342.2001 225.6000 ;
	    RECT 1379.4000 224.4000 1380.6000 225.6000 ;
	    RECT 1381.5000 224.4000 1381.8000 225.6000 ;
	    RECT 1384.2001 222.6000 1385.1000 226.5000 ;
	    RECT 1411.2001 222.6000 1412.1000 227.7000 ;
	    RECT 1413.0000 225.4500 1414.2001 225.6000 ;
	    RECT 1429.8000 225.4500 1431.0000 225.6000 ;
	    RECT 1413.0000 224.5500 1431.0000 225.4500 ;
	    RECT 1413.0000 224.4000 1414.2001 224.5500 ;
	    RECT 1429.8000 224.4000 1431.0000 224.5500 ;
	    RECT 1432.2001 223.5000 1433.4000 239.7000 ;
	    RECT 1446.6000 223.5000 1447.8000 239.7000 ;
	    RECT 1449.0000 233.7000 1450.2001 239.7000 ;
	    RECT 1473.0000 233.7000 1474.2001 239.7000 ;
	    RECT 1475.4000 233.7000 1476.6000 239.7000 ;
	    RECT 1477.8000 234.3000 1479.0000 239.7000 ;
	    RECT 1475.7001 233.4000 1476.6000 233.7000 ;
	    RECT 1480.2001 233.7000 1481.4000 239.7000 ;
	    RECT 1506.6000 233.7000 1507.8000 239.7000 ;
	    RECT 1509.0000 234.3000 1510.2001 239.7000 ;
	    RECT 1480.2001 233.4000 1481.1000 233.7000 ;
	    RECT 1475.7001 232.5000 1481.1000 233.4000 ;
	    RECT 1470.6000 231.4500 1471.8000 231.6000 ;
	    RECT 1477.8000 231.4500 1479.0000 231.6000 ;
	    RECT 1470.6000 230.5500 1479.0000 231.4500 ;
	    RECT 1470.6000 230.4000 1471.8000 230.5500 ;
	    RECT 1477.8000 230.4000 1479.0000 230.5500 ;
	    RECT 1480.2001 229.5000 1481.1000 232.5000 ;
	    RECT 1506.9000 233.4000 1507.8000 233.7000 ;
	    RECT 1511.4000 233.7000 1512.6000 239.7000 ;
	    RECT 1513.8000 233.7000 1515.0000 239.7000 ;
	    RECT 1540.2001 233.7000 1541.4000 239.7000 ;
	    RECT 1542.6000 234.3000 1543.8000 239.7000 ;
	    RECT 1511.4000 233.4000 1512.3000 233.7000 ;
	    RECT 1506.9000 232.5000 1512.3000 233.4000 ;
	    RECT 1540.5000 233.4000 1541.4000 233.7000 ;
	    RECT 1545.0000 233.7000 1546.2001 239.7000 ;
	    RECT 1547.4000 233.7000 1548.6000 239.7000 ;
	    RECT 1545.0000 233.4000 1545.9000 233.7000 ;
	    RECT 1540.5000 232.5000 1545.9000 233.4000 ;
	    RECT 1506.9000 229.5000 1507.8000 232.5000 ;
	    RECT 1509.0000 230.4000 1510.2001 231.6000 ;
	    RECT 1540.5000 229.5000 1541.4000 232.5000 ;
	    RECT 1542.6000 230.4000 1543.8000 231.6000 ;
	    RECT 1477.8000 229.2000 1479.0000 229.5000 ;
	    RECT 1509.0000 229.2000 1510.2001 229.5000 ;
	    RECT 1542.6000 229.2000 1543.8000 229.5000 ;
	    RECT 1473.0000 227.4000 1474.2001 228.6000 ;
	    RECT 1480.2001 227.4000 1481.4000 228.6000 ;
	    RECT 1494.6000 228.4500 1495.8000 228.6000 ;
	    RECT 1506.6000 228.4500 1507.8000 228.6000 ;
	    RECT 1494.6000 227.5500 1507.8000 228.4500 ;
	    RECT 1494.6000 227.4000 1495.8000 227.5500 ;
	    RECT 1506.6000 227.4000 1507.8000 227.5500 ;
	    RECT 1513.8000 227.4000 1515.0000 228.6000 ;
	    RECT 1530.6000 228.4500 1531.8000 228.6000 ;
	    RECT 1540.2001 228.4500 1541.4000 228.6000 ;
	    RECT 1530.6000 227.5500 1541.4000 228.4500 ;
	    RECT 1530.6000 227.4000 1531.8000 227.5500 ;
	    RECT 1540.2001 227.4000 1541.4000 227.5500 ;
	    RECT 1547.4000 227.4000 1548.6000 228.6000 ;
	    RECT 1473.0000 226.2000 1474.2001 226.5000 ;
	    RECT 1475.4000 224.4000 1476.6000 225.6000 ;
	    RECT 1477.5000 224.4000 1477.8000 225.6000 ;
	    RECT 1413.0000 223.2000 1414.2001 223.5000 ;
	    RECT 1480.2001 222.6000 1481.1000 226.5000 ;
	    RECT 1194.6000 222.4500 1195.8000 222.6000 ;
	    RECT 1185.1500 221.5500 1195.8000 222.4500 ;
	    RECT 1194.6000 221.4000 1195.8000 221.5500 ;
	    RECT 1196.7001 220.8000 1197.0000 222.3000 ;
	    RECT 1199.1000 221.4000 1200.9000 222.6000 ;
	    RECT 1201.8000 222.4500 1203.0000 222.6000 ;
	    RECT 1204.2001 222.4500 1205.4000 222.6000 ;
	    RECT 1201.8000 221.5500 1205.4000 222.4500 ;
	    RECT 1201.8000 221.4000 1203.0000 221.5500 ;
	    RECT 1204.2001 221.4000 1205.4000 221.5500 ;
	    RECT 1209.0000 222.4500 1210.2001 222.6000 ;
	    RECT 1228.2001 222.4500 1229.4000 222.6000 ;
	    RECT 1209.0000 221.5500 1229.4000 222.4500 ;
	    RECT 1209.0000 221.4000 1210.2001 221.5500 ;
	    RECT 1228.2001 221.4000 1229.4000 221.5500 ;
	    RECT 1230.3000 220.8000 1230.6000 222.3000 ;
	    RECT 1232.7001 221.4000 1234.5000 222.6000 ;
	    RECT 1235.4000 222.4500 1236.6000 222.6000 ;
	    RECT 1257.0000 222.4500 1258.2001 222.6000 ;
	    RECT 1235.4000 221.5500 1258.2001 222.4500 ;
	    RECT 1259.7001 222.3000 1262.1000 222.6000 ;
	    RECT 1296.3000 222.3000 1298.7001 222.6000 ;
	    RECT 1259.7001 221.7000 1262.4000 222.3000 ;
	    RECT 1235.4000 221.4000 1236.6000 221.5500 ;
	    RECT 1257.0000 221.4000 1258.2001 221.5500 ;
	    RECT 1194.9000 219.3000 1200.3000 219.9000 ;
	    RECT 1201.8000 219.3000 1202.7001 220.5000 ;
	    RECT 1228.5000 219.3000 1233.9000 219.9000 ;
	    RECT 1235.4000 219.3000 1236.3000 220.5000 ;
	    RECT 1002.6000 219.0000 1008.6000 219.3000 ;
	    RECT 1002.6000 213.3000 1003.8000 219.0000 ;
	    RECT 1005.0000 213.3000 1006.2000 218.1000 ;
	    RECT 1007.4000 213.3000 1008.6000 219.0000 ;
	    RECT 1009.8000 213.3000 1011.0000 219.3000 ;
	    RECT 1029.9000 218.4000 1032.6000 219.3000 ;
	    RECT 1029.9000 213.3000 1031.1000 218.4000 ;
	    RECT 1033.8000 213.3000 1035.0000 219.3000 ;
	    RECT 1057.8000 219.0000 1063.8000 219.3000 ;
	    RECT 1057.8000 213.3000 1059.0000 219.0000 ;
	    RECT 1060.2001 213.3000 1061.4000 218.1000 ;
	    RECT 1062.6000 213.3000 1063.8000 219.0000 ;
	    RECT 1065.0000 213.3000 1066.2001 219.3000 ;
	    RECT 1084.2001 213.3000 1085.4000 219.3000 ;
	    RECT 1086.6000 218.4000 1089.3000 219.3000 ;
	    RECT 1088.1000 213.3000 1089.3000 218.4000 ;
	    RECT 1108.2001 213.3000 1109.4000 219.3000 ;
	    RECT 1110.6000 218.4000 1113.3000 219.3000 ;
	    RECT 1112.1000 213.3000 1113.3000 218.4000 ;
	    RECT 1140.3000 218.4000 1143.0000 219.3000 ;
	    RECT 1140.3000 213.3000 1141.5000 218.4000 ;
	    RECT 1144.2001 213.3000 1145.4000 219.3000 ;
	    RECT 1163.4000 213.3000 1164.6000 219.3000 ;
	    RECT 1165.8000 218.4000 1168.5000 219.3000 ;
	    RECT 1167.3000 213.3000 1168.5000 218.4000 ;
	    RECT 1194.6000 219.0000 1200.6000 219.3000 ;
	    RECT 1170.6000 216.4500 1171.8000 216.6000 ;
	    RECT 1182.6000 216.4500 1183.8000 216.6000 ;
	    RECT 1170.6000 215.5500 1183.8000 216.4500 ;
	    RECT 1170.6000 215.4000 1171.8000 215.5500 ;
	    RECT 1182.6000 215.4000 1183.8000 215.5500 ;
	    RECT 1194.6000 213.3000 1195.8000 219.0000 ;
	    RECT 1197.0000 213.3000 1198.2001 218.1000 ;
	    RECT 1199.4000 213.3000 1200.6000 219.0000 ;
	    RECT 1201.8000 213.3000 1203.0000 219.3000 ;
	    RECT 1228.2001 219.0000 1234.2001 219.3000 ;
	    RECT 1228.2001 213.3000 1229.4000 219.0000 ;
	    RECT 1230.6000 213.3000 1231.8000 218.1000 ;
	    RECT 1233.0000 213.3000 1234.2001 219.0000 ;
	    RECT 1235.4000 213.3000 1236.6000 219.3000 ;
	    RECT 1249.8000 216.4500 1251.0000 216.6000 ;
	    RECT 1257.0000 216.4500 1258.2001 216.6000 ;
	    RECT 1249.8000 215.5500 1258.2001 216.4500 ;
	    RECT 1249.8000 215.4000 1251.0000 215.5500 ;
	    RECT 1257.0000 215.4000 1258.2001 215.5500 ;
	    RECT 1261.2001 213.3000 1262.4000 221.7000 ;
	    RECT 1266.6000 213.3000 1267.8000 222.3000 ;
	    RECT 1278.6000 219.4500 1279.8000 219.6000 ;
	    RECT 1288.2001 219.4500 1289.4000 219.6000 ;
	    RECT 1278.6000 218.5500 1289.4000 219.4500 ;
	    RECT 1278.6000 218.4000 1279.8000 218.5500 ;
	    RECT 1288.2001 218.4000 1289.4000 218.5500 ;
	    RECT 1283.4000 216.4500 1284.6000 216.6000 ;
	    RECT 1288.2001 216.4500 1289.4000 216.6000 ;
	    RECT 1283.4000 215.5500 1289.4000 216.4500 ;
	    RECT 1283.4000 215.4000 1284.6000 215.5500 ;
	    RECT 1288.2001 215.4000 1289.4000 215.5500 ;
	    RECT 1290.6000 213.3000 1291.8000 222.3000 ;
	    RECT 1296.0000 221.7000 1298.7001 222.3000 ;
	    RECT 1300.2001 222.4500 1301.4000 222.6000 ;
	    RECT 1309.8000 222.4500 1311.0000 222.6000 ;
	    RECT 1333.8000 222.4500 1335.0000 222.6000 ;
	    RECT 1296.0000 213.3000 1297.2001 221.7000 ;
	    RECT 1300.2001 221.5500 1335.0000 222.4500 ;
	    RECT 1336.5000 222.3000 1338.9000 222.6000 ;
	    RECT 1382.7001 222.3000 1385.1000 222.6000 ;
	    RECT 1336.5000 221.7000 1339.2001 222.3000 ;
	    RECT 1300.2001 221.4000 1301.4000 221.5500 ;
	    RECT 1309.8000 221.4000 1311.0000 221.5500 ;
	    RECT 1333.8000 221.4000 1335.0000 221.5500 ;
	    RECT 1309.8000 213.3000 1311.0000 220.5000 ;
	    RECT 1312.2001 218.4000 1313.4000 219.6000 ;
	    RECT 1312.2001 217.2000 1313.4000 217.5000 ;
	    RECT 1312.2001 213.3000 1313.4000 216.3000 ;
	    RECT 1338.0000 213.3000 1339.2001 221.7000 ;
	    RECT 1343.4000 213.3000 1344.6000 222.3000 ;
	    RECT 1377.0000 213.3000 1378.2001 222.3000 ;
	    RECT 1382.4000 221.7000 1385.1000 222.3000 ;
	    RECT 1386.6000 222.4500 1387.8000 222.6000 ;
	    RECT 1408.2001 222.4500 1409.4000 222.6000 ;
	    RECT 1382.4000 213.3000 1383.6000 221.7000 ;
	    RECT 1386.6000 221.5500 1409.4000 222.4500 ;
	    RECT 1386.6000 221.4000 1387.8000 221.5500 ;
	    RECT 1408.2001 221.4000 1409.4000 221.5500 ;
	    RECT 1410.3000 221.4000 1412.1000 222.6000 ;
	    RECT 1414.2001 220.8000 1414.5000 222.3000 ;
	    RECT 1415.4000 221.4000 1416.6000 222.6000 ;
	    RECT 1432.2001 222.4500 1433.4000 222.6000 ;
	    RECT 1444.2001 222.4500 1445.4000 222.6000 ;
	    RECT 1432.2001 221.5500 1445.4000 222.4500 ;
	    RECT 1432.2001 221.4000 1433.4000 221.5500 ;
	    RECT 1444.2001 221.4000 1445.4000 221.5500 ;
	    RECT 1446.6000 221.4000 1447.8000 222.6000 ;
	    RECT 1478.7001 222.3000 1481.1000 222.6000 ;
	    RECT 1408.5000 219.3000 1409.4000 220.5000 ;
	    RECT 1410.9000 219.3000 1416.3000 219.9000 ;
	    RECT 1408.2001 213.3000 1409.4000 219.3000 ;
	    RECT 1410.6000 219.0000 1416.6000 219.3000 ;
	    RECT 1410.6000 213.3000 1411.8000 219.0000 ;
	    RECT 1413.0000 213.3000 1414.2001 218.1000 ;
	    RECT 1415.4000 213.3000 1416.6000 219.0000 ;
	    RECT 1429.8000 218.4000 1431.0000 219.6000 ;
	    RECT 1429.8000 217.2000 1431.0000 217.5000 ;
	    RECT 1429.8000 213.3000 1431.0000 216.3000 ;
	    RECT 1432.2001 213.3000 1433.4000 220.5000 ;
	    RECT 1446.6000 213.3000 1447.8000 220.5000 ;
	    RECT 1449.0000 218.4000 1450.2001 219.6000 ;
	    RECT 1449.0000 217.2000 1450.2001 217.5000 ;
	    RECT 1449.0000 213.3000 1450.2001 216.3000 ;
	    RECT 1473.0000 213.3000 1474.2001 222.3000 ;
	    RECT 1478.4000 221.7000 1481.1000 222.3000 ;
	    RECT 1506.9000 222.6000 1507.8000 226.5000 ;
	    RECT 1513.8000 226.2000 1515.0000 226.5000 ;
	    RECT 1510.2001 224.4000 1510.5000 225.6000 ;
	    RECT 1511.4000 224.4000 1512.6000 225.6000 ;
	    RECT 1540.5000 222.6000 1541.4000 226.5000 ;
	    RECT 1547.4000 226.2000 1548.6000 226.5000 ;
	    RECT 1543.8000 224.4000 1544.1000 225.6000 ;
	    RECT 1545.0000 224.4000 1546.2001 225.6000 ;
	    RECT 1559.4000 223.5000 1560.6000 239.7000 ;
	    RECT 1561.8000 233.7000 1563.0000 239.7000 ;
	    RECT 1506.9000 222.3000 1509.3000 222.6000 ;
	    RECT 1540.5000 222.3000 1542.9000 222.6000 ;
	    RECT 1506.9000 221.7000 1509.6000 222.3000 ;
	    RECT 1478.4000 213.3000 1479.6000 221.7000 ;
	    RECT 1508.4000 213.3000 1509.6000 221.7000 ;
	    RECT 1513.8000 213.3000 1515.0000 222.3000 ;
	    RECT 1540.5000 221.7000 1543.2001 222.3000 ;
	    RECT 1542.0000 213.3000 1543.2001 221.7000 ;
	    RECT 1547.4000 213.3000 1548.6000 222.3000 ;
	    RECT 1559.4000 221.4000 1560.6000 222.6000 ;
	    RECT 1559.4000 213.3000 1560.6000 220.5000 ;
	    RECT 1561.8000 218.4000 1563.0000 219.6000 ;
	    RECT 1561.8000 217.2000 1563.0000 217.5000 ;
	    RECT 1561.8000 213.3000 1563.0000 216.3000 ;
	    RECT 1.2000 210.6000 1569.0000 212.4000 ;
	    RECT 19.5000 204.6000 20.7000 209.7000 ;
	    RECT 19.5000 203.7000 22.2000 204.6000 ;
	    RECT 23.4000 203.7000 24.6000 209.7000 ;
	    RECT 47.4000 203.7000 48.6000 209.7000 ;
	    RECT 49.8000 204.0000 51.0000 209.7000 ;
	    RECT 52.2000 204.9000 53.4000 209.7000 ;
	    RECT 54.6000 204.0000 55.8000 209.7000 ;
	    RECT 49.8000 203.7000 55.8000 204.0000 ;
	    RECT 21.0000 199.5000 22.2000 203.7000 ;
	    RECT 23.4000 202.5000 24.6000 202.8000 ;
	    RECT 47.7000 202.5000 48.6000 203.7000 ;
	    RECT 50.1000 203.1000 55.5000 203.7000 ;
	    RECT 69.0000 202.5000 70.2000 209.7000 ;
	    RECT 71.4000 206.7000 72.6000 209.7000 ;
	    RECT 71.4000 205.5000 72.6000 205.8000 ;
	    RECT 71.4000 204.4500 72.6000 204.6000 ;
	    RECT 73.8000 204.4500 75.0000 204.6000 ;
	    RECT 71.4000 203.5500 75.0000 204.4500 ;
	    RECT 95.4000 203.7000 96.6000 209.7000 ;
	    RECT 97.8000 204.0000 99.0000 209.7000 ;
	    RECT 100.2000 204.9000 101.4000 209.7000 ;
	    RECT 102.6000 204.0000 103.8000 209.7000 ;
	    RECT 97.8000 203.7000 103.8000 204.0000 ;
	    RECT 71.4000 203.4000 72.6000 203.5500 ;
	    RECT 73.8000 203.4000 75.0000 203.5500 ;
	    RECT 95.7000 202.5000 96.6000 203.7000 ;
	    RECT 98.1000 203.1000 103.5000 203.7000 ;
	    RECT 117.0000 202.5000 118.2000 209.7000 ;
	    RECT 119.4000 206.7000 120.6000 209.7000 ;
	    RECT 119.4000 205.5000 120.6000 205.8000 ;
	    RECT 119.4000 204.4500 120.6000 204.6000 ;
	    RECT 131.4000 204.4500 132.6000 204.6000 ;
	    RECT 136.2000 204.4500 137.4000 204.6000 ;
	    RECT 119.4000 203.5500 137.4000 204.4500 ;
	    RECT 138.6000 203.7000 139.8000 209.7000 ;
	    RECT 142.5000 204.6000 143.7000 209.7000 ;
	    RECT 141.0000 203.7000 143.7000 204.6000 ;
	    RECT 162.6000 203.7000 163.8000 209.7000 ;
	    RECT 166.5000 204.6000 167.7000 209.7000 ;
	    RECT 165.0000 203.7000 167.7000 204.6000 ;
	    RECT 119.4000 203.4000 120.6000 203.5500 ;
	    RECT 131.4000 203.4000 132.6000 203.5500 ;
	    RECT 136.2000 203.4000 137.4000 203.5500 ;
	    RECT 138.6000 202.5000 139.8000 202.8000 ;
	    RECT 23.4000 201.4500 24.6000 201.6000 ;
	    RECT 25.8000 201.4500 27.0000 201.6000 ;
	    RECT 23.4000 200.5500 27.0000 201.4500 ;
	    RECT 23.4000 200.4000 24.6000 200.5500 ;
	    RECT 25.8000 200.4000 27.0000 200.5500 ;
	    RECT 47.4000 200.4000 48.6000 201.6000 ;
	    RECT 49.5000 200.4000 51.3000 201.6000 ;
	    RECT 53.4000 200.7000 53.7000 202.2000 ;
	    RECT 54.6000 200.4000 55.8000 201.6000 ;
	    RECT 69.0000 201.4500 70.2000 201.6000 ;
	    RECT 57.1500 200.5500 70.2000 201.4500 ;
	    RECT 21.0000 198.4500 22.2000 198.6000 ;
	    RECT 40.2000 198.4500 41.4000 198.6000 ;
	    RECT 21.0000 197.5500 41.4000 198.4500 ;
	    RECT 21.0000 197.4000 22.2000 197.5500 ;
	    RECT 40.2000 197.4000 41.4000 197.5500 ;
	    RECT 18.6000 194.4000 19.8000 195.6000 ;
	    RECT 18.6000 193.2000 19.8000 193.5000 ;
	    RECT 18.6000 183.3000 19.8000 189.3000 ;
	    RECT 21.0000 183.3000 22.2000 196.5000 ;
	    RECT 45.0000 195.4500 46.2000 195.6000 ;
	    RECT 47.4000 195.4500 48.6000 195.6000 ;
	    RECT 45.0000 194.5500 48.6000 195.4500 ;
	    RECT 45.0000 194.4000 46.2000 194.5500 ;
	    RECT 47.4000 194.4000 48.6000 194.5500 ;
	    RECT 50.4000 195.3000 51.3000 200.4000 ;
	    RECT 52.2000 199.5000 53.4000 199.8000 ;
	    RECT 52.2000 198.4500 53.4000 198.6000 ;
	    RECT 57.1500 198.4500 58.0500 200.5500 ;
	    RECT 69.0000 200.4000 70.2000 200.5500 ;
	    RECT 93.0000 201.4500 94.2000 201.6000 ;
	    RECT 95.4000 201.4500 96.6000 201.6000 ;
	    RECT 93.0000 200.5500 96.6000 201.4500 ;
	    RECT 93.0000 200.4000 94.2000 200.5500 ;
	    RECT 95.4000 200.4000 96.6000 200.5500 ;
	    RECT 97.5000 200.4000 99.3000 201.6000 ;
	    RECT 101.4000 200.7000 101.7000 202.2000 ;
	    RECT 102.6000 200.4000 103.8000 201.6000 ;
	    RECT 117.0000 201.4500 118.2000 201.6000 ;
	    RECT 105.1500 200.5500 118.2000 201.4500 ;
	    RECT 52.2000 197.5500 58.0500 198.4500 ;
	    RECT 52.2000 197.4000 53.4000 197.5500 ;
	    RECT 50.4000 194.4000 51.9000 195.3000 ;
	    RECT 48.6000 192.6000 49.5000 193.5000 ;
	    RECT 48.6000 191.4000 49.8000 192.6000 ;
	    RECT 23.4000 183.3000 24.6000 189.3000 ;
	    RECT 48.3000 183.3000 49.5000 189.3000 ;
	    RECT 50.7000 183.3000 51.9000 194.4000 ;
	    RECT 54.6000 183.3000 55.8000 195.3000 ;
	    RECT 69.0000 183.3000 70.2000 199.5000 ;
	    RECT 95.4000 194.4000 96.6000 195.6000 ;
	    RECT 98.4000 195.3000 99.3000 200.4000 ;
	    RECT 100.2000 199.5000 101.4000 199.8000 ;
	    RECT 100.2000 198.4500 101.4000 198.6000 ;
	    RECT 105.1500 198.4500 106.0500 200.5500 ;
	    RECT 117.0000 200.4000 118.2000 200.5500 ;
	    RECT 124.2000 201.4500 125.4000 201.6000 ;
	    RECT 138.6000 201.4500 139.8000 201.6000 ;
	    RECT 124.2000 200.5500 139.8000 201.4500 ;
	    RECT 124.2000 200.4000 125.4000 200.5500 ;
	    RECT 138.6000 200.4000 139.8000 200.5500 ;
	    RECT 141.0000 199.5000 142.2000 203.7000 ;
	    RECT 162.6000 202.5000 163.8000 202.8000 ;
	    RECT 162.6000 200.4000 163.8000 201.6000 ;
	    RECT 165.0000 199.5000 166.2000 203.7000 ;
	    RECT 299.4000 200.7000 300.6000 209.7000 ;
	    RECT 304.2000 203.7000 305.4000 209.7000 ;
	    RECT 309.0000 204.9000 310.2000 209.7000 ;
	    RECT 311.4000 205.5000 312.6000 209.7000 ;
	    RECT 313.8000 205.5000 315.0000 209.7000 ;
	    RECT 316.2000 205.5000 317.4000 209.7000 ;
	    RECT 318.6000 206.7000 319.8000 209.7000 ;
	    RECT 321.0000 205.5000 322.2000 209.7000 ;
	    RECT 323.4000 206.7000 324.6000 209.7000 ;
	    RECT 325.8000 205.5000 327.0000 209.7000 ;
	    RECT 328.2000 205.5000 329.4000 209.7000 ;
	    RECT 330.6000 205.5000 331.8000 209.7000 ;
	    RECT 333.0000 205.5000 334.2000 209.7000 ;
	    RECT 306.3000 203.7000 310.2000 204.9000 ;
	    RECT 335.4000 204.9000 336.6000 209.7000 ;
	    RECT 315.3000 203.7000 322.2000 204.6000 ;
	    RECT 306.3000 202.8000 307.5000 203.7000 ;
	    RECT 303.0000 201.6000 307.5000 202.8000 ;
	    RECT 299.4000 199.5000 312.6000 200.7000 ;
	    RECT 315.3000 200.1000 316.5000 203.7000 ;
	    RECT 321.0000 203.4000 322.2000 203.7000 ;
	    RECT 323.4000 203.4000 324.6000 204.6000 ;
	    RECT 325.5000 203.4000 325.8000 204.6000 ;
	    RECT 330.3000 203.4000 331.8000 204.6000 ;
	    RECT 335.4000 203.7000 339.0000 204.9000 ;
	    RECT 340.2000 203.7000 341.4000 209.7000 ;
	    RECT 318.6000 202.5000 319.8000 202.8000 ;
	    RECT 321.0000 202.2000 322.2000 202.5000 ;
	    RECT 318.6000 200.4000 319.8000 201.6000 ;
	    RECT 321.0000 201.3000 327.6000 202.2000 ;
	    RECT 326.4000 201.0000 327.6000 201.3000 ;
	    RECT 100.2000 197.5500 106.0500 198.4500 ;
	    RECT 100.2000 197.4000 101.4000 197.5500 ;
	    RECT 98.4000 194.4000 99.9000 195.3000 ;
	    RECT 96.6000 192.6000 97.5000 193.5000 ;
	    RECT 96.6000 191.4000 97.8000 192.6000 ;
	    RECT 71.4000 183.3000 72.6000 189.3000 ;
	    RECT 96.3000 183.3000 97.5000 189.3000 ;
	    RECT 98.7000 183.3000 99.9000 194.4000 ;
	    RECT 102.6000 183.3000 103.8000 195.3000 ;
	    RECT 117.0000 183.3000 118.2000 199.5000 ;
	    RECT 119.4000 198.4500 120.6000 198.6000 ;
	    RECT 141.0000 198.4500 142.2000 198.6000 ;
	    RECT 119.4000 197.5500 142.2000 198.4500 ;
	    RECT 119.4000 197.4000 120.6000 197.5500 ;
	    RECT 141.0000 197.4000 142.2000 197.5500 ;
	    RECT 165.0000 198.4500 166.2000 198.6000 ;
	    RECT 205.8000 198.4500 207.0000 198.6000 ;
	    RECT 165.0000 197.5500 207.0000 198.4500 ;
	    RECT 165.0000 197.4000 166.2000 197.5500 ;
	    RECT 205.8000 197.4000 207.0000 197.5500 ;
	    RECT 119.4000 183.3000 120.6000 189.3000 ;
	    RECT 138.6000 183.3000 139.8000 189.3000 ;
	    RECT 141.0000 183.3000 142.2000 196.5000 ;
	    RECT 143.4000 195.4500 144.6000 195.6000 ;
	    RECT 153.0000 195.4500 154.2000 195.6000 ;
	    RECT 143.4000 194.5500 154.2000 195.4500 ;
	    RECT 143.4000 194.4000 144.6000 194.5500 ;
	    RECT 153.0000 194.4000 154.2000 194.5500 ;
	    RECT 143.4000 193.2000 144.6000 193.5000 ;
	    RECT 143.4000 183.3000 144.6000 189.3000 ;
	    RECT 162.6000 183.3000 163.8000 189.3000 ;
	    RECT 165.0000 183.3000 166.2000 196.5000 ;
	    RECT 167.4000 195.4500 168.6000 195.6000 ;
	    RECT 169.8000 195.4500 171.0000 195.6000 ;
	    RECT 220.2000 195.4500 221.4000 195.6000 ;
	    RECT 167.4000 194.5500 221.4000 195.4500 ;
	    RECT 167.4000 194.4000 168.6000 194.5500 ;
	    RECT 169.8000 194.4000 171.0000 194.5500 ;
	    RECT 220.2000 194.4000 221.4000 194.5500 ;
	    RECT 167.4000 193.2000 168.6000 193.5000 ;
	    RECT 299.4000 191.1000 300.6000 199.5000 ;
	    RECT 313.5000 198.9000 316.5000 200.1000 ;
	    RECT 322.2000 198.9000 327.0000 200.1000 ;
	    RECT 330.6000 199.2000 331.8000 203.4000 ;
	    RECT 337.8000 202.8000 339.0000 203.7000 ;
	    RECT 337.8000 201.9000 340.5000 202.8000 ;
	    RECT 339.3000 200.1000 340.5000 201.9000 ;
	    RECT 345.0000 201.9000 346.2000 209.7000 ;
	    RECT 347.4000 204.0000 348.6000 209.7000 ;
	    RECT 349.8000 206.7000 351.0000 209.7000 ;
	    RECT 364.2000 206.7000 365.4000 209.7000 ;
	    RECT 364.2000 205.5000 365.4000 205.8000 ;
	    RECT 347.4000 202.8000 348.9000 204.0000 ;
	    RECT 364.2000 203.4000 365.4000 204.6000 ;
	    RECT 345.0000 201.0000 346.8000 201.9000 ;
	    RECT 339.3000 198.9000 345.0000 200.1000 ;
	    RECT 301.5000 198.0000 302.7000 198.3000 ;
	    RECT 301.5000 197.1000 308.1000 198.0000 ;
	    RECT 309.0000 197.4000 310.2000 198.6000 ;
	    RECT 335.4000 198.0000 336.6000 198.9000 ;
	    RECT 345.9000 198.0000 346.8000 201.0000 ;
	    RECT 311.1000 197.1000 336.6000 198.0000 ;
	    RECT 345.6000 197.1000 346.8000 198.0000 ;
	    RECT 343.5000 196.2000 344.7000 196.5000 ;
	    RECT 304.2000 194.4000 305.4000 195.6000 ;
	    RECT 306.3000 195.3000 344.7000 196.2000 ;
	    RECT 309.3000 195.0000 310.5000 195.3000 ;
	    RECT 345.6000 194.4000 346.5000 197.1000 ;
	    RECT 347.7000 196.2000 348.9000 202.8000 ;
	    RECT 366.6000 202.5000 367.8000 209.7000 ;
	    RECT 381.0000 206.7000 382.2000 209.7000 ;
	    RECT 381.0000 205.5000 382.2000 205.8000 ;
	    RECT 381.0000 203.4000 382.2000 204.6000 ;
	    RECT 383.4000 202.5000 384.6000 209.7000 ;
	    RECT 397.8000 206.7000 399.0000 209.7000 ;
	    RECT 397.8000 205.5000 399.0000 205.8000 ;
	    RECT 397.8000 203.4000 399.0000 204.6000 ;
	    RECT 400.2000 202.5000 401.4000 209.7000 ;
	    RECT 532.2000 206.7000 533.4000 209.7000 ;
	    RECT 534.6000 204.0000 535.8000 209.7000 ;
	    RECT 534.3000 202.8000 535.8000 204.0000 ;
	    RECT 366.6000 201.4500 367.8000 201.6000 ;
	    RECT 381.0000 201.4500 382.2000 201.6000 ;
	    RECT 366.6000 200.5500 382.2000 201.4500 ;
	    RECT 366.6000 200.4000 367.8000 200.5500 ;
	    RECT 381.0000 200.4000 382.2000 200.5500 ;
	    RECT 383.4000 201.4500 384.6000 201.6000 ;
	    RECT 395.4000 201.4500 396.6000 201.6000 ;
	    RECT 383.4000 200.5500 396.6000 201.4500 ;
	    RECT 383.4000 200.4000 384.6000 200.5500 ;
	    RECT 395.4000 200.4000 396.6000 200.5500 ;
	    RECT 400.2000 201.4500 401.4000 201.6000 ;
	    RECT 529.8000 201.4500 531.0000 201.6000 ;
	    RECT 400.2000 200.5500 531.0000 201.4500 ;
	    RECT 400.2000 200.4000 401.4000 200.5500 ;
	    RECT 529.8000 200.4000 531.0000 200.5500 ;
	    RECT 313.8000 194.1000 315.0000 194.4000 ;
	    RECT 306.9000 193.5000 315.0000 194.1000 ;
	    RECT 305.7000 193.2000 315.0000 193.5000 ;
	    RECT 316.5000 193.5000 329.4000 194.4000 ;
	    RECT 301.8000 192.0000 304.2000 193.2000 ;
	    RECT 305.7000 192.3000 307.8000 193.2000 ;
	    RECT 316.5000 192.3000 317.4000 193.5000 ;
	    RECT 328.2000 193.2000 329.4000 193.5000 ;
	    RECT 333.0000 193.5000 346.5000 194.4000 ;
	    RECT 347.4000 195.0000 348.9000 196.2000 ;
	    RECT 347.4000 193.5000 348.6000 195.0000 ;
	    RECT 333.0000 193.2000 334.2000 193.5000 ;
	    RECT 303.3000 191.4000 304.2000 192.0000 ;
	    RECT 308.7000 191.4000 317.4000 192.3000 ;
	    RECT 318.3000 191.4000 322.2000 192.6000 ;
	    RECT 299.4000 190.2000 302.4000 191.1000 ;
	    RECT 303.3000 190.2000 309.6000 191.4000 ;
	    RECT 301.5000 189.3000 302.4000 190.2000 ;
	    RECT 167.4000 183.3000 168.6000 189.3000 ;
	    RECT 299.4000 183.3000 300.6000 189.3000 ;
	    RECT 301.5000 188.4000 303.0000 189.3000 ;
	    RECT 301.8000 183.3000 303.0000 188.4000 ;
	    RECT 304.2000 182.4000 305.4000 189.3000 ;
	    RECT 306.6000 183.3000 307.8000 190.2000 ;
	    RECT 309.0000 183.3000 310.2000 189.3000 ;
	    RECT 311.4000 183.3000 312.6000 187.5000 ;
	    RECT 313.8000 183.3000 315.0000 187.5000 ;
	    RECT 316.2000 183.3000 317.4000 190.5000 ;
	    RECT 318.6000 183.3000 319.8000 189.3000 ;
	    RECT 321.0000 183.3000 322.2000 190.5000 ;
	    RECT 323.4000 183.3000 324.6000 189.3000 ;
	    RECT 325.8000 183.3000 327.0000 192.6000 ;
	    RECT 337.8000 191.4000 341.7000 192.6000 ;
	    RECT 330.6000 190.2000 336.9000 191.4000 ;
	    RECT 328.2000 183.3000 329.4000 187.5000 ;
	    RECT 330.6000 183.3000 331.8000 187.5000 ;
	    RECT 333.0000 183.3000 334.2000 187.5000 ;
	    RECT 335.4000 183.3000 336.6000 189.3000 ;
	    RECT 337.8000 183.3000 339.0000 191.4000 ;
	    RECT 345.6000 191.1000 346.5000 193.5000 ;
	    RECT 347.4000 191.4000 348.6000 192.6000 ;
	    RECT 342.6000 190.2000 346.5000 191.1000 ;
	    RECT 340.2000 183.3000 341.4000 189.3000 ;
	    RECT 342.6000 183.3000 343.8000 190.2000 ;
	    RECT 345.0000 183.3000 346.2000 189.3000 ;
	    RECT 347.4000 183.3000 348.6000 190.5000 ;
	    RECT 349.8000 183.3000 351.0000 189.3000 ;
	    RECT 364.2000 183.3000 365.4000 189.3000 ;
	    RECT 366.6000 183.3000 367.8000 199.5000 ;
	    RECT 381.0000 183.3000 382.2000 189.3000 ;
	    RECT 383.4000 183.3000 384.6000 199.5000 ;
	    RECT 397.8000 183.3000 399.0000 189.3000 ;
	    RECT 400.2000 183.3000 401.4000 199.5000 ;
	    RECT 534.3000 196.2000 535.5000 202.8000 ;
	    RECT 537.0000 201.9000 538.2000 209.7000 ;
	    RECT 541.8000 203.7000 543.0000 209.7000 ;
	    RECT 546.6000 204.9000 547.8000 209.7000 ;
	    RECT 549.0000 205.5000 550.2000 209.7000 ;
	    RECT 551.4000 205.5000 552.6000 209.7000 ;
	    RECT 553.8000 205.5000 555.0000 209.7000 ;
	    RECT 556.2000 205.5000 557.4000 209.7000 ;
	    RECT 558.6000 206.7000 559.8000 209.7000 ;
	    RECT 561.0000 205.5000 562.2000 209.7000 ;
	    RECT 563.4000 206.7000 564.6000 209.7000 ;
	    RECT 565.8000 205.5000 567.0000 209.7000 ;
	    RECT 568.2000 205.5000 569.4000 209.7000 ;
	    RECT 570.6000 205.5000 571.8000 209.7000 ;
	    RECT 544.2000 203.7000 547.8000 204.9000 ;
	    RECT 573.0000 204.9000 574.2000 209.7000 ;
	    RECT 544.2000 202.8000 545.4000 203.7000 ;
	    RECT 536.4000 201.0000 538.2000 201.9000 ;
	    RECT 542.7000 201.9000 545.4000 202.8000 ;
	    RECT 551.4000 203.4000 552.9000 204.6000 ;
	    RECT 557.4000 203.4000 557.7000 204.6000 ;
	    RECT 558.6000 203.4000 559.8000 204.6000 ;
	    RECT 561.0000 203.7000 567.9000 204.6000 ;
	    RECT 573.0000 203.7000 576.9000 204.9000 ;
	    RECT 577.8000 203.7000 579.0000 209.7000 ;
	    RECT 561.0000 203.4000 562.2000 203.7000 ;
	    RECT 536.4000 198.0000 537.3000 201.0000 ;
	    RECT 542.7000 200.1000 543.9000 201.9000 ;
	    RECT 538.2000 198.9000 543.9000 200.1000 ;
	    RECT 551.4000 199.2000 552.6000 203.4000 ;
	    RECT 563.4000 202.5000 564.6000 202.8000 ;
	    RECT 561.0000 202.2000 562.2000 202.5000 ;
	    RECT 555.6000 201.3000 562.2000 202.2000 ;
	    RECT 555.6000 201.0000 556.8000 201.3000 ;
	    RECT 563.4000 200.4000 564.6000 201.6000 ;
	    RECT 566.7000 200.1000 567.9000 203.7000 ;
	    RECT 575.7000 202.8000 576.9000 203.7000 ;
	    RECT 575.7000 201.6000 580.2000 202.8000 ;
	    RECT 582.6000 200.7000 583.8000 209.7000 ;
	    RECT 606.6000 200.7000 607.8000 209.7000 ;
	    RECT 612.0000 201.3000 613.2000 209.7000 ;
	    RECT 633.0000 206.7000 634.2000 209.7000 ;
	    RECT 635.4000 206.7000 636.6000 209.7000 ;
	    RECT 637.8000 206.7000 639.0000 209.7000 ;
	    RECT 649.8000 206.7000 651.0000 209.7000 ;
	    RECT 633.0000 205.5000 634.2000 205.8000 ;
	    RECT 628.2000 204.4500 629.4000 204.6000 ;
	    RECT 633.0000 204.4500 634.2000 204.6000 ;
	    RECT 628.2000 203.5500 634.2000 204.4500 ;
	    RECT 628.2000 203.4000 629.4000 203.5500 ;
	    RECT 633.0000 203.4000 634.2000 203.5500 ;
	    RECT 635.7000 202.5000 636.6000 206.7000 ;
	    RECT 649.8000 205.5000 651.0000 205.8000 ;
	    RECT 637.8000 204.4500 639.0000 204.6000 ;
	    RECT 649.8000 204.4500 651.0000 204.6000 ;
	    RECT 637.8000 203.5500 651.0000 204.4500 ;
	    RECT 637.8000 203.4000 639.0000 203.5500 ;
	    RECT 649.8000 203.4000 651.0000 203.5500 ;
	    RECT 652.2000 202.5000 653.4000 209.7000 ;
	    RECT 684.3000 203.7000 685.5000 209.7000 ;
	    RECT 688.2000 203.7000 689.4000 209.7000 ;
	    RECT 690.6000 206.7000 691.8000 209.7000 ;
	    RECT 690.3000 205.5000 691.5000 205.8000 ;
	    RECT 690.6000 204.4500 691.8000 204.6000 ;
	    RECT 695.4000 204.4500 696.6000 204.6000 ;
	    RECT 635.4000 201.4500 636.6000 201.6000 ;
	    RECT 649.8000 201.4500 651.0000 201.6000 ;
	    RECT 612.0000 200.7000 614.7000 201.3000 ;
	    RECT 556.2000 198.9000 561.0000 200.1000 ;
	    RECT 566.7000 198.9000 569.7000 200.1000 ;
	    RECT 570.6000 199.5000 583.8000 200.7000 ;
	    RECT 612.3000 200.4000 614.7000 200.7000 ;
	    RECT 635.4000 200.5500 651.0000 201.4500 ;
	    RECT 635.4000 200.4000 636.6000 200.5500 ;
	    RECT 649.8000 200.4000 651.0000 200.5500 ;
	    RECT 652.2000 201.4500 653.4000 201.6000 ;
	    RECT 683.4000 201.4500 684.6000 201.6000 ;
	    RECT 652.2000 200.5500 684.6000 201.4500 ;
	    RECT 652.2000 200.4000 653.4000 200.5500 ;
	    RECT 683.4000 200.4000 684.6000 200.5500 ;
	    RECT 685.8000 200.4000 687.0000 201.6000 ;
	    RECT 546.6000 198.0000 547.8000 198.9000 ;
	    RECT 536.4000 197.1000 537.6000 198.0000 ;
	    RECT 546.6000 197.1000 572.1000 198.0000 ;
	    RECT 573.0000 197.4000 574.2000 198.6000 ;
	    RECT 580.5000 198.0000 581.7000 198.3000 ;
	    RECT 575.1000 197.1000 581.7000 198.0000 ;
	    RECT 534.3000 195.0000 535.8000 196.2000 ;
	    RECT 534.6000 193.5000 535.8000 195.0000 ;
	    RECT 536.7000 194.4000 537.6000 197.1000 ;
	    RECT 538.5000 196.2000 539.7000 196.5000 ;
	    RECT 538.5000 195.3000 576.9000 196.2000 ;
	    RECT 572.7000 195.0000 573.9000 195.3000 ;
	    RECT 577.8000 194.4000 579.0000 195.6000 ;
	    RECT 536.7000 193.5000 550.2000 194.4000 ;
	    RECT 484.2000 192.4500 485.4000 192.6000 ;
	    RECT 534.6000 192.4500 535.8000 192.6000 ;
	    RECT 484.2000 191.5500 535.8000 192.4500 ;
	    RECT 484.2000 191.4000 485.4000 191.5500 ;
	    RECT 534.6000 191.4000 535.8000 191.5500 ;
	    RECT 536.7000 191.1000 537.6000 193.5000 ;
	    RECT 549.0000 193.2000 550.2000 193.5000 ;
	    RECT 553.8000 193.5000 566.7000 194.4000 ;
	    RECT 553.8000 193.2000 555.0000 193.5000 ;
	    RECT 541.5000 191.4000 545.4000 192.6000 ;
	    RECT 532.2000 183.3000 533.4000 189.3000 ;
	    RECT 534.6000 183.3000 535.8000 190.5000 ;
	    RECT 536.7000 190.2000 540.6000 191.1000 ;
	    RECT 537.0000 183.3000 538.2000 189.3000 ;
	    RECT 539.4000 183.3000 540.6000 190.2000 ;
	    RECT 541.8000 183.3000 543.0000 189.3000 ;
	    RECT 544.2000 183.3000 545.4000 191.4000 ;
	    RECT 546.3000 190.2000 552.6000 191.4000 ;
	    RECT 546.6000 183.3000 547.8000 189.3000 ;
	    RECT 549.0000 183.3000 550.2000 187.5000 ;
	    RECT 551.4000 183.3000 552.6000 187.5000 ;
	    RECT 553.8000 183.3000 555.0000 187.5000 ;
	    RECT 556.2000 183.3000 557.4000 192.6000 ;
	    RECT 561.0000 191.4000 564.9000 192.6000 ;
	    RECT 565.8000 192.3000 566.7000 193.5000 ;
	    RECT 568.2000 194.1000 569.4000 194.4000 ;
	    RECT 568.2000 193.5000 576.3000 194.1000 ;
	    RECT 568.2000 193.2000 577.5000 193.5000 ;
	    RECT 575.4000 192.3000 577.5000 193.2000 ;
	    RECT 565.8000 191.4000 574.5000 192.3000 ;
	    RECT 579.0000 192.0000 581.4000 193.2000 ;
	    RECT 579.0000 191.4000 579.9000 192.0000 ;
	    RECT 558.6000 183.3000 559.8000 189.3000 ;
	    RECT 561.0000 183.3000 562.2000 190.5000 ;
	    RECT 563.4000 183.3000 564.6000 189.3000 ;
	    RECT 565.8000 183.3000 567.0000 190.5000 ;
	    RECT 573.6000 190.2000 579.9000 191.4000 ;
	    RECT 582.6000 191.1000 583.8000 199.5000 ;
	    RECT 609.0000 197.4000 610.2000 198.6000 ;
	    RECT 611.1000 197.4000 611.4000 198.6000 ;
	    RECT 606.6000 196.5000 607.8000 196.8000 ;
	    RECT 613.8000 196.5000 614.7000 200.4000 ;
	    RECT 606.6000 194.4000 607.8000 195.6000 ;
	    RECT 613.8000 195.4500 615.0000 195.6000 ;
	    RECT 628.2000 195.4500 629.4000 195.6000 ;
	    RECT 613.8000 194.5500 629.4000 195.4500 ;
	    RECT 635.7000 195.3000 636.6000 199.5000 ;
	    RECT 637.8000 198.4500 639.0000 198.6000 ;
	    RECT 645.0000 198.4500 646.2000 198.6000 ;
	    RECT 637.8000 197.5500 646.2000 198.4500 ;
	    RECT 637.8000 197.4000 639.0000 197.5500 ;
	    RECT 645.0000 197.4000 646.2000 197.5500 ;
	    RECT 637.8000 196.2000 639.0000 196.5000 ;
	    RECT 613.8000 194.4000 615.0000 194.5500 ;
	    RECT 628.2000 194.4000 629.4000 194.5500 ;
	    RECT 611.4000 193.5000 612.6000 193.8000 ;
	    RECT 604.2000 192.4500 605.4000 192.6000 ;
	    RECT 611.4000 192.4500 612.6000 192.6000 ;
	    RECT 604.2000 191.5500 612.6000 192.4500 ;
	    RECT 604.2000 191.4000 605.4000 191.5500 ;
	    RECT 611.4000 191.4000 612.6000 191.5500 ;
	    RECT 580.8000 190.2000 583.8000 191.1000 ;
	    RECT 613.8000 190.5000 614.7000 193.5000 ;
	    RECT 568.2000 183.3000 569.4000 187.5000 ;
	    RECT 570.6000 183.3000 571.8000 187.5000 ;
	    RECT 573.0000 183.3000 574.2000 189.3000 ;
	    RECT 575.4000 183.3000 576.6000 190.2000 ;
	    RECT 580.8000 189.3000 581.7000 190.2000 ;
	    RECT 609.3000 189.6000 614.7000 190.5000 ;
	    RECT 609.3000 189.3000 610.2000 189.6000 ;
	    RECT 577.8000 182.4000 579.0000 189.3000 ;
	    RECT 580.2000 188.4000 581.7000 189.3000 ;
	    RECT 580.2000 183.3000 581.4000 188.4000 ;
	    RECT 582.6000 183.3000 583.8000 189.3000 ;
	    RECT 606.6000 183.3000 607.8000 189.3000 ;
	    RECT 609.0000 183.3000 610.2000 189.3000 ;
	    RECT 613.8000 189.3000 614.7000 189.6000 ;
	    RECT 611.4000 183.3000 612.6000 188.7000 ;
	    RECT 613.8000 183.3000 615.0000 189.3000 ;
	    RECT 633.0000 183.3000 634.2000 195.3000 ;
	    RECT 635.4000 194.1000 638.1000 195.3000 ;
	    RECT 636.9000 183.3000 638.1000 194.1000 ;
	    RECT 649.8000 183.3000 651.0000 189.3000 ;
	    RECT 652.2000 183.3000 653.4000 199.5000 ;
	    RECT 683.5500 198.6000 684.4500 200.4000 ;
	    RECT 685.8000 199.2000 687.0000 199.5000 ;
	    RECT 683.4000 197.4000 684.6000 198.6000 ;
	    RECT 688.2000 198.3000 689.1000 203.7000 ;
	    RECT 690.6000 203.5500 696.6000 204.4500 ;
	    RECT 690.6000 203.4000 691.8000 203.5500 ;
	    RECT 695.4000 203.4000 696.6000 203.5500 ;
	    RECT 760.2000 203.1000 761.4000 209.7000 ;
	    RECT 762.6000 204.0000 763.8000 209.7000 ;
	    RECT 766.5000 207.6000 768.3000 209.7000 ;
	    RECT 766.5000 206.7000 768.6000 207.6000 ;
	    RECT 771.0000 206.7000 772.2000 209.7000 ;
	    RECT 773.4000 206.7000 774.6000 209.7000 ;
	    RECT 775.8000 206.7000 777.3000 209.7000 ;
	    RECT 780.0000 207.6000 781.2000 209.7000 ;
	    RECT 780.0000 206.7000 783.0000 207.6000 ;
	    RECT 767.4000 205.5000 768.6000 206.7000 ;
	    RECT 773.7000 205.8000 774.6000 206.7000 ;
	    RECT 773.7000 204.9000 777.9000 205.8000 ;
	    RECT 776.7000 204.6000 777.9000 204.9000 ;
	    RECT 779.4000 204.6000 780.6000 205.8000 ;
	    RECT 781.8000 205.5000 783.0000 206.7000 ;
	    RECT 764.7000 203.1000 765.9000 203.4000 ;
	    RECT 760.2000 202.2000 765.9000 203.1000 ;
	    RECT 760.2000 199.5000 761.4000 202.2000 ;
	    RECT 770.7000 201.3000 771.9000 201.6000 ;
	    RECT 779.4000 201.3000 780.3000 204.6000 ;
	    RECT 784.2000 203.7000 785.4000 209.7000 ;
	    RECT 786.6000 202.5000 787.8000 209.7000 ;
	    RECT 793.8000 209.4000 795.0000 210.6000 ;
	    RECT 805.8000 202.5000 807.0000 209.7000 ;
	    RECT 808.2000 203.7000 809.4000 209.7000 ;
	    RECT 810.6000 202.8000 811.8000 209.7000 ;
	    RECT 808.5000 201.9000 811.8000 202.8000 ;
	    RECT 829.8000 202.8000 831.0000 209.7000 ;
	    RECT 832.2000 203.7000 833.4000 209.7000 ;
	    RECT 829.8000 201.9000 833.1000 202.8000 ;
	    RECT 834.6000 202.5000 835.8000 209.7000 ;
	    RECT 853.8000 203.7000 855.0000 209.7000 ;
	    RECT 857.7000 204.6000 858.9000 209.7000 ;
	    RECT 856.2000 203.7000 858.9000 204.6000 ;
	    RECT 885.0000 203.7000 886.2000 209.7000 ;
	    RECT 887.4000 204.0000 888.6000 209.7000 ;
	    RECT 889.8000 204.9000 891.0000 209.7000 ;
	    RECT 892.2000 204.0000 893.4000 209.7000 ;
	    RECT 887.4000 203.7000 893.4000 204.0000 ;
	    RECT 853.8000 202.5000 855.0000 202.8000 ;
	    RECT 770.1000 200.4000 783.3000 201.3000 ;
	    RECT 784.2000 200.4000 785.4000 201.6000 ;
	    RECT 786.3000 200.4000 786.6000 201.6000 ;
	    RECT 805.8000 200.4000 807.0000 201.6000 ;
	    RECT 767.4000 199.2000 768.6000 199.5000 ;
	    RECT 690.6000 198.4500 691.8000 198.6000 ;
	    RECT 757.8000 198.4500 759.0000 198.6000 ;
	    RECT 685.5000 196.8000 685.8000 198.3000 ;
	    RECT 688.2000 197.4000 689.7000 198.3000 ;
	    RECT 690.6000 197.5500 759.0000 198.4500 ;
	    RECT 690.6000 197.4000 691.8000 197.5500 ;
	    RECT 757.8000 197.4000 759.0000 197.5500 ;
	    RECT 760.2000 197.4000 761.4000 198.6000 ;
	    RECT 762.9000 198.3000 768.6000 199.2000 ;
	    RECT 762.9000 198.0000 764.1000 198.3000 ;
	    RECT 765.3000 197.1000 766.5000 197.4000 ;
	    RECT 762.3000 196.5000 766.5000 197.1000 ;
	    RECT 690.6000 195.3000 691.5000 196.5000 ;
	    RECT 760.2000 196.2000 766.5000 196.5000 ;
	    RECT 683.4000 194.4000 689.4000 195.3000 ;
	    RECT 683.4000 183.3000 684.6000 194.4000 ;
	    RECT 685.8000 183.3000 687.0000 193.5000 ;
	    RECT 688.2000 183.3000 689.4000 194.4000 ;
	    RECT 690.6000 183.3000 691.8000 195.3000 ;
	    RECT 760.2000 183.3000 761.4000 196.2000 ;
	    RECT 770.1000 195.6000 771.0000 200.4000 ;
	    RECT 780.9000 200.1000 782.1000 200.4000 ;
	    RECT 783.3000 198.6000 784.5000 198.9000 ;
	    RECT 777.0000 197.4000 778.2000 198.6000 ;
	    RECT 779.1000 197.7000 784.5000 198.6000 ;
	    RECT 805.8000 198.6000 807.0000 199.5000 ;
	    RECT 779.4000 196.5000 787.8000 196.8000 ;
	    RECT 779.1000 196.2000 787.8000 196.5000 ;
	    RECT 762.6000 183.3000 763.8000 195.3000 ;
	    RECT 767.4000 194.7000 771.0000 195.6000 ;
	    RECT 773.1000 195.9000 787.8000 196.2000 ;
	    RECT 773.1000 195.3000 780.3000 195.9000 ;
	    RECT 767.4000 193.2000 768.3000 194.7000 ;
	    RECT 766.2000 192.0000 768.3000 193.2000 ;
	    RECT 770.7000 193.5000 771.9000 193.8000 ;
	    RECT 773.1000 193.5000 774.0000 195.3000 ;
	    RECT 770.7000 192.6000 774.0000 193.5000 ;
	    RECT 774.9000 193.5000 783.0000 194.4000 ;
	    RECT 774.9000 193.2000 776.1000 193.5000 ;
	    RECT 781.8000 193.2000 783.0000 193.5000 ;
	    RECT 772.5000 191.1000 773.7000 191.4000 ;
	    RECT 776.7000 191.1000 777.9000 191.4000 ;
	    RECT 767.4000 189.3000 768.6000 190.5000 ;
	    RECT 772.5000 190.2000 777.9000 191.1000 ;
	    RECT 773.7000 189.3000 774.6000 190.2000 ;
	    RECT 781.8000 189.3000 783.0000 190.5000 ;
	    RECT 766.5000 183.3000 768.3000 189.3000 ;
	    RECT 771.0000 183.3000 772.2000 189.3000 ;
	    RECT 773.4000 183.3000 774.6000 189.3000 ;
	    RECT 775.8000 183.3000 777.0000 189.3000 ;
	    RECT 780.0000 188.4000 783.0000 189.3000 ;
	    RECT 780.0000 183.3000 781.2000 188.4000 ;
	    RECT 784.2000 183.3000 785.4000 195.0000 ;
	    RECT 786.6000 183.3000 787.8000 195.9000 ;
	    RECT 805.8000 195.3000 806.7000 198.6000 ;
	    RECT 808.5000 197.4000 809.4000 201.9000 ;
	    RECT 810.6000 199.5000 811.8000 199.8000 ;
	    RECT 829.8000 199.5000 831.0000 199.8000 ;
	    RECT 810.6000 197.4000 811.8000 198.6000 ;
	    RECT 829.8000 197.4000 831.0000 198.6000 ;
	    RECT 832.2000 197.4000 833.1000 201.9000 ;
	    RECT 834.6000 200.4000 835.8000 201.6000 ;
	    RECT 853.8000 200.4000 855.0000 201.6000 ;
	    RECT 856.2000 199.5000 857.4000 203.7000 ;
	    RECT 885.3000 202.5000 886.2000 203.7000 ;
	    RECT 887.7000 203.1000 893.1000 203.7000 ;
	    RECT 911.4000 202.5000 912.6000 209.7000 ;
	    RECT 913.8000 206.7000 915.0000 209.7000 ;
	    RECT 913.8000 205.5000 915.0000 205.8000 ;
	    RECT 913.8000 204.4500 915.0000 204.6000 ;
	    RECT 930.6000 204.4500 931.8000 204.6000 ;
	    RECT 913.8000 203.5500 931.8000 204.4500 ;
	    RECT 933.0000 203.7000 934.2000 209.7000 ;
	    RECT 936.9000 204.6000 938.1000 209.7000 ;
	    RECT 940.2000 209.4000 941.4000 210.6000 ;
	    RECT 962.7000 205.2000 963.9000 209.7000 ;
	    RECT 935.4000 203.7000 938.1000 204.6000 ;
	    RECT 961.8000 203.7000 963.9000 205.2000 ;
	    RECT 965.1000 204.0000 966.3000 209.7000 ;
	    RECT 969.0000 203.7000 970.2000 209.7000 ;
	    RECT 995.4000 204.0000 996.6000 209.7000 ;
	    RECT 997.8000 204.9000 999.0000 209.7000 ;
	    RECT 1000.2000 204.0000 1001.4000 209.7000 ;
	    RECT 995.4000 203.7000 1001.4000 204.0000 ;
	    RECT 1002.6000 203.7000 1003.8000 209.7000 ;
	    RECT 1014.6000 206.7000 1015.8000 209.7000 ;
	    RECT 1014.6000 205.5000 1015.8000 205.8000 ;
	    RECT 913.8000 203.4000 915.0000 203.5500 ;
	    RECT 930.6000 203.4000 931.8000 203.5500 ;
	    RECT 933.0000 202.5000 934.2000 202.8000 ;
	    RECT 882.6000 201.4500 883.8000 201.6000 ;
	    RECT 885.0000 201.4500 886.2000 201.6000 ;
	    RECT 882.6000 200.5500 886.2000 201.4500 ;
	    RECT 882.6000 200.4000 883.8000 200.5500 ;
	    RECT 885.0000 200.4000 886.2000 200.5500 ;
	    RECT 887.1000 200.4000 888.9000 201.6000 ;
	    RECT 891.0000 200.7000 891.3000 202.2000 ;
	    RECT 892.2000 201.4500 893.4000 201.6000 ;
	    RECT 909.0000 201.4500 910.2000 201.6000 ;
	    RECT 892.2000 200.5500 910.2000 201.4500 ;
	    RECT 892.2000 200.4000 893.4000 200.5500 ;
	    RECT 909.0000 200.4000 910.2000 200.5500 ;
	    RECT 911.4000 200.4000 912.6000 201.6000 ;
	    RECT 921.0000 201.4500 922.2000 201.6000 ;
	    RECT 933.0000 201.4500 934.2000 201.6000 ;
	    RECT 921.0000 200.5500 934.2000 201.4500 ;
	    RECT 921.0000 200.4000 922.2000 200.5500 ;
	    RECT 933.0000 200.4000 934.2000 200.5500 ;
	    RECT 834.6000 198.6000 835.8000 199.5000 ;
	    RECT 807.6000 196.2000 809.4000 197.4000 ;
	    RECT 808.5000 195.3000 809.4000 196.2000 ;
	    RECT 832.2000 196.2000 834.0000 197.4000 ;
	    RECT 832.2000 195.3000 833.1000 196.2000 ;
	    RECT 834.9000 195.3000 835.8000 198.6000 ;
	    RECT 856.2000 197.4000 857.4000 198.6000 ;
	    RECT 805.8000 183.3000 807.0000 195.3000 ;
	    RECT 808.5000 194.4000 811.8000 195.3000 ;
	    RECT 808.2000 183.3000 809.4000 193.5000 ;
	    RECT 810.6000 183.3000 811.8000 194.4000 ;
	    RECT 829.8000 194.4000 833.1000 195.3000 ;
	    RECT 829.8000 183.3000 831.0000 194.4000 ;
	    RECT 832.2000 183.3000 833.4000 193.5000 ;
	    RECT 834.6000 183.3000 835.8000 195.3000 ;
	    RECT 853.8000 183.3000 855.0000 189.3000 ;
	    RECT 856.2000 183.3000 857.4000 196.5000 ;
	    RECT 858.6000 194.4000 859.8000 195.6000 ;
	    RECT 885.0000 194.4000 886.2000 195.6000 ;
	    RECT 888.0000 195.3000 888.9000 200.4000 ;
	    RECT 889.8000 199.5000 891.0000 199.8000 ;
	    RECT 935.4000 199.5000 936.6000 203.7000 ;
	    RECT 961.8000 199.5000 962.7000 203.7000 ;
	    RECT 969.0000 203.4000 969.9000 203.7000 ;
	    RECT 967.2000 202.8000 969.9000 203.4000 ;
	    RECT 995.7000 203.1000 1001.1000 203.7000 ;
	    RECT 963.6000 202.5000 969.9000 202.8000 ;
	    RECT 1002.6000 202.5000 1003.5000 203.7000 ;
	    RECT 1014.6000 203.4000 1015.8000 204.6000 ;
	    RECT 1017.0000 202.5000 1018.2000 209.7000 ;
	    RECT 963.6000 201.9000 968.1000 202.5000 ;
	    RECT 963.6000 201.6000 964.8000 201.9000 ;
	    RECT 889.8000 197.4000 891.0000 198.6000 ;
	    RECT 888.0000 194.4000 889.5000 195.3000 ;
	    RECT 858.6000 193.2000 859.8000 193.5000 ;
	    RECT 886.2000 192.6000 887.1000 193.5000 ;
	    RECT 886.2000 191.4000 887.4000 192.6000 ;
	    RECT 858.6000 183.3000 859.8000 189.3000 ;
	    RECT 885.9000 183.3000 887.1000 189.3000 ;
	    RECT 888.3000 183.3000 889.5000 194.4000 ;
	    RECT 892.2000 183.3000 893.4000 195.3000 ;
	    RECT 911.4000 183.3000 912.6000 199.5000 ;
	    RECT 935.4000 198.4500 936.6000 198.6000 ;
	    RECT 959.4000 198.4500 960.6000 198.6000 ;
	    RECT 935.4000 197.5500 960.6000 198.4500 ;
	    RECT 935.4000 197.4000 936.6000 197.5500 ;
	    RECT 959.4000 197.4000 960.6000 197.5500 ;
	    RECT 961.8000 197.4000 963.0000 198.6000 ;
	    RECT 963.9000 196.5000 964.8000 201.6000 ;
	    RECT 966.0000 200.7000 967.2000 201.0000 ;
	    RECT 966.0000 199.8000 967.5000 200.7000 ;
	    RECT 969.0000 200.4000 970.2000 201.6000 ;
	    RECT 995.4000 200.4000 996.6000 201.6000 ;
	    RECT 997.5000 200.7000 997.8000 202.2000 ;
	    RECT 999.9000 200.4000 1001.7000 201.6000 ;
	    RECT 1002.6000 201.4500 1003.8000 201.6000 ;
	    RECT 1014.6000 201.4500 1015.8000 201.6000 ;
	    RECT 1002.6000 200.5500 1015.8000 201.4500 ;
	    RECT 1002.6000 200.4000 1003.8000 200.5500 ;
	    RECT 1014.6000 200.4000 1015.8000 200.5500 ;
	    RECT 1017.0000 201.4500 1018.2000 201.6000 ;
	    RECT 1041.0000 201.4500 1042.2001 201.6000 ;
	    RECT 1017.0000 200.5500 1042.2001 201.4500 ;
	    RECT 1043.4000 200.7000 1044.6000 209.7000 ;
	    RECT 1048.8000 201.3000 1050.0000 209.7000 ;
	    RECT 1048.8000 200.7000 1051.5000 201.3000 ;
	    RECT 1074.6000 200.7000 1075.8000 209.7000 ;
	    RECT 1080.0000 201.3000 1081.2001 209.7000 ;
	    RECT 1080.0000 200.7000 1082.7001 201.3000 ;
	    RECT 1105.8000 200.7000 1107.0000 209.7000 ;
	    RECT 1111.2001 201.3000 1112.4000 209.7000 ;
	    RECT 1134.6000 206.7000 1135.8000 209.7000 ;
	    RECT 1134.6000 205.5000 1135.8000 205.8000 ;
	    RECT 1134.6000 203.4000 1135.8000 204.6000 ;
	    RECT 1137.0000 202.5000 1138.2001 209.7000 ;
	    RECT 1141.8000 204.4500 1143.0000 204.6000 ;
	    RECT 1158.6000 204.4500 1159.8000 204.6000 ;
	    RECT 1141.8000 203.5500 1159.8000 204.4500 ;
	    RECT 1161.0000 203.7000 1162.2001 209.7000 ;
	    RECT 1163.4000 204.0000 1164.6000 209.7000 ;
	    RECT 1165.8000 204.9000 1167.0000 209.7000 ;
	    RECT 1168.2001 204.0000 1169.4000 209.7000 ;
	    RECT 1163.4000 203.7000 1169.4000 204.0000 ;
	    RECT 1141.8000 203.4000 1143.0000 203.5500 ;
	    RECT 1158.6000 203.4000 1159.8000 203.5500 ;
	    RECT 1161.3000 202.5000 1162.2001 203.7000 ;
	    RECT 1163.7001 203.1000 1169.1000 203.7000 ;
	    RECT 1180.2001 202.5000 1181.4000 209.7000 ;
	    RECT 1182.6000 206.7000 1183.8000 209.7000 ;
	    RECT 1182.6000 205.5000 1183.8000 205.8000 ;
	    RECT 1182.6000 204.4500 1183.8000 204.6000 ;
	    RECT 1185.0000 204.4500 1186.2001 204.6000 ;
	    RECT 1182.6000 203.5500 1186.2001 204.4500 ;
	    RECT 1209.0000 204.0000 1210.2001 209.7000 ;
	    RECT 1211.4000 204.9000 1212.6000 209.7000 ;
	    RECT 1213.8000 204.0000 1215.0000 209.7000 ;
	    RECT 1209.0000 203.7000 1215.0000 204.0000 ;
	    RECT 1216.2001 203.7000 1217.4000 209.7000 ;
	    RECT 1182.6000 203.4000 1183.8000 203.5500 ;
	    RECT 1185.0000 203.4000 1186.2001 203.5500 ;
	    RECT 1209.3000 203.1000 1214.7001 203.7000 ;
	    RECT 1216.2001 202.5000 1217.1000 203.7000 ;
	    RECT 1230.6000 202.5000 1231.8000 209.7000 ;
	    RECT 1233.0000 206.7000 1234.2001 209.7000 ;
	    RECT 1233.0000 205.5000 1234.2001 205.8000 ;
	    RECT 1253.1000 204.6000 1254.3000 209.7000 ;
	    RECT 1233.0000 203.4000 1234.2001 204.6000 ;
	    RECT 1253.1000 203.7000 1255.8000 204.6000 ;
	    RECT 1257.0000 203.7000 1258.2001 209.7000 ;
	    RECT 1281.0000 203.7000 1282.2001 209.7000 ;
	    RECT 1283.4000 204.0000 1284.6000 209.7000 ;
	    RECT 1285.8000 204.9000 1287.0000 209.7000 ;
	    RECT 1288.2001 204.0000 1289.4000 209.7000 ;
	    RECT 1283.4000 203.7000 1289.4000 204.0000 ;
	    RECT 1308.3000 204.6000 1309.5000 209.7000 ;
	    RECT 1308.3000 203.7000 1311.0000 204.6000 ;
	    RECT 1312.2001 203.7000 1313.4000 209.7000 ;
	    RECT 1360.2001 203.7000 1361.4000 209.7000 ;
	    RECT 1362.6000 204.6000 1364.1000 209.7000 ;
	    RECT 1366.8000 204.3000 1369.2001 209.7000 ;
	    RECT 1371.9000 204.6000 1373.4000 209.7000 ;
	    RECT 1137.0000 201.4500 1138.2001 201.6000 ;
	    RECT 1158.6000 201.4500 1159.8000 201.6000 ;
	    RECT 1111.2001 200.7000 1113.9000 201.3000 ;
	    RECT 1017.0000 200.4000 1018.2000 200.5500 ;
	    RECT 1041.0000 200.4000 1042.2001 200.5500 ;
	    RECT 1049.1000 200.4000 1051.5000 200.7000 ;
	    RECT 1080.3000 200.4000 1082.7001 200.7000 ;
	    RECT 1111.5000 200.4000 1113.9000 200.7000 ;
	    RECT 1137.0000 200.5500 1159.8000 201.4500 ;
	    RECT 1137.0000 200.4000 1138.2001 200.5500 ;
	    RECT 1158.6000 200.4000 1159.8000 200.5500 ;
	    RECT 1161.0000 200.4000 1162.2001 201.6000 ;
	    RECT 1163.1000 200.4000 1164.9000 201.6000 ;
	    RECT 1167.0000 200.7000 1167.3000 202.2000 ;
	    RECT 1168.2001 200.4000 1169.4000 201.6000 ;
	    RECT 1180.2001 201.4500 1181.4000 201.6000 ;
	    RECT 1170.7500 200.5500 1207.6500 201.4500 ;
	    RECT 966.6000 199.5000 967.5000 199.8000 ;
	    RECT 997.8000 199.5000 999.0000 199.8000 ;
	    RECT 969.0000 199.2000 970.2000 199.5000 ;
	    RECT 966.6000 197.4000 967.8000 198.6000 ;
	    RECT 997.8000 197.4000 999.0000 198.6000 ;
	    RECT 913.8000 183.3000 915.0000 189.3000 ;
	    RECT 933.0000 183.3000 934.2000 189.3000 ;
	    RECT 935.4000 183.3000 936.6000 196.5000 ;
	    RECT 937.8000 195.4500 939.0000 195.6000 ;
	    RECT 940.2000 195.4500 941.4000 195.6000 ;
	    RECT 937.8000 194.5500 941.4000 195.4500 ;
	    RECT 937.8000 194.4000 939.0000 194.5500 ;
	    RECT 940.2000 194.4000 941.4000 194.5500 ;
	    RECT 961.8000 195.3000 962.7000 196.5000 ;
	    RECT 963.9000 195.6000 967.5000 196.5000 ;
	    RECT 937.8000 193.2000 939.0000 193.5000 ;
	    RECT 940.2000 192.4500 941.4000 192.6000 ;
	    RECT 942.6000 192.4500 943.8000 192.6000 ;
	    RECT 954.6000 192.4500 955.8000 192.6000 ;
	    RECT 940.2000 191.5500 955.8000 192.4500 ;
	    RECT 940.2000 191.4000 941.4000 191.5500 ;
	    RECT 942.6000 191.4000 943.8000 191.5500 ;
	    RECT 954.6000 191.4000 955.8000 191.5500 ;
	    RECT 937.8000 183.3000 939.0000 189.3000 ;
	    RECT 961.8000 183.3000 963.0000 195.3000 ;
	    RECT 964.2000 183.3000 965.4000 194.7000 ;
	    RECT 966.6000 189.3000 967.5000 195.6000 ;
	    RECT 999.9000 195.3000 1000.8000 200.4000 ;
	    RECT 966.6000 183.3000 967.8000 189.3000 ;
	    RECT 969.0000 183.3000 970.2000 189.3000 ;
	    RECT 995.4000 183.3000 996.6000 195.3000 ;
	    RECT 999.3000 194.4000 1000.8000 195.3000 ;
	    RECT 1002.6000 194.4000 1003.8000 195.6000 ;
	    RECT 999.3000 183.3000 1000.5000 194.4000 ;
	    RECT 1001.7000 192.6000 1002.6000 193.5000 ;
	    RECT 1001.4000 191.4000 1002.6000 192.6000 ;
	    RECT 1001.7000 183.3000 1002.9000 189.3000 ;
	    RECT 1014.6000 183.3000 1015.8000 189.3000 ;
	    RECT 1017.0000 183.3000 1018.2000 199.5000 ;
	    RECT 1045.8000 197.4000 1047.0000 198.6000 ;
	    RECT 1047.9000 197.4000 1048.2001 198.6000 ;
	    RECT 1043.4000 196.5000 1044.6000 196.8000 ;
	    RECT 1050.6000 196.5000 1051.5000 200.4000 ;
	    RECT 1077.0000 197.4000 1078.2001 198.6000 ;
	    RECT 1079.1000 197.4000 1079.4000 198.6000 ;
	    RECT 1074.6000 196.5000 1075.8000 196.8000 ;
	    RECT 1081.8000 196.5000 1082.7001 200.4000 ;
	    RECT 1108.2001 197.4000 1109.4000 198.6000 ;
	    RECT 1110.3000 197.4000 1110.6000 198.6000 ;
	    RECT 1105.8000 196.5000 1107.0000 196.8000 ;
	    RECT 1113.0000 196.5000 1113.9000 200.4000 ;
	    RECT 1041.0000 195.4500 1042.2001 195.6000 ;
	    RECT 1043.4000 195.4500 1044.6000 195.6000 ;
	    RECT 1041.0000 194.5500 1044.6000 195.4500 ;
	    RECT 1041.0000 194.4000 1042.2001 194.5500 ;
	    RECT 1043.4000 194.4000 1044.6000 194.5500 ;
	    RECT 1050.6000 195.4500 1051.8000 195.6000 ;
	    RECT 1074.6000 195.4500 1075.8000 195.6000 ;
	    RECT 1077.0000 195.4500 1078.2001 195.6000 ;
	    RECT 1050.6000 194.5500 1078.2001 195.4500 ;
	    RECT 1050.6000 194.4000 1051.8000 194.5500 ;
	    RECT 1074.6000 194.4000 1075.8000 194.5500 ;
	    RECT 1077.0000 194.4000 1078.2001 194.5500 ;
	    RECT 1081.8000 195.4500 1083.0000 195.6000 ;
	    RECT 1093.8000 195.4500 1095.0000 195.6000 ;
	    RECT 1081.8000 194.5500 1095.0000 195.4500 ;
	    RECT 1081.8000 194.4000 1083.0000 194.5500 ;
	    RECT 1093.8000 194.4000 1095.0000 194.5500 ;
	    RECT 1105.8000 194.4000 1107.0000 195.6000 ;
	    RECT 1113.0000 195.4500 1114.2001 195.6000 ;
	    RECT 1134.6000 195.4500 1135.8000 195.6000 ;
	    RECT 1113.0000 194.5500 1135.8000 195.4500 ;
	    RECT 1113.0000 194.4000 1114.2001 194.5500 ;
	    RECT 1134.6000 194.4000 1135.8000 194.5500 ;
	    RECT 1048.2001 193.5000 1049.4000 193.8000 ;
	    RECT 1079.4000 193.5000 1080.6000 193.8000 ;
	    RECT 1110.6000 193.5000 1111.8000 193.8000 ;
	    RECT 1048.2001 191.4000 1049.4000 192.6000 ;
	    RECT 1050.6000 190.5000 1051.5000 193.5000 ;
	    RECT 1079.4000 191.4000 1080.6000 192.6000 ;
	    RECT 1081.8000 190.5000 1082.7001 193.5000 ;
	    RECT 1110.6000 191.4000 1111.8000 192.6000 ;
	    RECT 1113.0000 190.5000 1113.9000 193.5000 ;
	    RECT 1046.1000 189.6000 1051.5000 190.5000 ;
	    RECT 1046.1000 189.3000 1047.0000 189.6000 ;
	    RECT 1043.4000 183.3000 1044.6000 189.3000 ;
	    RECT 1045.8000 183.3000 1047.0000 189.3000 ;
	    RECT 1050.6000 189.3000 1051.5000 189.6000 ;
	    RECT 1077.3000 189.6000 1082.7001 190.5000 ;
	    RECT 1077.3000 189.3000 1078.2001 189.6000 ;
	    RECT 1048.2001 183.3000 1049.4000 188.7000 ;
	    RECT 1050.6000 183.3000 1051.8000 189.3000 ;
	    RECT 1074.6000 183.3000 1075.8000 189.3000 ;
	    RECT 1077.0000 183.3000 1078.2001 189.3000 ;
	    RECT 1081.8000 189.3000 1082.7001 189.6000 ;
	    RECT 1108.5000 189.6000 1113.9000 190.5000 ;
	    RECT 1108.5000 189.3000 1109.4000 189.6000 ;
	    RECT 1079.4000 183.3000 1080.6000 188.7000 ;
	    RECT 1081.8000 183.3000 1083.0000 189.3000 ;
	    RECT 1105.8000 183.3000 1107.0000 189.3000 ;
	    RECT 1108.2001 183.3000 1109.4000 189.3000 ;
	    RECT 1113.0000 189.3000 1113.9000 189.6000 ;
	    RECT 1110.6000 183.3000 1111.8000 188.7000 ;
	    RECT 1113.0000 183.3000 1114.2001 189.3000 ;
	    RECT 1134.6000 183.3000 1135.8000 189.3000 ;
	    RECT 1137.0000 183.3000 1138.2001 199.5000 ;
	    RECT 1156.2001 195.4500 1157.4000 195.6000 ;
	    RECT 1161.0000 195.4500 1162.2001 195.6000 ;
	    RECT 1156.2001 194.5500 1162.2001 195.4500 ;
	    RECT 1156.2001 194.4000 1157.4000 194.5500 ;
	    RECT 1161.0000 194.4000 1162.2001 194.5500 ;
	    RECT 1164.0000 195.3000 1164.9000 200.4000 ;
	    RECT 1165.8000 199.5000 1167.0000 199.8000 ;
	    RECT 1165.8000 198.4500 1167.0000 198.6000 ;
	    RECT 1170.7500 198.4500 1171.6500 200.5500 ;
	    RECT 1180.2001 200.4000 1181.4000 200.5500 ;
	    RECT 1165.8000 197.5500 1171.6500 198.4500 ;
	    RECT 1165.8000 197.4000 1167.0000 197.5500 ;
	    RECT 1164.0000 194.4000 1165.5000 195.3000 ;
	    RECT 1162.2001 192.6000 1163.1000 193.5000 ;
	    RECT 1162.2001 191.4000 1163.4000 192.6000 ;
	    RECT 1146.6000 186.4500 1147.8000 186.6000 ;
	    RECT 1158.6000 186.4500 1159.8000 186.6000 ;
	    RECT 1146.6000 185.5500 1159.8000 186.4500 ;
	    RECT 1146.6000 185.4000 1147.8000 185.5500 ;
	    RECT 1158.6000 185.4000 1159.8000 185.5500 ;
	    RECT 1161.9000 183.3000 1163.1000 189.3000 ;
	    RECT 1164.3000 183.3000 1165.5000 194.4000 ;
	    RECT 1168.2001 183.3000 1169.4000 195.3000 ;
	    RECT 1180.2001 183.3000 1181.4000 199.5000 ;
	    RECT 1206.7500 198.4500 1207.6500 200.5500 ;
	    RECT 1209.0000 200.4000 1210.2001 201.6000 ;
	    RECT 1211.1000 200.7000 1211.4000 202.2000 ;
	    RECT 1213.5000 200.4000 1215.3000 201.6000 ;
	    RECT 1216.2001 201.4500 1217.4000 201.6000 ;
	    RECT 1221.0000 201.4500 1222.2001 201.6000 ;
	    RECT 1216.2001 200.5500 1222.2001 201.4500 ;
	    RECT 1216.2001 200.4000 1217.4000 200.5500 ;
	    RECT 1221.0000 200.4000 1222.2001 200.5500 ;
	    RECT 1230.6000 201.4500 1231.8000 201.6000 ;
	    RECT 1237.8000 201.4500 1239.0000 201.6000 ;
	    RECT 1230.6000 200.5500 1239.0000 201.4500 ;
	    RECT 1230.6000 200.4000 1231.8000 200.5500 ;
	    RECT 1237.8000 200.4000 1239.0000 200.5500 ;
	    RECT 1211.4000 199.5000 1212.6000 199.8000 ;
	    RECT 1211.4000 198.4500 1212.6000 198.6000 ;
	    RECT 1206.7500 197.5500 1212.6000 198.4500 ;
	    RECT 1211.4000 197.4000 1212.6000 197.5500 ;
	    RECT 1213.5000 195.3000 1214.4000 200.4000 ;
	    RECT 1254.6000 199.5000 1255.8000 203.7000 ;
	    RECT 1257.0000 202.5000 1258.2001 202.8000 ;
	    RECT 1281.3000 202.5000 1282.2001 203.7000 ;
	    RECT 1283.7001 203.1000 1289.1000 203.7000 ;
	    RECT 1257.0000 200.4000 1258.2001 201.6000 ;
	    RECT 1264.2001 201.4500 1265.4000 201.6000 ;
	    RECT 1278.6000 201.4500 1279.8000 201.6000 ;
	    RECT 1281.0000 201.4500 1282.2001 201.6000 ;
	    RECT 1264.2001 200.5500 1282.2001 201.4500 ;
	    RECT 1264.2001 200.4000 1265.4000 200.5500 ;
	    RECT 1278.6000 200.4000 1279.8000 200.5500 ;
	    RECT 1281.0000 200.4000 1282.2001 200.5500 ;
	    RECT 1283.1000 200.4000 1284.9000 201.6000 ;
	    RECT 1287.0000 200.7000 1287.3000 202.2000 ;
	    RECT 1288.2001 200.4000 1289.4000 201.6000 ;
	    RECT 1182.6000 183.3000 1183.8000 189.3000 ;
	    RECT 1209.0000 183.3000 1210.2001 195.3000 ;
	    RECT 1212.9000 194.4000 1214.4000 195.3000 ;
	    RECT 1216.2001 194.4000 1217.4000 195.6000 ;
	    RECT 1212.9000 183.3000 1214.1000 194.4000 ;
	    RECT 1215.3000 192.6000 1216.2001 193.5000 ;
	    RECT 1215.0000 191.4000 1216.2001 192.6000 ;
	    RECT 1215.3000 183.3000 1216.5000 189.3000 ;
	    RECT 1230.6000 183.3000 1231.8000 199.5000 ;
	    RECT 1254.6000 198.4500 1255.8000 198.6000 ;
	    RECT 1276.2001 198.4500 1277.4000 198.6000 ;
	    RECT 1254.6000 197.5500 1277.4000 198.4500 ;
	    RECT 1254.6000 197.4000 1255.8000 197.5500 ;
	    RECT 1276.2001 197.4000 1277.4000 197.5500 ;
	    RECT 1252.2001 194.4000 1253.4000 195.6000 ;
	    RECT 1252.2001 193.2000 1253.4000 193.5000 ;
	    RECT 1233.0000 183.3000 1234.2001 189.3000 ;
	    RECT 1252.2001 183.3000 1253.4000 189.3000 ;
	    RECT 1254.6000 183.3000 1255.8000 196.5000 ;
	    RECT 1281.0000 194.4000 1282.2001 195.6000 ;
	    RECT 1284.0000 195.3000 1284.9000 200.4000 ;
	    RECT 1285.8000 199.5000 1287.0000 199.8000 ;
	    RECT 1309.8000 199.5000 1311.0000 203.7000 ;
	    RECT 1360.2001 202.8000 1363.5000 203.7000 ;
	    RECT 1365.0000 203.1000 1367.4000 203.4000 ;
	    RECT 1312.2001 202.5000 1313.4000 202.8000 ;
	    RECT 1362.3000 202.5000 1363.5000 202.8000 ;
	    RECT 1364.4000 202.2000 1367.4000 203.1000 ;
	    RECT 1364.4000 201.6000 1365.3000 202.2000 ;
	    RECT 1312.2001 200.4000 1313.4000 201.6000 ;
	    RECT 1348.2001 201.4500 1349.4000 201.6000 ;
	    RECT 1360.2001 201.4500 1361.4000 201.6000 ;
	    RECT 1348.2001 200.5500 1361.4000 201.4500 ;
	    RECT 1348.2001 200.4000 1349.4000 200.5500 ;
	    RECT 1360.2001 200.4000 1361.4000 200.5500 ;
	    RECT 1362.3000 200.7000 1365.3000 201.6000 ;
	    RECT 1362.3000 200.4000 1362.6000 200.7000 ;
	    RECT 1366.2001 200.1000 1367.4000 201.3000 ;
	    RECT 1366.2001 199.2000 1367.1000 200.1000 ;
	    RECT 1285.8000 198.4500 1287.0000 198.6000 ;
	    RECT 1295.4000 198.4500 1296.6000 198.6000 ;
	    RECT 1285.8000 197.5500 1296.6000 198.4500 ;
	    RECT 1285.8000 197.4000 1287.0000 197.5500 ;
	    RECT 1295.4000 197.4000 1296.6000 197.5500 ;
	    RECT 1309.8000 198.4500 1311.0000 198.6000 ;
	    RECT 1360.2001 198.4500 1361.4000 198.6000 ;
	    RECT 1309.8000 197.5500 1361.4000 198.4500 ;
	    RECT 1363.2001 198.3000 1367.1000 199.2000 ;
	    RECT 1368.3000 199.5000 1369.2001 204.3000 ;
	    RECT 1374.6000 203.7000 1375.8000 209.7000 ;
	    RECT 1370.1000 202.2000 1371.3000 203.4000 ;
	    RECT 1372.2001 202.8000 1375.8000 203.7000 ;
	    RECT 1372.2001 202.5000 1373.4000 202.8000 ;
	    RECT 1370.4000 201.6000 1371.3000 202.2000 ;
	    RECT 1370.4000 200.4000 1371.6000 201.6000 ;
	    RECT 1373.4000 200.4000 1373.7001 201.6000 ;
	    RECT 1374.6000 200.4000 1375.8000 201.6000 ;
	    RECT 1398.6000 200.7000 1399.8000 209.7000 ;
	    RECT 1404.0000 201.3000 1405.2001 209.7000 ;
	    RECT 1420.2001 206.7000 1421.4000 209.7000 ;
	    RECT 1420.2001 205.5000 1421.4000 205.8000 ;
	    RECT 1408.2001 204.4500 1409.4000 204.6000 ;
	    RECT 1420.2001 204.4500 1421.4000 204.6000 ;
	    RECT 1408.2001 203.5500 1421.4000 204.4500 ;
	    RECT 1408.2001 203.4000 1409.4000 203.5500 ;
	    RECT 1420.2001 203.4000 1421.4000 203.5500 ;
	    RECT 1422.6000 202.5000 1423.8000 209.7000 ;
	    RECT 1422.6000 201.4500 1423.8000 201.6000 ;
	    RECT 1444.2001 201.4500 1445.4000 201.6000 ;
	    RECT 1404.0000 200.7000 1406.7001 201.3000 ;
	    RECT 1404.3000 200.4000 1406.7001 200.7000 ;
	    RECT 1422.6000 200.5500 1445.4000 201.4500 ;
	    RECT 1448.4000 201.3000 1449.6000 209.7000 ;
	    RECT 1422.6000 200.4000 1423.8000 200.5500 ;
	    RECT 1444.2001 200.4000 1445.4000 200.5500 ;
	    RECT 1446.9000 200.7000 1449.6000 201.3000 ;
	    RECT 1453.8000 200.7000 1455.0000 209.7000 ;
	    RECT 1477.8000 200.7000 1479.0000 209.7000 ;
	    RECT 1483.2001 201.3000 1484.4000 209.7000 ;
	    RECT 1510.8000 201.3000 1512.0000 209.7000 ;
	    RECT 1483.2001 200.7000 1485.9000 201.3000 ;
	    RECT 1446.9000 200.4000 1449.3000 200.7000 ;
	    RECT 1483.5000 200.4000 1485.9000 200.7000 ;
	    RECT 1368.3000 198.3000 1368.9000 199.5000 ;
	    RECT 1369.8000 198.4500 1371.0000 198.6000 ;
	    RECT 1363.2001 198.0000 1364.4000 198.3000 ;
	    RECT 1309.8000 197.4000 1311.0000 197.5500 ;
	    RECT 1360.2001 197.4000 1361.4000 197.5500 ;
	    RECT 1369.8000 197.5500 1397.2500 198.4500 ;
	    RECT 1369.8000 197.4000 1371.0000 197.5500 ;
	    RECT 1366.5000 197.1000 1367.7001 197.4000 ;
	    RECT 1302.6000 195.4500 1303.8000 195.6000 ;
	    RECT 1307.4000 195.4500 1308.6000 195.6000 ;
	    RECT 1284.0000 194.4000 1285.5000 195.3000 ;
	    RECT 1282.2001 192.6000 1283.1000 193.5000 ;
	    RECT 1282.2001 191.4000 1283.4000 192.6000 ;
	    RECT 1257.0000 183.3000 1258.2001 189.3000 ;
	    RECT 1281.9000 183.3000 1283.1000 189.3000 ;
	    RECT 1284.3000 183.3000 1285.5000 194.4000 ;
	    RECT 1288.2001 183.3000 1289.4000 195.3000 ;
	    RECT 1302.6000 194.5500 1308.6000 195.4500 ;
	    RECT 1302.6000 194.4000 1303.8000 194.5500 ;
	    RECT 1307.4000 194.4000 1308.6000 194.5500 ;
	    RECT 1307.4000 193.2000 1308.6000 193.5000 ;
	    RECT 1307.4000 183.3000 1308.6000 189.3000 ;
	    RECT 1309.8000 183.3000 1311.0000 196.5000 ;
	    RECT 1362.6000 196.2000 1367.7001 197.1000 ;
	    RECT 1362.6000 195.3000 1363.5000 196.2000 ;
	    RECT 1368.9000 195.3000 1369.8000 196.5000 ;
	    RECT 1396.3500 195.4500 1397.2500 197.5500 ;
	    RECT 1401.0000 197.4000 1402.2001 198.6000 ;
	    RECT 1403.1000 197.4000 1403.4000 198.6000 ;
	    RECT 1398.6000 196.5000 1399.8000 196.8000 ;
	    RECT 1405.8000 196.5000 1406.7001 200.4000 ;
	    RECT 1398.6000 195.4500 1399.8000 195.6000 ;
	    RECT 1360.2001 194.4000 1363.5000 195.3000 ;
	    RECT 1312.2001 183.3000 1313.4000 189.3000 ;
	    RECT 1360.2001 183.3000 1361.4000 194.4000 ;
	    RECT 1362.3000 194.1000 1363.5000 194.4000 ;
	    RECT 1366.8000 194.4000 1369.8000 195.3000 ;
	    RECT 1372.2001 194.4000 1375.8000 195.3000 ;
	    RECT 1396.3500 194.5500 1399.8000 195.4500 ;
	    RECT 1398.6000 194.4000 1399.8000 194.5500 ;
	    RECT 1405.8000 195.4500 1407.0000 195.6000 ;
	    RECT 1417.8000 195.4500 1419.0000 195.6000 ;
	    RECT 1405.8000 194.5500 1419.0000 195.4500 ;
	    RECT 1405.8000 194.4000 1407.0000 194.5500 ;
	    RECT 1417.8000 194.4000 1419.0000 194.5500 ;
	    RECT 1362.6000 183.3000 1364.1000 193.2000 ;
	    RECT 1366.8000 183.3000 1369.2001 194.4000 ;
	    RECT 1372.2001 194.1000 1373.4000 194.4000 ;
	    RECT 1371.9000 183.3000 1373.4000 193.2000 ;
	    RECT 1374.6000 183.3000 1375.8000 194.4000 ;
	    RECT 1403.4000 193.5000 1404.6000 193.8000 ;
	    RECT 1396.2001 192.4500 1397.4000 192.6000 ;
	    RECT 1403.4000 192.4500 1404.6000 192.6000 ;
	    RECT 1396.2001 191.5500 1404.6000 192.4500 ;
	    RECT 1396.2001 191.4000 1397.4000 191.5500 ;
	    RECT 1403.4000 191.4000 1404.6000 191.5500 ;
	    RECT 1405.8000 190.5000 1406.7001 193.5000 ;
	    RECT 1401.3000 189.6000 1406.7001 190.5000 ;
	    RECT 1401.3000 189.3000 1402.2001 189.6000 ;
	    RECT 1398.6000 183.3000 1399.8000 189.3000 ;
	    RECT 1401.0000 183.3000 1402.2001 189.3000 ;
	    RECT 1405.8000 189.3000 1406.7001 189.6000 ;
	    RECT 1403.4000 183.3000 1404.6000 188.7000 ;
	    RECT 1405.8000 183.3000 1407.0000 189.3000 ;
	    RECT 1420.2001 183.3000 1421.4000 189.3000 ;
	    RECT 1422.6000 183.3000 1423.8000 199.5000 ;
	    RECT 1446.9000 196.5000 1447.8000 200.4000 ;
	    RECT 1450.2001 197.4000 1450.5000 198.6000 ;
	    RECT 1451.4000 197.4000 1452.6000 198.6000 ;
	    RECT 1480.2001 197.4000 1481.4000 198.6000 ;
	    RECT 1482.3000 197.4000 1482.6000 198.6000 ;
	    RECT 1453.8000 196.5000 1455.0000 196.8000 ;
	    RECT 1477.8000 196.5000 1479.0000 196.8000 ;
	    RECT 1485.0000 196.5000 1485.9000 200.4000 ;
	    RECT 1509.3000 200.7000 1512.0000 201.3000 ;
	    RECT 1516.2001 200.7000 1517.4000 209.7000 ;
	    RECT 1542.6000 206.7000 1543.8000 209.7000 ;
	    RECT 1542.9000 205.5000 1544.1000 205.8000 ;
	    RECT 1542.6000 203.4000 1543.8000 204.6000 ;
	    RECT 1545.0000 203.7000 1546.2001 209.7000 ;
	    RECT 1548.9000 203.7000 1550.1000 209.7000 ;
	    RECT 1509.3000 200.4000 1511.7001 200.7000 ;
	    RECT 1509.3000 196.5000 1510.2001 200.4000 ;
	    RECT 1512.6000 197.4000 1512.9000 198.6000 ;
	    RECT 1513.8000 197.4000 1515.0000 198.6000 ;
	    RECT 1540.2001 198.4500 1541.4000 198.6000 ;
	    RECT 1542.6000 198.4500 1543.8000 198.6000 ;
	    RECT 1540.2001 197.5500 1543.8000 198.4500 ;
	    RECT 1545.3000 198.3000 1546.2001 203.7000 ;
	    RECT 1547.4000 201.4500 1548.6000 201.6000 ;
	    RECT 1557.0000 201.4500 1558.2001 201.6000 ;
	    RECT 1547.4000 200.5500 1558.2001 201.4500 ;
	    RECT 1547.4000 200.4000 1548.6000 200.5500 ;
	    RECT 1557.0000 200.4000 1558.2001 200.5500 ;
	    RECT 1547.4000 199.2000 1548.6000 199.5000 ;
	    RECT 1549.8000 198.4500 1551.0000 198.6000 ;
	    RECT 1554.6000 198.4500 1555.8000 198.6000 ;
	    RECT 1540.2001 197.4000 1541.4000 197.5500 ;
	    RECT 1542.6000 197.4000 1543.8000 197.5500 ;
	    RECT 1544.7001 197.4000 1546.2001 198.3000 ;
	    RECT 1548.6000 196.8000 1548.9000 198.3000 ;
	    RECT 1549.8000 197.5500 1555.8000 198.4500 ;
	    RECT 1549.8000 197.4000 1551.0000 197.5500 ;
	    RECT 1554.6000 197.4000 1555.8000 197.5500 ;
	    RECT 1516.2001 196.5000 1517.4000 196.8000 ;
	    RECT 1444.2001 195.4500 1445.4000 195.6000 ;
	    RECT 1446.6000 195.4500 1447.8000 195.6000 ;
	    RECT 1444.2001 194.5500 1447.8000 195.4500 ;
	    RECT 1444.2001 194.4000 1445.4000 194.5500 ;
	    RECT 1446.6000 194.4000 1447.8000 194.5500 ;
	    RECT 1453.8000 194.4000 1455.0000 195.6000 ;
	    RECT 1468.2001 195.4500 1469.4000 195.6000 ;
	    RECT 1477.8000 195.4500 1479.0000 195.6000 ;
	    RECT 1468.2001 194.5500 1479.0000 195.4500 ;
	    RECT 1468.2001 194.4000 1469.4000 194.5500 ;
	    RECT 1477.8000 194.4000 1479.0000 194.5500 ;
	    RECT 1485.0000 194.4000 1486.2001 195.6000 ;
	    RECT 1506.6000 195.4500 1507.8000 195.6000 ;
	    RECT 1509.0000 195.4500 1510.2001 195.6000 ;
	    RECT 1506.6000 194.5500 1510.2001 195.4500 ;
	    RECT 1506.6000 194.4000 1507.8000 194.5500 ;
	    RECT 1509.0000 194.4000 1510.2001 194.5500 ;
	    RECT 1516.2001 194.4000 1517.4000 195.6000 ;
	    RECT 1542.9000 195.3000 1543.8000 196.5000 ;
	    RECT 1449.0000 193.5000 1450.2001 193.8000 ;
	    RECT 1482.6000 193.5000 1483.8000 193.8000 ;
	    RECT 1511.4000 193.5000 1512.6000 193.8000 ;
	    RECT 1446.9000 190.5000 1447.8000 193.5000 ;
	    RECT 1449.0000 192.4500 1450.2001 192.6000 ;
	    RECT 1482.6000 192.4500 1483.8000 192.6000 ;
	    RECT 1449.0000 191.5500 1483.8000 192.4500 ;
	    RECT 1449.0000 191.4000 1450.2001 191.5500 ;
	    RECT 1482.6000 191.4000 1483.8000 191.5500 ;
	    RECT 1485.0000 190.5000 1485.9000 193.5000 ;
	    RECT 1446.9000 189.6000 1452.3000 190.5000 ;
	    RECT 1446.9000 189.3000 1447.8000 189.6000 ;
	    RECT 1446.6000 183.3000 1447.8000 189.3000 ;
	    RECT 1451.4000 189.3000 1452.3000 189.6000 ;
	    RECT 1480.5000 189.6000 1485.9000 190.5000 ;
	    RECT 1480.5000 189.3000 1481.4000 189.6000 ;
	    RECT 1449.0000 183.3000 1450.2001 188.7000 ;
	    RECT 1451.4000 183.3000 1452.6000 189.3000 ;
	    RECT 1453.8000 183.3000 1455.0000 189.3000 ;
	    RECT 1477.8000 183.3000 1479.0000 189.3000 ;
	    RECT 1480.2001 183.3000 1481.4000 189.3000 ;
	    RECT 1485.0000 189.3000 1485.9000 189.6000 ;
	    RECT 1509.3000 190.5000 1510.2001 193.5000 ;
	    RECT 1511.4000 192.4500 1512.6000 192.6000 ;
	    RECT 1528.2001 192.4500 1529.4000 192.6000 ;
	    RECT 1511.4000 191.5500 1529.4000 192.4500 ;
	    RECT 1511.4000 191.4000 1512.6000 191.5500 ;
	    RECT 1528.2001 191.4000 1529.4000 191.5500 ;
	    RECT 1509.3000 189.6000 1514.7001 190.5000 ;
	    RECT 1509.3000 189.3000 1510.2001 189.6000 ;
	    RECT 1482.6000 183.3000 1483.8000 188.7000 ;
	    RECT 1485.0000 183.3000 1486.2001 189.3000 ;
	    RECT 1509.0000 183.3000 1510.2001 189.3000 ;
	    RECT 1513.8000 189.3000 1514.7001 189.6000 ;
	    RECT 1511.4000 183.3000 1512.6000 188.7000 ;
	    RECT 1513.8000 183.3000 1515.0000 189.3000 ;
	    RECT 1516.2001 183.3000 1517.4000 189.3000 ;
	    RECT 1542.6000 183.3000 1543.8000 195.3000 ;
	    RECT 1545.0000 194.4000 1551.0000 195.3000 ;
	    RECT 1545.0000 183.3000 1546.2001 194.4000 ;
	    RECT 1547.4000 183.3000 1548.6000 193.5000 ;
	    RECT 1549.8000 183.3000 1551.0000 194.4000 ;
	    RECT 1.2000 180.6000 1569.0000 182.4000 ;
	    RECT 13.8000 173.7000 15.0000 179.7000 ;
	    RECT 16.2000 163.5000 17.4000 179.7000 ;
	    RECT 40.2000 167.7000 41.4000 179.7000 ;
	    RECT 44.1000 168.6000 45.3000 179.7000 ;
	    RECT 46.5000 173.7000 47.7000 179.7000 ;
	    RECT 172.2000 173.7000 173.4000 179.7000 ;
	    RECT 174.6000 174.6000 175.8000 179.7000 ;
	    RECT 174.3000 173.7000 175.8000 174.6000 ;
	    RECT 177.0000 173.7000 178.2000 180.6000 ;
	    RECT 174.3000 172.8000 175.2000 173.7000 ;
	    RECT 179.4000 172.8000 180.6000 179.7000 ;
	    RECT 181.8000 173.7000 183.0000 179.7000 ;
	    RECT 184.2000 175.5000 185.4000 179.7000 ;
	    RECT 186.6000 175.5000 187.8000 179.7000 ;
	    RECT 172.2000 171.9000 175.2000 172.8000 ;
	    RECT 46.2000 170.4000 47.4000 171.6000 ;
	    RECT 46.5000 169.5000 47.4000 170.4000 ;
	    RECT 44.1000 167.7000 45.6000 168.6000 ;
	    RECT 33.0000 165.4500 34.2000 165.6000 ;
	    RECT 42.6000 165.4500 43.8000 165.6000 ;
	    RECT 33.0000 164.5500 43.8000 165.4500 ;
	    RECT 33.0000 164.4000 34.2000 164.5500 ;
	    RECT 42.6000 164.4000 43.8000 164.5500 ;
	    RECT 42.6000 163.2000 43.8000 163.5000 ;
	    RECT 44.7000 162.6000 45.6000 167.7000 ;
	    RECT 47.4000 167.4000 48.6000 168.6000 ;
	    RECT 172.2000 163.5000 173.4000 171.9000 ;
	    RECT 176.1000 171.6000 182.4000 172.8000 ;
	    RECT 189.0000 172.5000 190.2000 179.7000 ;
	    RECT 191.4000 173.7000 192.6000 179.7000 ;
	    RECT 193.8000 172.5000 195.0000 179.7000 ;
	    RECT 196.2000 173.7000 197.4000 179.7000 ;
	    RECT 176.1000 171.0000 177.0000 171.6000 ;
	    RECT 174.6000 169.8000 177.0000 171.0000 ;
	    RECT 181.5000 170.7000 190.2000 171.6000 ;
	    RECT 178.5000 169.8000 180.6000 170.7000 ;
	    RECT 178.5000 169.5000 187.8000 169.8000 ;
	    RECT 179.7000 168.9000 187.8000 169.5000 ;
	    RECT 186.6000 168.6000 187.8000 168.9000 ;
	    RECT 189.3000 169.5000 190.2000 170.7000 ;
	    RECT 191.1000 170.4000 195.0000 171.6000 ;
	    RECT 198.6000 170.4000 199.8000 179.7000 ;
	    RECT 201.0000 175.5000 202.2000 179.7000 ;
	    RECT 203.4000 175.5000 204.6000 179.7000 ;
	    RECT 205.8000 175.5000 207.0000 179.7000 ;
	    RECT 208.2000 173.7000 209.4000 179.7000 ;
	    RECT 203.4000 171.6000 209.7000 172.8000 ;
	    RECT 210.6000 171.6000 211.8000 179.7000 ;
	    RECT 213.0000 173.7000 214.2000 179.7000 ;
	    RECT 215.4000 172.8000 216.6000 179.7000 ;
	    RECT 217.8000 173.7000 219.0000 179.7000 ;
	    RECT 215.4000 171.9000 219.3000 172.8000 ;
	    RECT 220.2000 172.5000 221.4000 179.7000 ;
	    RECT 222.6000 173.7000 223.8000 179.7000 ;
	    RECT 249.0000 173.7000 250.2000 179.7000 ;
	    RECT 210.6000 170.4000 214.5000 171.6000 ;
	    RECT 201.0000 169.5000 202.2000 169.8000 ;
	    RECT 189.3000 168.6000 202.2000 169.5000 ;
	    RECT 205.8000 169.5000 207.0000 169.8000 ;
	    RECT 218.4000 169.5000 219.3000 171.9000 ;
	    RECT 220.2000 170.4000 221.4000 171.6000 ;
	    RECT 205.8000 168.6000 219.3000 169.5000 ;
	    RECT 177.0000 167.4000 178.2000 168.6000 ;
	    RECT 182.1000 167.7000 183.3000 168.0000 ;
	    RECT 179.1000 166.8000 217.5000 167.7000 ;
	    RECT 216.3000 166.5000 217.5000 166.8000 ;
	    RECT 218.4000 165.9000 219.3000 168.6000 ;
	    RECT 220.2000 168.0000 221.4000 169.5000 ;
	    RECT 220.2000 166.8000 221.7000 168.0000 ;
	    RECT 174.3000 165.0000 180.9000 165.9000 ;
	    RECT 174.3000 164.7000 175.5000 165.0000 ;
	    RECT 181.8000 164.4000 183.0000 165.6000 ;
	    RECT 183.9000 165.0000 209.4000 165.9000 ;
	    RECT 218.4000 165.0000 219.6000 165.9000 ;
	    RECT 208.2000 164.1000 209.4000 165.0000 ;
	    RECT 16.2000 161.4000 17.4000 162.6000 ;
	    RECT 18.6000 162.4500 19.8000 162.6000 ;
	    RECT 40.2000 162.4500 41.4000 162.6000 ;
	    RECT 18.6000 161.5500 41.4000 162.4500 ;
	    RECT 18.6000 161.4000 19.8000 161.5500 ;
	    RECT 40.2000 161.4000 41.4000 161.5500 ;
	    RECT 42.3000 160.8000 42.6000 162.3000 ;
	    RECT 44.7000 161.4000 46.5000 162.6000 ;
	    RECT 47.4000 162.4500 48.6000 162.6000 ;
	    RECT 126.6000 162.4500 127.8000 162.6000 ;
	    RECT 47.4000 161.5500 127.8000 162.4500 ;
	    RECT 47.4000 161.4000 48.6000 161.5500 ;
	    RECT 126.6000 161.4000 127.8000 161.5500 ;
	    RECT 172.2000 162.3000 185.4000 163.5000 ;
	    RECT 186.3000 162.9000 189.3000 164.1000 ;
	    RECT 195.0000 162.9000 199.8000 164.1000 ;
	    RECT 13.8000 158.4000 15.0000 159.6000 ;
	    RECT 13.8000 157.2000 15.0000 157.5000 ;
	    RECT 13.8000 153.3000 15.0000 156.3000 ;
	    RECT 16.2000 153.3000 17.4000 160.5000 ;
	    RECT 40.5000 159.3000 45.9000 159.9000 ;
	    RECT 47.4000 159.3000 48.3000 160.5000 ;
	    RECT 40.2000 159.0000 46.2000 159.3000 ;
	    RECT 40.2000 153.3000 41.4000 159.0000 ;
	    RECT 42.6000 153.3000 43.8000 158.1000 ;
	    RECT 45.0000 153.3000 46.2000 159.0000 ;
	    RECT 47.4000 153.3000 48.6000 159.3000 ;
	    RECT 172.2000 153.3000 173.4000 162.3000 ;
	    RECT 175.8000 160.2000 180.3000 161.4000 ;
	    RECT 179.1000 159.3000 180.3000 160.2000 ;
	    RECT 188.1000 159.3000 189.3000 162.9000 ;
	    RECT 191.4000 161.4000 192.6000 162.6000 ;
	    RECT 199.2000 161.7000 200.4000 162.0000 ;
	    RECT 193.8000 160.8000 200.4000 161.7000 ;
	    RECT 193.8000 160.5000 195.0000 160.8000 ;
	    RECT 191.4000 160.2000 192.6000 160.5000 ;
	    RECT 203.4000 159.6000 204.6000 163.8000 ;
	    RECT 212.1000 162.9000 217.8000 164.1000 ;
	    RECT 212.1000 161.1000 213.3000 162.9000 ;
	    RECT 218.7000 162.0000 219.6000 165.0000 ;
	    RECT 193.8000 159.3000 195.0000 159.6000 ;
	    RECT 177.0000 153.3000 178.2000 159.3000 ;
	    RECT 179.1000 158.1000 183.0000 159.3000 ;
	    RECT 188.1000 158.4000 195.0000 159.3000 ;
	    RECT 196.2000 158.4000 197.4000 159.6000 ;
	    RECT 198.3000 158.4000 198.6000 159.6000 ;
	    RECT 203.1000 158.4000 204.6000 159.6000 ;
	    RECT 210.6000 160.2000 213.3000 161.1000 ;
	    RECT 217.8000 161.1000 219.6000 162.0000 ;
	    RECT 210.6000 159.3000 211.8000 160.2000 ;
	    RECT 181.8000 153.3000 183.0000 158.1000 ;
	    RECT 208.2000 158.1000 211.8000 159.3000 ;
	    RECT 184.2000 153.3000 185.4000 157.5000 ;
	    RECT 186.6000 153.3000 187.8000 157.5000 ;
	    RECT 189.0000 153.3000 190.2000 157.5000 ;
	    RECT 191.4000 153.3000 192.6000 156.3000 ;
	    RECT 193.8000 153.3000 195.0000 157.5000 ;
	    RECT 196.2000 153.3000 197.4000 156.3000 ;
	    RECT 198.6000 153.3000 199.8000 157.5000 ;
	    RECT 201.0000 153.3000 202.2000 157.5000 ;
	    RECT 203.4000 153.3000 204.6000 157.5000 ;
	    RECT 205.8000 153.3000 207.0000 157.5000 ;
	    RECT 208.2000 153.3000 209.4000 158.1000 ;
	    RECT 213.0000 153.3000 214.2000 159.3000 ;
	    RECT 217.8000 153.3000 219.0000 161.1000 ;
	    RECT 220.5000 160.2000 221.7000 166.8000 ;
	    RECT 251.4000 166.5000 252.6000 179.7000 ;
	    RECT 253.8000 173.7000 255.0000 179.7000 ;
	    RECT 273.0000 173.7000 274.2000 179.7000 ;
	    RECT 253.8000 169.5000 255.0000 169.8000 ;
	    RECT 253.8000 168.4500 255.0000 168.6000 ;
	    RECT 256.2000 168.4500 257.4000 168.6000 ;
	    RECT 253.8000 167.5500 257.4000 168.4500 ;
	    RECT 253.8000 167.4000 255.0000 167.5500 ;
	    RECT 256.2000 167.4000 257.4000 167.5500 ;
	    RECT 275.4000 166.5000 276.6000 179.7000 ;
	    RECT 277.8000 173.7000 279.0000 179.7000 ;
	    RECT 405.0000 173.7000 406.2000 179.7000 ;
	    RECT 407.4000 172.5000 408.6000 179.7000 ;
	    RECT 409.8000 173.7000 411.0000 179.7000 ;
	    RECT 412.2000 172.8000 413.4000 179.7000 ;
	    RECT 414.6000 173.7000 415.8000 179.7000 ;
	    RECT 409.5000 171.9000 413.4000 172.8000 ;
	    RECT 289.8000 171.4500 291.0000 171.6000 ;
	    RECT 407.4000 171.4500 408.6000 171.6000 ;
	    RECT 289.8000 170.5500 408.6000 171.4500 ;
	    RECT 289.8000 170.4000 291.0000 170.5500 ;
	    RECT 407.4000 170.4000 408.6000 170.5500 ;
	    RECT 277.8000 169.5000 279.0000 169.8000 ;
	    RECT 409.5000 169.5000 410.4000 171.9000 ;
	    RECT 417.0000 171.6000 418.2000 179.7000 ;
	    RECT 419.4000 173.7000 420.6000 179.7000 ;
	    RECT 421.8000 175.5000 423.0000 179.7000 ;
	    RECT 424.2000 175.5000 425.4000 179.7000 ;
	    RECT 426.6000 175.5000 427.8000 179.7000 ;
	    RECT 419.1000 171.6000 425.4000 172.8000 ;
	    RECT 414.3000 170.4000 418.2000 171.6000 ;
	    RECT 429.0000 170.4000 430.2000 179.7000 ;
	    RECT 431.4000 173.7000 432.6000 179.7000 ;
	    RECT 433.8000 172.5000 435.0000 179.7000 ;
	    RECT 436.2000 173.7000 437.4000 179.7000 ;
	    RECT 438.6000 172.5000 439.8000 179.7000 ;
	    RECT 441.0000 175.5000 442.2000 179.7000 ;
	    RECT 443.4000 175.5000 444.6000 179.7000 ;
	    RECT 445.8000 173.7000 447.0000 179.7000 ;
	    RECT 448.2000 172.8000 449.4000 179.7000 ;
	    RECT 450.6000 173.7000 451.8000 180.6000 ;
	    RECT 453.0000 174.6000 454.2000 179.7000 ;
	    RECT 453.0000 173.7000 454.5000 174.6000 ;
	    RECT 455.4000 173.7000 456.6000 179.7000 ;
	    RECT 487.5000 173.7000 488.7000 179.7000 ;
	    RECT 453.6000 172.8000 454.5000 173.7000 ;
	    RECT 446.4000 171.6000 452.7000 172.8000 ;
	    RECT 453.6000 171.9000 456.6000 172.8000 ;
	    RECT 433.8000 170.4000 437.7000 171.6000 ;
	    RECT 438.6000 170.7000 447.3000 171.6000 ;
	    RECT 451.8000 171.0000 452.7000 171.6000 ;
	    RECT 421.8000 169.5000 423.0000 169.8000 ;
	    RECT 277.8000 168.4500 279.0000 168.6000 ;
	    RECT 289.8000 168.4500 291.0000 168.6000 ;
	    RECT 277.8000 167.5500 291.0000 168.4500 ;
	    RECT 407.4000 168.0000 408.6000 169.5000 ;
	    RECT 277.8000 167.4000 279.0000 167.5500 ;
	    RECT 289.8000 167.4000 291.0000 167.5500 ;
	    RECT 407.1000 166.8000 408.6000 168.0000 ;
	    RECT 409.5000 168.6000 423.0000 169.5000 ;
	    RECT 426.6000 169.5000 427.8000 169.8000 ;
	    RECT 438.6000 169.5000 439.5000 170.7000 ;
	    RECT 448.2000 169.8000 450.3000 170.7000 ;
	    RECT 451.8000 169.8000 454.2000 171.0000 ;
	    RECT 426.6000 168.6000 439.5000 169.5000 ;
	    RECT 441.0000 169.5000 450.3000 169.8000 ;
	    RECT 441.0000 168.9000 449.1000 169.5000 ;
	    RECT 441.0000 168.6000 442.2000 168.9000 ;
	    RECT 251.4000 165.4500 252.6000 165.6000 ;
	    RECT 270.6000 165.4500 271.8000 165.6000 ;
	    RECT 251.4000 164.5500 271.8000 165.4500 ;
	    RECT 251.4000 164.4000 252.6000 164.5500 ;
	    RECT 270.6000 164.4000 271.8000 164.5500 ;
	    RECT 275.4000 165.4500 276.6000 165.6000 ;
	    RECT 285.0000 165.4500 286.2000 165.6000 ;
	    RECT 275.4000 164.5500 286.2000 165.4500 ;
	    RECT 275.4000 164.4000 276.6000 164.5500 ;
	    RECT 285.0000 164.4000 286.2000 164.5500 ;
	    RECT 249.0000 161.4000 250.2000 162.6000 ;
	    RECT 249.0000 160.2000 250.2000 160.5000 ;
	    RECT 220.2000 159.0000 221.7000 160.2000 ;
	    RECT 251.4000 159.3000 252.6000 163.5000 ;
	    RECT 273.0000 161.4000 274.2000 162.6000 ;
	    RECT 273.0000 160.2000 274.2000 160.5000 ;
	    RECT 275.4000 159.3000 276.6000 163.5000 ;
	    RECT 407.1000 160.2000 408.3000 166.8000 ;
	    RECT 409.5000 165.9000 410.4000 168.6000 ;
	    RECT 445.5000 167.7000 446.7000 168.0000 ;
	    RECT 411.3000 166.8000 449.7000 167.7000 ;
	    RECT 450.6000 167.4000 451.8000 168.6000 ;
	    RECT 411.3000 166.5000 412.5000 166.8000 ;
	    RECT 409.2000 165.0000 410.4000 165.9000 ;
	    RECT 419.4000 165.0000 444.9000 165.9000 ;
	    RECT 409.2000 162.0000 410.1000 165.0000 ;
	    RECT 419.4000 164.1000 420.6000 165.0000 ;
	    RECT 445.8000 164.4000 447.0000 165.6000 ;
	    RECT 447.9000 165.0000 454.5000 165.9000 ;
	    RECT 453.3000 164.7000 454.5000 165.0000 ;
	    RECT 411.0000 162.9000 416.7000 164.1000 ;
	    RECT 409.2000 161.1000 411.0000 162.0000 ;
	    RECT 220.2000 153.3000 221.4000 159.0000 ;
	    RECT 222.6000 153.3000 223.8000 156.3000 ;
	    RECT 249.0000 153.3000 250.2000 159.3000 ;
	    RECT 251.4000 158.4000 254.1000 159.3000 ;
	    RECT 252.9000 153.3000 254.1000 158.4000 ;
	    RECT 273.0000 153.3000 274.2000 159.3000 ;
	    RECT 275.4000 158.4000 278.1000 159.3000 ;
	    RECT 407.1000 159.0000 408.6000 160.2000 ;
	    RECT 276.9000 153.3000 278.1000 158.4000 ;
	    RECT 405.0000 153.3000 406.2000 156.3000 ;
	    RECT 407.4000 153.3000 408.6000 159.0000 ;
	    RECT 409.8000 153.3000 411.0000 161.1000 ;
	    RECT 415.5000 161.1000 416.7000 162.9000 ;
	    RECT 415.5000 160.2000 418.2000 161.1000 ;
	    RECT 417.0000 159.3000 418.2000 160.2000 ;
	    RECT 424.2000 159.6000 425.4000 163.8000 ;
	    RECT 429.0000 162.9000 433.8000 164.1000 ;
	    RECT 439.5000 162.9000 442.5000 164.1000 ;
	    RECT 455.4000 163.5000 456.6000 171.9000 ;
	    RECT 487.8000 170.4000 489.0000 171.6000 ;
	    RECT 487.8000 169.5000 488.7000 170.4000 ;
	    RECT 489.9000 168.6000 491.1000 179.7000 ;
	    RECT 457.8000 168.4500 459.0000 168.6000 ;
	    RECT 486.6000 168.4500 487.8000 168.6000 ;
	    RECT 457.8000 167.5500 487.8000 168.4500 ;
	    RECT 457.8000 167.4000 459.0000 167.5500 ;
	    RECT 486.6000 167.4000 487.8000 167.5500 ;
	    RECT 489.6000 167.7000 491.1000 168.6000 ;
	    RECT 493.8000 167.7000 495.0000 179.7000 ;
	    RECT 428.4000 161.7000 429.6000 162.0000 ;
	    RECT 428.4000 160.8000 435.0000 161.7000 ;
	    RECT 436.2000 161.4000 437.4000 162.6000 ;
	    RECT 433.8000 160.5000 435.0000 160.8000 ;
	    RECT 436.2000 160.2000 437.4000 160.5000 ;
	    RECT 414.6000 153.3000 415.8000 159.3000 ;
	    RECT 417.0000 158.1000 420.6000 159.3000 ;
	    RECT 424.2000 158.4000 425.7000 159.6000 ;
	    RECT 430.2000 158.4000 430.5000 159.6000 ;
	    RECT 431.4000 158.4000 432.6000 159.6000 ;
	    RECT 433.8000 159.3000 435.0000 159.6000 ;
	    RECT 439.5000 159.3000 440.7000 162.9000 ;
	    RECT 443.4000 162.3000 456.6000 163.5000 ;
	    RECT 489.6000 162.6000 490.5000 167.7000 ;
	    RECT 491.4000 165.4500 492.6000 165.6000 ;
	    RECT 491.4000 164.5500 497.2500 165.4500 ;
	    RECT 491.4000 164.4000 492.6000 164.5500 ;
	    RECT 491.4000 163.2000 492.6000 163.5000 ;
	    RECT 448.5000 160.2000 453.0000 161.4000 ;
	    RECT 448.5000 159.3000 449.7000 160.2000 ;
	    RECT 433.8000 158.4000 440.7000 159.3000 ;
	    RECT 419.4000 153.3000 420.6000 158.1000 ;
	    RECT 445.8000 158.1000 449.7000 159.3000 ;
	    RECT 421.8000 153.3000 423.0000 157.5000 ;
	    RECT 424.2000 153.3000 425.4000 157.5000 ;
	    RECT 426.6000 153.3000 427.8000 157.5000 ;
	    RECT 429.0000 153.3000 430.2000 157.5000 ;
	    RECT 431.4000 153.3000 432.6000 156.3000 ;
	    RECT 433.8000 153.3000 435.0000 157.5000 ;
	    RECT 436.2000 153.3000 437.4000 156.3000 ;
	    RECT 438.6000 153.3000 439.8000 157.5000 ;
	    RECT 441.0000 153.3000 442.2000 157.5000 ;
	    RECT 443.4000 153.3000 444.6000 157.5000 ;
	    RECT 445.8000 153.3000 447.0000 158.1000 ;
	    RECT 450.6000 153.3000 451.8000 159.3000 ;
	    RECT 455.4000 153.3000 456.6000 162.3000 ;
	    RECT 486.6000 161.4000 487.8000 162.6000 ;
	    RECT 488.7000 161.4000 490.5000 162.6000 ;
	    RECT 492.6000 160.8000 492.9000 162.3000 ;
	    RECT 493.8000 161.4000 495.0000 162.6000 ;
	    RECT 496.3500 162.4500 497.2500 164.5500 ;
	    RECT 508.2000 163.5000 509.4000 179.7000 ;
	    RECT 510.6000 173.7000 511.8000 179.7000 ;
	    RECT 580.2000 166.8000 581.4000 179.7000 ;
	    RECT 582.6000 167.7000 583.8000 179.7000 ;
	    RECT 586.5000 173.7000 588.3000 179.7000 ;
	    RECT 591.0000 173.7000 592.2000 179.7000 ;
	    RECT 593.4000 173.7000 594.6000 179.7000 ;
	    RECT 595.8000 173.7000 597.0000 179.7000 ;
	    RECT 600.0000 174.6000 601.2000 179.7000 ;
	    RECT 600.0000 173.7000 603.0000 174.6000 ;
	    RECT 587.4000 172.5000 588.6000 173.7000 ;
	    RECT 593.7000 172.8000 594.6000 173.7000 ;
	    RECT 592.5000 171.9000 597.9000 172.8000 ;
	    RECT 601.8000 172.5000 603.0000 173.7000 ;
	    RECT 592.5000 171.6000 593.7000 171.9000 ;
	    RECT 596.7000 171.6000 597.9000 171.9000 ;
	    RECT 586.2000 169.8000 588.3000 171.0000 ;
	    RECT 587.4000 168.3000 588.3000 169.8000 ;
	    RECT 590.7000 169.5000 594.0000 170.4000 ;
	    RECT 590.7000 169.2000 591.9000 169.5000 ;
	    RECT 587.4000 167.4000 591.0000 168.3000 ;
	    RECT 580.2000 166.5000 586.5000 166.8000 ;
	    RECT 582.3000 165.9000 586.5000 166.5000 ;
	    RECT 585.3000 165.6000 586.5000 165.9000 ;
	    RECT 510.6000 165.4500 511.8000 165.6000 ;
	    RECT 580.2000 165.4500 581.4000 165.6000 ;
	    RECT 510.6000 164.5500 581.4000 165.4500 ;
	    RECT 510.6000 164.4000 511.8000 164.5500 ;
	    RECT 580.2000 164.4000 581.4000 164.5500 ;
	    RECT 582.9000 164.7000 584.1000 165.0000 ;
	    RECT 582.9000 163.8000 588.6000 164.7000 ;
	    RECT 587.4000 163.5000 588.6000 163.8000 ;
	    RECT 508.2000 162.4500 509.4000 162.6000 ;
	    RECT 496.3500 161.5500 509.4000 162.4500 ;
	    RECT 508.2000 161.4000 509.4000 161.5500 ;
	    RECT 517.8000 162.4500 519.0000 162.6000 ;
	    RECT 558.6000 162.4500 559.8000 162.6000 ;
	    RECT 517.8000 161.5500 559.8000 162.4500 ;
	    RECT 517.8000 161.4000 519.0000 161.5500 ;
	    RECT 558.6000 161.4000 559.8000 161.5500 ;
	    RECT 580.2000 160.8000 581.4000 163.5000 ;
	    RECT 590.1000 162.6000 591.0000 167.4000 ;
	    RECT 593.1000 167.7000 594.0000 169.5000 ;
	    RECT 594.9000 169.5000 596.1000 169.8000 ;
	    RECT 601.8000 169.5000 603.0000 169.8000 ;
	    RECT 594.9000 168.6000 603.0000 169.5000 ;
	    RECT 604.2000 168.0000 605.4000 179.7000 ;
	    RECT 593.1000 167.1000 600.3000 167.7000 ;
	    RECT 606.6000 167.1000 607.8000 179.7000 ;
	    RECT 593.1000 166.8000 607.8000 167.1000 ;
	    RECT 599.1000 166.5000 607.8000 166.8000 ;
	    RECT 599.4000 166.2000 607.8000 166.5000 ;
	    RECT 625.8000 167.7000 627.0000 179.7000 ;
	    RECT 628.2000 169.5000 629.4000 179.7000 ;
	    RECT 630.6000 168.6000 631.8000 179.7000 ;
	    RECT 628.5000 167.7000 631.8000 168.6000 ;
	    RECT 597.0000 164.4000 598.2000 165.6000 ;
	    RECT 599.1000 164.4000 604.5000 165.3000 ;
	    RECT 603.3000 164.1000 604.5000 164.4000 ;
	    RECT 625.8000 164.4000 626.7000 167.7000 ;
	    RECT 628.5000 166.8000 629.4000 167.7000 ;
	    RECT 627.6000 165.6000 629.4000 166.8000 ;
	    RECT 707.4000 166.8000 708.6000 179.7000 ;
	    RECT 709.8000 167.7000 711.0000 179.7000 ;
	    RECT 713.7000 173.7000 715.5000 179.7000 ;
	    RECT 718.2000 173.7000 719.4000 179.7000 ;
	    RECT 720.6000 173.7000 721.8000 179.7000 ;
	    RECT 723.0000 173.7000 724.2000 179.7000 ;
	    RECT 727.2000 174.6000 728.4000 179.7000 ;
	    RECT 727.2000 173.7000 730.2000 174.6000 ;
	    RECT 714.6000 172.5000 715.8000 173.7000 ;
	    RECT 720.9000 172.8000 721.8000 173.7000 ;
	    RECT 719.7000 171.9000 725.1000 172.8000 ;
	    RECT 729.0000 172.5000 730.2000 173.7000 ;
	    RECT 719.7000 171.6000 720.9000 171.9000 ;
	    RECT 723.9000 171.6000 725.1000 171.9000 ;
	    RECT 713.4000 169.8000 715.5000 171.0000 ;
	    RECT 714.6000 168.3000 715.5000 169.8000 ;
	    RECT 717.9000 169.5000 721.2000 170.4000 ;
	    RECT 717.9000 169.2000 719.1000 169.5000 ;
	    RECT 714.6000 167.4000 718.2000 168.3000 ;
	    RECT 707.4000 166.5000 713.7000 166.8000 ;
	    RECT 709.5000 165.9000 713.7000 166.5000 ;
	    RECT 712.5000 165.6000 713.7000 165.9000 ;
	    RECT 625.8000 163.5000 627.0000 164.4000 ;
	    RECT 600.9000 162.6000 602.1000 162.9000 ;
	    RECT 590.1000 161.7000 603.3000 162.6000 ;
	    RECT 590.7000 161.4000 591.9000 161.7000 ;
	    RECT 486.9000 159.3000 487.8000 160.5000 ;
	    RECT 489.3000 159.3000 494.7000 159.9000 ;
	    RECT 486.6000 153.3000 487.8000 159.3000 ;
	    RECT 489.0000 159.0000 495.0000 159.3000 ;
	    RECT 489.0000 153.3000 490.2000 159.0000 ;
	    RECT 491.4000 153.3000 492.6000 158.1000 ;
	    RECT 493.8000 153.3000 495.0000 159.0000 ;
	    RECT 508.2000 153.3000 509.4000 160.5000 ;
	    RECT 580.2000 159.9000 585.9000 160.8000 ;
	    RECT 510.6000 159.4500 511.8000 159.6000 ;
	    RECT 532.2000 159.4500 533.4000 159.6000 ;
	    RECT 577.8000 159.4500 579.0000 159.6000 ;
	    RECT 510.6000 158.5500 579.0000 159.4500 ;
	    RECT 510.6000 158.4000 511.8000 158.5500 ;
	    RECT 532.2000 158.4000 533.4000 158.5500 ;
	    RECT 577.8000 158.4000 579.0000 158.5500 ;
	    RECT 510.6000 157.2000 511.8000 157.5000 ;
	    RECT 546.6000 156.4500 547.8000 156.6000 ;
	    RECT 575.4000 156.4500 576.6000 156.6000 ;
	    RECT 510.6000 153.3000 511.8000 156.3000 ;
	    RECT 546.6000 155.5500 576.6000 156.4500 ;
	    RECT 546.6000 155.4000 547.8000 155.5500 ;
	    RECT 575.4000 155.4000 576.6000 155.5500 ;
	    RECT 580.2000 153.3000 581.4000 159.9000 ;
	    RECT 584.7000 159.6000 585.9000 159.9000 ;
	    RECT 582.6000 153.3000 583.8000 159.0000 ;
	    RECT 599.4000 158.4000 600.3000 161.7000 ;
	    RECT 604.2000 161.4000 605.4000 162.6000 ;
	    RECT 606.3000 161.4000 606.6000 162.6000 ;
	    RECT 625.8000 161.4000 627.0000 162.6000 ;
	    RECT 628.5000 161.1000 629.4000 165.6000 ;
	    RECT 654.6000 165.4500 655.8000 165.6000 ;
	    RECT 707.4000 165.4500 708.6000 165.6000 ;
	    RECT 654.6000 164.5500 708.6000 165.4500 ;
	    RECT 654.6000 164.4000 655.8000 164.5500 ;
	    RECT 707.4000 164.4000 708.6000 164.5500 ;
	    RECT 710.1000 164.7000 711.3000 165.0000 ;
	    RECT 710.1000 163.8000 715.8000 164.7000 ;
	    RECT 714.6000 163.5000 715.8000 163.8000 ;
	    RECT 630.6000 163.2000 631.8000 163.5000 ;
	    RECT 596.7000 158.1000 597.9000 158.4000 ;
	    RECT 587.4000 156.3000 588.6000 157.5000 ;
	    RECT 593.7000 157.2000 597.9000 158.1000 ;
	    RECT 599.4000 157.2000 600.6000 158.4000 ;
	    RECT 593.7000 156.3000 594.6000 157.2000 ;
	    RECT 601.8000 156.3000 603.0000 157.5000 ;
	    RECT 586.5000 155.4000 588.6000 156.3000 ;
	    RECT 586.5000 153.3000 588.3000 155.4000 ;
	    RECT 591.0000 153.3000 592.2000 156.3000 ;
	    RECT 593.4000 153.3000 594.6000 156.3000 ;
	    RECT 595.8000 153.3000 597.3000 156.3000 ;
	    RECT 600.0000 155.4000 603.0000 156.3000 ;
	    RECT 600.0000 153.3000 601.2000 155.4000 ;
	    RECT 604.2000 153.3000 605.4000 159.3000 ;
	    RECT 606.6000 153.3000 607.8000 160.5000 ;
	    RECT 625.8000 153.3000 627.0000 160.5000 ;
	    RECT 628.5000 160.2000 631.8000 161.1000 ;
	    RECT 628.2000 153.3000 629.4000 159.3000 ;
	    RECT 630.6000 153.3000 631.8000 160.2000 ;
	    RECT 707.4000 160.8000 708.6000 163.5000 ;
	    RECT 717.3000 162.6000 718.2000 167.4000 ;
	    RECT 720.3000 167.7000 721.2000 169.5000 ;
	    RECT 722.1000 169.5000 723.3000 169.8000 ;
	    RECT 729.0000 169.5000 730.2000 169.8000 ;
	    RECT 722.1000 168.6000 730.2000 169.5000 ;
	    RECT 731.4000 168.0000 732.6000 179.7000 ;
	    RECT 720.3000 167.1000 727.5000 167.7000 ;
	    RECT 733.8000 167.1000 735.0000 179.7000 ;
	    RECT 757.8000 167.7000 759.0000 179.7000 ;
	    RECT 761.7000 168.6000 762.9000 179.7000 ;
	    RECT 764.1000 173.7000 765.3000 179.7000 ;
	    RECT 779.4000 173.7000 780.6000 179.7000 ;
	    RECT 763.8000 170.4000 765.0000 171.6000 ;
	    RECT 764.1000 169.5000 765.0000 170.4000 ;
	    RECT 761.7000 167.7000 763.2000 168.6000 ;
	    RECT 720.3000 166.8000 735.0000 167.1000 ;
	    RECT 726.3000 166.5000 735.0000 166.8000 ;
	    RECT 726.6000 166.2000 735.0000 166.5000 ;
	    RECT 724.2000 164.4000 725.4000 165.6000 ;
	    RECT 743.4000 165.4500 744.6000 165.6000 ;
	    RECT 760.2000 165.4500 761.4000 165.6000 ;
	    RECT 726.3000 164.4000 731.7000 165.3000 ;
	    RECT 743.4000 164.5500 761.4000 165.4500 ;
	    RECT 743.4000 164.4000 744.6000 164.5500 ;
	    RECT 760.2000 164.4000 761.4000 164.5500 ;
	    RECT 730.5000 164.1000 731.7000 164.4000 ;
	    RECT 760.2000 163.2000 761.4000 163.5000 ;
	    RECT 728.1000 162.6000 729.3000 162.9000 ;
	    RECT 762.3000 162.6000 763.2000 167.7000 ;
	    RECT 765.0000 168.4500 766.2000 168.6000 ;
	    RECT 779.4000 168.4500 780.6000 168.6000 ;
	    RECT 765.0000 167.5500 780.6000 168.4500 ;
	    RECT 765.0000 167.4000 766.2000 167.5500 ;
	    RECT 779.4000 167.4000 780.6000 167.5500 ;
	    RECT 781.8000 163.5000 783.0000 179.7000 ;
	    RECT 832.2000 179.4000 833.4000 180.6000 ;
	    RECT 916.2000 173.7000 917.4000 179.7000 ;
	    RECT 918.6000 174.6000 919.8000 179.7000 ;
	    RECT 918.3000 173.7000 919.8000 174.6000 ;
	    RECT 921.0000 173.7000 922.2000 180.6000 ;
	    RECT 918.3000 172.8000 919.2000 173.7000 ;
	    RECT 923.4000 172.8000 924.6000 179.7000 ;
	    RECT 925.8000 173.7000 927.0000 179.7000 ;
	    RECT 928.2000 175.5000 929.4000 179.7000 ;
	    RECT 930.6000 175.5000 931.8000 179.7000 ;
	    RECT 916.2000 171.9000 919.2000 172.8000 ;
	    RECT 916.2000 163.5000 917.4000 171.9000 ;
	    RECT 920.1000 171.6000 926.4000 172.8000 ;
	    RECT 933.0000 172.5000 934.2000 179.7000 ;
	    RECT 935.4000 173.7000 936.6000 179.7000 ;
	    RECT 937.8000 172.5000 939.0000 179.7000 ;
	    RECT 940.2000 173.7000 941.4000 179.7000 ;
	    RECT 920.1000 171.0000 921.0000 171.6000 ;
	    RECT 918.6000 169.8000 921.0000 171.0000 ;
	    RECT 925.5000 170.7000 934.2000 171.6000 ;
	    RECT 922.5000 169.8000 924.6000 170.7000 ;
	    RECT 922.5000 169.5000 931.8000 169.8000 ;
	    RECT 923.7000 168.9000 931.8000 169.5000 ;
	    RECT 930.6000 168.6000 931.8000 168.9000 ;
	    RECT 933.3000 169.5000 934.2000 170.7000 ;
	    RECT 935.1000 170.4000 939.0000 171.6000 ;
	    RECT 942.6000 170.4000 943.8000 179.7000 ;
	    RECT 945.0000 175.5000 946.2000 179.7000 ;
	    RECT 947.4000 175.5000 948.6000 179.7000 ;
	    RECT 949.8000 175.5000 951.0000 179.7000 ;
	    RECT 952.2000 173.7000 953.4000 179.7000 ;
	    RECT 947.4000 171.6000 953.7000 172.8000 ;
	    RECT 954.6000 171.6000 955.8000 179.7000 ;
	    RECT 957.0000 173.7000 958.2000 179.7000 ;
	    RECT 959.4000 172.8000 960.6000 179.7000 ;
	    RECT 961.8000 173.7000 963.0000 179.7000 ;
	    RECT 959.4000 171.9000 963.3000 172.8000 ;
	    RECT 964.2000 172.5000 965.4000 179.7000 ;
	    RECT 966.6000 173.7000 967.8000 179.7000 ;
	    RECT 993.9000 173.7000 995.1000 179.7000 ;
	    RECT 954.6000 170.4000 958.5000 171.6000 ;
	    RECT 945.0000 169.5000 946.2000 169.8000 ;
	    RECT 933.3000 168.6000 946.2000 169.5000 ;
	    RECT 949.8000 169.5000 951.0000 169.8000 ;
	    RECT 962.4000 169.5000 963.3000 171.9000 ;
	    RECT 964.2000 171.4500 965.4000 171.6000 ;
	    RECT 978.6000 171.4500 979.8000 171.6000 ;
	    RECT 983.4000 171.4500 984.6000 171.6000 ;
	    RECT 964.2000 170.5500 984.6000 171.4500 ;
	    RECT 964.2000 170.4000 965.4000 170.5500 ;
	    RECT 978.6000 170.4000 979.8000 170.5500 ;
	    RECT 983.4000 170.4000 984.6000 170.5500 ;
	    RECT 994.2000 170.4000 995.4000 171.6000 ;
	    RECT 994.2000 169.5000 995.1000 170.4000 ;
	    RECT 949.8000 168.6000 963.3000 169.5000 ;
	    RECT 921.0000 167.4000 922.2000 168.6000 ;
	    RECT 926.1000 167.7000 927.3000 168.0000 ;
	    RECT 923.1000 166.8000 961.5000 167.7000 ;
	    RECT 960.3000 166.5000 961.5000 166.8000 ;
	    RECT 962.4000 165.9000 963.3000 168.6000 ;
	    RECT 964.2000 168.0000 965.4000 169.5000 ;
	    RECT 996.3000 168.6000 997.5000 179.7000 ;
	    RECT 964.2000 166.8000 965.7000 168.0000 ;
	    RECT 993.0000 167.4000 994.2000 168.6000 ;
	    RECT 996.0000 167.7000 997.5000 168.6000 ;
	    RECT 1000.2000 167.7000 1001.4000 179.7000 ;
	    RECT 918.3000 165.0000 924.9000 165.9000 ;
	    RECT 918.3000 164.7000 919.5000 165.0000 ;
	    RECT 925.8000 164.4000 927.0000 165.6000 ;
	    RECT 927.9000 165.0000 953.4000 165.9000 ;
	    RECT 962.4000 165.0000 963.6000 165.9000 ;
	    RECT 952.2000 164.1000 953.4000 165.0000 ;
	    RECT 717.3000 161.7000 730.5000 162.6000 ;
	    RECT 717.9000 161.4000 719.1000 161.7000 ;
	    RECT 707.4000 159.9000 713.1000 160.8000 ;
	    RECT 707.4000 153.3000 708.6000 159.9000 ;
	    RECT 711.9000 159.6000 713.1000 159.9000 ;
	    RECT 709.8000 153.3000 711.0000 159.0000 ;
	    RECT 726.6000 158.4000 727.5000 161.7000 ;
	    RECT 731.4000 161.4000 732.6000 162.6000 ;
	    RECT 733.5000 161.4000 733.8000 162.6000 ;
	    RECT 753.0000 162.4500 754.2000 162.6000 ;
	    RECT 757.8000 162.4500 759.0000 162.6000 ;
	    RECT 753.0000 161.5500 759.0000 162.4500 ;
	    RECT 753.0000 161.4000 754.2000 161.5500 ;
	    RECT 757.8000 161.4000 759.0000 161.5500 ;
	    RECT 759.9000 160.8000 760.2000 162.3000 ;
	    RECT 762.3000 161.4000 764.1000 162.6000 ;
	    RECT 765.0000 162.4500 766.2000 162.6000 ;
	    RECT 774.6000 162.4500 775.8000 162.6000 ;
	    RECT 765.0000 161.5500 775.8000 162.4500 ;
	    RECT 765.0000 161.4000 766.2000 161.5500 ;
	    RECT 774.6000 161.4000 775.8000 161.5500 ;
	    RECT 781.8000 162.4500 783.0000 162.6000 ;
	    RECT 803.4000 162.4500 804.6000 162.6000 ;
	    RECT 781.8000 161.5500 804.6000 162.4500 ;
	    RECT 781.8000 161.4000 783.0000 161.5500 ;
	    RECT 803.4000 161.4000 804.6000 161.5500 ;
	    RECT 916.2000 162.3000 929.4000 163.5000 ;
	    RECT 930.3000 162.9000 933.3000 164.1000 ;
	    RECT 939.0000 162.9000 943.8000 164.1000 ;
	    RECT 723.9000 158.1000 725.1000 158.4000 ;
	    RECT 714.6000 156.3000 715.8000 157.5000 ;
	    RECT 720.9000 157.2000 725.1000 158.1000 ;
	    RECT 726.6000 157.2000 727.8000 158.4000 ;
	    RECT 720.9000 156.3000 721.8000 157.2000 ;
	    RECT 729.0000 156.3000 730.2000 157.5000 ;
	    RECT 713.7000 155.4000 715.8000 156.3000 ;
	    RECT 713.7000 153.3000 715.5000 155.4000 ;
	    RECT 718.2000 153.3000 719.4000 156.3000 ;
	    RECT 720.6000 153.3000 721.8000 156.3000 ;
	    RECT 723.0000 153.3000 724.5000 156.3000 ;
	    RECT 727.2000 155.4000 730.2000 156.3000 ;
	    RECT 727.2000 153.3000 728.4000 155.4000 ;
	    RECT 731.4000 153.3000 732.6000 159.3000 ;
	    RECT 733.8000 153.3000 735.0000 160.5000 ;
	    RECT 758.1000 159.3000 763.5000 159.9000 ;
	    RECT 765.0000 159.3000 765.9000 160.5000 ;
	    RECT 757.8000 159.0000 763.8000 159.3000 ;
	    RECT 757.8000 153.3000 759.0000 159.0000 ;
	    RECT 760.2000 153.3000 761.4000 158.1000 ;
	    RECT 762.6000 153.3000 763.8000 159.0000 ;
	    RECT 765.0000 153.3000 766.2000 159.3000 ;
	    RECT 779.4000 158.4000 780.6000 159.6000 ;
	    RECT 779.4000 157.2000 780.6000 157.5000 ;
	    RECT 779.4000 153.3000 780.6000 156.3000 ;
	    RECT 781.8000 153.3000 783.0000 160.5000 ;
	    RECT 916.2000 153.3000 917.4000 162.3000 ;
	    RECT 919.8000 160.2000 924.3000 161.4000 ;
	    RECT 923.1000 159.3000 924.3000 160.2000 ;
	    RECT 932.1000 159.3000 933.3000 162.9000 ;
	    RECT 935.4000 161.4000 936.6000 162.6000 ;
	    RECT 943.2000 161.7000 944.4000 162.0000 ;
	    RECT 937.8000 160.8000 944.4000 161.7000 ;
	    RECT 937.8000 160.5000 939.0000 160.8000 ;
	    RECT 935.4000 160.2000 936.6000 160.5000 ;
	    RECT 947.4000 159.6000 948.6000 163.8000 ;
	    RECT 956.1000 162.9000 961.8000 164.1000 ;
	    RECT 956.1000 161.1000 957.3000 162.9000 ;
	    RECT 962.7000 162.0000 963.6000 165.0000 ;
	    RECT 937.8000 159.3000 939.0000 159.6000 ;
	    RECT 921.0000 153.3000 922.2000 159.3000 ;
	    RECT 923.1000 158.1000 927.0000 159.3000 ;
	    RECT 932.1000 158.4000 939.0000 159.3000 ;
	    RECT 940.2000 158.4000 941.4000 159.6000 ;
	    RECT 942.3000 158.4000 942.6000 159.6000 ;
	    RECT 947.1000 158.4000 948.6000 159.6000 ;
	    RECT 954.6000 160.2000 957.3000 161.1000 ;
	    RECT 961.8000 161.1000 963.6000 162.0000 ;
	    RECT 954.6000 159.3000 955.8000 160.2000 ;
	    RECT 925.8000 153.3000 927.0000 158.1000 ;
	    RECT 952.2000 158.1000 955.8000 159.3000 ;
	    RECT 928.2000 153.3000 929.4000 157.5000 ;
	    RECT 930.6000 153.3000 931.8000 157.5000 ;
	    RECT 933.0000 153.3000 934.2000 157.5000 ;
	    RECT 935.4000 153.3000 936.6000 156.3000 ;
	    RECT 937.8000 153.3000 939.0000 157.5000 ;
	    RECT 940.2000 153.3000 941.4000 156.3000 ;
	    RECT 942.6000 153.3000 943.8000 157.5000 ;
	    RECT 945.0000 153.3000 946.2000 157.5000 ;
	    RECT 947.4000 153.3000 948.6000 157.5000 ;
	    RECT 949.8000 153.3000 951.0000 157.5000 ;
	    RECT 952.2000 153.3000 953.4000 158.1000 ;
	    RECT 957.0000 153.3000 958.2000 159.3000 ;
	    RECT 961.8000 153.3000 963.0000 161.1000 ;
	    RECT 964.5000 160.2000 965.7000 166.8000 ;
	    RECT 996.0000 162.6000 996.9000 167.7000 ;
	    RECT 997.8000 164.4000 999.0000 165.6000 ;
	    RECT 1014.6000 163.5000 1015.8000 179.7000 ;
	    RECT 1017.0000 173.7000 1018.2000 179.7000 ;
	    RECT 1036.2001 173.7000 1037.4000 179.7000 ;
	    RECT 1036.2001 169.5000 1037.4000 169.8000 ;
	    RECT 1033.8000 168.4500 1035.0000 168.6000 ;
	    RECT 1036.2001 168.4500 1037.4000 168.6000 ;
	    RECT 1033.8000 167.5500 1037.4000 168.4500 ;
	    RECT 1033.8000 167.4000 1035.0000 167.5500 ;
	    RECT 1036.2001 167.4000 1037.4000 167.5500 ;
	    RECT 1038.6000 166.5000 1039.8000 179.7000 ;
	    RECT 1041.0000 173.7000 1042.2001 179.7000 ;
	    RECT 1065.0000 173.7000 1066.2001 179.7000 ;
	    RECT 1067.4000 173.7000 1068.6000 179.7000 ;
	    RECT 1069.8000 174.3000 1071.0000 179.7000 ;
	    RECT 1067.7001 173.4000 1068.6000 173.7000 ;
	    RECT 1072.2001 173.7000 1073.4000 179.7000 ;
	    RECT 1096.2001 173.7000 1097.4000 179.7000 ;
	    RECT 1098.6000 173.7000 1099.8000 179.7000 ;
	    RECT 1101.0000 174.3000 1102.2001 179.7000 ;
	    RECT 1072.2001 173.4000 1073.1000 173.7000 ;
	    RECT 1067.7001 172.5000 1073.1000 173.4000 ;
	    RECT 1098.9000 173.4000 1099.8000 173.7000 ;
	    RECT 1103.4000 173.7000 1104.6000 179.7000 ;
	    RECT 1137.0000 173.7000 1138.2001 179.7000 ;
	    RECT 1139.4000 173.7000 1140.6000 179.7000 ;
	    RECT 1141.8000 174.3000 1143.0000 179.7000 ;
	    RECT 1103.4000 173.4000 1104.3000 173.7000 ;
	    RECT 1098.9000 172.5000 1104.3000 173.4000 ;
	    RECT 1139.7001 173.4000 1140.6000 173.7000 ;
	    RECT 1144.2001 173.7000 1145.4000 179.7000 ;
	    RECT 1146.6000 177.4500 1147.8000 177.6000 ;
	    RECT 1163.4000 177.4500 1164.6000 177.6000 ;
	    RECT 1146.6000 176.5500 1164.6000 177.4500 ;
	    RECT 1146.6000 176.4000 1147.8000 176.5500 ;
	    RECT 1163.4000 176.4000 1164.6000 176.5500 ;
	    RECT 1170.6000 173.7000 1171.8000 179.7000 ;
	    RECT 1173.0000 173.7000 1174.2001 179.7000 ;
	    RECT 1144.2001 173.4000 1145.1000 173.7000 ;
	    RECT 1139.7001 172.5000 1145.1000 173.4000 ;
	    RECT 1048.2001 171.4500 1049.4000 171.6000 ;
	    RECT 1069.8000 171.4500 1071.0000 171.6000 ;
	    RECT 1048.2001 170.5500 1071.0000 171.4500 ;
	    RECT 1048.2001 170.4000 1049.4000 170.5500 ;
	    RECT 1069.8000 170.4000 1071.0000 170.5500 ;
	    RECT 1072.2001 169.5000 1073.1000 172.5000 ;
	    RECT 1079.4000 171.4500 1080.6000 171.6000 ;
	    RECT 1101.0000 171.4500 1102.2001 171.6000 ;
	    RECT 1079.4000 170.5500 1102.2001 171.4500 ;
	    RECT 1079.4000 170.4000 1080.6000 170.5500 ;
	    RECT 1101.0000 170.4000 1102.2001 170.5500 ;
	    RECT 1103.4000 169.5000 1104.3000 172.5000 ;
	    RECT 1120.2001 171.4500 1121.4000 171.6000 ;
	    RECT 1139.4000 171.4500 1140.6000 171.6000 ;
	    RECT 1120.2001 170.5500 1140.6000 171.4500 ;
	    RECT 1120.2001 170.4000 1121.4000 170.5500 ;
	    RECT 1139.4000 170.4000 1140.6000 170.5500 ;
	    RECT 1141.8000 170.4000 1143.0000 171.6000 ;
	    RECT 1144.2001 169.5000 1145.1000 172.5000 ;
	    RECT 1069.8000 169.2000 1071.0000 169.5000 ;
	    RECT 1101.0000 169.2000 1102.2001 169.5000 ;
	    RECT 1141.8000 169.2000 1143.0000 169.5000 ;
	    RECT 1057.8000 168.4500 1059.0000 168.6000 ;
	    RECT 1065.0000 168.4500 1066.2001 168.6000 ;
	    RECT 1057.8000 167.5500 1066.2001 168.4500 ;
	    RECT 1057.8000 167.4000 1059.0000 167.5500 ;
	    RECT 1065.0000 167.4000 1066.2001 167.5500 ;
	    RECT 1072.2001 168.4500 1073.4000 168.6000 ;
	    RECT 1096.2001 168.4500 1097.4000 168.6000 ;
	    RECT 1072.2001 167.5500 1097.4000 168.4500 ;
	    RECT 1072.2001 167.4000 1073.4000 167.5500 ;
	    RECT 1096.2001 167.4000 1097.4000 167.5500 ;
	    RECT 1103.4000 167.4000 1104.6000 168.6000 ;
	    RECT 1108.2001 168.4500 1109.4000 168.6000 ;
	    RECT 1137.0000 168.4500 1138.2001 168.6000 ;
	    RECT 1108.2001 167.5500 1138.2001 168.4500 ;
	    RECT 1108.2001 167.4000 1109.4000 167.5500 ;
	    RECT 1137.0000 167.4000 1138.2001 167.5500 ;
	    RECT 1144.2001 168.4500 1145.4000 168.6000 ;
	    RECT 1149.0000 168.4500 1150.2001 168.6000 ;
	    RECT 1144.2001 167.5500 1150.2001 168.4500 ;
	    RECT 1144.2001 167.4000 1145.4000 167.5500 ;
	    RECT 1149.0000 167.4000 1150.2001 167.5500 ;
	    RECT 1151.4000 168.4500 1152.6000 168.6000 ;
	    RECT 1170.6000 168.4500 1171.8000 168.6000 ;
	    RECT 1151.4000 167.5500 1171.8000 168.4500 ;
	    RECT 1151.4000 167.4000 1152.6000 167.5500 ;
	    RECT 1170.6000 167.4000 1171.8000 167.5500 ;
	    RECT 1173.3000 167.4000 1174.2001 173.7000 ;
	    RECT 1175.4000 168.3000 1176.6000 179.7000 ;
	    RECT 1177.8000 167.7000 1179.0000 179.7000 ;
	    RECT 1197.0000 173.7000 1198.2001 179.7000 ;
	    RECT 1173.3000 166.5000 1176.9000 167.4000 ;
	    RECT 1178.1000 166.5000 1179.0000 167.7000 ;
	    RECT 1199.4000 166.5000 1200.6000 179.7000 ;
	    RECT 1201.8000 173.7000 1203.0000 179.7000 ;
	    RECT 1216.2001 173.7000 1217.4000 179.7000 ;
	    RECT 1201.8000 169.5000 1203.0000 169.8000 ;
	    RECT 1201.8000 167.4000 1203.0000 168.6000 ;
	    RECT 1065.0000 166.2000 1066.2001 166.5000 ;
	    RECT 1038.6000 165.4500 1039.8000 165.6000 ;
	    RECT 1050.6000 165.4500 1051.8000 165.6000 ;
	    RECT 1038.6000 164.5500 1051.8000 165.4500 ;
	    RECT 1038.6000 164.4000 1039.8000 164.5500 ;
	    RECT 1050.6000 164.4000 1051.8000 164.5500 ;
	    RECT 1067.4000 164.4000 1068.6000 165.6000 ;
	    RECT 1069.5000 164.4000 1069.8000 165.6000 ;
	    RECT 997.8000 163.2000 999.0000 163.5000 ;
	    RECT 993.0000 161.4000 994.2000 162.6000 ;
	    RECT 995.1000 161.4000 996.9000 162.6000 ;
	    RECT 999.0000 160.8000 999.3000 162.3000 ;
	    RECT 1000.2000 161.4000 1001.4000 162.6000 ;
	    RECT 1002.6000 162.4500 1003.8000 162.6000 ;
	    RECT 1014.6000 162.4500 1015.8000 162.6000 ;
	    RECT 1002.6000 161.5500 1015.8000 162.4500 ;
	    RECT 1002.6000 161.4000 1003.8000 161.5500 ;
	    RECT 1014.6000 161.4000 1015.8000 161.5500 ;
	    RECT 964.2000 159.0000 965.7000 160.2000 ;
	    RECT 993.3000 159.3000 994.2000 160.5000 ;
	    RECT 995.7000 159.3000 1001.1000 159.9000 ;
	    RECT 964.2000 153.3000 965.4000 159.0000 ;
	    RECT 966.6000 153.3000 967.8000 156.3000 ;
	    RECT 993.0000 153.3000 994.2000 159.3000 ;
	    RECT 995.4000 159.0000 1001.4000 159.3000 ;
	    RECT 995.4000 153.3000 996.6000 159.0000 ;
	    RECT 997.8000 153.3000 999.0000 158.1000 ;
	    RECT 1000.2000 153.3000 1001.4000 159.0000 ;
	    RECT 1014.6000 153.3000 1015.8000 160.5000 ;
	    RECT 1017.0000 158.4000 1018.2000 159.6000 ;
	    RECT 1038.6000 159.3000 1039.8000 163.5000 ;
	    RECT 1072.2001 162.6000 1073.1000 166.5000 ;
	    RECT 1096.2001 166.2000 1097.4000 166.5000 ;
	    RECT 1098.6000 164.4000 1099.8000 165.6000 ;
	    RECT 1100.7001 164.4000 1101.0000 165.6000 ;
	    RECT 1103.4000 162.6000 1104.3000 166.5000 ;
	    RECT 1137.0000 166.2000 1138.2001 166.5000 ;
	    RECT 1139.4000 164.4000 1140.6000 165.6000 ;
	    RECT 1141.5000 164.4000 1141.8000 165.6000 ;
	    RECT 1144.2001 162.6000 1145.1000 166.5000 ;
	    RECT 1173.0000 164.4000 1174.2001 165.6000 ;
	    RECT 1170.6000 163.5000 1171.8000 163.8000 ;
	    RECT 1173.3000 163.2000 1174.2001 163.5000 ;
	    RECT 1041.0000 161.4000 1042.2001 162.6000 ;
	    RECT 1070.7001 162.3000 1073.1000 162.6000 ;
	    RECT 1101.9000 162.3000 1104.3000 162.6000 ;
	    RECT 1142.7001 162.3000 1145.1000 162.6000 ;
	    RECT 1041.0000 160.2000 1042.2001 160.5000 ;
	    RECT 1037.1000 158.4000 1039.8000 159.3000 ;
	    RECT 1017.0000 157.2000 1018.2000 157.5000 ;
	    RECT 1017.0000 153.3000 1018.2000 156.3000 ;
	    RECT 1037.1000 153.3000 1038.3000 158.4000 ;
	    RECT 1041.0000 153.3000 1042.2001 159.3000 ;
	    RECT 1065.0000 153.3000 1066.2001 162.3000 ;
	    RECT 1070.4000 161.7000 1073.1000 162.3000 ;
	    RECT 1070.4000 153.3000 1071.6000 161.7000 ;
	    RECT 1096.2001 153.3000 1097.4000 162.3000 ;
	    RECT 1101.6000 161.7000 1104.3000 162.3000 ;
	    RECT 1101.6000 153.3000 1102.8000 161.7000 ;
	    RECT 1105.8000 156.4500 1107.0000 156.6000 ;
	    RECT 1132.2001 156.4500 1133.4000 156.6000 ;
	    RECT 1105.8000 155.5500 1133.4000 156.4500 ;
	    RECT 1105.8000 155.4000 1107.0000 155.5500 ;
	    RECT 1132.2001 155.4000 1133.4000 155.5500 ;
	    RECT 1137.0000 153.3000 1138.2001 162.3000 ;
	    RECT 1142.4000 161.7000 1145.1000 162.3000 ;
	    RECT 1158.6000 162.4500 1159.8000 162.6000 ;
	    RECT 1165.8000 162.4500 1167.0000 162.6000 ;
	    RECT 1170.6000 162.4500 1171.8000 162.6000 ;
	    RECT 1142.4000 153.3000 1143.6000 161.7000 ;
	    RECT 1158.6000 161.5500 1171.8000 162.4500 ;
	    RECT 1173.3000 162.3000 1174.8000 163.2000 ;
	    RECT 1173.6000 162.0000 1174.8000 162.3000 ;
	    RECT 1158.6000 161.4000 1159.8000 161.5500 ;
	    RECT 1165.8000 161.4000 1167.0000 161.5500 ;
	    RECT 1170.6000 161.4000 1171.8000 161.5500 ;
	    RECT 1176.0000 161.4000 1176.9000 166.5000 ;
	    RECT 1177.8000 165.4500 1179.0000 165.6000 ;
	    RECT 1180.2001 165.4500 1181.4000 165.6000 ;
	    RECT 1177.8000 164.5500 1181.4000 165.4500 ;
	    RECT 1177.8000 164.4000 1179.0000 164.5500 ;
	    RECT 1180.2001 164.4000 1181.4000 164.5500 ;
	    RECT 1199.4000 164.4000 1200.6000 165.6000 ;
	    RECT 1218.6000 163.5000 1219.8000 179.7000 ;
	    RECT 1350.6000 173.7000 1351.8000 179.7000 ;
	    RECT 1353.0000 174.6000 1354.2001 179.7000 ;
	    RECT 1352.7001 173.7000 1354.2001 174.6000 ;
	    RECT 1355.4000 173.7000 1356.6000 180.6000 ;
	    RECT 1352.7001 172.8000 1353.6000 173.7000 ;
	    RECT 1357.8000 172.8000 1359.0000 179.7000 ;
	    RECT 1360.2001 173.7000 1361.4000 179.7000 ;
	    RECT 1362.6000 175.5000 1363.8000 179.7000 ;
	    RECT 1365.0000 175.5000 1366.2001 179.7000 ;
	    RECT 1350.6000 171.9000 1353.6000 172.8000 ;
	    RECT 1350.6000 163.5000 1351.8000 171.9000 ;
	    RECT 1354.5000 171.6000 1360.8000 172.8000 ;
	    RECT 1367.4000 172.5000 1368.6000 179.7000 ;
	    RECT 1369.8000 173.7000 1371.0000 179.7000 ;
	    RECT 1372.2001 172.5000 1373.4000 179.7000 ;
	    RECT 1374.6000 173.7000 1375.8000 179.7000 ;
	    RECT 1354.5000 171.0000 1355.4000 171.6000 ;
	    RECT 1353.0000 169.8000 1355.4000 171.0000 ;
	    RECT 1359.9000 170.7000 1368.6000 171.6000 ;
	    RECT 1356.9000 169.8000 1359.0000 170.7000 ;
	    RECT 1356.9000 169.5000 1366.2001 169.8000 ;
	    RECT 1358.1000 168.9000 1366.2001 169.5000 ;
	    RECT 1365.0000 168.6000 1366.2001 168.9000 ;
	    RECT 1367.7001 169.5000 1368.6000 170.7000 ;
	    RECT 1369.5000 170.4000 1373.4000 171.6000 ;
	    RECT 1377.0000 170.4000 1378.2001 179.7000 ;
	    RECT 1379.4000 175.5000 1380.6000 179.7000 ;
	    RECT 1381.8000 175.5000 1383.0000 179.7000 ;
	    RECT 1384.2001 175.5000 1385.4000 179.7000 ;
	    RECT 1386.6000 173.7000 1387.8000 179.7000 ;
	    RECT 1381.8000 171.6000 1388.1000 172.8000 ;
	    RECT 1389.0000 171.6000 1390.2001 179.7000 ;
	    RECT 1391.4000 173.7000 1392.6000 179.7000 ;
	    RECT 1393.8000 172.8000 1395.0000 179.7000 ;
	    RECT 1396.2001 173.7000 1397.4000 179.7000 ;
	    RECT 1393.8000 171.9000 1397.7001 172.8000 ;
	    RECT 1398.6000 172.5000 1399.8000 179.7000 ;
	    RECT 1401.0000 173.7000 1402.2001 179.7000 ;
	    RECT 1389.0000 170.4000 1392.9000 171.6000 ;
	    RECT 1379.4000 169.5000 1380.6000 169.8000 ;
	    RECT 1367.7001 168.6000 1380.6000 169.5000 ;
	    RECT 1384.2001 169.5000 1385.4000 169.8000 ;
	    RECT 1396.8000 169.5000 1397.7001 171.9000 ;
	    RECT 1398.6000 170.4000 1399.8000 171.6000 ;
	    RECT 1384.2001 168.6000 1397.7001 169.5000 ;
	    RECT 1355.4000 167.4000 1356.6000 168.6000 ;
	    RECT 1360.5000 167.7000 1361.7001 168.0000 ;
	    RECT 1357.5000 166.8000 1395.9000 167.7000 ;
	    RECT 1394.7001 166.5000 1395.9000 166.8000 ;
	    RECT 1396.8000 165.9000 1397.7001 168.6000 ;
	    RECT 1398.6000 168.0000 1399.8000 169.5000 ;
	    RECT 1398.6000 166.8000 1400.1000 168.0000 ;
	    RECT 1420.2001 167.7000 1421.4000 179.7000 ;
	    RECT 1424.1000 168.9000 1425.3000 179.7000 ;
	    RECT 1429.8000 174.4500 1431.0000 174.6000 ;
	    RECT 1441.8000 174.4500 1443.0000 174.6000 ;
	    RECT 1429.8000 173.5500 1443.0000 174.4500 ;
	    RECT 1444.2001 173.7000 1445.4000 179.7000 ;
	    RECT 1429.8000 173.4000 1431.0000 173.5500 ;
	    RECT 1441.8000 173.4000 1443.0000 173.5500 ;
	    RECT 1444.2001 169.5000 1445.4000 169.8000 ;
	    RECT 1422.6000 167.7000 1425.3000 168.9000 ;
	    RECT 1352.7001 165.0000 1359.3000 165.9000 ;
	    RECT 1352.7001 164.7000 1353.9000 165.0000 ;
	    RECT 1360.2001 164.4000 1361.4000 165.6000 ;
	    RECT 1362.3000 165.0000 1387.8000 165.9000 ;
	    RECT 1396.8000 165.0000 1398.0000 165.9000 ;
	    RECT 1386.6000 164.1000 1387.8000 165.0000 ;
	    RECT 1176.0000 161.1000 1177.2001 161.4000 ;
	    RECT 1172.7001 160.5000 1177.2001 161.1000 ;
	    RECT 1170.9000 160.2000 1177.2001 160.5000 ;
	    RECT 1170.9000 159.6000 1173.6000 160.2000 ;
	    RECT 1170.9000 159.3000 1171.8000 159.6000 ;
	    RECT 1178.1000 159.3000 1179.0000 163.5000 ;
	    RECT 1197.0000 161.4000 1198.2001 162.6000 ;
	    RECT 1197.0000 160.2000 1198.2001 160.5000 ;
	    RECT 1199.4000 159.3000 1200.6000 163.5000 ;
	    RECT 1218.6000 162.4500 1219.8000 162.6000 ;
	    RECT 1288.2001 162.4500 1289.4000 162.6000 ;
	    RECT 1218.6000 161.5500 1289.4000 162.4500 ;
	    RECT 1218.6000 161.4000 1219.8000 161.5500 ;
	    RECT 1288.2001 161.4000 1289.4000 161.5500 ;
	    RECT 1350.6000 162.3000 1363.8000 163.5000 ;
	    RECT 1364.7001 162.9000 1367.7001 164.1000 ;
	    RECT 1373.4000 162.9000 1378.2001 164.1000 ;
	    RECT 1204.2001 159.4500 1205.4000 159.6000 ;
	    RECT 1216.2001 159.4500 1217.4000 159.6000 ;
	    RECT 1170.6000 153.3000 1171.8000 159.3000 ;
	    RECT 1174.5000 153.3000 1175.7001 159.0000 ;
	    RECT 1176.9000 157.8000 1179.0000 159.3000 ;
	    RECT 1176.9000 153.3000 1178.1000 157.8000 ;
	    RECT 1197.0000 153.3000 1198.2001 159.3000 ;
	    RECT 1199.4000 158.4000 1202.1000 159.3000 ;
	    RECT 1204.2001 158.5500 1217.4000 159.4500 ;
	    RECT 1204.2001 158.4000 1205.4000 158.5500 ;
	    RECT 1216.2001 158.4000 1217.4000 158.5500 ;
	    RECT 1200.9000 153.3000 1202.1000 158.4000 ;
	    RECT 1216.2001 157.2000 1217.4000 157.5000 ;
	    RECT 1216.2001 153.3000 1217.4000 156.3000 ;
	    RECT 1218.6000 153.3000 1219.8000 160.5000 ;
	    RECT 1350.6000 153.3000 1351.8000 162.3000 ;
	    RECT 1354.2001 160.2000 1358.7001 161.4000 ;
	    RECT 1357.5000 159.3000 1358.7001 160.2000 ;
	    RECT 1366.5000 159.3000 1367.7001 162.9000 ;
	    RECT 1369.8000 161.4000 1371.0000 162.6000 ;
	    RECT 1377.6000 161.7000 1378.8000 162.0000 ;
	    RECT 1372.2001 160.8000 1378.8000 161.7000 ;
	    RECT 1372.2001 160.5000 1373.4000 160.8000 ;
	    RECT 1369.8000 160.2000 1371.0000 160.5000 ;
	    RECT 1381.8000 159.6000 1383.0000 163.8000 ;
	    RECT 1390.5000 162.9000 1396.2001 164.1000 ;
	    RECT 1390.5000 161.1000 1391.7001 162.9000 ;
	    RECT 1397.1000 162.0000 1398.0000 165.0000 ;
	    RECT 1372.2001 159.3000 1373.4000 159.6000 ;
	    RECT 1355.4000 153.3000 1356.6000 159.3000 ;
	    RECT 1357.5000 158.1000 1361.4000 159.3000 ;
	    RECT 1366.5000 158.4000 1373.4000 159.3000 ;
	    RECT 1374.6000 158.4000 1375.8000 159.6000 ;
	    RECT 1376.7001 158.4000 1377.0000 159.6000 ;
	    RECT 1381.5000 158.4000 1383.0000 159.6000 ;
	    RECT 1389.0000 160.2000 1391.7001 161.1000 ;
	    RECT 1396.2001 161.1000 1398.0000 162.0000 ;
	    RECT 1389.0000 159.3000 1390.2001 160.2000 ;
	    RECT 1360.2001 153.3000 1361.4000 158.1000 ;
	    RECT 1386.6000 158.1000 1390.2001 159.3000 ;
	    RECT 1362.6000 153.3000 1363.8000 157.5000 ;
	    RECT 1365.0000 153.3000 1366.2001 157.5000 ;
	    RECT 1367.4000 153.3000 1368.6000 157.5000 ;
	    RECT 1369.8000 153.3000 1371.0000 156.3000 ;
	    RECT 1372.2001 153.3000 1373.4000 157.5000 ;
	    RECT 1374.6000 153.3000 1375.8000 156.3000 ;
	    RECT 1377.0000 153.3000 1378.2001 157.5000 ;
	    RECT 1379.4000 153.3000 1380.6000 157.5000 ;
	    RECT 1381.8000 153.3000 1383.0000 157.5000 ;
	    RECT 1384.2001 153.3000 1385.4000 157.5000 ;
	    RECT 1386.6000 153.3000 1387.8000 158.1000 ;
	    RECT 1391.4000 153.3000 1392.6000 159.3000 ;
	    RECT 1396.2001 153.3000 1397.4000 161.1000 ;
	    RECT 1398.9000 160.2000 1400.1000 166.8000 ;
	    RECT 1422.9000 163.5000 1423.8000 167.7000 ;
	    RECT 1444.2001 167.4000 1445.4000 168.6000 ;
	    RECT 1425.0000 166.5000 1426.2001 166.8000 ;
	    RECT 1446.6000 166.5000 1447.8000 179.7000 ;
	    RECT 1449.0000 173.7000 1450.2001 179.7000 ;
	    RECT 1425.0000 164.4000 1426.2001 165.6000 ;
	    RECT 1446.6000 165.4500 1447.8000 165.6000 ;
	    RECT 1461.0000 165.4500 1462.2001 165.6000 ;
	    RECT 1446.6000 164.5500 1462.2001 165.4500 ;
	    RECT 1446.6000 164.4000 1447.8000 164.5500 ;
	    RECT 1461.0000 164.4000 1462.2001 164.5500 ;
	    RECT 1463.4000 163.5000 1464.6000 179.7000 ;
	    RECT 1465.8000 173.7000 1467.0000 179.7000 ;
	    RECT 1492.2001 173.7000 1493.4000 179.7000 ;
	    RECT 1494.6000 173.7000 1495.8000 179.7000 ;
	    RECT 1497.0000 174.3000 1498.2001 179.7000 ;
	    RECT 1494.9000 173.4000 1495.8000 173.7000 ;
	    RECT 1499.4000 173.7000 1500.6000 179.7000 ;
	    RECT 1523.4000 173.7000 1524.6000 179.7000 ;
	    RECT 1525.8000 174.3000 1527.0000 179.7000 ;
	    RECT 1499.4000 173.4000 1500.3000 173.7000 ;
	    RECT 1494.9000 172.5000 1500.3000 173.4000 ;
	    RECT 1477.8000 171.4500 1479.0000 171.6000 ;
	    RECT 1497.0000 171.4500 1498.2001 171.6000 ;
	    RECT 1477.8000 170.5500 1498.2001 171.4500 ;
	    RECT 1477.8000 170.4000 1479.0000 170.5500 ;
	    RECT 1497.0000 170.4000 1498.2001 170.5500 ;
	    RECT 1499.4000 169.5000 1500.3000 172.5000 ;
	    RECT 1523.7001 173.4000 1524.6000 173.7000 ;
	    RECT 1528.2001 173.7000 1529.4000 179.7000 ;
	    RECT 1530.6000 173.7000 1531.8000 179.7000 ;
	    RECT 1554.6000 173.7000 1555.8000 179.7000 ;
	    RECT 1557.0000 173.7000 1558.2001 179.7000 ;
	    RECT 1559.4000 174.3000 1560.6000 179.7000 ;
	    RECT 1528.2001 173.4000 1529.1000 173.7000 ;
	    RECT 1523.7001 172.5000 1529.1000 173.4000 ;
	    RECT 1557.3000 173.4000 1558.2001 173.7000 ;
	    RECT 1561.8000 173.7000 1563.0000 179.7000 ;
	    RECT 1561.8000 173.4000 1562.7001 173.7000 ;
	    RECT 1557.3000 172.5000 1562.7001 173.4000 ;
	    RECT 1523.7001 169.5000 1524.6000 172.5000 ;
	    RECT 1525.8000 170.4000 1527.0000 171.6000 ;
	    RECT 1554.6000 171.4500 1555.8000 171.6000 ;
	    RECT 1559.4000 171.4500 1560.6000 171.6000 ;
	    RECT 1554.6000 170.5500 1560.6000 171.4500 ;
	    RECT 1554.6000 170.4000 1555.8000 170.5500 ;
	    RECT 1559.4000 170.4000 1560.6000 170.5500 ;
	    RECT 1561.8000 169.5000 1562.7001 172.5000 ;
	    RECT 1497.0000 169.2000 1498.2001 169.5000 ;
	    RECT 1525.8000 169.2000 1527.0000 169.5000 ;
	    RECT 1559.4000 169.2000 1560.6000 169.5000 ;
	    RECT 1473.0000 168.4500 1474.2001 168.6000 ;
	    RECT 1492.2001 168.4500 1493.4000 168.6000 ;
	    RECT 1473.0000 167.5500 1493.4000 168.4500 ;
	    RECT 1473.0000 167.4000 1474.2001 167.5500 ;
	    RECT 1492.2001 167.4000 1493.4000 167.5500 ;
	    RECT 1499.4000 167.4000 1500.6000 168.6000 ;
	    RECT 1518.6000 168.4500 1519.8000 168.6000 ;
	    RECT 1523.4000 168.4500 1524.6000 168.6000 ;
	    RECT 1518.6000 167.5500 1524.6000 168.4500 ;
	    RECT 1518.6000 167.4000 1519.8000 167.5500 ;
	    RECT 1523.4000 167.4000 1524.6000 167.5500 ;
	    RECT 1530.6000 167.4000 1531.8000 168.6000 ;
	    RECT 1542.6000 168.4500 1543.8000 168.6000 ;
	    RECT 1554.6000 168.4500 1555.8000 168.6000 ;
	    RECT 1542.6000 167.5500 1555.8000 168.4500 ;
	    RECT 1542.6000 167.4000 1543.8000 167.5500 ;
	    RECT 1554.6000 167.4000 1555.8000 167.5500 ;
	    RECT 1561.8000 167.4000 1563.0000 168.6000 ;
	    RECT 1492.2001 166.2000 1493.4000 166.5000 ;
	    RECT 1494.6000 164.4000 1495.8000 165.6000 ;
	    RECT 1496.7001 164.4000 1497.0000 165.6000 ;
	    RECT 1422.6000 162.4500 1423.8000 162.6000 ;
	    RECT 1444.2001 162.4500 1445.4000 162.6000 ;
	    RECT 1422.6000 161.5500 1445.4000 162.4500 ;
	    RECT 1422.6000 161.4000 1423.8000 161.5500 ;
	    RECT 1444.2001 161.4000 1445.4000 161.5500 ;
	    RECT 1398.6000 159.0000 1400.1000 160.2000 ;
	    RECT 1405.8000 159.4500 1407.0000 159.6000 ;
	    RECT 1420.2001 159.4500 1421.4000 159.6000 ;
	    RECT 1398.6000 153.3000 1399.8000 159.0000 ;
	    RECT 1405.8000 158.5500 1421.4000 159.4500 ;
	    RECT 1405.8000 158.4000 1407.0000 158.5500 ;
	    RECT 1420.2001 158.4000 1421.4000 158.5500 ;
	    RECT 1420.2001 157.2000 1421.4000 157.5000 ;
	    RECT 1422.9000 156.3000 1423.8000 160.5000 ;
	    RECT 1446.6000 159.3000 1447.8000 163.5000 ;
	    RECT 1499.4000 162.6000 1500.3000 166.5000 ;
	    RECT 1449.0000 162.4500 1450.2001 162.6000 ;
	    RECT 1453.8000 162.4500 1455.0000 162.6000 ;
	    RECT 1449.0000 161.5500 1455.0000 162.4500 ;
	    RECT 1449.0000 161.4000 1450.2001 161.5500 ;
	    RECT 1453.8000 161.4000 1455.0000 161.5500 ;
	    RECT 1463.4000 162.4500 1464.6000 162.6000 ;
	    RECT 1465.8000 162.4500 1467.0000 162.6000 ;
	    RECT 1463.4000 161.5500 1467.0000 162.4500 ;
	    RECT 1497.9000 162.3000 1500.3000 162.6000 ;
	    RECT 1463.4000 161.4000 1464.6000 161.5500 ;
	    RECT 1465.8000 161.4000 1467.0000 161.5500 ;
	    RECT 1449.0000 160.2000 1450.2001 160.5000 ;
	    RECT 1445.1000 158.4000 1447.8000 159.3000 ;
	    RECT 1401.0000 153.3000 1402.2001 156.3000 ;
	    RECT 1420.2001 153.3000 1421.4000 156.3000 ;
	    RECT 1422.6000 153.3000 1423.8000 156.3000 ;
	    RECT 1425.0000 153.3000 1426.2001 156.3000 ;
	    RECT 1445.1000 153.3000 1446.3000 158.4000 ;
	    RECT 1449.0000 153.3000 1450.2001 159.3000 ;
	    RECT 1463.4000 153.3000 1464.6000 160.5000 ;
	    RECT 1465.8000 159.4500 1467.0000 159.6000 ;
	    RECT 1468.2001 159.4500 1469.4000 159.6000 ;
	    RECT 1465.8000 158.5500 1469.4000 159.4500 ;
	    RECT 1465.8000 158.4000 1467.0000 158.5500 ;
	    RECT 1468.2001 158.4000 1469.4000 158.5500 ;
	    RECT 1465.8000 157.2000 1467.0000 157.5000 ;
	    RECT 1465.8000 153.3000 1467.0000 156.3000 ;
	    RECT 1492.2001 153.3000 1493.4000 162.3000 ;
	    RECT 1497.6000 161.7000 1500.3000 162.3000 ;
	    RECT 1523.7001 162.6000 1524.6000 166.5000 ;
	    RECT 1530.6000 166.2000 1531.8000 166.5000 ;
	    RECT 1554.6000 166.2000 1555.8000 166.5000 ;
	    RECT 1527.0000 164.4000 1527.3000 165.6000 ;
	    RECT 1528.2001 164.4000 1529.4000 165.6000 ;
	    RECT 1557.0000 164.4000 1558.2001 165.6000 ;
	    RECT 1559.1000 164.4000 1559.4000 165.6000 ;
	    RECT 1561.8000 162.6000 1562.7001 166.5000 ;
	    RECT 1523.7001 162.3000 1526.1000 162.6000 ;
	    RECT 1560.3000 162.3000 1562.7001 162.6000 ;
	    RECT 1523.7001 161.7000 1526.4000 162.3000 ;
	    RECT 1497.6000 153.3000 1498.8000 161.7000 ;
	    RECT 1525.2001 153.3000 1526.4000 161.7000 ;
	    RECT 1530.6000 153.3000 1531.8000 162.3000 ;
	    RECT 1554.6000 153.3000 1555.8000 162.3000 ;
	    RECT 1560.0000 161.7000 1562.7001 162.3000 ;
	    RECT 1560.0000 153.3000 1561.2001 161.7000 ;
	    RECT 1.2000 150.6000 1569.0000 152.4000 ;
	    RECT 126.6000 140.7000 127.8000 149.7000 ;
	    RECT 131.4000 143.7000 132.6000 149.7000 ;
	    RECT 136.2000 144.9000 137.4000 149.7000 ;
	    RECT 138.6000 145.5000 139.8000 149.7000 ;
	    RECT 141.0000 145.5000 142.2000 149.7000 ;
	    RECT 143.4000 145.5000 144.6000 149.7000 ;
	    RECT 145.8000 146.7000 147.0000 149.7000 ;
	    RECT 148.2000 145.5000 149.4000 149.7000 ;
	    RECT 150.6000 146.7000 151.8000 149.7000 ;
	    RECT 153.0000 145.5000 154.2000 149.7000 ;
	    RECT 155.4000 145.5000 156.6000 149.7000 ;
	    RECT 157.8000 145.5000 159.0000 149.7000 ;
	    RECT 160.2000 145.5000 161.4000 149.7000 ;
	    RECT 133.5000 143.7000 137.4000 144.9000 ;
	    RECT 162.6000 144.9000 163.8000 149.7000 ;
	    RECT 142.5000 143.7000 149.4000 144.6000 ;
	    RECT 133.5000 142.8000 134.7000 143.7000 ;
	    RECT 130.2000 141.6000 134.7000 142.8000 ;
	    RECT 126.6000 139.5000 139.8000 140.7000 ;
	    RECT 142.5000 140.1000 143.7000 143.7000 ;
	    RECT 148.2000 143.4000 149.4000 143.7000 ;
	    RECT 150.6000 143.4000 151.8000 144.6000 ;
	    RECT 152.7000 143.4000 153.0000 144.6000 ;
	    RECT 157.5000 143.4000 159.0000 144.6000 ;
	    RECT 162.6000 143.7000 166.2000 144.9000 ;
	    RECT 167.4000 143.7000 168.6000 149.7000 ;
	    RECT 145.8000 142.5000 147.0000 142.8000 ;
	    RECT 148.2000 142.2000 149.4000 142.5000 ;
	    RECT 145.8000 140.4000 147.0000 141.6000 ;
	    RECT 148.2000 141.3000 154.8000 142.2000 ;
	    RECT 153.6000 141.0000 154.8000 141.3000 ;
	    RECT 126.6000 131.1000 127.8000 139.5000 ;
	    RECT 140.7000 138.9000 143.7000 140.1000 ;
	    RECT 149.4000 138.9000 154.2000 140.1000 ;
	    RECT 157.8000 139.2000 159.0000 143.4000 ;
	    RECT 165.0000 142.8000 166.2000 143.7000 ;
	    RECT 165.0000 141.9000 167.7000 142.8000 ;
	    RECT 166.5000 140.1000 167.7000 141.9000 ;
	    RECT 172.2000 141.9000 173.4000 149.7000 ;
	    RECT 174.6000 144.0000 175.8000 149.7000 ;
	    RECT 177.0000 146.7000 178.2000 149.7000 ;
	    RECT 191.4000 146.7000 192.6000 149.7000 ;
	    RECT 191.4000 145.5000 192.6000 145.8000 ;
	    RECT 174.6000 142.8000 176.1000 144.0000 ;
	    RECT 191.4000 143.4000 192.6000 144.6000 ;
	    RECT 172.2000 141.0000 174.0000 141.9000 ;
	    RECT 166.5000 138.9000 172.2000 140.1000 ;
	    RECT 128.7000 138.0000 129.9000 138.3000 ;
	    RECT 128.7000 137.1000 135.3000 138.0000 ;
	    RECT 136.2000 137.4000 137.4000 138.6000 ;
	    RECT 162.6000 138.0000 163.8000 138.9000 ;
	    RECT 173.1000 138.0000 174.0000 141.0000 ;
	    RECT 138.3000 137.1000 163.8000 138.0000 ;
	    RECT 172.8000 137.1000 174.0000 138.0000 ;
	    RECT 170.7000 136.2000 171.9000 136.5000 ;
	    RECT 131.4000 134.4000 132.6000 135.6000 ;
	    RECT 133.5000 135.3000 171.9000 136.2000 ;
	    RECT 136.5000 135.0000 137.7000 135.3000 ;
	    RECT 172.8000 134.4000 173.7000 137.1000 ;
	    RECT 174.9000 136.2000 176.1000 142.8000 ;
	    RECT 193.8000 142.5000 195.0000 149.7000 ;
	    RECT 193.8000 141.4500 195.0000 141.6000 ;
	    RECT 280.2000 141.4500 281.4000 141.6000 ;
	    RECT 193.8000 140.5500 281.4000 141.4500 ;
	    RECT 193.8000 140.4000 195.0000 140.5500 ;
	    RECT 280.2000 140.4000 281.4000 140.5500 ;
	    RECT 328.2000 140.7000 329.4000 149.7000 ;
	    RECT 333.0000 143.7000 334.2000 149.7000 ;
	    RECT 337.8000 144.9000 339.0000 149.7000 ;
	    RECT 340.2000 145.5000 341.4000 149.7000 ;
	    RECT 342.6000 145.5000 343.8000 149.7000 ;
	    RECT 345.0000 145.5000 346.2000 149.7000 ;
	    RECT 347.4000 146.7000 348.6000 149.7000 ;
	    RECT 349.8000 145.5000 351.0000 149.7000 ;
	    RECT 352.2000 146.7000 353.4000 149.7000 ;
	    RECT 354.6000 145.5000 355.8000 149.7000 ;
	    RECT 357.0000 145.5000 358.2000 149.7000 ;
	    RECT 359.4000 145.5000 360.6000 149.7000 ;
	    RECT 361.8000 145.5000 363.0000 149.7000 ;
	    RECT 335.1000 143.7000 339.0000 144.9000 ;
	    RECT 364.2000 144.9000 365.4000 149.7000 ;
	    RECT 344.1000 143.7000 351.0000 144.6000 ;
	    RECT 335.1000 142.8000 336.3000 143.7000 ;
	    RECT 331.8000 141.6000 336.3000 142.8000 ;
	    RECT 328.2000 139.5000 341.4000 140.7000 ;
	    RECT 344.1000 140.1000 345.3000 143.7000 ;
	    RECT 349.8000 143.4000 351.0000 143.7000 ;
	    RECT 352.2000 143.4000 353.4000 144.6000 ;
	    RECT 354.3000 143.4000 354.6000 144.6000 ;
	    RECT 359.1000 143.4000 360.6000 144.6000 ;
	    RECT 364.2000 143.7000 367.8000 144.9000 ;
	    RECT 369.0000 143.7000 370.2000 149.7000 ;
	    RECT 347.4000 142.5000 348.6000 142.8000 ;
	    RECT 349.8000 142.2000 351.0000 142.5000 ;
	    RECT 347.4000 140.4000 348.6000 141.6000 ;
	    RECT 349.8000 141.3000 356.4000 142.2000 ;
	    RECT 355.2000 141.0000 356.4000 141.3000 ;
	    RECT 141.0000 134.1000 142.2000 134.4000 ;
	    RECT 134.1000 133.5000 142.2000 134.1000 ;
	    RECT 132.9000 133.2000 142.2000 133.5000 ;
	    RECT 143.7000 133.5000 156.6000 134.4000 ;
	    RECT 129.0000 132.0000 131.4000 133.2000 ;
	    RECT 132.9000 132.3000 135.0000 133.2000 ;
	    RECT 143.7000 132.3000 144.6000 133.5000 ;
	    RECT 155.4000 133.2000 156.6000 133.5000 ;
	    RECT 160.2000 133.5000 173.7000 134.4000 ;
	    RECT 174.6000 135.0000 176.1000 136.2000 ;
	    RECT 174.6000 133.5000 175.8000 135.0000 ;
	    RECT 160.2000 133.2000 161.4000 133.5000 ;
	    RECT 130.5000 131.4000 131.4000 132.0000 ;
	    RECT 135.9000 131.4000 144.6000 132.3000 ;
	    RECT 145.5000 131.4000 149.4000 132.6000 ;
	    RECT 126.6000 130.2000 129.6000 131.1000 ;
	    RECT 130.5000 130.2000 136.8000 131.4000 ;
	    RECT 128.7000 129.3000 129.6000 130.2000 ;
	    RECT 126.6000 123.3000 127.8000 129.3000 ;
	    RECT 128.7000 128.4000 130.2000 129.3000 ;
	    RECT 129.0000 123.3000 130.2000 128.4000 ;
	    RECT 131.4000 122.4000 132.6000 129.3000 ;
	    RECT 133.8000 123.3000 135.0000 130.2000 ;
	    RECT 136.2000 123.3000 137.4000 129.3000 ;
	    RECT 138.6000 123.3000 139.8000 127.5000 ;
	    RECT 141.0000 123.3000 142.2000 127.5000 ;
	    RECT 143.4000 123.3000 144.6000 130.5000 ;
	    RECT 145.8000 123.3000 147.0000 129.3000 ;
	    RECT 148.2000 123.3000 149.4000 130.5000 ;
	    RECT 150.6000 123.3000 151.8000 129.3000 ;
	    RECT 153.0000 123.3000 154.2000 132.6000 ;
	    RECT 165.0000 131.4000 168.9000 132.6000 ;
	    RECT 157.8000 130.2000 164.1000 131.4000 ;
	    RECT 155.4000 123.3000 156.6000 127.5000 ;
	    RECT 157.8000 123.3000 159.0000 127.5000 ;
	    RECT 160.2000 123.3000 161.4000 127.5000 ;
	    RECT 162.6000 123.3000 163.8000 129.3000 ;
	    RECT 165.0000 123.3000 166.2000 131.4000 ;
	    RECT 172.8000 131.1000 173.7000 133.5000 ;
	    RECT 174.6000 131.4000 175.8000 132.6000 ;
	    RECT 169.8000 130.2000 173.7000 131.1000 ;
	    RECT 167.4000 123.3000 168.6000 129.3000 ;
	    RECT 169.8000 123.3000 171.0000 130.2000 ;
	    RECT 172.2000 123.3000 173.4000 129.3000 ;
	    RECT 174.6000 123.3000 175.8000 130.5000 ;
	    RECT 177.0000 123.3000 178.2000 129.3000 ;
	    RECT 191.4000 123.3000 192.6000 129.3000 ;
	    RECT 193.8000 123.3000 195.0000 139.5000 ;
	    RECT 222.6000 138.4500 223.8000 138.6000 ;
	    RECT 321.0000 138.4500 322.2000 138.6000 ;
	    RECT 222.6000 137.5500 322.2000 138.4500 ;
	    RECT 222.6000 137.4000 223.8000 137.5500 ;
	    RECT 321.0000 137.4000 322.2000 137.5500 ;
	    RECT 328.2000 131.1000 329.4000 139.5000 ;
	    RECT 342.3000 138.9000 345.3000 140.1000 ;
	    RECT 351.0000 138.9000 355.8000 140.1000 ;
	    RECT 359.4000 139.2000 360.6000 143.4000 ;
	    RECT 366.6000 142.8000 367.8000 143.7000 ;
	    RECT 366.6000 141.9000 369.3000 142.8000 ;
	    RECT 368.1000 140.1000 369.3000 141.9000 ;
	    RECT 373.8000 141.9000 375.0000 149.7000 ;
	    RECT 376.2000 144.0000 377.4000 149.7000 ;
	    RECT 378.6000 146.7000 379.8000 149.7000 ;
	    RECT 376.2000 142.8000 377.7000 144.0000 ;
	    RECT 373.8000 141.0000 375.6000 141.9000 ;
	    RECT 368.1000 138.9000 373.8000 140.1000 ;
	    RECT 330.3000 138.0000 331.5000 138.3000 ;
	    RECT 330.3000 137.1000 336.9000 138.0000 ;
	    RECT 337.8000 137.4000 339.0000 138.6000 ;
	    RECT 364.2000 138.0000 365.4000 138.9000 ;
	    RECT 374.7000 138.0000 375.6000 141.0000 ;
	    RECT 339.9000 137.1000 365.4000 138.0000 ;
	    RECT 374.4000 137.1000 375.6000 138.0000 ;
	    RECT 372.3000 136.2000 373.5000 136.5000 ;
	    RECT 333.0000 134.4000 334.2000 135.6000 ;
	    RECT 335.1000 135.3000 373.5000 136.2000 ;
	    RECT 338.1000 135.0000 339.3000 135.3000 ;
	    RECT 374.4000 134.4000 375.3000 137.1000 ;
	    RECT 376.5000 136.2000 377.7000 142.8000 ;
	    RECT 393.0000 142.5000 394.2000 149.7000 ;
	    RECT 395.4000 146.7000 396.6000 149.7000 ;
	    RECT 395.4000 145.5000 396.6000 145.8000 ;
	    RECT 395.4000 144.4500 396.6000 144.6000 ;
	    RECT 424.2000 144.4500 425.4000 144.6000 ;
	    RECT 395.4000 143.5500 425.4000 144.4500 ;
	    RECT 395.4000 143.4000 396.6000 143.5500 ;
	    RECT 424.2000 143.4000 425.4000 143.5500 ;
	    RECT 393.0000 141.4500 394.2000 141.6000 ;
	    RECT 460.2000 141.4500 461.4000 141.6000 ;
	    RECT 393.0000 140.5500 461.4000 141.4500 ;
	    RECT 393.0000 140.4000 394.2000 140.5500 ;
	    RECT 460.2000 140.4000 461.4000 140.5500 ;
	    RECT 527.4000 140.7000 528.6000 149.7000 ;
	    RECT 532.2000 143.7000 533.4000 149.7000 ;
	    RECT 537.0000 144.9000 538.2000 149.7000 ;
	    RECT 539.4000 145.5000 540.6000 149.7000 ;
	    RECT 541.8000 145.5000 543.0000 149.7000 ;
	    RECT 544.2000 145.5000 545.4000 149.7000 ;
	    RECT 546.6000 146.7000 547.8000 149.7000 ;
	    RECT 549.0000 145.5000 550.2000 149.7000 ;
	    RECT 551.4000 146.7000 552.6000 149.7000 ;
	    RECT 553.8000 145.5000 555.0000 149.7000 ;
	    RECT 556.2000 145.5000 557.4000 149.7000 ;
	    RECT 558.6000 145.5000 559.8000 149.7000 ;
	    RECT 561.0000 145.5000 562.2000 149.7000 ;
	    RECT 534.3000 143.7000 538.2000 144.9000 ;
	    RECT 563.4000 144.9000 564.6000 149.7000 ;
	    RECT 543.3000 143.7000 550.2000 144.6000 ;
	    RECT 534.3000 142.8000 535.5000 143.7000 ;
	    RECT 531.0000 141.6000 535.5000 142.8000 ;
	    RECT 527.4000 139.5000 540.6000 140.7000 ;
	    RECT 543.3000 140.1000 544.5000 143.7000 ;
	    RECT 549.0000 143.4000 550.2000 143.7000 ;
	    RECT 551.4000 143.4000 552.6000 144.6000 ;
	    RECT 553.5000 143.4000 553.8000 144.6000 ;
	    RECT 558.3000 143.4000 559.8000 144.6000 ;
	    RECT 563.4000 143.7000 567.0000 144.9000 ;
	    RECT 568.2000 143.7000 569.4000 149.7000 ;
	    RECT 546.6000 142.5000 547.8000 142.8000 ;
	    RECT 549.0000 142.2000 550.2000 142.5000 ;
	    RECT 546.6000 140.4000 547.8000 141.6000 ;
	    RECT 549.0000 141.3000 555.6000 142.2000 ;
	    RECT 554.4000 141.0000 555.6000 141.3000 ;
	    RECT 342.6000 134.1000 343.8000 134.4000 ;
	    RECT 335.7000 133.5000 343.8000 134.1000 ;
	    RECT 334.5000 133.2000 343.8000 133.5000 ;
	    RECT 345.3000 133.5000 358.2000 134.4000 ;
	    RECT 330.6000 132.0000 333.0000 133.2000 ;
	    RECT 334.5000 132.3000 336.6000 133.2000 ;
	    RECT 345.3000 132.3000 346.2000 133.5000 ;
	    RECT 357.0000 133.2000 358.2000 133.5000 ;
	    RECT 361.8000 133.5000 375.3000 134.4000 ;
	    RECT 376.2000 135.0000 377.7000 136.2000 ;
	    RECT 376.2000 133.5000 377.4000 135.0000 ;
	    RECT 361.8000 133.2000 363.0000 133.5000 ;
	    RECT 332.1000 131.4000 333.0000 132.0000 ;
	    RECT 337.5000 131.4000 346.2000 132.3000 ;
	    RECT 347.1000 131.4000 351.0000 132.6000 ;
	    RECT 328.2000 130.2000 331.2000 131.1000 ;
	    RECT 332.1000 130.2000 338.4000 131.4000 ;
	    RECT 270.6000 129.4500 271.8000 129.6000 ;
	    RECT 292.2000 129.4500 293.4000 129.6000 ;
	    RECT 270.6000 128.5500 293.4000 129.4500 ;
	    RECT 330.3000 129.3000 331.2000 130.2000 ;
	    RECT 270.6000 128.4000 271.8000 128.5500 ;
	    RECT 292.2000 128.4000 293.4000 128.5500 ;
	    RECT 215.4000 126.4500 216.6000 126.6000 ;
	    RECT 277.8000 126.4500 279.0000 126.6000 ;
	    RECT 215.4000 125.5500 279.0000 126.4500 ;
	    RECT 215.4000 125.4000 216.6000 125.5500 ;
	    RECT 277.8000 125.4000 279.0000 125.5500 ;
	    RECT 328.2000 123.3000 329.4000 129.3000 ;
	    RECT 330.3000 128.4000 331.8000 129.3000 ;
	    RECT 330.6000 123.3000 331.8000 128.4000 ;
	    RECT 333.0000 122.4000 334.2000 129.3000 ;
	    RECT 335.4000 123.3000 336.6000 130.2000 ;
	    RECT 337.8000 123.3000 339.0000 129.3000 ;
	    RECT 340.2000 123.3000 341.4000 127.5000 ;
	    RECT 342.6000 123.3000 343.8000 127.5000 ;
	    RECT 345.0000 123.3000 346.2000 130.5000 ;
	    RECT 347.4000 123.3000 348.6000 129.3000 ;
	    RECT 349.8000 123.3000 351.0000 130.5000 ;
	    RECT 352.2000 123.3000 353.4000 129.3000 ;
	    RECT 354.6000 123.3000 355.8000 132.6000 ;
	    RECT 366.6000 131.4000 370.5000 132.6000 ;
	    RECT 359.4000 130.2000 365.7000 131.4000 ;
	    RECT 357.0000 123.3000 358.2000 127.5000 ;
	    RECT 359.4000 123.3000 360.6000 127.5000 ;
	    RECT 361.8000 123.3000 363.0000 127.5000 ;
	    RECT 364.2000 123.3000 365.4000 129.3000 ;
	    RECT 366.6000 123.3000 367.8000 131.4000 ;
	    RECT 374.4000 131.1000 375.3000 133.5000 ;
	    RECT 376.2000 131.4000 377.4000 132.6000 ;
	    RECT 371.4000 130.2000 375.3000 131.1000 ;
	    RECT 369.0000 123.3000 370.2000 129.3000 ;
	    RECT 371.4000 123.3000 372.6000 130.2000 ;
	    RECT 373.8000 123.3000 375.0000 129.3000 ;
	    RECT 376.2000 123.3000 377.4000 130.5000 ;
	    RECT 378.6000 123.3000 379.8000 129.3000 ;
	    RECT 393.0000 123.3000 394.2000 139.5000 ;
	    RECT 527.4000 131.1000 528.6000 139.5000 ;
	    RECT 541.5000 138.9000 544.5000 140.1000 ;
	    RECT 550.2000 138.9000 555.0000 140.1000 ;
	    RECT 558.6000 139.2000 559.8000 143.4000 ;
	    RECT 565.8000 142.8000 567.0000 143.7000 ;
	    RECT 565.8000 141.9000 568.5000 142.8000 ;
	    RECT 567.3000 140.1000 568.5000 141.9000 ;
	    RECT 573.0000 141.9000 574.2000 149.7000 ;
	    RECT 575.4000 144.0000 576.6000 149.7000 ;
	    RECT 577.8000 146.7000 579.0000 149.7000 ;
	    RECT 575.4000 142.8000 576.9000 144.0000 ;
	    RECT 597.0000 143.7000 598.2000 149.7000 ;
	    RECT 600.9000 144.6000 602.1000 149.7000 ;
	    RECT 621.0000 146.7000 622.2000 149.7000 ;
	    RECT 623.4000 146.7000 624.6000 149.7000 ;
	    RECT 625.8000 146.7000 627.0000 149.7000 ;
	    RECT 621.0000 145.5000 622.2000 145.8000 ;
	    RECT 599.4000 143.7000 602.1000 144.6000 ;
	    RECT 613.8000 144.4500 615.0000 144.6000 ;
	    RECT 621.0000 144.4500 622.2000 144.6000 ;
	    RECT 573.0000 141.0000 574.8000 141.9000 ;
	    RECT 567.3000 138.9000 573.0000 140.1000 ;
	    RECT 529.5000 138.0000 530.7000 138.3000 ;
	    RECT 529.5000 137.1000 536.1000 138.0000 ;
	    RECT 537.0000 137.4000 538.2000 138.6000 ;
	    RECT 563.4000 138.0000 564.6000 138.9000 ;
	    RECT 573.9000 138.0000 574.8000 141.0000 ;
	    RECT 539.1000 137.1000 564.6000 138.0000 ;
	    RECT 573.6000 137.1000 574.8000 138.0000 ;
	    RECT 571.5000 136.2000 572.7000 136.5000 ;
	    RECT 532.2000 134.4000 533.4000 135.6000 ;
	    RECT 534.3000 135.3000 572.7000 136.2000 ;
	    RECT 537.3000 135.0000 538.5000 135.3000 ;
	    RECT 573.6000 134.4000 574.5000 137.1000 ;
	    RECT 575.7000 136.2000 576.9000 142.8000 ;
	    RECT 597.0000 142.5000 598.2000 142.8000 ;
	    RECT 580.2000 141.4500 581.4000 141.6000 ;
	    RECT 597.0000 141.4500 598.2000 141.6000 ;
	    RECT 580.2000 140.5500 598.2000 141.4500 ;
	    RECT 580.2000 140.4000 581.4000 140.5500 ;
	    RECT 597.0000 140.4000 598.2000 140.5500 ;
	    RECT 599.4000 139.5000 600.6000 143.7000 ;
	    RECT 613.8000 143.5500 622.2000 144.4500 ;
	    RECT 613.8000 143.4000 615.0000 143.5500 ;
	    RECT 621.0000 143.4000 622.2000 143.5500 ;
	    RECT 623.7000 142.5000 624.6000 146.7000 ;
	    RECT 702.6000 143.1000 703.8000 149.7000 ;
	    RECT 705.0000 144.0000 706.2000 149.7000 ;
	    RECT 708.9000 147.6000 710.7000 149.7000 ;
	    RECT 708.9000 146.7000 711.0000 147.6000 ;
	    RECT 713.4000 146.7000 714.6000 149.7000 ;
	    RECT 715.8000 146.7000 717.0000 149.7000 ;
	    RECT 718.2000 146.7000 719.7000 149.7000 ;
	    RECT 722.4000 147.6000 723.6000 149.7000 ;
	    RECT 722.4000 146.7000 725.4000 147.6000 ;
	    RECT 709.8000 145.5000 711.0000 146.7000 ;
	    RECT 716.1000 145.8000 717.0000 146.7000 ;
	    RECT 716.1000 144.9000 720.3000 145.8000 ;
	    RECT 719.1000 144.6000 720.3000 144.9000 ;
	    RECT 721.8000 144.6000 723.0000 145.8000 ;
	    RECT 724.2000 145.5000 725.4000 146.7000 ;
	    RECT 707.1000 143.1000 708.3000 143.4000 ;
	    RECT 702.6000 142.2000 708.3000 143.1000 ;
	    RECT 623.4000 141.4500 624.6000 141.6000 ;
	    RECT 700.2000 141.4500 701.4000 141.6000 ;
	    RECT 623.4000 140.5500 701.4000 141.4500 ;
	    RECT 623.4000 140.4000 624.6000 140.5500 ;
	    RECT 700.2000 140.4000 701.4000 140.5500 ;
	    RECT 702.6000 139.5000 703.8000 142.2000 ;
	    RECT 713.1000 141.3000 714.3000 141.6000 ;
	    RECT 721.8000 141.3000 722.7000 144.6000 ;
	    RECT 726.6000 143.7000 727.8000 149.7000 ;
	    RECT 729.0000 142.5000 730.2000 149.7000 ;
	    RECT 798.6000 143.1000 799.8000 149.7000 ;
	    RECT 801.0000 144.0000 802.2000 149.7000 ;
	    RECT 804.9000 147.6000 806.7000 149.7000 ;
	    RECT 804.9000 146.7000 807.0000 147.6000 ;
	    RECT 809.4000 146.7000 810.6000 149.7000 ;
	    RECT 811.8000 146.7000 813.0000 149.7000 ;
	    RECT 814.2000 146.7000 815.7000 149.7000 ;
	    RECT 818.4000 147.6000 819.6000 149.7000 ;
	    RECT 818.4000 146.7000 821.4000 147.6000 ;
	    RECT 805.8000 145.5000 807.0000 146.7000 ;
	    RECT 812.1000 145.8000 813.0000 146.7000 ;
	    RECT 812.1000 144.9000 816.3000 145.8000 ;
	    RECT 815.1000 144.6000 816.3000 144.9000 ;
	    RECT 817.8000 144.6000 819.0000 145.8000 ;
	    RECT 820.2000 145.5000 821.4000 146.7000 ;
	    RECT 803.1000 143.1000 804.3000 143.4000 ;
	    RECT 798.6000 142.2000 804.3000 143.1000 ;
	    RECT 712.5000 140.4000 725.7000 141.3000 ;
	    RECT 726.6000 140.4000 727.8000 141.6000 ;
	    RECT 728.7000 140.4000 729.0000 141.6000 ;
	    RECT 599.4000 138.4500 600.6000 138.6000 ;
	    RECT 621.0000 138.4500 622.2000 138.6000 ;
	    RECT 599.4000 137.5500 622.2000 138.4500 ;
	    RECT 599.4000 137.4000 600.6000 137.5500 ;
	    RECT 621.0000 137.4000 622.2000 137.5500 ;
	    RECT 541.8000 134.1000 543.0000 134.4000 ;
	    RECT 534.9000 133.5000 543.0000 134.1000 ;
	    RECT 533.7000 133.2000 543.0000 133.5000 ;
	    RECT 544.5000 133.5000 557.4000 134.4000 ;
	    RECT 529.8000 132.0000 532.2000 133.2000 ;
	    RECT 533.7000 132.3000 535.8000 133.2000 ;
	    RECT 544.5000 132.3000 545.4000 133.5000 ;
	    RECT 556.2000 133.2000 557.4000 133.5000 ;
	    RECT 561.0000 133.5000 574.5000 134.4000 ;
	    RECT 575.4000 135.0000 576.9000 136.2000 ;
	    RECT 575.4000 133.5000 576.6000 135.0000 ;
	    RECT 561.0000 133.2000 562.2000 133.5000 ;
	    RECT 531.3000 131.4000 532.2000 132.0000 ;
	    RECT 536.7000 131.4000 545.4000 132.3000 ;
	    RECT 546.3000 131.4000 550.2000 132.6000 ;
	    RECT 527.4000 130.2000 530.4000 131.1000 ;
	    RECT 531.3000 130.2000 537.6000 131.4000 ;
	    RECT 529.5000 129.3000 530.4000 130.2000 ;
	    RECT 395.4000 123.3000 396.6000 129.3000 ;
	    RECT 527.4000 123.3000 528.6000 129.3000 ;
	    RECT 529.5000 128.4000 531.0000 129.3000 ;
	    RECT 529.8000 123.3000 531.0000 128.4000 ;
	    RECT 532.2000 122.4000 533.4000 129.3000 ;
	    RECT 534.6000 123.3000 535.8000 130.2000 ;
	    RECT 537.0000 123.3000 538.2000 129.3000 ;
	    RECT 539.4000 123.3000 540.6000 127.5000 ;
	    RECT 541.8000 123.3000 543.0000 127.5000 ;
	    RECT 544.2000 123.3000 545.4000 130.5000 ;
	    RECT 546.6000 123.3000 547.8000 129.3000 ;
	    RECT 549.0000 123.3000 550.2000 130.5000 ;
	    RECT 551.4000 123.3000 552.6000 129.3000 ;
	    RECT 553.8000 123.3000 555.0000 132.6000 ;
	    RECT 565.8000 131.4000 569.7000 132.6000 ;
	    RECT 558.6000 130.2000 564.9000 131.4000 ;
	    RECT 556.2000 123.3000 557.4000 127.5000 ;
	    RECT 558.6000 123.3000 559.8000 127.5000 ;
	    RECT 561.0000 123.3000 562.2000 127.5000 ;
	    RECT 563.4000 123.3000 564.6000 129.3000 ;
	    RECT 565.8000 123.3000 567.0000 131.4000 ;
	    RECT 573.6000 131.1000 574.5000 133.5000 ;
	    RECT 575.4000 131.4000 576.6000 132.6000 ;
	    RECT 570.6000 130.2000 574.5000 131.1000 ;
	    RECT 568.2000 123.3000 569.4000 129.3000 ;
	    RECT 570.6000 123.3000 571.8000 130.2000 ;
	    RECT 573.0000 123.3000 574.2000 129.3000 ;
	    RECT 575.4000 123.3000 576.6000 130.5000 ;
	    RECT 577.8000 123.3000 579.0000 129.3000 ;
	    RECT 597.0000 123.3000 598.2000 129.3000 ;
	    RECT 599.4000 123.3000 600.6000 136.5000 ;
	    RECT 601.8000 135.4500 603.0000 135.6000 ;
	    RECT 609.0000 135.4500 610.2000 135.6000 ;
	    RECT 601.8000 134.5500 610.2000 135.4500 ;
	    RECT 623.7000 135.3000 624.6000 139.5000 ;
	    RECT 709.8000 139.2000 711.0000 139.5000 ;
	    RECT 625.8000 137.4000 627.0000 138.6000 ;
	    RECT 676.2000 138.4500 677.4000 138.6000 ;
	    RECT 702.6000 138.4500 703.8000 138.6000 ;
	    RECT 676.2000 137.5500 703.8000 138.4500 ;
	    RECT 705.3000 138.3000 711.0000 139.2000 ;
	    RECT 705.3000 138.0000 706.5000 138.3000 ;
	    RECT 676.2000 137.4000 677.4000 137.5500 ;
	    RECT 702.6000 137.4000 703.8000 137.5500 ;
	    RECT 707.7000 137.1000 708.9000 137.4000 ;
	    RECT 704.7000 136.5000 708.9000 137.1000 ;
	    RECT 625.8000 136.2000 627.0000 136.5000 ;
	    RECT 702.6000 136.2000 708.9000 136.5000 ;
	    RECT 601.8000 134.4000 603.0000 134.5500 ;
	    RECT 609.0000 134.4000 610.2000 134.5500 ;
	    RECT 601.8000 133.2000 603.0000 133.5000 ;
	    RECT 601.8000 123.3000 603.0000 129.3000 ;
	    RECT 621.0000 123.3000 622.2000 135.3000 ;
	    RECT 623.4000 134.1000 626.1000 135.3000 ;
	    RECT 624.9000 123.3000 626.1000 134.1000 ;
	    RECT 702.6000 123.3000 703.8000 136.2000 ;
	    RECT 712.5000 135.6000 713.4000 140.4000 ;
	    RECT 723.3000 140.1000 724.5000 140.4000 ;
	    RECT 798.6000 139.5000 799.8000 142.2000 ;
	    RECT 809.1000 141.3000 810.3000 141.6000 ;
	    RECT 817.8000 141.3000 818.7000 144.6000 ;
	    RECT 822.6000 143.7000 823.8000 149.7000 ;
	    RECT 825.0000 142.5000 826.2000 149.7000 ;
	    RECT 851.4000 144.0000 852.6000 149.7000 ;
	    RECT 853.8000 144.9000 855.0000 149.7000 ;
	    RECT 856.2000 144.0000 857.4000 149.7000 ;
	    RECT 851.4000 143.7000 857.4000 144.0000 ;
	    RECT 858.6000 143.7000 859.8000 149.7000 ;
	    RECT 851.7000 143.1000 857.1000 143.7000 ;
	    RECT 858.6000 142.5000 859.5000 143.7000 ;
	    RECT 870.6000 142.5000 871.8000 149.7000 ;
	    RECT 873.0000 146.7000 874.2000 149.7000 ;
	    RECT 873.0000 145.5000 874.2000 145.8000 ;
	    RECT 873.0000 144.4500 874.2000 144.6000 ;
	    RECT 935.4000 144.4500 936.6000 144.6000 ;
	    RECT 873.0000 143.5500 936.6000 144.4500 ;
	    RECT 873.0000 143.4000 874.2000 143.5500 ;
	    RECT 935.4000 143.4000 936.6000 143.5500 ;
	    RECT 808.5000 140.4000 821.7000 141.3000 ;
	    RECT 822.6000 140.4000 823.8000 141.6000 ;
	    RECT 824.7000 140.4000 825.0000 141.6000 ;
	    RECT 832.2000 141.4500 833.4000 141.6000 ;
	    RECT 851.4000 141.4500 852.6000 141.6000 ;
	    RECT 832.2000 140.5500 852.6000 141.4500 ;
	    RECT 853.5000 140.7000 853.8000 142.2000 ;
	    RECT 832.2000 140.4000 833.4000 140.5500 ;
	    RECT 851.4000 140.4000 852.6000 140.5500 ;
	    RECT 855.9000 140.4000 857.7000 141.6000 ;
	    RECT 858.6000 140.4000 859.8000 141.6000 ;
	    RECT 861.0000 141.4500 862.2000 141.6000 ;
	    RECT 870.6000 141.4500 871.8000 141.6000 ;
	    RECT 861.0000 140.5500 871.8000 141.4500 ;
	    RECT 861.0000 140.4000 862.2000 140.5500 ;
	    RECT 870.6000 140.4000 871.8000 140.5500 ;
	    RECT 1005.0000 140.7000 1006.2000 149.7000 ;
	    RECT 1009.8000 143.7000 1011.0000 149.7000 ;
	    RECT 1014.6000 144.9000 1015.8000 149.7000 ;
	    RECT 1017.0000 145.5000 1018.2000 149.7000 ;
	    RECT 1019.4000 145.5000 1020.6000 149.7000 ;
	    RECT 1021.8000 145.5000 1023.0000 149.7000 ;
	    RECT 1024.2001 146.7000 1025.4000 149.7000 ;
	    RECT 1026.6000 145.5000 1027.8000 149.7000 ;
	    RECT 1029.0000 146.7000 1030.2001 149.7000 ;
	    RECT 1031.4000 145.5000 1032.6000 149.7000 ;
	    RECT 1033.8000 145.5000 1035.0000 149.7000 ;
	    RECT 1036.2001 145.5000 1037.4000 149.7000 ;
	    RECT 1038.6000 145.5000 1039.8000 149.7000 ;
	    RECT 1011.9000 143.7000 1015.8000 144.9000 ;
	    RECT 1041.0000 144.9000 1042.2001 149.7000 ;
	    RECT 1020.9000 143.7000 1027.8000 144.6000 ;
	    RECT 1011.9000 142.8000 1013.1000 143.7000 ;
	    RECT 1008.6000 141.6000 1013.1000 142.8000 ;
	    RECT 805.8000 139.2000 807.0000 139.5000 ;
	    RECT 725.7000 138.6000 726.9000 138.9000 ;
	    RECT 719.4000 137.4000 720.6000 138.6000 ;
	    RECT 721.5000 137.7000 726.9000 138.6000 ;
	    RECT 779.4000 138.4500 780.6000 138.6000 ;
	    RECT 798.6000 138.4500 799.8000 138.6000 ;
	    RECT 779.4000 137.5500 799.8000 138.4500 ;
	    RECT 801.3000 138.3000 807.0000 139.2000 ;
	    RECT 801.3000 138.0000 802.5000 138.3000 ;
	    RECT 779.4000 137.4000 780.6000 137.5500 ;
	    RECT 798.6000 137.4000 799.8000 137.5500 ;
	    RECT 803.7000 137.1000 804.9000 137.4000 ;
	    RECT 721.8000 136.5000 730.2000 136.8000 ;
	    RECT 800.7000 136.5000 804.9000 137.1000 ;
	    RECT 721.5000 136.2000 730.2000 136.5000 ;
	    RECT 705.0000 123.3000 706.2000 135.3000 ;
	    RECT 709.8000 134.7000 713.4000 135.6000 ;
	    RECT 715.5000 135.9000 730.2000 136.2000 ;
	    RECT 715.5000 135.3000 722.7000 135.9000 ;
	    RECT 709.8000 133.2000 710.7000 134.7000 ;
	    RECT 708.6000 132.0000 710.7000 133.2000 ;
	    RECT 713.1000 133.5000 714.3000 133.8000 ;
	    RECT 715.5000 133.5000 716.4000 135.3000 ;
	    RECT 713.1000 132.6000 716.4000 133.5000 ;
	    RECT 717.3000 133.5000 725.4000 134.4000 ;
	    RECT 717.3000 133.2000 718.5000 133.5000 ;
	    RECT 724.2000 133.2000 725.4000 133.5000 ;
	    RECT 714.9000 131.1000 716.1000 131.4000 ;
	    RECT 719.1000 131.1000 720.3000 131.4000 ;
	    RECT 709.8000 129.3000 711.0000 130.5000 ;
	    RECT 714.9000 130.2000 720.3000 131.1000 ;
	    RECT 716.1000 129.3000 717.0000 130.2000 ;
	    RECT 724.2000 129.3000 725.4000 130.5000 ;
	    RECT 708.9000 123.3000 710.7000 129.3000 ;
	    RECT 713.4000 123.3000 714.6000 129.3000 ;
	    RECT 715.8000 123.3000 717.0000 129.3000 ;
	    RECT 718.2000 123.3000 719.4000 129.3000 ;
	    RECT 722.4000 128.4000 725.4000 129.3000 ;
	    RECT 722.4000 123.3000 723.6000 128.4000 ;
	    RECT 726.6000 123.3000 727.8000 135.0000 ;
	    RECT 729.0000 123.3000 730.2000 135.9000 ;
	    RECT 798.6000 136.2000 804.9000 136.5000 ;
	    RECT 798.6000 123.3000 799.8000 136.2000 ;
	    RECT 808.5000 135.6000 809.4000 140.4000 ;
	    RECT 819.3000 140.1000 820.5000 140.4000 ;
	    RECT 853.8000 139.5000 855.0000 139.8000 ;
	    RECT 821.7000 138.6000 822.9000 138.9000 ;
	    RECT 815.4000 137.4000 816.6000 138.6000 ;
	    RECT 817.5000 137.7000 822.9000 138.6000 ;
	    RECT 853.8000 137.4000 855.0000 138.6000 ;
	    RECT 817.8000 136.5000 826.2000 136.8000 ;
	    RECT 817.5000 136.2000 826.2000 136.5000 ;
	    RECT 801.0000 123.3000 802.2000 135.3000 ;
	    RECT 805.8000 134.7000 809.4000 135.6000 ;
	    RECT 811.5000 135.9000 826.2000 136.2000 ;
	    RECT 811.5000 135.3000 818.7000 135.9000 ;
	    RECT 805.8000 133.2000 806.7000 134.7000 ;
	    RECT 804.6000 132.0000 806.7000 133.2000 ;
	    RECT 809.1000 133.5000 810.3000 133.8000 ;
	    RECT 811.5000 133.5000 812.4000 135.3000 ;
	    RECT 809.1000 132.6000 812.4000 133.5000 ;
	    RECT 813.3000 133.5000 821.4000 134.4000 ;
	    RECT 813.3000 133.2000 814.5000 133.5000 ;
	    RECT 820.2000 133.2000 821.4000 133.5000 ;
	    RECT 810.9000 131.1000 812.1000 131.4000 ;
	    RECT 815.1000 131.1000 816.3000 131.4000 ;
	    RECT 805.8000 129.3000 807.0000 130.5000 ;
	    RECT 810.9000 130.2000 816.3000 131.1000 ;
	    RECT 812.1000 129.3000 813.0000 130.2000 ;
	    RECT 820.2000 129.3000 821.4000 130.5000 ;
	    RECT 804.9000 123.3000 806.7000 129.3000 ;
	    RECT 809.4000 123.3000 810.6000 129.3000 ;
	    RECT 811.8000 123.3000 813.0000 129.3000 ;
	    RECT 814.2000 123.3000 815.4000 129.3000 ;
	    RECT 818.4000 128.4000 821.4000 129.3000 ;
	    RECT 818.4000 123.3000 819.6000 128.4000 ;
	    RECT 822.6000 123.3000 823.8000 135.0000 ;
	    RECT 825.0000 123.3000 826.2000 135.9000 ;
	    RECT 855.9000 135.3000 856.8000 140.4000 ;
	    RECT 858.7500 138.4500 859.6500 140.4000 ;
	    RECT 1005.0000 139.5000 1018.2000 140.7000 ;
	    RECT 1020.9000 140.1000 1022.1000 143.7000 ;
	    RECT 1026.6000 143.4000 1027.8000 143.7000 ;
	    RECT 1029.0000 143.4000 1030.2001 144.6000 ;
	    RECT 1031.1000 143.4000 1031.4000 144.6000 ;
	    RECT 1035.9000 143.4000 1037.4000 144.6000 ;
	    RECT 1041.0000 143.7000 1044.6000 144.9000 ;
	    RECT 1045.8000 143.7000 1047.0000 149.7000 ;
	    RECT 1024.2001 142.5000 1025.4000 142.8000 ;
	    RECT 1026.6000 142.2000 1027.8000 142.5000 ;
	    RECT 1024.2001 140.4000 1025.4000 141.6000 ;
	    RECT 1026.6000 141.3000 1033.2001 142.2000 ;
	    RECT 1032.0000 141.0000 1033.2001 141.3000 ;
	    RECT 868.2000 138.4500 869.4000 138.6000 ;
	    RECT 858.7500 137.5500 869.4000 138.4500 ;
	    RECT 868.2000 137.4000 869.4000 137.5500 ;
	    RECT 851.4000 123.3000 852.6000 135.3000 ;
	    RECT 855.3000 134.4000 856.8000 135.3000 ;
	    RECT 858.6000 134.4000 859.8000 135.6000 ;
	    RECT 855.3000 123.3000 856.5000 134.4000 ;
	    RECT 857.7000 132.6000 858.6000 133.5000 ;
	    RECT 857.4000 131.4000 858.6000 132.6000 ;
	    RECT 857.7000 123.3000 858.9000 129.3000 ;
	    RECT 870.6000 123.3000 871.8000 139.5000 ;
	    RECT 1005.0000 131.1000 1006.2000 139.5000 ;
	    RECT 1019.1000 138.9000 1022.1000 140.1000 ;
	    RECT 1027.8000 138.9000 1032.6000 140.1000 ;
	    RECT 1036.2001 139.2000 1037.4000 143.4000 ;
	    RECT 1043.4000 142.8000 1044.6000 143.7000 ;
	    RECT 1043.4000 141.9000 1046.1000 142.8000 ;
	    RECT 1044.9000 140.1000 1046.1000 141.9000 ;
	    RECT 1050.6000 141.9000 1051.8000 149.7000 ;
	    RECT 1053.0000 144.0000 1054.2001 149.7000 ;
	    RECT 1055.4000 146.7000 1056.6000 149.7000 ;
	    RECT 1053.0000 142.8000 1054.5000 144.0000 ;
	    RECT 1074.6000 143.7000 1075.8000 149.7000 ;
	    RECT 1078.5000 144.6000 1079.7001 149.7000 ;
	    RECT 1077.0000 143.7000 1079.7001 144.6000 ;
	    RECT 1099.5000 144.6000 1100.7001 149.7000 ;
	    RECT 1099.5000 143.7000 1102.2001 144.6000 ;
	    RECT 1103.4000 143.7000 1104.6000 149.7000 ;
	    RECT 1151.4000 143.7000 1152.6000 149.7000 ;
	    RECT 1153.8000 144.6000 1155.3000 149.7000 ;
	    RECT 1158.0000 144.3000 1160.4000 149.7000 ;
	    RECT 1163.1000 144.6000 1164.6000 149.7000 ;
	    RECT 1050.6000 141.0000 1052.4000 141.9000 ;
	    RECT 1044.9000 138.9000 1050.6000 140.1000 ;
	    RECT 1007.1000 138.0000 1008.3000 138.3000 ;
	    RECT 1007.1000 137.1000 1013.7000 138.0000 ;
	    RECT 1014.6000 137.4000 1015.8000 138.6000 ;
	    RECT 1041.0000 138.0000 1042.2001 138.9000 ;
	    RECT 1051.5000 138.0000 1052.4000 141.0000 ;
	    RECT 1016.7000 137.1000 1042.2001 138.0000 ;
	    RECT 1051.2001 137.1000 1052.4000 138.0000 ;
	    RECT 1049.1000 136.2000 1050.3000 136.5000 ;
	    RECT 1009.8000 134.4000 1011.0000 135.6000 ;
	    RECT 1011.9000 135.3000 1050.3000 136.2000 ;
	    RECT 1014.9000 135.0000 1016.1000 135.3000 ;
	    RECT 1051.2001 134.4000 1052.1000 137.1000 ;
	    RECT 1053.3000 136.2000 1054.5000 142.8000 ;
	    RECT 1074.6000 142.5000 1075.8000 142.8000 ;
	    RECT 1074.6000 140.4000 1075.8000 141.6000 ;
	    RECT 1077.0000 139.5000 1078.2001 143.7000 ;
	    RECT 1101.0000 139.5000 1102.2001 143.7000 ;
	    RECT 1151.4000 142.8000 1155.0000 143.7000 ;
	    RECT 1103.4000 142.5000 1104.6000 142.8000 ;
	    RECT 1153.8000 142.5000 1155.0000 142.8000 ;
	    RECT 1155.9000 142.2000 1157.1000 143.4000 ;
	    RECT 1155.9000 141.6000 1156.8000 142.2000 ;
	    RECT 1103.4000 140.4000 1104.6000 141.6000 ;
	    RECT 1151.4000 140.4000 1152.6000 141.6000 ;
	    RECT 1153.5000 140.4000 1153.8000 141.6000 ;
	    RECT 1155.6000 140.4000 1156.8000 141.6000 ;
	    RECT 1077.0000 138.4500 1078.2001 138.6000 ;
	    RECT 1098.6000 138.4500 1099.8000 138.6000 ;
	    RECT 1077.0000 137.5500 1099.8000 138.4500 ;
	    RECT 1077.0000 137.4000 1078.2001 137.5500 ;
	    RECT 1098.6000 137.4000 1099.8000 137.5500 ;
	    RECT 1101.0000 138.4500 1102.2001 138.6000 ;
	    RECT 1151.5500 138.4500 1152.4501 140.4000 ;
	    RECT 1158.0000 139.5000 1158.9000 144.3000 ;
	    RECT 1165.8000 143.7000 1167.0000 149.7000 ;
	    RECT 1180.2001 146.7000 1181.4000 149.7000 ;
	    RECT 1180.2001 145.5000 1181.4000 145.8000 ;
	    RECT 1159.8000 143.1000 1162.2001 143.4000 ;
	    RECT 1159.8000 142.2000 1162.8000 143.1000 ;
	    RECT 1163.7001 142.8000 1167.0000 143.7000 ;
	    RECT 1180.2001 143.4000 1181.4000 144.6000 ;
	    RECT 1163.7001 142.5000 1164.9000 142.8000 ;
	    RECT 1182.6000 142.5000 1183.8000 149.7000 ;
	    RECT 1213.8000 143.7000 1215.0000 149.7000 ;
	    RECT 1217.7001 143.7000 1220.1000 149.7000 ;
	    RECT 1222.8000 143.7000 1224.0000 149.7000 ;
	    RECT 1254.6000 143.7000 1255.8000 149.7000 ;
	    RECT 1258.5000 143.7000 1260.9000 149.7000 ;
	    RECT 1263.6000 143.7000 1264.8000 149.7000 ;
	    RECT 1278.6000 146.7000 1279.8000 149.7000 ;
	    RECT 1278.6000 145.5000 1279.8000 145.8000 ;
	    RECT 1271.4000 144.4500 1272.6000 144.6000 ;
	    RECT 1278.6000 144.4500 1279.8000 144.6000 ;
	    RECT 1161.9000 141.6000 1162.8000 142.2000 ;
	    RECT 1159.8000 140.1000 1161.0000 141.3000 ;
	    RECT 1161.9000 140.7000 1164.9000 141.6000 ;
	    RECT 1164.6000 140.4000 1164.9000 140.7000 ;
	    RECT 1165.8000 141.4500 1167.0000 141.6000 ;
	    RECT 1168.2001 141.4500 1169.4000 141.6000 ;
	    RECT 1165.8000 140.5500 1169.4000 141.4500 ;
	    RECT 1165.8000 140.4000 1167.0000 140.5500 ;
	    RECT 1168.2001 140.4000 1169.4000 140.5500 ;
	    RECT 1180.2001 141.4500 1181.4000 141.6000 ;
	    RECT 1182.6000 141.4500 1183.8000 141.6000 ;
	    RECT 1180.2001 140.5500 1183.8000 141.4500 ;
	    RECT 1180.2001 140.4000 1181.4000 140.5500 ;
	    RECT 1182.6000 140.4000 1183.8000 140.5500 ;
	    RECT 1211.4000 141.4500 1212.6000 141.6000 ;
	    RECT 1216.2001 141.4500 1217.4000 141.6000 ;
	    RECT 1211.4000 140.5500 1217.4000 141.4500 ;
	    RECT 1211.4000 140.4000 1212.6000 140.5500 ;
	    RECT 1216.2001 140.4000 1217.4000 140.5500 ;
	    RECT 1101.0000 137.5500 1152.4501 138.4500 ;
	    RECT 1101.0000 137.4000 1102.2001 137.5500 ;
	    RECT 1156.2001 137.4000 1157.4000 138.6000 ;
	    RECT 1158.3000 138.3000 1158.9000 139.5000 ;
	    RECT 1160.1000 139.2000 1161.0000 140.1000 ;
	    RECT 1218.6000 139.5000 1219.5000 143.7000 ;
	    RECT 1221.0000 141.4500 1222.2001 141.6000 ;
	    RECT 1242.6000 141.4500 1243.8000 141.6000 ;
	    RECT 1221.0000 140.5500 1243.8000 141.4500 ;
	    RECT 1221.0000 140.4000 1222.2001 140.5500 ;
	    RECT 1242.6000 140.4000 1243.8000 140.5500 ;
	    RECT 1252.2001 141.4500 1253.4000 141.6000 ;
	    RECT 1257.0000 141.4500 1258.2001 141.6000 ;
	    RECT 1252.2001 140.5500 1258.2001 141.4500 ;
	    RECT 1252.2001 140.4000 1253.4000 140.5500 ;
	    RECT 1257.0000 140.4000 1258.2001 140.5500 ;
	    RECT 1259.4000 139.5000 1260.3000 143.7000 ;
	    RECT 1271.4000 143.5500 1279.8000 144.4500 ;
	    RECT 1271.4000 143.4000 1272.6000 143.5500 ;
	    RECT 1278.6000 143.4000 1279.8000 143.5500 ;
	    RECT 1281.0000 142.5000 1282.2001 149.7000 ;
	    RECT 1307.4000 144.0000 1308.6000 149.7000 ;
	    RECT 1309.8000 144.9000 1311.0000 149.7000 ;
	    RECT 1312.2001 144.0000 1313.4000 149.7000 ;
	    RECT 1307.4000 143.7000 1313.4000 144.0000 ;
	    RECT 1314.6000 143.7000 1315.8000 149.7000 ;
	    RECT 1338.6000 144.0000 1339.8000 149.7000 ;
	    RECT 1341.0000 144.9000 1342.2001 149.7000 ;
	    RECT 1343.4000 144.0000 1344.6000 149.7000 ;
	    RECT 1338.6000 143.7000 1344.6000 144.0000 ;
	    RECT 1345.8000 143.7000 1347.0000 149.7000 ;
	    RECT 1379.4000 143.7000 1380.6000 149.7000 ;
	    RECT 1381.8000 144.0000 1383.0000 149.7000 ;
	    RECT 1384.2001 144.9000 1385.4000 149.7000 ;
	    RECT 1386.6000 144.0000 1387.8000 149.7000 ;
	    RECT 1381.8000 143.7000 1387.8000 144.0000 ;
	    RECT 1413.0000 144.0000 1414.2001 149.7000 ;
	    RECT 1415.4000 144.9000 1416.6000 149.7000 ;
	    RECT 1417.8000 144.0000 1419.0000 149.7000 ;
	    RECT 1413.0000 143.7000 1419.0000 144.0000 ;
	    RECT 1420.2001 143.7000 1421.4000 149.7000 ;
	    RECT 1444.2001 146.7000 1445.4000 149.7000 ;
	    RECT 1446.6000 146.7000 1447.8000 149.7000 ;
	    RECT 1444.2001 145.5000 1445.4000 145.8000 ;
	    RECT 1425.0000 144.4500 1426.2001 144.6000 ;
	    RECT 1444.2001 144.4500 1445.4000 144.6000 ;
	    RECT 1307.7001 143.1000 1313.1000 143.7000 ;
	    RECT 1314.6000 142.5000 1315.5000 143.7000 ;
	    RECT 1338.9000 143.1000 1344.3000 143.7000 ;
	    RECT 1345.8000 142.5000 1346.7001 143.7000 ;
	    RECT 1379.7001 142.5000 1380.6000 143.7000 ;
	    RECT 1382.1000 143.1000 1387.5000 143.7000 ;
	    RECT 1413.3000 143.1000 1418.7001 143.7000 ;
	    RECT 1420.2001 142.5000 1421.1000 143.7000 ;
	    RECT 1425.0000 143.5500 1445.4000 144.4500 ;
	    RECT 1425.0000 143.4000 1426.2001 143.5500 ;
	    RECT 1444.2001 143.4000 1445.4000 143.5500 ;
	    RECT 1446.9000 143.4000 1447.8000 146.7000 ;
	    RECT 1449.0000 144.3000 1450.2001 149.7000 ;
	    RECT 1451.4000 143.7000 1452.6000 149.7000 ;
	    RECT 1446.9000 142.5000 1450.5000 143.4000 ;
	    RECT 1261.8000 141.4500 1263.0000 141.6000 ;
	    RECT 1276.2001 141.4500 1277.4000 141.6000 ;
	    RECT 1278.6000 141.4500 1279.8000 141.6000 ;
	    RECT 1261.8000 140.5500 1279.8000 141.4500 ;
	    RECT 1261.8000 140.4000 1263.0000 140.5500 ;
	    RECT 1276.2001 140.4000 1277.4000 140.5500 ;
	    RECT 1278.6000 140.4000 1279.8000 140.5500 ;
	    RECT 1281.0000 141.4500 1282.2001 141.6000 ;
	    RECT 1305.0000 141.4500 1306.2001 141.6000 ;
	    RECT 1281.0000 140.5500 1306.2001 141.4500 ;
	    RECT 1281.0000 140.4000 1282.2001 140.5500 ;
	    RECT 1305.0000 140.4000 1306.2001 140.5500 ;
	    RECT 1307.4000 140.4000 1308.6000 141.6000 ;
	    RECT 1309.5000 140.7000 1309.8000 142.2000 ;
	    RECT 1311.9000 140.4000 1313.7001 141.6000 ;
	    RECT 1314.6000 141.4500 1315.8000 141.6000 ;
	    RECT 1336.2001 141.4500 1337.4000 141.6000 ;
	    RECT 1314.6000 140.5500 1337.4000 141.4500 ;
	    RECT 1314.6000 140.4000 1315.8000 140.5500 ;
	    RECT 1336.2001 140.4000 1337.4000 140.5500 ;
	    RECT 1338.6000 140.4000 1339.8000 141.6000 ;
	    RECT 1340.7001 140.7000 1341.0000 142.2000 ;
	    RECT 1343.1000 140.4000 1344.9000 141.6000 ;
	    RECT 1345.8000 141.4500 1347.0000 141.6000 ;
	    RECT 1348.2001 141.4500 1349.4000 141.6000 ;
	    RECT 1345.8000 140.5500 1349.4000 141.4500 ;
	    RECT 1345.8000 140.4000 1347.0000 140.5500 ;
	    RECT 1348.2001 140.4000 1349.4000 140.5500 ;
	    RECT 1379.4000 140.4000 1380.6000 141.6000 ;
	    RECT 1381.5000 140.4000 1383.3000 141.6000 ;
	    RECT 1385.4000 140.7000 1385.7001 142.2000 ;
	    RECT 1386.6000 141.4500 1387.8000 141.6000 ;
	    RECT 1413.0000 141.4500 1414.2001 141.6000 ;
	    RECT 1386.6000 140.5500 1414.2001 141.4500 ;
	    RECT 1415.1000 140.7000 1415.4000 142.2000 ;
	    RECT 1386.6000 140.4000 1387.8000 140.5500 ;
	    RECT 1413.0000 140.4000 1414.2001 140.5500 ;
	    RECT 1417.5000 140.4000 1419.3000 141.6000 ;
	    RECT 1420.2001 141.4500 1421.4000 141.6000 ;
	    RECT 1441.8000 141.4500 1443.0000 141.6000 ;
	    RECT 1420.2001 140.5500 1443.0000 141.4500 ;
	    RECT 1420.2001 140.4000 1421.4000 140.5500 ;
	    RECT 1441.8000 140.4000 1443.0000 140.5500 ;
	    RECT 1446.6000 140.4000 1447.8000 141.6000 ;
	    RECT 1309.8000 139.5000 1311.0000 139.8000 ;
	    RECT 1160.1000 138.3000 1164.0000 139.2000 ;
	    RECT 1162.8000 138.0000 1164.0000 138.3000 ;
	    RECT 1159.5000 137.1000 1160.7001 137.4000 ;
	    RECT 1019.4000 134.1000 1020.6000 134.4000 ;
	    RECT 1012.5000 133.5000 1020.6000 134.1000 ;
	    RECT 1011.3000 133.2000 1020.6000 133.5000 ;
	    RECT 1022.1000 133.5000 1035.0000 134.4000 ;
	    RECT 1007.4000 132.0000 1009.8000 133.2000 ;
	    RECT 1011.3000 132.3000 1013.4000 133.2000 ;
	    RECT 1022.1000 132.3000 1023.0000 133.5000 ;
	    RECT 1033.8000 133.2000 1035.0000 133.5000 ;
	    RECT 1038.6000 133.5000 1052.1000 134.4000 ;
	    RECT 1053.0000 135.0000 1054.5000 136.2000 ;
	    RECT 1053.0000 133.5000 1054.2001 135.0000 ;
	    RECT 1038.6000 133.2000 1039.8000 133.5000 ;
	    RECT 1008.9000 131.4000 1009.8000 132.0000 ;
	    RECT 1014.3000 131.4000 1023.0000 132.3000 ;
	    RECT 1023.9000 131.4000 1027.8000 132.6000 ;
	    RECT 1005.0000 130.2000 1008.0000 131.1000 ;
	    RECT 1008.9000 130.2000 1015.2000 131.4000 ;
	    RECT 1007.1000 129.3000 1008.0000 130.2000 ;
	    RECT 873.0000 123.3000 874.2000 129.3000 ;
	    RECT 1005.0000 123.3000 1006.2000 129.3000 ;
	    RECT 1007.1000 128.4000 1008.6000 129.3000 ;
	    RECT 1007.4000 123.3000 1008.6000 128.4000 ;
	    RECT 1009.8000 122.4000 1011.0000 129.3000 ;
	    RECT 1012.2000 123.3000 1013.4000 130.2000 ;
	    RECT 1014.6000 123.3000 1015.8000 129.3000 ;
	    RECT 1017.0000 123.3000 1018.2000 127.5000 ;
	    RECT 1019.4000 123.3000 1020.6000 127.5000 ;
	    RECT 1021.8000 123.3000 1023.0000 130.5000 ;
	    RECT 1024.2001 123.3000 1025.4000 129.3000 ;
	    RECT 1026.6000 123.3000 1027.8000 130.5000 ;
	    RECT 1029.0000 123.3000 1030.2001 129.3000 ;
	    RECT 1031.4000 123.3000 1032.6000 132.6000 ;
	    RECT 1043.4000 131.4000 1047.3000 132.6000 ;
	    RECT 1036.2001 130.2000 1042.5000 131.4000 ;
	    RECT 1033.8000 123.3000 1035.0000 127.5000 ;
	    RECT 1036.2001 123.3000 1037.4000 127.5000 ;
	    RECT 1038.6000 123.3000 1039.8000 127.5000 ;
	    RECT 1041.0000 123.3000 1042.2001 129.3000 ;
	    RECT 1043.4000 123.3000 1044.6000 131.4000 ;
	    RECT 1051.2001 131.1000 1052.1000 133.5000 ;
	    RECT 1053.0000 131.4000 1054.2001 132.6000 ;
	    RECT 1048.2001 130.2000 1052.1000 131.1000 ;
	    RECT 1045.8000 123.3000 1047.0000 129.3000 ;
	    RECT 1048.2001 123.3000 1049.4000 130.2000 ;
	    RECT 1050.6000 123.3000 1051.8000 129.3000 ;
	    RECT 1053.0000 123.3000 1054.2001 130.5000 ;
	    RECT 1055.4000 123.3000 1056.6000 129.3000 ;
	    RECT 1074.6000 123.3000 1075.8000 129.3000 ;
	    RECT 1077.0000 123.3000 1078.2001 136.5000 ;
	    RECT 1079.4000 134.4000 1080.6000 135.6000 ;
	    RECT 1081.8000 135.4500 1083.0000 135.6000 ;
	    RECT 1098.6000 135.4500 1099.8000 135.6000 ;
	    RECT 1081.8000 134.5500 1099.8000 135.4500 ;
	    RECT 1081.8000 134.4000 1083.0000 134.5500 ;
	    RECT 1098.6000 134.4000 1099.8000 134.5500 ;
	    RECT 1079.4000 133.2000 1080.6000 133.5000 ;
	    RECT 1098.6000 133.2000 1099.8000 133.5000 ;
	    RECT 1079.4000 123.3000 1080.6000 129.3000 ;
	    RECT 1098.6000 123.3000 1099.8000 129.3000 ;
	    RECT 1101.0000 123.3000 1102.2001 136.5000 ;
	    RECT 1157.4000 135.3000 1158.3000 136.5000 ;
	    RECT 1159.5000 136.2000 1164.6000 137.1000 ;
	    RECT 1163.7001 135.3000 1164.6000 136.2000 ;
	    RECT 1151.4000 134.4000 1155.0000 135.3000 ;
	    RECT 1157.4000 134.4000 1160.4000 135.3000 ;
	    RECT 1103.4000 123.3000 1104.6000 129.3000 ;
	    RECT 1151.4000 123.3000 1152.6000 134.4000 ;
	    RECT 1153.8000 134.1000 1155.0000 134.4000 ;
	    RECT 1153.8000 123.3000 1155.3000 133.2000 ;
	    RECT 1158.0000 123.3000 1160.4000 134.4000 ;
	    RECT 1163.7001 134.4000 1167.0000 135.3000 ;
	    RECT 1163.7001 134.1000 1164.9000 134.4000 ;
	    RECT 1163.1000 123.3000 1164.6000 133.2000 ;
	    RECT 1165.8000 123.3000 1167.0000 134.4000 ;
	    RECT 1180.2001 123.3000 1181.4000 129.3000 ;
	    RECT 1182.6000 123.3000 1183.8000 139.5000 ;
	    RECT 1216.5000 138.6000 1217.7001 139.5000 ;
	    RECT 1221.0000 139.2000 1222.2001 139.5000 ;
	    RECT 1257.3000 138.6000 1258.5000 139.5000 ;
	    RECT 1261.8000 139.2000 1263.0000 139.5000 ;
	    RECT 1187.4000 138.4500 1188.6000 138.6000 ;
	    RECT 1213.8000 138.4500 1215.0000 138.6000 ;
	    RECT 1187.4000 137.5500 1215.0000 138.4500 ;
	    RECT 1187.4000 137.4000 1188.6000 137.5500 ;
	    RECT 1213.8000 137.4000 1215.0000 137.5500 ;
	    RECT 1218.6000 137.4000 1219.8000 138.6000 ;
	    RECT 1216.5000 136.5000 1217.7001 137.1000 ;
	    RECT 1222.2001 136.8000 1222.5000 138.3000 ;
	    RECT 1223.4000 137.4000 1224.6000 138.6000 ;
	    RECT 1254.6000 137.4000 1255.8000 138.6000 ;
	    RECT 1259.4000 137.4000 1260.6000 138.6000 ;
	    RECT 1264.2001 138.4500 1265.4000 138.6000 ;
	    RECT 1278.6000 138.4500 1279.8000 138.6000 ;
	    RECT 1257.3000 136.5000 1258.5000 137.1000 ;
	    RECT 1263.0000 136.8000 1263.3000 138.3000 ;
	    RECT 1264.2001 137.5500 1279.8000 138.4500 ;
	    RECT 1264.2001 137.4000 1265.4000 137.5500 ;
	    RECT 1278.6000 137.4000 1279.8000 137.5500 ;
	    RECT 1213.8000 136.2000 1215.0000 136.5000 ;
	    RECT 1216.5000 136.2000 1219.5000 136.5000 ;
	    RECT 1254.6000 136.2000 1255.8000 136.5000 ;
	    RECT 1257.3000 136.2000 1260.3000 136.5000 ;
	    RECT 1216.5000 135.3000 1217.4000 136.2000 ;
	    RECT 1257.3000 135.3000 1258.2001 136.2000 ;
	    RECT 1213.8000 124.2000 1215.0000 135.3000 ;
	    RECT 1216.2001 125.1000 1217.4000 135.3000 ;
	    RECT 1218.6000 134.4000 1224.6000 135.3000 ;
	    RECT 1218.6000 124.2000 1219.8000 134.4000 ;
	    RECT 1213.8000 123.3000 1219.8000 124.2000 ;
	    RECT 1221.0000 123.3000 1222.2001 133.5000 ;
	    RECT 1223.4000 123.3000 1224.6000 134.4000 ;
	    RECT 1254.6000 124.2000 1255.8000 135.3000 ;
	    RECT 1257.0000 125.1000 1258.2001 135.3000 ;
	    RECT 1259.4000 134.4000 1265.4000 135.3000 ;
	    RECT 1259.4000 124.2000 1260.6000 134.4000 ;
	    RECT 1254.6000 123.3000 1260.6000 124.2000 ;
	    RECT 1261.8000 123.3000 1263.0000 133.5000 ;
	    RECT 1264.2001 123.3000 1265.4000 134.4000 ;
	    RECT 1278.6000 123.3000 1279.8000 129.3000 ;
	    RECT 1281.0000 123.3000 1282.2001 139.5000 ;
	    RECT 1309.8000 137.4000 1311.0000 138.6000 ;
	    RECT 1311.9000 135.3000 1312.8000 140.4000 ;
	    RECT 1341.0000 139.5000 1342.2001 139.8000 ;
	    RECT 1336.2001 138.4500 1337.4000 138.6000 ;
	    RECT 1341.0000 138.4500 1342.2001 138.6000 ;
	    RECT 1336.2001 137.5500 1342.2001 138.4500 ;
	    RECT 1336.2001 137.4000 1337.4000 137.5500 ;
	    RECT 1341.0000 137.4000 1342.2001 137.5500 ;
	    RECT 1307.4000 123.3000 1308.6000 135.3000 ;
	    RECT 1311.3000 134.4000 1312.8000 135.3000 ;
	    RECT 1314.6000 135.4500 1315.8000 135.6000 ;
	    RECT 1331.4000 135.4500 1332.6000 135.6000 ;
	    RECT 1314.6000 134.5500 1332.6000 135.4500 ;
	    RECT 1343.1000 135.3000 1344.0000 140.4000 ;
	    RECT 1314.6000 134.4000 1315.8000 134.5500 ;
	    RECT 1331.4000 134.4000 1332.6000 134.5500 ;
	    RECT 1311.3000 123.3000 1312.5000 134.4000 ;
	    RECT 1313.7001 132.6000 1314.6000 133.5000 ;
	    RECT 1313.4000 131.4000 1314.6000 132.6000 ;
	    RECT 1313.7001 123.3000 1314.9000 129.3000 ;
	    RECT 1338.6000 123.3000 1339.8000 135.3000 ;
	    RECT 1342.5000 134.4000 1344.0000 135.3000 ;
	    RECT 1345.8000 134.4000 1347.0000 135.6000 ;
	    RECT 1377.0000 135.4500 1378.2001 135.6000 ;
	    RECT 1379.4000 135.4500 1380.6000 135.6000 ;
	    RECT 1377.0000 134.5500 1380.6000 135.4500 ;
	    RECT 1377.0000 134.4000 1378.2001 134.5500 ;
	    RECT 1379.4000 134.4000 1380.6000 134.5500 ;
	    RECT 1382.4000 135.3000 1383.3000 140.4000 ;
	    RECT 1384.2001 139.5000 1385.4000 139.8000 ;
	    RECT 1415.4000 139.5000 1416.6000 139.8000 ;
	    RECT 1384.2001 138.4500 1385.4000 138.6000 ;
	    RECT 1415.4000 138.4500 1416.6000 138.6000 ;
	    RECT 1384.2001 137.5500 1416.6000 138.4500 ;
	    RECT 1384.2001 137.4000 1385.4000 137.5500 ;
	    RECT 1415.4000 137.4000 1416.6000 137.5500 ;
	    RECT 1417.5000 135.3000 1418.4000 140.4000 ;
	    RECT 1447.2001 139.2000 1448.4000 139.5000 ;
	    RECT 1449.6000 138.0000 1450.5000 142.5000 ;
	    RECT 1451.7001 139.5000 1452.6000 143.7000 ;
	    RECT 1475.4000 140.7000 1476.6000 149.7000 ;
	    RECT 1480.8000 141.3000 1482.0000 149.7000 ;
	    RECT 1509.0000 143.7000 1510.2001 149.7000 ;
	    RECT 1511.4000 144.0000 1512.6000 149.7000 ;
	    RECT 1513.8000 144.9000 1515.0000 149.7000 ;
	    RECT 1516.2001 144.0000 1517.4000 149.7000 ;
	    RECT 1511.4000 143.7000 1517.4000 144.0000 ;
	    RECT 1540.2001 144.0000 1541.4000 149.7000 ;
	    RECT 1542.6000 144.9000 1543.8000 149.7000 ;
	    RECT 1545.0000 144.0000 1546.2001 149.7000 ;
	    RECT 1540.2001 143.7000 1546.2001 144.0000 ;
	    RECT 1547.4000 143.7000 1548.6000 149.7000 ;
	    RECT 1509.3000 142.5000 1510.2001 143.7000 ;
	    RECT 1511.7001 143.1000 1517.1000 143.7000 ;
	    RECT 1540.5000 143.1000 1545.9000 143.7000 ;
	    RECT 1547.4000 142.5000 1548.3000 143.7000 ;
	    RECT 1480.8000 140.7000 1483.5000 141.3000 ;
	    RECT 1481.1000 140.4000 1483.5000 140.7000 ;
	    RECT 1509.0000 140.4000 1510.2001 141.6000 ;
	    RECT 1511.1000 140.4000 1512.9000 141.6000 ;
	    RECT 1515.0000 140.7000 1515.3000 142.2000 ;
	    RECT 1516.2001 141.4500 1517.4000 141.6000 ;
	    RECT 1540.2001 141.4500 1541.4000 141.6000 ;
	    RECT 1516.2001 140.5500 1541.4000 141.4500 ;
	    RECT 1542.3000 140.7000 1542.6000 142.2000 ;
	    RECT 1516.2001 140.4000 1517.4000 140.5500 ;
	    RECT 1540.2001 140.4000 1541.4000 140.5500 ;
	    RECT 1544.7001 140.4000 1546.5000 141.6000 ;
	    RECT 1547.4000 141.4500 1548.6000 141.6000 ;
	    RECT 1554.6000 141.4500 1555.8000 141.6000 ;
	    RECT 1547.4000 140.5500 1555.8000 141.4500 ;
	    RECT 1547.4000 140.4000 1548.6000 140.5500 ;
	    RECT 1554.6000 140.4000 1555.8000 140.5500 ;
	    RECT 1449.3000 137.1000 1450.5000 138.0000 ;
	    RECT 1451.4000 138.4500 1452.6000 138.6000 ;
	    RECT 1473.0000 138.4500 1474.2001 138.6000 ;
	    RECT 1451.4000 137.5500 1474.2001 138.4500 ;
	    RECT 1451.4000 137.4000 1452.6000 137.5500 ;
	    RECT 1473.0000 137.4000 1474.2001 137.5500 ;
	    RECT 1477.8000 137.4000 1479.0000 138.6000 ;
	    RECT 1479.9000 137.4000 1480.2001 138.6000 ;
	    RECT 1444.2001 136.8000 1450.5000 137.1000 ;
	    RECT 1444.2001 136.2000 1450.2001 136.8000 ;
	    RECT 1475.4000 136.5000 1476.6000 136.8000 ;
	    RECT 1482.6000 136.5000 1483.5000 140.4000 ;
	    RECT 1382.4000 134.4000 1383.9000 135.3000 ;
	    RECT 1342.5000 123.3000 1343.7001 134.4000 ;
	    RECT 1344.9000 132.6000 1345.8000 133.5000 ;
	    RECT 1344.6000 131.4000 1345.8000 132.6000 ;
	    RECT 1380.6000 132.6000 1381.5000 133.5000 ;
	    RECT 1380.6000 131.4000 1381.8000 132.6000 ;
	    RECT 1344.9000 123.3000 1346.1000 129.3000 ;
	    RECT 1380.3000 123.3000 1381.5000 129.3000 ;
	    RECT 1382.7001 123.3000 1383.9000 134.4000 ;
	    RECT 1386.6000 123.3000 1387.8000 135.3000 ;
	    RECT 1413.0000 123.3000 1414.2001 135.3000 ;
	    RECT 1416.9000 134.4000 1418.4000 135.3000 ;
	    RECT 1420.2001 134.4000 1421.4000 135.6000 ;
	    RECT 1416.9000 123.3000 1418.1000 134.4000 ;
	    RECT 1419.3000 132.6000 1420.2001 133.5000 ;
	    RECT 1419.0000 131.4000 1420.2001 132.6000 ;
	    RECT 1419.3000 123.3000 1420.5000 129.3000 ;
	    RECT 1444.2001 123.3000 1445.4000 136.2000 ;
	    RECT 1451.7001 135.3000 1452.6000 136.5000 ;
	    RECT 1448.1000 123.3000 1449.3000 135.3000 ;
	    RECT 1450.5000 134.4000 1452.6000 135.3000 ;
	    RECT 1475.4000 135.4500 1476.6000 135.6000 ;
	    RECT 1477.8000 135.4500 1479.0000 135.6000 ;
	    RECT 1475.4000 134.5500 1479.0000 135.4500 ;
	    RECT 1475.4000 134.4000 1476.6000 134.5500 ;
	    RECT 1477.8000 134.4000 1479.0000 134.5500 ;
	    RECT 1482.6000 135.4500 1483.8000 135.6000 ;
	    RECT 1485.0000 135.4500 1486.2001 135.6000 ;
	    RECT 1482.6000 134.5500 1486.2001 135.4500 ;
	    RECT 1482.6000 134.4000 1483.8000 134.5500 ;
	    RECT 1485.0000 134.4000 1486.2001 134.5500 ;
	    RECT 1494.6000 135.4500 1495.8000 135.6000 ;
	    RECT 1509.0000 135.4500 1510.2001 135.6000 ;
	    RECT 1494.6000 134.5500 1510.2001 135.4500 ;
	    RECT 1494.6000 134.4000 1495.8000 134.5500 ;
	    RECT 1509.0000 134.4000 1510.2001 134.5500 ;
	    RECT 1512.0000 135.3000 1512.9000 140.4000 ;
	    RECT 1513.8000 139.5000 1515.0000 139.8000 ;
	    RECT 1542.6000 139.5000 1543.8000 139.8000 ;
	    RECT 1513.8000 138.4500 1515.0000 138.6000 ;
	    RECT 1516.2001 138.4500 1517.4000 138.6000 ;
	    RECT 1542.6000 138.4500 1543.8000 138.6000 ;
	    RECT 1513.8000 137.5500 1543.8000 138.4500 ;
	    RECT 1513.8000 137.4000 1515.0000 137.5500 ;
	    RECT 1516.2001 137.4000 1517.4000 137.5500 ;
	    RECT 1542.6000 137.4000 1543.8000 137.5500 ;
	    RECT 1544.7001 135.3000 1545.6000 140.4000 ;
	    RECT 1512.0000 134.4000 1513.5000 135.3000 ;
	    RECT 1450.5000 123.3000 1451.7001 134.4000 ;
	    RECT 1480.2001 133.5000 1481.4000 133.8000 ;
	    RECT 1473.0000 132.4500 1474.2001 132.6000 ;
	    RECT 1480.2001 132.4500 1481.4000 132.6000 ;
	    RECT 1473.0000 131.5500 1481.4000 132.4500 ;
	    RECT 1473.0000 131.4000 1474.2001 131.5500 ;
	    RECT 1480.2001 131.4000 1481.4000 131.5500 ;
	    RECT 1482.6000 130.5000 1483.5000 133.5000 ;
	    RECT 1510.2001 132.6000 1511.1000 133.5000 ;
	    RECT 1510.2001 131.4000 1511.4000 132.6000 ;
	    RECT 1478.1000 129.6000 1483.5000 130.5000 ;
	    RECT 1478.1000 129.3000 1479.0000 129.6000 ;
	    RECT 1475.4000 123.3000 1476.6000 129.3000 ;
	    RECT 1477.8000 123.3000 1479.0000 129.3000 ;
	    RECT 1482.6000 129.3000 1483.5000 129.6000 ;
	    RECT 1480.2001 123.3000 1481.4000 128.7000 ;
	    RECT 1482.6000 123.3000 1483.8000 129.3000 ;
	    RECT 1509.9000 123.3000 1511.1000 129.3000 ;
	    RECT 1512.3000 123.3000 1513.5000 134.4000 ;
	    RECT 1516.2001 123.3000 1517.4000 135.3000 ;
	    RECT 1540.2001 123.3000 1541.4000 135.3000 ;
	    RECT 1544.1000 134.4000 1545.6000 135.3000 ;
	    RECT 1547.4000 135.4500 1548.6000 135.6000 ;
	    RECT 1557.0000 135.4500 1558.2001 135.6000 ;
	    RECT 1547.4000 134.5500 1558.2001 135.4500 ;
	    RECT 1547.4000 134.4000 1548.6000 134.5500 ;
	    RECT 1557.0000 134.4000 1558.2001 134.5500 ;
	    RECT 1544.1000 123.3000 1545.3000 134.4000 ;
	    RECT 1546.5000 132.6000 1547.4000 133.5000 ;
	    RECT 1546.2001 131.4000 1547.4000 132.6000 ;
	    RECT 1546.5000 123.3000 1547.7001 129.3000 ;
	    RECT 1.2000 120.6000 1569.0000 122.4000 ;
	    RECT 18.6000 113.7000 19.8000 119.7000 ;
	    RECT 18.6000 109.5000 19.8000 109.8000 ;
	    RECT 18.6000 107.4000 19.8000 108.6000 ;
	    RECT 21.0000 106.5000 22.2000 119.7000 ;
	    RECT 23.4000 113.7000 24.6000 119.7000 ;
	    RECT 48.3000 113.7000 49.5000 119.7000 ;
	    RECT 48.6000 110.4000 49.8000 111.6000 ;
	    RECT 48.6000 109.5000 49.5000 110.4000 ;
	    RECT 50.7000 108.6000 51.9000 119.7000 ;
	    RECT 47.4000 107.4000 48.6000 108.6000 ;
	    RECT 50.4000 107.7000 51.9000 108.6000 ;
	    RECT 54.6000 107.7000 55.8000 119.7000 ;
	    RECT 21.0000 105.4500 22.2000 105.6000 ;
	    RECT 47.5500 105.4500 48.4500 107.4000 ;
	    RECT 21.0000 104.5500 48.4500 105.4500 ;
	    RECT 21.0000 104.4000 22.2000 104.5500 ;
	    RECT 21.0000 99.3000 22.2000 103.5000 ;
	    RECT 50.4000 102.6000 51.3000 107.7000 ;
	    RECT 52.2000 105.4500 53.4000 105.6000 ;
	    RECT 52.2000 104.5500 58.0500 105.4500 ;
	    RECT 52.2000 104.4000 53.4000 104.5500 ;
	    RECT 52.2000 103.2000 53.4000 103.5000 ;
	    RECT 23.4000 101.4000 24.6000 102.6000 ;
	    RECT 47.4000 101.4000 48.6000 102.6000 ;
	    RECT 49.5000 101.4000 51.3000 102.6000 ;
	    RECT 53.4000 100.8000 53.7000 102.3000 ;
	    RECT 54.6000 101.4000 55.8000 102.6000 ;
	    RECT 57.1500 102.4500 58.0500 104.5500 ;
	    RECT 69.0000 103.5000 70.2000 119.7000 ;
	    RECT 71.4000 113.7000 72.6000 119.7000 ;
	    RECT 203.4000 113.7000 204.6000 119.7000 ;
	    RECT 205.8000 112.5000 207.0000 119.7000 ;
	    RECT 208.2000 113.7000 209.4000 119.7000 ;
	    RECT 210.6000 112.8000 211.8000 119.7000 ;
	    RECT 213.0000 113.7000 214.2000 119.7000 ;
	    RECT 207.9000 111.9000 211.8000 112.8000 ;
	    RECT 179.4000 111.4500 180.6000 111.6000 ;
	    RECT 205.8000 111.4500 207.0000 111.6000 ;
	    RECT 179.4000 110.5500 207.0000 111.4500 ;
	    RECT 179.4000 110.4000 180.6000 110.5500 ;
	    RECT 205.8000 110.4000 207.0000 110.5500 ;
	    RECT 207.9000 109.5000 208.8000 111.9000 ;
	    RECT 215.4000 111.6000 216.6000 119.7000 ;
	    RECT 217.8000 113.7000 219.0000 119.7000 ;
	    RECT 220.2000 115.5000 221.4000 119.7000 ;
	    RECT 222.6000 115.5000 223.8000 119.7000 ;
	    RECT 225.0000 115.5000 226.2000 119.7000 ;
	    RECT 217.5000 111.6000 223.8000 112.8000 ;
	    RECT 212.7000 110.4000 216.6000 111.6000 ;
	    RECT 227.4000 110.4000 228.6000 119.7000 ;
	    RECT 229.8000 113.7000 231.0000 119.7000 ;
	    RECT 232.2000 112.5000 233.4000 119.7000 ;
	    RECT 234.6000 113.7000 235.8000 119.7000 ;
	    RECT 237.0000 112.5000 238.2000 119.7000 ;
	    RECT 239.4000 115.5000 240.6000 119.7000 ;
	    RECT 241.8000 115.5000 243.0000 119.7000 ;
	    RECT 244.2000 113.7000 245.4000 119.7000 ;
	    RECT 246.6000 112.8000 247.8000 119.7000 ;
	    RECT 249.0000 113.7000 250.2000 120.6000 ;
	    RECT 251.4000 114.6000 252.6000 119.7000 ;
	    RECT 251.4000 113.7000 252.9000 114.6000 ;
	    RECT 253.8000 113.7000 255.0000 119.7000 ;
	    RECT 252.0000 112.8000 252.9000 113.7000 ;
	    RECT 244.8000 111.6000 251.1000 112.8000 ;
	    RECT 252.0000 111.9000 255.0000 112.8000 ;
	    RECT 232.2000 110.4000 236.1000 111.6000 ;
	    RECT 237.0000 110.7000 245.7000 111.6000 ;
	    RECT 250.2000 111.0000 251.1000 111.6000 ;
	    RECT 220.2000 109.5000 221.4000 109.8000 ;
	    RECT 205.8000 108.0000 207.0000 109.5000 ;
	    RECT 205.5000 106.8000 207.0000 108.0000 ;
	    RECT 207.9000 108.6000 221.4000 109.5000 ;
	    RECT 225.0000 109.5000 226.2000 109.8000 ;
	    RECT 237.0000 109.5000 237.9000 110.7000 ;
	    RECT 246.6000 109.8000 248.7000 110.7000 ;
	    RECT 250.2000 109.8000 252.6000 111.0000 ;
	    RECT 225.0000 108.6000 237.9000 109.5000 ;
	    RECT 239.4000 109.5000 248.7000 109.8000 ;
	    RECT 239.4000 108.9000 247.5000 109.5000 ;
	    RECT 239.4000 108.6000 240.6000 108.9000 ;
	    RECT 69.0000 102.4500 70.2000 102.6000 ;
	    RECT 57.1500 101.5500 70.2000 102.4500 ;
	    RECT 69.0000 101.4000 70.2000 101.5500 ;
	    RECT 23.4000 100.2000 24.6000 100.5000 ;
	    RECT 47.7000 99.3000 48.6000 100.5000 ;
	    RECT 50.1000 99.3000 55.5000 99.9000 ;
	    RECT 19.5000 98.4000 22.2000 99.3000 ;
	    RECT 19.5000 93.3000 20.7000 98.4000 ;
	    RECT 23.4000 93.3000 24.6000 99.3000 ;
	    RECT 47.4000 93.3000 48.6000 99.3000 ;
	    RECT 49.8000 99.0000 55.8000 99.3000 ;
	    RECT 49.8000 93.3000 51.0000 99.0000 ;
	    RECT 52.2000 93.3000 53.4000 98.1000 ;
	    RECT 54.6000 93.3000 55.8000 99.0000 ;
	    RECT 69.0000 93.3000 70.2000 100.5000 ;
	    RECT 205.5000 100.2000 206.7000 106.8000 ;
	    RECT 207.9000 105.9000 208.8000 108.6000 ;
	    RECT 243.9000 107.7000 245.1000 108.0000 ;
	    RECT 209.7000 106.8000 248.1000 107.7000 ;
	    RECT 249.0000 107.4000 250.2000 108.6000 ;
	    RECT 209.7000 106.5000 210.9000 106.8000 ;
	    RECT 207.6000 105.0000 208.8000 105.9000 ;
	    RECT 217.8000 105.0000 243.3000 105.9000 ;
	    RECT 207.6000 102.0000 208.5000 105.0000 ;
	    RECT 217.8000 104.1000 219.0000 105.0000 ;
	    RECT 244.2000 104.4000 245.4000 105.6000 ;
	    RECT 246.3000 105.0000 252.9000 105.9000 ;
	    RECT 251.7000 104.7000 252.9000 105.0000 ;
	    RECT 209.4000 102.9000 215.1000 104.1000 ;
	    RECT 207.6000 101.1000 209.4000 102.0000 ;
	    RECT 71.4000 99.4500 72.6000 99.6000 ;
	    RECT 172.2000 99.4500 173.4000 99.6000 ;
	    RECT 71.4000 98.5500 173.4000 99.4500 ;
	    RECT 205.5000 99.0000 207.0000 100.2000 ;
	    RECT 71.4000 98.4000 72.6000 98.5500 ;
	    RECT 172.2000 98.4000 173.4000 98.5500 ;
	    RECT 71.4000 97.2000 72.6000 97.5000 ;
	    RECT 71.4000 93.3000 72.6000 96.3000 ;
	    RECT 203.4000 93.3000 204.6000 96.3000 ;
	    RECT 205.8000 93.3000 207.0000 99.0000 ;
	    RECT 208.2000 93.3000 209.4000 101.1000 ;
	    RECT 213.9000 101.1000 215.1000 102.9000 ;
	    RECT 213.9000 100.2000 216.6000 101.1000 ;
	    RECT 215.4000 99.3000 216.6000 100.2000 ;
	    RECT 222.6000 99.6000 223.8000 103.8000 ;
	    RECT 227.4000 102.9000 232.2000 104.1000 ;
	    RECT 237.9000 102.9000 240.9000 104.1000 ;
	    RECT 253.8000 103.5000 255.0000 111.9000 ;
	    RECT 277.8000 107.7000 279.0000 119.7000 ;
	    RECT 281.7000 108.6000 282.9000 119.7000 ;
	    RECT 284.1000 113.7000 285.3000 119.7000 ;
	    RECT 312.3000 113.7000 313.5000 119.7000 ;
	    RECT 283.8000 110.4000 285.0000 111.6000 ;
	    RECT 284.1000 109.5000 285.0000 110.4000 ;
	    RECT 312.6000 110.4000 313.8000 111.6000 ;
	    RECT 312.6000 109.5000 313.5000 110.4000 ;
	    RECT 314.7000 108.6000 315.9000 119.7000 ;
	    RECT 281.7000 107.7000 283.2000 108.6000 ;
	    RECT 280.2000 104.4000 281.4000 105.6000 ;
	    RECT 226.8000 101.7000 228.0000 102.0000 ;
	    RECT 226.8000 100.8000 233.4000 101.7000 ;
	    RECT 234.6000 101.4000 235.8000 102.6000 ;
	    RECT 232.2000 100.5000 233.4000 100.8000 ;
	    RECT 234.6000 100.2000 235.8000 100.5000 ;
	    RECT 213.0000 93.3000 214.2000 99.3000 ;
	    RECT 215.4000 98.1000 219.0000 99.3000 ;
	    RECT 222.6000 98.4000 224.1000 99.6000 ;
	    RECT 228.6000 98.4000 228.9000 99.6000 ;
	    RECT 229.8000 98.4000 231.0000 99.6000 ;
	    RECT 232.2000 99.3000 233.4000 99.6000 ;
	    RECT 237.9000 99.3000 239.1000 102.9000 ;
	    RECT 241.8000 102.3000 255.0000 103.5000 ;
	    RECT 280.2000 103.2000 281.4000 103.5000 ;
	    RECT 282.3000 102.6000 283.2000 107.7000 ;
	    RECT 285.0000 107.4000 286.2000 108.6000 ;
	    RECT 292.2000 108.4500 293.4000 108.6000 ;
	    RECT 311.4000 108.4500 312.6000 108.6000 ;
	    RECT 292.2000 107.5500 312.6000 108.4500 ;
	    RECT 292.2000 107.4000 293.4000 107.5500 ;
	    RECT 311.4000 107.4000 312.6000 107.5500 ;
	    RECT 314.4000 107.7000 315.9000 108.6000 ;
	    RECT 318.6000 107.7000 319.8000 119.7000 ;
	    RECT 330.6000 113.7000 331.8000 119.7000 ;
	    RECT 314.4000 102.6000 315.3000 107.7000 ;
	    RECT 316.2000 105.4500 317.4000 105.6000 ;
	    RECT 316.2000 104.5500 322.0500 105.4500 ;
	    RECT 316.2000 104.4000 317.4000 104.5500 ;
	    RECT 316.2000 103.2000 317.4000 103.5000 ;
	    RECT 246.9000 100.2000 251.4000 101.4000 ;
	    RECT 246.9000 99.3000 248.1000 100.2000 ;
	    RECT 232.2000 98.4000 239.1000 99.3000 ;
	    RECT 217.8000 93.3000 219.0000 98.1000 ;
	    RECT 244.2000 98.1000 248.1000 99.3000 ;
	    RECT 220.2000 93.3000 221.4000 97.5000 ;
	    RECT 222.6000 93.3000 223.8000 97.5000 ;
	    RECT 225.0000 93.3000 226.2000 97.5000 ;
	    RECT 227.4000 93.3000 228.6000 97.5000 ;
	    RECT 229.8000 93.3000 231.0000 96.3000 ;
	    RECT 232.2000 93.3000 233.4000 97.5000 ;
	    RECT 234.6000 93.3000 235.8000 96.3000 ;
	    RECT 237.0000 93.3000 238.2000 97.5000 ;
	    RECT 239.4000 93.3000 240.6000 97.5000 ;
	    RECT 241.8000 93.3000 243.0000 97.5000 ;
	    RECT 244.2000 93.3000 245.4000 98.1000 ;
	    RECT 249.0000 93.3000 250.2000 99.3000 ;
	    RECT 253.8000 93.3000 255.0000 102.3000 ;
	    RECT 277.8000 101.4000 279.0000 102.6000 ;
	    RECT 279.9000 100.8000 280.2000 102.3000 ;
	    RECT 282.3000 101.4000 284.1000 102.6000 ;
	    RECT 285.0000 102.4500 286.2000 102.6000 ;
	    RECT 309.0000 102.4500 310.2000 102.6000 ;
	    RECT 285.0000 101.5500 310.2000 102.4500 ;
	    RECT 285.0000 101.4000 286.2000 101.5500 ;
	    RECT 309.0000 101.4000 310.2000 101.5500 ;
	    RECT 311.4000 101.4000 312.6000 102.6000 ;
	    RECT 313.5000 101.4000 315.3000 102.6000 ;
	    RECT 317.4000 100.8000 317.7000 102.3000 ;
	    RECT 318.6000 101.4000 319.8000 102.6000 ;
	    RECT 321.1500 102.4500 322.0500 104.5500 ;
	    RECT 333.0000 103.5000 334.2000 119.7000 ;
	    RECT 393.1500 117.4500 394.0500 120.6000 ;
	    RECT 397.8000 117.4500 399.0000 117.6000 ;
	    RECT 429.0000 117.4500 430.2000 117.6000 ;
	    RECT 393.1500 116.5500 430.2000 117.4500 ;
	    RECT 397.8000 116.4000 399.0000 116.5500 ;
	    RECT 429.0000 116.4000 430.2000 116.5500 ;
	    RECT 465.0000 113.7000 466.2000 119.7000 ;
	    RECT 467.4000 114.6000 468.6000 119.7000 ;
	    RECT 467.1000 113.7000 468.6000 114.6000 ;
	    RECT 469.8000 113.7000 471.0000 120.6000 ;
	    RECT 467.1000 112.8000 468.0000 113.7000 ;
	    RECT 472.2000 112.8000 473.4000 119.7000 ;
	    RECT 474.6000 113.7000 475.8000 119.7000 ;
	    RECT 477.0000 115.5000 478.2000 119.7000 ;
	    RECT 479.4000 115.5000 480.6000 119.7000 ;
	    RECT 465.0000 111.9000 468.0000 112.8000 ;
	    RECT 465.0000 103.5000 466.2000 111.9000 ;
	    RECT 468.9000 111.6000 475.2000 112.8000 ;
	    RECT 481.8000 112.5000 483.0000 119.7000 ;
	    RECT 484.2000 113.7000 485.4000 119.7000 ;
	    RECT 486.6000 112.5000 487.8000 119.7000 ;
	    RECT 489.0000 113.7000 490.2000 119.7000 ;
	    RECT 468.9000 111.0000 469.8000 111.6000 ;
	    RECT 467.4000 109.8000 469.8000 111.0000 ;
	    RECT 474.3000 110.7000 483.0000 111.6000 ;
	    RECT 471.3000 109.8000 473.4000 110.7000 ;
	    RECT 471.3000 109.5000 480.6000 109.8000 ;
	    RECT 472.5000 108.9000 480.6000 109.5000 ;
	    RECT 479.4000 108.6000 480.6000 108.9000 ;
	    RECT 482.1000 109.5000 483.0000 110.7000 ;
	    RECT 483.9000 110.4000 487.8000 111.6000 ;
	    RECT 491.4000 110.4000 492.6000 119.7000 ;
	    RECT 493.8000 115.5000 495.0000 119.7000 ;
	    RECT 496.2000 115.5000 497.4000 119.7000 ;
	    RECT 498.6000 115.5000 499.8000 119.7000 ;
	    RECT 501.0000 113.7000 502.2000 119.7000 ;
	    RECT 496.2000 111.6000 502.5000 112.8000 ;
	    RECT 503.4000 111.6000 504.6000 119.7000 ;
	    RECT 505.8000 113.7000 507.0000 119.7000 ;
	    RECT 508.2000 112.8000 509.4000 119.7000 ;
	    RECT 510.6000 113.7000 511.8000 119.7000 ;
	    RECT 508.2000 111.9000 512.1000 112.8000 ;
	    RECT 513.0000 112.5000 514.2000 119.7000 ;
	    RECT 515.4000 113.7000 516.6000 119.7000 ;
	    RECT 647.4000 113.7000 648.6000 119.7000 ;
	    RECT 649.8000 112.5000 651.0000 119.7000 ;
	    RECT 652.2000 113.7000 653.4000 119.7000 ;
	    RECT 654.6000 112.8000 655.8000 119.7000 ;
	    RECT 657.0000 113.7000 658.2000 119.7000 ;
	    RECT 503.4000 110.4000 507.3000 111.6000 ;
	    RECT 493.8000 109.5000 495.0000 109.8000 ;
	    RECT 482.1000 108.6000 495.0000 109.5000 ;
	    RECT 498.6000 109.5000 499.8000 109.8000 ;
	    RECT 511.2000 109.5000 512.1000 111.9000 ;
	    RECT 651.9000 111.9000 655.8000 112.8000 ;
	    RECT 513.0000 110.4000 514.2000 111.6000 ;
	    RECT 577.8000 111.4500 579.0000 111.6000 ;
	    RECT 649.8000 111.4500 651.0000 111.6000 ;
	    RECT 577.8000 110.5500 651.0000 111.4500 ;
	    RECT 577.8000 110.4000 579.0000 110.5500 ;
	    RECT 649.8000 110.4000 651.0000 110.5500 ;
	    RECT 651.9000 109.5000 652.8000 111.9000 ;
	    RECT 659.4000 111.6000 660.6000 119.7000 ;
	    RECT 661.8000 113.7000 663.0000 119.7000 ;
	    RECT 664.2000 115.5000 665.4000 119.7000 ;
	    RECT 666.6000 115.5000 667.8000 119.7000 ;
	    RECT 669.0000 115.5000 670.2000 119.7000 ;
	    RECT 661.5000 111.6000 667.8000 112.8000 ;
	    RECT 656.7000 110.4000 660.6000 111.6000 ;
	    RECT 671.4000 110.4000 672.6000 119.7000 ;
	    RECT 673.8000 113.7000 675.0000 119.7000 ;
	    RECT 676.2000 112.5000 677.4000 119.7000 ;
	    RECT 678.6000 113.7000 679.8000 119.7000 ;
	    RECT 681.0000 112.5000 682.2000 119.7000 ;
	    RECT 683.4000 115.5000 684.6000 119.7000 ;
	    RECT 685.8000 115.5000 687.0000 119.7000 ;
	    RECT 688.2000 113.7000 689.4000 119.7000 ;
	    RECT 690.6000 112.8000 691.8000 119.7000 ;
	    RECT 693.0000 113.7000 694.2000 120.6000 ;
	    RECT 695.4000 114.6000 696.6000 119.7000 ;
	    RECT 695.4000 113.7000 696.9000 114.6000 ;
	    RECT 697.8000 113.7000 699.0000 119.7000 ;
	    RECT 722.7000 113.7000 723.9000 119.7000 ;
	    RECT 696.0000 112.8000 696.9000 113.7000 ;
	    RECT 688.8000 111.6000 695.1000 112.8000 ;
	    RECT 696.0000 111.9000 699.0000 112.8000 ;
	    RECT 676.2000 110.4000 680.1000 111.6000 ;
	    RECT 681.0000 110.7000 689.7000 111.6000 ;
	    RECT 694.2000 111.0000 695.1000 111.6000 ;
	    RECT 664.2000 109.5000 665.4000 109.8000 ;
	    RECT 498.6000 108.6000 512.1000 109.5000 ;
	    RECT 469.8000 107.4000 471.0000 108.6000 ;
	    RECT 474.9000 107.7000 476.1000 108.0000 ;
	    RECT 471.9000 106.8000 510.3000 107.7000 ;
	    RECT 509.1000 106.5000 510.3000 106.8000 ;
	    RECT 511.2000 105.9000 512.1000 108.6000 ;
	    RECT 513.0000 108.0000 514.2000 109.5000 ;
	    RECT 649.8000 108.0000 651.0000 109.5000 ;
	    RECT 513.0000 106.8000 514.5000 108.0000 ;
	    RECT 467.1000 105.0000 473.7000 105.9000 ;
	    RECT 467.1000 104.7000 468.3000 105.0000 ;
	    RECT 474.6000 104.4000 475.8000 105.6000 ;
	    RECT 476.7000 105.0000 502.2000 105.9000 ;
	    RECT 511.2000 105.0000 512.4000 105.9000 ;
	    RECT 501.0000 104.1000 502.2000 105.0000 ;
	    RECT 333.0000 102.4500 334.2000 102.6000 ;
	    RECT 321.1500 101.5500 334.2000 102.4500 ;
	    RECT 333.0000 101.4000 334.2000 101.5500 ;
	    RECT 465.0000 102.3000 478.2000 103.5000 ;
	    RECT 479.1000 102.9000 482.1000 104.1000 ;
	    RECT 487.8000 102.9000 492.6000 104.1000 ;
	    RECT 278.1000 99.3000 283.5000 99.9000 ;
	    RECT 285.0000 99.3000 285.9000 100.5000 ;
	    RECT 311.7000 99.3000 312.6000 100.5000 ;
	    RECT 314.1000 99.3000 319.5000 99.9000 ;
	    RECT 321.0000 99.4500 322.2000 99.6000 ;
	    RECT 330.6000 99.4500 331.8000 99.6000 ;
	    RECT 277.8000 99.0000 283.8000 99.3000 ;
	    RECT 277.8000 93.3000 279.0000 99.0000 ;
	    RECT 280.2000 93.3000 281.4000 98.1000 ;
	    RECT 282.6000 93.3000 283.8000 99.0000 ;
	    RECT 285.0000 93.3000 286.2000 99.3000 ;
	    RECT 311.4000 93.3000 312.6000 99.3000 ;
	    RECT 313.8000 99.0000 319.8000 99.3000 ;
	    RECT 313.8000 93.3000 315.0000 99.0000 ;
	    RECT 316.2000 93.3000 317.4000 98.1000 ;
	    RECT 318.6000 93.3000 319.8000 99.0000 ;
	    RECT 321.0000 98.5500 331.8000 99.4500 ;
	    RECT 321.0000 98.4000 322.2000 98.5500 ;
	    RECT 330.6000 98.4000 331.8000 98.5500 ;
	    RECT 330.6000 97.2000 331.8000 97.5000 ;
	    RECT 330.6000 93.3000 331.8000 96.3000 ;
	    RECT 333.0000 93.3000 334.2000 100.5000 ;
	    RECT 465.0000 93.3000 466.2000 102.3000 ;
	    RECT 468.6000 100.2000 473.1000 101.4000 ;
	    RECT 471.9000 99.3000 473.1000 100.2000 ;
	    RECT 480.9000 99.3000 482.1000 102.9000 ;
	    RECT 484.2000 101.4000 485.4000 102.6000 ;
	    RECT 492.0000 101.7000 493.2000 102.0000 ;
	    RECT 486.6000 100.8000 493.2000 101.7000 ;
	    RECT 486.6000 100.5000 487.8000 100.8000 ;
	    RECT 484.2000 100.2000 485.4000 100.5000 ;
	    RECT 496.2000 99.6000 497.4000 103.8000 ;
	    RECT 504.9000 102.9000 510.6000 104.1000 ;
	    RECT 504.9000 101.1000 506.1000 102.9000 ;
	    RECT 511.5000 102.0000 512.4000 105.0000 ;
	    RECT 486.6000 99.3000 487.8000 99.6000 ;
	    RECT 469.8000 93.3000 471.0000 99.3000 ;
	    RECT 471.9000 98.1000 475.8000 99.3000 ;
	    RECT 480.9000 98.4000 487.8000 99.3000 ;
	    RECT 489.0000 98.4000 490.2000 99.6000 ;
	    RECT 491.1000 98.4000 491.4000 99.6000 ;
	    RECT 495.9000 98.4000 497.4000 99.6000 ;
	    RECT 503.4000 100.2000 506.1000 101.1000 ;
	    RECT 510.6000 101.1000 512.4000 102.0000 ;
	    RECT 503.4000 99.3000 504.6000 100.2000 ;
	    RECT 474.6000 93.3000 475.8000 98.1000 ;
	    RECT 501.0000 98.1000 504.6000 99.3000 ;
	    RECT 477.0000 93.3000 478.2000 97.5000 ;
	    RECT 479.4000 93.3000 480.6000 97.5000 ;
	    RECT 481.8000 93.3000 483.0000 97.5000 ;
	    RECT 484.2000 93.3000 485.4000 96.3000 ;
	    RECT 486.6000 93.3000 487.8000 97.5000 ;
	    RECT 489.0000 93.3000 490.2000 96.3000 ;
	    RECT 491.4000 93.3000 492.6000 97.5000 ;
	    RECT 493.8000 93.3000 495.0000 97.5000 ;
	    RECT 496.2000 93.3000 497.4000 97.5000 ;
	    RECT 498.6000 93.3000 499.8000 97.5000 ;
	    RECT 501.0000 93.3000 502.2000 98.1000 ;
	    RECT 505.8000 93.3000 507.0000 99.3000 ;
	    RECT 510.6000 93.3000 511.8000 101.1000 ;
	    RECT 513.3000 100.2000 514.5000 106.8000 ;
	    RECT 513.0000 99.0000 514.5000 100.2000 ;
	    RECT 649.5000 106.8000 651.0000 108.0000 ;
	    RECT 651.9000 108.6000 665.4000 109.5000 ;
	    RECT 669.0000 109.5000 670.2000 109.8000 ;
	    RECT 681.0000 109.5000 681.9000 110.7000 ;
	    RECT 690.6000 109.8000 692.7000 110.7000 ;
	    RECT 694.2000 109.8000 696.6000 111.0000 ;
	    RECT 669.0000 108.6000 681.9000 109.5000 ;
	    RECT 683.4000 109.5000 692.7000 109.8000 ;
	    RECT 683.4000 108.9000 691.5000 109.5000 ;
	    RECT 683.4000 108.6000 684.6000 108.9000 ;
	    RECT 649.5000 100.2000 650.7000 106.8000 ;
	    RECT 651.9000 105.9000 652.8000 108.6000 ;
	    RECT 687.9000 107.7000 689.1000 108.0000 ;
	    RECT 653.7000 106.8000 692.1000 107.7000 ;
	    RECT 693.0000 107.4000 694.2000 108.6000 ;
	    RECT 653.7000 106.5000 654.9000 106.8000 ;
	    RECT 651.6000 105.0000 652.8000 105.9000 ;
	    RECT 661.8000 105.0000 687.3000 105.9000 ;
	    RECT 651.6000 102.0000 652.5000 105.0000 ;
	    RECT 661.8000 104.1000 663.0000 105.0000 ;
	    RECT 688.2000 104.4000 689.4000 105.6000 ;
	    RECT 690.3000 105.0000 696.9000 105.9000 ;
	    RECT 695.7000 104.7000 696.9000 105.0000 ;
	    RECT 653.4000 102.9000 659.1000 104.1000 ;
	    RECT 651.6000 101.1000 653.4000 102.0000 ;
	    RECT 649.5000 99.0000 651.0000 100.2000 ;
	    RECT 513.0000 93.3000 514.2000 99.0000 ;
	    RECT 515.4000 93.3000 516.6000 96.3000 ;
	    RECT 647.4000 93.3000 648.6000 96.3000 ;
	    RECT 649.8000 93.3000 651.0000 99.0000 ;
	    RECT 652.2000 93.3000 653.4000 101.1000 ;
	    RECT 657.9000 101.1000 659.1000 102.9000 ;
	    RECT 657.9000 100.2000 660.6000 101.1000 ;
	    RECT 659.4000 99.3000 660.6000 100.2000 ;
	    RECT 666.6000 99.6000 667.8000 103.8000 ;
	    RECT 671.4000 102.9000 676.2000 104.1000 ;
	    RECT 681.9000 102.9000 684.9000 104.1000 ;
	    RECT 697.8000 103.5000 699.0000 111.9000 ;
	    RECT 723.0000 110.4000 724.2000 111.6000 ;
	    RECT 723.0000 109.5000 723.9000 110.4000 ;
	    RECT 725.1000 108.6000 726.3000 119.7000 ;
	    RECT 721.8000 107.4000 723.0000 108.6000 ;
	    RECT 724.8000 107.7000 726.3000 108.6000 ;
	    RECT 729.0000 107.7000 730.2000 119.7000 ;
	    RECT 670.8000 101.7000 672.0000 102.0000 ;
	    RECT 670.8000 100.8000 677.4000 101.7000 ;
	    RECT 678.6000 101.4000 679.8000 102.6000 ;
	    RECT 676.2000 100.5000 677.4000 100.8000 ;
	    RECT 678.6000 100.2000 679.8000 100.5000 ;
	    RECT 657.0000 93.3000 658.2000 99.3000 ;
	    RECT 659.4000 98.1000 663.0000 99.3000 ;
	    RECT 666.6000 98.4000 668.1000 99.6000 ;
	    RECT 672.6000 98.4000 672.9000 99.6000 ;
	    RECT 673.8000 98.4000 675.0000 99.6000 ;
	    RECT 676.2000 99.3000 677.4000 99.6000 ;
	    RECT 681.9000 99.3000 683.1000 102.9000 ;
	    RECT 685.8000 102.3000 699.0000 103.5000 ;
	    RECT 724.8000 102.6000 725.7000 107.7000 ;
	    RECT 726.6000 105.4500 727.8000 105.6000 ;
	    RECT 726.6000 104.5500 732.4500 105.4500 ;
	    RECT 726.6000 104.4000 727.8000 104.5500 ;
	    RECT 726.6000 103.2000 727.8000 103.5000 ;
	    RECT 690.9000 100.2000 695.4000 101.4000 ;
	    RECT 690.9000 99.3000 692.1000 100.2000 ;
	    RECT 676.2000 98.4000 683.1000 99.3000 ;
	    RECT 661.8000 93.3000 663.0000 98.1000 ;
	    RECT 688.2000 98.1000 692.1000 99.3000 ;
	    RECT 664.2000 93.3000 665.4000 97.5000 ;
	    RECT 666.6000 93.3000 667.8000 97.5000 ;
	    RECT 669.0000 93.3000 670.2000 97.5000 ;
	    RECT 671.4000 93.3000 672.6000 97.5000 ;
	    RECT 673.8000 93.3000 675.0000 96.3000 ;
	    RECT 676.2000 93.3000 677.4000 97.5000 ;
	    RECT 678.6000 93.3000 679.8000 96.3000 ;
	    RECT 681.0000 93.3000 682.2000 97.5000 ;
	    RECT 683.4000 93.3000 684.6000 97.5000 ;
	    RECT 685.8000 93.3000 687.0000 97.5000 ;
	    RECT 688.2000 93.3000 689.4000 98.1000 ;
	    RECT 693.0000 93.3000 694.2000 99.3000 ;
	    RECT 697.8000 93.3000 699.0000 102.3000 ;
	    RECT 721.8000 101.4000 723.0000 102.6000 ;
	    RECT 723.9000 101.4000 725.7000 102.6000 ;
	    RECT 727.8000 100.8000 728.1000 102.3000 ;
	    RECT 729.0000 101.4000 730.2000 102.6000 ;
	    RECT 731.5500 102.4500 732.4500 104.5500 ;
	    RECT 743.4000 103.5000 744.6000 119.7000 ;
	    RECT 745.8000 113.7000 747.0000 119.7000 ;
	    RECT 772.2000 108.6000 773.4000 119.7000 ;
	    RECT 774.6000 109.5000 775.8000 119.7000 ;
	    RECT 777.0000 108.6000 778.2000 119.7000 ;
	    RECT 772.2000 107.7000 778.2000 108.6000 ;
	    RECT 779.4000 107.7000 780.6000 119.7000 ;
	    RECT 798.6000 113.7000 799.8000 119.7000 ;
	    RECT 779.4000 106.5000 780.3000 107.7000 ;
	    RECT 801.0000 106.5000 802.2000 119.7000 ;
	    RECT 803.4000 113.7000 804.6000 119.7000 ;
	    RECT 805.8000 119.4000 807.0000 120.6000 ;
	    RECT 935.4000 113.7000 936.6000 119.7000 ;
	    RECT 937.8000 114.6000 939.0000 119.7000 ;
	    RECT 937.5000 113.7000 939.0000 114.6000 ;
	    RECT 940.2000 113.7000 941.4000 120.6000 ;
	    RECT 937.5000 112.8000 938.4000 113.7000 ;
	    RECT 942.6000 112.8000 943.8000 119.7000 ;
	    RECT 945.0000 113.7000 946.2000 119.7000 ;
	    RECT 947.4000 115.5000 948.6000 119.7000 ;
	    RECT 949.8000 115.5000 951.0000 119.7000 ;
	    RECT 935.4000 111.9000 938.4000 112.8000 ;
	    RECT 803.4000 109.5000 804.6000 109.8000 ;
	    RECT 803.4000 108.4500 804.6000 108.6000 ;
	    RECT 805.8000 108.4500 807.0000 108.6000 ;
	    RECT 803.4000 107.5500 807.0000 108.4500 ;
	    RECT 803.4000 107.4000 804.6000 107.5500 ;
	    RECT 805.8000 107.4000 807.0000 107.5500 ;
	    RECT 772.2000 104.4000 773.4000 105.6000 ;
	    RECT 774.3000 104.7000 774.6000 106.2000 ;
	    RECT 777.0000 104.7000 778.5000 105.6000 ;
	    RECT 779.4000 105.4500 780.6000 105.6000 ;
	    RECT 791.4000 105.4500 792.6000 105.6000 ;
	    RECT 774.6000 103.5000 775.8000 103.8000 ;
	    RECT 743.4000 102.4500 744.6000 102.6000 ;
	    RECT 731.5500 101.5500 744.6000 102.4500 ;
	    RECT 743.4000 101.4000 744.6000 101.5500 ;
	    RECT 774.6000 101.4000 775.8000 102.6000 ;
	    RECT 722.1000 99.3000 723.0000 100.5000 ;
	    RECT 724.5000 99.3000 729.9000 99.9000 ;
	    RECT 721.8000 93.3000 723.0000 99.3000 ;
	    RECT 724.2000 99.0000 730.2000 99.3000 ;
	    RECT 724.2000 93.3000 725.4000 99.0000 ;
	    RECT 726.6000 93.3000 727.8000 98.1000 ;
	    RECT 729.0000 93.3000 730.2000 99.0000 ;
	    RECT 743.4000 93.3000 744.6000 100.5000 ;
	    RECT 745.8000 99.4500 747.0000 99.6000 ;
	    RECT 769.8000 99.4500 771.0000 99.6000 ;
	    RECT 745.8000 98.5500 771.0000 99.4500 ;
	    RECT 777.0000 99.3000 777.9000 104.7000 ;
	    RECT 779.4000 104.5500 792.6000 105.4500 ;
	    RECT 779.4000 104.4000 780.6000 104.5500 ;
	    RECT 791.4000 104.4000 792.6000 104.5500 ;
	    RECT 793.8000 105.4500 795.0000 105.6000 ;
	    RECT 801.0000 105.4500 802.2000 105.6000 ;
	    RECT 793.8000 104.5500 802.2000 105.4500 ;
	    RECT 793.8000 104.4000 795.0000 104.5500 ;
	    RECT 801.0000 104.4000 802.2000 104.5500 ;
	    RECT 935.4000 103.5000 936.6000 111.9000 ;
	    RECT 939.3000 111.6000 945.6000 112.8000 ;
	    RECT 952.2000 112.5000 953.4000 119.7000 ;
	    RECT 954.6000 113.7000 955.8000 119.7000 ;
	    RECT 957.0000 112.5000 958.2000 119.7000 ;
	    RECT 959.4000 113.7000 960.6000 119.7000 ;
	    RECT 939.3000 111.0000 940.2000 111.6000 ;
	    RECT 937.8000 109.8000 940.2000 111.0000 ;
	    RECT 944.7000 110.7000 953.4000 111.6000 ;
	    RECT 941.7000 109.8000 943.8000 110.7000 ;
	    RECT 941.7000 109.5000 951.0000 109.8000 ;
	    RECT 942.9000 108.9000 951.0000 109.5000 ;
	    RECT 949.8000 108.6000 951.0000 108.9000 ;
	    RECT 952.5000 109.5000 953.4000 110.7000 ;
	    RECT 954.3000 110.4000 958.2000 111.6000 ;
	    RECT 961.8000 110.4000 963.0000 119.7000 ;
	    RECT 964.2000 115.5000 965.4000 119.7000 ;
	    RECT 966.6000 115.5000 967.8000 119.7000 ;
	    RECT 969.0000 115.5000 970.2000 119.7000 ;
	    RECT 971.4000 113.7000 972.6000 119.7000 ;
	    RECT 966.6000 111.6000 972.9000 112.8000 ;
	    RECT 973.8000 111.6000 975.0000 119.7000 ;
	    RECT 976.2000 113.7000 977.4000 119.7000 ;
	    RECT 978.6000 112.8000 979.8000 119.7000 ;
	    RECT 981.0000 113.7000 982.2000 119.7000 ;
	    RECT 978.6000 111.9000 982.5000 112.8000 ;
	    RECT 983.4000 112.5000 984.6000 119.7000 ;
	    RECT 985.8000 113.7000 987.0000 119.7000 ;
	    RECT 973.8000 110.4000 977.7000 111.6000 ;
	    RECT 964.2000 109.5000 965.4000 109.8000 ;
	    RECT 952.5000 108.6000 965.4000 109.5000 ;
	    RECT 969.0000 109.5000 970.2000 109.8000 ;
	    RECT 981.6000 109.5000 982.5000 111.9000 ;
	    RECT 983.4000 110.4000 984.6000 111.6000 ;
	    RECT 969.0000 108.6000 982.5000 109.5000 ;
	    RECT 940.2000 107.4000 941.4000 108.6000 ;
	    RECT 945.3000 107.7000 946.5000 108.0000 ;
	    RECT 942.3000 106.8000 980.7000 107.7000 ;
	    RECT 979.5000 106.5000 980.7000 106.8000 ;
	    RECT 981.6000 105.9000 982.5000 108.6000 ;
	    RECT 983.4000 108.0000 984.6000 109.5000 ;
	    RECT 983.4000 106.8000 984.9000 108.0000 ;
	    RECT 937.5000 105.0000 944.1000 105.9000 ;
	    RECT 937.5000 104.7000 938.7000 105.0000 ;
	    RECT 945.0000 104.4000 946.2000 105.6000 ;
	    RECT 947.1000 105.0000 972.6000 105.9000 ;
	    RECT 981.6000 105.0000 982.8000 105.9000 ;
	    RECT 971.4000 104.1000 972.6000 105.0000 ;
	    RECT 798.6000 101.4000 799.8000 102.6000 ;
	    RECT 798.6000 100.2000 799.8000 100.5000 ;
	    RECT 779.4000 99.4500 780.6000 99.6000 ;
	    RECT 781.8000 99.4500 783.0000 99.6000 ;
	    RECT 745.8000 98.4000 747.0000 98.5500 ;
	    RECT 769.8000 98.4000 771.0000 98.5500 ;
	    RECT 745.8000 97.2000 747.0000 97.5000 ;
	    RECT 745.8000 93.3000 747.0000 96.3000 ;
	    RECT 773.1000 93.3000 774.3000 99.3000 ;
	    RECT 777.0000 93.3000 778.2000 99.3000 ;
	    RECT 779.4000 98.5500 783.0000 99.4500 ;
	    RECT 801.0000 99.3000 802.2000 103.5000 ;
	    RECT 935.4000 102.3000 948.6000 103.5000 ;
	    RECT 949.5000 102.9000 952.5000 104.1000 ;
	    RECT 958.2000 102.9000 963.0000 104.1000 ;
	    RECT 779.4000 98.4000 780.6000 98.5500 ;
	    RECT 781.8000 98.4000 783.0000 98.5500 ;
	    RECT 779.1000 97.2000 780.3000 97.5000 ;
	    RECT 779.4000 93.3000 780.6000 96.3000 ;
	    RECT 798.6000 93.3000 799.8000 99.3000 ;
	    RECT 801.0000 98.4000 803.7000 99.3000 ;
	    RECT 802.5000 93.3000 803.7000 98.4000 ;
	    RECT 935.4000 93.3000 936.6000 102.3000 ;
	    RECT 939.0000 100.2000 943.5000 101.4000 ;
	    RECT 942.3000 99.3000 943.5000 100.2000 ;
	    RECT 951.3000 99.3000 952.5000 102.9000 ;
	    RECT 954.6000 101.4000 955.8000 102.6000 ;
	    RECT 962.4000 101.7000 963.6000 102.0000 ;
	    RECT 957.0000 100.8000 963.6000 101.7000 ;
	    RECT 957.0000 100.5000 958.2000 100.8000 ;
	    RECT 954.6000 100.2000 955.8000 100.5000 ;
	    RECT 966.6000 99.6000 967.8000 103.8000 ;
	    RECT 975.3000 102.9000 981.0000 104.1000 ;
	    RECT 975.3000 101.1000 976.5000 102.9000 ;
	    RECT 981.9000 102.0000 982.8000 105.0000 ;
	    RECT 957.0000 99.3000 958.2000 99.6000 ;
	    RECT 940.2000 93.3000 941.4000 99.3000 ;
	    RECT 942.3000 98.1000 946.2000 99.3000 ;
	    RECT 951.3000 98.4000 958.2000 99.3000 ;
	    RECT 959.4000 98.4000 960.6000 99.6000 ;
	    RECT 961.5000 98.4000 961.8000 99.6000 ;
	    RECT 966.3000 98.4000 967.8000 99.6000 ;
	    RECT 973.8000 100.2000 976.5000 101.1000 ;
	    RECT 981.0000 101.1000 982.8000 102.0000 ;
	    RECT 973.8000 99.3000 975.0000 100.2000 ;
	    RECT 945.0000 93.3000 946.2000 98.1000 ;
	    RECT 971.4000 98.1000 975.0000 99.3000 ;
	    RECT 947.4000 93.3000 948.6000 97.5000 ;
	    RECT 949.8000 93.3000 951.0000 97.5000 ;
	    RECT 952.2000 93.3000 953.4000 97.5000 ;
	    RECT 954.6000 93.3000 955.8000 96.3000 ;
	    RECT 957.0000 93.3000 958.2000 97.5000 ;
	    RECT 959.4000 93.3000 960.6000 96.3000 ;
	    RECT 961.8000 93.3000 963.0000 97.5000 ;
	    RECT 964.2000 93.3000 965.4000 97.5000 ;
	    RECT 966.6000 93.3000 967.8000 97.5000 ;
	    RECT 969.0000 93.3000 970.2000 97.5000 ;
	    RECT 971.4000 93.3000 972.6000 98.1000 ;
	    RECT 976.2000 93.3000 977.4000 99.3000 ;
	    RECT 981.0000 93.3000 982.2000 101.1000 ;
	    RECT 983.7000 100.2000 984.9000 106.8000 ;
	    RECT 1000.2000 103.5000 1001.4000 119.7000 ;
	    RECT 1002.6000 113.7000 1003.8000 119.7000 ;
	    RECT 1072.2001 107.1000 1073.4000 119.7000 ;
	    RECT 1074.6000 108.0000 1075.8000 119.7000 ;
	    RECT 1078.8000 114.6000 1080.0000 119.7000 ;
	    RECT 1077.0000 113.7000 1080.0000 114.6000 ;
	    RECT 1083.0000 113.7000 1084.2001 119.7000 ;
	    RECT 1085.4000 113.7000 1086.6000 119.7000 ;
	    RECT 1087.8000 113.7000 1089.0000 119.7000 ;
	    RECT 1091.7001 113.7000 1093.5000 119.7000 ;
	    RECT 1077.0000 112.5000 1078.2001 113.7000 ;
	    RECT 1085.4000 112.8000 1086.3000 113.7000 ;
	    RECT 1082.1000 111.9000 1087.5000 112.8000 ;
	    RECT 1091.4000 112.5000 1092.6000 113.7000 ;
	    RECT 1082.1000 111.6000 1083.3000 111.9000 ;
	    RECT 1086.3000 111.6000 1087.5000 111.9000 ;
	    RECT 1077.0000 109.5000 1078.2001 109.8000 ;
	    RECT 1083.9000 109.5000 1085.1000 109.8000 ;
	    RECT 1077.0000 108.6000 1085.1000 109.5000 ;
	    RECT 1086.0000 109.5000 1089.3000 110.4000 ;
	    RECT 1086.0000 107.7000 1086.9000 109.5000 ;
	    RECT 1088.1000 109.2000 1089.3000 109.5000 ;
	    RECT 1091.7001 109.8000 1093.8000 111.0000 ;
	    RECT 1091.7001 108.3000 1092.6000 109.8000 ;
	    RECT 1079.7001 107.1000 1086.9000 107.7000 ;
	    RECT 1072.2001 106.8000 1086.9000 107.1000 ;
	    RECT 1089.0000 107.4000 1092.6000 108.3000 ;
	    RECT 1096.2001 107.7000 1097.4000 119.7000 ;
	    RECT 1072.2001 106.5000 1080.9000 106.8000 ;
	    RECT 1072.2001 106.2000 1080.6000 106.5000 ;
	    RECT 1075.5000 104.4000 1080.9000 105.3000 ;
	    RECT 1081.8000 104.4000 1083.0000 105.6000 ;
	    RECT 1075.5000 104.1000 1076.7001 104.4000 ;
	    RECT 1077.9000 102.6000 1079.1000 102.9000 ;
	    RECT 1089.0000 102.6000 1089.9000 107.4000 ;
	    RECT 1098.6000 106.8000 1099.8000 119.7000 ;
	    RECT 1113.0000 113.7000 1114.2001 119.7000 ;
	    RECT 1093.5000 106.5000 1099.8000 106.8000 ;
	    RECT 1093.5000 105.9000 1097.7001 106.5000 ;
	    RECT 1093.5000 105.6000 1094.7001 105.9000 ;
	    RECT 1098.6000 105.4500 1099.8000 105.6000 ;
	    RECT 1110.6000 105.4500 1111.8000 105.6000 ;
	    RECT 1095.9000 104.7000 1097.1000 105.0000 ;
	    RECT 1091.4000 103.8000 1097.1000 104.7000 ;
	    RECT 1098.6000 104.5500 1111.8000 105.4500 ;
	    RECT 1098.6000 104.4000 1099.8000 104.5500 ;
	    RECT 1110.6000 104.4000 1111.8000 104.5500 ;
	    RECT 1091.4000 103.5000 1092.6000 103.8000 ;
	    RECT 1115.4000 103.5000 1116.6000 119.7000 ;
	    RECT 1139.4000 108.4500 1140.6000 108.6000 ;
	    RECT 1144.2001 108.4500 1145.4000 108.6000 ;
	    RECT 1139.4000 107.5500 1145.4000 108.4500 ;
	    RECT 1146.6000 107.7000 1147.8000 119.7000 ;
	    RECT 1150.5000 108.6000 1151.7001 119.7000 ;
	    RECT 1152.9000 113.7000 1154.1000 119.7000 ;
	    RECT 1152.6000 110.4000 1153.8000 111.6000 ;
	    RECT 1152.9000 109.5000 1153.8000 110.4000 ;
	    RECT 1150.5000 107.7000 1152.0000 108.6000 ;
	    RECT 1139.4000 107.4000 1140.6000 107.5500 ;
	    RECT 1144.2001 107.4000 1145.4000 107.5500 ;
	    RECT 1149.0000 105.4500 1150.2001 105.6000 ;
	    RECT 1144.3500 104.5500 1150.2001 105.4500 ;
	    RECT 1000.2000 102.4500 1001.4000 102.6000 ;
	    RECT 1012.2000 102.4500 1013.4000 102.6000 ;
	    RECT 1000.2000 101.5500 1013.4000 102.4500 ;
	    RECT 1000.2000 101.4000 1001.4000 101.5500 ;
	    RECT 1012.2000 101.4000 1013.4000 101.5500 ;
	    RECT 1073.4000 101.4000 1073.7001 102.6000 ;
	    RECT 1074.6000 101.4000 1075.8000 102.6000 ;
	    RECT 1076.7001 101.7000 1089.9000 102.6000 ;
	    RECT 983.4000 99.0000 984.9000 100.2000 ;
	    RECT 983.4000 93.3000 984.6000 99.0000 ;
	    RECT 985.8000 93.3000 987.0000 96.3000 ;
	    RECT 1000.2000 93.3000 1001.4000 100.5000 ;
	    RECT 1002.6000 99.4500 1003.8000 99.6000 ;
	    RECT 1069.8000 99.4500 1071.0000 99.6000 ;
	    RECT 1002.6000 98.5500 1071.0000 99.4500 ;
	    RECT 1002.6000 98.4000 1003.8000 98.5500 ;
	    RECT 1069.8000 98.4000 1071.0000 98.5500 ;
	    RECT 1002.6000 97.2000 1003.8000 97.5000 ;
	    RECT 1002.6000 93.3000 1003.8000 96.3000 ;
	    RECT 1072.2001 93.3000 1073.4000 100.5000 ;
	    RECT 1074.6000 93.3000 1075.8000 99.3000 ;
	    RECT 1079.7001 98.4000 1080.6000 101.7000 ;
	    RECT 1088.1000 101.4000 1089.3000 101.7000 ;
	    RECT 1098.6000 100.8000 1099.8000 103.5000 ;
	    RECT 1115.4000 102.4500 1116.6000 102.6000 ;
	    RECT 1144.3500 102.4500 1145.2500 104.5500 ;
	    RECT 1149.0000 104.4000 1150.2001 104.5500 ;
	    RECT 1149.0000 103.2000 1150.2001 103.5000 ;
	    RECT 1151.1000 102.6000 1152.0000 107.7000 ;
	    RECT 1153.8000 108.4500 1155.0000 108.6000 ;
	    RECT 1170.6000 108.4500 1171.8000 108.6000 ;
	    RECT 1153.8000 107.5500 1171.8000 108.4500 ;
	    RECT 1177.8000 107.7000 1179.0000 119.7000 ;
	    RECT 1181.7001 108.6000 1182.9000 119.7000 ;
	    RECT 1184.1000 113.7000 1185.3000 119.7000 ;
	    RECT 1209.9000 113.7000 1211.1000 119.7000 ;
	    RECT 1183.8000 110.4000 1185.0000 111.6000 ;
	    RECT 1184.1000 109.5000 1185.0000 110.4000 ;
	    RECT 1210.2001 110.4000 1211.4000 111.6000 ;
	    RECT 1210.2001 109.5000 1211.1000 110.4000 ;
	    RECT 1212.3000 108.6000 1213.5000 119.7000 ;
	    RECT 1181.7001 107.7000 1183.2001 108.6000 ;
	    RECT 1153.8000 107.4000 1155.0000 107.5500 ;
	    RECT 1170.6000 107.4000 1171.8000 107.5500 ;
	    RECT 1156.2001 105.4500 1157.4000 105.6000 ;
	    RECT 1177.8000 105.4500 1179.0000 105.6000 ;
	    RECT 1156.2001 104.5500 1179.0000 105.4500 ;
	    RECT 1156.2001 104.4000 1157.4000 104.5500 ;
	    RECT 1177.8000 104.4000 1179.0000 104.5500 ;
	    RECT 1180.2001 104.4000 1181.4000 105.6000 ;
	    RECT 1180.2001 103.2000 1181.4000 103.5000 ;
	    RECT 1182.3000 102.6000 1183.2001 107.7000 ;
	    RECT 1185.0000 107.4000 1186.2001 108.6000 ;
	    RECT 1209.0000 107.4000 1210.2001 108.6000 ;
	    RECT 1212.0000 107.7000 1213.5000 108.6000 ;
	    RECT 1216.2001 107.7000 1217.4000 119.7000 ;
	    RECT 1235.4000 113.7000 1236.6000 119.7000 ;
	    RECT 1212.0000 102.6000 1212.9000 107.7000 ;
	    RECT 1237.8000 106.5000 1239.0000 119.7000 ;
	    RECT 1240.2001 113.7000 1241.4000 119.7000 ;
	    RECT 1269.0000 118.8000 1275.0000 119.7000 ;
	    RECT 1240.2001 109.5000 1241.4000 109.8000 ;
	    RECT 1240.2001 107.4000 1241.4000 108.6000 ;
	    RECT 1245.0000 108.4500 1246.2001 108.6000 ;
	    RECT 1266.6000 108.4500 1267.8000 108.6000 ;
	    RECT 1245.0000 107.5500 1267.8000 108.4500 ;
	    RECT 1269.0000 107.7000 1270.2001 118.8000 ;
	    RECT 1271.4000 107.7000 1272.6000 117.9000 ;
	    RECT 1273.8000 108.6000 1275.0000 118.8000 ;
	    RECT 1276.2001 109.5000 1277.4000 119.7000 ;
	    RECT 1278.6000 108.6000 1279.8000 119.7000 ;
	    RECT 1273.8000 107.7000 1279.8000 108.6000 ;
	    RECT 1321.8000 108.6000 1323.0000 119.7000 ;
	    RECT 1324.2001 109.8000 1325.7001 119.7000 ;
	    RECT 1324.2001 108.6000 1325.4000 108.9000 ;
	    RECT 1321.8000 107.7000 1325.4000 108.6000 ;
	    RECT 1328.4000 107.7000 1330.8000 119.7000 ;
	    RECT 1333.5000 109.8000 1335.0000 119.7000 ;
	    RECT 1333.5000 108.6000 1334.7001 108.9000 ;
	    RECT 1336.2001 108.6000 1337.4000 119.7000 ;
	    RECT 1444.2001 119.4000 1445.4000 120.6000 ;
	    RECT 1468.2001 113.7000 1469.4000 119.7000 ;
	    RECT 1470.6000 112.5000 1471.8000 119.7000 ;
	    RECT 1473.0000 113.7000 1474.2001 119.7000 ;
	    RECT 1475.4000 112.8000 1476.6000 119.7000 ;
	    RECT 1477.8000 113.7000 1479.0000 119.7000 ;
	    RECT 1472.7001 111.9000 1476.6000 112.8000 ;
	    RECT 1453.8000 111.4500 1455.0000 111.6000 ;
	    RECT 1470.6000 111.4500 1471.8000 111.6000 ;
	    RECT 1453.8000 110.5500 1471.8000 111.4500 ;
	    RECT 1453.8000 110.4000 1455.0000 110.5500 ;
	    RECT 1470.6000 110.4000 1471.8000 110.5500 ;
	    RECT 1472.7001 109.5000 1473.6000 111.9000 ;
	    RECT 1480.2001 111.6000 1481.4000 119.7000 ;
	    RECT 1482.6000 113.7000 1483.8000 119.7000 ;
	    RECT 1485.0000 115.5000 1486.2001 119.7000 ;
	    RECT 1487.4000 115.5000 1488.6000 119.7000 ;
	    RECT 1489.8000 115.5000 1491.0000 119.7000 ;
	    RECT 1482.3000 111.6000 1488.6000 112.8000 ;
	    RECT 1477.5000 110.4000 1481.4000 111.6000 ;
	    RECT 1492.2001 110.4000 1493.4000 119.7000 ;
	    RECT 1494.6000 113.7000 1495.8000 119.7000 ;
	    RECT 1497.0000 112.5000 1498.2001 119.7000 ;
	    RECT 1499.4000 113.7000 1500.6000 119.7000 ;
	    RECT 1501.8000 112.5000 1503.0000 119.7000 ;
	    RECT 1504.2001 115.5000 1505.4000 119.7000 ;
	    RECT 1506.6000 115.5000 1507.8000 119.7000 ;
	    RECT 1509.0000 113.7000 1510.2001 119.7000 ;
	    RECT 1511.4000 112.8000 1512.6000 119.7000 ;
	    RECT 1513.8000 113.7000 1515.0000 120.6000 ;
	    RECT 1516.2001 114.6000 1517.4000 119.7000 ;
	    RECT 1516.2001 113.7000 1517.7001 114.6000 ;
	    RECT 1518.6000 113.7000 1519.8000 119.7000 ;
	    RECT 1516.8000 112.8000 1517.7001 113.7000 ;
	    RECT 1509.6000 111.6000 1515.9000 112.8000 ;
	    RECT 1516.8000 111.9000 1519.8000 112.8000 ;
	    RECT 1497.0000 110.4000 1500.9000 111.6000 ;
	    RECT 1501.8000 110.7000 1510.5000 111.6000 ;
	    RECT 1515.0000 111.0000 1515.9000 111.6000 ;
	    RECT 1485.0000 109.5000 1486.2001 109.8000 ;
	    RECT 1333.5000 107.7000 1337.4000 108.6000 ;
	    RECT 1470.6000 108.0000 1471.8000 109.5000 ;
	    RECT 1245.0000 107.4000 1246.2001 107.5500 ;
	    RECT 1266.6000 107.4000 1267.8000 107.5500 ;
	    RECT 1271.7001 106.8000 1272.6000 107.7000 ;
	    RECT 1269.0000 106.5000 1270.2001 106.8000 ;
	    RECT 1271.7001 106.5000 1274.7001 106.8000 ;
	    RECT 1329.0000 106.5000 1329.9000 107.7000 ;
	    RECT 1470.3000 106.8000 1471.8000 108.0000 ;
	    RECT 1472.7001 108.6000 1486.2001 109.5000 ;
	    RECT 1489.8000 109.5000 1491.0000 109.8000 ;
	    RECT 1501.8000 109.5000 1502.7001 110.7000 ;
	    RECT 1511.4000 109.8000 1513.5000 110.7000 ;
	    RECT 1515.0000 109.8000 1517.4000 111.0000 ;
	    RECT 1489.8000 108.6000 1502.7001 109.5000 ;
	    RECT 1504.2001 109.5000 1513.5000 109.8000 ;
	    RECT 1504.2001 108.9000 1512.3000 109.5000 ;
	    RECT 1504.2001 108.6000 1505.4000 108.9000 ;
	    RECT 1271.7001 105.9000 1272.9000 106.5000 ;
	    RECT 1213.8000 104.4000 1215.0000 105.6000 ;
	    RECT 1237.8000 105.4500 1239.0000 105.6000 ;
	    RECT 1266.6000 105.4500 1267.8000 105.6000 ;
	    RECT 1237.8000 104.5500 1267.8000 105.4500 ;
	    RECT 1237.8000 104.4000 1239.0000 104.5500 ;
	    RECT 1266.6000 104.4000 1267.8000 104.5500 ;
	    RECT 1269.0000 104.4000 1270.2001 105.6000 ;
	    RECT 1273.8000 104.4000 1275.0000 105.6000 ;
	    RECT 1277.4000 104.7000 1277.7001 106.2000 ;
	    RECT 1331.7001 105.6000 1332.9000 105.9000 ;
	    RECT 1278.6000 104.4000 1279.8000 105.6000 ;
	    RECT 1329.0000 104.4000 1330.2001 105.6000 ;
	    RECT 1331.7001 104.7000 1334.1000 105.6000 ;
	    RECT 1332.9000 104.4000 1334.1000 104.7000 ;
	    RECT 1271.7001 103.5000 1272.9000 104.4000 ;
	    RECT 1276.2001 103.5000 1277.4000 103.8000 ;
	    RECT 1213.8000 103.2000 1215.0000 103.5000 ;
	    RECT 1115.4000 101.5500 1145.2500 102.4500 ;
	    RECT 1115.4000 101.4000 1116.6000 101.5500 ;
	    RECT 1146.6000 101.4000 1147.8000 102.6000 ;
	    RECT 1148.7001 100.8000 1149.0000 102.3000 ;
	    RECT 1151.1000 101.4000 1152.9000 102.6000 ;
	    RECT 1153.8000 102.4500 1155.0000 102.6000 ;
	    RECT 1158.6000 102.4500 1159.8000 102.6000 ;
	    RECT 1153.8000 101.5500 1159.8000 102.4500 ;
	    RECT 1153.8000 101.4000 1155.0000 101.5500 ;
	    RECT 1158.6000 101.4000 1159.8000 101.5500 ;
	    RECT 1168.2001 102.4500 1169.4000 102.6000 ;
	    RECT 1175.4000 102.4500 1176.6000 102.6000 ;
	    RECT 1177.8000 102.4500 1179.0000 102.6000 ;
	    RECT 1168.2001 101.5500 1179.0000 102.4500 ;
	    RECT 1168.2001 101.4000 1169.4000 101.5500 ;
	    RECT 1175.4000 101.4000 1176.6000 101.5500 ;
	    RECT 1177.8000 101.4000 1179.0000 101.5500 ;
	    RECT 1179.9000 100.8000 1180.2001 102.3000 ;
	    RECT 1182.3000 101.4000 1184.1000 102.6000 ;
	    RECT 1185.0000 102.4500 1186.2001 102.6000 ;
	    RECT 1206.6000 102.4500 1207.8000 102.6000 ;
	    RECT 1185.0000 101.5500 1207.8000 102.4500 ;
	    RECT 1185.0000 101.4000 1186.2001 101.5500 ;
	    RECT 1206.6000 101.4000 1207.8000 101.5500 ;
	    RECT 1209.0000 101.4000 1210.2001 102.6000 ;
	    RECT 1211.1000 101.4000 1212.9000 102.6000 ;
	    RECT 1216.2001 102.4500 1217.4000 102.6000 ;
	    RECT 1233.0000 102.4500 1234.2001 102.6000 ;
	    RECT 1215.0000 100.8000 1215.3000 102.3000 ;
	    RECT 1216.2001 101.5500 1234.2001 102.4500 ;
	    RECT 1216.2001 101.4000 1217.4000 101.5500 ;
	    RECT 1233.0000 101.4000 1234.2001 101.5500 ;
	    RECT 1235.4000 101.4000 1236.6000 102.6000 ;
	    RECT 1094.1000 99.9000 1099.8000 100.8000 ;
	    RECT 1094.1000 99.6000 1095.3000 99.9000 ;
	    RECT 1077.0000 96.3000 1078.2001 97.5000 ;
	    RECT 1079.4000 97.2000 1080.6000 98.4000 ;
	    RECT 1082.1000 98.1000 1083.3000 98.4000 ;
	    RECT 1082.1000 97.2000 1086.3000 98.1000 ;
	    RECT 1085.4000 96.3000 1086.3000 97.2000 ;
	    RECT 1091.4000 96.3000 1092.6000 97.5000 ;
	    RECT 1077.0000 95.4000 1080.0000 96.3000 ;
	    RECT 1078.8000 93.3000 1080.0000 95.4000 ;
	    RECT 1082.7001 93.3000 1084.2001 96.3000 ;
	    RECT 1085.4000 93.3000 1086.6000 96.3000 ;
	    RECT 1087.8000 93.3000 1089.0000 96.3000 ;
	    RECT 1091.4000 95.4000 1093.5000 96.3000 ;
	    RECT 1091.7001 93.3000 1093.5000 95.4000 ;
	    RECT 1096.2001 93.3000 1097.4000 99.0000 ;
	    RECT 1098.6000 93.3000 1099.8000 99.9000 ;
	    RECT 1113.0000 98.4000 1114.2001 99.6000 ;
	    RECT 1113.0000 97.2000 1114.2001 97.5000 ;
	    RECT 1113.0000 93.3000 1114.2001 96.3000 ;
	    RECT 1115.4000 93.3000 1116.6000 100.5000 ;
	    RECT 1146.9000 99.3000 1152.3000 99.9000 ;
	    RECT 1153.8000 99.3000 1154.7001 100.5000 ;
	    RECT 1178.1000 99.3000 1183.5000 99.9000 ;
	    RECT 1185.0000 99.3000 1185.9000 100.5000 ;
	    RECT 1209.3000 99.3000 1210.2001 100.5000 ;
	    RECT 1235.4000 100.2000 1236.6000 100.5000 ;
	    RECT 1211.7001 99.3000 1217.1000 99.9000 ;
	    RECT 1237.8000 99.3000 1239.0000 103.5000 ;
	    RECT 1247.4000 102.4500 1248.6000 102.6000 ;
	    RECT 1271.4000 102.4500 1272.6000 102.6000 ;
	    RECT 1247.4000 101.5500 1272.6000 102.4500 ;
	    RECT 1247.4000 101.4000 1248.6000 101.5500 ;
	    RECT 1271.4000 101.4000 1272.6000 101.5500 ;
	    RECT 1273.8000 99.3000 1274.7001 103.5000 ;
	    RECT 1329.0000 102.6000 1329.9000 103.5000 ;
	    RECT 1276.2001 101.4000 1277.4000 102.6000 ;
	    RECT 1307.4000 102.4500 1308.6000 102.6000 ;
	    RECT 1321.8000 102.4500 1323.0000 102.6000 ;
	    RECT 1307.4000 101.5500 1323.0000 102.4500 ;
	    RECT 1307.4000 101.4000 1308.6000 101.5500 ;
	    RECT 1321.8000 101.4000 1323.0000 101.5500 ;
	    RECT 1323.9000 101.4000 1324.2001 102.6000 ;
	    RECT 1326.0000 101.4000 1327.2001 102.6000 ;
	    RECT 1326.3000 100.8000 1327.2001 101.4000 ;
	    RECT 1328.4000 101.7000 1329.9000 102.6000 ;
	    RECT 1330.8000 102.9000 1332.0000 103.2000 ;
	    RECT 1330.8000 102.6000 1335.0000 102.9000 ;
	    RECT 1330.8000 102.0000 1335.3000 102.6000 ;
	    RECT 1334.1000 101.7000 1335.3000 102.0000 ;
	    RECT 1324.2001 100.2000 1325.4000 100.5000 ;
	    RECT 1321.8000 99.3000 1325.4000 100.2000 ;
	    RECT 1326.3000 99.6000 1327.5000 100.8000 ;
	    RECT 1146.6000 99.0000 1152.6000 99.3000 ;
	    RECT 1146.6000 93.3000 1147.8000 99.0000 ;
	    RECT 1149.0000 93.3000 1150.2001 98.1000 ;
	    RECT 1151.4000 93.3000 1152.6000 99.0000 ;
	    RECT 1153.8000 93.3000 1155.0000 99.3000 ;
	    RECT 1177.8000 99.0000 1183.8000 99.3000 ;
	    RECT 1156.2001 96.4500 1157.4000 96.6000 ;
	    RECT 1168.2001 96.4500 1169.4000 96.6000 ;
	    RECT 1156.2001 95.5500 1169.4000 96.4500 ;
	    RECT 1156.2001 95.4000 1157.4000 95.5500 ;
	    RECT 1168.2001 95.4000 1169.4000 95.5500 ;
	    RECT 1177.8000 93.3000 1179.0000 99.0000 ;
	    RECT 1180.2001 93.3000 1181.4000 98.1000 ;
	    RECT 1182.6000 93.3000 1183.8000 99.0000 ;
	    RECT 1185.0000 93.3000 1186.2001 99.3000 ;
	    RECT 1209.0000 93.3000 1210.2001 99.3000 ;
	    RECT 1211.4000 99.0000 1217.4000 99.3000 ;
	    RECT 1211.4000 93.3000 1212.6000 99.0000 ;
	    RECT 1213.8000 93.3000 1215.0000 98.1000 ;
	    RECT 1216.2001 93.3000 1217.4000 99.0000 ;
	    RECT 1235.4000 93.3000 1236.6000 99.3000 ;
	    RECT 1237.8000 98.4000 1240.5000 99.3000 ;
	    RECT 1239.3000 93.3000 1240.5000 98.4000 ;
	    RECT 1242.6000 96.4500 1243.8000 96.6000 ;
	    RECT 1249.8000 96.4500 1251.0000 96.6000 ;
	    RECT 1242.6000 95.5500 1251.0000 96.4500 ;
	    RECT 1242.6000 95.4000 1243.8000 95.5500 ;
	    RECT 1249.8000 95.4000 1251.0000 95.5500 ;
	    RECT 1269.0000 93.3000 1270.2001 99.3000 ;
	    RECT 1272.9000 93.3000 1275.3000 99.3000 ;
	    RECT 1278.0000 93.3000 1279.2001 99.3000 ;
	    RECT 1321.8000 93.3000 1323.0000 99.3000 ;
	    RECT 1328.4000 98.7000 1329.3000 101.7000 ;
	    RECT 1335.0000 101.4000 1335.3000 101.7000 ;
	    RECT 1336.2001 101.4000 1337.4000 102.6000 ;
	    RECT 1330.2001 99.6000 1332.6000 100.8000 ;
	    RECT 1333.5000 100.2000 1334.7001 100.5000 ;
	    RECT 1470.3000 100.2000 1471.5000 106.8000 ;
	    RECT 1472.7001 105.9000 1473.6000 108.6000 ;
	    RECT 1508.7001 107.7000 1509.9000 108.0000 ;
	    RECT 1474.5000 106.8000 1512.9000 107.7000 ;
	    RECT 1513.8000 107.4000 1515.0000 108.6000 ;
	    RECT 1474.5000 106.5000 1475.7001 106.8000 ;
	    RECT 1472.4000 105.0000 1473.6000 105.9000 ;
	    RECT 1482.6000 105.0000 1508.1000 105.9000 ;
	    RECT 1472.4000 102.0000 1473.3000 105.0000 ;
	    RECT 1482.6000 104.1000 1483.8000 105.0000 ;
	    RECT 1509.0000 104.4000 1510.2001 105.6000 ;
	    RECT 1511.1000 105.0000 1517.7001 105.9000 ;
	    RECT 1516.5000 104.7000 1517.7001 105.0000 ;
	    RECT 1474.2001 102.9000 1479.9000 104.1000 ;
	    RECT 1472.4000 101.1000 1474.2001 102.0000 ;
	    RECT 1333.5000 99.3000 1337.4000 100.2000 ;
	    RECT 1324.2001 93.3000 1325.7001 98.4000 ;
	    RECT 1328.4000 93.3000 1330.8000 98.7000 ;
	    RECT 1333.5000 93.3000 1335.0000 98.4000 ;
	    RECT 1336.2001 93.3000 1337.4000 99.3000 ;
	    RECT 1470.3000 99.0000 1471.8000 100.2000 ;
	    RECT 1468.2001 93.3000 1469.4000 96.3000 ;
	    RECT 1470.6000 93.3000 1471.8000 99.0000 ;
	    RECT 1473.0000 93.3000 1474.2001 101.1000 ;
	    RECT 1478.7001 101.1000 1479.9000 102.9000 ;
	    RECT 1478.7001 100.2000 1481.4000 101.1000 ;
	    RECT 1480.2001 99.3000 1481.4000 100.2000 ;
	    RECT 1487.4000 99.6000 1488.6000 103.8000 ;
	    RECT 1492.2001 102.9000 1497.0000 104.1000 ;
	    RECT 1502.7001 102.9000 1505.7001 104.1000 ;
	    RECT 1518.6000 103.5000 1519.8000 111.9000 ;
	    RECT 1542.6000 107.7000 1543.8000 119.7000 ;
	    RECT 1545.0000 108.6000 1546.2001 119.7000 ;
	    RECT 1547.4000 109.5000 1548.6000 119.7000 ;
	    RECT 1549.8000 108.6000 1551.0000 119.7000 ;
	    RECT 1545.0000 107.7000 1551.0000 108.6000 ;
	    RECT 1542.9000 106.5000 1543.8000 107.7000 ;
	    RECT 1540.2001 105.4500 1541.4000 105.6000 ;
	    RECT 1542.6000 105.4500 1543.8000 105.6000 ;
	    RECT 1540.2001 104.5500 1543.8000 105.4500 ;
	    RECT 1544.7001 104.7000 1546.2001 105.6000 ;
	    RECT 1548.6000 104.7000 1548.9000 106.2000 ;
	    RECT 1540.2001 104.4000 1541.4000 104.5500 ;
	    RECT 1542.6000 104.4000 1543.8000 104.5500 ;
	    RECT 1491.6000 101.7000 1492.8000 102.0000 ;
	    RECT 1491.6000 100.8000 1498.2001 101.7000 ;
	    RECT 1499.4000 101.4000 1500.6000 102.6000 ;
	    RECT 1497.0000 100.5000 1498.2001 100.8000 ;
	    RECT 1499.4000 100.2000 1500.6000 100.5000 ;
	    RECT 1477.8000 93.3000 1479.0000 99.3000 ;
	    RECT 1480.2001 98.1000 1483.8000 99.3000 ;
	    RECT 1487.4000 98.4000 1488.9000 99.6000 ;
	    RECT 1493.4000 98.4000 1493.7001 99.6000 ;
	    RECT 1494.6000 98.4000 1495.8000 99.6000 ;
	    RECT 1497.0000 99.3000 1498.2001 99.6000 ;
	    RECT 1502.7001 99.3000 1503.9000 102.9000 ;
	    RECT 1506.6000 102.3000 1519.8000 103.5000 ;
	    RECT 1511.7001 100.2000 1516.2001 101.4000 ;
	    RECT 1511.7001 99.3000 1512.9000 100.2000 ;
	    RECT 1497.0000 98.4000 1503.9000 99.3000 ;
	    RECT 1482.6000 93.3000 1483.8000 98.1000 ;
	    RECT 1509.0000 98.1000 1512.9000 99.3000 ;
	    RECT 1485.0000 93.3000 1486.2001 97.5000 ;
	    RECT 1487.4000 93.3000 1488.6000 97.5000 ;
	    RECT 1489.8000 93.3000 1491.0000 97.5000 ;
	    RECT 1492.2001 93.3000 1493.4000 97.5000 ;
	    RECT 1494.6000 93.3000 1495.8000 96.3000 ;
	    RECT 1497.0000 93.3000 1498.2001 97.5000 ;
	    RECT 1499.4000 93.3000 1500.6000 96.3000 ;
	    RECT 1501.8000 93.3000 1503.0000 97.5000 ;
	    RECT 1504.2001 93.3000 1505.4000 97.5000 ;
	    RECT 1506.6000 93.3000 1507.8000 97.5000 ;
	    RECT 1509.0000 93.3000 1510.2001 98.1000 ;
	    RECT 1513.8000 93.3000 1515.0000 99.3000 ;
	    RECT 1518.6000 93.3000 1519.8000 102.3000 ;
	    RECT 1523.4000 99.4500 1524.6000 99.6000 ;
	    RECT 1542.6000 99.4500 1543.8000 99.6000 ;
	    RECT 1523.4000 98.5500 1543.8000 99.4500 ;
	    RECT 1545.3000 99.3000 1546.2001 104.7000 ;
	    RECT 1549.8000 104.4000 1551.0000 105.6000 ;
	    RECT 1547.4000 103.5000 1548.6000 103.8000 ;
	    RECT 1547.4000 101.4000 1548.6000 102.6000 ;
	    RECT 1523.4000 98.4000 1524.6000 98.5500 ;
	    RECT 1542.6000 98.4000 1543.8000 98.5500 ;
	    RECT 1542.9000 97.2000 1544.1000 97.5000 ;
	    RECT 1542.6000 93.3000 1543.8000 96.3000 ;
	    RECT 1545.0000 93.3000 1546.2001 99.3000 ;
	    RECT 1548.9000 93.3000 1550.1000 99.3000 ;
	    RECT 1.2000 90.6000 1569.0000 92.4000 ;
	    RECT 124.2000 80.7000 125.4000 89.7000 ;
	    RECT 129.0000 83.7000 130.2000 89.7000 ;
	    RECT 133.8000 84.9000 135.0000 89.7000 ;
	    RECT 136.2000 85.5000 137.4000 89.7000 ;
	    RECT 138.6000 85.5000 139.8000 89.7000 ;
	    RECT 141.0000 85.5000 142.2000 89.7000 ;
	    RECT 143.4000 86.7000 144.6000 89.7000 ;
	    RECT 145.8000 85.5000 147.0000 89.7000 ;
	    RECT 148.2000 86.7000 149.4000 89.7000 ;
	    RECT 150.6000 85.5000 151.8000 89.7000 ;
	    RECT 153.0000 85.5000 154.2000 89.7000 ;
	    RECT 155.4000 85.5000 156.6000 89.7000 ;
	    RECT 157.8000 85.5000 159.0000 89.7000 ;
	    RECT 131.1000 83.7000 135.0000 84.9000 ;
	    RECT 160.2000 84.9000 161.4000 89.7000 ;
	    RECT 140.1000 83.7000 147.0000 84.6000 ;
	    RECT 131.1000 82.8000 132.3000 83.7000 ;
	    RECT 127.8000 81.6000 132.3000 82.8000 ;
	    RECT 124.2000 79.5000 137.4000 80.7000 ;
	    RECT 140.1000 80.1000 141.3000 83.7000 ;
	    RECT 145.8000 83.4000 147.0000 83.7000 ;
	    RECT 148.2000 83.4000 149.4000 84.6000 ;
	    RECT 150.3000 83.4000 150.6000 84.6000 ;
	    RECT 155.1000 83.4000 156.6000 84.6000 ;
	    RECT 160.2000 83.7000 163.8000 84.9000 ;
	    RECT 165.0000 83.7000 166.2000 89.7000 ;
	    RECT 143.4000 82.5000 144.6000 82.8000 ;
	    RECT 145.8000 82.2000 147.0000 82.5000 ;
	    RECT 143.4000 80.4000 144.6000 81.6000 ;
	    RECT 145.8000 81.3000 152.4000 82.2000 ;
	    RECT 151.2000 81.0000 152.4000 81.3000 ;
	    RECT 124.2000 71.1000 125.4000 79.5000 ;
	    RECT 138.3000 78.9000 141.3000 80.1000 ;
	    RECT 147.0000 78.9000 151.8000 80.1000 ;
	    RECT 155.4000 79.2000 156.6000 83.4000 ;
	    RECT 162.6000 82.8000 163.8000 83.7000 ;
	    RECT 162.6000 81.9000 165.3000 82.8000 ;
	    RECT 164.1000 80.1000 165.3000 81.9000 ;
	    RECT 169.8000 81.9000 171.0000 89.7000 ;
	    RECT 172.2000 84.0000 173.4000 89.7000 ;
	    RECT 174.6000 86.7000 175.8000 89.7000 ;
	    RECT 309.0000 86.7000 310.2000 89.7000 ;
	    RECT 311.4000 84.0000 312.6000 89.7000 ;
	    RECT 172.2000 82.8000 173.7000 84.0000 ;
	    RECT 169.8000 81.0000 171.6000 81.9000 ;
	    RECT 164.1000 78.9000 169.8000 80.1000 ;
	    RECT 126.3000 78.0000 127.5000 78.3000 ;
	    RECT 126.3000 77.1000 132.9000 78.0000 ;
	    RECT 133.8000 77.4000 135.0000 78.6000 ;
	    RECT 160.2000 78.0000 161.4000 78.9000 ;
	    RECT 170.7000 78.0000 171.6000 81.0000 ;
	    RECT 135.9000 77.1000 161.4000 78.0000 ;
	    RECT 170.4000 77.1000 171.6000 78.0000 ;
	    RECT 168.3000 76.2000 169.5000 76.5000 ;
	    RECT 129.0000 74.4000 130.2000 75.6000 ;
	    RECT 131.1000 75.3000 169.5000 76.2000 ;
	    RECT 134.1000 75.0000 135.3000 75.3000 ;
	    RECT 170.4000 74.4000 171.3000 77.1000 ;
	    RECT 172.5000 76.2000 173.7000 82.8000 ;
	    RECT 138.6000 74.1000 139.8000 74.4000 ;
	    RECT 131.7000 73.5000 139.8000 74.1000 ;
	    RECT 130.5000 73.2000 139.8000 73.5000 ;
	    RECT 141.3000 73.5000 154.2000 74.4000 ;
	    RECT 126.6000 72.0000 129.0000 73.2000 ;
	    RECT 130.5000 72.3000 132.6000 73.2000 ;
	    RECT 141.3000 72.3000 142.2000 73.5000 ;
	    RECT 153.0000 73.2000 154.2000 73.5000 ;
	    RECT 157.8000 73.5000 171.3000 74.4000 ;
	    RECT 172.2000 75.0000 173.7000 76.2000 ;
	    RECT 311.1000 82.8000 312.6000 84.0000 ;
	    RECT 311.1000 76.2000 312.3000 82.8000 ;
	    RECT 313.8000 81.9000 315.0000 89.7000 ;
	    RECT 318.6000 83.7000 319.8000 89.7000 ;
	    RECT 323.4000 84.9000 324.6000 89.7000 ;
	    RECT 325.8000 85.5000 327.0000 89.7000 ;
	    RECT 328.2000 85.5000 329.4000 89.7000 ;
	    RECT 330.6000 85.5000 331.8000 89.7000 ;
	    RECT 333.0000 85.5000 334.2000 89.7000 ;
	    RECT 335.4000 86.7000 336.6000 89.7000 ;
	    RECT 337.8000 85.5000 339.0000 89.7000 ;
	    RECT 340.2000 86.7000 341.4000 89.7000 ;
	    RECT 342.6000 85.5000 343.8000 89.7000 ;
	    RECT 345.0000 85.5000 346.2000 89.7000 ;
	    RECT 347.4000 85.5000 348.6000 89.7000 ;
	    RECT 321.0000 83.7000 324.6000 84.9000 ;
	    RECT 349.8000 84.9000 351.0000 89.7000 ;
	    RECT 321.0000 82.8000 322.2000 83.7000 ;
	    RECT 313.2000 81.0000 315.0000 81.9000 ;
	    RECT 319.5000 81.9000 322.2000 82.8000 ;
	    RECT 328.2000 83.4000 329.7000 84.6000 ;
	    RECT 334.2000 83.4000 334.5000 84.6000 ;
	    RECT 335.4000 83.4000 336.6000 84.6000 ;
	    RECT 337.8000 83.7000 344.7000 84.6000 ;
	    RECT 349.8000 83.7000 353.7000 84.9000 ;
	    RECT 354.6000 83.7000 355.8000 89.7000 ;
	    RECT 337.8000 83.4000 339.0000 83.7000 ;
	    RECT 313.2000 78.0000 314.1000 81.0000 ;
	    RECT 319.5000 80.1000 320.7000 81.9000 ;
	    RECT 315.0000 78.9000 320.7000 80.1000 ;
	    RECT 328.2000 79.2000 329.4000 83.4000 ;
	    RECT 340.2000 82.5000 341.4000 82.8000 ;
	    RECT 337.8000 82.2000 339.0000 82.5000 ;
	    RECT 332.4000 81.3000 339.0000 82.2000 ;
	    RECT 332.4000 81.0000 333.6000 81.3000 ;
	    RECT 340.2000 80.4000 341.4000 81.6000 ;
	    RECT 343.5000 80.1000 344.7000 83.7000 ;
	    RECT 352.5000 82.8000 353.7000 83.7000 ;
	    RECT 352.5000 81.6000 357.0000 82.8000 ;
	    RECT 359.4000 80.7000 360.6000 89.7000 ;
	    RECT 491.4000 86.7000 492.6000 89.7000 ;
	    RECT 493.8000 84.0000 495.0000 89.7000 ;
	    RECT 333.0000 78.9000 337.8000 80.1000 ;
	    RECT 343.5000 78.9000 346.5000 80.1000 ;
	    RECT 347.4000 79.5000 360.6000 80.7000 ;
	    RECT 323.4000 78.0000 324.6000 78.9000 ;
	    RECT 313.2000 77.1000 314.4000 78.0000 ;
	    RECT 323.4000 77.1000 348.9000 78.0000 ;
	    RECT 349.8000 77.4000 351.0000 78.6000 ;
	    RECT 357.3000 78.0000 358.5000 78.3000 ;
	    RECT 351.9000 77.1000 358.5000 78.0000 ;
	    RECT 311.1000 75.0000 312.6000 76.2000 ;
	    RECT 172.2000 73.5000 173.4000 75.0000 ;
	    RECT 311.4000 73.5000 312.6000 75.0000 ;
	    RECT 313.5000 74.4000 314.4000 77.1000 ;
	    RECT 315.3000 76.2000 316.5000 76.5000 ;
	    RECT 315.3000 75.3000 353.7000 76.2000 ;
	    RECT 349.5000 75.0000 350.7000 75.3000 ;
	    RECT 354.6000 74.4000 355.8000 75.6000 ;
	    RECT 313.5000 73.5000 327.0000 74.4000 ;
	    RECT 157.8000 73.2000 159.0000 73.5000 ;
	    RECT 128.1000 71.4000 129.0000 72.0000 ;
	    RECT 133.5000 71.4000 142.2000 72.3000 ;
	    RECT 143.1000 71.4000 147.0000 72.6000 ;
	    RECT 124.2000 70.2000 127.2000 71.1000 ;
	    RECT 128.1000 70.2000 134.4000 71.4000 ;
	    RECT 126.3000 69.3000 127.2000 70.2000 ;
	    RECT 124.2000 63.3000 125.4000 69.3000 ;
	    RECT 126.3000 68.4000 127.8000 69.3000 ;
	    RECT 126.6000 63.3000 127.8000 68.4000 ;
	    RECT 129.0000 62.4000 130.2000 69.3000 ;
	    RECT 131.4000 63.3000 132.6000 70.2000 ;
	    RECT 133.8000 63.3000 135.0000 69.3000 ;
	    RECT 136.2000 63.3000 137.4000 67.5000 ;
	    RECT 138.6000 63.3000 139.8000 67.5000 ;
	    RECT 141.0000 63.3000 142.2000 70.5000 ;
	    RECT 143.4000 63.3000 144.6000 69.3000 ;
	    RECT 145.8000 63.3000 147.0000 70.5000 ;
	    RECT 148.2000 63.3000 149.4000 69.3000 ;
	    RECT 150.6000 63.3000 151.8000 72.6000 ;
	    RECT 162.6000 71.4000 166.5000 72.6000 ;
	    RECT 155.4000 70.2000 161.7000 71.4000 ;
	    RECT 153.0000 63.3000 154.2000 67.5000 ;
	    RECT 155.4000 63.3000 156.6000 67.5000 ;
	    RECT 157.8000 63.3000 159.0000 67.5000 ;
	    RECT 160.2000 63.3000 161.4000 69.3000 ;
	    RECT 162.6000 63.3000 163.8000 71.4000 ;
	    RECT 170.4000 71.1000 171.3000 73.5000 ;
	    RECT 172.2000 71.4000 173.4000 72.6000 ;
	    RECT 311.4000 71.4000 312.6000 72.6000 ;
	    RECT 167.4000 70.2000 171.3000 71.1000 ;
	    RECT 313.5000 71.1000 314.4000 73.5000 ;
	    RECT 325.8000 73.2000 327.0000 73.5000 ;
	    RECT 330.6000 73.5000 343.5000 74.4000 ;
	    RECT 330.6000 73.2000 331.8000 73.5000 ;
	    RECT 318.3000 71.4000 322.2000 72.6000 ;
	    RECT 165.0000 63.3000 166.2000 69.3000 ;
	    RECT 167.4000 63.3000 168.6000 70.2000 ;
	    RECT 169.8000 63.3000 171.0000 69.3000 ;
	    RECT 172.2000 63.3000 173.4000 70.5000 ;
	    RECT 174.6000 63.3000 175.8000 69.3000 ;
	    RECT 309.0000 63.3000 310.2000 69.3000 ;
	    RECT 311.4000 63.3000 312.6000 70.5000 ;
	    RECT 313.5000 70.2000 317.4000 71.1000 ;
	    RECT 313.8000 63.3000 315.0000 69.3000 ;
	    RECT 316.2000 63.3000 317.4000 70.2000 ;
	    RECT 318.6000 63.3000 319.8000 69.3000 ;
	    RECT 321.0000 63.3000 322.2000 71.4000 ;
	    RECT 323.1000 70.2000 329.4000 71.4000 ;
	    RECT 323.4000 63.3000 324.6000 69.3000 ;
	    RECT 325.8000 63.3000 327.0000 67.5000 ;
	    RECT 328.2000 63.3000 329.4000 67.5000 ;
	    RECT 330.6000 63.3000 331.8000 67.5000 ;
	    RECT 333.0000 63.3000 334.2000 72.6000 ;
	    RECT 337.8000 71.4000 341.7000 72.6000 ;
	    RECT 342.6000 72.3000 343.5000 73.5000 ;
	    RECT 345.0000 74.1000 346.2000 74.4000 ;
	    RECT 345.0000 73.5000 353.1000 74.1000 ;
	    RECT 345.0000 73.2000 354.3000 73.5000 ;
	    RECT 352.2000 72.3000 354.3000 73.2000 ;
	    RECT 342.6000 71.4000 351.3000 72.3000 ;
	    RECT 355.8000 72.0000 358.2000 73.2000 ;
	    RECT 355.8000 71.4000 356.7000 72.0000 ;
	    RECT 335.4000 63.3000 336.6000 69.3000 ;
	    RECT 337.8000 63.3000 339.0000 70.5000 ;
	    RECT 340.2000 63.3000 341.4000 69.3000 ;
	    RECT 342.6000 63.3000 343.8000 70.5000 ;
	    RECT 350.4000 70.2000 356.7000 71.4000 ;
	    RECT 359.4000 71.1000 360.6000 79.5000 ;
	    RECT 493.5000 82.8000 495.0000 84.0000 ;
	    RECT 493.5000 76.2000 494.7000 82.8000 ;
	    RECT 496.2000 81.9000 497.4000 89.7000 ;
	    RECT 501.0000 83.7000 502.2000 89.7000 ;
	    RECT 505.8000 84.9000 507.0000 89.7000 ;
	    RECT 508.2000 85.5000 509.4000 89.7000 ;
	    RECT 510.6000 85.5000 511.8000 89.7000 ;
	    RECT 513.0000 85.5000 514.2000 89.7000 ;
	    RECT 515.4000 85.5000 516.6000 89.7000 ;
	    RECT 517.8000 86.7000 519.0000 89.7000 ;
	    RECT 520.2000 85.5000 521.4000 89.7000 ;
	    RECT 522.6000 86.7000 523.8000 89.7000 ;
	    RECT 525.0000 85.5000 526.2000 89.7000 ;
	    RECT 527.4000 85.5000 528.6000 89.7000 ;
	    RECT 529.8000 85.5000 531.0000 89.7000 ;
	    RECT 503.4000 83.7000 507.0000 84.9000 ;
	    RECT 532.2000 84.9000 533.4000 89.7000 ;
	    RECT 503.4000 82.8000 504.6000 83.7000 ;
	    RECT 495.6000 81.0000 497.4000 81.9000 ;
	    RECT 501.9000 81.9000 504.6000 82.8000 ;
	    RECT 510.6000 83.4000 512.1000 84.6000 ;
	    RECT 516.6000 83.4000 516.9000 84.6000 ;
	    RECT 517.8000 83.4000 519.0000 84.6000 ;
	    RECT 520.2000 83.7000 527.1000 84.6000 ;
	    RECT 532.2000 83.7000 536.1000 84.9000 ;
	    RECT 537.0000 83.7000 538.2000 89.7000 ;
	    RECT 520.2000 83.4000 521.4000 83.7000 ;
	    RECT 495.6000 78.0000 496.5000 81.0000 ;
	    RECT 501.9000 80.1000 503.1000 81.9000 ;
	    RECT 497.4000 78.9000 503.1000 80.1000 ;
	    RECT 510.6000 79.2000 511.8000 83.4000 ;
	    RECT 522.6000 82.5000 523.8000 82.8000 ;
	    RECT 520.2000 82.2000 521.4000 82.5000 ;
	    RECT 514.8000 81.3000 521.4000 82.2000 ;
	    RECT 514.8000 81.0000 516.0000 81.3000 ;
	    RECT 522.6000 80.4000 523.8000 81.6000 ;
	    RECT 525.9000 80.1000 527.1000 83.7000 ;
	    RECT 534.9000 82.8000 536.1000 83.7000 ;
	    RECT 534.9000 81.6000 539.4000 82.8000 ;
	    RECT 541.8000 80.7000 543.0000 89.7000 ;
	    RECT 561.9000 84.6000 563.1000 89.7000 ;
	    RECT 561.9000 83.7000 564.6000 84.6000 ;
	    RECT 565.8000 83.7000 567.0000 89.7000 ;
	    RECT 515.4000 78.9000 520.2000 80.1000 ;
	    RECT 525.9000 78.9000 528.9000 80.1000 ;
	    RECT 529.8000 79.5000 543.0000 80.7000 ;
	    RECT 563.4000 79.5000 564.6000 83.7000 ;
	    RECT 565.8000 82.5000 567.0000 82.8000 ;
	    RECT 580.2000 82.5000 581.4000 89.7000 ;
	    RECT 582.6000 86.7000 583.8000 89.7000 ;
	    RECT 597.0000 86.7000 598.2000 89.7000 ;
	    RECT 582.6000 85.5000 583.8000 85.8000 ;
	    RECT 597.0000 85.5000 598.2000 85.8000 ;
	    RECT 582.6000 84.4500 583.8000 84.6000 ;
	    RECT 597.0000 84.4500 598.2000 84.6000 ;
	    RECT 582.6000 83.5500 598.2000 84.4500 ;
	    RECT 582.6000 83.4000 583.8000 83.5500 ;
	    RECT 597.0000 83.4000 598.2000 83.5500 ;
	    RECT 599.4000 82.5000 600.6000 89.7000 ;
	    RECT 717.0000 84.4500 718.2000 84.6000 ;
	    RECT 729.0000 84.4500 730.2000 84.6000 ;
	    RECT 717.0000 83.5500 730.2000 84.4500 ;
	    RECT 717.0000 83.4000 718.2000 83.5500 ;
	    RECT 729.0000 83.4000 730.2000 83.5500 ;
	    RECT 565.8000 80.4000 567.0000 81.6000 ;
	    RECT 580.2000 81.4500 581.4000 81.6000 ;
	    RECT 594.6000 81.4500 595.8000 81.6000 ;
	    RECT 580.2000 80.5500 595.8000 81.4500 ;
	    RECT 580.2000 80.4000 581.4000 80.5500 ;
	    RECT 594.6000 80.4000 595.8000 80.5500 ;
	    RECT 599.4000 81.4500 600.6000 81.6000 ;
	    RECT 729.0000 81.4500 730.2000 81.6000 ;
	    RECT 599.4000 80.5500 730.2000 81.4500 ;
	    RECT 599.4000 80.4000 600.6000 80.5500 ;
	    RECT 729.0000 80.4000 730.2000 80.5500 ;
	    RECT 731.4000 80.7000 732.6000 89.7000 ;
	    RECT 736.2000 83.7000 737.4000 89.7000 ;
	    RECT 741.0000 84.9000 742.2000 89.7000 ;
	    RECT 743.4000 85.5000 744.6000 89.7000 ;
	    RECT 745.8000 85.5000 747.0000 89.7000 ;
	    RECT 748.2000 85.5000 749.4000 89.7000 ;
	    RECT 750.6000 86.7000 751.8000 89.7000 ;
	    RECT 753.0000 85.5000 754.2000 89.7000 ;
	    RECT 755.4000 86.7000 756.6000 89.7000 ;
	    RECT 757.8000 85.5000 759.0000 89.7000 ;
	    RECT 760.2000 85.5000 761.4000 89.7000 ;
	    RECT 762.6000 85.5000 763.8000 89.7000 ;
	    RECT 765.0000 85.5000 766.2000 89.7000 ;
	    RECT 738.3000 83.7000 742.2000 84.9000 ;
	    RECT 767.4000 84.9000 768.6000 89.7000 ;
	    RECT 747.3000 83.7000 754.2000 84.6000 ;
	    RECT 738.3000 82.8000 739.5000 83.7000 ;
	    RECT 735.0000 81.6000 739.5000 82.8000 ;
	    RECT 731.4000 79.5000 744.6000 80.7000 ;
	    RECT 747.3000 80.1000 748.5000 83.7000 ;
	    RECT 753.0000 83.4000 754.2000 83.7000 ;
	    RECT 755.4000 83.4000 756.6000 84.6000 ;
	    RECT 757.5000 83.4000 757.8000 84.6000 ;
	    RECT 762.3000 83.4000 763.8000 84.6000 ;
	    RECT 767.4000 83.7000 771.0000 84.9000 ;
	    RECT 772.2000 83.7000 773.4000 89.7000 ;
	    RECT 750.6000 82.5000 751.8000 82.8000 ;
	    RECT 753.0000 82.2000 754.2000 82.5000 ;
	    RECT 750.6000 80.4000 751.8000 81.6000 ;
	    RECT 753.0000 81.3000 759.6000 82.2000 ;
	    RECT 758.4000 81.0000 759.6000 81.3000 ;
	    RECT 505.8000 78.0000 507.0000 78.9000 ;
	    RECT 495.6000 77.1000 496.8000 78.0000 ;
	    RECT 505.8000 77.1000 531.3000 78.0000 ;
	    RECT 532.2000 77.4000 533.4000 78.6000 ;
	    RECT 539.7000 78.0000 540.9000 78.3000 ;
	    RECT 534.3000 77.1000 540.9000 78.0000 ;
	    RECT 493.5000 75.0000 495.0000 76.2000 ;
	    RECT 493.8000 73.5000 495.0000 75.0000 ;
	    RECT 495.9000 74.4000 496.8000 77.1000 ;
	    RECT 497.7000 76.2000 498.9000 76.5000 ;
	    RECT 497.7000 75.3000 536.1000 76.2000 ;
	    RECT 531.9000 75.0000 533.1000 75.3000 ;
	    RECT 537.0000 74.4000 538.2000 75.6000 ;
	    RECT 495.9000 73.5000 509.4000 74.4000 ;
	    RECT 493.8000 71.4000 495.0000 72.6000 ;
	    RECT 357.6000 70.2000 360.6000 71.1000 ;
	    RECT 495.9000 71.1000 496.8000 73.5000 ;
	    RECT 508.2000 73.2000 509.4000 73.5000 ;
	    RECT 513.0000 73.5000 525.9000 74.4000 ;
	    RECT 513.0000 73.2000 514.2000 73.5000 ;
	    RECT 500.7000 71.4000 504.6000 72.6000 ;
	    RECT 345.0000 63.3000 346.2000 67.5000 ;
	    RECT 347.4000 63.3000 348.6000 67.5000 ;
	    RECT 349.8000 63.3000 351.0000 69.3000 ;
	    RECT 352.2000 63.3000 353.4000 70.2000 ;
	    RECT 357.6000 69.3000 358.5000 70.2000 ;
	    RECT 354.6000 62.4000 355.8000 69.3000 ;
	    RECT 357.0000 68.4000 358.5000 69.3000 ;
	    RECT 357.0000 63.3000 358.2000 68.4000 ;
	    RECT 359.4000 63.3000 360.6000 69.3000 ;
	    RECT 491.4000 63.3000 492.6000 69.3000 ;
	    RECT 493.8000 63.3000 495.0000 70.5000 ;
	    RECT 495.9000 70.2000 499.8000 71.1000 ;
	    RECT 496.2000 63.3000 497.4000 69.3000 ;
	    RECT 498.6000 63.3000 499.8000 70.2000 ;
	    RECT 501.0000 63.3000 502.2000 69.3000 ;
	    RECT 503.4000 63.3000 504.6000 71.4000 ;
	    RECT 505.5000 70.2000 511.8000 71.4000 ;
	    RECT 505.8000 63.3000 507.0000 69.3000 ;
	    RECT 508.2000 63.3000 509.4000 67.5000 ;
	    RECT 510.6000 63.3000 511.8000 67.5000 ;
	    RECT 513.0000 63.3000 514.2000 67.5000 ;
	    RECT 515.4000 63.3000 516.6000 72.6000 ;
	    RECT 520.2000 71.4000 524.1000 72.6000 ;
	    RECT 525.0000 72.3000 525.9000 73.5000 ;
	    RECT 527.4000 74.1000 528.6000 74.4000 ;
	    RECT 527.4000 73.5000 535.5000 74.1000 ;
	    RECT 527.4000 73.2000 536.7000 73.5000 ;
	    RECT 534.6000 72.3000 536.7000 73.2000 ;
	    RECT 525.0000 71.4000 533.7000 72.3000 ;
	    RECT 538.2000 72.0000 540.6000 73.2000 ;
	    RECT 538.2000 71.4000 539.1000 72.0000 ;
	    RECT 517.8000 63.3000 519.0000 69.3000 ;
	    RECT 520.2000 63.3000 521.4000 70.5000 ;
	    RECT 522.6000 63.3000 523.8000 69.3000 ;
	    RECT 525.0000 63.3000 526.2000 70.5000 ;
	    RECT 532.8000 70.2000 539.1000 71.4000 ;
	    RECT 541.8000 71.1000 543.0000 79.5000 ;
	    RECT 563.4000 78.4500 564.6000 78.6000 ;
	    RECT 573.0000 78.4500 574.2000 78.6000 ;
	    RECT 563.4000 77.5500 574.2000 78.4500 ;
	    RECT 563.4000 77.4000 564.6000 77.5500 ;
	    RECT 573.0000 77.4000 574.2000 77.5500 ;
	    RECT 544.2000 75.4500 545.4000 75.6000 ;
	    RECT 561.0000 75.4500 562.2000 75.6000 ;
	    RECT 544.2000 74.5500 562.2000 75.4500 ;
	    RECT 544.2000 74.4000 545.4000 74.5500 ;
	    RECT 561.0000 74.4000 562.2000 74.5500 ;
	    RECT 561.0000 73.2000 562.2000 73.5000 ;
	    RECT 540.0000 70.2000 543.0000 71.1000 ;
	    RECT 527.4000 63.3000 528.6000 67.5000 ;
	    RECT 529.8000 63.3000 531.0000 67.5000 ;
	    RECT 532.2000 63.3000 533.4000 69.3000 ;
	    RECT 534.6000 63.3000 535.8000 70.2000 ;
	    RECT 540.0000 69.3000 540.9000 70.2000 ;
	    RECT 537.0000 62.4000 538.2000 69.3000 ;
	    RECT 539.4000 68.4000 540.9000 69.3000 ;
	    RECT 539.4000 63.3000 540.6000 68.4000 ;
	    RECT 541.8000 63.3000 543.0000 69.3000 ;
	    RECT 561.0000 63.3000 562.2000 69.3000 ;
	    RECT 563.4000 63.3000 564.6000 76.5000 ;
	    RECT 565.8000 63.3000 567.0000 69.3000 ;
	    RECT 580.2000 63.3000 581.4000 79.5000 ;
	    RECT 582.6000 63.3000 583.8000 69.3000 ;
	    RECT 597.0000 63.3000 598.2000 69.3000 ;
	    RECT 599.4000 63.3000 600.6000 79.5000 ;
	    RECT 731.4000 71.1000 732.6000 79.5000 ;
	    RECT 745.5000 78.9000 748.5000 80.1000 ;
	    RECT 754.2000 78.9000 759.0000 80.1000 ;
	    RECT 762.6000 79.2000 763.8000 83.4000 ;
	    RECT 769.8000 82.8000 771.0000 83.7000 ;
	    RECT 769.8000 81.9000 772.5000 82.8000 ;
	    RECT 771.3000 80.1000 772.5000 81.9000 ;
	    RECT 777.0000 81.9000 778.2000 89.7000 ;
	    RECT 779.4000 84.0000 780.6000 89.7000 ;
	    RECT 781.8000 86.7000 783.0000 89.7000 ;
	    RECT 779.4000 82.8000 780.9000 84.0000 ;
	    RECT 832.2000 83.7000 833.4000 89.7000 ;
	    RECT 834.6000 82.8000 835.8000 89.7000 ;
	    RECT 837.0000 83.7000 838.2000 89.7000 ;
	    RECT 839.4000 82.8000 840.6000 89.7000 ;
	    RECT 841.8000 83.7000 843.0000 89.7000 ;
	    RECT 844.2000 82.8000 845.4000 89.7000 ;
	    RECT 846.6000 83.7000 847.8000 89.7000 ;
	    RECT 849.0000 82.8000 850.2000 89.7000 ;
	    RECT 851.4000 83.7000 852.6000 89.7000 ;
	    RECT 911.4000 83.7000 912.6000 89.7000 ;
	    RECT 777.0000 81.0000 778.8000 81.9000 ;
	    RECT 771.3000 78.9000 777.0000 80.1000 ;
	    RECT 733.5000 78.0000 734.7000 78.3000 ;
	    RECT 733.5000 77.1000 740.1000 78.0000 ;
	    RECT 741.0000 77.4000 742.2000 78.6000 ;
	    RECT 767.4000 78.0000 768.6000 78.9000 ;
	    RECT 777.9000 78.0000 778.8000 81.0000 ;
	    RECT 743.1000 77.1000 768.6000 78.0000 ;
	    RECT 777.6000 77.1000 778.8000 78.0000 ;
	    RECT 775.5000 76.2000 776.7000 76.5000 ;
	    RECT 736.2000 74.4000 737.4000 75.6000 ;
	    RECT 738.3000 75.3000 776.7000 76.2000 ;
	    RECT 741.3000 75.0000 742.5000 75.3000 ;
	    RECT 777.6000 74.4000 778.5000 77.1000 ;
	    RECT 779.7000 76.2000 780.9000 82.8000 ;
	    RECT 832.2000 81.6000 835.8000 82.8000 ;
	    RECT 837.3000 81.6000 840.6000 82.8000 ;
	    RECT 842.1000 81.6000 845.4000 82.8000 ;
	    RECT 847.5000 81.6000 850.2000 82.8000 ;
	    RECT 913.8000 82.8000 915.0000 89.7000 ;
	    RECT 916.2000 83.7000 917.4000 89.7000 ;
	    RECT 918.6000 82.8000 919.8000 89.7000 ;
	    RECT 921.0000 83.7000 922.2000 89.7000 ;
	    RECT 923.4000 82.8000 924.6000 89.7000 ;
	    RECT 925.8000 83.7000 927.0000 89.7000 ;
	    RECT 928.2000 82.8000 929.4000 89.7000 ;
	    RECT 930.6000 83.7000 931.8000 89.7000 ;
	    RECT 950.7000 84.6000 951.9000 89.7000 ;
	    RECT 950.7000 83.7000 953.4000 84.6000 ;
	    RECT 954.6000 83.7000 955.8000 89.7000 ;
	    RECT 973.8000 83.7000 975.0000 89.7000 ;
	    RECT 977.7000 84.6000 978.9000 89.7000 ;
	    RECT 990.6000 86.7000 991.8000 89.7000 ;
	    RECT 990.6000 85.5000 991.8000 85.8000 ;
	    RECT 976.2000 83.7000 978.9000 84.6000 ;
	    RECT 913.8000 81.6000 916.5000 82.8000 ;
	    RECT 918.6000 81.6000 921.9000 82.8000 ;
	    RECT 923.4000 81.6000 926.7000 82.8000 ;
	    RECT 928.2000 81.6000 931.8000 82.8000 ;
	    RECT 832.2000 79.5000 833.4000 81.6000 ;
	    RECT 837.3000 80.7000 838.5000 81.6000 ;
	    RECT 842.1000 80.7000 843.3000 81.6000 ;
	    RECT 847.5000 80.7000 848.7000 81.6000 ;
	    RECT 851.4000 81.4500 852.6000 81.6000 ;
	    RECT 911.4000 81.4500 912.6000 81.6000 ;
	    RECT 834.6000 79.5000 838.5000 80.7000 ;
	    RECT 839.7000 79.5000 843.3000 80.7000 ;
	    RECT 844.8000 79.5000 848.7000 80.7000 ;
	    RECT 849.9000 79.5000 850.5000 80.7000 ;
	    RECT 851.4000 80.5500 912.6000 81.4500 ;
	    RECT 915.3000 80.7000 916.5000 81.6000 ;
	    RECT 920.7000 80.7000 921.9000 81.6000 ;
	    RECT 925.5000 80.7000 926.7000 81.6000 ;
	    RECT 851.4000 80.4000 852.6000 80.5500 ;
	    RECT 911.4000 80.4000 912.6000 80.5500 ;
	    RECT 913.5000 79.5000 914.1000 80.7000 ;
	    RECT 915.3000 79.5000 919.2000 80.7000 ;
	    RECT 920.7000 79.5000 924.3000 80.7000 ;
	    RECT 925.5000 79.5000 929.4000 80.7000 ;
	    RECT 930.6000 79.5000 931.8000 81.6000 ;
	    RECT 952.2000 79.5000 953.4000 83.7000 ;
	    RECT 954.6000 82.5000 955.8000 82.8000 ;
	    RECT 973.8000 82.5000 975.0000 82.8000 ;
	    RECT 954.6000 81.4500 955.8000 81.6000 ;
	    RECT 971.4000 81.4500 972.6000 81.6000 ;
	    RECT 954.6000 80.5500 972.6000 81.4500 ;
	    RECT 954.6000 80.4000 955.8000 80.5500 ;
	    RECT 971.4000 80.4000 972.6000 80.5500 ;
	    RECT 973.8000 80.4000 975.0000 81.6000 ;
	    RECT 976.2000 79.5000 977.4000 83.7000 ;
	    RECT 990.6000 83.4000 991.8000 84.6000 ;
	    RECT 993.0000 82.5000 994.2000 89.7000 ;
	    RECT 1127.4000 86.7000 1128.6000 89.7000 ;
	    RECT 1129.8000 84.0000 1131.0000 89.7000 ;
	    RECT 1129.5000 82.8000 1131.0000 84.0000 ;
	    RECT 993.0000 81.4500 994.2000 81.6000 ;
	    RECT 997.8000 81.4500 999.0000 81.6000 ;
	    RECT 993.0000 80.5500 999.0000 81.4500 ;
	    RECT 993.0000 80.4000 994.2000 80.5500 ;
	    RECT 997.8000 80.4000 999.0000 80.5500 ;
	    RECT 808.2000 78.4500 809.4000 78.6000 ;
	    RECT 832.2000 78.4500 833.4000 78.6000 ;
	    RECT 808.2000 77.5500 833.4000 78.4500 ;
	    RECT 808.2000 77.4000 809.4000 77.5500 ;
	    RECT 832.2000 77.4000 833.4000 77.5500 ;
	    RECT 837.3000 77.4000 838.5000 79.5000 ;
	    RECT 842.1000 77.4000 843.3000 79.5000 ;
	    RECT 847.5000 77.4000 848.7000 79.5000 ;
	    RECT 915.3000 77.4000 916.5000 79.5000 ;
	    RECT 920.7000 77.4000 921.9000 79.5000 ;
	    RECT 925.5000 77.4000 926.7000 79.5000 ;
	    RECT 930.6000 78.4500 931.8000 78.6000 ;
	    RECT 942.6000 78.4500 943.8000 78.6000 ;
	    RECT 947.4000 78.4500 948.6000 78.6000 ;
	    RECT 930.6000 77.5500 948.6000 78.4500 ;
	    RECT 930.6000 77.4000 931.8000 77.5500 ;
	    RECT 942.6000 77.4000 943.8000 77.5500 ;
	    RECT 947.4000 77.4000 948.6000 77.5500 ;
	    RECT 952.2000 78.4500 953.4000 78.6000 ;
	    RECT 964.2000 78.4500 965.4000 78.6000 ;
	    RECT 952.2000 77.5500 965.4000 78.4500 ;
	    RECT 952.2000 77.4000 953.4000 77.5500 ;
	    RECT 964.2000 77.4000 965.4000 77.5500 ;
	    RECT 976.2000 78.4500 977.4000 78.6000 ;
	    RECT 990.6000 78.4500 991.8000 78.6000 ;
	    RECT 976.2000 77.5500 991.8000 78.4500 ;
	    RECT 976.2000 77.4000 977.4000 77.5500 ;
	    RECT 990.6000 77.4000 991.8000 77.5500 ;
	    RECT 834.3000 76.5000 835.8000 77.4000 ;
	    RECT 832.2000 76.2000 835.8000 76.5000 ;
	    RECT 837.3000 76.2000 840.6000 77.4000 ;
	    RECT 842.1000 76.2000 845.4000 77.4000 ;
	    RECT 847.5000 76.2000 850.2000 77.4000 ;
	    RECT 745.8000 74.1000 747.0000 74.4000 ;
	    RECT 738.9000 73.5000 747.0000 74.1000 ;
	    RECT 737.7000 73.2000 747.0000 73.5000 ;
	    RECT 748.5000 73.5000 761.4000 74.4000 ;
	    RECT 733.8000 72.0000 736.2000 73.2000 ;
	    RECT 737.7000 72.3000 739.8000 73.2000 ;
	    RECT 748.5000 72.3000 749.4000 73.5000 ;
	    RECT 760.2000 73.2000 761.4000 73.5000 ;
	    RECT 765.0000 73.5000 778.5000 74.4000 ;
	    RECT 779.4000 75.0000 780.9000 76.2000 ;
	    RECT 779.4000 73.5000 780.6000 75.0000 ;
	    RECT 765.0000 73.2000 766.2000 73.5000 ;
	    RECT 735.3000 71.4000 736.2000 72.0000 ;
	    RECT 740.7000 71.4000 749.4000 72.3000 ;
	    RECT 750.3000 71.4000 754.2000 72.6000 ;
	    RECT 731.4000 70.2000 734.4000 71.1000 ;
	    RECT 735.3000 70.2000 741.6000 71.4000 ;
	    RECT 733.5000 69.3000 734.4000 70.2000 ;
	    RECT 731.4000 63.3000 732.6000 69.3000 ;
	    RECT 733.5000 68.4000 735.0000 69.3000 ;
	    RECT 733.8000 63.3000 735.0000 68.4000 ;
	    RECT 736.2000 62.4000 737.4000 69.3000 ;
	    RECT 738.6000 63.3000 739.8000 70.2000 ;
	    RECT 741.0000 63.3000 742.2000 69.3000 ;
	    RECT 743.4000 63.3000 744.6000 67.5000 ;
	    RECT 745.8000 63.3000 747.0000 67.5000 ;
	    RECT 748.2000 63.3000 749.4000 70.5000 ;
	    RECT 750.6000 63.3000 751.8000 69.3000 ;
	    RECT 753.0000 63.3000 754.2000 70.5000 ;
	    RECT 755.4000 63.3000 756.6000 69.3000 ;
	    RECT 757.8000 63.3000 759.0000 72.6000 ;
	    RECT 769.8000 71.4000 773.7000 72.6000 ;
	    RECT 762.6000 70.2000 768.9000 71.4000 ;
	    RECT 760.2000 63.3000 761.4000 67.5000 ;
	    RECT 762.6000 63.3000 763.8000 67.5000 ;
	    RECT 765.0000 63.3000 766.2000 67.5000 ;
	    RECT 767.4000 63.3000 768.6000 69.3000 ;
	    RECT 769.8000 63.3000 771.0000 71.4000 ;
	    RECT 777.6000 71.1000 778.5000 73.5000 ;
	    RECT 779.4000 71.4000 780.6000 72.6000 ;
	    RECT 774.6000 70.2000 778.5000 71.1000 ;
	    RECT 772.2000 63.3000 773.4000 69.3000 ;
	    RECT 774.6000 63.3000 775.8000 70.2000 ;
	    RECT 777.0000 63.3000 778.2000 69.3000 ;
	    RECT 779.4000 63.3000 780.6000 70.5000 ;
	    RECT 781.8000 63.3000 783.0000 69.3000 ;
	    RECT 832.2000 63.3000 833.4000 75.3000 ;
	    RECT 834.6000 63.3000 835.8000 76.2000 ;
	    RECT 837.0000 63.3000 838.2000 75.3000 ;
	    RECT 839.4000 63.3000 840.6000 76.2000 ;
	    RECT 841.8000 63.3000 843.0000 75.3000 ;
	    RECT 844.2000 63.3000 845.4000 76.2000 ;
	    RECT 846.6000 63.3000 847.8000 75.3000 ;
	    RECT 849.0000 63.3000 850.2000 76.2000 ;
	    RECT 913.8000 76.2000 916.5000 77.4000 ;
	    RECT 918.6000 76.2000 921.9000 77.4000 ;
	    RECT 923.4000 76.2000 926.7000 77.4000 ;
	    RECT 928.2000 76.5000 929.7000 77.4000 ;
	    RECT 928.2000 76.2000 931.8000 76.5000 ;
	    RECT 851.4000 63.3000 852.6000 75.3000 ;
	    RECT 911.4000 63.3000 912.6000 75.3000 ;
	    RECT 913.8000 63.3000 915.0000 76.2000 ;
	    RECT 916.2000 63.3000 917.4000 75.3000 ;
	    RECT 918.6000 63.3000 919.8000 76.2000 ;
	    RECT 921.0000 63.3000 922.2000 75.3000 ;
	    RECT 923.4000 63.3000 924.6000 76.2000 ;
	    RECT 925.8000 63.3000 927.0000 75.3000 ;
	    RECT 928.2000 63.3000 929.4000 76.2000 ;
	    RECT 935.4000 75.4500 936.6000 75.6000 ;
	    RECT 949.8000 75.4500 951.0000 75.6000 ;
	    RECT 930.6000 63.3000 931.8000 75.3000 ;
	    RECT 935.4000 74.5500 951.0000 75.4500 ;
	    RECT 935.4000 74.4000 936.6000 74.5500 ;
	    RECT 949.8000 74.4000 951.0000 74.5500 ;
	    RECT 949.8000 73.2000 951.0000 73.5000 ;
	    RECT 949.8000 63.3000 951.0000 69.3000 ;
	    RECT 952.2000 63.3000 953.4000 76.5000 ;
	    RECT 954.6000 63.3000 955.8000 69.3000 ;
	    RECT 973.8000 63.3000 975.0000 69.3000 ;
	    RECT 976.2000 63.3000 977.4000 76.5000 ;
	    RECT 978.6000 74.4000 979.8000 75.6000 ;
	    RECT 978.6000 73.2000 979.8000 73.5000 ;
	    RECT 978.6000 63.3000 979.8000 69.3000 ;
	    RECT 990.6000 63.3000 991.8000 69.3000 ;
	    RECT 993.0000 63.3000 994.2000 79.5000 ;
	    RECT 1129.5000 76.2000 1130.7001 82.8000 ;
	    RECT 1132.2001 81.9000 1133.4000 89.7000 ;
	    RECT 1137.0000 83.7000 1138.2001 89.7000 ;
	    RECT 1141.8000 84.9000 1143.0000 89.7000 ;
	    RECT 1144.2001 85.5000 1145.4000 89.7000 ;
	    RECT 1146.6000 85.5000 1147.8000 89.7000 ;
	    RECT 1149.0000 85.5000 1150.2001 89.7000 ;
	    RECT 1151.4000 85.5000 1152.6000 89.7000 ;
	    RECT 1153.8000 86.7000 1155.0000 89.7000 ;
	    RECT 1156.2001 85.5000 1157.4000 89.7000 ;
	    RECT 1158.6000 86.7000 1159.8000 89.7000 ;
	    RECT 1161.0000 85.5000 1162.2001 89.7000 ;
	    RECT 1163.4000 85.5000 1164.6000 89.7000 ;
	    RECT 1165.8000 85.5000 1167.0000 89.7000 ;
	    RECT 1139.4000 83.7000 1143.0000 84.9000 ;
	    RECT 1168.2001 84.9000 1169.4000 89.7000 ;
	    RECT 1139.4000 82.8000 1140.6000 83.7000 ;
	    RECT 1131.6000 81.0000 1133.4000 81.9000 ;
	    RECT 1137.9000 81.9000 1140.6000 82.8000 ;
	    RECT 1146.6000 83.4000 1148.1000 84.6000 ;
	    RECT 1152.6000 83.4000 1152.9000 84.6000 ;
	    RECT 1153.8000 83.4000 1155.0000 84.6000 ;
	    RECT 1156.2001 83.7000 1163.1000 84.6000 ;
	    RECT 1168.2001 83.7000 1172.1000 84.9000 ;
	    RECT 1173.0000 83.7000 1174.2001 89.7000 ;
	    RECT 1156.2001 83.4000 1157.4000 83.7000 ;
	    RECT 1131.6000 78.0000 1132.5000 81.0000 ;
	    RECT 1137.9000 80.1000 1139.1000 81.9000 ;
	    RECT 1133.4000 78.9000 1139.1000 80.1000 ;
	    RECT 1146.6000 79.2000 1147.8000 83.4000 ;
	    RECT 1158.6000 82.5000 1159.8000 82.8000 ;
	    RECT 1156.2001 82.2000 1157.4000 82.5000 ;
	    RECT 1150.8000 81.3000 1157.4000 82.2000 ;
	    RECT 1150.8000 81.0000 1152.0000 81.3000 ;
	    RECT 1158.6000 80.4000 1159.8000 81.6000 ;
	    RECT 1161.9000 80.1000 1163.1000 83.7000 ;
	    RECT 1170.9000 82.8000 1172.1000 83.7000 ;
	    RECT 1170.9000 81.6000 1175.4000 82.8000 ;
	    RECT 1177.8000 80.7000 1179.0000 89.7000 ;
	    RECT 1204.2001 84.0000 1205.4000 89.7000 ;
	    RECT 1206.6000 84.9000 1207.8000 89.7000 ;
	    RECT 1209.0000 84.0000 1210.2001 89.7000 ;
	    RECT 1204.2001 83.7000 1210.2001 84.0000 ;
	    RECT 1211.4000 83.7000 1212.6000 89.7000 ;
	    RECT 1240.8000 83.7000 1242.0000 89.7000 ;
	    RECT 1244.7001 83.7000 1247.1000 89.7000 ;
	    RECT 1249.8000 83.7000 1251.0000 89.7000 ;
	    RECT 1276.2001 83.7000 1277.4000 89.7000 ;
	    RECT 1278.6000 84.0000 1279.8000 89.7000 ;
	    RECT 1281.0000 84.9000 1282.2001 89.7000 ;
	    RECT 1283.4000 84.0000 1284.6000 89.7000 ;
	    RECT 1278.6000 83.7000 1284.6000 84.0000 ;
	    RECT 1303.5000 84.6000 1304.7001 89.7000 ;
	    RECT 1303.5000 83.7000 1306.2001 84.6000 ;
	    RECT 1307.4000 83.7000 1308.6000 89.7000 ;
	    RECT 1326.6000 83.7000 1327.8000 89.7000 ;
	    RECT 1330.5000 84.6000 1331.7001 89.7000 ;
	    RECT 1329.0000 83.7000 1331.7001 84.6000 ;
	    RECT 1362.6000 83.7000 1363.8000 89.7000 ;
	    RECT 1365.0000 84.0000 1366.2001 89.7000 ;
	    RECT 1367.4000 84.9000 1368.6000 89.7000 ;
	    RECT 1369.8000 84.0000 1371.0000 89.7000 ;
	    RECT 1365.0000 83.7000 1371.0000 84.0000 ;
	    RECT 1204.5000 83.1000 1209.9000 83.7000 ;
	    RECT 1211.4000 82.5000 1212.3000 83.7000 ;
	    RECT 1151.4000 78.9000 1156.2001 80.1000 ;
	    RECT 1161.9000 78.9000 1164.9000 80.1000 ;
	    RECT 1165.8000 79.5000 1179.0000 80.7000 ;
	    RECT 1180.2001 81.4500 1181.4000 81.6000 ;
	    RECT 1204.2001 81.4500 1205.4000 81.6000 ;
	    RECT 1180.2001 80.5500 1205.4000 81.4500 ;
	    RECT 1206.3000 80.7000 1206.6000 82.2000 ;
	    RECT 1180.2001 80.4000 1181.4000 80.5500 ;
	    RECT 1204.2001 80.4000 1205.4000 80.5500 ;
	    RECT 1208.7001 80.4000 1210.5000 81.6000 ;
	    RECT 1211.4000 81.4500 1212.6000 81.6000 ;
	    RECT 1237.8000 81.4500 1239.0000 81.6000 ;
	    RECT 1211.4000 80.5500 1239.0000 81.4500 ;
	    RECT 1211.4000 80.4000 1212.6000 80.5500 ;
	    RECT 1237.8000 80.4000 1239.0000 80.5500 ;
	    RECT 1242.6000 80.4000 1243.8000 81.6000 ;
	    RECT 1206.6000 79.5000 1207.8000 79.8000 ;
	    RECT 1141.8000 78.0000 1143.0000 78.9000 ;
	    RECT 1131.6000 77.1000 1132.8000 78.0000 ;
	    RECT 1141.8000 77.1000 1167.3000 78.0000 ;
	    RECT 1168.2001 77.4000 1169.4000 78.6000 ;
	    RECT 1175.7001 78.0000 1176.9000 78.3000 ;
	    RECT 1170.3000 77.1000 1176.9000 78.0000 ;
	    RECT 1129.5000 75.0000 1131.0000 76.2000 ;
	    RECT 1129.8000 73.5000 1131.0000 75.0000 ;
	    RECT 1131.9000 74.4000 1132.8000 77.1000 ;
	    RECT 1133.7001 76.2000 1134.9000 76.5000 ;
	    RECT 1133.7001 75.3000 1172.1000 76.2000 ;
	    RECT 1167.9000 75.0000 1169.1000 75.3000 ;
	    RECT 1173.0000 74.4000 1174.2001 75.6000 ;
	    RECT 1131.9000 73.5000 1145.4000 74.4000 ;
	    RECT 1089.0000 72.4500 1090.2001 72.6000 ;
	    RECT 1113.0000 72.4500 1114.2001 72.6000 ;
	    RECT 1129.8000 72.4500 1131.0000 72.6000 ;
	    RECT 1089.0000 71.5500 1131.0000 72.4500 ;
	    RECT 1089.0000 71.4000 1090.2001 71.5500 ;
	    RECT 1113.0000 71.4000 1114.2001 71.5500 ;
	    RECT 1129.8000 71.4000 1131.0000 71.5500 ;
	    RECT 1131.9000 71.1000 1132.8000 73.5000 ;
	    RECT 1144.2001 73.2000 1145.4000 73.5000 ;
	    RECT 1149.0000 73.5000 1161.9000 74.4000 ;
	    RECT 1149.0000 73.2000 1150.2001 73.5000 ;
	    RECT 1136.7001 71.4000 1140.6000 72.6000 ;
	    RECT 1127.4000 63.3000 1128.6000 69.3000 ;
	    RECT 1129.8000 63.3000 1131.0000 70.5000 ;
	    RECT 1131.9000 70.2000 1135.8000 71.1000 ;
	    RECT 1132.2001 63.3000 1133.4000 69.3000 ;
	    RECT 1134.6000 63.3000 1135.8000 70.2000 ;
	    RECT 1137.0000 63.3000 1138.2001 69.3000 ;
	    RECT 1139.4000 63.3000 1140.6000 71.4000 ;
	    RECT 1141.5000 70.2000 1147.8000 71.4000 ;
	    RECT 1141.8000 63.3000 1143.0000 69.3000 ;
	    RECT 1144.2001 63.3000 1145.4000 67.5000 ;
	    RECT 1146.6000 63.3000 1147.8000 67.5000 ;
	    RECT 1149.0000 63.3000 1150.2001 67.5000 ;
	    RECT 1151.4000 63.3000 1152.6000 72.6000 ;
	    RECT 1156.2001 71.4000 1160.1000 72.6000 ;
	    RECT 1161.0000 72.3000 1161.9000 73.5000 ;
	    RECT 1163.4000 74.1000 1164.6000 74.4000 ;
	    RECT 1163.4000 73.5000 1171.5000 74.1000 ;
	    RECT 1163.4000 73.2000 1172.7001 73.5000 ;
	    RECT 1170.6000 72.3000 1172.7001 73.2000 ;
	    RECT 1161.0000 71.4000 1169.7001 72.3000 ;
	    RECT 1174.2001 72.0000 1176.6000 73.2000 ;
	    RECT 1174.2001 71.4000 1175.1000 72.0000 ;
	    RECT 1153.8000 63.3000 1155.0000 69.3000 ;
	    RECT 1156.2001 63.3000 1157.4000 70.5000 ;
	    RECT 1158.6000 63.3000 1159.8000 69.3000 ;
	    RECT 1161.0000 63.3000 1162.2001 70.5000 ;
	    RECT 1168.8000 70.2000 1175.1000 71.4000 ;
	    RECT 1177.8000 71.1000 1179.0000 79.5000 ;
	    RECT 1185.0000 78.4500 1186.2001 78.6000 ;
	    RECT 1206.6000 78.4500 1207.8000 78.6000 ;
	    RECT 1185.0000 77.5500 1207.8000 78.4500 ;
	    RECT 1185.0000 77.4000 1186.2001 77.5500 ;
	    RECT 1206.6000 77.4000 1207.8000 77.5500 ;
	    RECT 1208.7001 75.3000 1209.6000 80.4000 ;
	    RECT 1245.3000 79.5000 1246.2001 83.7000 ;
	    RECT 1276.5000 82.5000 1277.4000 83.7000 ;
	    RECT 1278.9000 83.1000 1284.3000 83.7000 ;
	    RECT 1247.4000 80.4000 1248.6000 81.6000 ;
	    RECT 1249.8000 81.4500 1251.0000 81.6000 ;
	    RECT 1276.2001 81.4500 1277.4000 81.6000 ;
	    RECT 1249.8000 80.5500 1277.4000 81.4500 ;
	    RECT 1249.8000 80.4000 1251.0000 80.5500 ;
	    RECT 1276.2001 80.4000 1277.4000 80.5500 ;
	    RECT 1278.3000 80.4000 1280.1000 81.6000 ;
	    RECT 1282.2001 80.7000 1282.5000 82.2000 ;
	    RECT 1283.4000 81.4500 1284.6000 81.6000 ;
	    RECT 1288.2001 81.4500 1289.4000 81.6000 ;
	    RECT 1283.4000 80.5500 1289.4000 81.4500 ;
	    RECT 1283.4000 80.4000 1284.6000 80.5500 ;
	    RECT 1288.2001 80.4000 1289.4000 80.5500 ;
	    RECT 1242.6000 79.2000 1243.8000 79.5000 ;
	    RECT 1247.1000 78.6000 1248.3000 79.5000 ;
	    RECT 1223.4000 78.4500 1224.6000 78.6000 ;
	    RECT 1240.2001 78.4500 1241.4000 78.6000 ;
	    RECT 1211.5500 77.5500 1241.4000 78.4500 ;
	    RECT 1211.5500 75.6000 1212.4501 77.5500 ;
	    RECT 1223.4000 77.4000 1224.6000 77.5500 ;
	    RECT 1240.2001 77.4000 1241.4000 77.5500 ;
	    RECT 1242.3000 76.8000 1242.6000 78.3000 ;
	    RECT 1245.0000 77.4000 1246.2001 78.6000 ;
	    RECT 1249.8000 78.4500 1251.0000 78.6000 ;
	    RECT 1269.0000 78.4500 1270.2001 78.6000 ;
	    RECT 1249.8000 77.5500 1270.2001 78.4500 ;
	    RECT 1249.8000 77.4000 1251.0000 77.5500 ;
	    RECT 1269.0000 77.4000 1270.2001 77.5500 ;
	    RECT 1247.1000 76.5000 1248.3000 77.1000 ;
	    RECT 1245.3000 76.2000 1248.3000 76.5000 ;
	    RECT 1249.8000 76.2000 1251.0000 76.5000 ;
	    RECT 1176.0000 70.2000 1179.0000 71.1000 ;
	    RECT 1163.4000 63.3000 1164.6000 67.5000 ;
	    RECT 1165.8000 63.3000 1167.0000 67.5000 ;
	    RECT 1168.2001 63.3000 1169.4000 69.3000 ;
	    RECT 1170.6000 63.3000 1171.8000 70.2000 ;
	    RECT 1176.0000 69.3000 1176.9000 70.2000 ;
	    RECT 1173.0000 62.4000 1174.2001 69.3000 ;
	    RECT 1175.4000 68.4000 1176.9000 69.3000 ;
	    RECT 1175.4000 63.3000 1176.6000 68.4000 ;
	    RECT 1177.8000 63.3000 1179.0000 69.3000 ;
	    RECT 1204.2001 63.3000 1205.4000 75.3000 ;
	    RECT 1208.1000 74.4000 1209.6000 75.3000 ;
	    RECT 1211.4000 74.4000 1212.6000 75.6000 ;
	    RECT 1247.4000 75.3000 1248.3000 76.2000 ;
	    RECT 1257.0000 75.4500 1258.2001 75.6000 ;
	    RECT 1276.2001 75.4500 1277.4000 75.6000 ;
	    RECT 1240.2001 74.4000 1246.2001 75.3000 ;
	    RECT 1208.1000 63.3000 1209.3000 74.4000 ;
	    RECT 1210.5000 72.6000 1211.4000 73.5000 ;
	    RECT 1210.2001 71.4000 1211.4000 72.6000 ;
	    RECT 1210.5000 63.3000 1211.7001 69.3000 ;
	    RECT 1240.2001 63.3000 1241.4000 74.4000 ;
	    RECT 1242.6000 63.3000 1243.8000 73.5000 ;
	    RECT 1245.0000 64.2000 1246.2001 74.4000 ;
	    RECT 1247.4000 65.1000 1248.6000 75.3000 ;
	    RECT 1249.8000 64.2000 1251.0000 75.3000 ;
	    RECT 1257.0000 74.5500 1277.4000 75.4500 ;
	    RECT 1257.0000 74.4000 1258.2001 74.5500 ;
	    RECT 1276.2001 74.4000 1277.4000 74.5500 ;
	    RECT 1279.2001 75.3000 1280.1000 80.4000 ;
	    RECT 1281.0000 79.5000 1282.2001 79.8000 ;
	    RECT 1305.0000 79.5000 1306.2001 83.7000 ;
	    RECT 1307.4000 82.5000 1308.6000 82.8000 ;
	    RECT 1326.6000 82.5000 1327.8000 82.8000 ;
	    RECT 1307.4000 81.4500 1308.6000 81.6000 ;
	    RECT 1314.6000 81.4500 1315.8000 81.6000 ;
	    RECT 1307.4000 80.5500 1315.8000 81.4500 ;
	    RECT 1307.4000 80.4000 1308.6000 80.5500 ;
	    RECT 1314.6000 80.4000 1315.8000 80.5500 ;
	    RECT 1321.8000 81.4500 1323.0000 81.6000 ;
	    RECT 1326.6000 81.4500 1327.8000 81.6000 ;
	    RECT 1321.8000 80.5500 1327.8000 81.4500 ;
	    RECT 1321.8000 80.4000 1323.0000 80.5500 ;
	    RECT 1326.6000 80.4000 1327.8000 80.5500 ;
	    RECT 1329.0000 79.5000 1330.2001 83.7000 ;
	    RECT 1362.9000 82.5000 1363.8000 83.7000 ;
	    RECT 1365.3000 83.1000 1370.7001 83.7000 ;
	    RECT 1384.2001 82.5000 1385.4000 89.7000 ;
	    RECT 1386.6000 86.7000 1387.8000 89.7000 ;
	    RECT 1401.0000 86.7000 1402.2001 89.7000 ;
	    RECT 1386.6000 85.5000 1387.8000 85.8000 ;
	    RECT 1401.0000 85.5000 1402.2001 85.8000 ;
	    RECT 1386.6000 84.4500 1387.8000 84.6000 ;
	    RECT 1398.6000 84.4500 1399.8000 84.6000 ;
	    RECT 1386.6000 83.5500 1399.8000 84.4500 ;
	    RECT 1386.6000 83.4000 1387.8000 83.5500 ;
	    RECT 1398.6000 83.4000 1399.8000 83.5500 ;
	    RECT 1401.0000 83.4000 1402.2001 84.6000 ;
	    RECT 1403.4000 82.5000 1404.6000 89.7000 ;
	    RECT 1427.4000 84.0000 1428.6000 89.7000 ;
	    RECT 1429.8000 84.9000 1431.0000 89.7000 ;
	    RECT 1432.2001 84.0000 1433.4000 89.7000 ;
	    RECT 1427.4000 83.7000 1433.4000 84.0000 ;
	    RECT 1434.6000 83.7000 1435.8000 89.7000 ;
	    RECT 1458.6000 86.7000 1459.8000 89.7000 ;
	    RECT 1458.9000 85.5000 1460.1000 85.8000 ;
	    RECT 1456.2001 84.4500 1457.4000 84.6000 ;
	    RECT 1458.6000 84.4500 1459.8000 84.6000 ;
	    RECT 1427.7001 83.1000 1433.1000 83.7000 ;
	    RECT 1434.6000 82.5000 1435.5000 83.7000 ;
	    RECT 1456.2001 83.5500 1459.8000 84.4500 ;
	    RECT 1461.0000 83.7000 1462.2001 89.7000 ;
	    RECT 1464.9000 83.7000 1466.1000 89.7000 ;
	    RECT 1456.2001 83.4000 1457.4000 83.5500 ;
	    RECT 1458.6000 83.4000 1459.8000 83.5500 ;
	    RECT 1362.6000 80.4000 1363.8000 81.6000 ;
	    RECT 1364.7001 80.4000 1366.5000 81.6000 ;
	    RECT 1368.6000 80.7000 1368.9000 82.2000 ;
	    RECT 1369.8000 80.4000 1371.0000 81.6000 ;
	    RECT 1384.2001 81.4500 1385.4000 81.6000 ;
	    RECT 1372.3500 80.5500 1385.4000 81.4500 ;
	    RECT 1281.0000 77.4000 1282.2001 78.6000 ;
	    RECT 1283.4000 78.4500 1284.6000 78.6000 ;
	    RECT 1305.0000 78.4500 1306.2001 78.6000 ;
	    RECT 1283.4000 77.5500 1306.2001 78.4500 ;
	    RECT 1283.4000 77.4000 1284.6000 77.5500 ;
	    RECT 1305.0000 77.4000 1306.2001 77.5500 ;
	    RECT 1329.0000 78.4500 1330.2001 78.6000 ;
	    RECT 1329.0000 77.5500 1363.6500 78.4500 ;
	    RECT 1329.0000 77.4000 1330.2001 77.5500 ;
	    RECT 1279.2001 74.4000 1280.7001 75.3000 ;
	    RECT 1277.4000 72.6000 1278.3000 73.5000 ;
	    RECT 1277.4000 71.4000 1278.6000 72.6000 ;
	    RECT 1245.0000 63.3000 1251.0000 64.2000 ;
	    RECT 1277.1000 63.3000 1278.3000 69.3000 ;
	    RECT 1279.5000 63.3000 1280.7001 74.4000 ;
	    RECT 1283.4000 63.3000 1284.6000 75.3000 ;
	    RECT 1302.6000 74.4000 1303.8000 75.6000 ;
	    RECT 1302.6000 73.2000 1303.8000 73.5000 ;
	    RECT 1302.6000 63.3000 1303.8000 69.3000 ;
	    RECT 1305.0000 63.3000 1306.2001 76.5000 ;
	    RECT 1307.4000 63.3000 1308.6000 69.3000 ;
	    RECT 1326.6000 63.3000 1327.8000 69.3000 ;
	    RECT 1329.0000 63.3000 1330.2001 76.5000 ;
	    RECT 1362.7500 75.6000 1363.6500 77.5500 ;
	    RECT 1331.4000 75.4500 1332.6000 75.6000 ;
	    RECT 1350.6000 75.4500 1351.8000 75.6000 ;
	    RECT 1331.4000 74.5500 1351.8000 75.4500 ;
	    RECT 1331.4000 74.4000 1332.6000 74.5500 ;
	    RECT 1350.6000 74.4000 1351.8000 74.5500 ;
	    RECT 1362.6000 74.4000 1363.8000 75.6000 ;
	    RECT 1365.6000 75.3000 1366.5000 80.4000 ;
	    RECT 1367.4000 79.5000 1368.6000 79.8000 ;
	    RECT 1367.4000 78.4500 1368.6000 78.6000 ;
	    RECT 1372.3500 78.4500 1373.2500 80.5500 ;
	    RECT 1384.2001 80.4000 1385.4000 80.5500 ;
	    RECT 1403.4000 81.4500 1404.6000 81.6000 ;
	    RECT 1403.4000 80.5500 1426.0500 81.4500 ;
	    RECT 1403.4000 80.4000 1404.6000 80.5500 ;
	    RECT 1367.4000 77.5500 1373.2500 78.4500 ;
	    RECT 1367.4000 77.4000 1368.6000 77.5500 ;
	    RECT 1365.6000 74.4000 1367.1000 75.3000 ;
	    RECT 1331.4000 73.2000 1332.6000 73.5000 ;
	    RECT 1363.8000 72.6000 1364.7001 73.5000 ;
	    RECT 1363.8000 71.4000 1365.0000 72.6000 ;
	    RECT 1331.4000 63.3000 1332.6000 69.3000 ;
	    RECT 1363.5000 63.3000 1364.7001 69.3000 ;
	    RECT 1365.9000 63.3000 1367.1000 74.4000 ;
	    RECT 1369.8000 63.3000 1371.0000 75.3000 ;
	    RECT 1384.2001 63.3000 1385.4000 79.5000 ;
	    RECT 1386.6000 63.3000 1387.8000 69.3000 ;
	    RECT 1401.0000 63.3000 1402.2001 69.3000 ;
	    RECT 1403.4000 63.3000 1404.6000 79.5000 ;
	    RECT 1425.1500 78.4500 1426.0500 80.5500 ;
	    RECT 1427.4000 80.4000 1428.6000 81.6000 ;
	    RECT 1429.5000 80.7000 1429.8000 82.2000 ;
	    RECT 1431.9000 80.4000 1433.7001 81.6000 ;
	    RECT 1434.6000 81.4500 1435.8000 81.6000 ;
	    RECT 1458.6000 81.4500 1459.8000 81.6000 ;
	    RECT 1434.6000 80.5500 1459.8000 81.4500 ;
	    RECT 1434.6000 80.4000 1435.8000 80.5500 ;
	    RECT 1458.6000 80.4000 1459.8000 80.5500 ;
	    RECT 1429.8000 79.5000 1431.0000 79.8000 ;
	    RECT 1429.8000 78.4500 1431.0000 78.6000 ;
	    RECT 1425.1500 77.5500 1431.0000 78.4500 ;
	    RECT 1429.8000 77.4000 1431.0000 77.5500 ;
	    RECT 1431.9000 75.3000 1432.8000 80.4000 ;
	    RECT 1458.6000 77.4000 1459.8000 78.6000 ;
	    RECT 1461.3000 78.3000 1462.2001 83.7000 ;
	    RECT 1463.4000 81.4500 1464.6000 81.6000 ;
	    RECT 1485.0000 81.4500 1486.2001 81.6000 ;
	    RECT 1463.4000 80.5500 1486.2001 81.4500 ;
	    RECT 1489.8000 80.7000 1491.0000 89.7000 ;
	    RECT 1495.2001 81.3000 1496.4000 89.7000 ;
	    RECT 1495.2001 80.7000 1497.9000 81.3000 ;
	    RECT 1521.0000 80.7000 1522.2001 89.7000 ;
	    RECT 1526.4000 81.3000 1527.6000 89.7000 ;
	    RECT 1526.4000 80.7000 1529.1000 81.3000 ;
	    RECT 1552.2001 80.7000 1553.4000 89.7000 ;
	    RECT 1557.6000 81.3000 1558.8000 89.7000 ;
	    RECT 1557.6000 80.7000 1560.3000 81.3000 ;
	    RECT 1463.4000 80.4000 1464.6000 80.5500 ;
	    RECT 1485.0000 80.4000 1486.2001 80.5500 ;
	    RECT 1495.5000 80.4000 1497.9000 80.7000 ;
	    RECT 1526.7001 80.4000 1529.1000 80.7000 ;
	    RECT 1557.9000 80.4000 1560.3000 80.7000 ;
	    RECT 1463.4000 79.2000 1464.6000 79.5000 ;
	    RECT 1460.7001 77.4000 1462.2001 78.3000 ;
	    RECT 1464.6000 76.8000 1464.9000 78.3000 ;
	    RECT 1465.8000 77.4000 1467.0000 78.6000 ;
	    RECT 1492.2001 77.4000 1493.4000 78.6000 ;
	    RECT 1494.3000 77.4000 1494.6000 78.6000 ;
	    RECT 1489.8000 76.5000 1491.0000 76.8000 ;
	    RECT 1497.0000 76.5000 1497.9000 80.4000 ;
	    RECT 1523.4000 77.4000 1524.6000 78.6000 ;
	    RECT 1525.5000 77.4000 1525.8000 78.6000 ;
	    RECT 1521.0000 76.5000 1522.2001 76.8000 ;
	    RECT 1528.2001 76.5000 1529.1000 80.4000 ;
	    RECT 1554.6000 77.4000 1555.8000 78.6000 ;
	    RECT 1556.7001 77.4000 1557.0000 78.6000 ;
	    RECT 1552.2001 76.5000 1553.4000 76.8000 ;
	    RECT 1559.4000 76.5000 1560.3000 80.4000 ;
	    RECT 1427.4000 63.3000 1428.6000 75.3000 ;
	    RECT 1431.3000 74.4000 1432.8000 75.3000 ;
	    RECT 1434.6000 74.4000 1435.8000 75.6000 ;
	    RECT 1458.9000 75.3000 1459.8000 76.5000 ;
	    RECT 1431.3000 63.3000 1432.5000 74.4000 ;
	    RECT 1433.7001 72.6000 1434.6000 73.5000 ;
	    RECT 1433.4000 71.4000 1434.6000 72.6000 ;
	    RECT 1433.7001 63.3000 1434.9000 69.3000 ;
	    RECT 1458.6000 63.3000 1459.8000 75.3000 ;
	    RECT 1461.0000 74.4000 1467.0000 75.3000 ;
	    RECT 1489.8000 74.4000 1491.0000 75.6000 ;
	    RECT 1497.0000 75.4500 1498.2001 75.6000 ;
	    RECT 1497.0000 74.5500 1519.6500 75.4500 ;
	    RECT 1497.0000 74.4000 1498.2001 74.5500 ;
	    RECT 1461.0000 63.3000 1462.2001 74.4000 ;
	    RECT 1463.4000 63.3000 1464.6000 73.5000 ;
	    RECT 1465.8000 63.3000 1467.0000 74.4000 ;
	    RECT 1494.6000 73.5000 1495.8000 73.8000 ;
	    RECT 1480.2001 72.4500 1481.4000 72.6000 ;
	    RECT 1494.6000 72.4500 1495.8000 72.6000 ;
	    RECT 1480.2001 71.5500 1495.8000 72.4500 ;
	    RECT 1480.2001 71.4000 1481.4000 71.5500 ;
	    RECT 1494.6000 71.4000 1495.8000 71.5500 ;
	    RECT 1497.0000 70.5000 1497.9000 73.5000 ;
	    RECT 1518.7500 72.4500 1519.6500 74.5500 ;
	    RECT 1521.0000 74.4000 1522.2001 75.6000 ;
	    RECT 1528.2001 75.4500 1529.4000 75.6000 ;
	    RECT 1545.0000 75.4500 1546.2001 75.6000 ;
	    RECT 1528.2001 74.5500 1546.2001 75.4500 ;
	    RECT 1528.2001 74.4000 1529.4000 74.5500 ;
	    RECT 1545.0000 74.4000 1546.2001 74.5500 ;
	    RECT 1547.4000 75.4500 1548.6000 75.6000 ;
	    RECT 1552.2001 75.4500 1553.4000 75.6000 ;
	    RECT 1547.4000 74.5500 1553.4000 75.4500 ;
	    RECT 1547.4000 74.4000 1548.6000 74.5500 ;
	    RECT 1552.2001 74.4000 1553.4000 74.5500 ;
	    RECT 1559.4000 75.4500 1560.6000 75.6000 ;
	    RECT 1564.2001 75.4500 1565.4000 75.6000 ;
	    RECT 1559.4000 74.5500 1565.4000 75.4500 ;
	    RECT 1559.4000 74.4000 1560.6000 74.5500 ;
	    RECT 1564.2001 74.4000 1565.4000 74.5500 ;
	    RECT 1525.8000 73.5000 1527.0000 73.8000 ;
	    RECT 1557.0000 73.5000 1558.2001 73.8000 ;
	    RECT 1525.8000 72.4500 1527.0000 72.6000 ;
	    RECT 1518.7500 71.5500 1527.0000 72.4500 ;
	    RECT 1525.8000 71.4000 1527.0000 71.5500 ;
	    RECT 1528.2001 70.5000 1529.1000 73.5000 ;
	    RECT 1557.0000 71.4000 1558.2001 72.6000 ;
	    RECT 1559.4000 70.5000 1560.3000 73.5000 ;
	    RECT 1492.5000 69.6000 1497.9000 70.5000 ;
	    RECT 1492.5000 69.3000 1493.4000 69.6000 ;
	    RECT 1489.8000 63.3000 1491.0000 69.3000 ;
	    RECT 1492.2001 63.3000 1493.4000 69.3000 ;
	    RECT 1497.0000 69.3000 1497.9000 69.6000 ;
	    RECT 1523.7001 69.6000 1529.1000 70.5000 ;
	    RECT 1523.7001 69.3000 1524.6000 69.6000 ;
	    RECT 1494.6000 63.3000 1495.8000 68.7000 ;
	    RECT 1497.0000 63.3000 1498.2001 69.3000 ;
	    RECT 1521.0000 63.3000 1522.2001 69.3000 ;
	    RECT 1523.4000 63.3000 1524.6000 69.3000 ;
	    RECT 1528.2001 69.3000 1529.1000 69.6000 ;
	    RECT 1554.9000 69.6000 1560.3000 70.5000 ;
	    RECT 1554.9000 69.3000 1555.8000 69.6000 ;
	    RECT 1525.8000 63.3000 1527.0000 68.7000 ;
	    RECT 1528.2001 63.3000 1529.4000 69.3000 ;
	    RECT 1552.2001 63.3000 1553.4000 69.3000 ;
	    RECT 1554.6000 63.3000 1555.8000 69.3000 ;
	    RECT 1559.4000 69.3000 1560.3000 69.6000 ;
	    RECT 1557.0000 63.3000 1558.2001 68.7000 ;
	    RECT 1559.4000 63.3000 1560.6000 69.3000 ;
	    RECT 1.2000 60.6000 1569.0000 62.4000 ;
	    RECT 124.2000 53.7000 125.4000 59.7000 ;
	    RECT 126.6000 52.5000 127.8000 59.7000 ;
	    RECT 129.0000 53.7000 130.2000 59.7000 ;
	    RECT 131.4000 52.8000 132.6000 59.7000 ;
	    RECT 133.8000 53.7000 135.0000 59.7000 ;
	    RECT 128.7000 51.9000 132.6000 52.8000 ;
	    RECT 23.4000 51.4500 24.6000 51.6000 ;
	    RECT 126.6000 51.4500 127.8000 51.6000 ;
	    RECT 23.4000 50.5500 127.8000 51.4500 ;
	    RECT 23.4000 50.4000 24.6000 50.5500 ;
	    RECT 126.6000 50.4000 127.8000 50.5500 ;
	    RECT 128.7000 49.5000 129.6000 51.9000 ;
	    RECT 136.2000 51.6000 137.4000 59.7000 ;
	    RECT 138.6000 53.7000 139.8000 59.7000 ;
	    RECT 141.0000 55.5000 142.2000 59.7000 ;
	    RECT 143.4000 55.5000 144.6000 59.7000 ;
	    RECT 145.8000 55.5000 147.0000 59.7000 ;
	    RECT 138.3000 51.6000 144.6000 52.8000 ;
	    RECT 133.5000 50.4000 137.4000 51.6000 ;
	    RECT 148.2000 50.4000 149.4000 59.7000 ;
	    RECT 150.6000 53.7000 151.8000 59.7000 ;
	    RECT 153.0000 52.5000 154.2000 59.7000 ;
	    RECT 155.4000 53.7000 156.6000 59.7000 ;
	    RECT 157.8000 52.5000 159.0000 59.7000 ;
	    RECT 160.2000 55.5000 161.4000 59.7000 ;
	    RECT 162.6000 55.5000 163.8000 59.7000 ;
	    RECT 165.0000 53.7000 166.2000 59.7000 ;
	    RECT 167.4000 52.8000 168.6000 59.7000 ;
	    RECT 169.8000 53.7000 171.0000 60.6000 ;
	    RECT 172.2000 54.6000 173.4000 59.7000 ;
	    RECT 172.2000 53.7000 173.7000 54.6000 ;
	    RECT 174.6000 53.7000 175.8000 59.7000 ;
	    RECT 306.6000 53.7000 307.8000 59.7000 ;
	    RECT 172.8000 52.8000 173.7000 53.7000 ;
	    RECT 165.6000 51.6000 171.9000 52.8000 ;
	    RECT 172.8000 51.9000 175.8000 52.8000 ;
	    RECT 309.0000 52.5000 310.2000 59.7000 ;
	    RECT 311.4000 53.7000 312.6000 59.7000 ;
	    RECT 313.8000 52.8000 315.0000 59.7000 ;
	    RECT 316.2000 53.7000 317.4000 59.7000 ;
	    RECT 153.0000 50.4000 156.9000 51.6000 ;
	    RECT 157.8000 50.7000 166.5000 51.6000 ;
	    RECT 171.0000 51.0000 171.9000 51.6000 ;
	    RECT 141.0000 49.5000 142.2000 49.8000 ;
	    RECT 126.6000 48.0000 127.8000 49.5000 ;
	    RECT 126.3000 46.8000 127.8000 48.0000 ;
	    RECT 128.7000 48.6000 142.2000 49.5000 ;
	    RECT 145.8000 49.5000 147.0000 49.8000 ;
	    RECT 157.8000 49.5000 158.7000 50.7000 ;
	    RECT 167.4000 49.8000 169.5000 50.7000 ;
	    RECT 171.0000 49.8000 173.4000 51.0000 ;
	    RECT 145.8000 48.6000 158.7000 49.5000 ;
	    RECT 160.2000 49.5000 169.5000 49.8000 ;
	    RECT 160.2000 48.9000 168.3000 49.5000 ;
	    RECT 160.2000 48.6000 161.4000 48.9000 ;
	    RECT 126.3000 40.2000 127.5000 46.8000 ;
	    RECT 128.7000 45.9000 129.6000 48.6000 ;
	    RECT 164.7000 47.7000 165.9000 48.0000 ;
	    RECT 130.5000 46.8000 168.9000 47.7000 ;
	    RECT 169.8000 47.4000 171.0000 48.6000 ;
	    RECT 130.5000 46.5000 131.7000 46.8000 ;
	    RECT 128.4000 45.0000 129.6000 45.9000 ;
	    RECT 138.6000 45.0000 164.1000 45.9000 ;
	    RECT 128.4000 42.0000 129.3000 45.0000 ;
	    RECT 138.6000 44.1000 139.8000 45.0000 ;
	    RECT 165.0000 44.4000 166.2000 45.6000 ;
	    RECT 167.1000 45.0000 173.7000 45.9000 ;
	    RECT 172.5000 44.7000 173.7000 45.0000 ;
	    RECT 130.2000 42.9000 135.9000 44.1000 ;
	    RECT 128.4000 41.1000 130.2000 42.0000 ;
	    RECT 126.3000 39.0000 127.8000 40.2000 ;
	    RECT 124.2000 33.3000 125.4000 36.3000 ;
	    RECT 126.6000 33.3000 127.8000 39.0000 ;
	    RECT 129.0000 33.3000 130.2000 41.1000 ;
	    RECT 134.7000 41.1000 135.9000 42.9000 ;
	    RECT 134.7000 40.2000 137.4000 41.1000 ;
	    RECT 136.2000 39.3000 137.4000 40.2000 ;
	    RECT 143.4000 39.6000 144.6000 43.8000 ;
	    RECT 148.2000 42.9000 153.0000 44.1000 ;
	    RECT 158.7000 42.9000 161.7000 44.1000 ;
	    RECT 174.6000 43.5000 175.8000 51.9000 ;
	    RECT 311.1000 51.9000 315.0000 52.8000 ;
	    RECT 253.8000 51.4500 255.0000 51.6000 ;
	    RECT 309.0000 51.4500 310.2000 51.6000 ;
	    RECT 253.8000 50.5500 310.2000 51.4500 ;
	    RECT 253.8000 50.4000 255.0000 50.5500 ;
	    RECT 309.0000 50.4000 310.2000 50.5500 ;
	    RECT 311.1000 49.5000 312.0000 51.9000 ;
	    RECT 318.6000 51.6000 319.8000 59.7000 ;
	    RECT 321.0000 53.7000 322.2000 59.7000 ;
	    RECT 323.4000 55.5000 324.6000 59.7000 ;
	    RECT 325.8000 55.5000 327.0000 59.7000 ;
	    RECT 328.2000 55.5000 329.4000 59.7000 ;
	    RECT 320.7000 51.6000 327.0000 52.8000 ;
	    RECT 315.9000 50.4000 319.8000 51.6000 ;
	    RECT 330.6000 50.4000 331.8000 59.7000 ;
	    RECT 333.0000 53.7000 334.2000 59.7000 ;
	    RECT 335.4000 52.5000 336.6000 59.7000 ;
	    RECT 337.8000 53.7000 339.0000 59.7000 ;
	    RECT 340.2000 52.5000 341.4000 59.7000 ;
	    RECT 342.6000 55.5000 343.8000 59.7000 ;
	    RECT 345.0000 55.5000 346.2000 59.7000 ;
	    RECT 347.4000 53.7000 348.6000 59.7000 ;
	    RECT 349.8000 52.8000 351.0000 59.7000 ;
	    RECT 352.2000 53.7000 353.4000 60.6000 ;
	    RECT 354.6000 54.6000 355.8000 59.7000 ;
	    RECT 354.6000 53.7000 356.1000 54.6000 ;
	    RECT 357.0000 53.7000 358.2000 59.7000 ;
	    RECT 371.4000 53.7000 372.6000 59.7000 ;
	    RECT 355.2000 52.8000 356.1000 53.7000 ;
	    RECT 348.0000 51.6000 354.3000 52.8000 ;
	    RECT 355.2000 51.9000 358.2000 52.8000 ;
	    RECT 335.4000 50.4000 339.3000 51.6000 ;
	    RECT 340.2000 50.7000 348.9000 51.6000 ;
	    RECT 353.4000 51.0000 354.3000 51.6000 ;
	    RECT 323.4000 49.5000 324.6000 49.8000 ;
	    RECT 309.0000 48.0000 310.2000 49.5000 ;
	    RECT 147.6000 41.7000 148.8000 42.0000 ;
	    RECT 147.6000 40.8000 154.2000 41.7000 ;
	    RECT 155.4000 41.4000 156.6000 42.6000 ;
	    RECT 153.0000 40.5000 154.2000 40.8000 ;
	    RECT 155.4000 40.2000 156.6000 40.5000 ;
	    RECT 133.8000 33.3000 135.0000 39.3000 ;
	    RECT 136.2000 38.1000 139.8000 39.3000 ;
	    RECT 143.4000 38.4000 144.9000 39.6000 ;
	    RECT 149.4000 38.4000 149.7000 39.6000 ;
	    RECT 150.6000 38.4000 151.8000 39.6000 ;
	    RECT 153.0000 39.3000 154.2000 39.6000 ;
	    RECT 158.7000 39.3000 159.9000 42.9000 ;
	    RECT 162.6000 42.3000 175.8000 43.5000 ;
	    RECT 167.7000 40.2000 172.2000 41.4000 ;
	    RECT 167.7000 39.3000 168.9000 40.2000 ;
	    RECT 153.0000 38.4000 159.9000 39.3000 ;
	    RECT 138.6000 33.3000 139.8000 38.1000 ;
	    RECT 165.0000 38.1000 168.9000 39.3000 ;
	    RECT 141.0000 33.3000 142.2000 37.5000 ;
	    RECT 143.4000 33.3000 144.6000 37.5000 ;
	    RECT 145.8000 33.3000 147.0000 37.5000 ;
	    RECT 148.2000 33.3000 149.4000 37.5000 ;
	    RECT 150.6000 33.3000 151.8000 36.3000 ;
	    RECT 153.0000 33.3000 154.2000 37.5000 ;
	    RECT 155.4000 33.3000 156.6000 36.3000 ;
	    RECT 157.8000 33.3000 159.0000 37.5000 ;
	    RECT 160.2000 33.3000 161.4000 37.5000 ;
	    RECT 162.6000 33.3000 163.8000 37.5000 ;
	    RECT 165.0000 33.3000 166.2000 38.1000 ;
	    RECT 169.8000 33.3000 171.0000 39.3000 ;
	    RECT 174.6000 33.3000 175.8000 42.3000 ;
	    RECT 308.7000 46.8000 310.2000 48.0000 ;
	    RECT 311.1000 48.6000 324.6000 49.5000 ;
	    RECT 328.2000 49.5000 329.4000 49.8000 ;
	    RECT 340.2000 49.5000 341.1000 50.7000 ;
	    RECT 349.8000 49.8000 351.9000 50.7000 ;
	    RECT 353.4000 49.8000 355.8000 51.0000 ;
	    RECT 328.2000 48.6000 341.1000 49.5000 ;
	    RECT 342.6000 49.5000 351.9000 49.8000 ;
	    RECT 342.6000 48.9000 350.7000 49.5000 ;
	    RECT 342.6000 48.6000 343.8000 48.9000 ;
	    RECT 308.7000 40.2000 309.9000 46.8000 ;
	    RECT 311.1000 45.9000 312.0000 48.6000 ;
	    RECT 347.1000 47.7000 348.3000 48.0000 ;
	    RECT 312.9000 46.8000 351.3000 47.7000 ;
	    RECT 352.2000 47.4000 353.4000 48.6000 ;
	    RECT 312.9000 46.5000 314.1000 46.8000 ;
	    RECT 310.8000 45.0000 312.0000 45.9000 ;
	    RECT 321.0000 45.0000 346.5000 45.9000 ;
	    RECT 310.8000 42.0000 311.7000 45.0000 ;
	    RECT 321.0000 44.1000 322.2000 45.0000 ;
	    RECT 347.4000 44.4000 348.6000 45.6000 ;
	    RECT 349.5000 45.0000 356.1000 45.9000 ;
	    RECT 354.9000 44.7000 356.1000 45.0000 ;
	    RECT 312.6000 42.9000 318.3000 44.1000 ;
	    RECT 310.8000 41.1000 312.6000 42.0000 ;
	    RECT 308.7000 39.0000 310.2000 40.2000 ;
	    RECT 306.6000 33.3000 307.8000 36.3000 ;
	    RECT 309.0000 33.3000 310.2000 39.0000 ;
	    RECT 311.4000 33.3000 312.6000 41.1000 ;
	    RECT 317.1000 41.1000 318.3000 42.9000 ;
	    RECT 317.1000 40.2000 319.8000 41.1000 ;
	    RECT 318.6000 39.3000 319.8000 40.2000 ;
	    RECT 325.8000 39.6000 327.0000 43.8000 ;
	    RECT 330.6000 42.9000 335.4000 44.1000 ;
	    RECT 341.1000 42.9000 344.1000 44.1000 ;
	    RECT 357.0000 43.5000 358.2000 51.9000 ;
	    RECT 373.8000 43.5000 375.0000 59.7000 ;
	    RECT 397.8000 47.7000 399.0000 59.7000 ;
	    RECT 401.7000 48.6000 402.9000 59.7000 ;
	    RECT 404.1000 53.7000 405.3000 59.7000 ;
	    RECT 424.2000 53.7000 425.4000 59.7000 ;
	    RECT 403.8000 50.4000 405.0000 51.6000 ;
	    RECT 404.1000 49.5000 405.0000 50.4000 ;
	    RECT 401.7000 47.7000 403.2000 48.6000 ;
	    RECT 400.2000 45.4500 401.4000 45.6000 ;
	    RECT 395.5500 44.5500 401.4000 45.4500 ;
	    RECT 330.0000 41.7000 331.2000 42.0000 ;
	    RECT 330.0000 40.8000 336.6000 41.7000 ;
	    RECT 337.8000 41.4000 339.0000 42.6000 ;
	    RECT 335.4000 40.5000 336.6000 40.8000 ;
	    RECT 337.8000 40.2000 339.0000 40.5000 ;
	    RECT 316.2000 33.3000 317.4000 39.3000 ;
	    RECT 318.6000 38.1000 322.2000 39.3000 ;
	    RECT 325.8000 38.4000 327.3000 39.6000 ;
	    RECT 331.8000 38.4000 332.1000 39.6000 ;
	    RECT 333.0000 38.4000 334.2000 39.6000 ;
	    RECT 335.4000 39.3000 336.6000 39.6000 ;
	    RECT 341.1000 39.3000 342.3000 42.9000 ;
	    RECT 345.0000 42.3000 358.2000 43.5000 ;
	    RECT 350.1000 40.2000 354.6000 41.4000 ;
	    RECT 350.1000 39.3000 351.3000 40.2000 ;
	    RECT 335.4000 38.4000 342.3000 39.3000 ;
	    RECT 321.0000 33.3000 322.2000 38.1000 ;
	    RECT 347.4000 38.1000 351.3000 39.3000 ;
	    RECT 323.4000 33.3000 324.6000 37.5000 ;
	    RECT 325.8000 33.3000 327.0000 37.5000 ;
	    RECT 328.2000 33.3000 329.4000 37.5000 ;
	    RECT 330.6000 33.3000 331.8000 37.5000 ;
	    RECT 333.0000 33.3000 334.2000 36.3000 ;
	    RECT 335.4000 33.3000 336.6000 37.5000 ;
	    RECT 337.8000 33.3000 339.0000 36.3000 ;
	    RECT 340.2000 33.3000 341.4000 37.5000 ;
	    RECT 342.6000 33.3000 343.8000 37.5000 ;
	    RECT 345.0000 33.3000 346.2000 37.5000 ;
	    RECT 347.4000 33.3000 348.6000 38.1000 ;
	    RECT 352.2000 33.3000 353.4000 39.3000 ;
	    RECT 357.0000 33.3000 358.2000 42.3000 ;
	    RECT 373.8000 42.4500 375.0000 42.6000 ;
	    RECT 395.5500 42.4500 396.4500 44.5500 ;
	    RECT 400.2000 44.4000 401.4000 44.5500 ;
	    RECT 400.2000 43.2000 401.4000 43.5000 ;
	    RECT 402.3000 42.6000 403.2000 47.7000 ;
	    RECT 405.0000 47.4000 406.2000 48.6000 ;
	    RECT 405.1500 45.4500 406.0500 47.4000 ;
	    RECT 426.6000 46.5000 427.8000 59.7000 ;
	    RECT 429.0000 53.7000 430.2000 59.7000 ;
	    RECT 429.0000 49.5000 430.2000 49.8000 ;
	    RECT 429.0000 47.4000 430.2000 48.6000 ;
	    RECT 460.2000 47.7000 461.4000 59.7000 ;
	    RECT 464.1000 48.6000 465.3000 59.7000 ;
	    RECT 466.5000 53.7000 467.7000 59.7000 ;
	    RECT 494.7000 53.7000 495.9000 59.7000 ;
	    RECT 466.2000 50.4000 467.4000 51.6000 ;
	    RECT 466.5000 49.5000 467.4000 50.4000 ;
	    RECT 495.0000 50.4000 496.2000 51.6000 ;
	    RECT 495.0000 49.5000 495.9000 50.4000 ;
	    RECT 497.1000 48.6000 498.3000 59.7000 ;
	    RECT 464.1000 47.7000 465.6000 48.6000 ;
	    RECT 426.6000 45.4500 427.8000 45.6000 ;
	    RECT 405.1500 44.5500 427.8000 45.4500 ;
	    RECT 426.6000 44.4000 427.8000 44.5500 ;
	    RECT 460.2000 45.4500 461.4000 45.6000 ;
	    RECT 462.6000 45.4500 463.8000 45.6000 ;
	    RECT 460.2000 44.5500 463.8000 45.4500 ;
	    RECT 460.2000 44.4000 461.4000 44.5500 ;
	    RECT 462.6000 44.4000 463.8000 44.5500 ;
	    RECT 373.8000 41.5500 396.4500 42.4500 ;
	    RECT 373.8000 41.4000 375.0000 41.5500 ;
	    RECT 397.8000 41.4000 399.0000 42.6000 ;
	    RECT 399.9000 40.8000 400.2000 42.3000 ;
	    RECT 402.3000 41.4000 404.1000 42.6000 ;
	    RECT 405.0000 42.4500 406.2000 42.6000 ;
	    RECT 421.8000 42.4500 423.0000 42.6000 ;
	    RECT 405.0000 41.5500 423.0000 42.4500 ;
	    RECT 405.0000 41.4000 406.2000 41.5500 ;
	    RECT 421.8000 41.4000 423.0000 41.5500 ;
	    RECT 424.2000 41.4000 425.4000 42.6000 ;
	    RECT 369.0000 39.4500 370.2000 39.6000 ;
	    RECT 371.4000 39.4500 372.6000 39.6000 ;
	    RECT 369.0000 38.5500 372.6000 39.4500 ;
	    RECT 369.0000 38.4000 370.2000 38.5500 ;
	    RECT 371.4000 38.4000 372.6000 38.5500 ;
	    RECT 371.4000 37.2000 372.6000 37.5000 ;
	    RECT 371.4000 33.3000 372.6000 36.3000 ;
	    RECT 373.8000 33.3000 375.0000 40.5000 ;
	    RECT 398.1000 39.3000 403.5000 39.9000 ;
	    RECT 405.0000 39.3000 405.9000 40.5000 ;
	    RECT 424.2000 40.2000 425.4000 40.5000 ;
	    RECT 426.6000 39.3000 427.8000 43.5000 ;
	    RECT 462.6000 43.2000 463.8000 43.5000 ;
	    RECT 464.7000 42.6000 465.6000 47.7000 ;
	    RECT 467.4000 48.4500 468.6000 48.6000 ;
	    RECT 469.8000 48.4500 471.0000 48.6000 ;
	    RECT 467.4000 47.5500 471.0000 48.4500 ;
	    RECT 467.4000 47.4000 468.6000 47.5500 ;
	    RECT 469.8000 47.4000 471.0000 47.5500 ;
	    RECT 493.8000 47.4000 495.0000 48.6000 ;
	    RECT 496.8000 47.7000 498.3000 48.6000 ;
	    RECT 501.0000 47.7000 502.2000 59.7000 ;
	    RECT 503.4000 59.4000 504.6000 60.6000 ;
	    RECT 520.2000 53.7000 521.4000 59.7000 ;
	    RECT 496.8000 42.6000 497.7000 47.7000 ;
	    RECT 522.6000 46.5000 523.8000 59.7000 ;
	    RECT 525.0000 53.7000 526.2000 59.7000 ;
	    RECT 525.0000 49.5000 526.2000 49.8000 ;
	    RECT 498.6000 44.4000 499.8000 45.6000 ;
	    RECT 501.0000 45.4500 502.2000 45.6000 ;
	    RECT 522.6000 45.4500 523.8000 45.6000 ;
	    RECT 501.0000 44.5500 523.8000 45.4500 ;
	    RECT 501.0000 44.4000 502.2000 44.5500 ;
	    RECT 522.6000 44.4000 523.8000 44.5500 ;
	    RECT 537.0000 43.5000 538.2000 59.7000 ;
	    RECT 539.4000 53.7000 540.6000 59.7000 ;
	    RECT 671.4000 53.7000 672.6000 59.7000 ;
	    RECT 673.8000 52.5000 675.0000 59.7000 ;
	    RECT 676.2000 53.7000 677.4000 59.7000 ;
	    RECT 678.6000 52.8000 679.8000 59.7000 ;
	    RECT 681.0000 53.7000 682.2000 59.7000 ;
	    RECT 675.9000 51.9000 679.8000 52.8000 ;
	    RECT 585.0000 51.4500 586.2000 51.6000 ;
	    RECT 673.8000 51.4500 675.0000 51.6000 ;
	    RECT 585.0000 50.5500 675.0000 51.4500 ;
	    RECT 585.0000 50.4000 586.2000 50.5500 ;
	    RECT 673.8000 50.4000 675.0000 50.5500 ;
	    RECT 675.9000 49.5000 676.8000 51.9000 ;
	    RECT 683.4000 51.6000 684.6000 59.7000 ;
	    RECT 685.8000 53.7000 687.0000 59.7000 ;
	    RECT 688.2000 55.5000 689.4000 59.7000 ;
	    RECT 690.6000 55.5000 691.8000 59.7000 ;
	    RECT 693.0000 55.5000 694.2000 59.7000 ;
	    RECT 685.5000 51.6000 691.8000 52.8000 ;
	    RECT 680.7000 50.4000 684.6000 51.6000 ;
	    RECT 695.4000 50.4000 696.6000 59.7000 ;
	    RECT 697.8000 53.7000 699.0000 59.7000 ;
	    RECT 700.2000 52.5000 701.4000 59.7000 ;
	    RECT 702.6000 53.7000 703.8000 59.7000 ;
	    RECT 705.0000 52.5000 706.2000 59.7000 ;
	    RECT 707.4000 55.5000 708.6000 59.7000 ;
	    RECT 709.8000 55.5000 711.0000 59.7000 ;
	    RECT 712.2000 53.7000 713.4000 59.7000 ;
	    RECT 714.6000 52.8000 715.8000 59.7000 ;
	    RECT 717.0000 53.7000 718.2000 60.6000 ;
	    RECT 719.4000 54.6000 720.6000 59.7000 ;
	    RECT 719.4000 53.7000 720.9000 54.6000 ;
	    RECT 721.8000 53.7000 723.0000 59.7000 ;
	    RECT 736.2000 53.7000 737.4000 59.7000 ;
	    RECT 720.0000 52.8000 720.9000 53.7000 ;
	    RECT 712.8000 51.6000 719.1000 52.8000 ;
	    RECT 720.0000 51.9000 723.0000 52.8000 ;
	    RECT 700.2000 50.4000 704.1000 51.6000 ;
	    RECT 705.0000 50.7000 713.7000 51.6000 ;
	    RECT 718.2000 51.0000 719.1000 51.6000 ;
	    RECT 688.2000 49.5000 689.4000 49.8000 ;
	    RECT 673.8000 48.0000 675.0000 49.5000 ;
	    RECT 673.5000 46.8000 675.0000 48.0000 ;
	    RECT 675.9000 48.6000 689.4000 49.5000 ;
	    RECT 693.0000 49.5000 694.2000 49.8000 ;
	    RECT 705.0000 49.5000 705.9000 50.7000 ;
	    RECT 714.6000 49.8000 716.7000 50.7000 ;
	    RECT 718.2000 49.8000 720.6000 51.0000 ;
	    RECT 693.0000 48.6000 705.9000 49.5000 ;
	    RECT 707.4000 49.5000 716.7000 49.8000 ;
	    RECT 707.4000 48.9000 715.5000 49.5000 ;
	    RECT 707.4000 48.6000 708.6000 48.9000 ;
	    RECT 498.6000 43.2000 499.8000 43.5000 ;
	    RECT 457.8000 42.4500 459.0000 42.6000 ;
	    RECT 460.2000 42.4500 461.4000 42.6000 ;
	    RECT 457.8000 41.5500 461.4000 42.4500 ;
	    RECT 457.8000 41.4000 459.0000 41.5500 ;
	    RECT 460.2000 41.4000 461.4000 41.5500 ;
	    RECT 462.3000 40.8000 462.6000 42.3000 ;
	    RECT 464.7000 41.4000 466.5000 42.6000 ;
	    RECT 467.4000 42.4500 468.6000 42.6000 ;
	    RECT 486.6000 42.4500 487.8000 42.6000 ;
	    RECT 467.4000 41.5500 487.8000 42.4500 ;
	    RECT 467.4000 41.4000 468.6000 41.5500 ;
	    RECT 486.6000 41.4000 487.8000 41.5500 ;
	    RECT 491.4000 42.4500 492.6000 42.6000 ;
	    RECT 493.8000 42.4500 495.0000 42.6000 ;
	    RECT 491.4000 41.5500 495.0000 42.4500 ;
	    RECT 491.4000 41.4000 492.6000 41.5500 ;
	    RECT 493.8000 41.4000 495.0000 41.5500 ;
	    RECT 495.9000 41.4000 497.7000 42.6000 ;
	    RECT 501.0000 42.4500 502.2000 42.6000 ;
	    RECT 503.4000 42.4500 504.6000 42.6000 ;
	    RECT 499.8000 40.8000 500.1000 42.3000 ;
	    RECT 501.0000 41.5500 504.6000 42.4500 ;
	    RECT 501.0000 41.4000 502.2000 41.5500 ;
	    RECT 503.4000 41.4000 504.6000 41.5500 ;
	    RECT 520.2000 41.4000 521.4000 42.6000 ;
	    RECT 460.5000 39.3000 465.9000 39.9000 ;
	    RECT 467.4000 39.3000 468.3000 40.5000 ;
	    RECT 494.1000 39.3000 495.0000 40.5000 ;
	    RECT 520.2000 40.2000 521.4000 40.5000 ;
	    RECT 496.5000 39.3000 501.9000 39.9000 ;
	    RECT 522.6000 39.3000 523.8000 43.5000 ;
	    RECT 525.0000 42.4500 526.2000 42.6000 ;
	    RECT 537.0000 42.4500 538.2000 42.6000 ;
	    RECT 525.0000 41.5500 538.2000 42.4500 ;
	    RECT 525.0000 41.4000 526.2000 41.5500 ;
	    RECT 537.0000 41.4000 538.2000 41.5500 ;
	    RECT 397.8000 39.0000 403.8000 39.3000 ;
	    RECT 397.8000 33.3000 399.0000 39.0000 ;
	    RECT 400.2000 33.3000 401.4000 38.1000 ;
	    RECT 402.6000 33.3000 403.8000 39.0000 ;
	    RECT 405.0000 33.3000 406.2000 39.3000 ;
	    RECT 424.2000 33.3000 425.4000 39.3000 ;
	    RECT 426.6000 38.4000 429.3000 39.3000 ;
	    RECT 428.1000 33.3000 429.3000 38.4000 ;
	    RECT 460.2000 39.0000 466.2000 39.3000 ;
	    RECT 460.2000 33.3000 461.4000 39.0000 ;
	    RECT 462.6000 33.3000 463.8000 38.1000 ;
	    RECT 465.0000 33.3000 466.2000 39.0000 ;
	    RECT 467.4000 33.3000 468.6000 39.3000 ;
	    RECT 493.8000 33.3000 495.0000 39.3000 ;
	    RECT 496.2000 39.0000 502.2000 39.3000 ;
	    RECT 496.2000 33.3000 497.4000 39.0000 ;
	    RECT 498.6000 33.3000 499.8000 38.1000 ;
	    RECT 501.0000 33.3000 502.2000 39.0000 ;
	    RECT 520.2000 33.3000 521.4000 39.3000 ;
	    RECT 522.6000 38.4000 525.3000 39.3000 ;
	    RECT 524.1000 33.3000 525.3000 38.4000 ;
	    RECT 537.0000 33.3000 538.2000 40.5000 ;
	    RECT 673.5000 40.2000 674.7000 46.8000 ;
	    RECT 675.9000 45.9000 676.8000 48.6000 ;
	    RECT 711.9000 47.7000 713.1000 48.0000 ;
	    RECT 677.7000 46.8000 716.1000 47.7000 ;
	    RECT 717.0000 47.4000 718.2000 48.6000 ;
	    RECT 677.7000 46.5000 678.9000 46.8000 ;
	    RECT 675.6000 45.0000 676.8000 45.9000 ;
	    RECT 685.8000 45.0000 711.3000 45.9000 ;
	    RECT 675.6000 42.0000 676.5000 45.0000 ;
	    RECT 685.8000 44.1000 687.0000 45.0000 ;
	    RECT 712.2000 44.4000 713.4000 45.6000 ;
	    RECT 714.3000 45.0000 720.9000 45.9000 ;
	    RECT 719.7000 44.7000 720.9000 45.0000 ;
	    RECT 677.4000 42.9000 683.1000 44.1000 ;
	    RECT 675.6000 41.1000 677.4000 42.0000 ;
	    RECT 539.4000 39.4500 540.6000 39.6000 ;
	    RECT 544.2000 39.4500 545.4000 39.6000 ;
	    RECT 539.4000 38.5500 545.4000 39.4500 ;
	    RECT 673.5000 39.0000 675.0000 40.2000 ;
	    RECT 539.4000 38.4000 540.6000 38.5500 ;
	    RECT 544.2000 38.4000 545.4000 38.5500 ;
	    RECT 539.4000 37.2000 540.6000 37.5000 ;
	    RECT 539.4000 33.3000 540.6000 36.3000 ;
	    RECT 671.4000 33.3000 672.6000 36.3000 ;
	    RECT 673.8000 33.3000 675.0000 39.0000 ;
	    RECT 676.2000 33.3000 677.4000 41.1000 ;
	    RECT 681.9000 41.1000 683.1000 42.9000 ;
	    RECT 681.9000 40.2000 684.6000 41.1000 ;
	    RECT 683.4000 39.3000 684.6000 40.2000 ;
	    RECT 690.6000 39.6000 691.8000 43.8000 ;
	    RECT 695.4000 42.9000 700.2000 44.1000 ;
	    RECT 705.9000 42.9000 708.9000 44.1000 ;
	    RECT 721.8000 43.5000 723.0000 51.9000 ;
	    RECT 738.6000 43.5000 739.8000 59.7000 ;
	    RECT 760.2000 59.4000 761.4000 60.6000 ;
	    RECT 762.6000 47.7000 763.8000 59.7000 ;
	    RECT 766.5000 48.6000 767.7000 59.7000 ;
	    RECT 768.9000 53.7000 770.1000 59.7000 ;
	    RECT 794.7000 53.7000 795.9000 59.7000 ;
	    RECT 768.6000 50.4000 769.8000 51.6000 ;
	    RECT 768.9000 49.5000 769.8000 50.4000 ;
	    RECT 795.0000 50.4000 796.2000 51.6000 ;
	    RECT 795.0000 49.5000 795.9000 50.4000 ;
	    RECT 797.1000 48.6000 798.3000 59.7000 ;
	    RECT 766.5000 47.7000 768.0000 48.6000 ;
	    RECT 765.0000 44.4000 766.2000 45.6000 ;
	    RECT 694.8000 41.7000 696.0000 42.0000 ;
	    RECT 694.8000 40.8000 701.4000 41.7000 ;
	    RECT 702.6000 41.4000 703.8000 42.6000 ;
	    RECT 700.2000 40.5000 701.4000 40.8000 ;
	    RECT 702.6000 40.2000 703.8000 40.5000 ;
	    RECT 681.0000 33.3000 682.2000 39.3000 ;
	    RECT 683.4000 38.1000 687.0000 39.3000 ;
	    RECT 690.6000 38.4000 692.1000 39.6000 ;
	    RECT 696.6000 38.4000 696.9000 39.6000 ;
	    RECT 697.8000 38.4000 699.0000 39.6000 ;
	    RECT 700.2000 39.3000 701.4000 39.6000 ;
	    RECT 705.9000 39.3000 707.1000 42.9000 ;
	    RECT 709.8000 42.3000 723.0000 43.5000 ;
	    RECT 765.0000 43.2000 766.2000 43.5000 ;
	    RECT 767.1000 42.6000 768.0000 47.7000 ;
	    RECT 769.8000 48.4500 771.0000 48.6000 ;
	    RECT 774.6000 48.4500 775.8000 48.6000 ;
	    RECT 769.8000 47.5500 775.8000 48.4500 ;
	    RECT 769.8000 47.4000 771.0000 47.5500 ;
	    RECT 774.6000 47.4000 775.8000 47.5500 ;
	    RECT 793.8000 47.4000 795.0000 48.6000 ;
	    RECT 796.8000 47.7000 798.3000 48.6000 ;
	    RECT 801.0000 47.7000 802.2000 59.7000 ;
	    RECT 832.2000 59.4000 833.4000 60.6000 ;
	    RECT 839.4000 59.4000 840.6000 60.6000 ;
	    RECT 885.0000 57.4500 886.2000 57.6000 ;
	    RECT 911.5500 57.4500 912.4500 60.6000 ;
	    RECT 885.0000 56.5500 912.4500 57.4500 ;
	    RECT 885.0000 56.4000 886.2000 56.5500 ;
	    RECT 933.0000 53.7000 934.2000 59.7000 ;
	    RECT 935.4000 52.5000 936.6000 59.7000 ;
	    RECT 937.8000 53.7000 939.0000 59.7000 ;
	    RECT 940.2000 52.8000 941.4000 59.7000 ;
	    RECT 942.6000 53.7000 943.8000 59.7000 ;
	    RECT 937.5000 51.9000 941.4000 52.8000 ;
	    RECT 856.2000 51.4500 857.4000 51.6000 ;
	    RECT 935.4000 51.4500 936.6000 51.6000 ;
	    RECT 856.2000 50.5500 936.6000 51.4500 ;
	    RECT 856.2000 50.4000 857.4000 50.5500 ;
	    RECT 935.4000 50.4000 936.6000 50.5500 ;
	    RECT 937.5000 49.5000 938.4000 51.9000 ;
	    RECT 945.0000 51.6000 946.2000 59.7000 ;
	    RECT 947.4000 53.7000 948.6000 59.7000 ;
	    RECT 949.8000 55.5000 951.0000 59.7000 ;
	    RECT 952.2000 55.5000 953.4000 59.7000 ;
	    RECT 954.6000 55.5000 955.8000 59.7000 ;
	    RECT 947.1000 51.6000 953.4000 52.8000 ;
	    RECT 942.3000 50.4000 946.2000 51.6000 ;
	    RECT 957.0000 50.4000 958.2000 59.7000 ;
	    RECT 959.4000 53.7000 960.6000 59.7000 ;
	    RECT 961.8000 52.5000 963.0000 59.7000 ;
	    RECT 964.2000 53.7000 965.4000 59.7000 ;
	    RECT 966.6000 52.5000 967.8000 59.7000 ;
	    RECT 969.0000 55.5000 970.2000 59.7000 ;
	    RECT 971.4000 55.5000 972.6000 59.7000 ;
	    RECT 973.8000 53.7000 975.0000 59.7000 ;
	    RECT 976.2000 52.8000 977.4000 59.7000 ;
	    RECT 978.6000 53.7000 979.8000 60.6000 ;
	    RECT 981.0000 54.6000 982.2000 59.7000 ;
	    RECT 981.0000 53.7000 982.5000 54.6000 ;
	    RECT 983.4000 53.7000 984.6000 59.7000 ;
	    RECT 1008.3000 53.7000 1009.5000 59.7000 ;
	    RECT 981.6000 52.8000 982.5000 53.7000 ;
	    RECT 974.4000 51.6000 980.7000 52.8000 ;
	    RECT 981.6000 51.9000 984.6000 52.8000 ;
	    RECT 961.8000 50.4000 965.7000 51.6000 ;
	    RECT 966.6000 50.7000 975.3000 51.6000 ;
	    RECT 979.8000 51.0000 980.7000 51.6000 ;
	    RECT 949.8000 49.5000 951.0000 49.8000 ;
	    RECT 935.4000 48.0000 936.6000 49.5000 ;
	    RECT 796.8000 42.6000 797.7000 47.7000 ;
	    RECT 935.1000 46.8000 936.6000 48.0000 ;
	    RECT 937.5000 48.6000 951.0000 49.5000 ;
	    RECT 954.6000 49.5000 955.8000 49.8000 ;
	    RECT 966.6000 49.5000 967.5000 50.7000 ;
	    RECT 976.2000 49.8000 978.3000 50.7000 ;
	    RECT 979.8000 49.8000 982.2000 51.0000 ;
	    RECT 954.6000 48.6000 967.5000 49.5000 ;
	    RECT 969.0000 49.5000 978.3000 49.8000 ;
	    RECT 969.0000 48.9000 977.1000 49.5000 ;
	    RECT 969.0000 48.6000 970.2000 48.9000 ;
	    RECT 798.6000 44.4000 799.8000 45.6000 ;
	    RECT 798.6000 43.2000 799.8000 43.5000 ;
	    RECT 714.9000 40.2000 719.4000 41.4000 ;
	    RECT 714.9000 39.3000 716.1000 40.2000 ;
	    RECT 700.2000 38.4000 707.1000 39.3000 ;
	    RECT 685.8000 33.3000 687.0000 38.1000 ;
	    RECT 712.2000 38.1000 716.1000 39.3000 ;
	    RECT 688.2000 33.3000 689.4000 37.5000 ;
	    RECT 690.6000 33.3000 691.8000 37.5000 ;
	    RECT 693.0000 33.3000 694.2000 37.5000 ;
	    RECT 695.4000 33.3000 696.6000 37.5000 ;
	    RECT 697.8000 33.3000 699.0000 36.3000 ;
	    RECT 700.2000 33.3000 701.4000 37.5000 ;
	    RECT 702.6000 33.3000 703.8000 36.3000 ;
	    RECT 705.0000 33.3000 706.2000 37.5000 ;
	    RECT 707.4000 33.3000 708.6000 37.5000 ;
	    RECT 709.8000 33.3000 711.0000 37.5000 ;
	    RECT 712.2000 33.3000 713.4000 38.1000 ;
	    RECT 717.0000 33.3000 718.2000 39.3000 ;
	    RECT 721.8000 33.3000 723.0000 42.3000 ;
	    RECT 724.2000 42.4500 725.4000 42.6000 ;
	    RECT 738.6000 42.4500 739.8000 42.6000 ;
	    RECT 724.2000 41.5500 739.8000 42.4500 ;
	    RECT 724.2000 41.4000 725.4000 41.5500 ;
	    RECT 738.6000 41.4000 739.8000 41.5500 ;
	    RECT 760.2000 42.4500 761.4000 42.6000 ;
	    RECT 762.6000 42.4500 763.8000 42.6000 ;
	    RECT 760.2000 41.5500 763.8000 42.4500 ;
	    RECT 760.2000 41.4000 761.4000 41.5500 ;
	    RECT 762.6000 41.4000 763.8000 41.5500 ;
	    RECT 764.7000 40.8000 765.0000 42.3000 ;
	    RECT 767.1000 41.4000 768.9000 42.6000 ;
	    RECT 769.8000 41.4000 771.0000 42.6000 ;
	    RECT 772.2000 42.4500 773.4000 42.6000 ;
	    RECT 793.8000 42.4500 795.0000 42.6000 ;
	    RECT 772.2000 41.5500 795.0000 42.4500 ;
	    RECT 772.2000 41.4000 773.4000 41.5500 ;
	    RECT 793.8000 41.4000 795.0000 41.5500 ;
	    RECT 795.9000 41.4000 797.7000 42.6000 ;
	    RECT 801.0000 42.4500 802.2000 42.6000 ;
	    RECT 832.2000 42.4500 833.4000 42.6000 ;
	    RECT 799.8000 40.8000 800.1000 42.3000 ;
	    RECT 801.0000 41.5500 833.4000 42.4500 ;
	    RECT 801.0000 41.4000 802.2000 41.5500 ;
	    RECT 832.2000 41.4000 833.4000 41.5500 ;
	    RECT 731.4000 39.4500 732.6000 39.6000 ;
	    RECT 736.2000 39.4500 737.4000 39.6000 ;
	    RECT 731.4000 38.5500 737.4000 39.4500 ;
	    RECT 731.4000 38.4000 732.6000 38.5500 ;
	    RECT 736.2000 38.4000 737.4000 38.5500 ;
	    RECT 736.2000 37.2000 737.4000 37.5000 ;
	    RECT 736.2000 33.3000 737.4000 36.3000 ;
	    RECT 738.6000 33.3000 739.8000 40.5000 ;
	    RECT 762.9000 39.3000 768.3000 39.9000 ;
	    RECT 769.8000 39.3000 770.7000 40.5000 ;
	    RECT 794.1000 39.3000 795.0000 40.5000 ;
	    RECT 935.1000 40.2000 936.3000 46.8000 ;
	    RECT 937.5000 45.9000 938.4000 48.6000 ;
	    RECT 973.5000 47.7000 974.7000 48.0000 ;
	    RECT 939.3000 46.8000 977.7000 47.7000 ;
	    RECT 978.6000 47.4000 979.8000 48.6000 ;
	    RECT 939.3000 46.5000 940.5000 46.8000 ;
	    RECT 937.2000 45.0000 938.4000 45.9000 ;
	    RECT 947.4000 45.0000 972.9000 45.9000 ;
	    RECT 937.2000 42.0000 938.1000 45.0000 ;
	    RECT 947.4000 44.1000 948.6000 45.0000 ;
	    RECT 973.8000 44.4000 975.0000 45.6000 ;
	    RECT 975.9000 45.0000 982.5000 45.9000 ;
	    RECT 981.3000 44.7000 982.5000 45.0000 ;
	    RECT 939.0000 42.9000 944.7000 44.1000 ;
	    RECT 937.2000 41.1000 939.0000 42.0000 ;
	    RECT 796.5000 39.3000 801.9000 39.9000 ;
	    RECT 762.6000 39.0000 768.6000 39.3000 ;
	    RECT 762.6000 33.3000 763.8000 39.0000 ;
	    RECT 765.0000 33.3000 766.2000 38.1000 ;
	    RECT 767.4000 33.3000 768.6000 39.0000 ;
	    RECT 769.8000 33.3000 771.0000 39.3000 ;
	    RECT 793.8000 33.3000 795.0000 39.3000 ;
	    RECT 796.2000 39.0000 802.2000 39.3000 ;
	    RECT 935.1000 39.0000 936.6000 40.2000 ;
	    RECT 796.2000 33.3000 797.4000 39.0000 ;
	    RECT 798.6000 33.3000 799.8000 38.1000 ;
	    RECT 801.0000 33.3000 802.2000 39.0000 ;
	    RECT 933.0000 33.3000 934.2000 36.3000 ;
	    RECT 935.4000 33.3000 936.6000 39.0000 ;
	    RECT 937.8000 33.3000 939.0000 41.1000 ;
	    RECT 943.5000 41.1000 944.7000 42.9000 ;
	    RECT 943.5000 40.2000 946.2000 41.1000 ;
	    RECT 945.0000 39.3000 946.2000 40.2000 ;
	    RECT 952.2000 39.6000 953.4000 43.8000 ;
	    RECT 957.0000 42.9000 961.8000 44.1000 ;
	    RECT 967.5000 42.9000 970.5000 44.1000 ;
	    RECT 983.4000 43.5000 984.6000 51.9000 ;
	    RECT 1008.6000 50.4000 1009.8000 51.6000 ;
	    RECT 1008.6000 49.5000 1009.5000 50.4000 ;
	    RECT 1010.7000 48.6000 1011.9000 59.7000 ;
	    RECT 990.6000 48.4500 991.8000 48.6000 ;
	    RECT 1007.4000 48.4500 1008.6000 48.6000 ;
	    RECT 990.6000 47.5500 1008.6000 48.4500 ;
	    RECT 990.6000 47.4000 991.8000 47.5500 ;
	    RECT 1007.4000 47.4000 1008.6000 47.5500 ;
	    RECT 1010.4000 47.7000 1011.9000 48.6000 ;
	    RECT 1014.6000 47.7000 1015.8000 59.7000 ;
	    RECT 1055.4000 48.6000 1056.6000 59.7000 ;
	    RECT 1057.8000 49.8000 1059.3000 59.7000 ;
	    RECT 1058.1000 48.6000 1059.3000 48.9000 ;
	    RECT 1055.4000 47.7000 1059.3000 48.6000 ;
	    RECT 1062.0000 47.7000 1064.4000 59.7000 ;
	    RECT 1067.1000 49.8000 1068.6000 59.7000 ;
	    RECT 1067.4000 48.6000 1068.6000 48.9000 ;
	    RECT 1069.8000 48.6000 1071.0000 59.7000 ;
	    RECT 1067.4000 47.7000 1071.0000 48.6000 ;
	    RECT 1089.0000 48.6000 1090.2001 59.7000 ;
	    RECT 1091.4000 49.5000 1092.6000 59.7000 ;
	    RECT 1089.0000 47.7000 1092.3000 48.6000 ;
	    RECT 1093.8000 47.7000 1095.0000 59.7000 ;
	    RECT 1139.4000 59.4000 1140.6000 60.6000 ;
	    RECT 1141.8000 48.6000 1143.0000 59.7000 ;
	    RECT 1144.2001 49.8000 1145.7001 59.7000 ;
	    RECT 1144.5000 48.6000 1145.7001 48.9000 ;
	    RECT 1141.8000 47.7000 1145.7001 48.6000 ;
	    RECT 1148.4000 47.7000 1150.8000 59.7000 ;
	    RECT 1153.5000 49.8000 1155.0000 59.7000 ;
	    RECT 1153.8000 48.6000 1155.0000 48.9000 ;
	    RECT 1156.2001 48.6000 1157.4000 59.7000 ;
	    RECT 1175.4000 53.7000 1176.6000 59.7000 ;
	    RECT 1175.4000 49.5000 1176.6000 49.8000 ;
	    RECT 1153.8000 47.7000 1157.4000 48.6000 ;
	    RECT 956.4000 41.7000 957.6000 42.0000 ;
	    RECT 956.4000 40.8000 963.0000 41.7000 ;
	    RECT 964.2000 41.4000 965.4000 42.6000 ;
	    RECT 961.8000 40.5000 963.0000 40.8000 ;
	    RECT 964.2000 40.2000 965.4000 40.5000 ;
	    RECT 942.6000 33.3000 943.8000 39.3000 ;
	    RECT 945.0000 38.1000 948.6000 39.3000 ;
	    RECT 952.2000 38.4000 953.7000 39.6000 ;
	    RECT 958.2000 38.4000 958.5000 39.6000 ;
	    RECT 959.4000 38.4000 960.6000 39.6000 ;
	    RECT 961.8000 39.3000 963.0000 39.6000 ;
	    RECT 967.5000 39.3000 968.7000 42.9000 ;
	    RECT 971.4000 42.3000 984.6000 43.5000 ;
	    RECT 1010.4000 42.6000 1011.3000 47.7000 ;
	    RECT 1062.9000 46.5000 1063.8000 47.7000 ;
	    RECT 1091.4000 46.8000 1092.3000 47.7000 ;
	    RECT 1059.9000 45.6000 1061.1000 45.9000 ;
	    RECT 1091.4000 45.6000 1093.2001 46.8000 ;
	    RECT 1012.2000 44.4000 1013.4000 45.6000 ;
	    RECT 1058.7001 44.7000 1061.1000 45.6000 ;
	    RECT 1062.6000 45.4500 1063.8000 45.6000 ;
	    RECT 1086.6000 45.4500 1087.8000 45.6000 ;
	    RECT 1058.7001 44.4000 1059.9000 44.7000 ;
	    RECT 1062.6000 44.5500 1087.8000 45.4500 ;
	    RECT 1062.6000 44.4000 1063.8000 44.5500 ;
	    RECT 1086.6000 44.4000 1087.8000 44.5500 ;
	    RECT 1089.0000 44.4000 1090.2001 45.6000 ;
	    RECT 1012.2000 43.2000 1013.4000 43.5000 ;
	    RECT 1060.8000 42.9000 1062.0000 43.2000 ;
	    RECT 1057.8000 42.6000 1062.0000 42.9000 ;
	    RECT 976.5000 40.2000 981.0000 41.4000 ;
	    RECT 976.5000 39.3000 977.7000 40.2000 ;
	    RECT 961.8000 38.4000 968.7000 39.3000 ;
	    RECT 947.4000 33.3000 948.6000 38.1000 ;
	    RECT 973.8000 38.1000 977.7000 39.3000 ;
	    RECT 949.8000 33.3000 951.0000 37.5000 ;
	    RECT 952.2000 33.3000 953.4000 37.5000 ;
	    RECT 954.6000 33.3000 955.8000 37.5000 ;
	    RECT 957.0000 33.3000 958.2000 37.5000 ;
	    RECT 959.4000 33.3000 960.6000 36.3000 ;
	    RECT 961.8000 33.3000 963.0000 37.5000 ;
	    RECT 964.2000 33.3000 965.4000 36.3000 ;
	    RECT 966.6000 33.3000 967.8000 37.5000 ;
	    RECT 969.0000 33.3000 970.2000 37.5000 ;
	    RECT 971.4000 33.3000 972.6000 37.5000 ;
	    RECT 973.8000 33.3000 975.0000 38.1000 ;
	    RECT 978.6000 33.3000 979.8000 39.3000 ;
	    RECT 983.4000 33.3000 984.6000 42.3000 ;
	    RECT 1007.4000 41.4000 1008.6000 42.6000 ;
	    RECT 1009.5000 41.4000 1011.3000 42.6000 ;
	    RECT 1014.6000 42.4500 1015.8000 42.6000 ;
	    RECT 1026.6000 42.4500 1027.8000 42.6000 ;
	    RECT 1013.4000 40.8000 1013.7000 42.3000 ;
	    RECT 1014.6000 41.5500 1027.8000 42.4500 ;
	    RECT 1014.6000 41.4000 1015.8000 41.5500 ;
	    RECT 1026.6000 41.4000 1027.8000 41.5500 ;
	    RECT 1055.4000 41.4000 1056.6000 42.6000 ;
	    RECT 1057.5000 42.0000 1062.0000 42.6000 ;
	    RECT 1062.9000 42.6000 1063.8000 43.5000 ;
	    RECT 1089.0000 43.2000 1090.2001 43.5000 ;
	    RECT 1057.5000 41.7000 1058.7001 42.0000 ;
	    RECT 1062.9000 41.7000 1064.4000 42.6000 ;
	    RECT 1057.5000 41.4000 1057.8000 41.7000 ;
	    RECT 1007.7000 39.3000 1008.6000 40.5000 ;
	    RECT 1058.1000 40.2000 1059.3000 40.5000 ;
	    RECT 1010.1000 39.3000 1015.5000 39.9000 ;
	    RECT 1055.4000 39.3000 1059.3000 40.2000 ;
	    RECT 1060.2001 39.6000 1062.6000 40.8000 ;
	    RECT 1007.4000 33.3000 1008.6000 39.3000 ;
	    RECT 1009.8000 39.0000 1015.8000 39.3000 ;
	    RECT 1009.8000 33.3000 1011.0000 39.0000 ;
	    RECT 1012.2000 33.3000 1013.4000 38.1000 ;
	    RECT 1014.6000 33.3000 1015.8000 39.0000 ;
	    RECT 1055.4000 33.3000 1056.6000 39.3000 ;
	    RECT 1063.5000 38.7000 1064.4000 41.7000 ;
	    RECT 1065.6000 41.4000 1066.8000 42.6000 ;
	    RECT 1068.6000 41.4000 1068.9000 42.6000 ;
	    RECT 1069.8000 41.4000 1071.0000 42.6000 ;
	    RECT 1065.6000 40.8000 1066.5000 41.4000 ;
	    RECT 1091.4000 41.1000 1092.3000 45.6000 ;
	    RECT 1094.1000 44.4000 1095.0000 47.7000 ;
	    RECT 1149.3000 46.5000 1150.2001 47.7000 ;
	    RECT 1175.4000 47.4000 1176.6000 48.6000 ;
	    RECT 1177.8000 46.5000 1179.0000 59.7000 ;
	    RECT 1180.2001 53.7000 1181.4000 59.7000 ;
	    RECT 1194.6000 53.7000 1195.8000 59.7000 ;
	    RECT 1146.3000 45.6000 1147.5000 45.9000 ;
	    RECT 1145.1000 44.7000 1147.5000 45.6000 ;
	    RECT 1149.0000 45.4500 1150.2001 45.6000 ;
	    RECT 1173.0000 45.4500 1174.2001 45.6000 ;
	    RECT 1145.1000 44.4000 1146.3000 44.7000 ;
	    RECT 1149.0000 44.5500 1174.2001 45.4500 ;
	    RECT 1149.0000 44.4000 1150.2001 44.5500 ;
	    RECT 1173.0000 44.4000 1174.2001 44.5500 ;
	    RECT 1177.8000 44.4000 1179.0000 45.6000 ;
	    RECT 1093.8000 43.5000 1095.0000 44.4000 ;
	    RECT 1197.0000 43.5000 1198.2001 59.7000 ;
	    RECT 1237.8000 48.6000 1239.0000 59.7000 ;
	    RECT 1240.2001 49.8000 1241.7001 59.7000 ;
	    RECT 1240.2001 48.6000 1241.4000 48.9000 ;
	    RECT 1237.8000 47.7000 1241.4000 48.6000 ;
	    RECT 1244.4000 47.7000 1246.8000 59.7000 ;
	    RECT 1249.5000 49.8000 1251.0000 59.7000 ;
	    RECT 1249.5000 48.6000 1250.7001 48.9000 ;
	    RECT 1252.2001 48.6000 1253.4000 59.7000 ;
	    RECT 1386.6000 53.7000 1387.8000 59.7000 ;
	    RECT 1389.0000 54.6000 1390.2001 59.7000 ;
	    RECT 1388.7001 53.7000 1390.2001 54.6000 ;
	    RECT 1391.4000 53.7000 1392.6000 60.6000 ;
	    RECT 1388.7001 52.8000 1389.6000 53.7000 ;
	    RECT 1393.8000 52.8000 1395.0000 59.7000 ;
	    RECT 1396.2001 53.7000 1397.4000 59.7000 ;
	    RECT 1398.6000 55.5000 1399.8000 59.7000 ;
	    RECT 1401.0000 55.5000 1402.2001 59.7000 ;
	    RECT 1249.5000 47.7000 1253.4000 48.6000 ;
	    RECT 1386.6000 51.9000 1389.6000 52.8000 ;
	    RECT 1245.0000 46.5000 1245.9000 47.7000 ;
	    RECT 1247.7001 45.6000 1248.9000 45.9000 ;
	    RECT 1213.8000 45.4500 1215.0000 45.6000 ;
	    RECT 1204.3500 44.5500 1215.0000 45.4500 ;
	    RECT 1147.2001 42.9000 1148.4000 43.2000 ;
	    RECT 1144.2001 42.6000 1148.4000 42.9000 ;
	    RECT 1141.8000 41.4000 1143.0000 42.6000 ;
	    RECT 1143.9000 42.0000 1148.4000 42.6000 ;
	    RECT 1149.3000 42.6000 1150.2001 43.5000 ;
	    RECT 1143.9000 41.7000 1145.1000 42.0000 ;
	    RECT 1149.3000 41.7000 1150.8000 42.6000 ;
	    RECT 1143.9000 41.4000 1144.2001 41.7000 ;
	    RECT 1065.3000 39.6000 1066.5000 40.8000 ;
	    RECT 1067.4000 40.2000 1068.6000 40.5000 ;
	    RECT 1089.0000 40.2000 1092.3000 41.1000 ;
	    RECT 1067.4000 39.3000 1071.0000 40.2000 ;
	    RECT 1057.8000 33.3000 1059.3000 38.4000 ;
	    RECT 1062.0000 33.3000 1064.4000 38.7000 ;
	    RECT 1067.1000 33.3000 1068.6000 38.4000 ;
	    RECT 1069.8000 33.3000 1071.0000 39.3000 ;
	    RECT 1089.0000 33.3000 1090.2001 40.2000 ;
	    RECT 1091.4000 33.3000 1092.6000 39.3000 ;
	    RECT 1093.8000 33.3000 1095.0000 40.5000 ;
	    RECT 1144.5000 40.2000 1145.7001 40.5000 ;
	    RECT 1141.8000 39.3000 1145.7001 40.2000 ;
	    RECT 1146.6000 39.6000 1149.0000 40.8000 ;
	    RECT 1141.8000 33.3000 1143.0000 39.3000 ;
	    RECT 1149.9000 38.7000 1150.8000 41.7000 ;
	    RECT 1152.0000 41.4000 1153.2001 42.6000 ;
	    RECT 1155.0000 41.4000 1155.3000 42.6000 ;
	    RECT 1156.2001 41.4000 1157.4000 42.6000 ;
	    RECT 1152.0000 40.8000 1152.9000 41.4000 ;
	    RECT 1151.7001 39.6000 1152.9000 40.8000 ;
	    RECT 1153.8000 40.2000 1155.0000 40.5000 ;
	    RECT 1153.8000 39.3000 1157.4000 40.2000 ;
	    RECT 1177.8000 39.3000 1179.0000 43.5000 ;
	    RECT 1180.2001 41.4000 1181.4000 42.6000 ;
	    RECT 1197.0000 42.4500 1198.2001 42.6000 ;
	    RECT 1204.3500 42.4500 1205.2500 44.5500 ;
	    RECT 1213.8000 44.4000 1215.0000 44.5500 ;
	    RECT 1245.0000 44.4000 1246.2001 45.6000 ;
	    RECT 1247.7001 44.7000 1250.1000 45.6000 ;
	    RECT 1248.9000 44.4000 1250.1000 44.7000 ;
	    RECT 1386.6000 43.5000 1387.8000 51.9000 ;
	    RECT 1390.5000 51.6000 1396.8000 52.8000 ;
	    RECT 1403.4000 52.5000 1404.6000 59.7000 ;
	    RECT 1405.8000 53.7000 1407.0000 59.7000 ;
	    RECT 1408.2001 52.5000 1409.4000 59.7000 ;
	    RECT 1410.6000 53.7000 1411.8000 59.7000 ;
	    RECT 1390.5000 51.0000 1391.4000 51.6000 ;
	    RECT 1389.0000 49.8000 1391.4000 51.0000 ;
	    RECT 1395.9000 50.7000 1404.6000 51.6000 ;
	    RECT 1392.9000 49.8000 1395.0000 50.7000 ;
	    RECT 1392.9000 49.5000 1402.2001 49.8000 ;
	    RECT 1394.1000 48.9000 1402.2001 49.5000 ;
	    RECT 1401.0000 48.6000 1402.2001 48.9000 ;
	    RECT 1403.7001 49.5000 1404.6000 50.7000 ;
	    RECT 1405.5000 50.4000 1409.4000 51.6000 ;
	    RECT 1413.0000 50.4000 1414.2001 59.7000 ;
	    RECT 1415.4000 55.5000 1416.6000 59.7000 ;
	    RECT 1417.8000 55.5000 1419.0000 59.7000 ;
	    RECT 1420.2001 55.5000 1421.4000 59.7000 ;
	    RECT 1422.6000 53.7000 1423.8000 59.7000 ;
	    RECT 1417.8000 51.6000 1424.1000 52.8000 ;
	    RECT 1425.0000 51.6000 1426.2001 59.7000 ;
	    RECT 1427.4000 53.7000 1428.6000 59.7000 ;
	    RECT 1429.8000 52.8000 1431.0000 59.7000 ;
	    RECT 1432.2001 53.7000 1433.4000 59.7000 ;
	    RECT 1429.8000 51.9000 1433.7001 52.8000 ;
	    RECT 1434.6000 52.5000 1435.8000 59.7000 ;
	    RECT 1437.0000 53.7000 1438.2001 59.7000 ;
	    RECT 1425.0000 50.4000 1428.9000 51.6000 ;
	    RECT 1415.4000 49.5000 1416.6000 49.8000 ;
	    RECT 1403.7001 48.6000 1416.6000 49.5000 ;
	    RECT 1420.2001 49.5000 1421.4000 49.8000 ;
	    RECT 1432.8000 49.5000 1433.7001 51.9000 ;
	    RECT 1434.6000 50.4000 1435.8000 51.6000 ;
	    RECT 1420.2001 48.6000 1433.7001 49.5000 ;
	    RECT 1391.4000 47.4000 1392.6000 48.6000 ;
	    RECT 1396.5000 47.7000 1397.7001 48.0000 ;
	    RECT 1393.5000 46.8000 1431.9000 47.7000 ;
	    RECT 1430.7001 46.5000 1431.9000 46.8000 ;
	    RECT 1432.8000 45.9000 1433.7001 48.6000 ;
	    RECT 1434.6000 48.0000 1435.8000 49.5000 ;
	    RECT 1456.2001 48.6000 1457.4000 59.7000 ;
	    RECT 1458.6000 49.5000 1459.8000 59.7000 ;
	    RECT 1434.6000 46.8000 1436.1000 48.0000 ;
	    RECT 1456.2001 47.7000 1459.5000 48.6000 ;
	    RECT 1461.0000 47.7000 1462.2001 59.7000 ;
	    RECT 1487.4000 53.7000 1488.6000 59.7000 ;
	    RECT 1489.8000 53.7000 1491.0000 59.7000 ;
	    RECT 1492.2001 54.3000 1493.4000 59.7000 ;
	    RECT 1490.1000 53.4000 1491.0000 53.7000 ;
	    RECT 1494.6000 53.7000 1495.8000 59.7000 ;
	    RECT 1513.8000 53.7000 1515.0000 59.7000 ;
	    RECT 1494.6000 53.4000 1495.5000 53.7000 ;
	    RECT 1490.1000 52.5000 1495.5000 53.4000 ;
	    RECT 1465.8000 51.4500 1467.0000 51.6000 ;
	    RECT 1492.2001 51.4500 1493.4000 51.6000 ;
	    RECT 1465.8000 50.5500 1493.4000 51.4500 ;
	    RECT 1465.8000 50.4000 1467.0000 50.5500 ;
	    RECT 1492.2001 50.4000 1493.4000 50.5500 ;
	    RECT 1494.6000 49.5000 1495.5000 52.5000 ;
	    RECT 1513.8000 49.5000 1515.0000 49.8000 ;
	    RECT 1492.2001 49.2000 1493.4000 49.5000 ;
	    RECT 1388.7001 45.0000 1395.3000 45.9000 ;
	    RECT 1388.7001 44.7000 1389.9000 45.0000 ;
	    RECT 1396.2001 44.4000 1397.4000 45.6000 ;
	    RECT 1398.3000 45.0000 1423.8000 45.9000 ;
	    RECT 1432.8000 45.0000 1434.0000 45.9000 ;
	    RECT 1422.6000 44.1000 1423.8000 45.0000 ;
	    RECT 1245.0000 42.6000 1245.9000 43.5000 ;
	    RECT 1197.0000 41.5500 1205.2500 42.4500 ;
	    RECT 1206.6000 42.4500 1207.8000 42.6000 ;
	    RECT 1237.8000 42.4500 1239.0000 42.6000 ;
	    RECT 1206.6000 41.5500 1239.0000 42.4500 ;
	    RECT 1197.0000 41.4000 1198.2001 41.5500 ;
	    RECT 1206.6000 41.4000 1207.8000 41.5500 ;
	    RECT 1237.8000 41.4000 1239.0000 41.5500 ;
	    RECT 1239.9000 41.4000 1240.2001 42.6000 ;
	    RECT 1242.0000 41.4000 1243.2001 42.6000 ;
	    RECT 1242.3000 40.8000 1243.2001 41.4000 ;
	    RECT 1244.4000 41.7000 1245.9000 42.6000 ;
	    RECT 1246.8000 42.9000 1248.0000 43.2000 ;
	    RECT 1246.8000 42.6000 1251.0000 42.9000 ;
	    RECT 1246.8000 42.0000 1251.3000 42.6000 ;
	    RECT 1250.1000 41.7000 1251.3000 42.0000 ;
	    RECT 1180.2001 40.2000 1181.4000 40.5000 ;
	    RECT 1182.6000 39.4500 1183.8000 39.6000 ;
	    RECT 1194.6000 39.4500 1195.8000 39.6000 ;
	    RECT 1144.2001 33.3000 1145.7001 38.4000 ;
	    RECT 1148.4000 33.3000 1150.8000 38.7000 ;
	    RECT 1153.5000 33.3000 1155.0000 38.4000 ;
	    RECT 1156.2001 33.3000 1157.4000 39.3000 ;
	    RECT 1176.3000 38.4000 1179.0000 39.3000 ;
	    RECT 1176.3000 33.3000 1177.5000 38.4000 ;
	    RECT 1180.2001 33.3000 1181.4000 39.3000 ;
	    RECT 1182.6000 38.5500 1195.8000 39.4500 ;
	    RECT 1182.6000 38.4000 1183.8000 38.5500 ;
	    RECT 1194.6000 38.4000 1195.8000 38.5500 ;
	    RECT 1194.6000 37.2000 1195.8000 37.5000 ;
	    RECT 1194.6000 33.3000 1195.8000 36.3000 ;
	    RECT 1197.0000 33.3000 1198.2001 40.5000 ;
	    RECT 1240.2001 40.2000 1241.4000 40.5000 ;
	    RECT 1237.8000 39.3000 1241.4000 40.2000 ;
	    RECT 1242.3000 39.6000 1243.5000 40.8000 ;
	    RECT 1237.8000 33.3000 1239.0000 39.3000 ;
	    RECT 1244.4000 38.7000 1245.3000 41.7000 ;
	    RECT 1251.0000 41.4000 1251.3000 41.7000 ;
	    RECT 1252.2001 41.4000 1253.4000 42.6000 ;
	    RECT 1386.6000 42.3000 1399.8000 43.5000 ;
	    RECT 1400.7001 42.9000 1403.7001 44.1000 ;
	    RECT 1409.4000 42.9000 1414.2001 44.1000 ;
	    RECT 1246.2001 39.6000 1248.6000 40.8000 ;
	    RECT 1249.5000 40.2000 1250.7001 40.5000 ;
	    RECT 1249.5000 39.3000 1253.4000 40.2000 ;
	    RECT 1240.2001 33.3000 1241.7001 38.4000 ;
	    RECT 1244.4000 33.3000 1246.8000 38.7000 ;
	    RECT 1249.5000 33.3000 1251.0000 38.4000 ;
	    RECT 1252.2001 33.3000 1253.4000 39.3000 ;
	    RECT 1386.6000 33.3000 1387.8000 42.3000 ;
	    RECT 1390.2001 40.2000 1394.7001 41.4000 ;
	    RECT 1393.5000 39.3000 1394.7001 40.2000 ;
	    RECT 1402.5000 39.3000 1403.7001 42.9000 ;
	    RECT 1405.8000 41.4000 1407.0000 42.6000 ;
	    RECT 1413.6000 41.7000 1414.8000 42.0000 ;
	    RECT 1408.2001 40.8000 1414.8000 41.7000 ;
	    RECT 1408.2001 40.5000 1409.4000 40.8000 ;
	    RECT 1405.8000 40.2000 1407.0000 40.5000 ;
	    RECT 1417.8000 39.6000 1419.0000 43.8000 ;
	    RECT 1426.5000 42.9000 1432.2001 44.1000 ;
	    RECT 1426.5000 41.1000 1427.7001 42.9000 ;
	    RECT 1433.1000 42.0000 1434.0000 45.0000 ;
	    RECT 1408.2001 39.3000 1409.4000 39.6000 ;
	    RECT 1391.4000 33.3000 1392.6000 39.3000 ;
	    RECT 1393.5000 38.1000 1397.4000 39.3000 ;
	    RECT 1402.5000 38.4000 1409.4000 39.3000 ;
	    RECT 1410.6000 38.4000 1411.8000 39.6000 ;
	    RECT 1412.7001 38.4000 1413.0000 39.6000 ;
	    RECT 1417.5000 38.4000 1419.0000 39.6000 ;
	    RECT 1425.0000 40.2000 1427.7001 41.1000 ;
	    RECT 1432.2001 41.1000 1434.0000 42.0000 ;
	    RECT 1425.0000 39.3000 1426.2001 40.2000 ;
	    RECT 1396.2001 33.3000 1397.4000 38.1000 ;
	    RECT 1422.6000 38.1000 1426.2001 39.3000 ;
	    RECT 1398.6000 33.3000 1399.8000 37.5000 ;
	    RECT 1401.0000 33.3000 1402.2001 37.5000 ;
	    RECT 1403.4000 33.3000 1404.6000 37.5000 ;
	    RECT 1405.8000 33.3000 1407.0000 36.3000 ;
	    RECT 1408.2001 33.3000 1409.4000 37.5000 ;
	    RECT 1410.6000 33.3000 1411.8000 36.3000 ;
	    RECT 1413.0000 33.3000 1414.2001 37.5000 ;
	    RECT 1415.4000 33.3000 1416.6000 37.5000 ;
	    RECT 1417.8000 33.3000 1419.0000 37.5000 ;
	    RECT 1420.2001 33.3000 1421.4000 37.5000 ;
	    RECT 1422.6000 33.3000 1423.8000 38.1000 ;
	    RECT 1427.4000 33.3000 1428.6000 39.3000 ;
	    RECT 1432.2001 33.3000 1433.4000 41.1000 ;
	    RECT 1434.9000 40.2000 1436.1000 46.8000 ;
	    RECT 1458.6000 46.8000 1459.5000 47.7000 ;
	    RECT 1458.6000 45.6000 1460.4000 46.8000 ;
	    RECT 1453.8000 45.4500 1455.0000 45.6000 ;
	    RECT 1456.2001 45.4500 1457.4000 45.6000 ;
	    RECT 1453.8000 44.5500 1457.4000 45.4500 ;
	    RECT 1453.8000 44.4000 1455.0000 44.5500 ;
	    RECT 1456.2001 44.4000 1457.4000 44.5500 ;
	    RECT 1456.2001 43.2000 1457.4000 43.5000 ;
	    RECT 1458.6000 41.1000 1459.5000 45.6000 ;
	    RECT 1461.3000 44.4000 1462.2001 47.7000 ;
	    RECT 1487.4000 47.4000 1488.6000 48.6000 ;
	    RECT 1494.6000 48.4500 1495.8000 48.6000 ;
	    RECT 1511.4000 48.4500 1512.6000 48.6000 ;
	    RECT 1494.6000 47.5500 1512.6000 48.4500 ;
	    RECT 1494.6000 47.4000 1495.8000 47.5500 ;
	    RECT 1511.4000 47.4000 1512.6000 47.5500 ;
	    RECT 1513.8000 47.4000 1515.0000 48.6000 ;
	    RECT 1516.2001 46.5000 1517.4000 59.7000 ;
	    RECT 1518.6000 53.7000 1519.8000 59.7000 ;
	    RECT 1525.8000 59.4000 1527.0000 60.6000 ;
	    RECT 1537.8000 47.7000 1539.0000 59.7000 ;
	    RECT 1540.2001 49.5000 1541.4000 59.7000 ;
	    RECT 1542.6000 48.6000 1543.8000 59.7000 ;
	    RECT 1554.6000 53.7000 1555.8000 59.7000 ;
	    RECT 1540.5000 47.7000 1543.8000 48.6000 ;
	    RECT 1487.4000 46.2000 1488.6000 46.5000 ;
	    RECT 1489.8000 44.4000 1491.0000 45.6000 ;
	    RECT 1491.9000 44.4000 1492.2001 45.6000 ;
	    RECT 1461.0000 43.5000 1462.2001 44.4000 ;
	    RECT 1494.6000 42.6000 1495.5000 46.5000 ;
	    RECT 1516.2001 45.4500 1517.4000 45.6000 ;
	    RECT 1530.6000 45.4500 1531.8000 45.6000 ;
	    RECT 1516.2001 44.5500 1531.8000 45.4500 ;
	    RECT 1516.2001 44.4000 1517.4000 44.5500 ;
	    RECT 1530.6000 44.4000 1531.8000 44.5500 ;
	    RECT 1537.8000 44.4000 1538.7001 47.7000 ;
	    RECT 1540.5000 46.8000 1541.4000 47.7000 ;
	    RECT 1539.6000 45.6000 1541.4000 46.8000 ;
	    RECT 1537.8000 43.5000 1539.0000 44.4000 ;
	    RECT 1493.1000 42.3000 1495.5000 42.6000 ;
	    RECT 1434.6000 39.0000 1436.1000 40.2000 ;
	    RECT 1456.2001 40.2000 1459.5000 41.1000 ;
	    RECT 1434.6000 33.3000 1435.8000 39.0000 ;
	    RECT 1437.0000 33.3000 1438.2001 36.3000 ;
	    RECT 1456.2001 33.3000 1457.4000 40.2000 ;
	    RECT 1458.6000 33.3000 1459.8000 39.3000 ;
	    RECT 1461.0000 33.3000 1462.2001 40.5000 ;
	    RECT 1487.4000 33.3000 1488.6000 42.3000 ;
	    RECT 1492.8000 41.7000 1495.5000 42.3000 ;
	    RECT 1492.8000 33.3000 1494.0000 41.7000 ;
	    RECT 1516.2001 39.3000 1517.4000 43.5000 ;
	    RECT 1518.6000 42.4500 1519.8000 42.6000 ;
	    RECT 1525.8000 42.4500 1527.0000 42.6000 ;
	    RECT 1518.6000 41.5500 1527.0000 42.4500 ;
	    RECT 1518.6000 41.4000 1519.8000 41.5500 ;
	    RECT 1525.8000 41.4000 1527.0000 41.5500 ;
	    RECT 1540.5000 41.1000 1541.4000 45.6000 ;
	    RECT 1542.6000 45.4500 1543.8000 45.6000 ;
	    RECT 1552.2001 45.4500 1553.4000 45.6000 ;
	    RECT 1542.6000 44.5500 1553.4000 45.4500 ;
	    RECT 1542.6000 44.4000 1543.8000 44.5500 ;
	    RECT 1552.2001 44.4000 1553.4000 44.5500 ;
	    RECT 1557.0000 43.5000 1558.2001 59.7000 ;
	    RECT 1542.6000 43.2000 1543.8000 43.5000 ;
	    RECT 1557.0000 41.4000 1558.2001 42.6000 ;
	    RECT 1518.6000 40.2000 1519.8000 40.5000 ;
	    RECT 1514.7001 38.4000 1517.4000 39.3000 ;
	    RECT 1514.7001 33.3000 1515.9000 38.4000 ;
	    RECT 1518.6000 33.3000 1519.8000 39.3000 ;
	    RECT 1537.8000 33.3000 1539.0000 40.5000 ;
	    RECT 1540.5000 40.2000 1543.8000 41.1000 ;
	    RECT 1540.2001 33.3000 1541.4000 39.3000 ;
	    RECT 1542.6000 33.3000 1543.8000 40.2000 ;
	    RECT 1554.6000 38.4000 1555.8000 39.6000 ;
	    RECT 1554.6000 37.2000 1555.8000 37.5000 ;
	    RECT 1554.6000 33.3000 1555.8000 36.3000 ;
	    RECT 1557.0000 33.3000 1558.2001 40.5000 ;
	    RECT 1.2000 30.6000 1569.0000 32.4000 ;
	    RECT 124.2000 26.7000 125.4000 29.7000 ;
	    RECT 126.6000 24.0000 127.8000 29.7000 ;
	    RECT 126.3000 22.8000 127.8000 24.0000 ;
	    RECT 126.3000 16.2000 127.5000 22.8000 ;
	    RECT 129.0000 21.9000 130.2000 29.7000 ;
	    RECT 133.8000 23.7000 135.0000 29.7000 ;
	    RECT 138.6000 24.9000 139.8000 29.7000 ;
	    RECT 141.0000 25.5000 142.2000 29.7000 ;
	    RECT 143.4000 25.5000 144.6000 29.7000 ;
	    RECT 145.8000 25.5000 147.0000 29.7000 ;
	    RECT 148.2000 25.5000 149.4000 29.7000 ;
	    RECT 150.6000 26.7000 151.8000 29.7000 ;
	    RECT 153.0000 25.5000 154.2000 29.7000 ;
	    RECT 155.4000 26.7000 156.6000 29.7000 ;
	    RECT 157.8000 25.5000 159.0000 29.7000 ;
	    RECT 160.2000 25.5000 161.4000 29.7000 ;
	    RECT 162.6000 25.5000 163.8000 29.7000 ;
	    RECT 136.2000 23.7000 139.8000 24.9000 ;
	    RECT 165.0000 24.9000 166.2000 29.7000 ;
	    RECT 136.2000 22.8000 137.4000 23.7000 ;
	    RECT 128.4000 21.0000 130.2000 21.9000 ;
	    RECT 134.7000 21.9000 137.4000 22.8000 ;
	    RECT 143.4000 23.4000 144.9000 24.6000 ;
	    RECT 149.4000 23.4000 149.7000 24.6000 ;
	    RECT 150.6000 23.4000 151.8000 24.6000 ;
	    RECT 153.0000 23.7000 159.9000 24.6000 ;
	    RECT 165.0000 23.7000 168.9000 24.9000 ;
	    RECT 169.8000 23.7000 171.0000 29.7000 ;
	    RECT 153.0000 23.4000 154.2000 23.7000 ;
	    RECT 128.4000 18.0000 129.3000 21.0000 ;
	    RECT 134.7000 20.1000 135.9000 21.9000 ;
	    RECT 130.2000 18.9000 135.9000 20.1000 ;
	    RECT 143.4000 19.2000 144.6000 23.4000 ;
	    RECT 155.4000 22.5000 156.6000 22.8000 ;
	    RECT 153.0000 22.2000 154.2000 22.5000 ;
	    RECT 147.6000 21.3000 154.2000 22.2000 ;
	    RECT 147.6000 21.0000 148.8000 21.3000 ;
	    RECT 155.4000 20.4000 156.6000 21.6000 ;
	    RECT 158.7000 20.1000 159.9000 23.7000 ;
	    RECT 167.7000 22.8000 168.9000 23.7000 ;
	    RECT 167.7000 21.6000 172.2000 22.8000 ;
	    RECT 174.6000 20.7000 175.8000 29.7000 ;
	    RECT 306.6000 26.7000 307.8000 29.7000 ;
	    RECT 309.0000 24.0000 310.2000 29.7000 ;
	    RECT 148.2000 18.9000 153.0000 20.1000 ;
	    RECT 158.7000 18.9000 161.7000 20.1000 ;
	    RECT 162.6000 19.5000 175.8000 20.7000 ;
	    RECT 138.6000 18.0000 139.8000 18.9000 ;
	    RECT 128.4000 17.1000 129.6000 18.0000 ;
	    RECT 138.6000 17.1000 164.1000 18.0000 ;
	    RECT 165.0000 17.4000 166.2000 18.6000 ;
	    RECT 172.5000 18.0000 173.7000 18.3000 ;
	    RECT 167.1000 17.1000 173.7000 18.0000 ;
	    RECT 126.3000 15.0000 127.8000 16.2000 ;
	    RECT 126.6000 13.5000 127.8000 15.0000 ;
	    RECT 128.7000 14.4000 129.6000 17.1000 ;
	    RECT 130.5000 16.2000 131.7000 16.5000 ;
	    RECT 130.5000 15.3000 168.9000 16.2000 ;
	    RECT 164.7000 15.0000 165.9000 15.3000 ;
	    RECT 169.8000 14.4000 171.0000 15.6000 ;
	    RECT 128.7000 13.5000 142.2000 14.4000 ;
	    RECT 73.8000 12.4500 75.0000 12.6000 ;
	    RECT 126.6000 12.4500 127.8000 12.6000 ;
	    RECT 73.8000 11.5500 127.8000 12.4500 ;
	    RECT 73.8000 11.4000 75.0000 11.5500 ;
	    RECT 126.6000 11.4000 127.8000 11.5500 ;
	    RECT 128.7000 11.1000 129.6000 13.5000 ;
	    RECT 141.0000 13.2000 142.2000 13.5000 ;
	    RECT 145.8000 13.5000 158.7000 14.4000 ;
	    RECT 145.8000 13.2000 147.0000 13.5000 ;
	    RECT 133.5000 11.4000 137.4000 12.6000 ;
	    RECT 124.2000 3.3000 125.4000 9.3000 ;
	    RECT 126.6000 3.3000 127.8000 10.5000 ;
	    RECT 128.7000 10.2000 132.6000 11.1000 ;
	    RECT 129.0000 3.3000 130.2000 9.3000 ;
	    RECT 131.4000 3.3000 132.6000 10.2000 ;
	    RECT 133.8000 3.3000 135.0000 9.3000 ;
	    RECT 136.2000 3.3000 137.4000 11.4000 ;
	    RECT 138.3000 10.2000 144.6000 11.4000 ;
	    RECT 138.6000 3.3000 139.8000 9.3000 ;
	    RECT 141.0000 3.3000 142.2000 7.5000 ;
	    RECT 143.4000 3.3000 144.6000 7.5000 ;
	    RECT 145.8000 3.3000 147.0000 7.5000 ;
	    RECT 148.2000 3.3000 149.4000 12.6000 ;
	    RECT 153.0000 11.4000 156.9000 12.6000 ;
	    RECT 157.8000 12.3000 158.7000 13.5000 ;
	    RECT 160.2000 14.1000 161.4000 14.4000 ;
	    RECT 160.2000 13.5000 168.3000 14.1000 ;
	    RECT 160.2000 13.2000 169.5000 13.5000 ;
	    RECT 167.4000 12.3000 169.5000 13.2000 ;
	    RECT 157.8000 11.4000 166.5000 12.3000 ;
	    RECT 171.0000 12.0000 173.4000 13.2000 ;
	    RECT 171.0000 11.4000 171.9000 12.0000 ;
	    RECT 150.6000 3.3000 151.8000 9.3000 ;
	    RECT 153.0000 3.3000 154.2000 10.5000 ;
	    RECT 155.4000 3.3000 156.6000 9.3000 ;
	    RECT 157.8000 3.3000 159.0000 10.5000 ;
	    RECT 165.6000 10.2000 171.9000 11.4000 ;
	    RECT 174.6000 11.1000 175.8000 19.5000 ;
	    RECT 308.7000 22.8000 310.2000 24.0000 ;
	    RECT 308.7000 16.2000 309.9000 22.8000 ;
	    RECT 311.4000 21.9000 312.6000 29.7000 ;
	    RECT 316.2000 23.7000 317.4000 29.7000 ;
	    RECT 321.0000 24.9000 322.2000 29.7000 ;
	    RECT 323.4000 25.5000 324.6000 29.7000 ;
	    RECT 325.8000 25.5000 327.0000 29.7000 ;
	    RECT 328.2000 25.5000 329.4000 29.7000 ;
	    RECT 330.6000 25.5000 331.8000 29.7000 ;
	    RECT 333.0000 26.7000 334.2000 29.7000 ;
	    RECT 335.4000 25.5000 336.6000 29.7000 ;
	    RECT 337.8000 26.7000 339.0000 29.7000 ;
	    RECT 340.2000 25.5000 341.4000 29.7000 ;
	    RECT 342.6000 25.5000 343.8000 29.7000 ;
	    RECT 345.0000 25.5000 346.2000 29.7000 ;
	    RECT 318.6000 23.7000 322.2000 24.9000 ;
	    RECT 347.4000 24.9000 348.6000 29.7000 ;
	    RECT 318.6000 22.8000 319.8000 23.7000 ;
	    RECT 310.8000 21.0000 312.6000 21.9000 ;
	    RECT 317.1000 21.9000 319.8000 22.8000 ;
	    RECT 325.8000 23.4000 327.3000 24.6000 ;
	    RECT 331.8000 23.4000 332.1000 24.6000 ;
	    RECT 333.0000 23.4000 334.2000 24.6000 ;
	    RECT 335.4000 23.7000 342.3000 24.6000 ;
	    RECT 347.4000 23.7000 351.3000 24.9000 ;
	    RECT 352.2000 23.7000 353.4000 29.7000 ;
	    RECT 335.4000 23.4000 336.6000 23.7000 ;
	    RECT 310.8000 18.0000 311.7000 21.0000 ;
	    RECT 317.1000 20.1000 318.3000 21.9000 ;
	    RECT 312.6000 18.9000 318.3000 20.1000 ;
	    RECT 325.8000 19.2000 327.0000 23.4000 ;
	    RECT 337.8000 22.5000 339.0000 22.8000 ;
	    RECT 335.4000 22.2000 336.6000 22.5000 ;
	    RECT 330.0000 21.3000 336.6000 22.2000 ;
	    RECT 330.0000 21.0000 331.2000 21.3000 ;
	    RECT 337.8000 20.4000 339.0000 21.6000 ;
	    RECT 341.1000 20.1000 342.3000 23.7000 ;
	    RECT 350.1000 22.8000 351.3000 23.7000 ;
	    RECT 350.1000 21.6000 354.6000 22.8000 ;
	    RECT 357.0000 20.7000 358.2000 29.7000 ;
	    RECT 489.0000 26.7000 490.2000 29.7000 ;
	    RECT 491.4000 24.0000 492.6000 29.7000 ;
	    RECT 330.6000 18.9000 335.4000 20.1000 ;
	    RECT 341.1000 18.9000 344.1000 20.1000 ;
	    RECT 345.0000 19.5000 358.2000 20.7000 ;
	    RECT 321.0000 18.0000 322.2000 18.9000 ;
	    RECT 310.8000 17.1000 312.0000 18.0000 ;
	    RECT 321.0000 17.1000 346.5000 18.0000 ;
	    RECT 347.4000 17.4000 348.6000 18.6000 ;
	    RECT 354.9000 18.0000 356.1000 18.3000 ;
	    RECT 349.5000 17.1000 356.1000 18.0000 ;
	    RECT 308.7000 15.0000 310.2000 16.2000 ;
	    RECT 309.0000 13.5000 310.2000 15.0000 ;
	    RECT 311.1000 14.4000 312.0000 17.1000 ;
	    RECT 312.9000 16.2000 314.1000 16.5000 ;
	    RECT 312.9000 15.3000 351.3000 16.2000 ;
	    RECT 347.1000 15.0000 348.3000 15.3000 ;
	    RECT 352.2000 14.4000 353.4000 15.6000 ;
	    RECT 311.1000 13.5000 324.6000 14.4000 ;
	    RECT 256.2000 12.4500 257.4000 12.6000 ;
	    RECT 309.0000 12.4500 310.2000 12.6000 ;
	    RECT 256.2000 11.5500 310.2000 12.4500 ;
	    RECT 256.2000 11.4000 257.4000 11.5500 ;
	    RECT 309.0000 11.4000 310.2000 11.5500 ;
	    RECT 172.8000 10.2000 175.8000 11.1000 ;
	    RECT 311.1000 11.1000 312.0000 13.5000 ;
	    RECT 323.4000 13.2000 324.6000 13.5000 ;
	    RECT 328.2000 13.5000 341.1000 14.4000 ;
	    RECT 328.2000 13.2000 329.4000 13.5000 ;
	    RECT 315.9000 11.4000 319.8000 12.6000 ;
	    RECT 160.2000 3.3000 161.4000 7.5000 ;
	    RECT 162.6000 3.3000 163.8000 7.5000 ;
	    RECT 165.0000 3.3000 166.2000 9.3000 ;
	    RECT 167.4000 3.3000 168.6000 10.2000 ;
	    RECT 172.8000 9.3000 173.7000 10.2000 ;
	    RECT 169.8000 2.4000 171.0000 9.3000 ;
	    RECT 172.2000 8.4000 173.7000 9.3000 ;
	    RECT 172.2000 3.3000 173.4000 8.4000 ;
	    RECT 174.6000 3.3000 175.8000 9.3000 ;
	    RECT 306.6000 3.3000 307.8000 9.3000 ;
	    RECT 309.0000 3.3000 310.2000 10.5000 ;
	    RECT 311.1000 10.2000 315.0000 11.1000 ;
	    RECT 311.4000 3.3000 312.6000 9.3000 ;
	    RECT 313.8000 3.3000 315.0000 10.2000 ;
	    RECT 316.2000 3.3000 317.4000 9.3000 ;
	    RECT 318.6000 3.3000 319.8000 11.4000 ;
	    RECT 320.7000 10.2000 327.0000 11.4000 ;
	    RECT 321.0000 3.3000 322.2000 9.3000 ;
	    RECT 323.4000 3.3000 324.6000 7.5000 ;
	    RECT 325.8000 3.3000 327.0000 7.5000 ;
	    RECT 328.2000 3.3000 329.4000 7.5000 ;
	    RECT 330.6000 3.3000 331.8000 12.6000 ;
	    RECT 335.4000 11.4000 339.3000 12.6000 ;
	    RECT 340.2000 12.3000 341.1000 13.5000 ;
	    RECT 342.6000 14.1000 343.8000 14.4000 ;
	    RECT 342.6000 13.5000 350.7000 14.1000 ;
	    RECT 342.6000 13.2000 351.9000 13.5000 ;
	    RECT 349.8000 12.3000 351.9000 13.2000 ;
	    RECT 340.2000 11.4000 348.9000 12.3000 ;
	    RECT 353.4000 12.0000 355.8000 13.2000 ;
	    RECT 353.4000 11.4000 354.3000 12.0000 ;
	    RECT 333.0000 3.3000 334.2000 9.3000 ;
	    RECT 335.4000 3.3000 336.6000 10.5000 ;
	    RECT 337.8000 3.3000 339.0000 9.3000 ;
	    RECT 340.2000 3.3000 341.4000 10.5000 ;
	    RECT 348.0000 10.2000 354.3000 11.4000 ;
	    RECT 357.0000 11.1000 358.2000 19.5000 ;
	    RECT 491.1000 22.8000 492.6000 24.0000 ;
	    RECT 491.1000 16.2000 492.3000 22.8000 ;
	    RECT 493.8000 21.9000 495.0000 29.7000 ;
	    RECT 498.6000 23.7000 499.8000 29.7000 ;
	    RECT 503.4000 24.9000 504.6000 29.7000 ;
	    RECT 505.8000 25.5000 507.0000 29.7000 ;
	    RECT 508.2000 25.5000 509.4000 29.7000 ;
	    RECT 510.6000 25.5000 511.8000 29.7000 ;
	    RECT 513.0000 25.5000 514.2000 29.7000 ;
	    RECT 515.4000 26.7000 516.6000 29.7000 ;
	    RECT 517.8000 25.5000 519.0000 29.7000 ;
	    RECT 520.2000 26.7000 521.4000 29.7000 ;
	    RECT 522.6000 25.5000 523.8000 29.7000 ;
	    RECT 525.0000 25.5000 526.2000 29.7000 ;
	    RECT 527.4000 25.5000 528.6000 29.7000 ;
	    RECT 501.0000 23.7000 504.6000 24.9000 ;
	    RECT 529.8000 24.9000 531.0000 29.7000 ;
	    RECT 501.0000 22.8000 502.2000 23.7000 ;
	    RECT 493.2000 21.0000 495.0000 21.9000 ;
	    RECT 499.5000 21.9000 502.2000 22.8000 ;
	    RECT 508.2000 23.4000 509.7000 24.6000 ;
	    RECT 514.2000 23.4000 514.5000 24.6000 ;
	    RECT 515.4000 23.4000 516.6000 24.6000 ;
	    RECT 517.8000 23.7000 524.7000 24.6000 ;
	    RECT 529.8000 23.7000 533.7000 24.9000 ;
	    RECT 534.6000 23.7000 535.8000 29.7000 ;
	    RECT 517.8000 23.4000 519.0000 23.7000 ;
	    RECT 493.2000 18.0000 494.1000 21.0000 ;
	    RECT 499.5000 20.1000 500.7000 21.9000 ;
	    RECT 495.0000 18.9000 500.7000 20.1000 ;
	    RECT 508.2000 19.2000 509.4000 23.4000 ;
	    RECT 520.2000 22.5000 521.4000 22.8000 ;
	    RECT 517.8000 22.2000 519.0000 22.5000 ;
	    RECT 512.4000 21.3000 519.0000 22.2000 ;
	    RECT 512.4000 21.0000 513.6000 21.3000 ;
	    RECT 520.2000 20.4000 521.4000 21.6000 ;
	    RECT 523.5000 20.1000 524.7000 23.7000 ;
	    RECT 532.5000 22.8000 533.7000 23.7000 ;
	    RECT 532.5000 21.6000 537.0000 22.8000 ;
	    RECT 539.4000 20.7000 540.6000 29.7000 ;
	    RECT 559.5000 24.6000 560.7000 29.7000 ;
	    RECT 559.5000 23.7000 562.2000 24.6000 ;
	    RECT 563.4000 23.7000 564.6000 29.7000 ;
	    RECT 577.8000 26.7000 579.0000 29.7000 ;
	    RECT 577.8000 25.5000 579.0000 25.8000 ;
	    RECT 513.0000 18.9000 517.8000 20.1000 ;
	    RECT 523.5000 18.9000 526.5000 20.1000 ;
	    RECT 527.4000 19.5000 540.6000 20.7000 ;
	    RECT 561.0000 19.5000 562.2000 23.7000 ;
	    RECT 577.8000 23.4000 579.0000 24.6000 ;
	    RECT 563.4000 22.5000 564.6000 22.8000 ;
	    RECT 580.2000 22.5000 581.4000 29.7000 ;
	    RECT 594.6000 26.7000 595.8000 29.7000 ;
	    RECT 594.6000 25.5000 595.8000 25.8000 ;
	    RECT 585.0000 24.4500 586.2000 24.6000 ;
	    RECT 594.6000 24.4500 595.8000 24.6000 ;
	    RECT 585.0000 23.5500 595.8000 24.4500 ;
	    RECT 585.0000 23.4000 586.2000 23.5500 ;
	    RECT 594.6000 23.4000 595.8000 23.5500 ;
	    RECT 597.0000 22.5000 598.2000 29.7000 ;
	    RECT 563.4000 20.4000 564.6000 21.6000 ;
	    RECT 580.2000 21.4500 581.4000 21.6000 ;
	    RECT 594.6000 21.4500 595.8000 21.6000 ;
	    RECT 580.2000 20.5500 595.8000 21.4500 ;
	    RECT 580.2000 20.4000 581.4000 20.5500 ;
	    RECT 594.6000 20.4000 595.8000 20.5500 ;
	    RECT 597.0000 21.4500 598.2000 21.6000 ;
	    RECT 726.6000 21.4500 727.8000 21.6000 ;
	    RECT 597.0000 20.5500 727.8000 21.4500 ;
	    RECT 597.0000 20.4000 598.2000 20.5500 ;
	    RECT 726.6000 20.4000 727.8000 20.5500 ;
	    RECT 729.0000 20.7000 730.2000 29.7000 ;
	    RECT 733.8000 23.7000 735.0000 29.7000 ;
	    RECT 738.6000 24.9000 739.8000 29.7000 ;
	    RECT 741.0000 25.5000 742.2000 29.7000 ;
	    RECT 743.4000 25.5000 744.6000 29.7000 ;
	    RECT 745.8000 25.5000 747.0000 29.7000 ;
	    RECT 748.2000 26.7000 749.4000 29.7000 ;
	    RECT 750.6000 25.5000 751.8000 29.7000 ;
	    RECT 753.0000 26.7000 754.2000 29.7000 ;
	    RECT 755.4000 25.5000 756.6000 29.7000 ;
	    RECT 757.8000 25.5000 759.0000 29.7000 ;
	    RECT 760.2000 25.5000 761.4000 29.7000 ;
	    RECT 762.6000 25.5000 763.8000 29.7000 ;
	    RECT 735.9000 23.7000 739.8000 24.9000 ;
	    RECT 765.0000 24.9000 766.2000 29.7000 ;
	    RECT 744.9000 23.7000 751.8000 24.6000 ;
	    RECT 735.9000 22.8000 737.1000 23.7000 ;
	    RECT 732.6000 21.6000 737.1000 22.8000 ;
	    RECT 729.0000 19.5000 742.2000 20.7000 ;
	    RECT 744.9000 20.1000 746.1000 23.7000 ;
	    RECT 750.6000 23.4000 751.8000 23.7000 ;
	    RECT 753.0000 23.4000 754.2000 24.6000 ;
	    RECT 755.1000 23.4000 755.4000 24.6000 ;
	    RECT 759.9000 23.4000 761.4000 24.6000 ;
	    RECT 765.0000 23.7000 768.6000 24.9000 ;
	    RECT 769.8000 23.7000 771.0000 29.7000 ;
	    RECT 748.2000 22.5000 749.4000 22.8000 ;
	    RECT 750.6000 22.2000 751.8000 22.5000 ;
	    RECT 748.2000 20.4000 749.4000 21.6000 ;
	    RECT 750.6000 21.3000 757.2000 22.2000 ;
	    RECT 756.0000 21.0000 757.2000 21.3000 ;
	    RECT 503.4000 18.0000 504.6000 18.9000 ;
	    RECT 493.2000 17.1000 494.4000 18.0000 ;
	    RECT 503.4000 17.1000 528.9000 18.0000 ;
	    RECT 529.8000 17.4000 531.0000 18.6000 ;
	    RECT 537.3000 18.0000 538.5000 18.3000 ;
	    RECT 531.9000 17.1000 538.5000 18.0000 ;
	    RECT 491.1000 15.0000 492.6000 16.2000 ;
	    RECT 491.4000 13.5000 492.6000 15.0000 ;
	    RECT 493.5000 14.4000 494.4000 17.1000 ;
	    RECT 495.3000 16.2000 496.5000 16.5000 ;
	    RECT 495.3000 15.3000 533.7000 16.2000 ;
	    RECT 529.5000 15.0000 530.7000 15.3000 ;
	    RECT 534.6000 14.4000 535.8000 15.6000 ;
	    RECT 493.5000 13.5000 507.0000 14.4000 ;
	    RECT 424.2000 12.4500 425.4000 12.6000 ;
	    RECT 491.4000 12.4500 492.6000 12.6000 ;
	    RECT 424.2000 11.5500 492.6000 12.4500 ;
	    RECT 424.2000 11.4000 425.4000 11.5500 ;
	    RECT 491.4000 11.4000 492.6000 11.5500 ;
	    RECT 355.2000 10.2000 358.2000 11.1000 ;
	    RECT 493.5000 11.1000 494.4000 13.5000 ;
	    RECT 505.8000 13.2000 507.0000 13.5000 ;
	    RECT 510.6000 13.5000 523.5000 14.4000 ;
	    RECT 510.6000 13.2000 511.8000 13.5000 ;
	    RECT 498.3000 11.4000 502.2000 12.6000 ;
	    RECT 342.6000 3.3000 343.8000 7.5000 ;
	    RECT 345.0000 3.3000 346.2000 7.5000 ;
	    RECT 347.4000 3.3000 348.6000 9.3000 ;
	    RECT 349.8000 3.3000 351.0000 10.2000 ;
	    RECT 355.2000 9.3000 356.1000 10.2000 ;
	    RECT 352.2000 2.4000 353.4000 9.3000 ;
	    RECT 354.6000 8.4000 356.1000 9.3000 ;
	    RECT 354.6000 3.3000 355.8000 8.4000 ;
	    RECT 357.0000 3.3000 358.2000 9.3000 ;
	    RECT 489.0000 3.3000 490.2000 9.3000 ;
	    RECT 491.4000 3.3000 492.6000 10.5000 ;
	    RECT 493.5000 10.2000 497.4000 11.1000 ;
	    RECT 493.8000 3.3000 495.0000 9.3000 ;
	    RECT 496.2000 3.3000 497.4000 10.2000 ;
	    RECT 498.6000 3.3000 499.8000 9.3000 ;
	    RECT 501.0000 3.3000 502.2000 11.4000 ;
	    RECT 503.1000 10.2000 509.4000 11.4000 ;
	    RECT 503.4000 3.3000 504.6000 9.3000 ;
	    RECT 505.8000 3.3000 507.0000 7.5000 ;
	    RECT 508.2000 3.3000 509.4000 7.5000 ;
	    RECT 510.6000 3.3000 511.8000 7.5000 ;
	    RECT 513.0000 3.3000 514.2000 12.6000 ;
	    RECT 517.8000 11.4000 521.7000 12.6000 ;
	    RECT 522.6000 12.3000 523.5000 13.5000 ;
	    RECT 525.0000 14.1000 526.2000 14.4000 ;
	    RECT 525.0000 13.5000 533.1000 14.1000 ;
	    RECT 525.0000 13.2000 534.3000 13.5000 ;
	    RECT 532.2000 12.3000 534.3000 13.2000 ;
	    RECT 522.6000 11.4000 531.3000 12.3000 ;
	    RECT 535.8000 12.0000 538.2000 13.2000 ;
	    RECT 535.8000 11.4000 536.7000 12.0000 ;
	    RECT 515.4000 3.3000 516.6000 9.3000 ;
	    RECT 517.8000 3.3000 519.0000 10.5000 ;
	    RECT 520.2000 3.3000 521.4000 9.3000 ;
	    RECT 522.6000 3.3000 523.8000 10.5000 ;
	    RECT 530.4000 10.2000 536.7000 11.4000 ;
	    RECT 539.4000 11.1000 540.6000 19.5000 ;
	    RECT 541.8000 18.4500 543.0000 18.6000 ;
	    RECT 561.0000 18.4500 562.2000 18.6000 ;
	    RECT 541.8000 17.5500 562.2000 18.4500 ;
	    RECT 541.8000 17.4000 543.0000 17.5500 ;
	    RECT 561.0000 17.4000 562.2000 17.5500 ;
	    RECT 558.6000 14.4000 559.8000 15.6000 ;
	    RECT 558.6000 13.2000 559.8000 13.5000 ;
	    RECT 537.6000 10.2000 540.6000 11.1000 ;
	    RECT 525.0000 3.3000 526.2000 7.5000 ;
	    RECT 527.4000 3.3000 528.6000 7.5000 ;
	    RECT 529.8000 3.3000 531.0000 9.3000 ;
	    RECT 532.2000 3.3000 533.4000 10.2000 ;
	    RECT 537.6000 9.3000 538.5000 10.2000 ;
	    RECT 534.6000 2.4000 535.8000 9.3000 ;
	    RECT 537.0000 8.4000 538.5000 9.3000 ;
	    RECT 537.0000 3.3000 538.2000 8.4000 ;
	    RECT 539.4000 3.3000 540.6000 9.3000 ;
	    RECT 558.6000 3.3000 559.8000 9.3000 ;
	    RECT 561.0000 3.3000 562.2000 16.5000 ;
	    RECT 563.4000 3.3000 564.6000 9.3000 ;
	    RECT 577.8000 3.3000 579.0000 9.3000 ;
	    RECT 580.2000 3.3000 581.4000 19.5000 ;
	    RECT 594.6000 3.3000 595.8000 9.3000 ;
	    RECT 597.0000 3.3000 598.2000 19.5000 ;
	    RECT 729.0000 11.1000 730.2000 19.5000 ;
	    RECT 743.1000 18.9000 746.1000 20.1000 ;
	    RECT 751.8000 18.9000 756.6000 20.1000 ;
	    RECT 760.2000 19.2000 761.4000 23.4000 ;
	    RECT 767.4000 22.8000 768.6000 23.7000 ;
	    RECT 767.4000 21.9000 770.1000 22.8000 ;
	    RECT 768.9000 20.1000 770.1000 21.9000 ;
	    RECT 774.6000 21.9000 775.8000 29.7000 ;
	    RECT 777.0000 24.0000 778.2000 29.7000 ;
	    RECT 779.4000 26.7000 780.6000 29.7000 ;
	    RECT 777.0000 22.8000 778.5000 24.0000 ;
	    RECT 774.6000 21.0000 776.4000 21.9000 ;
	    RECT 768.9000 18.9000 774.6000 20.1000 ;
	    RECT 731.1000 18.0000 732.3000 18.3000 ;
	    RECT 731.1000 17.1000 737.7000 18.0000 ;
	    RECT 738.6000 17.4000 739.8000 18.6000 ;
	    RECT 765.0000 18.0000 766.2000 18.9000 ;
	    RECT 775.5000 18.0000 776.4000 21.0000 ;
	    RECT 740.7000 17.1000 766.2000 18.0000 ;
	    RECT 775.2000 17.1000 776.4000 18.0000 ;
	    RECT 773.1000 16.2000 774.3000 16.5000 ;
	    RECT 733.8000 14.4000 735.0000 15.6000 ;
	    RECT 735.9000 15.3000 774.3000 16.2000 ;
	    RECT 738.9000 15.0000 740.1000 15.3000 ;
	    RECT 775.2000 14.4000 776.1000 17.1000 ;
	    RECT 777.3000 16.2000 778.5000 22.8000 ;
	    RECT 793.8000 22.5000 795.0000 29.7000 ;
	    RECT 796.2000 26.7000 797.4000 29.7000 ;
	    RECT 796.2000 25.5000 797.4000 25.8000 ;
	    RECT 796.2000 24.4500 797.4000 24.6000 ;
	    RECT 796.2000 23.5500 814.0500 24.4500 ;
	    RECT 815.4000 23.7000 816.6000 29.7000 ;
	    RECT 819.3000 24.6000 820.5000 29.7000 ;
	    RECT 817.8000 23.7000 820.5000 24.6000 ;
	    RECT 839.4000 23.7000 840.6000 29.7000 ;
	    RECT 843.3000 24.6000 844.5000 29.7000 ;
	    RECT 856.2000 26.7000 857.4000 29.7000 ;
	    RECT 856.2000 25.5000 857.4000 25.8000 ;
	    RECT 841.8000 23.7000 844.5000 24.6000 ;
	    RECT 796.2000 23.4000 797.4000 23.5500 ;
	    RECT 793.8000 21.4500 795.0000 21.6000 ;
	    RECT 798.6000 21.4500 799.8000 21.6000 ;
	    RECT 793.8000 20.5500 799.8000 21.4500 ;
	    RECT 813.1500 21.4500 814.0500 23.5500 ;
	    RECT 815.4000 22.5000 816.6000 22.8000 ;
	    RECT 815.4000 21.4500 816.6000 21.6000 ;
	    RECT 813.1500 20.5500 816.6000 21.4500 ;
	    RECT 793.8000 20.4000 795.0000 20.5500 ;
	    RECT 798.6000 20.4000 799.8000 20.5500 ;
	    RECT 815.4000 20.4000 816.6000 20.5500 ;
	    RECT 817.8000 19.5000 819.0000 23.7000 ;
	    RECT 839.4000 22.5000 840.6000 22.8000 ;
	    RECT 839.4000 20.4000 840.6000 21.6000 ;
	    RECT 841.8000 19.5000 843.0000 23.7000 ;
	    RECT 856.2000 23.4000 857.4000 24.6000 ;
	    RECT 858.6000 22.5000 859.8000 29.7000 ;
	    RECT 885.0000 24.0000 886.2000 29.7000 ;
	    RECT 887.4000 24.9000 888.6000 29.7000 ;
	    RECT 889.8000 24.0000 891.0000 29.7000 ;
	    RECT 885.0000 23.7000 891.0000 24.0000 ;
	    RECT 892.2000 23.7000 893.4000 29.7000 ;
	    RECT 885.3000 23.1000 890.7000 23.7000 ;
	    RECT 892.2000 22.5000 893.1000 23.7000 ;
	    RECT 858.6000 21.4500 859.8000 21.6000 ;
	    RECT 858.6000 20.5500 883.6500 21.4500 ;
	    RECT 858.6000 20.4000 859.8000 20.5500 ;
	    RECT 743.4000 14.1000 744.6000 14.4000 ;
	    RECT 736.5000 13.5000 744.6000 14.1000 ;
	    RECT 735.3000 13.2000 744.6000 13.5000 ;
	    RECT 746.1000 13.5000 759.0000 14.4000 ;
	    RECT 731.4000 12.0000 733.8000 13.2000 ;
	    RECT 735.3000 12.3000 737.4000 13.2000 ;
	    RECT 746.1000 12.3000 747.0000 13.5000 ;
	    RECT 757.8000 13.2000 759.0000 13.5000 ;
	    RECT 762.6000 13.5000 776.1000 14.4000 ;
	    RECT 777.0000 15.0000 778.5000 16.2000 ;
	    RECT 777.0000 13.5000 778.2000 15.0000 ;
	    RECT 762.6000 13.2000 763.8000 13.5000 ;
	    RECT 732.9000 11.4000 733.8000 12.0000 ;
	    RECT 738.3000 11.4000 747.0000 12.3000 ;
	    RECT 747.9000 11.4000 751.8000 12.6000 ;
	    RECT 729.0000 10.2000 732.0000 11.1000 ;
	    RECT 732.9000 10.2000 739.2000 11.4000 ;
	    RECT 731.1000 9.3000 732.0000 10.2000 ;
	    RECT 729.0000 3.3000 730.2000 9.3000 ;
	    RECT 731.1000 8.4000 732.6000 9.3000 ;
	    RECT 731.4000 3.3000 732.6000 8.4000 ;
	    RECT 733.8000 2.4000 735.0000 9.3000 ;
	    RECT 736.2000 3.3000 737.4000 10.2000 ;
	    RECT 738.6000 3.3000 739.8000 9.3000 ;
	    RECT 741.0000 3.3000 742.2000 7.5000 ;
	    RECT 743.4000 3.3000 744.6000 7.5000 ;
	    RECT 745.8000 3.3000 747.0000 10.5000 ;
	    RECT 748.2000 3.3000 749.4000 9.3000 ;
	    RECT 750.6000 3.3000 751.8000 10.5000 ;
	    RECT 753.0000 3.3000 754.2000 9.3000 ;
	    RECT 755.4000 3.3000 756.6000 12.6000 ;
	    RECT 767.4000 11.4000 771.3000 12.6000 ;
	    RECT 760.2000 10.2000 766.5000 11.4000 ;
	    RECT 757.8000 3.3000 759.0000 7.5000 ;
	    RECT 760.2000 3.3000 761.4000 7.5000 ;
	    RECT 762.6000 3.3000 763.8000 7.5000 ;
	    RECT 765.0000 3.3000 766.2000 9.3000 ;
	    RECT 767.4000 3.3000 768.6000 11.4000 ;
	    RECT 775.2000 11.1000 776.1000 13.5000 ;
	    RECT 777.0000 11.4000 778.2000 12.6000 ;
	    RECT 772.2000 10.2000 776.1000 11.1000 ;
	    RECT 769.8000 3.3000 771.0000 9.3000 ;
	    RECT 772.2000 3.3000 773.4000 10.2000 ;
	    RECT 774.6000 3.3000 775.8000 9.3000 ;
	    RECT 777.0000 3.3000 778.2000 10.5000 ;
	    RECT 779.4000 3.3000 780.6000 9.3000 ;
	    RECT 793.8000 3.3000 795.0000 19.5000 ;
	    RECT 801.0000 18.4500 802.2000 18.6000 ;
	    RECT 817.8000 18.4500 819.0000 18.6000 ;
	    RECT 801.0000 17.5500 819.0000 18.4500 ;
	    RECT 801.0000 17.4000 802.2000 17.5500 ;
	    RECT 817.8000 17.4000 819.0000 17.5500 ;
	    RECT 841.8000 18.4500 843.0000 18.6000 ;
	    RECT 856.2000 18.4500 857.4000 18.6000 ;
	    RECT 841.8000 17.5500 857.4000 18.4500 ;
	    RECT 841.8000 17.4000 843.0000 17.5500 ;
	    RECT 856.2000 17.4000 857.4000 17.5500 ;
	    RECT 796.2000 3.3000 797.4000 9.3000 ;
	    RECT 815.4000 3.3000 816.6000 9.3000 ;
	    RECT 817.8000 3.3000 819.0000 16.5000 ;
	    RECT 820.2000 15.4500 821.4000 15.6000 ;
	    RECT 829.8000 15.4500 831.0000 15.6000 ;
	    RECT 820.2000 14.5500 831.0000 15.4500 ;
	    RECT 820.2000 14.4000 821.4000 14.5500 ;
	    RECT 829.8000 14.4000 831.0000 14.5500 ;
	    RECT 820.2000 13.2000 821.4000 13.5000 ;
	    RECT 820.2000 3.3000 821.4000 9.3000 ;
	    RECT 839.4000 3.3000 840.6000 9.3000 ;
	    RECT 841.8000 3.3000 843.0000 16.5000 ;
	    RECT 844.2000 13.2000 845.4000 13.5000 ;
	    RECT 844.2000 3.3000 845.4000 9.3000 ;
	    RECT 856.2000 3.3000 857.4000 9.3000 ;
	    RECT 858.6000 3.3000 859.8000 19.5000 ;
	    RECT 882.7500 18.4500 883.6500 20.5500 ;
	    RECT 885.0000 20.4000 886.2000 21.6000 ;
	    RECT 887.1000 20.7000 887.4000 22.2000 ;
	    RECT 889.5000 20.4000 891.3000 21.6000 ;
	    RECT 892.2000 21.4500 893.4000 21.6000 ;
	    RECT 964.2000 21.4500 965.4000 21.6000 ;
	    RECT 892.2000 20.5500 965.4000 21.4500 ;
	    RECT 892.2000 20.4000 893.4000 20.5500 ;
	    RECT 964.2000 20.4000 965.4000 20.5500 ;
	    RECT 1024.2001 20.7000 1025.4000 29.7000 ;
	    RECT 1029.0000 23.7000 1030.2001 29.7000 ;
	    RECT 1033.8000 24.9000 1035.0000 29.7000 ;
	    RECT 1036.2001 25.5000 1037.4000 29.7000 ;
	    RECT 1038.6000 25.5000 1039.8000 29.7000 ;
	    RECT 1041.0000 25.5000 1042.2001 29.7000 ;
	    RECT 1043.4000 26.7000 1044.6000 29.7000 ;
	    RECT 1045.8000 25.5000 1047.0000 29.7000 ;
	    RECT 1048.2001 26.7000 1049.4000 29.7000 ;
	    RECT 1050.6000 25.5000 1051.8000 29.7000 ;
	    RECT 1053.0000 25.5000 1054.2001 29.7000 ;
	    RECT 1055.4000 25.5000 1056.6000 29.7000 ;
	    RECT 1057.8000 25.5000 1059.0000 29.7000 ;
	    RECT 1031.1000 23.7000 1035.0000 24.9000 ;
	    RECT 1060.2001 24.9000 1061.4000 29.7000 ;
	    RECT 1040.1000 23.7000 1047.0000 24.6000 ;
	    RECT 1031.1000 22.8000 1032.3000 23.7000 ;
	    RECT 1027.8000 21.6000 1032.3000 22.8000 ;
	    RECT 887.4000 19.5000 888.6000 19.8000 ;
	    RECT 887.4000 18.4500 888.6000 18.6000 ;
	    RECT 882.7500 17.5500 888.6000 18.4500 ;
	    RECT 887.4000 17.4000 888.6000 17.5500 ;
	    RECT 889.5000 15.3000 890.4000 20.4000 ;
	    RECT 1024.2001 19.5000 1037.4000 20.7000 ;
	    RECT 1040.1000 20.1000 1041.3000 23.7000 ;
	    RECT 1045.8000 23.4000 1047.0000 23.7000 ;
	    RECT 1048.2001 23.4000 1049.4000 24.6000 ;
	    RECT 1050.3000 23.4000 1050.6000 24.6000 ;
	    RECT 1055.1000 23.4000 1056.6000 24.6000 ;
	    RECT 1060.2001 23.7000 1063.8000 24.9000 ;
	    RECT 1065.0000 23.7000 1066.2001 29.7000 ;
	    RECT 1043.4000 22.5000 1044.6000 22.8000 ;
	    RECT 1045.8000 22.2000 1047.0000 22.5000 ;
	    RECT 1043.4000 20.4000 1044.6000 21.6000 ;
	    RECT 1045.8000 21.3000 1052.4000 22.2000 ;
	    RECT 1051.2001 21.0000 1052.4000 21.3000 ;
	    RECT 885.0000 3.3000 886.2000 15.3000 ;
	    RECT 888.9000 14.4000 890.4000 15.3000 ;
	    RECT 892.2000 14.4000 893.4000 15.6000 ;
	    RECT 888.9000 3.3000 890.1000 14.4000 ;
	    RECT 891.3000 12.6000 892.2000 13.5000 ;
	    RECT 891.0000 11.4000 892.2000 12.6000 ;
	    RECT 1024.2001 11.1000 1025.4000 19.5000 ;
	    RECT 1038.3000 18.9000 1041.3000 20.1000 ;
	    RECT 1047.0000 18.9000 1051.8000 20.1000 ;
	    RECT 1055.4000 19.2000 1056.6000 23.4000 ;
	    RECT 1062.6000 22.8000 1063.8000 23.7000 ;
	    RECT 1062.6000 21.9000 1065.3000 22.8000 ;
	    RECT 1064.1000 20.1000 1065.3000 21.9000 ;
	    RECT 1069.8000 21.9000 1071.0000 29.7000 ;
	    RECT 1072.2001 24.0000 1073.4000 29.7000 ;
	    RECT 1074.6000 26.7000 1075.8000 29.7000 ;
	    RECT 1072.2001 22.8000 1073.7001 24.0000 ;
	    RECT 1069.8000 21.0000 1071.6000 21.9000 ;
	    RECT 1064.1000 18.9000 1069.8000 20.1000 ;
	    RECT 1026.3000 18.0000 1027.5000 18.3000 ;
	    RECT 1026.3000 17.1000 1032.9000 18.0000 ;
	    RECT 1033.8000 17.4000 1035.0000 18.6000 ;
	    RECT 1060.2001 18.0000 1061.4000 18.9000 ;
	    RECT 1070.7001 18.0000 1071.6000 21.0000 ;
	    RECT 1035.9000 17.1000 1061.4000 18.0000 ;
	    RECT 1070.4000 17.1000 1071.6000 18.0000 ;
	    RECT 1068.3000 16.2000 1069.5000 16.5000 ;
	    RECT 1026.6000 15.4500 1027.8000 15.6000 ;
	    RECT 1029.0000 15.4500 1030.2001 15.6000 ;
	    RECT 1026.6000 14.5500 1030.2001 15.4500 ;
	    RECT 1031.1000 15.3000 1069.5000 16.2000 ;
	    RECT 1034.1000 15.0000 1035.3000 15.3000 ;
	    RECT 1026.6000 14.4000 1027.8000 14.5500 ;
	    RECT 1029.0000 14.4000 1030.2001 14.5500 ;
	    RECT 1070.4000 14.4000 1071.3000 17.1000 ;
	    RECT 1072.5000 16.2000 1073.7001 22.8000 ;
	    RECT 1038.6000 14.1000 1039.8000 14.4000 ;
	    RECT 1031.7001 13.5000 1039.8000 14.1000 ;
	    RECT 1030.5000 13.2000 1039.8000 13.5000 ;
	    RECT 1041.3000 13.5000 1054.2001 14.4000 ;
	    RECT 1026.6000 12.0000 1029.0000 13.2000 ;
	    RECT 1030.5000 12.3000 1032.6000 13.2000 ;
	    RECT 1041.3000 12.3000 1042.2001 13.5000 ;
	    RECT 1053.0000 13.2000 1054.2001 13.5000 ;
	    RECT 1057.8000 13.5000 1071.3000 14.4000 ;
	    RECT 1072.2001 15.0000 1073.7001 16.2000 ;
	    RECT 1206.6000 20.7000 1207.8000 29.7000 ;
	    RECT 1211.4000 23.7000 1212.6000 29.7000 ;
	    RECT 1216.2001 24.9000 1217.4000 29.7000 ;
	    RECT 1218.6000 25.5000 1219.8000 29.7000 ;
	    RECT 1221.0000 25.5000 1222.2001 29.7000 ;
	    RECT 1223.4000 25.5000 1224.6000 29.7000 ;
	    RECT 1225.8000 26.7000 1227.0000 29.7000 ;
	    RECT 1228.2001 25.5000 1229.4000 29.7000 ;
	    RECT 1230.6000 26.7000 1231.8000 29.7000 ;
	    RECT 1233.0000 25.5000 1234.2001 29.7000 ;
	    RECT 1235.4000 25.5000 1236.6000 29.7000 ;
	    RECT 1237.8000 25.5000 1239.0000 29.7000 ;
	    RECT 1240.2001 25.5000 1241.4000 29.7000 ;
	    RECT 1213.5000 23.7000 1217.4000 24.9000 ;
	    RECT 1242.6000 24.9000 1243.8000 29.7000 ;
	    RECT 1222.5000 23.7000 1229.4000 24.6000 ;
	    RECT 1213.5000 22.8000 1214.7001 23.7000 ;
	    RECT 1210.2001 21.6000 1214.7001 22.8000 ;
	    RECT 1206.6000 19.5000 1219.8000 20.7000 ;
	    RECT 1222.5000 20.1000 1223.7001 23.7000 ;
	    RECT 1228.2001 23.4000 1229.4000 23.7000 ;
	    RECT 1230.6000 23.4000 1231.8000 24.6000 ;
	    RECT 1232.7001 23.4000 1233.0000 24.6000 ;
	    RECT 1237.5000 23.4000 1239.0000 24.6000 ;
	    RECT 1242.6000 23.7000 1246.2001 24.9000 ;
	    RECT 1247.4000 23.7000 1248.6000 29.7000 ;
	    RECT 1225.8000 22.5000 1227.0000 22.8000 ;
	    RECT 1228.2001 22.2000 1229.4000 22.5000 ;
	    RECT 1225.8000 20.4000 1227.0000 21.6000 ;
	    RECT 1228.2001 21.3000 1234.8000 22.2000 ;
	    RECT 1233.6000 21.0000 1234.8000 21.3000 ;
	    RECT 1072.2001 13.5000 1073.4000 15.0000 ;
	    RECT 1057.8000 13.2000 1059.0000 13.5000 ;
	    RECT 1028.1000 11.4000 1029.0000 12.0000 ;
	    RECT 1033.5000 11.4000 1042.2001 12.3000 ;
	    RECT 1043.1000 11.4000 1047.0000 12.6000 ;
	    RECT 1024.2001 10.2000 1027.2001 11.1000 ;
	    RECT 1028.1000 10.2000 1034.4000 11.4000 ;
	    RECT 1026.3000 9.3000 1027.2001 10.2000 ;
	    RECT 891.3000 3.3000 892.5000 9.3000 ;
	    RECT 1024.2001 3.3000 1025.4000 9.3000 ;
	    RECT 1026.3000 8.4000 1027.8000 9.3000 ;
	    RECT 1026.6000 3.3000 1027.8000 8.4000 ;
	    RECT 1029.0000 2.4000 1030.2001 9.3000 ;
	    RECT 1031.4000 3.3000 1032.6000 10.2000 ;
	    RECT 1033.8000 3.3000 1035.0000 9.3000 ;
	    RECT 1036.2001 3.3000 1037.4000 7.5000 ;
	    RECT 1038.6000 3.3000 1039.8000 7.5000 ;
	    RECT 1041.0000 3.3000 1042.2001 10.5000 ;
	    RECT 1043.4000 3.3000 1044.6000 9.3000 ;
	    RECT 1045.8000 3.3000 1047.0000 10.5000 ;
	    RECT 1048.2001 3.3000 1049.4000 9.3000 ;
	    RECT 1050.6000 3.3000 1051.8000 12.6000 ;
	    RECT 1062.6000 11.4000 1066.5000 12.6000 ;
	    RECT 1055.4000 10.2000 1061.7001 11.4000 ;
	    RECT 1053.0000 3.3000 1054.2001 7.5000 ;
	    RECT 1055.4000 3.3000 1056.6000 7.5000 ;
	    RECT 1057.8000 3.3000 1059.0000 7.5000 ;
	    RECT 1060.2001 3.3000 1061.4000 9.3000 ;
	    RECT 1062.6000 3.3000 1063.8000 11.4000 ;
	    RECT 1070.4000 11.1000 1071.3000 13.5000 ;
	    RECT 1072.2001 11.4000 1073.4000 12.6000 ;
	    RECT 1067.4000 10.2000 1071.3000 11.1000 ;
	    RECT 1206.6000 11.1000 1207.8000 19.5000 ;
	    RECT 1220.7001 18.9000 1223.7001 20.1000 ;
	    RECT 1229.4000 18.9000 1234.2001 20.1000 ;
	    RECT 1237.8000 19.2000 1239.0000 23.4000 ;
	    RECT 1245.0000 22.8000 1246.2001 23.7000 ;
	    RECT 1245.0000 21.9000 1247.7001 22.8000 ;
	    RECT 1246.5000 20.1000 1247.7001 21.9000 ;
	    RECT 1252.2001 21.9000 1253.4000 29.7000 ;
	    RECT 1254.6000 24.0000 1255.8000 29.7000 ;
	    RECT 1257.0000 26.7000 1258.2001 29.7000 ;
	    RECT 1271.4000 26.7000 1272.6000 29.7000 ;
	    RECT 1271.4000 25.5000 1272.6000 25.8000 ;
	    RECT 1254.6000 22.8000 1256.1000 24.0000 ;
	    RECT 1271.4000 23.4000 1272.6000 24.6000 ;
	    RECT 1252.2001 21.0000 1254.0000 21.9000 ;
	    RECT 1246.5000 18.9000 1252.2001 20.1000 ;
	    RECT 1208.7001 18.0000 1209.9000 18.3000 ;
	    RECT 1208.7001 17.1000 1215.3000 18.0000 ;
	    RECT 1216.2001 17.4000 1217.4000 18.6000 ;
	    RECT 1242.6000 18.0000 1243.8000 18.9000 ;
	    RECT 1253.1000 18.0000 1254.0000 21.0000 ;
	    RECT 1218.3000 17.1000 1243.8000 18.0000 ;
	    RECT 1252.8000 17.1000 1254.0000 18.0000 ;
	    RECT 1250.7001 16.2000 1251.9000 16.5000 ;
	    RECT 1211.4000 14.4000 1212.6000 15.6000 ;
	    RECT 1213.5000 15.3000 1251.9000 16.2000 ;
	    RECT 1216.5000 15.0000 1217.7001 15.3000 ;
	    RECT 1252.8000 14.4000 1253.7001 17.1000 ;
	    RECT 1254.9000 16.2000 1256.1000 22.8000 ;
	    RECT 1273.8000 22.5000 1275.0000 29.7000 ;
	    RECT 1297.8000 23.7000 1299.0000 29.7000 ;
	    RECT 1300.2001 24.0000 1301.4000 29.7000 ;
	    RECT 1302.6000 24.9000 1303.8000 29.7000 ;
	    RECT 1305.0000 24.0000 1306.2001 29.7000 ;
	    RECT 1324.2001 26.7000 1325.4000 29.7000 ;
	    RECT 1326.6000 26.7000 1327.8000 29.7000 ;
	    RECT 1329.0000 26.7000 1330.2001 29.7000 ;
	    RECT 1300.2001 23.7000 1306.2001 24.0000 ;
	    RECT 1298.1000 22.5000 1299.0000 23.7000 ;
	    RECT 1300.5000 23.1000 1305.9000 23.7000 ;
	    RECT 1326.6000 22.5000 1327.5000 26.7000 ;
	    RECT 1329.0000 25.5000 1330.2001 25.8000 ;
	    RECT 1329.0000 23.4000 1330.2001 24.6000 ;
	    RECT 1273.8000 21.4500 1275.0000 21.6000 ;
	    RECT 1276.2001 21.4500 1277.4000 21.6000 ;
	    RECT 1273.8000 20.5500 1277.4000 21.4500 ;
	    RECT 1273.8000 20.4000 1275.0000 20.5500 ;
	    RECT 1276.2001 20.4000 1277.4000 20.5500 ;
	    RECT 1278.6000 21.4500 1279.8000 21.6000 ;
	    RECT 1297.8000 21.4500 1299.0000 21.6000 ;
	    RECT 1278.6000 20.5500 1299.0000 21.4500 ;
	    RECT 1278.6000 20.4000 1279.8000 20.5500 ;
	    RECT 1297.8000 20.4000 1299.0000 20.5500 ;
	    RECT 1299.9000 20.4000 1301.7001 21.6000 ;
	    RECT 1303.8000 20.7000 1304.1000 22.2000 ;
	    RECT 1305.0000 20.4000 1306.2001 21.6000 ;
	    RECT 1307.4000 21.4500 1308.6000 21.6000 ;
	    RECT 1326.6000 21.4500 1327.8000 21.6000 ;
	    RECT 1307.4000 20.5500 1327.8000 21.4500 ;
	    RECT 1307.4000 20.4000 1308.6000 20.5500 ;
	    RECT 1326.6000 20.4000 1327.8000 20.5500 ;
	    RECT 1461.0000 20.7000 1462.2001 29.7000 ;
	    RECT 1465.8000 23.7000 1467.0000 29.7000 ;
	    RECT 1470.6000 24.9000 1471.8000 29.7000 ;
	    RECT 1473.0000 25.5000 1474.2001 29.7000 ;
	    RECT 1475.4000 25.5000 1476.6000 29.7000 ;
	    RECT 1477.8000 25.5000 1479.0000 29.7000 ;
	    RECT 1480.2001 26.7000 1481.4000 29.7000 ;
	    RECT 1482.6000 25.5000 1483.8000 29.7000 ;
	    RECT 1485.0000 26.7000 1486.2001 29.7000 ;
	    RECT 1487.4000 25.5000 1488.6000 29.7000 ;
	    RECT 1489.8000 25.5000 1491.0000 29.7000 ;
	    RECT 1492.2001 25.5000 1493.4000 29.7000 ;
	    RECT 1494.6000 25.5000 1495.8000 29.7000 ;
	    RECT 1467.9000 23.7000 1471.8000 24.9000 ;
	    RECT 1497.0000 24.9000 1498.2001 29.7000 ;
	    RECT 1476.9000 23.7000 1483.8000 24.6000 ;
	    RECT 1467.9000 22.8000 1469.1000 23.7000 ;
	    RECT 1464.6000 21.6000 1469.1000 22.8000 ;
	    RECT 1221.0000 14.1000 1222.2001 14.4000 ;
	    RECT 1214.1000 13.5000 1222.2001 14.1000 ;
	    RECT 1212.9000 13.2000 1222.2001 13.5000 ;
	    RECT 1223.7001 13.5000 1236.6000 14.4000 ;
	    RECT 1209.0000 12.0000 1211.4000 13.2000 ;
	    RECT 1212.9000 12.3000 1215.0000 13.2000 ;
	    RECT 1223.7001 12.3000 1224.6000 13.5000 ;
	    RECT 1235.4000 13.2000 1236.6000 13.5000 ;
	    RECT 1240.2001 13.5000 1253.7001 14.4000 ;
	    RECT 1254.6000 15.0000 1256.1000 16.2000 ;
	    RECT 1254.6000 13.5000 1255.8000 15.0000 ;
	    RECT 1240.2001 13.2000 1241.4000 13.5000 ;
	    RECT 1210.5000 11.4000 1211.4000 12.0000 ;
	    RECT 1215.9000 11.4000 1224.6000 12.3000 ;
	    RECT 1225.5000 11.4000 1229.4000 12.6000 ;
	    RECT 1065.0000 3.3000 1066.2001 9.3000 ;
	    RECT 1067.4000 3.3000 1068.6000 10.2000 ;
	    RECT 1069.8000 3.3000 1071.0000 9.3000 ;
	    RECT 1072.2001 3.3000 1073.4000 10.5000 ;
	    RECT 1206.6000 10.2000 1209.6000 11.1000 ;
	    RECT 1210.5000 10.2000 1216.8000 11.4000 ;
	    RECT 1208.7001 9.3000 1209.6000 10.2000 ;
	    RECT 1074.6000 3.3000 1075.8000 9.3000 ;
	    RECT 1206.6000 3.3000 1207.8000 9.3000 ;
	    RECT 1208.7001 8.4000 1210.2001 9.3000 ;
	    RECT 1209.0000 3.3000 1210.2001 8.4000 ;
	    RECT 1211.4000 2.4000 1212.6000 9.3000 ;
	    RECT 1213.8000 3.3000 1215.0000 10.2000 ;
	    RECT 1216.2001 3.3000 1217.4000 9.3000 ;
	    RECT 1218.6000 3.3000 1219.8000 7.5000 ;
	    RECT 1221.0000 3.3000 1222.2001 7.5000 ;
	    RECT 1223.4000 3.3000 1224.6000 10.5000 ;
	    RECT 1225.8000 3.3000 1227.0000 9.3000 ;
	    RECT 1228.2001 3.3000 1229.4000 10.5000 ;
	    RECT 1230.6000 3.3000 1231.8000 9.3000 ;
	    RECT 1233.0000 3.3000 1234.2001 12.6000 ;
	    RECT 1245.0000 11.4000 1248.9000 12.6000 ;
	    RECT 1237.8000 10.2000 1244.1000 11.4000 ;
	    RECT 1235.4000 3.3000 1236.6000 7.5000 ;
	    RECT 1237.8000 3.3000 1239.0000 7.5000 ;
	    RECT 1240.2001 3.3000 1241.4000 7.5000 ;
	    RECT 1242.6000 3.3000 1243.8000 9.3000 ;
	    RECT 1245.0000 3.3000 1246.2001 11.4000 ;
	    RECT 1252.8000 11.1000 1253.7001 13.5000 ;
	    RECT 1254.6000 11.4000 1255.8000 12.6000 ;
	    RECT 1249.8000 10.2000 1253.7001 11.1000 ;
	    RECT 1247.4000 3.3000 1248.6000 9.3000 ;
	    RECT 1249.8000 3.3000 1251.0000 10.2000 ;
	    RECT 1252.2001 3.3000 1253.4000 9.3000 ;
	    RECT 1254.6000 3.3000 1255.8000 10.5000 ;
	    RECT 1257.0000 3.3000 1258.2001 9.3000 ;
	    RECT 1271.4000 3.3000 1272.6000 9.3000 ;
	    RECT 1273.8000 3.3000 1275.0000 19.5000 ;
	    RECT 1297.8000 14.4000 1299.0000 15.6000 ;
	    RECT 1300.8000 15.3000 1301.7001 20.4000 ;
	    RECT 1302.6000 19.5000 1303.8000 19.8000 ;
	    RECT 1461.0000 19.5000 1474.2001 20.7000 ;
	    RECT 1476.9000 20.1000 1478.1000 23.7000 ;
	    RECT 1482.6000 23.4000 1483.8000 23.7000 ;
	    RECT 1485.0000 23.4000 1486.2001 24.6000 ;
	    RECT 1487.1000 23.4000 1487.4000 24.6000 ;
	    RECT 1491.9000 23.4000 1493.4000 24.6000 ;
	    RECT 1497.0000 23.7000 1500.6000 24.9000 ;
	    RECT 1501.8000 23.7000 1503.0000 29.7000 ;
	    RECT 1480.2001 22.5000 1481.4000 22.8000 ;
	    RECT 1482.6000 22.2000 1483.8000 22.5000 ;
	    RECT 1480.2001 20.4000 1481.4000 21.6000 ;
	    RECT 1482.6000 21.3000 1489.2001 22.2000 ;
	    RECT 1488.0000 21.0000 1489.2001 21.3000 ;
	    RECT 1302.6000 18.4500 1303.8000 18.6000 ;
	    RECT 1324.2001 18.4500 1325.4000 18.6000 ;
	    RECT 1302.6000 17.5500 1325.4000 18.4500 ;
	    RECT 1302.6000 17.4000 1303.8000 17.5500 ;
	    RECT 1324.2001 17.4000 1325.4000 17.5500 ;
	    RECT 1324.2001 16.2000 1325.4000 16.5000 ;
	    RECT 1326.6000 15.3000 1327.5000 19.5000 ;
	    RECT 1300.8000 14.4000 1302.3000 15.3000 ;
	    RECT 1299.0000 12.6000 1299.9000 13.5000 ;
	    RECT 1299.0000 11.4000 1300.2001 12.6000 ;
	    RECT 1298.7001 3.3000 1299.9000 9.3000 ;
	    RECT 1301.1000 3.3000 1302.3000 14.4000 ;
	    RECT 1305.0000 3.3000 1306.2001 15.3000 ;
	    RECT 1325.1000 14.1000 1327.8000 15.3000 ;
	    RECT 1325.1000 3.3000 1326.3000 14.1000 ;
	    RECT 1329.0000 3.3000 1330.2001 15.3000 ;
	    RECT 1461.0000 11.1000 1462.2001 19.5000 ;
	    RECT 1475.1000 18.9000 1478.1000 20.1000 ;
	    RECT 1483.8000 18.9000 1488.6000 20.1000 ;
	    RECT 1492.2001 19.2000 1493.4000 23.4000 ;
	    RECT 1499.4000 22.8000 1500.6000 23.7000 ;
	    RECT 1499.4000 21.9000 1502.1000 22.8000 ;
	    RECT 1500.9000 20.1000 1502.1000 21.9000 ;
	    RECT 1506.6000 21.9000 1507.8000 29.7000 ;
	    RECT 1509.0000 24.0000 1510.2001 29.7000 ;
	    RECT 1511.4000 26.7000 1512.6000 29.7000 ;
	    RECT 1509.0000 22.8000 1510.5000 24.0000 ;
	    RECT 1535.4000 23.7000 1536.6000 29.7000 ;
	    RECT 1537.8000 24.0000 1539.0000 29.7000 ;
	    RECT 1540.2001 24.9000 1541.4000 29.7000 ;
	    RECT 1542.6000 24.0000 1543.8000 29.7000 ;
	    RECT 1557.0000 26.7000 1558.2001 29.7000 ;
	    RECT 1557.0000 25.5000 1558.2001 25.8000 ;
	    RECT 1537.8000 23.7000 1543.8000 24.0000 ;
	    RECT 1552.2001 24.4500 1553.4000 24.6000 ;
	    RECT 1557.0000 24.4500 1558.2001 24.6000 ;
	    RECT 1506.6000 21.0000 1508.4000 21.9000 ;
	    RECT 1500.9000 18.9000 1506.6000 20.1000 ;
	    RECT 1463.1000 18.0000 1464.3000 18.3000 ;
	    RECT 1463.1000 17.1000 1469.7001 18.0000 ;
	    RECT 1470.6000 17.4000 1471.8000 18.6000 ;
	    RECT 1497.0000 18.0000 1498.2001 18.9000 ;
	    RECT 1507.5000 18.0000 1508.4000 21.0000 ;
	    RECT 1472.7001 17.1000 1498.2001 18.0000 ;
	    RECT 1507.2001 17.1000 1508.4000 18.0000 ;
	    RECT 1505.1000 16.2000 1506.3000 16.5000 ;
	    RECT 1465.8000 14.4000 1467.0000 15.6000 ;
	    RECT 1467.9000 15.3000 1506.3000 16.2000 ;
	    RECT 1470.9000 15.0000 1472.1000 15.3000 ;
	    RECT 1507.2001 14.4000 1508.1000 17.1000 ;
	    RECT 1509.3000 16.2000 1510.5000 22.8000 ;
	    RECT 1535.7001 22.5000 1536.6000 23.7000 ;
	    RECT 1538.1000 23.1000 1543.5000 23.7000 ;
	    RECT 1552.2001 23.5500 1558.2001 24.4500 ;
	    RECT 1552.2001 23.4000 1553.4000 23.5500 ;
	    RECT 1557.0000 23.4000 1558.2001 23.5500 ;
	    RECT 1559.4000 22.5000 1560.6000 29.7000 ;
	    RECT 1511.4000 21.4500 1512.6000 21.6000 ;
	    RECT 1535.4000 21.4500 1536.6000 21.6000 ;
	    RECT 1511.4000 20.5500 1536.6000 21.4500 ;
	    RECT 1511.4000 20.4000 1512.6000 20.5500 ;
	    RECT 1535.4000 20.4000 1536.6000 20.5500 ;
	    RECT 1537.5000 20.4000 1539.3000 21.6000 ;
	    RECT 1541.4000 20.7000 1541.7001 22.2000 ;
	    RECT 1542.6000 20.4000 1543.8000 21.6000 ;
	    RECT 1559.4000 21.4500 1560.6000 21.6000 ;
	    RECT 1545.1500 20.5500 1560.6000 21.4500 ;
	    RECT 1475.4000 14.1000 1476.6000 14.4000 ;
	    RECT 1468.5000 13.5000 1476.6000 14.1000 ;
	    RECT 1467.3000 13.2000 1476.6000 13.5000 ;
	    RECT 1478.1000 13.5000 1491.0000 14.4000 ;
	    RECT 1463.4000 12.0000 1465.8000 13.2000 ;
	    RECT 1467.3000 12.3000 1469.4000 13.2000 ;
	    RECT 1478.1000 12.3000 1479.0000 13.5000 ;
	    RECT 1489.8000 13.2000 1491.0000 13.5000 ;
	    RECT 1494.6000 13.5000 1508.1000 14.4000 ;
	    RECT 1509.0000 15.0000 1510.5000 16.2000 ;
	    RECT 1530.6000 15.4500 1531.8000 15.6000 ;
	    RECT 1535.4000 15.4500 1536.6000 15.6000 ;
	    RECT 1509.0000 13.5000 1510.2001 15.0000 ;
	    RECT 1530.6000 14.5500 1536.6000 15.4500 ;
	    RECT 1530.6000 14.4000 1531.8000 14.5500 ;
	    RECT 1535.4000 14.4000 1536.6000 14.5500 ;
	    RECT 1538.4000 15.3000 1539.3000 20.4000 ;
	    RECT 1540.2001 19.5000 1541.4000 19.8000 ;
	    RECT 1540.2001 18.4500 1541.4000 18.6000 ;
	    RECT 1545.1500 18.4500 1546.0500 20.5500 ;
	    RECT 1559.4000 20.4000 1560.6000 20.5500 ;
	    RECT 1540.2001 17.5500 1546.0500 18.4500 ;
	    RECT 1540.2001 17.4000 1541.4000 17.5500 ;
	    RECT 1538.4000 14.4000 1539.9000 15.3000 ;
	    RECT 1494.6000 13.2000 1495.8000 13.5000 ;
	    RECT 1464.9000 11.4000 1465.8000 12.0000 ;
	    RECT 1470.3000 11.4000 1479.0000 12.3000 ;
	    RECT 1479.9000 11.4000 1483.8000 12.6000 ;
	    RECT 1461.0000 10.2000 1464.0000 11.1000 ;
	    RECT 1464.9000 10.2000 1471.2001 11.4000 ;
	    RECT 1463.1000 9.3000 1464.0000 10.2000 ;
	    RECT 1461.0000 3.3000 1462.2001 9.3000 ;
	    RECT 1463.1000 8.4000 1464.6000 9.3000 ;
	    RECT 1463.4000 3.3000 1464.6000 8.4000 ;
	    RECT 1465.8000 2.4000 1467.0000 9.3000 ;
	    RECT 1468.2001 3.3000 1469.4000 10.2000 ;
	    RECT 1470.6000 3.3000 1471.8000 9.3000 ;
	    RECT 1473.0000 3.3000 1474.2001 7.5000 ;
	    RECT 1475.4000 3.3000 1476.6000 7.5000 ;
	    RECT 1477.8000 3.3000 1479.0000 10.5000 ;
	    RECT 1480.2001 3.3000 1481.4000 9.3000 ;
	    RECT 1482.6000 3.3000 1483.8000 10.5000 ;
	    RECT 1485.0000 3.3000 1486.2001 9.3000 ;
	    RECT 1487.4000 3.3000 1488.6000 12.6000 ;
	    RECT 1499.4000 11.4000 1503.3000 12.6000 ;
	    RECT 1492.2001 10.2000 1498.5000 11.4000 ;
	    RECT 1489.8000 3.3000 1491.0000 7.5000 ;
	    RECT 1492.2001 3.3000 1493.4000 7.5000 ;
	    RECT 1494.6000 3.3000 1495.8000 7.5000 ;
	    RECT 1497.0000 3.3000 1498.2001 9.3000 ;
	    RECT 1499.4000 3.3000 1500.6000 11.4000 ;
	    RECT 1507.2001 11.1000 1508.1000 13.5000 ;
	    RECT 1536.6000 12.6000 1537.5000 13.5000 ;
	    RECT 1509.0000 12.4500 1510.2001 12.6000 ;
	    RECT 1516.2001 12.4500 1517.4000 12.6000 ;
	    RECT 1509.0000 11.5500 1517.4000 12.4500 ;
	    RECT 1509.0000 11.4000 1510.2001 11.5500 ;
	    RECT 1516.2001 11.4000 1517.4000 11.5500 ;
	    RECT 1536.6000 11.4000 1537.8000 12.6000 ;
	    RECT 1504.2001 10.2000 1508.1000 11.1000 ;
	    RECT 1501.8000 3.3000 1503.0000 9.3000 ;
	    RECT 1504.2001 3.3000 1505.4000 10.2000 ;
	    RECT 1506.6000 3.3000 1507.8000 9.3000 ;
	    RECT 1509.0000 3.3000 1510.2001 10.5000 ;
	    RECT 1511.4000 3.3000 1512.6000 9.3000 ;
	    RECT 1536.3000 3.3000 1537.5000 9.3000 ;
	    RECT 1538.7001 3.3000 1539.9000 14.4000 ;
	    RECT 1542.6000 3.3000 1543.8000 15.3000 ;
	    RECT 1557.0000 3.3000 1558.2001 9.3000 ;
	    RECT 1559.4000 3.3000 1560.6000 19.5000 ;
	    RECT 1566.6000 2.4000 1567.8000 3.6000 ;
	    RECT 1.2000 0.6000 1569.0000 2.4000 ;
         LAYER metal2 ;
	    RECT 136.2000 1457.4000 137.4000 1458.6000 ;
	    RECT 131.4000 1454.4000 132.6000 1455.6000 ;
	    RECT 131.5500 1446.6000 132.4500 1454.4000 ;
	    RECT 131.4000 1445.4000 132.6000 1446.6000 ;
	    RECT 138.6000 1446.3000 139.8000 1466.7001 ;
	    RECT 141.0000 1446.3000 142.2000 1466.7001 ;
	    RECT 143.4000 1449.3000 144.6000 1466.7001 ;
	    RECT 145.8000 1463.4000 147.0000 1464.6000 ;
	    RECT 145.9500 1461.6000 146.8500 1463.4000 ;
	    RECT 145.8000 1460.4000 147.0000 1461.6000 ;
	    RECT 148.2000 1449.3000 149.4000 1466.7001 ;
	    RECT 150.6000 1463.4000 151.8000 1464.6000 ;
	    RECT 150.7500 1446.4501 151.6500 1463.4000 ;
	    RECT 153.0000 1449.3000 154.2000 1466.7001 ;
	    RECT 148.3500 1445.5500 151.6500 1446.4501 ;
	    RECT 155.4000 1446.3000 156.6000 1466.7001 ;
	    RECT 157.8000 1446.3000 159.0000 1466.7001 ;
	    RECT 160.2000 1446.3000 161.4000 1466.7001 ;
	    RECT 177.0000 1463.4000 178.2000 1464.6000 ;
	    RECT 191.4000 1463.4000 192.6000 1464.6000 ;
	    RECT 225.0000 1463.4000 226.2000 1464.6000 ;
	    RECT 268.2000 1463.4000 269.4000 1464.6000 ;
	    RECT 165.0000 1457.4000 166.2000 1458.6000 ;
	    RECT 129.0000 1436.4000 130.2000 1437.6000 ;
	    RECT 129.1500 1428.6000 130.0500 1436.4000 ;
	    RECT 129.0000 1427.4000 130.2000 1428.6000 ;
	    RECT 133.8000 1427.4000 135.0000 1428.6000 ;
	    RECT 133.9500 1425.6000 134.8500 1427.4000 ;
	    RECT 133.8000 1424.4000 135.0000 1425.6000 ;
	    RECT 49.8000 1421.4000 51.0000 1422.6000 ;
	    RECT 23.4000 1379.4000 24.6000 1380.6000 ;
	    RECT 23.5500 1308.6000 24.4500 1379.4000 ;
	    RECT 23.4000 1307.4000 24.6000 1308.6000 ;
	    RECT 49.9500 1302.6000 50.8500 1421.4000 ;
	    RECT 126.6000 1391.4000 127.8000 1392.6000 ;
	    RECT 126.7500 1380.6000 127.6500 1391.4000 ;
	    RECT 126.6000 1379.4000 127.8000 1380.6000 ;
	    RECT 131.4000 1376.4000 132.6000 1377.6000 ;
	    RECT 76.2000 1373.4000 77.4000 1374.6000 ;
	    RECT 54.6000 1304.4000 55.8000 1305.6000 ;
	    RECT 18.6000 1301.4000 19.8000 1302.6000 ;
	    RECT 49.8000 1301.4000 51.0000 1302.6000 ;
	    RECT 18.7500 1281.6000 19.6500 1301.4000 ;
	    RECT 54.7500 1281.6000 55.6500 1304.4000 ;
	    RECT 76.3500 1284.6000 77.2500 1373.4000 ;
	    RECT 131.5500 1368.6000 132.4500 1376.4000 ;
	    RECT 131.4000 1367.4000 132.6000 1368.6000 ;
	    RECT 105.0000 1355.4000 106.2000 1356.6000 ;
	    RECT 78.6000 1325.4000 79.8000 1326.6000 ;
	    RECT 57.0000 1283.4000 58.2000 1284.6000 ;
	    RECT 76.2000 1283.4000 77.4000 1284.6000 ;
	    RECT 18.6000 1280.4000 19.8000 1281.6000 ;
	    RECT 33.0000 1280.4000 34.2000 1281.6000 ;
	    RECT 35.4000 1280.4000 36.6000 1281.6000 ;
	    RECT 54.6000 1280.4000 55.8000 1281.6000 ;
	    RECT 28.2000 1277.4000 29.4000 1278.6000 ;
	    RECT 33.1500 1248.6000 34.0500 1280.4000 ;
	    RECT 35.5500 1278.6000 36.4500 1280.4000 ;
	    RECT 35.4000 1277.4000 36.6000 1278.6000 ;
	    RECT 35.4000 1274.4000 36.6000 1275.6000 ;
	    RECT 35.5500 1272.6000 36.4500 1274.4000 ;
	    RECT 35.4000 1271.4000 36.6000 1272.6000 ;
	    RECT 47.4000 1271.4000 48.6000 1272.6000 ;
	    RECT 33.0000 1247.4000 34.2000 1248.6000 ;
	    RECT 23.4000 1187.4000 24.6000 1188.6000 ;
	    RECT 23.5500 1185.6000 24.4500 1187.4000 ;
	    RECT 23.4000 1185.4501 24.6000 1185.6000 ;
	    RECT 23.4000 1184.5500 26.8500 1185.4501 ;
	    RECT 23.4000 1184.4000 24.6000 1184.5500 ;
	    RECT 18.6000 1181.4000 19.8000 1182.6000 ;
	    RECT 13.8000 1163.4000 15.0000 1164.6000 ;
	    RECT 13.9500 1152.6000 14.8500 1163.4000 ;
	    RECT 13.8000 1151.4000 15.0000 1152.6000 ;
	    RECT 18.7500 1044.6000 19.6500 1181.4000 ;
	    RECT 23.4000 1133.4000 24.6000 1134.6000 ;
	    RECT 18.6000 1043.4000 19.8000 1044.6000 ;
	    RECT 18.7500 1041.6000 19.6500 1043.4000 ;
	    RECT 18.6000 1040.4000 19.8000 1041.6000 ;
	    RECT 23.5500 1035.6000 24.4500 1133.4000 ;
	    RECT 23.4000 1034.4000 24.6000 1035.6000 ;
	    RECT 25.9500 945.6000 26.8500 1184.5500 ;
	    RECT 33.0000 1181.4000 34.2000 1182.6000 ;
	    RECT 35.4000 983.4000 36.6000 984.6000 ;
	    RECT 33.0000 947.4000 34.2000 948.6000 ;
	    RECT 18.6000 944.4000 19.8000 945.6000 ;
	    RECT 25.8000 944.4000 27.0000 945.6000 ;
	    RECT 28.2000 944.4000 29.4000 945.6000 ;
	    RECT 18.7500 918.6000 19.6500 944.4000 ;
	    RECT 28.3500 942.6000 29.2500 944.4000 ;
	    RECT 25.8000 941.4000 27.0000 942.6000 ;
	    RECT 28.2000 941.4000 29.4000 942.6000 ;
	    RECT 25.9500 921.6000 26.8500 941.4000 ;
	    RECT 25.8000 920.4000 27.0000 921.6000 ;
	    RECT 18.6000 917.4000 19.8000 918.6000 ;
	    RECT 18.7500 858.6000 19.6500 917.4000 ;
	    RECT 25.9500 864.6000 26.8500 920.4000 ;
	    RECT 33.1500 918.6000 34.0500 947.4000 ;
	    RECT 35.5500 942.6000 36.4500 983.4000 ;
	    RECT 35.4000 941.4000 36.6000 942.6000 ;
	    RECT 37.8000 941.4000 39.0000 942.6000 ;
	    RECT 47.5500 918.6000 48.4500 1271.4000 ;
	    RECT 57.1500 1260.6000 58.0500 1283.4000 ;
	    RECT 57.0000 1259.4000 58.2000 1260.6000 ;
	    RECT 54.6000 1187.4000 55.8000 1188.6000 ;
	    RECT 59.4000 1187.4000 60.6000 1188.6000 ;
	    RECT 54.7500 1185.6000 55.6500 1187.4000 ;
	    RECT 49.8000 1184.4000 51.0000 1185.6000 ;
	    RECT 54.6000 1184.4000 55.8000 1185.6000 ;
	    RECT 49.9500 1161.6000 50.8500 1184.4000 ;
	    RECT 59.5500 1182.6000 60.4500 1187.4000 ;
	    RECT 59.4000 1181.4000 60.6000 1182.6000 ;
	    RECT 71.4000 1181.4000 72.6000 1182.6000 ;
	    RECT 71.5500 1170.6000 72.4500 1181.4000 ;
	    RECT 71.4000 1169.4000 72.6000 1170.6000 ;
	    RECT 49.8000 1160.4000 51.0000 1161.6000 ;
	    RECT 49.8000 1097.4000 51.0000 1098.6000 ;
	    RECT 49.9500 1041.6000 50.8500 1097.4000 ;
	    RECT 57.0000 1079.4000 58.2000 1080.6000 ;
	    RECT 57.1500 1044.6000 58.0500 1079.4000 ;
	    RECT 57.0000 1043.4000 58.2000 1044.6000 ;
	    RECT 57.1500 1041.6000 58.0500 1043.4000 ;
	    RECT 49.8000 1040.4000 51.0000 1041.6000 ;
	    RECT 57.0000 1040.4000 58.2000 1041.6000 ;
	    RECT 66.6000 948.4500 67.8000 948.6000 ;
	    RECT 64.3500 947.5500 67.8000 948.4500 ;
	    RECT 64.3500 939.6000 65.2500 947.5500 ;
	    RECT 66.6000 947.4000 67.8000 947.5500 ;
	    RECT 71.4000 941.4000 72.6000 942.6000 ;
	    RECT 64.2000 938.4000 65.4000 939.6000 ;
	    RECT 71.5500 924.6000 72.4500 941.4000 ;
	    RECT 66.6000 923.4000 67.8000 924.6000 ;
	    RECT 71.4000 923.4000 72.6000 924.6000 ;
	    RECT 66.7500 921.6000 67.6500 923.4000 ;
	    RECT 54.6000 920.4000 55.8000 921.6000 ;
	    RECT 66.6000 920.4000 67.8000 921.6000 ;
	    RECT 33.0000 917.4000 34.2000 918.6000 ;
	    RECT 47.4000 917.4000 48.6000 918.6000 ;
	    RECT 47.4000 914.4000 48.6000 915.6000 ;
	    RECT 47.5500 912.6000 48.4500 914.4000 ;
	    RECT 47.4000 911.4000 48.6000 912.6000 ;
	    RECT 49.8000 881.4000 51.0000 882.6000 ;
	    RECT 52.2000 881.4000 53.4000 882.6000 ;
	    RECT 25.8000 863.4000 27.0000 864.6000 ;
	    RECT 25.9500 861.6000 26.8500 863.4000 ;
	    RECT 25.8000 860.4000 27.0000 861.6000 ;
	    RECT 47.4000 860.4000 48.6000 861.6000 ;
	    RECT 18.6000 857.4000 19.8000 858.6000 ;
	    RECT 23.4000 857.4000 24.6000 858.6000 ;
	    RECT 18.6000 854.4000 19.8000 855.6000 ;
	    RECT 18.7500 852.6000 19.6500 854.4000 ;
	    RECT 18.6000 851.4000 19.8000 852.6000 ;
	    RECT 18.6000 713.4000 19.8000 714.6000 ;
	    RECT 18.7500 648.6000 19.6500 713.4000 ;
	    RECT 18.6000 647.4000 19.8000 648.6000 ;
	    RECT 18.6000 563.4000 19.8000 564.6000 ;
	    RECT 18.7500 561.6000 19.6500 563.4000 ;
	    RECT 18.6000 560.4000 19.8000 561.6000 ;
	    RECT 23.5500 558.6000 24.4500 857.4000 ;
	    RECT 47.5500 798.6000 48.4500 860.4000 ;
	    RECT 47.4000 797.4000 48.6000 798.6000 ;
	    RECT 49.9500 762.6000 50.8500 881.4000 ;
	    RECT 52.3500 852.6000 53.2500 881.4000 ;
	    RECT 54.7500 864.6000 55.6500 920.4000 ;
	    RECT 71.4000 911.4000 72.6000 912.6000 ;
	    RECT 71.5500 864.6000 72.4500 911.4000 ;
	    RECT 78.7500 885.6000 79.6500 1325.4000 ;
	    RECT 83.4000 1307.4000 84.6000 1308.6000 ;
	    RECT 83.5500 1305.6000 84.4500 1307.4000 ;
	    RECT 83.4000 1304.4000 84.6000 1305.6000 ;
	    RECT 105.1500 1302.6000 106.0500 1355.4000 ;
	    RECT 126.6000 1331.4000 127.8000 1332.6000 ;
	    RECT 114.6000 1307.4000 115.8000 1308.6000 ;
	    RECT 81.0000 1301.4000 82.2000 1302.6000 ;
	    RECT 105.0000 1301.4000 106.2000 1302.6000 ;
	    RECT 107.4000 1301.4000 108.6000 1302.6000 ;
	    RECT 107.5500 1290.6000 108.4500 1301.4000 ;
	    RECT 107.4000 1289.4000 108.6000 1290.6000 ;
	    RECT 107.5500 1281.6000 108.4500 1289.4000 ;
	    RECT 83.4000 1280.4000 84.6000 1281.6000 ;
	    RECT 107.4000 1280.4000 108.6000 1281.6000 ;
	    RECT 112.2000 1280.4000 113.4000 1281.6000 ;
	    RECT 83.5500 1230.6000 84.4500 1280.4000 ;
	    RECT 93.0000 1277.4000 94.2000 1278.6000 ;
	    RECT 95.4000 1277.4000 96.6000 1278.6000 ;
	    RECT 85.8000 1274.4000 87.0000 1275.6000 ;
	    RECT 85.9500 1272.6000 86.8500 1274.4000 ;
	    RECT 85.8000 1271.4000 87.0000 1272.6000 ;
	    RECT 83.4000 1229.4000 84.6000 1230.6000 ;
	    RECT 93.1500 1182.6000 94.0500 1277.4000 ;
	    RECT 95.5500 1272.6000 96.4500 1277.4000 ;
	    RECT 95.4000 1271.4000 96.6000 1272.6000 ;
	    RECT 95.4000 1184.4000 96.6000 1185.6000 ;
	    RECT 81.0000 1181.4000 82.2000 1182.6000 ;
	    RECT 90.6000 1181.4000 91.8000 1182.6000 ;
	    RECT 93.0000 1181.4000 94.2000 1182.6000 ;
	    RECT 81.1500 1179.6000 82.0500 1181.4000 ;
	    RECT 81.0000 1178.4000 82.2000 1179.6000 ;
	    RECT 90.6000 1179.4501 91.8000 1179.6000 ;
	    RECT 95.5500 1179.4501 96.4500 1184.4000 ;
	    RECT 112.3500 1182.4501 113.2500 1280.4000 ;
	    RECT 114.7500 1266.6000 115.6500 1307.4000 ;
	    RECT 126.7500 1299.6000 127.6500 1331.4000 ;
	    RECT 126.6000 1298.4000 127.8000 1299.6000 ;
	    RECT 133.9500 1299.4501 134.8500 1424.4000 ;
	    RECT 136.2000 1416.3000 137.4000 1436.7001 ;
	    RECT 138.6000 1416.3000 139.8000 1436.7001 ;
	    RECT 141.0000 1416.3000 142.2000 1433.7001 ;
	    RECT 143.4000 1421.4000 144.6000 1422.6000 ;
	    RECT 145.8000 1416.3000 147.0000 1433.7001 ;
	    RECT 148.3500 1419.6000 149.2500 1445.5500 ;
	    RECT 148.2000 1418.4000 149.4000 1419.6000 ;
	    RECT 148.3500 1413.4501 149.2500 1418.4000 ;
	    RECT 150.6000 1416.3000 151.8000 1433.7001 ;
	    RECT 153.0000 1416.3000 154.2000 1436.7001 ;
	    RECT 155.4000 1416.3000 156.6000 1436.7001 ;
	    RECT 157.8000 1416.3000 159.0000 1436.7001 ;
	    RECT 160.2000 1415.4000 161.4000 1416.6000 ;
	    RECT 160.3500 1413.4501 161.2500 1415.4000 ;
	    RECT 148.3500 1412.5500 151.6500 1413.4501 ;
	    RECT 141.0000 1386.3000 142.2000 1406.7001 ;
	    RECT 143.4000 1386.3000 144.6000 1406.7001 ;
	    RECT 145.8000 1386.3000 147.0000 1406.7001 ;
	    RECT 148.2000 1389.3000 149.4000 1406.7001 ;
	    RECT 150.7500 1404.6000 151.6500 1412.5500 ;
	    RECT 157.9500 1412.5500 161.2500 1413.4501 ;
	    RECT 157.9500 1410.4501 158.8500 1412.5500 ;
	    RECT 155.5500 1409.5500 158.8500 1410.4501 ;
	    RECT 150.6000 1403.4000 151.8000 1404.6000 ;
	    RECT 136.2000 1364.4000 137.4000 1365.6000 ;
	    RECT 136.3500 1362.6000 137.2500 1364.4000 ;
	    RECT 136.2000 1361.4000 137.4000 1362.6000 ;
	    RECT 138.6000 1356.3000 139.8000 1376.7001 ;
	    RECT 141.0000 1356.3000 142.2000 1376.7001 ;
	    RECT 143.4000 1356.3000 144.6000 1373.7001 ;
	    RECT 145.8000 1361.4000 147.0000 1362.6000 ;
	    RECT 145.9500 1356.6000 146.8500 1361.4000 ;
	    RECT 145.8000 1355.4000 147.0000 1356.6000 ;
	    RECT 148.2000 1356.3000 149.4000 1373.7001 ;
	    RECT 150.7500 1359.6000 151.6500 1403.4000 ;
	    RECT 153.0000 1389.3000 154.2000 1406.7001 ;
	    RECT 155.5500 1401.6000 156.4500 1409.5500 ;
	    RECT 155.4000 1400.4000 156.6000 1401.6000 ;
	    RECT 157.8000 1389.3000 159.0000 1406.7001 ;
	    RECT 160.2000 1386.3000 161.4000 1406.7001 ;
	    RECT 162.6000 1386.3000 163.8000 1406.7001 ;
	    RECT 165.1500 1398.6000 166.0500 1457.4000 ;
	    RECT 177.1500 1452.6000 178.0500 1463.4000 ;
	    RECT 191.5500 1452.6000 192.4500 1463.4000 ;
	    RECT 225.1500 1461.6000 226.0500 1463.4000 ;
	    RECT 222.6000 1460.4000 223.8000 1461.6000 ;
	    RECT 225.0000 1460.4000 226.2000 1461.6000 ;
	    RECT 232.2000 1460.4000 233.4000 1461.6000 ;
	    RECT 256.2000 1460.4000 257.4000 1461.6000 ;
	    RECT 222.7500 1458.6000 223.6500 1460.4000 ;
	    RECT 232.3500 1458.6000 233.2500 1460.4000 ;
	    RECT 256.3500 1458.6000 257.2500 1460.4000 ;
	    RECT 222.6000 1457.4000 223.8000 1458.6000 ;
	    RECT 227.4000 1458.4501 228.6000 1458.6000 ;
	    RECT 229.8000 1458.4501 231.0000 1458.6000 ;
	    RECT 227.4000 1457.5500 231.0000 1458.4501 ;
	    RECT 227.4000 1457.4000 228.6000 1457.5500 ;
	    RECT 229.8000 1457.4000 231.0000 1457.5500 ;
	    RECT 232.2000 1457.4000 233.4000 1458.6000 ;
	    RECT 256.2000 1457.4000 257.4000 1458.6000 ;
	    RECT 265.8000 1457.4000 267.0000 1458.6000 ;
	    RECT 225.0000 1454.4000 226.2000 1455.6000 ;
	    RECT 177.0000 1451.4000 178.2000 1452.6000 ;
	    RECT 191.4000 1451.4000 192.6000 1452.6000 ;
	    RECT 172.2000 1430.4000 173.4000 1431.6000 ;
	    RECT 165.0000 1397.4000 166.2000 1398.6000 ;
	    RECT 169.8000 1397.4000 171.0000 1398.6000 ;
	    RECT 165.1500 1392.6000 166.0500 1397.4000 ;
	    RECT 169.9500 1395.6000 170.8500 1397.4000 ;
	    RECT 169.8000 1394.4000 171.0000 1395.6000 ;
	    RECT 165.0000 1391.4000 166.2000 1392.6000 ;
	    RECT 169.8000 1391.4000 171.0000 1392.6000 ;
	    RECT 150.6000 1358.4000 151.8000 1359.6000 ;
	    RECT 150.7500 1353.4501 151.6500 1358.4000 ;
	    RECT 153.0000 1356.3000 154.2000 1373.7001 ;
	    RECT 155.4000 1356.3000 156.6000 1376.7001 ;
	    RECT 157.8000 1356.3000 159.0000 1376.7001 ;
	    RECT 160.2000 1356.3000 161.4000 1376.7001 ;
	    RECT 167.4000 1361.4000 168.6000 1362.6000 ;
	    RECT 150.7500 1352.5500 154.0500 1353.4501 ;
	    RECT 143.4000 1326.3000 144.6000 1346.7001 ;
	    RECT 145.8000 1326.3000 147.0000 1346.7001 ;
	    RECT 148.2000 1326.3000 149.4000 1346.7001 ;
	    RECT 150.6000 1329.3000 151.8000 1346.7001 ;
	    RECT 153.1500 1344.6000 154.0500 1352.5500 ;
	    RECT 153.0000 1343.4000 154.2000 1344.6000 ;
	    RECT 153.1500 1326.6000 154.0500 1343.4000 ;
	    RECT 155.4000 1329.3000 156.6000 1346.7001 ;
	    RECT 157.8000 1340.4000 159.0000 1341.6000 ;
	    RECT 153.0000 1325.4000 154.2000 1326.6000 ;
	    RECT 157.9500 1326.4501 158.8500 1340.4000 ;
	    RECT 160.2000 1329.3000 161.4000 1346.7001 ;
	    RECT 157.9500 1325.5500 161.2500 1326.4501 ;
	    RECT 162.6000 1326.3000 163.8000 1346.7001 ;
	    RECT 165.0000 1326.3000 166.2000 1346.7001 ;
	    RECT 167.5500 1338.6000 168.4500 1361.4000 ;
	    RECT 167.4000 1337.4000 168.6000 1338.6000 ;
	    RECT 153.1500 1314.6000 154.0500 1325.4000 ;
	    RECT 153.0000 1313.4000 154.2000 1314.6000 ;
	    RECT 160.3500 1302.6000 161.2500 1325.5500 ;
	    RECT 162.6000 1307.4000 163.8000 1308.6000 ;
	    RECT 153.0000 1301.4000 154.2000 1302.6000 ;
	    RECT 160.2000 1301.4000 161.4000 1302.6000 ;
	    RECT 133.9500 1298.5500 137.2500 1299.4501 ;
	    RECT 114.6000 1265.4000 115.8000 1266.6000 ;
	    RECT 121.8000 1259.4000 123.0000 1260.6000 ;
	    RECT 119.4000 1187.4000 120.6000 1188.6000 ;
	    RECT 114.6000 1182.4501 115.8000 1182.6000 ;
	    RECT 112.3500 1181.5500 115.8000 1182.4501 ;
	    RECT 114.6000 1181.4000 115.8000 1181.5500 ;
	    RECT 90.6000 1178.5500 96.4500 1179.4501 ;
	    RECT 90.6000 1178.4000 91.8000 1178.5500 ;
	    RECT 100.2000 1178.4000 101.4000 1179.6000 ;
	    RECT 112.2000 1178.4000 113.4000 1179.6000 ;
	    RECT 85.8000 1151.4000 87.0000 1152.6000 ;
	    RECT 83.4000 1049.4000 84.6000 1050.6000 ;
	    RECT 83.5500 1044.6000 84.4500 1049.4000 ;
	    RECT 85.9500 1044.6000 86.8500 1151.4000 ;
	    RECT 100.3500 1044.6000 101.2500 1178.4000 ;
	    RECT 112.3500 1176.6000 113.2500 1178.4000 ;
	    RECT 119.5500 1176.6000 120.4500 1187.4000 ;
	    RECT 112.2000 1175.4000 113.4000 1176.6000 ;
	    RECT 119.4000 1175.4000 120.6000 1176.6000 ;
	    RECT 114.6000 1151.4000 115.8000 1152.6000 ;
	    RECT 83.4000 1043.4000 84.6000 1044.6000 ;
	    RECT 85.8000 1043.4000 87.0000 1044.6000 ;
	    RECT 100.2000 1043.4000 101.4000 1044.6000 ;
	    RECT 81.0000 929.4000 82.2000 930.6000 ;
	    RECT 78.6000 884.4000 79.8000 885.6000 ;
	    RECT 54.6000 863.4000 55.8000 864.6000 ;
	    RECT 71.4000 863.4000 72.6000 864.6000 ;
	    RECT 54.7500 861.6000 55.6500 863.4000 ;
	    RECT 54.6000 860.4000 55.8000 861.6000 ;
	    RECT 52.2000 851.4000 53.4000 852.6000 ;
	    RECT 71.5500 792.6000 72.4500 863.4000 ;
	    RECT 71.4000 791.4000 72.6000 792.6000 ;
	    RECT 49.8000 761.4000 51.0000 762.6000 ;
	    RECT 49.9500 702.6000 50.8500 761.4000 ;
	    RECT 52.2000 749.4000 53.4000 750.6000 ;
	    RECT 49.8000 701.4000 51.0000 702.6000 ;
	    RECT 49.9500 681.6000 50.8500 701.4000 ;
	    RECT 49.8000 680.4000 51.0000 681.6000 ;
	    RECT 42.6000 653.4000 43.8000 654.6000 ;
	    RECT 40.2000 647.4000 41.4000 648.6000 ;
	    RECT 40.3500 642.6000 41.2500 647.4000 ;
	    RECT 42.7500 645.6000 43.6500 653.4000 ;
	    RECT 42.6000 644.4000 43.8000 645.6000 ;
	    RECT 47.4000 644.4000 48.6000 645.6000 ;
	    RECT 40.2000 641.4000 41.4000 642.6000 ;
	    RECT 23.4000 557.4000 24.6000 558.6000 ;
	    RECT 40.2000 557.4000 41.4000 558.6000 ;
	    RECT 13.8000 491.4000 15.0000 492.6000 ;
	    RECT 13.9500 444.6000 14.8500 491.4000 ;
	    RECT 13.8000 443.4000 15.0000 444.6000 ;
	    RECT 13.9500 360.6000 14.8500 443.4000 ;
	    RECT 16.2000 398.4000 17.4000 399.6000 ;
	    RECT 13.8000 359.4000 15.0000 360.6000 ;
	    RECT 16.3500 354.4500 17.2500 398.4000 ;
	    RECT 13.9500 353.5500 17.2500 354.4500 ;
	    RECT 13.9500 159.6000 14.8500 353.5500 ;
	    RECT 23.5500 348.6000 24.4500 557.4000 ;
	    RECT 40.3500 441.6000 41.2500 557.4000 ;
	    RECT 47.5500 555.6000 48.4500 644.4000 ;
	    RECT 52.3500 642.6000 53.2500 749.4000 ;
	    RECT 71.5500 699.6000 72.4500 791.4000 ;
	    RECT 81.1500 705.6000 82.0500 929.4000 ;
	    RECT 85.9500 888.6000 86.8500 1043.4000 ;
	    RECT 100.2000 1040.4000 101.4000 1041.6000 ;
	    RECT 100.3500 1032.6000 101.2500 1040.4000 ;
	    RECT 100.2000 1031.4000 101.4000 1032.6000 ;
	    RECT 95.4000 959.4000 96.6000 960.6000 ;
	    RECT 95.5500 942.6000 96.4500 959.4000 ;
	    RECT 95.4000 941.4000 96.6000 942.6000 ;
	    RECT 102.6000 941.4000 103.8000 942.6000 ;
	    RECT 85.8000 887.4000 87.0000 888.6000 ;
	    RECT 88.2000 884.4000 89.4000 885.6000 ;
	    RECT 81.0000 704.4000 82.2000 705.6000 ;
	    RECT 71.4000 698.4000 72.6000 699.6000 ;
	    RECT 88.3500 675.6000 89.2500 884.4000 ;
	    RECT 102.7500 882.6000 103.6500 941.4000 ;
	    RECT 109.8000 914.4000 111.0000 915.6000 ;
	    RECT 102.6000 881.4000 103.8000 882.6000 ;
	    RECT 102.7500 864.6000 103.6500 881.4000 ;
	    RECT 109.9500 879.6000 110.8500 914.4000 ;
	    RECT 121.9500 882.6000 122.8500 1259.4000 ;
	    RECT 124.2000 1247.4000 125.4000 1248.6000 ;
	    RECT 126.7500 1134.6000 127.6500 1298.4000 ;
	    RECT 133.8000 1295.4000 135.0000 1296.6000 ;
	    RECT 131.4000 1256.4000 132.6000 1257.6000 ;
	    RECT 131.5500 1248.6000 132.4500 1256.4000 ;
	    RECT 131.4000 1247.4000 132.6000 1248.6000 ;
	    RECT 133.9500 1218.6000 134.8500 1295.4000 ;
	    RECT 136.3500 1245.6000 137.2500 1298.5500 ;
	    RECT 153.1500 1290.6000 154.0500 1301.4000 ;
	    RECT 153.0000 1289.4000 154.2000 1290.6000 ;
	    RECT 136.2000 1244.4000 137.4000 1245.6000 ;
	    RECT 138.6000 1236.3000 139.8000 1256.7001 ;
	    RECT 141.0000 1236.3000 142.2000 1256.7001 ;
	    RECT 143.4000 1236.3000 144.6000 1253.7001 ;
	    RECT 145.8000 1247.4000 147.0000 1248.6000 ;
	    RECT 145.9500 1242.6000 146.8500 1247.4000 ;
	    RECT 145.8000 1241.4000 147.0000 1242.6000 ;
	    RECT 148.2000 1236.3000 149.4000 1253.7001 ;
	    RECT 150.6000 1238.4000 151.8000 1239.6000 ;
	    RECT 150.7500 1233.4501 151.6500 1238.4000 ;
	    RECT 153.0000 1236.3000 154.2000 1253.7001 ;
	    RECT 155.4000 1236.3000 156.6000 1256.7001 ;
	    RECT 157.8000 1236.3000 159.0000 1256.7001 ;
	    RECT 160.2000 1236.3000 161.4000 1256.7001 ;
	    RECT 162.7500 1248.6000 163.6500 1307.4000 ;
	    RECT 167.5500 1284.6000 168.4500 1337.4000 ;
	    RECT 169.9500 1326.6000 170.8500 1391.4000 ;
	    RECT 172.3500 1374.6000 173.2500 1430.4000 ;
	    RECT 177.0000 1415.4000 178.2000 1416.6000 ;
	    RECT 177.1500 1401.6000 178.0500 1415.4000 ;
	    RECT 177.0000 1400.4000 178.2000 1401.6000 ;
	    RECT 220.2000 1400.4000 221.4000 1401.6000 ;
	    RECT 174.6000 1397.4000 175.8000 1398.6000 ;
	    RECT 203.4000 1397.4000 204.6000 1398.6000 ;
	    RECT 172.2000 1373.4000 173.4000 1374.6000 ;
	    RECT 172.2000 1334.4000 173.4000 1335.6000 ;
	    RECT 172.3500 1326.6000 173.2500 1334.4000 ;
	    RECT 169.8000 1325.4000 171.0000 1326.6000 ;
	    RECT 172.2000 1326.4501 173.4000 1326.6000 ;
	    RECT 174.7500 1326.4501 175.6500 1397.4000 ;
	    RECT 198.6000 1394.4000 199.8000 1395.6000 ;
	    RECT 196.2000 1391.4000 197.4000 1392.6000 ;
	    RECT 189.0000 1379.4000 190.2000 1380.6000 ;
	    RECT 179.4000 1370.4000 180.6000 1371.6000 ;
	    RECT 179.5500 1344.6000 180.4500 1370.4000 ;
	    RECT 189.1500 1359.6000 190.0500 1379.4000 ;
	    RECT 196.3500 1362.6000 197.2500 1391.4000 ;
	    RECT 198.7500 1386.6000 199.6500 1394.4000 ;
	    RECT 203.5500 1392.6000 204.4500 1397.4000 ;
	    RECT 203.4000 1391.4000 204.6000 1392.6000 ;
	    RECT 198.6000 1385.4000 199.8000 1386.6000 ;
	    RECT 217.8000 1373.4000 219.0000 1374.6000 ;
	    RECT 196.2000 1361.4000 197.4000 1362.6000 ;
	    RECT 189.0000 1358.4000 190.2000 1359.6000 ;
	    RECT 179.4000 1343.4000 180.6000 1344.6000 ;
	    RECT 172.2000 1325.5500 175.6500 1326.4501 ;
	    RECT 172.2000 1325.4000 173.4000 1325.5500 ;
	    RECT 167.4000 1283.4000 168.6000 1284.6000 ;
	    RECT 162.6000 1247.4000 163.8000 1248.6000 ;
	    RECT 148.3500 1232.5500 151.6500 1233.4501 ;
	    RECT 143.4000 1229.4000 144.6000 1230.6000 ;
	    RECT 133.8000 1217.4000 135.0000 1218.6000 ;
	    RECT 129.0000 1214.4000 130.2000 1215.6000 ;
	    RECT 129.1500 1206.6000 130.0500 1214.4000 ;
	    RECT 129.0000 1205.4000 130.2000 1206.6000 ;
	    RECT 133.9500 1179.4501 134.8500 1217.4000 ;
	    RECT 136.2000 1206.3000 137.4000 1226.7001 ;
	    RECT 138.6000 1206.3000 139.8000 1226.7001 ;
	    RECT 141.0000 1209.3000 142.2000 1226.7001 ;
	    RECT 143.5500 1221.6000 144.4500 1229.4000 ;
	    RECT 143.4000 1220.4000 144.6000 1221.6000 ;
	    RECT 145.8000 1209.3000 147.0000 1226.7001 ;
	    RECT 148.3500 1224.6000 149.2500 1232.5500 ;
	    RECT 148.2000 1223.4000 149.4000 1224.6000 ;
	    RECT 133.9500 1178.5500 137.2500 1179.4501 ;
	    RECT 133.8000 1175.4000 135.0000 1176.6000 ;
	    RECT 126.6000 1134.4501 127.8000 1134.6000 ;
	    RECT 124.3500 1133.5500 127.8000 1134.4501 ;
	    RECT 124.3500 1119.4501 125.2500 1133.5500 ;
	    RECT 126.6000 1133.4000 127.8000 1133.5500 ;
	    RECT 126.6000 1130.4000 127.8000 1131.6000 ;
	    RECT 126.7500 1128.6000 127.6500 1130.4000 ;
	    RECT 126.6000 1127.4000 127.8000 1128.6000 ;
	    RECT 131.4000 1127.4000 132.6000 1128.6000 ;
	    RECT 131.5500 1122.6000 132.4500 1127.4000 ;
	    RECT 131.4000 1121.4000 132.6000 1122.6000 ;
	    RECT 124.3500 1118.5500 127.6500 1119.4501 ;
	    RECT 124.2000 959.4000 125.4000 960.6000 ;
	    RECT 124.3500 954.6000 125.2500 959.4000 ;
	    RECT 124.2000 953.4000 125.4000 954.6000 ;
	    RECT 126.7500 924.6000 127.6500 1118.5500 ;
	    RECT 133.9500 1098.6000 134.8500 1175.4000 ;
	    RECT 136.3500 1110.6000 137.2500 1178.5500 ;
	    RECT 148.3500 1164.4501 149.2500 1223.4000 ;
	    RECT 150.6000 1209.3000 151.8000 1226.7001 ;
	    RECT 153.0000 1206.3000 154.2000 1226.7001 ;
	    RECT 155.4000 1206.3000 156.6000 1226.7001 ;
	    RECT 157.8000 1206.3000 159.0000 1226.7001 ;
	    RECT 169.9500 1200.6000 170.8500 1325.4000 ;
	    RECT 179.5500 1308.6000 180.4500 1343.4000 ;
	    RECT 181.8000 1340.4000 183.0000 1341.6000 ;
	    RECT 181.9500 1308.6000 182.8500 1340.4000 ;
	    RECT 179.4000 1307.4000 180.6000 1308.6000 ;
	    RECT 181.8000 1307.4000 183.0000 1308.6000 ;
	    RECT 174.6000 1259.4000 175.8000 1260.6000 ;
	    RECT 174.7500 1251.6000 175.6500 1259.4000 ;
	    RECT 174.6000 1250.4000 175.8000 1251.6000 ;
	    RECT 179.5500 1239.6000 180.4500 1307.4000 ;
	    RECT 184.2000 1301.4000 185.4000 1302.6000 ;
	    RECT 184.3500 1290.6000 185.2500 1301.4000 ;
	    RECT 184.2000 1289.4000 185.4000 1290.6000 ;
	    RECT 179.4000 1238.4000 180.6000 1239.6000 ;
	    RECT 189.1500 1224.6000 190.0500 1358.4000 ;
	    RECT 196.2000 1307.4000 197.4000 1308.6000 ;
	    RECT 196.3500 1305.6000 197.2500 1307.4000 ;
	    RECT 196.2000 1304.4000 197.4000 1305.6000 ;
	    RECT 196.2000 1298.4000 197.4000 1299.6000 ;
	    RECT 196.3500 1275.6000 197.2500 1298.4000 ;
	    RECT 196.2000 1274.4000 197.4000 1275.6000 ;
	    RECT 196.3500 1272.6000 197.2500 1274.4000 ;
	    RECT 196.2000 1271.4000 197.4000 1272.6000 ;
	    RECT 213.0000 1271.4000 214.2000 1272.6000 ;
	    RECT 213.1500 1224.6000 214.0500 1271.4000 ;
	    RECT 189.0000 1223.4000 190.2000 1224.6000 ;
	    RECT 213.0000 1223.4000 214.2000 1224.6000 ;
	    RECT 198.6000 1220.4000 199.8000 1221.6000 ;
	    RECT 172.2000 1211.4000 173.4000 1212.6000 ;
	    RECT 155.4000 1199.4000 156.6000 1200.6000 ;
	    RECT 169.8000 1199.4000 171.0000 1200.6000 ;
	    RECT 150.6000 1175.4000 151.8000 1176.6000 ;
	    RECT 150.7500 1170.6000 151.6500 1175.4000 ;
	    RECT 150.6000 1169.4000 151.8000 1170.6000 ;
	    RECT 150.6000 1164.4501 151.8000 1164.6000 ;
	    RECT 148.3500 1163.5500 151.8000 1164.4501 ;
	    RECT 150.6000 1163.4000 151.8000 1163.5500 ;
	    RECT 141.0000 1116.3000 142.2000 1136.7001 ;
	    RECT 143.4000 1116.3000 144.6000 1136.7001 ;
	    RECT 145.8000 1116.3000 147.0000 1136.7001 ;
	    RECT 148.2000 1116.3000 149.4000 1133.7001 ;
	    RECT 150.7500 1119.6000 151.6500 1163.4000 ;
	    RECT 155.5500 1140.6000 156.4500 1199.4000 ;
	    RECT 172.3500 1188.6000 173.2500 1211.4000 ;
	    RECT 172.2000 1187.4000 173.4000 1188.6000 ;
	    RECT 189.0000 1187.4000 190.2000 1188.6000 ;
	    RECT 172.2000 1175.4000 173.4000 1176.6000 ;
	    RECT 157.8000 1146.3000 159.0000 1166.7001 ;
	    RECT 160.2000 1146.3000 161.4000 1166.7001 ;
	    RECT 162.6000 1146.3000 163.8000 1166.7001 ;
	    RECT 165.0000 1149.3000 166.2000 1166.7001 ;
	    RECT 167.4000 1163.4000 168.6000 1164.6000 ;
	    RECT 169.8000 1149.3000 171.0000 1166.7001 ;
	    RECT 172.3500 1161.6000 173.2500 1175.4000 ;
	    RECT 172.2000 1160.4000 173.4000 1161.6000 ;
	    RECT 174.6000 1149.3000 175.8000 1166.7001 ;
	    RECT 177.0000 1146.3000 178.2000 1166.7001 ;
	    RECT 179.4000 1146.3000 180.6000 1166.7001 ;
	    RECT 181.8000 1157.4000 183.0000 1158.6000 ;
	    RECT 181.9500 1152.6000 182.8500 1157.4000 ;
	    RECT 186.6000 1154.4000 187.8000 1155.6000 ;
	    RECT 181.8000 1151.4000 183.0000 1152.6000 ;
	    RECT 155.4000 1139.4000 156.6000 1140.6000 ;
	    RECT 165.0000 1139.4000 166.2000 1140.6000 ;
	    RECT 150.6000 1118.4000 151.8000 1119.6000 ;
	    RECT 150.7500 1113.4501 151.6500 1118.4000 ;
	    RECT 153.0000 1116.3000 154.2000 1133.7001 ;
	    RECT 155.4000 1121.4000 156.6000 1122.6000 ;
	    RECT 155.5500 1116.6000 156.4500 1121.4000 ;
	    RECT 155.4000 1115.4000 156.6000 1116.6000 ;
	    RECT 157.8000 1116.3000 159.0000 1133.7001 ;
	    RECT 160.2000 1116.3000 161.4000 1136.7001 ;
	    RECT 162.6000 1116.3000 163.8000 1136.7001 ;
	    RECT 165.1500 1125.6000 166.0500 1139.4000 ;
	    RECT 169.8000 1136.4000 171.0000 1137.6000 ;
	    RECT 169.9500 1128.6000 170.8500 1136.4000 ;
	    RECT 181.9500 1128.6000 182.8500 1151.4000 ;
	    RECT 186.7500 1146.6000 187.6500 1154.4000 ;
	    RECT 189.1500 1146.6000 190.0500 1187.4000 ;
	    RECT 193.8000 1175.4000 195.0000 1176.6000 ;
	    RECT 196.2000 1154.4000 197.4000 1155.6000 ;
	    RECT 186.6000 1145.4000 187.8000 1146.6000 ;
	    RECT 189.0000 1145.4000 190.2000 1146.6000 ;
	    RECT 169.8000 1127.4000 171.0000 1128.6000 ;
	    RECT 181.8000 1127.4000 183.0000 1128.6000 ;
	    RECT 193.8000 1127.4000 195.0000 1128.6000 ;
	    RECT 165.0000 1124.4000 166.2000 1125.6000 ;
	    RECT 148.3500 1112.5500 151.6500 1113.4501 ;
	    RECT 136.2000 1109.4000 137.4000 1110.6000 ;
	    RECT 133.8000 1098.4501 135.0000 1098.6000 ;
	    RECT 131.5500 1097.5500 135.0000 1098.4501 ;
	    RECT 129.0000 1094.4000 130.2000 1095.6000 ;
	    RECT 129.1500 1086.6000 130.0500 1094.4000 ;
	    RECT 129.0000 1085.4000 130.2000 1086.6000 ;
	    RECT 129.0000 1076.4000 130.2000 1077.6000 ;
	    RECT 129.1500 1068.6000 130.0500 1076.4000 ;
	    RECT 129.0000 1067.4000 130.2000 1068.6000 ;
	    RECT 131.5500 1020.6000 132.4500 1097.5500 ;
	    RECT 133.8000 1097.4000 135.0000 1097.5500 ;
	    RECT 136.2000 1086.3000 137.4000 1106.7001 ;
	    RECT 138.6000 1086.3000 139.8000 1106.7001 ;
	    RECT 141.0000 1089.3000 142.2000 1106.7001 ;
	    RECT 143.4000 1100.4000 144.6000 1101.6000 ;
	    RECT 143.5500 1098.6000 144.4500 1100.4000 ;
	    RECT 143.4000 1097.4000 144.6000 1098.6000 ;
	    RECT 143.4000 1091.4000 144.6000 1092.6000 ;
	    RECT 133.8000 1073.4000 135.0000 1074.6000 ;
	    RECT 133.9500 1065.6000 134.8500 1073.4000 ;
	    RECT 133.8000 1064.4000 135.0000 1065.6000 ;
	    RECT 133.8000 1061.4000 135.0000 1062.6000 ;
	    RECT 131.4000 1019.4000 132.6000 1020.6000 ;
	    RECT 131.4000 1016.4000 132.6000 1017.6000 ;
	    RECT 131.5500 1008.6000 132.4500 1016.4000 ;
	    RECT 131.4000 1007.4000 132.6000 1008.6000 ;
	    RECT 133.9500 978.4500 134.8500 1061.4000 ;
	    RECT 136.2000 1056.3000 137.4000 1076.7001 ;
	    RECT 138.6000 1056.3000 139.8000 1076.7001 ;
	    RECT 141.0000 1056.3000 142.2000 1073.7001 ;
	    RECT 143.5500 1068.6000 144.4500 1091.4000 ;
	    RECT 145.8000 1089.3000 147.0000 1106.7001 ;
	    RECT 148.3500 1104.6000 149.2500 1112.5500 ;
	    RECT 160.2000 1109.4000 161.4000 1110.6000 ;
	    RECT 148.2000 1103.4000 149.4000 1104.6000 ;
	    RECT 143.4000 1067.4000 144.6000 1068.6000 ;
	    RECT 143.4000 1061.4000 144.6000 1062.6000 ;
	    RECT 143.5500 1044.6000 144.4500 1061.4000 ;
	    RECT 145.8000 1056.3000 147.0000 1073.7001 ;
	    RECT 148.3500 1059.6000 149.2500 1103.4000 ;
	    RECT 150.6000 1089.3000 151.8000 1106.7001 ;
	    RECT 153.0000 1086.3000 154.2000 1106.7001 ;
	    RECT 155.4000 1086.3000 156.6000 1106.7001 ;
	    RECT 157.8000 1086.3000 159.0000 1106.7001 ;
	    RECT 160.3500 1092.6000 161.2500 1109.4000 ;
	    RECT 165.1500 1098.6000 166.0500 1124.4000 ;
	    RECT 177.0000 1121.4000 178.2000 1122.6000 ;
	    RECT 177.1500 1119.6000 178.0500 1121.4000 ;
	    RECT 177.0000 1118.4000 178.2000 1119.6000 ;
	    RECT 179.4000 1118.4000 180.6000 1119.6000 ;
	    RECT 165.0000 1097.4000 166.2000 1098.6000 ;
	    RECT 169.8000 1097.4000 171.0000 1098.6000 ;
	    RECT 160.2000 1091.4000 161.4000 1092.6000 ;
	    RECT 162.6000 1085.4000 163.8000 1086.6000 ;
	    RECT 148.2000 1058.4000 149.4000 1059.6000 ;
	    RECT 143.4000 1043.4000 144.6000 1044.6000 ;
	    RECT 138.6000 1040.4000 139.8000 1041.6000 ;
	    RECT 145.8000 1040.4000 147.0000 1041.6000 ;
	    RECT 136.2000 1037.4000 137.4000 1038.6000 ;
	    RECT 136.3500 1023.4500 137.2500 1037.4000 ;
	    RECT 138.7500 1026.6000 139.6500 1040.4000 ;
	    RECT 141.0000 1037.4000 142.2000 1038.6000 ;
	    RECT 143.4000 1037.4000 144.6000 1038.6000 ;
	    RECT 138.6000 1025.4000 139.8000 1026.6000 ;
	    RECT 141.1500 1023.4500 142.0500 1037.4000 ;
	    RECT 136.3500 1022.5500 142.0500 1023.4500 ;
	    RECT 143.5500 1020.6000 144.4500 1037.4000 ;
	    RECT 145.9500 1032.6000 146.8500 1040.4000 ;
	    RECT 145.8000 1031.4000 147.0000 1032.6000 ;
	    RECT 148.3500 1023.4500 149.2500 1058.4000 ;
	    RECT 150.6000 1056.3000 151.8000 1073.7001 ;
	    RECT 153.0000 1056.3000 154.2000 1076.7001 ;
	    RECT 155.4000 1056.3000 156.6000 1076.7001 ;
	    RECT 157.8000 1056.3000 159.0000 1076.7001 ;
	    RECT 162.7500 1050.6000 163.6500 1085.4000 ;
	    RECT 165.0000 1073.4000 166.2000 1074.6000 ;
	    RECT 162.6000 1049.4000 163.8000 1050.6000 ;
	    RECT 150.6000 1031.4000 151.8000 1032.6000 ;
	    RECT 150.7500 1026.6000 151.6500 1031.4000 ;
	    RECT 150.6000 1025.4000 151.8000 1026.6000 ;
	    RECT 148.3500 1022.5500 151.6500 1023.4500 ;
	    RECT 136.2000 1019.4000 137.4000 1020.6000 ;
	    RECT 143.4000 1019.4000 144.6000 1020.6000 ;
	    RECT 136.3500 1005.6000 137.2500 1019.4000 ;
	    RECT 136.2000 1004.4000 137.4000 1005.6000 ;
	    RECT 138.6000 996.3000 139.8000 1016.7000 ;
	    RECT 141.0000 996.3000 142.2000 1016.7000 ;
	    RECT 143.4000 996.3000 144.6000 1013.7000 ;
	    RECT 145.8000 1001.4000 147.0000 1002.6000 ;
	    RECT 145.9500 993.4500 146.8500 1001.4000 ;
	    RECT 148.2000 996.3000 149.4000 1013.7000 ;
	    RECT 150.7500 999.6000 151.6500 1022.5500 ;
	    RECT 150.6000 998.4000 151.8000 999.6000 ;
	    RECT 143.5500 992.5500 146.8500 993.4500 ;
	    RECT 143.5500 990.6000 144.4500 992.5500 ;
	    RECT 136.2000 989.4000 137.4000 990.6000 ;
	    RECT 143.4000 989.4000 144.6000 990.6000 ;
	    RECT 136.3500 984.6000 137.2500 989.4000 ;
	    RECT 136.2000 983.4000 137.4000 984.6000 ;
	    RECT 136.2000 978.4500 137.4000 978.6000 ;
	    RECT 133.9500 977.5500 137.4000 978.4500 ;
	    RECT 136.2000 977.4000 137.4000 977.5500 ;
	    RECT 131.4000 974.4000 132.6000 975.6000 ;
	    RECT 131.5500 966.6000 132.4500 974.4000 ;
	    RECT 131.4000 965.4000 132.6000 966.6000 ;
	    RECT 131.4000 959.4000 132.6000 960.6000 ;
	    RECT 131.5500 939.6000 132.4500 959.4000 ;
	    RECT 133.8000 947.4000 135.0000 948.6000 ;
	    RECT 133.9500 939.6000 134.8500 947.4000 ;
	    RECT 131.4000 938.4000 132.6000 939.6000 ;
	    RECT 133.8000 938.4000 135.0000 939.6000 ;
	    RECT 126.6000 923.4000 127.8000 924.6000 ;
	    RECT 117.0000 881.4000 118.2000 882.6000 ;
	    RECT 121.8000 881.4000 123.0000 882.6000 ;
	    RECT 109.8000 878.4000 111.0000 879.6000 ;
	    RECT 102.6000 863.4000 103.8000 864.6000 ;
	    RECT 102.7500 861.6000 103.6500 863.4000 ;
	    RECT 102.6000 860.4000 103.8000 861.6000 ;
	    RECT 90.6000 854.4000 91.8000 855.6000 ;
	    RECT 90.7500 786.6000 91.6500 854.4000 ;
	    RECT 109.9500 831.6000 110.8500 878.4000 ;
	    RECT 117.1500 858.6000 118.0500 881.4000 ;
	    RECT 121.8000 878.4000 123.0000 879.6000 ;
	    RECT 119.4000 860.4000 120.6000 861.6000 ;
	    RECT 117.0000 857.4000 118.2000 858.6000 ;
	    RECT 109.8000 830.4000 111.0000 831.6000 ;
	    RECT 119.5500 822.6000 120.4500 860.4000 ;
	    RECT 119.4000 821.4000 120.6000 822.6000 ;
	    RECT 90.6000 785.4000 91.8000 786.6000 ;
	    RECT 90.7500 732.6000 91.6500 785.4000 ;
	    RECT 114.6000 773.4000 115.8000 774.6000 ;
	    RECT 105.0000 761.4000 106.2000 762.6000 ;
	    RECT 90.6000 731.4000 91.8000 732.6000 ;
	    RECT 97.8000 731.4000 99.0000 732.6000 ;
	    RECT 95.4000 701.4000 96.6000 702.6000 ;
	    RECT 95.5500 696.6000 96.4500 701.4000 ;
	    RECT 97.9500 699.6000 98.8500 731.4000 ;
	    RECT 102.6000 701.4000 103.8000 702.6000 ;
	    RECT 97.8000 698.4000 99.0000 699.6000 ;
	    RECT 95.4000 695.4000 96.6000 696.6000 ;
	    RECT 102.7500 681.6000 103.6500 701.4000 ;
	    RECT 95.4000 680.4000 96.6000 681.6000 ;
	    RECT 102.6000 680.4000 103.8000 681.6000 ;
	    RECT 93.0000 677.4000 94.2000 678.6000 ;
	    RECT 88.2000 674.4000 89.4000 675.6000 ;
	    RECT 66.6000 653.4000 67.8000 654.6000 ;
	    RECT 66.7500 648.6000 67.6500 653.4000 ;
	    RECT 66.6000 647.4000 67.8000 648.6000 ;
	    RECT 52.2000 641.4000 53.4000 642.6000 ;
	    RECT 71.4000 641.4000 72.6000 642.6000 ;
	    RECT 78.6000 641.4000 79.8000 642.6000 ;
	    RECT 71.5500 636.6000 72.4500 641.4000 ;
	    RECT 71.4000 635.4000 72.6000 636.6000 ;
	    RECT 78.7500 564.6000 79.6500 641.4000 ;
	    RECT 95.5500 600.6000 96.4500 680.4000 ;
	    RECT 102.7500 642.6000 103.6500 680.4000 ;
	    RECT 102.6000 641.4000 103.8000 642.6000 ;
	    RECT 95.4000 599.4000 96.6000 600.6000 ;
	    RECT 90.6000 587.4000 91.8000 588.6000 ;
	    RECT 57.0000 563.4000 58.2000 564.6000 ;
	    RECT 78.6000 563.4000 79.8000 564.6000 ;
	    RECT 57.1500 561.6000 58.0500 563.4000 ;
	    RECT 49.8000 560.4000 51.0000 561.6000 ;
	    RECT 57.0000 560.4000 58.2000 561.6000 ;
	    RECT 47.4000 554.4000 48.6000 555.6000 ;
	    RECT 49.9500 504.6000 50.8500 560.4000 ;
	    RECT 90.7500 555.6000 91.6500 587.4000 ;
	    RECT 93.0000 563.4000 94.2000 564.6000 ;
	    RECT 102.6000 563.4000 103.8000 564.6000 ;
	    RECT 93.1500 558.6000 94.0500 563.4000 ;
	    RECT 102.7500 561.6000 103.6500 563.4000 ;
	    RECT 95.4000 560.4000 96.6000 561.6000 ;
	    RECT 102.6000 560.4000 103.8000 561.6000 ;
	    RECT 93.0000 557.4000 94.2000 558.6000 ;
	    RECT 90.6000 554.4000 91.8000 555.6000 ;
	    RECT 95.5500 534.6000 96.4500 560.4000 ;
	    RECT 95.4000 533.4000 96.6000 534.6000 ;
	    RECT 49.8000 503.4000 51.0000 504.6000 ;
	    RECT 42.6000 491.4000 43.8000 492.6000 ;
	    RECT 35.4000 440.4000 36.6000 441.6000 ;
	    RECT 40.2000 440.4000 41.4000 441.6000 ;
	    RECT 35.5500 438.6000 36.4500 440.4000 ;
	    RECT 35.4000 437.4000 36.6000 438.6000 ;
	    RECT 35.4000 434.4000 36.6000 435.6000 ;
	    RECT 35.5500 420.6000 36.4500 434.4000 ;
	    RECT 35.4000 419.4000 36.6000 420.6000 ;
	    RECT 33.0000 413.4000 34.2000 414.6000 ;
	    RECT 33.1500 402.6000 34.0500 413.4000 ;
	    RECT 35.5500 408.6000 36.4500 419.4000 ;
	    RECT 35.4000 407.4000 36.6000 408.6000 ;
	    RECT 42.7500 402.6000 43.6500 491.4000 ;
	    RECT 85.8000 455.4000 87.0000 456.6000 ;
	    RECT 85.9500 441.6000 86.8500 455.4000 ;
	    RECT 64.2000 440.4000 65.4000 441.6000 ;
	    RECT 85.8000 440.4000 87.0000 441.6000 ;
	    RECT 88.2000 440.4000 89.4000 441.6000 ;
	    RECT 45.0000 437.4000 46.2000 438.6000 ;
	    RECT 33.0000 401.4000 34.2000 402.6000 ;
	    RECT 42.6000 401.4000 43.8000 402.6000 ;
	    RECT 40.2000 359.4000 41.4000 360.6000 ;
	    RECT 40.3500 348.6000 41.2500 359.4000 ;
	    RECT 23.4000 347.4000 24.6000 348.6000 ;
	    RECT 40.2000 347.4000 41.4000 348.6000 ;
	    RECT 23.5500 345.6000 24.4500 347.4000 ;
	    RECT 23.4000 344.4000 24.6000 345.6000 ;
	    RECT 30.6000 344.4000 31.8000 345.6000 ;
	    RECT 18.6000 341.4000 19.8000 342.6000 ;
	    RECT 25.8000 341.4000 27.0000 342.6000 ;
	    RECT 18.7500 282.6000 19.6500 341.4000 ;
	    RECT 25.9500 321.6000 26.8500 341.4000 ;
	    RECT 25.8000 320.4000 27.0000 321.6000 ;
	    RECT 28.2000 317.4000 29.4000 318.6000 ;
	    RECT 30.7500 288.6000 31.6500 344.4000 ;
	    RECT 33.0000 320.4000 34.2000 321.6000 ;
	    RECT 35.4000 320.4000 36.6000 321.6000 ;
	    RECT 25.8000 287.4000 27.0000 288.6000 ;
	    RECT 30.6000 287.4000 31.8000 288.6000 ;
	    RECT 25.9500 285.6000 26.8500 287.4000 ;
	    RECT 25.8000 284.4000 27.0000 285.6000 ;
	    RECT 18.6000 281.4000 19.8000 282.6000 ;
	    RECT 18.7500 198.6000 19.6500 281.4000 ;
	    RECT 25.8000 230.4000 27.0000 231.6000 ;
	    RECT 25.9500 201.6000 26.8500 230.4000 ;
	    RECT 33.1500 228.6000 34.0500 320.4000 ;
	    RECT 35.5500 318.6000 36.4500 320.4000 ;
	    RECT 35.4000 317.4000 36.6000 318.6000 ;
	    RECT 40.2000 317.4000 41.4000 318.6000 ;
	    RECT 40.3500 315.6000 41.2500 317.4000 ;
	    RECT 40.2000 314.4000 41.4000 315.6000 ;
	    RECT 33.0000 227.4000 34.2000 228.6000 ;
	    RECT 42.7500 216.6000 43.6500 401.4000 ;
	    RECT 42.6000 215.4000 43.8000 216.6000 ;
	    RECT 25.8000 200.4000 27.0000 201.6000 ;
	    RECT 18.6000 197.4000 19.8000 198.6000 ;
	    RECT 40.2000 197.4000 41.4000 198.6000 ;
	    RECT 18.7500 195.6000 19.6500 197.4000 ;
	    RECT 18.6000 194.4000 19.8000 195.6000 ;
	    RECT 18.7500 162.6000 19.6500 194.4000 ;
	    RECT 40.3500 168.6000 41.2500 197.4000 ;
	    RECT 45.1500 195.6000 46.0500 437.4000 ;
	    RECT 64.3500 420.6000 65.2500 440.4000 ;
	    RECT 66.6000 437.4000 67.8000 438.6000 ;
	    RECT 88.3500 420.6000 89.2500 440.4000 ;
	    RECT 64.2000 419.4000 65.4000 420.6000 ;
	    RECT 71.4000 419.4000 72.6000 420.6000 ;
	    RECT 88.2000 419.4000 89.4000 420.6000 ;
	    RECT 71.5500 402.6000 72.4500 419.4000 ;
	    RECT 64.2000 401.4000 65.4000 402.6000 ;
	    RECT 71.4000 401.4000 72.6000 402.6000 ;
	    RECT 64.3500 384.6000 65.2500 401.4000 ;
	    RECT 64.2000 383.4000 65.4000 384.6000 ;
	    RECT 66.6000 347.4000 67.8000 348.6000 ;
	    RECT 66.7500 345.6000 67.6500 347.4000 ;
	    RECT 66.6000 344.4000 67.8000 345.6000 ;
	    RECT 71.5500 342.6000 72.4500 401.4000 ;
	    RECT 88.2000 398.4000 89.4000 399.6000 ;
	    RECT 90.6000 398.4000 91.8000 399.6000 ;
	    RECT 88.3500 396.6000 89.2500 398.4000 ;
	    RECT 88.2000 395.4000 89.4000 396.6000 ;
	    RECT 47.4000 341.4000 48.6000 342.6000 ;
	    RECT 66.6000 341.4000 67.8000 342.6000 ;
	    RECT 71.4000 341.4000 72.6000 342.6000 ;
	    RECT 64.2000 329.4000 65.4000 330.6000 ;
	    RECT 64.3500 324.6000 65.2500 329.4000 ;
	    RECT 64.2000 323.4000 65.4000 324.6000 ;
	    RECT 47.4000 317.4000 48.6000 318.6000 ;
	    RECT 64.3500 231.6000 65.2500 323.4000 ;
	    RECT 66.7500 315.6000 67.6500 341.4000 ;
	    RECT 71.5500 336.6000 72.4500 341.4000 ;
	    RECT 73.8000 338.4000 75.0000 339.6000 ;
	    RECT 71.4000 335.4000 72.6000 336.6000 ;
	    RECT 73.9500 330.6000 74.8500 338.4000 ;
	    RECT 73.8000 329.4000 75.0000 330.6000 ;
	    RECT 73.8000 320.4000 75.0000 321.6000 ;
	    RECT 76.2000 320.4000 77.4000 321.6000 ;
	    RECT 73.9500 318.6000 74.8500 320.4000 ;
	    RECT 73.8000 317.4000 75.0000 318.6000 ;
	    RECT 66.6000 314.4000 67.8000 315.6000 ;
	    RECT 64.2000 230.4000 65.4000 231.6000 ;
	    RECT 71.4000 215.4000 72.6000 216.6000 ;
	    RECT 47.4000 200.4000 48.6000 201.6000 ;
	    RECT 54.6000 200.4000 55.8000 201.6000 ;
	    RECT 45.0000 194.4000 46.2000 195.6000 ;
	    RECT 47.5500 171.4500 48.4500 200.4000 ;
	    RECT 54.7500 198.6000 55.6500 200.4000 ;
	    RECT 54.6000 197.4000 55.8000 198.6000 ;
	    RECT 47.5500 170.5500 50.8500 171.4500 ;
	    RECT 40.2000 167.4000 41.4000 168.6000 ;
	    RECT 47.4000 167.4000 48.6000 168.6000 ;
	    RECT 33.0000 164.4000 34.2000 165.6000 ;
	    RECT 33.1500 162.6000 34.0500 164.4000 ;
	    RECT 16.2000 161.4000 17.4000 162.6000 ;
	    RECT 18.6000 161.4000 19.8000 162.6000 ;
	    RECT 33.0000 161.4000 34.2000 162.6000 ;
	    RECT 13.8000 158.4000 15.0000 159.6000 ;
	    RECT 13.9500 114.6000 14.8500 158.4000 ;
	    RECT 13.8000 113.4000 15.0000 114.6000 ;
	    RECT 18.7500 108.6000 19.6500 161.4000 ;
	    RECT 23.4000 113.4000 24.6000 114.6000 ;
	    RECT 18.6000 107.4000 19.8000 108.6000 ;
	    RECT 18.7500 102.6000 19.6500 107.4000 ;
	    RECT 23.5500 102.6000 24.4500 113.4000 ;
	    RECT 18.6000 101.4000 19.8000 102.6000 ;
	    RECT 23.4000 101.4000 24.6000 102.6000 ;
	    RECT 47.4000 101.4000 48.6000 102.6000 ;
	    RECT 23.5500 51.6000 24.4500 101.4000 ;
	    RECT 47.5500 84.6000 48.4500 101.4000 ;
	    RECT 47.4000 83.4000 48.6000 84.6000 ;
	    RECT 23.4000 50.4000 24.6000 51.6000 ;
	    RECT 49.9500 24.6000 50.8500 170.5500 ;
	    RECT 54.6000 101.4000 55.8000 102.6000 ;
	    RECT 71.5500 99.6000 72.4500 215.4000 ;
	    RECT 73.9500 204.6000 74.8500 317.4000 ;
	    RECT 76.3500 288.6000 77.2500 320.4000 ;
	    RECT 90.7500 318.6000 91.6500 398.4000 ;
	    RECT 105.1500 321.6000 106.0500 761.4000 ;
	    RECT 114.7500 648.6000 115.6500 773.4000 ;
	    RECT 121.9500 684.6000 122.8500 878.4000 ;
	    RECT 124.2000 869.4000 125.4000 870.6000 ;
	    RECT 124.3500 771.6000 125.2500 869.4000 ;
	    RECT 126.6000 863.4000 127.8000 864.6000 ;
	    RECT 126.7500 861.6000 127.6500 863.4000 ;
	    RECT 126.6000 860.4000 127.8000 861.6000 ;
	    RECT 126.6000 857.4000 127.8000 858.6000 ;
	    RECT 126.6000 830.4000 127.8000 831.6000 ;
	    RECT 126.7500 804.4500 127.6500 830.4000 ;
	    RECT 129.0000 804.4500 130.2000 804.6000 ;
	    RECT 126.7500 803.5500 130.2000 804.4500 ;
	    RECT 129.0000 803.4000 130.2000 803.5500 ;
	    RECT 124.2000 770.4000 125.4000 771.6000 ;
	    RECT 124.3500 720.6000 125.2500 770.4000 ;
	    RECT 124.2000 719.4000 125.4000 720.6000 ;
	    RECT 124.3500 714.6000 125.2500 719.4000 ;
	    RECT 124.2000 713.4000 125.4000 714.6000 ;
	    RECT 124.2000 701.4000 125.4000 702.6000 ;
	    RECT 121.8000 683.4000 123.0000 684.6000 ;
	    RECT 129.0000 680.4000 130.2000 681.6000 ;
	    RECT 114.6000 647.4000 115.8000 648.6000 ;
	    RECT 121.8000 644.4000 123.0000 645.6000 ;
	    RECT 119.4000 641.4000 120.6000 642.6000 ;
	    RECT 112.2000 638.4000 113.4000 639.6000 ;
	    RECT 112.3500 612.6000 113.2500 638.4000 ;
	    RECT 112.2000 611.4000 113.4000 612.6000 ;
	    RECT 107.4000 575.4000 108.6000 576.6000 ;
	    RECT 107.5500 558.6000 108.4500 575.4000 ;
	    RECT 117.0000 563.4000 118.2000 564.6000 ;
	    RECT 107.4000 557.4000 108.6000 558.6000 ;
	    RECT 117.1500 492.6000 118.0500 563.4000 ;
	    RECT 117.0000 491.4000 118.2000 492.6000 ;
	    RECT 117.1500 486.6000 118.0500 491.4000 ;
	    RECT 117.0000 485.4000 118.2000 486.6000 ;
	    RECT 119.4000 419.4000 120.6000 420.6000 ;
	    RECT 119.5500 402.6000 120.4500 419.4000 ;
	    RECT 119.4000 401.4000 120.6000 402.6000 ;
	    RECT 119.4000 398.4000 120.6000 399.6000 ;
	    RECT 119.5500 396.6000 120.4500 398.4000 ;
	    RECT 119.4000 395.4000 120.6000 396.6000 ;
	    RECT 107.4000 389.4000 108.6000 390.6000 ;
	    RECT 107.5500 342.6000 108.4500 389.4000 ;
	    RECT 121.9500 348.6000 122.8500 644.4000 ;
	    RECT 124.2000 638.4000 125.4000 639.6000 ;
	    RECT 124.3500 435.6000 125.2500 638.4000 ;
	    RECT 129.1500 561.6000 130.0500 680.4000 ;
	    RECT 131.5500 639.6000 132.4500 938.4000 ;
	    RECT 133.8000 926.4000 135.0000 927.6000 ;
	    RECT 133.9500 882.6000 134.8500 926.4000 ;
	    RECT 136.3500 906.6000 137.2500 977.4000 ;
	    RECT 138.6000 966.3000 139.8000 986.7000 ;
	    RECT 141.0000 966.3000 142.2000 986.7000 ;
	    RECT 143.4000 969.3000 144.6000 986.7000 ;
	    RECT 145.8000 980.4000 147.0000 981.6000 ;
	    RECT 145.9500 954.6000 146.8500 980.4000 ;
	    RECT 148.2000 969.3000 149.4000 986.7000 ;
	    RECT 150.7500 984.6000 151.6500 998.4000 ;
	    RECT 153.0000 996.3000 154.2000 1013.7000 ;
	    RECT 155.4000 996.3000 156.6000 1016.7000 ;
	    RECT 157.8000 996.3000 159.0000 1016.7000 ;
	    RECT 160.2000 996.3000 161.4000 1016.7000 ;
	    RECT 162.7500 990.6000 163.6500 1049.4000 ;
	    RECT 162.6000 989.4000 163.8000 990.6000 ;
	    RECT 150.6000 983.4000 151.8000 984.6000 ;
	    RECT 145.8000 953.4000 147.0000 954.6000 ;
	    RECT 138.6000 941.4000 139.8000 942.6000 ;
	    RECT 136.2000 905.4000 137.4000 906.6000 ;
	    RECT 133.8000 881.4000 135.0000 882.6000 ;
	    RECT 138.7500 819.4500 139.6500 941.4000 ;
	    RECT 150.7500 930.6000 151.6500 983.4000 ;
	    RECT 153.0000 969.3000 154.2000 986.7000 ;
	    RECT 153.0000 965.4000 154.2000 966.6000 ;
	    RECT 155.4000 966.3000 156.6000 986.7000 ;
	    RECT 157.8000 966.3000 159.0000 986.7000 ;
	    RECT 160.2000 966.3000 161.4000 986.7000 ;
	    RECT 162.6000 977.4000 163.8000 978.6000 ;
	    RECT 153.1500 948.6000 154.0500 965.4000 ;
	    RECT 153.0000 947.4000 154.2000 948.6000 ;
	    RECT 157.8000 944.4000 159.0000 945.6000 ;
	    RECT 150.6000 929.4000 151.8000 930.6000 ;
	    RECT 150.6000 893.4000 151.8000 894.6000 ;
	    RECT 141.0000 881.4000 142.2000 882.6000 ;
	    RECT 141.1500 879.6000 142.0500 881.4000 ;
	    RECT 141.0000 878.4000 142.2000 879.6000 ;
	    RECT 136.3500 818.5500 139.6500 819.4500 ;
	    RECT 136.3500 705.6000 137.2500 818.5500 ;
	    RECT 138.6000 815.4000 139.8000 816.6000 ;
	    RECT 141.0000 816.3000 142.2000 836.7000 ;
	    RECT 143.4000 816.3000 144.6000 836.7000 ;
	    RECT 145.8000 816.3000 147.0000 836.7000 ;
	    RECT 148.2000 816.3000 149.4000 833.7000 ;
	    RECT 150.7500 819.6000 151.6500 893.4000 ;
	    RECT 155.4000 881.4000 156.6000 882.6000 ;
	    RECT 153.0000 857.4000 154.2000 858.6000 ;
	    RECT 150.6000 818.4000 151.8000 819.6000 ;
	    RECT 136.2000 704.4000 137.4000 705.6000 ;
	    RECT 133.8000 683.4000 135.0000 684.6000 ;
	    RECT 131.4000 638.4000 132.6000 639.6000 ;
	    RECT 131.4000 614.4000 132.6000 615.6000 ;
	    RECT 131.5500 606.6000 132.4500 614.4000 ;
	    RECT 131.4000 605.4000 132.6000 606.6000 ;
	    RECT 131.4000 596.4000 132.6000 597.6000 ;
	    RECT 131.5500 588.6000 132.4500 596.4000 ;
	    RECT 133.9500 594.6000 134.8500 683.4000 ;
	    RECT 138.7500 657.6000 139.6500 815.4000 ;
	    RECT 141.0000 786.3000 142.2000 806.7000 ;
	    RECT 143.4000 786.3000 144.6000 806.7000 ;
	    RECT 145.8000 786.3000 147.0000 806.7000 ;
	    RECT 148.2000 789.3000 149.4000 806.7000 ;
	    RECT 150.7500 804.6000 151.6500 818.4000 ;
	    RECT 153.0000 816.3000 154.2000 833.7000 ;
	    RECT 155.5500 828.6000 156.4500 881.4000 ;
	    RECT 157.9500 855.6000 158.8500 944.4000 ;
	    RECT 162.7500 942.6000 163.6500 977.4000 ;
	    RECT 162.6000 941.4000 163.8000 942.6000 ;
	    RECT 162.6000 938.4000 163.8000 939.6000 ;
	    RECT 160.2000 860.4000 161.4000 861.6000 ;
	    RECT 160.3500 858.6000 161.2500 860.4000 ;
	    RECT 160.2000 857.4000 161.4000 858.6000 ;
	    RECT 157.8000 854.4000 159.0000 855.6000 ;
	    RECT 162.7500 843.4500 163.6500 938.4000 ;
	    RECT 165.1500 846.6000 166.0500 1073.4000 ;
	    RECT 167.4000 1037.4000 168.6000 1038.6000 ;
	    RECT 167.5500 1014.6000 168.4500 1037.4000 ;
	    RECT 167.4000 1013.4000 168.6000 1014.6000 ;
	    RECT 169.9500 939.6000 170.8500 1097.4000 ;
	    RECT 172.2000 1091.4000 173.4000 1092.6000 ;
	    RECT 172.3500 1086.6000 173.2500 1091.4000 ;
	    RECT 172.2000 1085.4000 173.4000 1086.6000 ;
	    RECT 172.2000 1070.4000 173.4000 1071.6000 ;
	    RECT 172.3500 1044.6000 173.2500 1070.4000 ;
	    RECT 177.0000 1055.4000 178.2000 1056.6000 ;
	    RECT 172.2000 1043.4000 173.4000 1044.6000 ;
	    RECT 172.3500 1002.6000 173.2500 1043.4000 ;
	    RECT 177.1500 1032.6000 178.0500 1055.4000 ;
	    RECT 177.0000 1031.4000 178.2000 1032.6000 ;
	    RECT 177.0000 1010.4000 178.2000 1011.6000 ;
	    RECT 172.2000 1001.4000 173.4000 1002.6000 ;
	    RECT 174.6000 971.4000 175.8000 972.6000 ;
	    RECT 174.7500 960.6000 175.6500 971.4000 ;
	    RECT 174.6000 959.4000 175.8000 960.6000 ;
	    RECT 177.1500 948.6000 178.0500 1010.4000 ;
	    RECT 179.5500 954.6000 180.4500 1118.4000 ;
	    RECT 191.4000 1085.4000 192.6000 1086.6000 ;
	    RECT 191.5500 1080.6000 192.4500 1085.4000 ;
	    RECT 191.4000 1079.4000 192.6000 1080.6000 ;
	    RECT 184.2000 1043.4000 185.4000 1044.6000 ;
	    RECT 184.3500 1041.6000 185.2500 1043.4000 ;
	    RECT 191.5500 1041.6000 192.4500 1079.4000 ;
	    RECT 181.8000 1040.4000 183.0000 1041.6000 ;
	    RECT 184.2000 1040.4000 185.4000 1041.6000 ;
	    RECT 191.4000 1040.4000 192.6000 1041.6000 ;
	    RECT 181.9500 1038.6000 182.8500 1040.4000 ;
	    RECT 181.8000 1037.4000 183.0000 1038.6000 ;
	    RECT 189.0000 1037.4000 190.2000 1038.6000 ;
	    RECT 191.4000 1037.4000 192.6000 1038.6000 ;
	    RECT 184.2000 1035.4501 185.4000 1035.6000 ;
	    RECT 191.5500 1035.4501 192.4500 1037.4000 ;
	    RECT 184.2000 1034.5500 192.4500 1035.4501 ;
	    RECT 184.2000 1034.4000 185.4000 1034.5500 ;
	    RECT 181.8000 1019.4000 183.0000 1020.6000 ;
	    RECT 179.4000 953.4000 180.6000 954.6000 ;
	    RECT 177.0000 947.4000 178.2000 948.6000 ;
	    RECT 179.4000 944.4000 180.6000 945.6000 ;
	    RECT 174.6000 941.4000 175.8000 942.6000 ;
	    RECT 169.8000 938.4000 171.0000 939.6000 ;
	    RECT 167.4000 888.4500 168.6000 888.6000 ;
	    RECT 167.4000 887.5500 170.8500 888.4500 ;
	    RECT 167.4000 887.4000 168.6000 887.5500 ;
	    RECT 167.4000 881.4000 168.6000 882.6000 ;
	    RECT 169.9500 876.6000 170.8500 887.5500 ;
	    RECT 174.7500 882.6000 175.6500 941.4000 ;
	    RECT 177.0000 884.4000 178.2000 885.6000 ;
	    RECT 174.6000 881.4000 175.8000 882.6000 ;
	    RECT 169.8000 875.4000 171.0000 876.6000 ;
	    RECT 174.6000 869.4000 175.8000 870.6000 ;
	    RECT 174.7500 864.6000 175.6500 869.4000 ;
	    RECT 174.6000 863.4000 175.8000 864.6000 ;
	    RECT 177.1500 861.6000 178.0500 884.4000 ;
	    RECT 177.0000 860.4000 178.2000 861.6000 ;
	    RECT 167.4000 857.4000 168.6000 858.6000 ;
	    RECT 165.0000 845.4000 166.2000 846.6000 ;
	    RECT 162.7500 842.5500 166.0500 843.4500 ;
	    RECT 155.4000 827.4000 156.6000 828.6000 ;
	    RECT 155.4000 821.4000 156.6000 822.6000 ;
	    RECT 157.8000 816.3000 159.0000 833.7000 ;
	    RECT 160.2000 816.3000 161.4000 836.7000 ;
	    RECT 162.6000 816.3000 163.8000 836.7000 ;
	    RECT 165.1500 825.6000 166.0500 842.5500 ;
	    RECT 165.0000 824.4000 166.2000 825.6000 ;
	    RECT 165.1500 816.6000 166.0500 824.4000 ;
	    RECT 165.0000 815.4000 166.2000 816.6000 ;
	    RECT 150.6000 803.4000 151.8000 804.6000 ;
	    RECT 141.0000 756.3000 142.2000 776.7000 ;
	    RECT 143.4000 756.3000 144.6000 776.7000 ;
	    RECT 145.8000 756.3000 147.0000 776.7000 ;
	    RECT 148.2000 756.3000 149.4000 773.7000 ;
	    RECT 150.7500 759.6000 151.6500 803.4000 ;
	    RECT 153.0000 789.3000 154.2000 806.7000 ;
	    RECT 155.4000 800.4000 156.6000 801.6000 ;
	    RECT 155.5500 798.6000 156.4500 800.4000 ;
	    RECT 155.4000 797.4000 156.6000 798.6000 ;
	    RECT 157.8000 789.3000 159.0000 806.7000 ;
	    RECT 160.2000 786.3000 161.4000 806.7000 ;
	    RECT 162.6000 786.3000 163.8000 806.7000 ;
	    RECT 165.0000 797.4000 166.2000 798.6000 ;
	    RECT 150.6000 758.4000 151.8000 759.6000 ;
	    RECT 141.0000 726.3000 142.2000 746.7000 ;
	    RECT 143.4000 726.3000 144.6000 746.7000 ;
	    RECT 145.8000 726.3000 147.0000 746.7000 ;
	    RECT 148.2000 729.3000 149.4000 746.7000 ;
	    RECT 150.7500 744.6000 151.6500 758.4000 ;
	    RECT 153.0000 756.3000 154.2000 773.7000 ;
	    RECT 155.4000 767.4000 156.6000 768.6000 ;
	    RECT 155.5500 762.6000 156.4500 767.4000 ;
	    RECT 155.4000 761.4000 156.6000 762.6000 ;
	    RECT 157.8000 756.3000 159.0000 773.7000 ;
	    RECT 160.2000 756.3000 161.4000 776.7000 ;
	    RECT 162.6000 756.3000 163.8000 776.7000 ;
	    RECT 167.5500 768.6000 168.4500 857.4000 ;
	    RECT 169.8000 836.4000 171.0000 837.6000 ;
	    RECT 169.9500 828.6000 170.8500 836.4000 ;
	    RECT 169.8000 827.4000 171.0000 828.6000 ;
	    RECT 174.6000 827.4000 175.8000 828.6000 ;
	    RECT 169.8000 794.4000 171.0000 795.6000 ;
	    RECT 169.9500 786.6000 170.8500 794.4000 ;
	    RECT 169.8000 785.4000 171.0000 786.6000 ;
	    RECT 169.8000 776.4000 171.0000 777.6000 ;
	    RECT 169.9500 768.6000 170.8500 776.4000 ;
	    RECT 167.4000 767.4000 168.6000 768.6000 ;
	    RECT 169.8000 767.4000 171.0000 768.6000 ;
	    RECT 165.0000 764.4000 166.2000 765.6000 ;
	    RECT 165.1500 756.6000 166.0500 764.4000 ;
	    RECT 165.0000 755.4000 166.2000 756.6000 ;
	    RECT 172.2000 755.4000 173.4000 756.6000 ;
	    RECT 150.6000 743.4000 151.8000 744.6000 ;
	    RECT 141.0000 713.4000 142.2000 714.6000 ;
	    RECT 141.1500 708.6000 142.0500 713.4000 ;
	    RECT 141.0000 707.4000 142.2000 708.6000 ;
	    RECT 148.2000 701.4000 149.4000 702.6000 ;
	    RECT 148.3500 696.6000 149.2500 701.4000 ;
	    RECT 148.2000 695.4000 149.4000 696.6000 ;
	    RECT 150.7500 678.6000 151.6500 743.4000 ;
	    RECT 153.0000 729.3000 154.2000 746.7000 ;
	    RECT 155.4000 740.4000 156.6000 741.6000 ;
	    RECT 155.5500 702.6000 156.4500 740.4000 ;
	    RECT 157.8000 729.3000 159.0000 746.7000 ;
	    RECT 157.8000 725.4000 159.0000 726.6000 ;
	    RECT 160.2000 726.3000 161.4000 746.7000 ;
	    RECT 162.6000 726.3000 163.8000 746.7000 ;
	    RECT 167.4000 743.4000 168.6000 744.6000 ;
	    RECT 165.0000 737.4000 166.2000 738.6000 ;
	    RECT 157.9500 723.4500 158.8500 725.4000 ;
	    RECT 157.9500 722.5500 161.2500 723.4500 ;
	    RECT 155.4000 701.4000 156.6000 702.6000 ;
	    RECT 155.4000 695.4000 156.6000 696.6000 ;
	    RECT 155.5500 681.6000 156.4500 695.4000 ;
	    RECT 155.4000 680.4000 156.6000 681.6000 ;
	    RECT 150.6000 677.4000 151.8000 678.6000 ;
	    RECT 153.0000 677.4000 154.2000 678.6000 ;
	    RECT 157.8000 677.4000 159.0000 678.6000 ;
	    RECT 138.6000 656.4000 139.8000 657.6000 ;
	    RECT 145.8000 635.4000 147.0000 636.6000 ;
	    RECT 136.2000 617.4000 137.4000 618.6000 ;
	    RECT 133.8000 593.4000 135.0000 594.6000 ;
	    RECT 131.4000 587.4000 132.6000 588.6000 ;
	    RECT 136.3500 585.6000 137.2500 617.4000 ;
	    RECT 138.6000 606.3000 139.8000 626.7000 ;
	    RECT 141.0000 606.3000 142.2000 626.7000 ;
	    RECT 143.4000 609.3000 144.6000 626.7000 ;
	    RECT 145.9500 621.6000 146.8500 635.4000 ;
	    RECT 145.8000 620.4000 147.0000 621.6000 ;
	    RECT 148.2000 609.3000 149.4000 626.7000 ;
	    RECT 150.7500 624.6000 151.6500 677.4000 ;
	    RECT 153.1500 672.6000 154.0500 677.4000 ;
	    RECT 153.0000 671.4000 154.2000 672.6000 ;
	    RECT 160.3500 636.6000 161.2500 722.5500 ;
	    RECT 162.6000 719.4000 163.8000 720.6000 ;
	    RECT 162.7500 684.6000 163.6500 719.4000 ;
	    RECT 167.5500 711.4500 168.4500 743.4000 ;
	    RECT 169.8000 734.4000 171.0000 735.6000 ;
	    RECT 169.9500 726.6000 170.8500 734.4000 ;
	    RECT 172.3500 726.6000 173.2500 755.4000 ;
	    RECT 169.8000 725.4000 171.0000 726.6000 ;
	    RECT 172.2000 725.4000 173.4000 726.6000 ;
	    RECT 165.1500 710.5500 168.4500 711.4500 ;
	    RECT 165.1500 705.6000 166.0500 710.5500 ;
	    RECT 167.5500 707.5500 173.2500 708.4500 ;
	    RECT 165.0000 704.4000 166.2000 705.6000 ;
	    RECT 167.5500 702.6000 168.4500 707.5500 ;
	    RECT 172.3500 705.6000 173.2500 707.5500 ;
	    RECT 169.8000 704.4000 171.0000 705.6000 ;
	    RECT 172.2000 704.4000 173.4000 705.6000 ;
	    RECT 169.9500 702.6000 170.8500 704.4000 ;
	    RECT 165.0000 701.4000 166.2000 702.6000 ;
	    RECT 167.4000 701.4000 168.6000 702.6000 ;
	    RECT 169.8000 701.4000 171.0000 702.6000 ;
	    RECT 172.2000 701.4000 173.4000 702.6000 ;
	    RECT 165.1500 699.4500 166.0500 701.4000 ;
	    RECT 172.3500 699.4500 173.2500 701.4000 ;
	    RECT 165.1500 698.5500 173.2500 699.4500 ;
	    RECT 169.8000 689.4000 171.0000 690.6000 ;
	    RECT 162.6000 683.4000 163.8000 684.6000 ;
	    RECT 162.6000 656.4000 163.8000 657.6000 ;
	    RECT 160.2000 635.4000 161.4000 636.6000 ;
	    RECT 150.6000 623.4000 151.8000 624.6000 ;
	    RECT 145.8000 599.4000 147.0000 600.6000 ;
	    RECT 136.2000 584.4000 137.4000 585.6000 ;
	    RECT 136.3500 582.6000 137.2500 584.4000 ;
	    RECT 136.2000 581.4000 137.4000 582.6000 ;
	    RECT 138.6000 576.3000 139.8000 596.7000 ;
	    RECT 141.0000 576.3000 142.2000 596.7000 ;
	    RECT 143.4000 576.3000 144.6000 593.7000 ;
	    RECT 145.9500 582.6000 146.8500 599.4000 ;
	    RECT 145.8000 581.4000 147.0000 582.6000 ;
	    RECT 148.2000 576.3000 149.4000 593.7000 ;
	    RECT 150.7500 579.6000 151.6500 623.4000 ;
	    RECT 153.0000 609.3000 154.2000 626.7000 ;
	    RECT 155.4000 606.3000 156.6000 626.7000 ;
	    RECT 157.8000 606.3000 159.0000 626.7000 ;
	    RECT 160.2000 606.3000 161.4000 626.7000 ;
	    RECT 150.6000 578.4000 151.8000 579.6000 ;
	    RECT 153.0000 576.3000 154.2000 593.7000 ;
	    RECT 155.4000 576.3000 156.6000 596.7000 ;
	    RECT 157.8000 576.3000 159.0000 596.7000 ;
	    RECT 160.2000 576.3000 161.4000 596.7000 ;
	    RECT 162.7500 573.4500 163.6500 656.4000 ;
	    RECT 167.4000 653.4000 168.6000 654.6000 ;
	    RECT 167.5500 645.6000 168.4500 653.4000 ;
	    RECT 167.4000 644.4000 168.6000 645.6000 ;
	    RECT 169.9500 642.6000 170.8500 689.4000 ;
	    RECT 174.7500 681.6000 175.6500 827.4000 ;
	    RECT 177.0000 758.4000 178.2000 759.6000 ;
	    RECT 177.1500 750.6000 178.0500 758.4000 ;
	    RECT 177.0000 749.4000 178.2000 750.6000 ;
	    RECT 177.0000 701.4000 178.2000 702.6000 ;
	    RECT 174.6000 680.4000 175.8000 681.6000 ;
	    RECT 177.1500 672.6000 178.0500 701.4000 ;
	    RECT 179.5500 684.6000 180.4500 944.4000 ;
	    RECT 181.9500 852.6000 182.8500 1019.4000 ;
	    RECT 191.4000 1001.4000 192.6000 1002.6000 ;
	    RECT 191.5500 999.6000 192.4500 1001.4000 ;
	    RECT 191.4000 998.4000 192.6000 999.6000 ;
	    RECT 189.0000 989.4000 190.2000 990.6000 ;
	    RECT 184.2000 953.4000 185.4000 954.6000 ;
	    RECT 181.8000 851.4000 183.0000 852.6000 ;
	    RECT 184.3500 849.4500 185.2500 953.4000 ;
	    RECT 181.9500 848.5500 185.2500 849.4500 ;
	    RECT 181.9500 759.6000 182.8500 848.5500 ;
	    RECT 184.2000 845.4000 185.4000 846.6000 ;
	    RECT 181.8000 758.4000 183.0000 759.6000 ;
	    RECT 179.4000 683.4000 180.6000 684.6000 ;
	    RECT 177.0000 671.4000 178.2000 672.6000 ;
	    RECT 179.5500 645.6000 180.4500 683.4000 ;
	    RECT 179.4000 644.4000 180.6000 645.6000 ;
	    RECT 169.8000 641.4000 171.0000 642.6000 ;
	    RECT 177.0000 641.4000 178.2000 642.6000 ;
	    RECT 169.8000 635.4000 171.0000 636.6000 ;
	    RECT 165.0000 581.4000 166.2000 582.6000 ;
	    RECT 160.3500 572.5500 163.6500 573.4500 ;
	    RECT 131.4000 563.4000 132.6000 564.6000 ;
	    RECT 129.0000 560.4000 130.2000 561.6000 ;
	    RECT 131.5500 558.6000 132.4500 563.4000 ;
	    RECT 131.4000 557.4000 132.6000 558.6000 ;
	    RECT 129.0000 536.4000 130.2000 537.6000 ;
	    RECT 129.1500 528.6000 130.0500 536.4000 ;
	    RECT 129.0000 527.4000 130.2000 528.6000 ;
	    RECT 131.5500 510.6000 132.4500 557.4000 ;
	    RECT 133.8000 527.4000 135.0000 528.6000 ;
	    RECT 133.9500 525.6000 134.8500 527.4000 ;
	    RECT 133.8000 524.4000 135.0000 525.6000 ;
	    RECT 136.2000 516.3000 137.4000 536.7000 ;
	    RECT 138.6000 516.3000 139.8000 536.7000 ;
	    RECT 141.0000 516.3000 142.2000 533.7000 ;
	    RECT 143.4000 533.4000 144.6000 534.6000 ;
	    RECT 143.5500 522.6000 144.4500 533.4000 ;
	    RECT 143.4000 521.4000 144.6000 522.6000 ;
	    RECT 145.8000 516.3000 147.0000 533.7000 ;
	    RECT 148.2000 518.4000 149.4000 519.6000 ;
	    RECT 148.3500 513.4500 149.2500 518.4000 ;
	    RECT 150.6000 516.3000 151.8000 533.7000 ;
	    RECT 153.0000 516.3000 154.2000 536.7000 ;
	    RECT 155.4000 516.3000 156.6000 536.7000 ;
	    RECT 157.8000 516.3000 159.0000 536.7000 ;
	    RECT 160.3500 528.6000 161.2500 572.5500 ;
	    RECT 162.6000 557.4000 163.8000 558.6000 ;
	    RECT 160.2000 527.4000 161.4000 528.6000 ;
	    RECT 148.3500 512.5500 151.6500 513.4500 ;
	    RECT 131.4000 509.4000 132.6000 510.6000 ;
	    RECT 136.2000 497.4000 137.4000 498.6000 ;
	    RECT 131.4000 494.4000 132.6000 495.6000 ;
	    RECT 131.5500 486.6000 132.4500 494.4000 ;
	    RECT 131.4000 485.4000 132.6000 486.6000 ;
	    RECT 138.6000 486.3000 139.8000 506.7000 ;
	    RECT 141.0000 486.3000 142.2000 506.7000 ;
	    RECT 143.4000 489.3000 144.6000 506.7000 ;
	    RECT 145.8000 503.4000 147.0000 504.6000 ;
	    RECT 145.9500 501.6000 146.8500 503.4000 ;
	    RECT 145.8000 500.4000 147.0000 501.6000 ;
	    RECT 148.2000 489.3000 149.4000 506.7000 ;
	    RECT 150.7500 504.6000 151.6500 512.5500 ;
	    RECT 150.6000 503.4000 151.8000 504.6000 ;
	    RECT 150.7500 486.4500 151.6500 503.4000 ;
	    RECT 153.0000 489.3000 154.2000 506.7000 ;
	    RECT 148.3500 485.5500 151.6500 486.4500 ;
	    RECT 155.4000 486.3000 156.6000 506.7000 ;
	    RECT 157.8000 486.3000 159.0000 506.7000 ;
	    RECT 160.2000 486.3000 161.4000 506.7000 ;
	    RECT 162.7500 498.6000 163.6500 557.4000 ;
	    RECT 162.6000 497.4000 163.8000 498.6000 ;
	    RECT 129.0000 476.4000 130.2000 477.6000 ;
	    RECT 129.1500 468.6000 130.0500 476.4000 ;
	    RECT 131.4000 473.4000 132.6000 474.6000 ;
	    RECT 129.0000 467.4000 130.2000 468.6000 ;
	    RECT 131.5500 447.4500 132.4500 473.4000 ;
	    RECT 133.8000 464.4000 135.0000 465.6000 ;
	    RECT 133.9500 462.6000 134.8500 464.4000 ;
	    RECT 133.8000 461.4000 135.0000 462.6000 ;
	    RECT 136.2000 456.3000 137.4000 476.7000 ;
	    RECT 138.6000 456.3000 139.8000 476.7000 ;
	    RECT 141.0000 456.3000 142.2000 473.7000 ;
	    RECT 143.4000 461.4000 144.6000 462.6000 ;
	    RECT 143.5500 456.6000 144.4500 461.4000 ;
	    RECT 143.4000 455.4000 144.6000 456.6000 ;
	    RECT 145.8000 456.3000 147.0000 473.7000 ;
	    RECT 148.3500 459.6000 149.2500 485.5500 ;
	    RECT 148.2000 458.4000 149.4000 459.6000 ;
	    RECT 129.1500 446.5500 132.4500 447.4500 ;
	    RECT 126.6000 440.4000 127.8000 441.6000 ;
	    RECT 124.2000 434.4000 125.4000 435.6000 ;
	    RECT 126.7500 414.6000 127.6500 440.4000 ;
	    RECT 129.1500 438.6000 130.0500 446.5500 ;
	    RECT 131.4000 443.4000 132.6000 444.6000 ;
	    RECT 131.5500 441.6000 132.4500 443.4000 ;
	    RECT 131.4000 440.4000 132.6000 441.6000 ;
	    RECT 136.2000 440.4000 137.4000 441.6000 ;
	    RECT 129.0000 437.4000 130.2000 438.6000 ;
	    RECT 126.6000 413.4000 127.8000 414.6000 ;
	    RECT 133.8000 413.4000 135.0000 414.6000 ;
	    RECT 131.4000 398.4000 132.6000 399.6000 ;
	    RECT 129.0000 374.4000 130.2000 375.6000 ;
	    RECT 129.1500 366.6000 130.0500 374.4000 ;
	    RECT 129.0000 365.4000 130.2000 366.6000 ;
	    RECT 121.8000 347.4000 123.0000 348.6000 ;
	    RECT 112.2000 344.4000 113.4000 345.6000 ;
	    RECT 112.3500 342.6000 113.2500 344.4000 ;
	    RECT 107.4000 341.4000 108.6000 342.6000 ;
	    RECT 109.8000 341.4000 111.0000 342.6000 ;
	    RECT 112.2000 341.4000 113.4000 342.6000 ;
	    RECT 117.0000 341.4000 118.2000 342.6000 ;
	    RECT 119.4000 341.4000 120.6000 342.6000 ;
	    RECT 109.9500 336.6000 110.8500 341.4000 ;
	    RECT 109.8000 335.4000 111.0000 336.6000 ;
	    RECT 105.0000 320.4000 106.2000 321.6000 ;
	    RECT 90.6000 317.4000 91.8000 318.6000 ;
	    RECT 76.2000 287.4000 77.4000 288.6000 ;
	    RECT 73.8000 203.4000 75.0000 204.6000 ;
	    RECT 71.4000 98.4000 72.6000 99.6000 ;
	    RECT 49.8000 23.4000 51.0000 24.6000 ;
	    RECT 73.9500 12.6000 74.8500 203.4000 ;
	    RECT 93.0000 200.4000 94.2000 201.6000 ;
	    RECT 102.6000 200.4000 103.8000 201.6000 ;
	    RECT 93.1500 144.6000 94.0500 200.4000 ;
	    RECT 102.7500 198.6000 103.6500 200.4000 ;
	    RECT 102.6000 197.4000 103.8000 198.6000 ;
	    RECT 95.4000 194.4000 96.6000 195.6000 ;
	    RECT 95.5500 192.6000 96.4500 194.4000 ;
	    RECT 95.4000 191.4000 96.6000 192.6000 ;
	    RECT 117.1500 162.6000 118.0500 341.4000 ;
	    RECT 129.0000 254.4000 130.2000 255.6000 ;
	    RECT 129.1500 246.6000 130.0500 254.4000 ;
	    RECT 129.0000 245.4000 130.2000 246.6000 ;
	    RECT 131.5500 204.6000 132.4500 398.4000 ;
	    RECT 133.9500 378.6000 134.8500 413.4000 ;
	    RECT 136.3500 402.6000 137.2500 440.4000 ;
	    RECT 148.3500 408.6000 149.2500 458.4000 ;
	    RECT 150.6000 456.3000 151.8000 473.7000 ;
	    RECT 153.0000 456.3000 154.2000 476.7000 ;
	    RECT 155.4000 456.3000 156.6000 476.7000 ;
	    RECT 157.8000 456.3000 159.0000 476.7000 ;
	    RECT 162.6000 449.4000 163.8000 450.6000 ;
	    RECT 162.7500 444.6000 163.6500 449.4000 ;
	    RECT 162.6000 443.4000 163.8000 444.6000 ;
	    RECT 160.2000 440.4000 161.4000 441.6000 ;
	    RECT 148.2000 407.4000 149.4000 408.6000 ;
	    RECT 136.2000 401.4000 137.4000 402.6000 ;
	    RECT 133.8000 377.4000 135.0000 378.6000 ;
	    RECT 133.9500 258.6000 134.8500 377.4000 ;
	    RECT 136.2000 366.3000 137.4000 386.7000 ;
	    RECT 138.6000 366.3000 139.8000 386.7000 ;
	    RECT 141.0000 369.3000 142.2000 386.7000 ;
	    RECT 143.4000 383.4000 144.6000 384.6000 ;
	    RECT 143.5500 381.6000 144.4500 383.4000 ;
	    RECT 143.4000 380.4000 144.6000 381.6000 ;
	    RECT 145.8000 369.3000 147.0000 386.7000 ;
	    RECT 148.3500 384.6000 149.2500 407.4000 ;
	    RECT 160.3500 390.6000 161.2500 440.4000 ;
	    RECT 162.6000 437.4000 163.8000 438.6000 ;
	    RECT 162.7500 426.6000 163.6500 437.4000 ;
	    RECT 162.6000 425.4000 163.8000 426.6000 ;
	    RECT 165.1500 414.6000 166.0500 581.4000 ;
	    RECT 169.9500 462.6000 170.8500 635.4000 ;
	    RECT 177.1500 621.6000 178.0500 641.4000 ;
	    RECT 177.0000 620.4000 178.2000 621.6000 ;
	    RECT 174.6000 611.4000 175.8000 612.6000 ;
	    RECT 174.6000 593.4000 175.8000 594.6000 ;
	    RECT 174.7500 591.6000 175.6500 593.4000 ;
	    RECT 174.6000 590.4000 175.8000 591.6000 ;
	    RECT 181.8000 587.4000 183.0000 588.6000 ;
	    RECT 177.0000 581.4000 178.2000 582.6000 ;
	    RECT 177.1500 576.6000 178.0500 581.4000 ;
	    RECT 181.9500 576.6000 182.8500 587.4000 ;
	    RECT 184.3500 582.6000 185.2500 845.4000 ;
	    RECT 189.1500 834.6000 190.0500 989.4000 ;
	    RECT 191.4000 977.4000 192.6000 978.6000 ;
	    RECT 191.5500 945.6000 192.4500 977.4000 ;
	    RECT 191.4000 944.4000 192.6000 945.6000 ;
	    RECT 191.4000 941.4000 192.6000 942.6000 ;
	    RECT 191.5500 927.6000 192.4500 941.4000 ;
	    RECT 191.4000 926.4000 192.6000 927.6000 ;
	    RECT 193.9500 912.4500 194.8500 1127.4000 ;
	    RECT 196.3500 1104.6000 197.2500 1154.4000 ;
	    RECT 196.2000 1103.4000 197.4000 1104.6000 ;
	    RECT 196.2000 1100.4000 197.4000 1101.6000 ;
	    RECT 196.3500 1062.6000 197.2500 1100.4000 ;
	    RECT 198.7500 1068.6000 199.6500 1220.4000 ;
	    RECT 217.9500 1155.6000 218.8500 1373.4000 ;
	    RECT 220.3500 1362.6000 221.2500 1400.4000 ;
	    RECT 225.1500 1365.6000 226.0500 1454.4000 ;
	    RECT 232.3500 1401.6000 233.2500 1457.4000 ;
	    RECT 251.4000 1454.4000 252.6000 1455.6000 ;
	    RECT 251.5500 1452.6000 252.4500 1454.4000 ;
	    RECT 265.9500 1452.6000 266.8500 1457.4000 ;
	    RECT 251.4000 1451.4000 252.6000 1452.6000 ;
	    RECT 265.8000 1451.4000 267.0000 1452.6000 ;
	    RECT 237.0000 1430.4000 238.2000 1431.6000 ;
	    RECT 232.2000 1400.4000 233.4000 1401.6000 ;
	    RECT 237.1500 1395.6000 238.0500 1430.4000 ;
	    RECT 237.0000 1394.4000 238.2000 1395.6000 ;
	    RECT 234.6000 1385.4000 235.8000 1386.6000 ;
	    RECT 225.0000 1364.4000 226.2000 1365.6000 ;
	    RECT 220.2000 1361.4000 221.4000 1362.6000 ;
	    RECT 232.2000 1307.4000 233.4000 1308.6000 ;
	    RECT 229.8000 1301.4000 231.0000 1302.6000 ;
	    RECT 232.2000 1301.4000 233.4000 1302.6000 ;
	    RECT 232.3500 1272.6000 233.2500 1301.4000 ;
	    RECT 232.2000 1271.4000 233.4000 1272.6000 ;
	    RECT 222.6000 1160.4000 223.8000 1161.6000 ;
	    RECT 222.7500 1158.6000 223.6500 1160.4000 ;
	    RECT 222.6000 1157.4000 223.8000 1158.6000 ;
	    RECT 217.8000 1154.4000 219.0000 1155.6000 ;
	    RECT 222.7500 1122.6000 223.6500 1157.4000 ;
	    RECT 229.8000 1139.4000 231.0000 1140.6000 ;
	    RECT 229.9500 1128.6000 230.8500 1139.4000 ;
	    RECT 229.8000 1127.4000 231.0000 1128.6000 ;
	    RECT 234.7500 1125.6000 235.6500 1385.4000 ;
	    RECT 244.2000 1367.4000 245.4000 1368.6000 ;
	    RECT 241.8000 1361.4000 243.0000 1362.6000 ;
	    RECT 237.0000 1304.4000 238.2000 1305.6000 ;
	    RECT 237.1500 1302.6000 238.0500 1304.4000 ;
	    RECT 237.0000 1301.4000 238.2000 1302.6000 ;
	    RECT 239.4000 1301.4000 240.6000 1302.6000 ;
	    RECT 239.5500 1290.6000 240.4500 1301.4000 ;
	    RECT 239.4000 1289.4000 240.6000 1290.6000 ;
	    RECT 241.9500 1284.6000 242.8500 1361.4000 ;
	    RECT 244.3500 1332.6000 245.2500 1367.4000 ;
	    RECT 244.2000 1331.4000 245.4000 1332.6000 ;
	    RECT 244.3500 1299.6000 245.2500 1331.4000 ;
	    RECT 244.2000 1298.4000 245.4000 1299.6000 ;
	    RECT 241.8000 1283.4000 243.0000 1284.6000 ;
	    RECT 239.4000 1199.4000 240.6000 1200.6000 ;
	    RECT 237.0000 1196.4000 238.2000 1197.6000 ;
	    RECT 234.6000 1124.4000 235.8000 1125.6000 ;
	    RECT 222.6000 1121.4000 223.8000 1122.6000 ;
	    RECT 229.8000 1121.4000 231.0000 1122.6000 ;
	    RECT 232.2000 1121.4000 233.4000 1122.6000 ;
	    RECT 210.6000 1103.4000 211.8000 1104.6000 ;
	    RECT 220.2000 1097.4000 221.4000 1098.6000 ;
	    RECT 198.6000 1067.4000 199.8000 1068.6000 ;
	    RECT 220.3500 1065.6000 221.2500 1097.4000 ;
	    RECT 222.7500 1086.6000 223.6500 1121.4000 ;
	    RECT 229.9500 1116.6000 230.8500 1121.4000 ;
	    RECT 229.8000 1115.4000 231.0000 1116.6000 ;
	    RECT 232.2000 1103.4000 233.4000 1104.6000 ;
	    RECT 225.0000 1100.4000 226.2000 1101.6000 ;
	    RECT 222.6000 1085.4000 223.8000 1086.6000 ;
	    RECT 222.6000 1067.4000 223.8000 1068.6000 ;
	    RECT 215.4000 1064.4000 216.6000 1065.6000 ;
	    RECT 220.2000 1064.4000 221.4000 1065.6000 ;
	    RECT 196.2000 1061.4000 197.4000 1062.6000 ;
	    RECT 196.2000 1037.4000 197.4000 1038.6000 ;
	    RECT 196.3500 942.6000 197.2500 1037.4000 ;
	    RECT 210.6000 1001.4000 211.8000 1002.6000 ;
	    RECT 210.7500 981.6000 211.6500 1001.4000 ;
	    RECT 210.6000 980.4000 211.8000 981.6000 ;
	    RECT 198.6000 953.4000 199.8000 954.6000 ;
	    RECT 198.7500 945.6000 199.6500 953.4000 ;
	    RECT 198.6000 944.4000 199.8000 945.6000 ;
	    RECT 196.2000 941.4000 197.4000 942.6000 ;
	    RECT 196.2000 912.4500 197.4000 912.6000 ;
	    RECT 193.9500 911.5500 197.4000 912.4500 ;
	    RECT 196.2000 911.4000 197.4000 911.5500 ;
	    RECT 189.0000 834.4500 190.2000 834.6000 ;
	    RECT 189.0000 833.5500 192.4500 834.4500 ;
	    RECT 189.0000 833.4000 190.2000 833.5500 ;
	    RECT 189.0000 821.4000 190.2000 822.6000 ;
	    RECT 186.6000 803.4000 187.8000 804.6000 ;
	    RECT 189.1500 708.6000 190.0500 821.4000 ;
	    RECT 191.5500 774.6000 192.4500 833.5500 ;
	    RECT 191.4000 773.4000 192.6000 774.6000 ;
	    RECT 196.3500 756.6000 197.2500 911.4000 ;
	    RECT 198.7500 897.6000 199.6500 944.4000 ;
	    RECT 215.5500 942.6000 216.4500 1064.4000 ;
	    RECT 222.7500 1062.6000 223.6500 1067.4000 ;
	    RECT 217.8000 1061.4000 219.0000 1062.6000 ;
	    RECT 222.6000 1061.4000 223.8000 1062.6000 ;
	    RECT 217.9500 1059.4501 218.8500 1061.4000 ;
	    RECT 217.9500 1058.5500 221.2500 1059.4501 ;
	    RECT 217.8000 1055.4000 219.0000 1056.6000 ;
	    RECT 217.9500 1050.6000 218.8500 1055.4000 ;
	    RECT 217.8000 1049.4000 219.0000 1050.6000 ;
	    RECT 220.3500 1032.6000 221.2500 1058.5500 ;
	    RECT 222.6000 1055.4000 223.8000 1056.6000 ;
	    RECT 222.7500 1035.6000 223.6500 1055.4000 ;
	    RECT 222.6000 1034.4000 223.8000 1035.6000 ;
	    RECT 220.2000 1031.4000 221.4000 1032.6000 ;
	    RECT 225.1500 1002.6000 226.0500 1100.4000 ;
	    RECT 232.3500 1068.6000 233.2500 1103.4000 ;
	    RECT 232.2000 1067.4000 233.4000 1068.6000 ;
	    RECT 227.4000 1061.4000 228.6000 1062.6000 ;
	    RECT 232.2000 1061.4000 233.4000 1062.6000 ;
	    RECT 225.0000 1001.4000 226.2000 1002.6000 ;
	    RECT 222.6000 995.4000 223.8000 996.6000 ;
	    RECT 217.8000 989.4000 219.0000 990.6000 ;
	    RECT 217.9500 978.6000 218.8500 989.4000 ;
	    RECT 220.2000 980.4000 221.4000 981.6000 ;
	    RECT 217.8000 977.4000 219.0000 978.6000 ;
	    RECT 220.3500 972.6000 221.2500 980.4000 ;
	    RECT 222.7500 978.6000 223.6500 995.4000 ;
	    RECT 227.5500 981.6000 228.4500 1061.4000 ;
	    RECT 229.8000 1037.4000 231.0000 1038.6000 ;
	    RECT 232.3500 1005.6000 233.2500 1061.4000 ;
	    RECT 237.1500 1056.4501 238.0500 1196.4000 ;
	    RECT 239.5500 1101.6000 240.4500 1199.4000 ;
	    RECT 241.9500 1182.6000 242.8500 1283.4000 ;
	    RECT 251.5500 1224.6000 252.4500 1451.4000 ;
	    RECT 268.3500 1431.6000 269.2500 1463.4000 ;
	    RECT 294.6000 1460.4000 295.8000 1461.6000 ;
	    RECT 304.2000 1460.4000 305.4000 1461.6000 ;
	    RECT 385.8000 1460.4000 387.0000 1461.6000 ;
	    RECT 270.6000 1457.4000 271.8000 1458.6000 ;
	    RECT 292.2000 1457.4000 293.4000 1458.6000 ;
	    RECT 294.7500 1458.4501 295.6500 1460.4000 ;
	    RECT 304.3500 1458.6000 305.2500 1460.4000 ;
	    RECT 301.8000 1458.4501 303.0000 1458.6000 ;
	    RECT 294.7500 1457.5500 303.0000 1458.4501 ;
	    RECT 301.8000 1457.4000 303.0000 1457.5500 ;
	    RECT 304.2000 1457.4000 305.4000 1458.6000 ;
	    RECT 268.2000 1430.4000 269.4000 1431.6000 ;
	    RECT 270.7500 1401.6000 271.6500 1457.4000 ;
	    RECT 292.3500 1434.6000 293.2500 1457.4000 ;
	    RECT 297.0000 1454.4000 298.2000 1455.6000 ;
	    RECT 297.1500 1452.6000 298.0500 1454.4000 ;
	    RECT 297.0000 1451.4000 298.2000 1452.6000 ;
	    RECT 292.2000 1433.4000 293.4000 1434.6000 ;
	    RECT 280.2000 1430.4000 281.4000 1431.6000 ;
	    RECT 280.3500 1404.6000 281.2500 1430.4000 ;
	    RECT 311.4000 1421.4000 312.6000 1422.6000 ;
	    RECT 311.5500 1404.6000 312.4500 1421.4000 ;
	    RECT 323.4000 1416.3000 324.6000 1436.7001 ;
	    RECT 325.8000 1416.3000 327.0000 1436.7001 ;
	    RECT 328.2000 1416.3000 329.4000 1436.7001 ;
	    RECT 330.6000 1416.3000 331.8000 1433.7001 ;
	    RECT 333.0000 1418.4000 334.2000 1419.6000 ;
	    RECT 316.2000 1409.4000 317.4000 1410.6000 ;
	    RECT 316.3500 1404.6000 317.2500 1409.4000 ;
	    RECT 280.2000 1403.4000 281.4000 1404.6000 ;
	    RECT 311.4000 1403.4000 312.6000 1404.6000 ;
	    RECT 316.2000 1403.4000 317.4000 1404.6000 ;
	    RECT 330.6000 1403.4000 331.8000 1404.6000 ;
	    RECT 261.0000 1400.4000 262.2000 1401.6000 ;
	    RECT 270.6000 1400.4000 271.8000 1401.6000 ;
	    RECT 282.6000 1400.4000 283.8000 1401.6000 ;
	    RECT 285.0000 1400.4000 286.2000 1401.6000 ;
	    RECT 261.1500 1380.6000 262.0500 1400.4000 ;
	    RECT 265.8000 1397.4000 267.0000 1398.6000 ;
	    RECT 261.0000 1379.4000 262.2000 1380.6000 ;
	    RECT 263.4000 1331.4000 264.6000 1332.6000 ;
	    RECT 261.0000 1259.4000 262.2000 1260.6000 ;
	    RECT 253.8000 1241.4000 255.0000 1242.6000 ;
	    RECT 251.4000 1223.4000 252.6000 1224.6000 ;
	    RECT 253.9500 1221.6000 254.8500 1241.4000 ;
	    RECT 258.6000 1235.4000 259.8000 1236.6000 ;
	    RECT 249.0000 1220.4000 250.2000 1221.6000 ;
	    RECT 253.8000 1220.4000 255.0000 1221.6000 ;
	    RECT 256.2000 1220.4000 257.4000 1221.6000 ;
	    RECT 246.6000 1217.4000 247.8000 1218.6000 ;
	    RECT 246.7500 1212.6000 247.6500 1217.4000 ;
	    RECT 246.6000 1211.4000 247.8000 1212.6000 ;
	    RECT 246.7500 1197.6000 247.6500 1211.4000 ;
	    RECT 246.6000 1196.4000 247.8000 1197.6000 ;
	    RECT 246.6000 1193.4000 247.8000 1194.6000 ;
	    RECT 241.8000 1181.4000 243.0000 1182.6000 ;
	    RECT 239.4000 1100.4000 240.6000 1101.6000 ;
	    RECT 239.4000 1073.4000 240.6000 1074.6000 ;
	    RECT 239.5500 1059.6000 240.4500 1073.4000 ;
	    RECT 239.4000 1058.4000 240.6000 1059.6000 ;
	    RECT 237.1500 1055.5500 240.4500 1056.4501 ;
	    RECT 234.6000 1019.4000 235.8000 1020.6000 ;
	    RECT 232.2000 1004.4000 233.4000 1005.6000 ;
	    RECT 227.4000 980.4000 228.6000 981.6000 ;
	    RECT 222.6000 977.4000 223.8000 978.6000 ;
	    RECT 220.2000 971.4000 221.4000 972.6000 ;
	    RECT 222.7500 954.6000 223.6500 977.4000 ;
	    RECT 222.6000 953.4000 223.8000 954.6000 ;
	    RECT 215.4000 941.4000 216.6000 942.6000 ;
	    RECT 232.3500 936.6000 233.2500 1004.4000 ;
	    RECT 234.7500 996.6000 235.6500 1019.4000 ;
	    RECT 239.5500 1005.6000 240.4500 1055.5500 ;
	    RECT 239.4000 1004.4000 240.6000 1005.6000 ;
	    RECT 237.0000 1001.4000 238.2000 1002.6000 ;
	    RECT 234.6000 995.4000 235.8000 996.6000 ;
	    RECT 237.1500 984.6000 238.0500 1001.4000 ;
	    RECT 237.0000 983.4000 238.2000 984.6000 ;
	    RECT 232.2000 935.4000 233.4000 936.6000 ;
	    RECT 213.0000 917.4000 214.2000 918.6000 ;
	    RECT 208.2000 914.4000 209.4000 915.6000 ;
	    RECT 208.3500 906.6000 209.2500 914.4000 ;
	    RECT 213.1500 912.6000 214.0500 917.4000 ;
	    RECT 213.0000 911.4000 214.2000 912.6000 ;
	    RECT 208.2000 905.4000 209.4000 906.6000 ;
	    RECT 215.4000 906.3000 216.6000 926.7000 ;
	    RECT 217.8000 906.3000 219.0000 926.7000 ;
	    RECT 220.2000 909.3000 221.4000 926.7000 ;
	    RECT 222.6000 920.4000 223.8000 921.6000 ;
	    RECT 198.6000 896.4000 199.8000 897.6000 ;
	    RECT 222.7500 882.6000 223.6500 920.4000 ;
	    RECT 225.0000 909.3000 226.2000 926.7000 ;
	    RECT 227.4000 923.4000 228.6000 924.6000 ;
	    RECT 225.0000 905.4000 226.2000 906.6000 ;
	    RECT 225.1500 888.6000 226.0500 905.4000 ;
	    RECT 227.5500 894.6000 228.4500 923.4000 ;
	    RECT 229.8000 909.3000 231.0000 926.7000 ;
	    RECT 232.2000 906.3000 233.4000 926.7000 ;
	    RECT 234.6000 906.3000 235.8000 926.7000 ;
	    RECT 237.0000 906.3000 238.2000 926.7000 ;
	    RECT 239.5500 906.6000 240.4500 1004.4000 ;
	    RECT 239.4000 905.4000 240.6000 906.6000 ;
	    RECT 237.0000 896.4000 238.2000 897.6000 ;
	    RECT 227.4000 893.4000 228.6000 894.6000 ;
	    RECT 225.0000 887.4000 226.2000 888.6000 ;
	    RECT 222.6000 881.4000 223.8000 882.6000 ;
	    RECT 227.4000 881.4000 228.6000 882.6000 ;
	    RECT 217.8000 875.4000 219.0000 876.6000 ;
	    RECT 210.6000 863.4000 211.8000 864.6000 ;
	    RECT 215.4000 863.4000 216.6000 864.6000 ;
	    RECT 213.0000 860.4000 214.2000 861.6000 ;
	    RECT 213.1500 822.6000 214.0500 860.4000 ;
	    RECT 217.9500 858.6000 218.8500 875.4000 ;
	    RECT 227.5500 861.6000 228.4500 881.4000 ;
	    RECT 227.4000 860.4000 228.6000 861.6000 ;
	    RECT 217.8000 857.4000 219.0000 858.6000 ;
	    RECT 220.2000 857.4000 221.4000 858.6000 ;
	    RECT 215.4000 851.4000 216.6000 852.6000 ;
	    RECT 215.5500 825.6000 216.4500 851.4000 ;
	    RECT 220.3500 825.6000 221.2500 857.4000 ;
	    RECT 222.6000 827.4000 223.8000 828.6000 ;
	    RECT 215.4000 824.4000 216.6000 825.6000 ;
	    RECT 220.2000 824.4000 221.4000 825.6000 ;
	    RECT 213.0000 821.4000 214.2000 822.6000 ;
	    RECT 203.4000 803.4000 204.6000 804.6000 ;
	    RECT 210.6000 803.4000 211.8000 804.6000 ;
	    RECT 203.5500 786.6000 204.4500 803.4000 ;
	    RECT 210.7500 801.6000 211.6500 803.4000 ;
	    RECT 210.6000 800.4000 211.8000 801.6000 ;
	    RECT 203.4000 785.4000 204.6000 786.6000 ;
	    RECT 196.2000 755.4000 197.4000 756.6000 ;
	    RECT 193.8000 749.4000 195.0000 750.6000 ;
	    RECT 193.9500 744.6000 194.8500 749.4000 ;
	    RECT 193.8000 743.4000 195.0000 744.6000 ;
	    RECT 215.5500 741.4500 216.4500 824.4000 ;
	    RECT 217.8000 821.4000 219.0000 822.6000 ;
	    RECT 217.9500 750.6000 218.8500 821.4000 ;
	    RECT 217.8000 749.4000 219.0000 750.6000 ;
	    RECT 215.5500 740.5500 218.8500 741.4500 ;
	    RECT 215.4000 737.4000 216.6000 738.6000 ;
	    RECT 191.4000 714.4500 192.6000 714.6000 ;
	    RECT 191.4000 713.5500 194.8500 714.4500 ;
	    RECT 191.4000 713.4000 192.6000 713.5500 ;
	    RECT 193.9500 708.6000 194.8500 713.5500 ;
	    RECT 205.8000 713.4000 207.0000 714.6000 ;
	    RECT 205.9500 708.6000 206.8500 713.4000 ;
	    RECT 189.0000 708.4500 190.2000 708.6000 ;
	    RECT 186.7500 707.5500 190.2000 708.4500 ;
	    RECT 184.2000 581.4000 185.4000 582.6000 ;
	    RECT 177.0000 575.4000 178.2000 576.6000 ;
	    RECT 181.8000 575.4000 183.0000 576.6000 ;
	    RECT 174.6000 509.4000 175.8000 510.6000 ;
	    RECT 174.7500 492.6000 175.6500 509.4000 ;
	    RECT 184.2000 503.4000 185.4000 504.6000 ;
	    RECT 177.0000 497.4000 178.2000 498.6000 ;
	    RECT 174.6000 491.4000 175.8000 492.6000 ;
	    RECT 172.2000 485.4000 173.4000 486.6000 ;
	    RECT 172.3500 471.6000 173.2500 485.4000 ;
	    RECT 172.2000 470.4000 173.4000 471.6000 ;
	    RECT 169.8000 461.4000 171.0000 462.6000 ;
	    RECT 169.8000 443.4000 171.0000 444.6000 ;
	    RECT 169.9500 441.6000 170.8500 443.4000 ;
	    RECT 169.8000 440.4000 171.0000 441.6000 ;
	    RECT 174.6000 440.4000 175.8000 441.6000 ;
	    RECT 167.4000 437.4000 168.6000 438.6000 ;
	    RECT 167.5500 417.6000 168.4500 437.4000 ;
	    RECT 174.7500 420.6000 175.6500 440.4000 ;
	    RECT 174.6000 419.4000 175.8000 420.6000 ;
	    RECT 167.4000 416.4000 168.6000 417.6000 ;
	    RECT 165.0000 413.4000 166.2000 414.6000 ;
	    RECT 172.2000 395.4000 173.4000 396.6000 ;
	    RECT 160.2000 389.4000 161.4000 390.6000 ;
	    RECT 148.2000 383.4000 149.4000 384.6000 ;
	    RECT 138.6000 341.4000 139.8000 342.6000 ;
	    RECT 138.7500 336.6000 139.6500 341.4000 ;
	    RECT 138.6000 335.4000 139.8000 336.6000 ;
	    RECT 143.4000 329.4000 144.6000 330.6000 ;
	    RECT 141.0000 323.4000 142.2000 324.6000 ;
	    RECT 141.1500 276.6000 142.0500 323.4000 ;
	    RECT 143.5500 321.6000 144.4500 329.4000 ;
	    RECT 143.4000 320.4000 144.6000 321.6000 ;
	    RECT 148.3500 294.6000 149.2500 383.4000 ;
	    RECT 150.6000 369.3000 151.8000 386.7000 ;
	    RECT 153.0000 366.3000 154.2000 386.7000 ;
	    RECT 155.4000 366.3000 156.6000 386.7000 ;
	    RECT 157.8000 366.3000 159.0000 386.7000 ;
	    RECT 172.3500 372.6000 173.2500 395.4000 ;
	    RECT 174.6000 377.4000 175.8000 378.6000 ;
	    RECT 172.2000 371.4000 173.4000 372.6000 ;
	    RECT 174.7500 360.6000 175.6500 377.4000 ;
	    RECT 160.2000 359.4000 161.4000 360.6000 ;
	    RECT 174.6000 359.4000 175.8000 360.6000 ;
	    RECT 160.3500 348.6000 161.2500 359.4000 ;
	    RECT 160.2000 347.4000 161.4000 348.6000 ;
	    RECT 160.2000 341.4000 161.4000 342.6000 ;
	    RECT 167.4000 341.4000 168.6000 342.6000 ;
	    RECT 157.8000 338.4000 159.0000 339.6000 ;
	    RECT 157.9500 324.6000 158.8500 338.4000 ;
	    RECT 157.8000 323.4000 159.0000 324.6000 ;
	    RECT 148.2000 293.4000 149.4000 294.6000 ;
	    RECT 143.4000 281.4000 144.6000 282.6000 ;
	    RECT 141.0000 275.4000 142.2000 276.6000 ;
	    RECT 133.8000 257.4000 135.0000 258.6000 ;
	    RECT 133.9500 246.6000 134.8500 257.4000 ;
	    RECT 133.8000 245.4000 135.0000 246.6000 ;
	    RECT 136.2000 246.3000 137.4000 266.7000 ;
	    RECT 138.6000 246.3000 139.8000 266.7000 ;
	    RECT 141.0000 249.3000 142.2000 266.7000 ;
	    RECT 143.5500 261.6000 144.4500 281.4000 ;
	    RECT 143.4000 260.4000 144.6000 261.6000 ;
	    RECT 145.8000 249.3000 147.0000 266.7000 ;
	    RECT 148.3500 264.6000 149.2500 293.4000 ;
	    RECT 160.3500 282.6000 161.2500 341.4000 ;
	    RECT 165.0000 323.4000 166.2000 324.6000 ;
	    RECT 174.6000 323.4000 175.8000 324.6000 ;
	    RECT 162.6000 287.4000 163.8000 288.6000 ;
	    RECT 160.2000 281.4000 161.4000 282.6000 ;
	    RECT 148.2000 263.4000 149.4000 264.6000 ;
	    RECT 150.6000 249.3000 151.8000 266.7000 ;
	    RECT 153.0000 246.3000 154.2000 266.7000 ;
	    RECT 155.4000 246.3000 156.6000 266.7000 ;
	    RECT 157.8000 246.3000 159.0000 266.7000 ;
	    RECT 162.7500 252.6000 163.6500 287.4000 ;
	    RECT 162.6000 251.4000 163.8000 252.6000 ;
	    RECT 131.4000 203.4000 132.6000 204.6000 ;
	    RECT 124.2000 200.4000 125.4000 201.6000 ;
	    RECT 124.3500 198.6000 125.2500 200.4000 ;
	    RECT 119.4000 197.4000 120.6000 198.6000 ;
	    RECT 124.2000 197.4000 125.4000 198.6000 ;
	    RECT 119.5500 192.6000 120.4500 197.4000 ;
	    RECT 119.4000 191.4000 120.6000 192.6000 ;
	    RECT 117.0000 161.4000 118.2000 162.6000 ;
	    RECT 126.6000 161.4000 127.8000 162.6000 ;
	    RECT 93.0000 143.4000 94.2000 144.6000 ;
	    RECT 126.7500 42.6000 127.6500 161.4000 ;
	    RECT 133.9500 138.4500 134.8500 245.4000 ;
	    RECT 165.1500 240.6000 166.0500 323.4000 ;
	    RECT 167.4000 317.4000 168.6000 318.6000 ;
	    RECT 167.5500 294.6000 168.4500 317.4000 ;
	    RECT 167.4000 293.4000 168.6000 294.6000 ;
	    RECT 167.4000 287.4000 168.6000 288.6000 ;
	    RECT 167.5500 285.6000 168.4500 287.4000 ;
	    RECT 167.4000 284.4000 168.6000 285.6000 ;
	    RECT 169.8000 276.3000 171.0000 296.7000 ;
	    RECT 172.2000 276.3000 173.4000 296.7000 ;
	    RECT 174.6000 276.3000 175.8000 293.7000 ;
	    RECT 177.1500 288.6000 178.0500 497.4000 ;
	    RECT 184.3500 492.6000 185.2500 503.4000 ;
	    RECT 186.7500 498.6000 187.6500 707.5500 ;
	    RECT 189.0000 707.4000 190.2000 707.5500 ;
	    RECT 193.8000 707.4000 195.0000 708.6000 ;
	    RECT 205.8000 707.4000 207.0000 708.6000 ;
	    RECT 189.0000 701.4000 190.2000 702.6000 ;
	    RECT 196.2000 702.4500 197.4000 702.6000 ;
	    RECT 191.5500 701.5500 197.4000 702.4500 ;
	    RECT 189.1500 687.6000 190.0500 701.4000 ;
	    RECT 191.5500 696.6000 192.4500 701.5500 ;
	    RECT 196.2000 701.4000 197.4000 701.5500 ;
	    RECT 196.2000 698.4000 197.4000 699.6000 ;
	    RECT 191.4000 695.4000 192.6000 696.6000 ;
	    RECT 196.3500 690.6000 197.2500 698.4000 ;
	    RECT 198.6000 695.4000 199.8000 696.6000 ;
	    RECT 213.0000 695.4000 214.2000 696.6000 ;
	    RECT 196.2000 689.4000 197.4000 690.6000 ;
	    RECT 189.0000 686.4000 190.2000 687.6000 ;
	    RECT 198.7500 654.6000 199.6500 695.4000 ;
	    RECT 213.1500 687.6000 214.0500 695.4000 ;
	    RECT 213.0000 686.4000 214.2000 687.6000 ;
	    RECT 213.0000 683.4000 214.2000 684.6000 ;
	    RECT 215.5500 681.4500 216.4500 737.4000 ;
	    RECT 217.9500 702.6000 218.8500 740.5500 ;
	    RECT 217.8000 701.4000 219.0000 702.6000 ;
	    RECT 213.1500 680.5500 216.4500 681.4500 ;
	    RECT 213.1500 660.6000 214.0500 680.5500 ;
	    RECT 217.9500 678.6000 218.8500 701.4000 ;
	    RECT 220.3500 696.6000 221.2500 824.4000 ;
	    RECT 222.7500 801.6000 223.6500 827.4000 ;
	    RECT 225.0000 803.4000 226.2000 804.6000 ;
	    RECT 225.1500 801.6000 226.0500 803.4000 ;
	    RECT 222.6000 800.4000 223.8000 801.6000 ;
	    RECT 225.0000 800.4000 226.2000 801.6000 ;
	    RECT 232.2000 797.4000 233.4000 798.6000 ;
	    RECT 232.3500 765.6000 233.2500 797.4000 ;
	    RECT 237.1500 780.6000 238.0500 896.4000 ;
	    RECT 239.4000 890.4000 240.6000 891.6000 ;
	    RECT 239.5500 855.6000 240.4500 890.4000 ;
	    RECT 239.4000 854.4000 240.6000 855.6000 ;
	    RECT 239.5500 819.6000 240.4500 854.4000 ;
	    RECT 239.4000 818.4000 240.6000 819.6000 ;
	    RECT 237.0000 779.4000 238.2000 780.6000 ;
	    RECT 237.1500 765.6000 238.0500 779.4000 ;
	    RECT 232.2000 764.4000 233.4000 765.6000 ;
	    RECT 237.0000 764.4000 238.2000 765.6000 ;
	    RECT 232.3500 756.6000 233.2500 764.4000 ;
	    RECT 234.6000 761.4000 235.8000 762.6000 ;
	    RECT 232.2000 755.4000 233.4000 756.6000 ;
	    RECT 232.2000 749.4000 233.4000 750.6000 ;
	    RECT 227.4000 737.4000 228.6000 738.6000 ;
	    RECT 227.5500 732.6000 228.4500 737.4000 ;
	    RECT 229.8000 734.4000 231.0000 735.6000 ;
	    RECT 227.4000 731.4000 228.6000 732.6000 ;
	    RECT 220.2000 695.4000 221.4000 696.6000 ;
	    RECT 225.0000 689.4000 226.2000 690.6000 ;
	    RECT 222.6000 683.4000 223.8000 684.6000 ;
	    RECT 220.2000 680.4000 221.4000 681.6000 ;
	    RECT 220.3500 678.6000 221.2500 680.4000 ;
	    RECT 222.7500 678.6000 223.6500 683.4000 ;
	    RECT 225.1500 678.6000 226.0500 689.4000 ;
	    RECT 229.9500 684.6000 230.8500 734.4000 ;
	    RECT 232.3500 705.6000 233.2500 749.4000 ;
	    RECT 232.2000 704.4000 233.4000 705.6000 ;
	    RECT 232.2000 701.4000 233.4000 702.6000 ;
	    RECT 229.8000 683.4000 231.0000 684.6000 ;
	    RECT 227.4000 680.4000 228.6000 681.6000 ;
	    RECT 215.4000 677.4000 216.6000 678.6000 ;
	    RECT 217.8000 677.4000 219.0000 678.6000 ;
	    RECT 220.2000 677.4000 221.4000 678.6000 ;
	    RECT 222.6000 677.4000 223.8000 678.6000 ;
	    RECT 225.0000 677.4000 226.2000 678.6000 ;
	    RECT 215.5500 672.6000 216.4500 677.4000 ;
	    RECT 215.4000 671.4000 216.6000 672.6000 ;
	    RECT 213.0000 659.4000 214.2000 660.6000 ;
	    RECT 198.6000 653.4000 199.8000 654.6000 ;
	    RECT 189.0000 641.4000 190.2000 642.6000 ;
	    RECT 186.6000 497.4000 187.8000 498.6000 ;
	    RECT 184.2000 491.4000 185.4000 492.6000 ;
	    RECT 186.7500 438.6000 187.6500 497.4000 ;
	    RECT 186.6000 437.4000 187.8000 438.6000 ;
	    RECT 184.2000 431.4000 185.4000 432.6000 ;
	    RECT 184.3500 321.6000 185.2500 431.4000 ;
	    RECT 186.6000 380.4000 187.8000 381.6000 ;
	    RECT 186.7500 342.6000 187.6500 380.4000 ;
	    RECT 189.1500 342.6000 190.0500 641.4000 ;
	    RECT 196.2000 623.4000 197.4000 624.6000 ;
	    RECT 193.8000 578.4000 195.0000 579.6000 ;
	    RECT 191.4000 531.4500 192.6000 531.6000 ;
	    RECT 193.9500 531.4500 194.8500 578.4000 ;
	    RECT 191.4000 530.5500 194.8500 531.4500 ;
	    RECT 191.4000 530.4000 192.6000 530.5500 ;
	    RECT 191.5500 378.6000 192.4500 530.4000 ;
	    RECT 193.8000 527.4000 195.0000 528.6000 ;
	    RECT 193.9500 504.6000 194.8500 527.4000 ;
	    RECT 193.8000 503.4000 195.0000 504.6000 ;
	    RECT 193.8000 464.4000 195.0000 465.6000 ;
	    RECT 193.9500 444.6000 194.8500 464.4000 ;
	    RECT 193.8000 443.4000 195.0000 444.6000 ;
	    RECT 193.8000 437.4000 195.0000 438.6000 ;
	    RECT 193.9500 426.6000 194.8500 437.4000 ;
	    RECT 193.8000 425.4000 195.0000 426.6000 ;
	    RECT 191.4000 377.4000 192.6000 378.6000 ;
	    RECT 186.6000 341.4000 187.8000 342.6000 ;
	    RECT 189.0000 341.4000 190.2000 342.6000 ;
	    RECT 186.7500 321.6000 187.6500 341.4000 ;
	    RECT 193.8000 338.4000 195.0000 339.6000 ;
	    RECT 193.9500 336.6000 194.8500 338.4000 ;
	    RECT 193.8000 335.4000 195.0000 336.6000 ;
	    RECT 184.2000 320.4000 185.4000 321.6000 ;
	    RECT 186.6000 320.4000 187.8000 321.6000 ;
	    RECT 177.0000 287.4000 178.2000 288.6000 ;
	    RECT 177.0000 281.4000 178.2000 282.6000 ;
	    RECT 177.0000 275.4000 178.2000 276.6000 ;
	    RECT 179.4000 276.3000 180.6000 293.7000 ;
	    RECT 181.8000 293.4000 183.0000 294.6000 ;
	    RECT 181.9500 279.6000 182.8500 293.4000 ;
	    RECT 181.8000 278.4000 183.0000 279.6000 ;
	    RECT 184.2000 276.3000 185.4000 293.7000 ;
	    RECT 186.6000 276.3000 187.8000 296.7000 ;
	    RECT 189.0000 276.3000 190.2000 296.7000 ;
	    RECT 191.4000 276.3000 192.6000 296.7000 ;
	    RECT 177.1500 270.6000 178.0500 275.4000 ;
	    RECT 196.3500 270.6000 197.2500 623.4000 ;
	    RECT 198.7500 606.6000 199.6500 653.4000 ;
	    RECT 215.5500 645.6000 216.4500 671.4000 ;
	    RECT 217.8000 659.4000 219.0000 660.6000 ;
	    RECT 222.6000 659.4000 223.8000 660.6000 ;
	    RECT 215.4000 644.4000 216.6000 645.6000 ;
	    RECT 217.9500 642.6000 218.8500 659.4000 ;
	    RECT 220.2000 645.4500 221.4000 645.6000 ;
	    RECT 222.7500 645.4500 223.6500 659.4000 ;
	    RECT 220.2000 644.5500 223.6500 645.4500 ;
	    RECT 220.2000 644.4000 221.4000 644.5500 ;
	    RECT 217.8000 641.4000 219.0000 642.6000 ;
	    RECT 222.6000 641.4000 223.8000 642.6000 ;
	    RECT 217.8000 635.4000 219.0000 636.6000 ;
	    RECT 215.4000 623.4000 216.6000 624.6000 ;
	    RECT 215.5500 612.6000 216.4500 623.4000 ;
	    RECT 215.4000 611.4000 216.6000 612.6000 ;
	    RECT 198.6000 605.4000 199.8000 606.6000 ;
	    RECT 210.6000 581.4000 211.8000 582.6000 ;
	    RECT 215.4000 581.4000 216.6000 582.6000 ;
	    RECT 210.7500 579.6000 211.6500 581.4000 ;
	    RECT 215.5500 579.6000 216.4500 581.4000 ;
	    RECT 210.6000 578.4000 211.8000 579.6000 ;
	    RECT 215.4000 578.4000 216.6000 579.6000 ;
	    RECT 213.0000 569.4000 214.2000 570.6000 ;
	    RECT 198.6000 563.4000 199.8000 564.6000 ;
	    RECT 198.7500 462.6000 199.6500 563.4000 ;
	    RECT 213.1500 501.6000 214.0500 569.4000 ;
	    RECT 215.4000 503.4000 216.6000 504.6000 ;
	    RECT 213.0000 500.4000 214.2000 501.6000 ;
	    RECT 198.6000 461.4000 199.8000 462.6000 ;
	    RECT 198.6000 458.4000 199.8000 459.6000 ;
	    RECT 213.0000 458.4000 214.2000 459.6000 ;
	    RECT 198.7500 450.6000 199.6500 458.4000 ;
	    RECT 198.6000 449.4000 199.8000 450.6000 ;
	    RECT 198.6000 440.4000 199.8000 441.6000 ;
	    RECT 198.7500 402.6000 199.6500 440.4000 ;
	    RECT 198.6000 401.4000 199.8000 402.6000 ;
	    RECT 198.6000 377.4000 199.8000 378.6000 ;
	    RECT 198.7500 375.6000 199.6500 377.4000 ;
	    RECT 198.6000 374.4000 199.8000 375.6000 ;
	    RECT 198.6000 339.4500 199.8000 339.6000 ;
	    RECT 198.6000 338.5500 202.0500 339.4500 ;
	    RECT 198.6000 338.4000 199.8000 338.5500 ;
	    RECT 198.7500 336.6000 199.6500 338.4000 ;
	    RECT 198.6000 335.4000 199.8000 336.6000 ;
	    RECT 198.7500 294.6000 199.6500 335.4000 ;
	    RECT 201.1500 315.6000 202.0500 338.5500 ;
	    RECT 201.0000 314.4000 202.2000 315.6000 ;
	    RECT 198.6000 293.4000 199.8000 294.6000 ;
	    RECT 205.8000 293.4000 207.0000 294.6000 ;
	    RECT 205.9500 291.6000 206.8500 293.4000 ;
	    RECT 205.8000 290.4000 207.0000 291.6000 ;
	    RECT 177.0000 269.4000 178.2000 270.6000 ;
	    RECT 196.2000 269.4000 197.4000 270.6000 ;
	    RECT 177.1500 252.6000 178.0500 269.4000 ;
	    RECT 172.2000 251.4000 173.4000 252.6000 ;
	    RECT 177.0000 251.4000 178.2000 252.6000 ;
	    RECT 181.8000 251.4000 183.0000 252.6000 ;
	    RECT 172.3500 240.6000 173.2500 251.4000 ;
	    RECT 165.0000 239.4000 166.2000 240.6000 ;
	    RECT 169.8000 239.4000 171.0000 240.6000 ;
	    RECT 172.2000 239.4000 173.4000 240.6000 ;
	    RECT 143.4000 216.3000 144.6000 236.7000 ;
	    RECT 145.8000 216.3000 147.0000 236.7000 ;
	    RECT 148.2000 216.3000 149.4000 236.7000 ;
	    RECT 150.6000 216.3000 151.8000 233.7000 ;
	    RECT 153.0000 218.4000 154.2000 219.6000 ;
	    RECT 153.1500 213.4500 154.0500 218.4000 ;
	    RECT 155.4000 216.3000 156.6000 233.7000 ;
	    RECT 157.8000 227.4000 159.0000 228.6000 ;
	    RECT 157.9500 222.6000 158.8500 227.4000 ;
	    RECT 157.8000 221.4000 159.0000 222.6000 ;
	    RECT 160.2000 216.3000 161.4000 233.7000 ;
	    RECT 162.6000 216.3000 163.8000 236.7000 ;
	    RECT 165.0000 216.3000 166.2000 236.7000 ;
	    RECT 167.4000 224.4000 168.6000 225.6000 ;
	    RECT 150.7500 212.5500 154.0500 213.4500 ;
	    RECT 136.2000 203.4000 137.4000 204.6000 ;
	    RECT 136.3500 150.6000 137.2500 203.4000 ;
	    RECT 136.2000 149.4000 137.4000 150.6000 ;
	    RECT 136.2000 138.4500 137.4000 138.6000 ;
	    RECT 133.9500 137.5500 137.4000 138.4500 ;
	    RECT 136.2000 137.4000 137.4000 137.5500 ;
	    RECT 131.4000 134.4000 132.6000 135.6000 ;
	    RECT 131.5500 126.6000 132.4500 134.4000 ;
	    RECT 131.4000 125.4000 132.6000 126.6000 ;
	    RECT 138.6000 126.3000 139.8000 146.7000 ;
	    RECT 141.0000 126.3000 142.2000 146.7000 ;
	    RECT 143.4000 129.3000 144.6000 146.7000 ;
	    RECT 145.8000 143.4000 147.0000 144.6000 ;
	    RECT 145.9500 141.6000 146.8500 143.4000 ;
	    RECT 145.8000 140.4000 147.0000 141.6000 ;
	    RECT 148.2000 129.3000 149.4000 146.7000 ;
	    RECT 150.7500 144.6000 151.6500 212.5500 ;
	    RECT 167.5500 210.6000 168.4500 224.4000 ;
	    RECT 167.4000 209.4000 168.6000 210.6000 ;
	    RECT 153.0000 203.4000 154.2000 204.6000 ;
	    RECT 153.1500 195.6000 154.0500 203.4000 ;
	    RECT 162.6000 200.4000 163.8000 201.6000 ;
	    RECT 162.7500 198.6000 163.6500 200.4000 ;
	    RECT 162.6000 197.4000 163.8000 198.6000 ;
	    RECT 169.9500 195.6000 170.8500 239.4000 ;
	    RECT 172.2000 236.4000 173.4000 237.6000 ;
	    RECT 172.3500 228.6000 173.2500 236.4000 ;
	    RECT 172.2000 227.4000 173.4000 228.6000 ;
	    RECT 179.4000 203.4000 180.6000 204.6000 ;
	    RECT 153.0000 194.4000 154.2000 195.6000 ;
	    RECT 169.8000 194.4000 171.0000 195.6000 ;
	    RECT 177.0000 176.4000 178.2000 177.6000 ;
	    RECT 177.1500 168.6000 178.0500 176.4000 ;
	    RECT 177.0000 167.4000 178.2000 168.6000 ;
	    RECT 174.6000 149.4000 175.8000 150.6000 ;
	    RECT 150.6000 143.4000 151.8000 144.6000 ;
	    RECT 150.7500 90.4500 151.6500 143.4000 ;
	    RECT 153.0000 129.3000 154.2000 146.7000 ;
	    RECT 155.4000 126.3000 156.6000 146.7000 ;
	    RECT 157.8000 126.3000 159.0000 146.7000 ;
	    RECT 160.2000 126.3000 161.4000 146.7000 ;
	    RECT 174.7500 132.6000 175.6500 149.4000 ;
	    RECT 174.6000 131.4000 175.8000 132.6000 ;
	    RECT 179.5500 111.6000 180.4500 203.4000 ;
	    RECT 181.9500 165.6000 182.8500 251.4000 ;
	    RECT 205.8000 227.4000 207.0000 228.6000 ;
	    RECT 193.8000 215.4000 195.0000 216.6000 ;
	    RECT 193.9500 204.6000 194.8500 215.4000 ;
	    RECT 193.8000 203.4000 195.0000 204.6000 ;
	    RECT 205.9500 198.6000 206.8500 227.4000 ;
	    RECT 208.2000 221.4000 209.4000 222.6000 ;
	    RECT 205.8000 197.4000 207.0000 198.6000 ;
	    RECT 208.3500 186.6000 209.2500 221.4000 ;
	    RECT 213.1500 216.6000 214.0500 458.4000 ;
	    RECT 217.9500 441.6000 218.8500 635.4000 ;
	    RECT 220.2000 605.4000 221.4000 606.6000 ;
	    RECT 220.3500 486.6000 221.2500 605.4000 ;
	    RECT 222.7500 582.6000 223.6500 641.4000 ;
	    RECT 227.5500 621.6000 228.4500 680.4000 ;
	    RECT 232.3500 666.6000 233.2500 701.4000 ;
	    RECT 232.2000 665.4000 233.4000 666.6000 ;
	    RECT 227.4000 620.4000 228.6000 621.6000 ;
	    RECT 232.3500 585.6000 233.2500 665.4000 ;
	    RECT 234.7500 630.6000 235.6500 761.4000 ;
	    RECT 237.0000 755.4000 238.2000 756.6000 ;
	    RECT 237.1500 660.6000 238.0500 755.4000 ;
	    RECT 239.5500 744.6000 240.4500 818.4000 ;
	    RECT 241.9500 798.6000 242.8500 1181.4000 ;
	    RECT 246.7500 1161.6000 247.6500 1193.4000 ;
	    RECT 246.6000 1160.4000 247.8000 1161.6000 ;
	    RECT 249.1500 1116.6000 250.0500 1220.4000 ;
	    RECT 251.4000 1217.4000 252.6000 1218.6000 ;
	    RECT 251.5500 1206.6000 252.4500 1217.4000 ;
	    RECT 251.4000 1205.4000 252.6000 1206.6000 ;
	    RECT 256.3500 1191.4501 257.2500 1220.4000 ;
	    RECT 253.9500 1190.5500 257.2500 1191.4501 ;
	    RECT 253.9500 1167.4501 254.8500 1190.5500 ;
	    RECT 256.2000 1187.4000 257.4000 1188.6000 ;
	    RECT 253.9500 1166.5500 257.2500 1167.4501 ;
	    RECT 253.8000 1163.4000 255.0000 1164.6000 ;
	    RECT 253.9500 1161.6000 254.8500 1163.4000 ;
	    RECT 253.8000 1160.4000 255.0000 1161.6000 ;
	    RECT 253.9500 1158.6000 254.8500 1160.4000 ;
	    RECT 253.8000 1157.4000 255.0000 1158.6000 ;
	    RECT 256.3500 1146.6000 257.2500 1166.5500 ;
	    RECT 258.7500 1146.6000 259.6500 1235.4000 ;
	    RECT 261.1500 1188.6000 262.0500 1259.4000 ;
	    RECT 263.5500 1224.6000 264.4500 1331.4000 ;
	    RECT 275.4000 1319.4000 276.6000 1320.6000 ;
	    RECT 275.5500 1314.6000 276.4500 1319.4000 ;
	    RECT 275.4000 1313.4000 276.6000 1314.6000 ;
	    RECT 273.0000 1301.4000 274.2000 1302.6000 ;
	    RECT 273.1500 1290.6000 274.0500 1301.4000 ;
	    RECT 273.0000 1289.4000 274.2000 1290.6000 ;
	    RECT 265.8000 1266.3000 267.0000 1286.7001 ;
	    RECT 268.2000 1266.3000 269.4000 1286.7001 ;
	    RECT 270.6000 1266.3000 271.8000 1286.7001 ;
	    RECT 273.0000 1269.3000 274.2000 1286.7001 ;
	    RECT 275.5500 1284.6000 276.4500 1313.4000 ;
	    RECT 280.2000 1301.4000 281.4000 1302.6000 ;
	    RECT 282.7500 1290.6000 283.6500 1400.4000 ;
	    RECT 285.1500 1398.6000 286.0500 1400.4000 ;
	    RECT 285.0000 1397.4000 286.2000 1398.6000 ;
	    RECT 287.4000 1307.4000 288.6000 1308.6000 ;
	    RECT 311.5500 1290.6000 312.4500 1403.4000 ;
	    RECT 313.8000 1400.4000 315.0000 1401.6000 ;
	    RECT 282.6000 1289.4000 283.8000 1290.6000 ;
	    RECT 292.2000 1289.4000 293.4000 1290.6000 ;
	    RECT 311.4000 1289.4000 312.6000 1290.6000 ;
	    RECT 275.4000 1283.4000 276.6000 1284.6000 ;
	    RECT 263.4000 1223.4000 264.6000 1224.6000 ;
	    RECT 273.0000 1220.4000 274.2000 1221.6000 ;
	    RECT 273.1500 1200.6000 274.0500 1220.4000 ;
	    RECT 273.0000 1199.4000 274.2000 1200.6000 ;
	    RECT 261.0000 1187.4000 262.2000 1188.6000 ;
	    RECT 261.0000 1184.4000 262.2000 1185.6000 ;
	    RECT 261.1500 1182.6000 262.0500 1184.4000 ;
	    RECT 261.0000 1181.4000 262.2000 1182.6000 ;
	    RECT 263.4000 1176.3000 264.6000 1196.7001 ;
	    RECT 265.8000 1176.3000 267.0000 1196.7001 ;
	    RECT 268.2000 1176.3000 269.4000 1193.7001 ;
	    RECT 270.6000 1193.4000 271.8000 1194.6000 ;
	    RECT 270.7500 1182.6000 271.6500 1193.4000 ;
	    RECT 270.6000 1181.4000 271.8000 1182.6000 ;
	    RECT 273.0000 1176.3000 274.2000 1193.7001 ;
	    RECT 275.5500 1179.6000 276.4500 1283.4000 ;
	    RECT 277.8000 1269.3000 279.0000 1286.7001 ;
	    RECT 280.2000 1280.4000 281.4000 1281.6000 ;
	    RECT 280.3500 1272.6000 281.2500 1280.4000 ;
	    RECT 280.2000 1271.4000 281.4000 1272.6000 ;
	    RECT 282.6000 1269.3000 283.8000 1286.7001 ;
	    RECT 285.0000 1266.3000 286.2000 1286.7001 ;
	    RECT 287.4000 1266.3000 288.6000 1286.7001 ;
	    RECT 289.8000 1277.4000 291.0000 1278.6000 ;
	    RECT 287.4000 1247.4000 288.6000 1248.6000 ;
	    RECT 285.0000 1223.4000 286.2000 1224.6000 ;
	    RECT 287.5500 1218.6000 288.4500 1247.4000 ;
	    RECT 287.4000 1217.4000 288.6000 1218.6000 ;
	    RECT 277.8000 1211.4000 279.0000 1212.6000 ;
	    RECT 277.9500 1200.6000 278.8500 1211.4000 ;
	    RECT 287.4000 1205.4000 288.6000 1206.6000 ;
	    RECT 277.8000 1199.4000 279.0000 1200.6000 ;
	    RECT 275.4000 1178.4000 276.6000 1179.6000 ;
	    RECT 275.4000 1175.4000 276.6000 1176.6000 ;
	    RECT 277.8000 1176.3000 279.0000 1193.7001 ;
	    RECT 280.2000 1176.3000 281.4000 1196.7001 ;
	    RECT 282.6000 1176.3000 283.8000 1196.7001 ;
	    RECT 285.0000 1176.3000 286.2000 1196.7001 ;
	    RECT 275.5500 1167.6000 276.4500 1175.4000 ;
	    RECT 275.4000 1166.4000 276.6000 1167.6000 ;
	    RECT 277.8000 1163.4000 279.0000 1164.6000 ;
	    RECT 265.8000 1157.4000 267.0000 1158.6000 ;
	    RECT 275.4000 1157.4000 276.6000 1158.6000 ;
	    RECT 265.9500 1152.6000 266.8500 1157.4000 ;
	    RECT 265.8000 1151.4000 267.0000 1152.6000 ;
	    RECT 273.0000 1151.4000 274.2000 1152.6000 ;
	    RECT 256.2000 1145.4000 257.4000 1146.6000 ;
	    RECT 258.6000 1145.4000 259.8000 1146.6000 ;
	    RECT 263.4000 1145.4000 264.6000 1146.6000 ;
	    RECT 256.2000 1139.4000 257.4000 1140.6000 ;
	    RECT 253.8000 1127.4000 255.0000 1128.6000 ;
	    RECT 244.2000 1115.4000 245.4000 1116.6000 ;
	    RECT 249.0000 1115.4000 250.2000 1116.6000 ;
	    RECT 244.3500 1044.4501 245.2500 1115.4000 ;
	    RECT 246.6000 1109.4000 247.8000 1110.6000 ;
	    RECT 246.7500 1098.6000 247.6500 1109.4000 ;
	    RECT 249.0000 1100.4000 250.2000 1101.6000 ;
	    RECT 246.6000 1097.4000 247.8000 1098.6000 ;
	    RECT 249.1500 1092.6000 250.0500 1100.4000 ;
	    RECT 251.4000 1097.4000 252.6000 1098.6000 ;
	    RECT 249.0000 1091.4000 250.2000 1092.6000 ;
	    RECT 246.6000 1044.4501 247.8000 1044.6000 ;
	    RECT 244.3500 1043.5500 247.8000 1044.4501 ;
	    RECT 246.6000 1043.4000 247.8000 1043.5500 ;
	    RECT 244.2000 1025.4000 245.4000 1026.6000 ;
	    RECT 244.3500 939.6000 245.2500 1025.4000 ;
	    RECT 251.5500 1020.6000 252.4500 1097.4000 ;
	    RECT 253.9500 1074.6000 254.8500 1127.4000 ;
	    RECT 256.3500 1125.6000 257.2500 1139.4000 ;
	    RECT 256.2000 1124.4000 257.4000 1125.6000 ;
	    RECT 256.2000 1091.4000 257.4000 1092.6000 ;
	    RECT 258.7500 1092.4501 259.6500 1145.4000 ;
	    RECT 261.0000 1109.4000 262.2000 1110.6000 ;
	    RECT 261.1500 1098.6000 262.0500 1109.4000 ;
	    RECT 263.5500 1101.6000 264.4500 1145.4000 ;
	    RECT 273.1500 1122.6000 274.0500 1151.4000 ;
	    RECT 270.6000 1121.4000 271.8000 1122.6000 ;
	    RECT 273.0000 1121.4000 274.2000 1122.6000 ;
	    RECT 263.4000 1100.4000 264.6000 1101.6000 ;
	    RECT 261.0000 1097.4000 262.2000 1098.6000 ;
	    RECT 270.7500 1092.6000 271.6500 1121.4000 ;
	    RECT 273.0000 1097.4000 274.2000 1098.6000 ;
	    RECT 273.1500 1092.6000 274.0500 1097.4000 ;
	    RECT 258.7500 1091.5500 262.0500 1092.4501 ;
	    RECT 253.8000 1073.4000 255.0000 1074.6000 ;
	    RECT 256.3500 1062.6000 257.2500 1091.4000 ;
	    RECT 258.6000 1085.4000 259.8000 1086.6000 ;
	    RECT 258.7500 1068.6000 259.6500 1085.4000 ;
	    RECT 258.6000 1067.4000 259.8000 1068.6000 ;
	    RECT 261.1500 1065.6000 262.0500 1091.5500 ;
	    RECT 270.6000 1091.4000 271.8000 1092.6000 ;
	    RECT 273.0000 1091.4000 274.2000 1092.6000 ;
	    RECT 261.0000 1064.4000 262.2000 1065.6000 ;
	    RECT 275.5500 1062.6000 276.4500 1157.4000 ;
	    RECT 277.9500 1140.6000 278.8500 1163.4000 ;
	    RECT 287.5500 1158.6000 288.4500 1205.4000 ;
	    RECT 289.9500 1167.6000 290.8500 1277.4000 ;
	    RECT 289.8000 1166.4000 291.0000 1167.6000 ;
	    RECT 287.4000 1157.4000 288.6000 1158.6000 ;
	    RECT 287.4000 1151.4000 288.6000 1152.6000 ;
	    RECT 277.8000 1139.4000 279.0000 1140.6000 ;
	    RECT 277.9500 1128.6000 278.8500 1139.4000 ;
	    RECT 277.8000 1127.4000 279.0000 1128.6000 ;
	    RECT 280.2000 1118.4000 281.4000 1119.6000 ;
	    RECT 277.8000 1103.4000 279.0000 1104.6000 ;
	    RECT 256.2000 1062.4501 257.4000 1062.6000 ;
	    RECT 253.9500 1061.5500 257.4000 1062.4501 ;
	    RECT 251.4000 1019.4000 252.6000 1020.6000 ;
	    RECT 253.9500 978.6000 254.8500 1061.5500 ;
	    RECT 256.2000 1061.4000 257.4000 1061.5500 ;
	    RECT 275.4000 1061.4000 276.6000 1062.6000 ;
	    RECT 268.2000 1058.4000 269.4000 1059.6000 ;
	    RECT 268.3500 1050.6000 269.2500 1058.4000 ;
	    RECT 268.2000 1049.4000 269.4000 1050.6000 ;
	    RECT 270.6000 1043.4000 271.8000 1044.6000 ;
	    RECT 273.0000 1043.4000 274.2000 1044.6000 ;
	    RECT 263.4000 1040.4000 264.6000 1041.6000 ;
	    RECT 268.2000 1040.4000 269.4000 1041.6000 ;
	    RECT 263.5500 1020.6000 264.4500 1040.4000 ;
	    RECT 265.8000 1037.4000 267.0000 1038.6000 ;
	    RECT 265.9500 1032.6000 266.8500 1037.4000 ;
	    RECT 265.8000 1031.4000 267.0000 1032.6000 ;
	    RECT 263.4000 1019.4000 264.6000 1020.6000 ;
	    RECT 265.8000 983.4000 267.0000 984.6000 ;
	    RECT 265.9500 981.6000 266.8500 983.4000 ;
	    RECT 268.3500 981.6000 269.2500 1040.4000 ;
	    RECT 270.7500 999.6000 271.6500 1043.4000 ;
	    RECT 273.1500 1038.6000 274.0500 1043.4000 ;
	    RECT 273.0000 1037.4000 274.2000 1038.6000 ;
	    RECT 273.0000 1034.4000 274.2000 1035.6000 ;
	    RECT 273.1500 1020.6000 274.0500 1034.4000 ;
	    RECT 277.9500 1032.6000 278.8500 1103.4000 ;
	    RECT 277.8000 1031.4000 279.0000 1032.6000 ;
	    RECT 280.3500 1029.4501 281.2500 1118.4000 ;
	    RECT 285.0000 1049.4000 286.2000 1050.6000 ;
	    RECT 277.9500 1028.5500 281.2500 1029.4501 ;
	    RECT 273.0000 1019.4000 274.2000 1020.6000 ;
	    RECT 270.6000 998.4000 271.8000 999.6000 ;
	    RECT 275.4000 989.4000 276.6000 990.6000 ;
	    RECT 273.0000 983.4000 274.2000 984.6000 ;
	    RECT 265.8000 980.4000 267.0000 981.6000 ;
	    RECT 268.2000 980.4000 269.4000 981.6000 ;
	    RECT 249.0000 977.4000 250.2000 978.6000 ;
	    RECT 253.8000 977.4000 255.0000 978.6000 ;
	    RECT 258.6000 977.4000 259.8000 978.6000 ;
	    RECT 270.6000 977.4000 271.8000 978.6000 ;
	    RECT 249.1500 972.6000 250.0500 977.4000 ;
	    RECT 249.0000 971.4000 250.2000 972.6000 ;
	    RECT 258.7500 966.6000 259.6500 977.4000 ;
	    RECT 258.6000 965.4000 259.8000 966.6000 ;
	    RECT 256.2000 953.4000 257.4000 954.6000 ;
	    RECT 249.0000 947.4000 250.2000 948.6000 ;
	    RECT 249.1500 942.6000 250.0500 947.4000 ;
	    RECT 253.8000 945.4500 255.0000 945.6000 ;
	    RECT 256.3500 945.4500 257.2500 953.4000 ;
	    RECT 270.7500 948.4500 271.6500 977.4000 ;
	    RECT 273.1500 975.6000 274.0500 983.4000 ;
	    RECT 275.5500 975.6000 276.4500 989.4000 ;
	    RECT 273.0000 974.4000 274.2000 975.6000 ;
	    RECT 275.4000 974.4000 276.6000 975.6000 ;
	    RECT 275.4000 950.4000 276.6000 951.6000 ;
	    RECT 270.7500 947.5500 274.0500 948.4500 ;
	    RECT 253.8000 944.5500 257.2500 945.4500 ;
	    RECT 253.8000 944.4000 255.0000 944.5500 ;
	    RECT 249.0000 941.4000 250.2000 942.6000 ;
	    RECT 244.2000 938.4000 245.4000 939.6000 ;
	    RECT 253.8000 935.4000 255.0000 936.6000 ;
	    RECT 244.2000 929.4000 245.4000 930.6000 ;
	    RECT 244.3500 924.6000 245.2500 929.4000 ;
	    RECT 253.9500 924.6000 254.8500 935.4000 ;
	    RECT 265.8000 929.4000 267.0000 930.6000 ;
	    RECT 265.9500 924.6000 266.8500 929.4000 ;
	    RECT 244.2000 923.4000 245.4000 924.6000 ;
	    RECT 253.8000 923.4000 255.0000 924.6000 ;
	    RECT 265.8000 923.4000 267.0000 924.6000 ;
	    RECT 251.4000 911.4000 252.6000 912.6000 ;
	    RECT 251.5500 864.6000 252.4500 911.4000 ;
	    RECT 261.0000 866.4000 262.2000 867.6000 ;
	    RECT 251.4000 863.4000 252.6000 864.6000 ;
	    RECT 246.6000 839.4000 247.8000 840.6000 ;
	    RECT 244.2000 833.4000 245.4000 834.6000 ;
	    RECT 244.3500 819.6000 245.2500 833.4000 ;
	    RECT 244.2000 818.4000 245.4000 819.6000 ;
	    RECT 246.7500 798.6000 247.6500 839.4000 ;
	    RECT 253.8000 827.4000 255.0000 828.6000 ;
	    RECT 253.9500 801.6000 254.8500 827.4000 ;
	    RECT 249.0000 800.4000 250.2000 801.6000 ;
	    RECT 253.8000 800.4000 255.0000 801.6000 ;
	    RECT 256.2000 800.4000 257.4000 801.6000 ;
	    RECT 241.8000 797.4000 243.0000 798.6000 ;
	    RECT 246.6000 797.4000 247.8000 798.6000 ;
	    RECT 239.4000 743.4000 240.6000 744.6000 ;
	    RECT 239.4000 701.4000 240.6000 702.6000 ;
	    RECT 239.4000 677.4000 240.6000 678.6000 ;
	    RECT 237.0000 659.4000 238.2000 660.6000 ;
	    RECT 239.5500 654.6000 240.4500 677.4000 ;
	    RECT 239.4000 653.4000 240.6000 654.6000 ;
	    RECT 239.4000 638.4000 240.6000 639.6000 ;
	    RECT 239.5500 636.6000 240.4500 638.4000 ;
	    RECT 239.4000 635.4000 240.6000 636.6000 ;
	    RECT 234.6000 629.4000 235.8000 630.6000 ;
	    RECT 239.4000 629.4000 240.6000 630.6000 ;
	    RECT 234.6000 623.4000 235.8000 624.6000 ;
	    RECT 234.7500 606.6000 235.6500 623.4000 ;
	    RECT 237.0000 620.4000 238.2000 621.6000 ;
	    RECT 234.6000 605.4000 235.8000 606.6000 ;
	    RECT 237.1500 600.6000 238.0500 620.4000 ;
	    RECT 239.5500 618.6000 240.4500 629.4000 ;
	    RECT 241.9500 618.6000 242.8500 797.4000 ;
	    RECT 249.1500 750.6000 250.0500 800.4000 ;
	    RECT 251.4000 797.4000 252.6000 798.6000 ;
	    RECT 251.5500 780.6000 252.4500 797.4000 ;
	    RECT 251.4000 779.4000 252.6000 780.6000 ;
	    RECT 251.5500 777.6000 252.4500 779.4000 ;
	    RECT 251.4000 776.4000 252.6000 777.6000 ;
	    RECT 251.4000 764.4000 252.6000 765.6000 ;
	    RECT 249.0000 749.4000 250.2000 750.6000 ;
	    RECT 251.5500 744.6000 252.4500 764.4000 ;
	    RECT 256.3500 762.6000 257.2500 800.4000 ;
	    RECT 256.2000 761.4000 257.4000 762.6000 ;
	    RECT 251.4000 743.4000 252.6000 744.6000 ;
	    RECT 244.2000 740.4000 245.4000 741.6000 ;
	    RECT 244.3500 678.6000 245.2500 740.4000 ;
	    RECT 249.0000 734.4000 250.2000 735.6000 ;
	    RECT 249.1500 732.6000 250.0500 734.4000 ;
	    RECT 249.0000 731.4000 250.2000 732.6000 ;
	    RECT 253.8000 719.4000 255.0000 720.6000 ;
	    RECT 251.4000 707.4000 252.6000 708.6000 ;
	    RECT 251.5500 702.6000 252.4500 707.4000 ;
	    RECT 246.6000 701.4000 247.8000 702.6000 ;
	    RECT 251.4000 701.4000 252.6000 702.6000 ;
	    RECT 246.7500 696.6000 247.6500 701.4000 ;
	    RECT 246.6000 695.4000 247.8000 696.6000 ;
	    RECT 251.4000 683.4000 252.6000 684.6000 ;
	    RECT 249.0000 680.4000 250.2000 681.6000 ;
	    RECT 249.1500 678.6000 250.0500 680.4000 ;
	    RECT 244.2000 677.4000 245.4000 678.6000 ;
	    RECT 249.0000 677.4000 250.2000 678.6000 ;
	    RECT 246.6000 659.4000 247.8000 660.6000 ;
	    RECT 239.4000 617.4000 240.6000 618.6000 ;
	    RECT 241.8000 617.4000 243.0000 618.6000 ;
	    RECT 237.0000 599.4000 238.2000 600.6000 ;
	    RECT 232.2000 584.4000 233.4000 585.6000 ;
	    RECT 222.6000 581.4000 223.8000 582.6000 ;
	    RECT 225.0000 581.4000 226.2000 582.6000 ;
	    RECT 225.1500 570.6000 226.0500 581.4000 ;
	    RECT 225.0000 569.4000 226.2000 570.6000 ;
	    RECT 241.8000 545.4000 243.0000 546.6000 ;
	    RECT 222.6000 503.4000 223.8000 504.6000 ;
	    RECT 227.4000 503.4000 228.6000 504.6000 ;
	    RECT 220.2000 485.4000 221.4000 486.6000 ;
	    RECT 220.3500 474.6000 221.2500 485.4000 ;
	    RECT 220.2000 473.4000 221.4000 474.6000 ;
	    RECT 217.8000 440.4000 219.0000 441.6000 ;
	    RECT 220.3500 438.6000 221.2500 473.4000 ;
	    RECT 215.4000 437.4000 216.6000 438.6000 ;
	    RECT 220.2000 437.4000 221.4000 438.6000 ;
	    RECT 220.2000 410.4000 221.4000 411.6000 ;
	    RECT 220.3500 384.6000 221.2500 410.4000 ;
	    RECT 220.2000 383.4000 221.4000 384.6000 ;
	    RECT 215.4000 221.4000 216.6000 222.6000 ;
	    RECT 213.0000 215.4000 214.2000 216.6000 ;
	    RECT 215.5500 198.6000 216.4500 221.4000 ;
	    RECT 215.4000 197.4000 216.6000 198.6000 ;
	    RECT 208.2000 185.4000 209.4000 186.6000 ;
	    RECT 181.8000 164.4000 183.0000 165.6000 ;
	    RECT 179.4000 110.4000 180.6000 111.6000 ;
	    RECT 172.2000 98.4000 173.4000 99.6000 ;
	    RECT 148.3500 89.5500 151.6500 90.4500 ;
	    RECT 133.8000 77.4000 135.0000 78.6000 ;
	    RECT 129.0000 74.4000 130.2000 75.6000 ;
	    RECT 129.1500 66.6000 130.0500 74.4000 ;
	    RECT 129.0000 65.4000 130.2000 66.6000 ;
	    RECT 136.2000 66.3000 137.4000 86.7000 ;
	    RECT 138.6000 66.3000 139.8000 86.7000 ;
	    RECT 141.0000 69.3000 142.2000 86.7000 ;
	    RECT 143.4000 83.4000 144.6000 84.6000 ;
	    RECT 143.5500 81.6000 144.4500 83.4000 ;
	    RECT 143.4000 80.4000 144.6000 81.6000 ;
	    RECT 145.8000 69.3000 147.0000 86.7000 ;
	    RECT 148.3500 84.6000 149.2500 89.5500 ;
	    RECT 148.2000 83.4000 149.4000 84.6000 ;
	    RECT 148.3500 57.4500 149.2500 83.4000 ;
	    RECT 150.6000 69.3000 151.8000 86.7000 ;
	    RECT 153.0000 66.3000 154.2000 86.7000 ;
	    RECT 155.4000 66.3000 156.6000 86.7000 ;
	    RECT 157.8000 66.3000 159.0000 86.7000 ;
	    RECT 172.3500 72.6000 173.2500 98.4000 ;
	    RECT 172.2000 71.4000 173.4000 72.6000 ;
	    RECT 126.6000 41.4000 127.8000 42.6000 ;
	    RECT 141.0000 36.3000 142.2000 56.7000 ;
	    RECT 143.4000 36.3000 144.6000 56.7000 ;
	    RECT 145.8000 36.3000 147.0000 56.7000 ;
	    RECT 148.3500 56.5500 151.6500 57.4500 ;
	    RECT 148.2000 36.3000 149.4000 53.7000 ;
	    RECT 150.7500 39.6000 151.6500 56.5500 ;
	    RECT 150.6000 38.4000 151.8000 39.6000 ;
	    RECT 73.8000 11.4000 75.0000 12.6000 ;
	    RECT 141.0000 6.3000 142.2000 26.7000 ;
	    RECT 143.4000 6.3000 144.6000 26.7000 ;
	    RECT 145.8000 6.3000 147.0000 26.7000 ;
	    RECT 148.2000 9.3000 149.4000 26.7000 ;
	    RECT 150.7500 24.6000 151.6500 38.4000 ;
	    RECT 153.0000 36.3000 154.2000 53.7000 ;
	    RECT 155.4000 41.4000 156.6000 42.6000 ;
	    RECT 157.8000 36.3000 159.0000 53.7000 ;
	    RECT 160.2000 36.3000 161.4000 56.7000 ;
	    RECT 162.6000 36.3000 163.8000 56.7000 ;
	    RECT 169.8000 56.4000 171.0000 57.6000 ;
	    RECT 169.9500 48.6000 170.8500 56.4000 ;
	    RECT 181.9500 48.6000 182.8500 164.4000 ;
	    RECT 184.2000 156.3000 185.4000 176.7000 ;
	    RECT 186.6000 156.3000 187.8000 176.7000 ;
	    RECT 189.0000 156.3000 190.2000 173.7000 ;
	    RECT 191.4000 161.4000 192.6000 162.6000 ;
	    RECT 191.4000 155.4000 192.6000 156.6000 ;
	    RECT 193.8000 156.3000 195.0000 173.7000 ;
	    RECT 196.2000 167.4000 197.4000 168.6000 ;
	    RECT 196.3500 159.6000 197.2500 167.4000 ;
	    RECT 196.2000 158.4000 197.4000 159.6000 ;
	    RECT 191.5500 144.6000 192.4500 155.4000 ;
	    RECT 196.3500 144.6000 197.2500 158.4000 ;
	    RECT 198.6000 156.3000 199.8000 173.7000 ;
	    RECT 201.0000 156.3000 202.2000 176.7000 ;
	    RECT 203.4000 156.3000 204.6000 176.7000 ;
	    RECT 205.8000 156.3000 207.0000 176.7000 ;
	    RECT 191.4000 143.4000 192.6000 144.6000 ;
	    RECT 196.2000 143.4000 197.4000 144.6000 ;
	    RECT 215.5500 126.6000 216.4500 197.4000 ;
	    RECT 220.2000 194.4000 221.4000 195.6000 ;
	    RECT 220.3500 171.6000 221.2500 194.4000 ;
	    RECT 220.2000 170.4000 221.4000 171.6000 ;
	    RECT 222.7500 138.6000 223.6500 503.4000 ;
	    RECT 225.0000 440.4000 226.2000 441.6000 ;
	    RECT 225.1500 432.6000 226.0500 440.4000 ;
	    RECT 225.0000 431.4000 226.2000 432.6000 ;
	    RECT 227.5500 366.6000 228.4500 503.4000 ;
	    RECT 229.8000 500.4000 231.0000 501.6000 ;
	    RECT 229.9500 492.6000 230.8500 500.4000 ;
	    RECT 229.8000 491.4000 231.0000 492.6000 ;
	    RECT 241.9500 462.6000 242.8500 545.4000 ;
	    RECT 246.7500 525.6000 247.6500 659.4000 ;
	    RECT 249.1500 642.6000 250.0500 677.4000 ;
	    RECT 249.0000 641.4000 250.2000 642.6000 ;
	    RECT 251.5500 621.6000 252.4500 683.4000 ;
	    RECT 253.9500 645.6000 254.8500 719.4000 ;
	    RECT 256.2000 713.4000 257.4000 714.6000 ;
	    RECT 256.3500 705.6000 257.2500 713.4000 ;
	    RECT 256.2000 704.4000 257.4000 705.6000 ;
	    RECT 261.1500 681.6000 262.0500 866.4000 ;
	    RECT 270.6000 851.4000 271.8000 852.6000 ;
	    RECT 270.7500 804.6000 271.6500 851.4000 ;
	    RECT 273.1500 834.6000 274.0500 947.5500 ;
	    RECT 275.5500 918.6000 276.4500 950.4000 ;
	    RECT 275.4000 917.4000 276.6000 918.6000 ;
	    RECT 273.0000 833.4000 274.2000 834.6000 ;
	    RECT 270.6000 803.4000 271.8000 804.6000 ;
	    RECT 275.4000 755.4000 276.6000 756.6000 ;
	    RECT 263.4000 743.4000 264.6000 744.6000 ;
	    RECT 261.0000 680.4000 262.2000 681.6000 ;
	    RECT 256.2000 674.4000 257.4000 675.6000 ;
	    RECT 256.3500 660.6000 257.2500 674.4000 ;
	    RECT 261.0000 671.4000 262.2000 672.6000 ;
	    RECT 261.1500 660.6000 262.0500 671.4000 ;
	    RECT 256.2000 659.4000 257.4000 660.6000 ;
	    RECT 261.0000 659.4000 262.2000 660.6000 ;
	    RECT 256.2000 653.4000 257.4000 654.6000 ;
	    RECT 253.8000 644.4000 255.0000 645.6000 ;
	    RECT 251.4000 620.4000 252.6000 621.6000 ;
	    RECT 249.0000 617.4000 250.2000 618.6000 ;
	    RECT 246.6000 524.4000 247.8000 525.6000 ;
	    RECT 234.6000 461.4000 235.8000 462.6000 ;
	    RECT 241.8000 461.4000 243.0000 462.6000 ;
	    RECT 244.2000 461.4000 245.4000 462.6000 ;
	    RECT 232.2000 443.4000 233.4000 444.6000 ;
	    RECT 232.3500 411.6000 233.2500 443.4000 ;
	    RECT 232.2000 410.4000 233.4000 411.6000 ;
	    RECT 227.4000 365.4000 228.6000 366.6000 ;
	    RECT 229.8000 341.4000 231.0000 342.6000 ;
	    RECT 229.9500 330.6000 230.8500 341.4000 ;
	    RECT 229.8000 329.4000 231.0000 330.6000 ;
	    RECT 229.9500 261.6000 230.8500 329.4000 ;
	    RECT 232.2000 320.4000 233.4000 321.6000 ;
	    RECT 229.8000 260.4000 231.0000 261.6000 ;
	    RECT 227.4000 167.4000 228.6000 168.6000 ;
	    RECT 222.6000 137.4000 223.8000 138.6000 ;
	    RECT 215.4000 125.4000 216.6000 126.6000 ;
	    RECT 227.5500 117.4500 228.4500 167.4000 ;
	    RECT 229.9500 126.6000 230.8500 260.4000 ;
	    RECT 232.3500 234.6000 233.2500 320.4000 ;
	    RECT 232.2000 233.4000 233.4000 234.6000 ;
	    RECT 232.2000 218.4000 233.4000 219.6000 ;
	    RECT 232.3500 216.6000 233.2500 218.4000 ;
	    RECT 232.2000 215.4000 233.4000 216.6000 ;
	    RECT 232.2000 209.4000 233.4000 210.6000 ;
	    RECT 232.3500 180.6000 233.2500 209.4000 ;
	    RECT 232.2000 179.4000 233.4000 180.6000 ;
	    RECT 229.8000 125.4000 231.0000 126.6000 ;
	    RECT 220.2000 96.3000 221.4000 116.7000 ;
	    RECT 222.6000 96.3000 223.8000 116.7000 ;
	    RECT 225.0000 96.3000 226.2000 116.7000 ;
	    RECT 227.5500 116.5500 230.8500 117.4500 ;
	    RECT 227.4000 96.3000 228.6000 113.7000 ;
	    RECT 229.9500 99.6000 230.8500 116.5500 ;
	    RECT 234.7500 114.6000 235.6500 461.4000 ;
	    RECT 239.4000 323.4000 240.6000 324.6000 ;
	    RECT 239.5500 321.6000 240.4500 323.4000 ;
	    RECT 239.4000 320.4000 240.6000 321.6000 ;
	    RECT 244.3500 222.6000 245.2500 461.4000 ;
	    RECT 246.6000 380.4000 247.8000 381.6000 ;
	    RECT 246.7500 378.6000 247.6500 380.4000 ;
	    RECT 246.6000 377.4000 247.8000 378.6000 ;
	    RECT 249.1500 222.6000 250.0500 617.4000 ;
	    RECT 253.8000 611.4000 255.0000 612.6000 ;
	    RECT 251.4000 605.4000 252.6000 606.6000 ;
	    RECT 251.5500 582.6000 252.4500 605.4000 ;
	    RECT 253.9500 585.6000 254.8500 611.4000 ;
	    RECT 253.8000 584.4000 255.0000 585.6000 ;
	    RECT 251.4000 581.4000 252.6000 582.6000 ;
	    RECT 251.4000 497.4000 252.6000 498.6000 ;
	    RECT 256.3500 465.6000 257.2500 653.4000 ;
	    RECT 258.6000 623.4000 259.8000 624.6000 ;
	    RECT 258.7500 591.6000 259.6500 623.4000 ;
	    RECT 261.1500 612.6000 262.0500 659.4000 ;
	    RECT 261.0000 611.4000 262.2000 612.6000 ;
	    RECT 258.6000 590.4000 259.8000 591.6000 ;
	    RECT 258.6000 581.4000 259.8000 582.6000 ;
	    RECT 258.7500 561.6000 259.6500 581.4000 ;
	    RECT 258.6000 560.4000 259.8000 561.6000 ;
	    RECT 263.5500 498.6000 264.4500 743.4000 ;
	    RECT 270.6000 740.4000 271.8000 741.6000 ;
	    RECT 268.2000 720.4500 269.4000 720.6000 ;
	    RECT 270.7500 720.4500 271.6500 740.4000 ;
	    RECT 275.5500 738.6000 276.4500 755.4000 ;
	    RECT 275.4000 737.4000 276.6000 738.6000 ;
	    RECT 268.2000 719.5500 271.6500 720.4500 ;
	    RECT 268.2000 719.4000 269.4000 719.5500 ;
	    RECT 265.8000 713.4000 267.0000 714.6000 ;
	    RECT 265.9500 708.6000 266.8500 713.4000 ;
	    RECT 265.8000 707.4000 267.0000 708.6000 ;
	    RECT 270.6000 701.4000 271.8000 702.6000 ;
	    RECT 277.9500 690.6000 278.8500 1028.5500 ;
	    RECT 285.1500 1002.6000 286.0500 1049.4000 ;
	    RECT 285.0000 1001.4000 286.2000 1002.6000 ;
	    RECT 282.6000 965.4000 283.8000 966.6000 ;
	    RECT 280.2000 947.4000 281.4000 948.6000 ;
	    RECT 282.7500 945.6000 283.6500 965.4000 ;
	    RECT 285.0000 953.4000 286.2000 954.6000 ;
	    RECT 285.1500 951.6000 286.0500 953.4000 ;
	    RECT 285.0000 950.4000 286.2000 951.6000 ;
	    RECT 287.5500 951.4500 288.4500 1151.4000 ;
	    RECT 289.9500 1146.6000 290.8500 1166.4000 ;
	    RECT 289.8000 1145.4000 291.0000 1146.6000 ;
	    RECT 289.8000 1103.4000 291.0000 1104.6000 ;
	    RECT 289.9500 1098.6000 290.8500 1103.4000 ;
	    RECT 289.8000 1097.4000 291.0000 1098.6000 ;
	    RECT 292.3500 1050.6000 293.2500 1289.4000 ;
	    RECT 311.4000 1283.4000 312.6000 1284.6000 ;
	    RECT 294.6000 1274.4000 295.8000 1275.6000 ;
	    RECT 294.7500 1266.6000 295.6500 1274.4000 ;
	    RECT 311.5500 1266.6000 312.4500 1283.4000 ;
	    RECT 294.6000 1265.4000 295.8000 1266.6000 ;
	    RECT 311.4000 1265.4000 312.6000 1266.6000 ;
	    RECT 294.6000 1262.4000 295.8000 1263.6000 ;
	    RECT 294.7500 1260.6000 295.6500 1262.4000 ;
	    RECT 294.6000 1259.4000 295.8000 1260.6000 ;
	    RECT 297.0000 1253.4000 298.2000 1254.6000 ;
	    RECT 297.1500 1161.6000 298.0500 1253.4000 ;
	    RECT 311.5500 1251.6000 312.4500 1265.4000 ;
	    RECT 311.4000 1250.4000 312.6000 1251.6000 ;
	    RECT 309.0000 1220.4000 310.2000 1221.6000 ;
	    RECT 309.1500 1218.6000 310.0500 1220.4000 ;
	    RECT 309.0000 1217.4000 310.2000 1218.6000 ;
	    RECT 304.2000 1214.4000 305.4000 1215.6000 ;
	    RECT 304.3500 1197.6000 305.2500 1214.4000 ;
	    RECT 309.0000 1199.4000 310.2000 1200.6000 ;
	    RECT 304.2000 1196.4000 305.4000 1197.6000 ;
	    RECT 299.4000 1190.4000 300.6000 1191.6000 ;
	    RECT 299.5500 1164.6000 300.4500 1190.4000 ;
	    RECT 304.2000 1184.4000 305.4000 1185.6000 ;
	    RECT 299.4000 1163.4000 300.6000 1164.6000 ;
	    RECT 297.0000 1160.4000 298.2000 1161.6000 ;
	    RECT 299.5500 1128.6000 300.4500 1163.4000 ;
	    RECT 304.3500 1152.6000 305.2500 1184.4000 ;
	    RECT 306.6000 1160.4000 307.8000 1161.6000 ;
	    RECT 304.2000 1151.4000 305.4000 1152.6000 ;
	    RECT 299.4000 1127.4000 300.6000 1128.6000 ;
	    RECT 304.2000 1127.4000 305.4000 1128.6000 ;
	    RECT 299.4000 1121.4000 300.6000 1122.6000 ;
	    RECT 301.8000 1121.4000 303.0000 1122.6000 ;
	    RECT 294.6000 1100.4000 295.8000 1101.6000 ;
	    RECT 299.5500 1101.4501 300.4500 1121.4000 ;
	    RECT 301.8000 1101.4501 303.0000 1101.6000 ;
	    RECT 299.5500 1100.5500 303.0000 1101.4501 ;
	    RECT 301.8000 1100.4000 303.0000 1100.5500 ;
	    RECT 294.7500 1095.6000 295.6500 1100.4000 ;
	    RECT 299.4000 1097.4000 300.6000 1098.6000 ;
	    RECT 301.8000 1097.4000 303.0000 1098.6000 ;
	    RECT 294.6000 1094.4000 295.8000 1095.6000 ;
	    RECT 299.5500 1080.6000 300.4500 1097.4000 ;
	    RECT 299.4000 1079.4000 300.6000 1080.6000 ;
	    RECT 294.6000 1061.4000 295.8000 1062.6000 ;
	    RECT 292.2000 1049.4000 293.4000 1050.6000 ;
	    RECT 294.7500 1041.6000 295.6500 1061.4000 ;
	    RECT 294.6000 1040.4000 295.8000 1041.6000 ;
	    RECT 292.2000 1037.4000 293.4000 1038.6000 ;
	    RECT 292.3500 1008.6000 293.2500 1037.4000 ;
	    RECT 294.6000 1031.4000 295.8000 1032.6000 ;
	    RECT 292.2000 1007.4000 293.4000 1008.6000 ;
	    RECT 292.2000 1004.4000 293.4000 1005.6000 ;
	    RECT 292.3500 990.6000 293.2500 1004.4000 ;
	    RECT 294.7500 1002.6000 295.6500 1031.4000 ;
	    RECT 294.6000 1001.4000 295.8000 1002.6000 ;
	    RECT 301.9500 990.6000 302.8500 1097.4000 ;
	    RECT 304.3500 1086.6000 305.2500 1127.4000 ;
	    RECT 306.7500 1125.6000 307.6500 1160.4000 ;
	    RECT 309.1500 1158.6000 310.0500 1199.4000 ;
	    RECT 313.9500 1161.6000 314.8500 1400.4000 ;
	    RECT 330.7500 1392.6000 331.6500 1403.4000 ;
	    RECT 316.2000 1391.4000 317.4000 1392.6000 ;
	    RECT 330.6000 1391.4000 331.8000 1392.6000 ;
	    RECT 313.8000 1160.4000 315.0000 1161.6000 ;
	    RECT 309.0000 1157.4000 310.2000 1158.6000 ;
	    RECT 311.4000 1139.4000 312.6000 1140.6000 ;
	    RECT 306.6000 1124.4000 307.8000 1125.6000 ;
	    RECT 304.2000 1085.4000 305.4000 1086.6000 ;
	    RECT 306.6000 1085.4000 307.8000 1086.6000 ;
	    RECT 304.3500 1068.6000 305.2500 1085.4000 ;
	    RECT 304.2000 1067.4000 305.4000 1068.6000 ;
	    RECT 304.2000 1065.4501 305.4000 1065.6000 ;
	    RECT 306.7500 1065.4501 307.6500 1085.4000 ;
	    RECT 304.2000 1064.5500 307.6500 1065.4501 ;
	    RECT 304.2000 1064.4000 305.4000 1064.5500 ;
	    RECT 311.5500 1062.6000 312.4500 1139.4000 ;
	    RECT 313.8000 1109.4000 315.0000 1110.6000 ;
	    RECT 313.9500 1086.6000 314.8500 1109.4000 ;
	    RECT 313.8000 1085.4000 315.0000 1086.6000 ;
	    RECT 311.4000 1061.4000 312.6000 1062.6000 ;
	    RECT 309.0000 1055.4000 310.2000 1056.6000 ;
	    RECT 309.1500 1050.6000 310.0500 1055.4000 ;
	    RECT 309.0000 1049.4000 310.2000 1050.6000 ;
	    RECT 309.1500 1044.6000 310.0500 1049.4000 ;
	    RECT 309.0000 1043.4000 310.2000 1044.6000 ;
	    RECT 313.8000 1043.4000 315.0000 1044.6000 ;
	    RECT 313.9500 1038.6000 314.8500 1043.4000 ;
	    RECT 313.8000 1037.4000 315.0000 1038.6000 ;
	    RECT 304.2000 1025.4000 305.4000 1026.6000 ;
	    RECT 311.4000 1025.4000 312.6000 1026.6000 ;
	    RECT 304.3500 1020.6000 305.2500 1025.4000 ;
	    RECT 304.2000 1019.4000 305.4000 1020.6000 ;
	    RECT 306.6000 1013.4000 307.8000 1014.6000 ;
	    RECT 306.7500 1005.6000 307.6500 1013.4000 ;
	    RECT 311.5500 1005.6000 312.4500 1025.4000 ;
	    RECT 306.6000 1004.4000 307.8000 1005.6000 ;
	    RECT 311.4000 1004.4000 312.6000 1005.6000 ;
	    RECT 292.2000 989.4000 293.4000 990.6000 ;
	    RECT 301.8000 989.4000 303.0000 990.6000 ;
	    RECT 287.5500 950.5500 290.8500 951.4500 ;
	    RECT 282.6000 944.4000 283.8000 945.6000 ;
	    RECT 285.1500 936.6000 286.0500 950.4000 ;
	    RECT 287.4000 947.4000 288.6000 948.6000 ;
	    RECT 285.0000 935.4000 286.2000 936.6000 ;
	    RECT 285.0000 920.4000 286.2000 921.6000 ;
	    RECT 285.1500 846.6000 286.0500 920.4000 ;
	    RECT 287.5500 852.6000 288.4500 947.4000 ;
	    RECT 289.9500 852.6000 290.8500 950.5500 ;
	    RECT 292.3500 942.6000 293.2500 989.4000 ;
	    RECT 301.8000 977.4000 303.0000 978.6000 ;
	    RECT 301.9500 948.6000 302.8500 977.4000 ;
	    RECT 304.2000 974.4000 305.4000 975.6000 ;
	    RECT 297.0000 947.4000 298.2000 948.6000 ;
	    RECT 301.8000 947.4000 303.0000 948.6000 ;
	    RECT 292.2000 941.4000 293.4000 942.6000 ;
	    RECT 292.2000 936.4500 293.4000 936.6000 ;
	    RECT 292.2000 935.5500 295.6500 936.4500 ;
	    RECT 292.2000 935.4000 293.4000 935.5500 ;
	    RECT 294.7500 930.6000 295.6500 935.5500 ;
	    RECT 294.6000 929.4000 295.8000 930.6000 ;
	    RECT 292.2000 923.4000 293.4000 924.6000 ;
	    RECT 292.3500 915.6000 293.2500 923.4000 ;
	    RECT 297.1500 918.6000 298.0500 947.4000 ;
	    RECT 301.8000 920.4000 303.0000 921.6000 ;
	    RECT 294.6000 917.4000 295.8000 918.6000 ;
	    RECT 297.0000 917.4000 298.2000 918.6000 ;
	    RECT 299.4000 917.4000 300.6000 918.6000 ;
	    RECT 292.2000 914.4000 293.4000 915.6000 ;
	    RECT 287.4000 851.4000 288.6000 852.6000 ;
	    RECT 289.8000 851.4000 291.0000 852.6000 ;
	    RECT 287.4000 848.4000 288.6000 849.6000 ;
	    RECT 285.0000 845.4000 286.2000 846.6000 ;
	    RECT 287.5500 825.6000 288.4500 848.4000 ;
	    RECT 292.3500 825.6000 293.2500 914.4000 ;
	    RECT 294.7500 912.6000 295.6500 917.4000 ;
	    RECT 299.5500 915.6000 300.4500 917.4000 ;
	    RECT 299.4000 914.4000 300.6000 915.6000 ;
	    RECT 301.9500 912.6000 302.8500 920.4000 ;
	    RECT 304.3500 918.6000 305.2500 974.4000 ;
	    RECT 304.2000 917.4000 305.4000 918.6000 ;
	    RECT 294.6000 911.4000 295.8000 912.6000 ;
	    RECT 301.8000 911.4000 303.0000 912.6000 ;
	    RECT 299.4000 893.4000 300.6000 894.6000 ;
	    RECT 299.5500 870.6000 300.4500 893.4000 ;
	    RECT 304.2000 887.4000 305.4000 888.6000 ;
	    RECT 299.4000 869.4000 300.6000 870.6000 ;
	    RECT 301.8000 863.4000 303.0000 864.6000 ;
	    RECT 294.6000 845.4000 295.8000 846.6000 ;
	    RECT 287.4000 824.4000 288.6000 825.6000 ;
	    RECT 292.2000 824.4000 293.4000 825.6000 ;
	    RECT 285.0000 800.4000 286.2000 801.6000 ;
	    RECT 280.2000 776.4000 281.4000 777.6000 ;
	    RECT 277.8000 689.4000 279.0000 690.6000 ;
	    RECT 273.0000 683.4000 274.2000 684.6000 ;
	    RECT 270.6000 641.4000 271.8000 642.6000 ;
	    RECT 270.7500 630.6000 271.6500 641.4000 ;
	    RECT 270.6000 629.4000 271.8000 630.6000 ;
	    RECT 268.2000 599.4000 269.4000 600.6000 ;
	    RECT 268.3500 594.6000 269.2500 599.4000 ;
	    RECT 270.6000 596.4000 271.8000 597.6000 ;
	    RECT 268.2000 593.4000 269.4000 594.6000 ;
	    RECT 268.2000 590.4000 269.4000 591.6000 ;
	    RECT 268.3500 501.6000 269.2500 590.4000 ;
	    RECT 270.7500 555.6000 271.6500 596.4000 ;
	    RECT 270.6000 554.4000 271.8000 555.6000 ;
	    RECT 273.1500 546.6000 274.0500 683.4000 ;
	    RECT 275.4000 680.4000 276.6000 681.6000 ;
	    RECT 275.5500 678.6000 276.4500 680.4000 ;
	    RECT 275.4000 677.4000 276.6000 678.6000 ;
	    RECT 277.8000 677.4000 279.0000 678.6000 ;
	    RECT 275.4000 647.4000 276.6000 648.6000 ;
	    RECT 275.5500 642.6000 276.4500 647.4000 ;
	    RECT 275.4000 641.4000 276.6000 642.6000 ;
	    RECT 277.9500 615.6000 278.8500 677.4000 ;
	    RECT 280.3500 645.6000 281.2500 776.4000 ;
	    RECT 285.1500 762.6000 286.0500 800.4000 ;
	    RECT 287.5500 765.6000 288.4500 824.4000 ;
	    RECT 292.3500 822.6000 293.2500 824.4000 ;
	    RECT 294.7500 822.6000 295.6500 845.4000 ;
	    RECT 301.9500 828.6000 302.8500 863.4000 ;
	    RECT 301.8000 827.4000 303.0000 828.6000 ;
	    RECT 289.8000 821.4000 291.0000 822.6000 ;
	    RECT 292.2000 821.4000 293.4000 822.6000 ;
	    RECT 294.6000 821.4000 295.8000 822.6000 ;
	    RECT 287.4000 764.4000 288.6000 765.6000 ;
	    RECT 285.0000 761.4000 286.2000 762.6000 ;
	    RECT 285.0000 758.4000 286.2000 759.6000 ;
	    RECT 285.1500 744.6000 286.0500 758.4000 ;
	    RECT 285.0000 743.4000 286.2000 744.6000 ;
	    RECT 285.0000 740.4000 286.2000 741.6000 ;
	    RECT 287.4000 740.4000 288.6000 741.6000 ;
	    RECT 285.1500 702.6000 286.0500 740.4000 ;
	    RECT 285.0000 701.4000 286.2000 702.6000 ;
	    RECT 285.0000 653.4000 286.2000 654.6000 ;
	    RECT 285.1500 645.6000 286.0500 653.4000 ;
	    RECT 280.2000 644.4000 281.4000 645.6000 ;
	    RECT 285.0000 644.4000 286.2000 645.6000 ;
	    RECT 287.5500 642.6000 288.4500 740.4000 ;
	    RECT 289.9500 720.6000 290.8500 821.4000 ;
	    RECT 299.4000 761.4000 300.6000 762.6000 ;
	    RECT 299.5500 744.6000 300.4500 761.4000 ;
	    RECT 299.4000 743.4000 300.6000 744.6000 ;
	    RECT 292.2000 737.4000 293.4000 738.6000 ;
	    RECT 289.8000 719.4000 291.0000 720.6000 ;
	    RECT 289.8000 647.4000 291.0000 648.6000 ;
	    RECT 289.9500 642.6000 290.8500 647.4000 ;
	    RECT 282.6000 641.4000 283.8000 642.6000 ;
	    RECT 287.4000 641.4000 288.6000 642.6000 ;
	    RECT 289.8000 641.4000 291.0000 642.6000 ;
	    RECT 282.7500 618.6000 283.6500 641.4000 ;
	    RECT 285.0000 620.4000 286.2000 621.6000 ;
	    RECT 282.6000 617.4000 283.8000 618.6000 ;
	    RECT 277.8000 614.4000 279.0000 615.6000 ;
	    RECT 280.2000 593.4000 281.4000 594.6000 ;
	    RECT 280.3500 588.6000 281.2500 593.4000 ;
	    RECT 280.2000 587.4000 281.4000 588.6000 ;
	    RECT 277.8000 584.4000 279.0000 585.6000 ;
	    RECT 280.2000 584.4000 281.4000 585.6000 ;
	    RECT 277.9500 582.6000 278.8500 584.4000 ;
	    RECT 275.4000 581.4000 276.6000 582.6000 ;
	    RECT 277.8000 581.4000 279.0000 582.6000 ;
	    RECT 275.5500 564.6000 276.4500 581.4000 ;
	    RECT 280.3500 576.6000 281.2500 584.4000 ;
	    RECT 280.2000 575.4000 281.4000 576.6000 ;
	    RECT 275.4000 563.4000 276.6000 564.6000 ;
	    RECT 275.4000 557.4000 276.6000 558.6000 ;
	    RECT 273.0000 545.4000 274.2000 546.6000 ;
	    RECT 277.8000 546.3000 279.0000 566.7000 ;
	    RECT 280.2000 546.3000 281.4000 566.7000 ;
	    RECT 282.6000 549.3000 283.8000 566.7000 ;
	    RECT 285.1500 561.6000 286.0500 620.4000 ;
	    RECT 292.3500 600.6000 293.2500 737.4000 ;
	    RECT 301.8000 707.4000 303.0000 708.6000 ;
	    RECT 301.9500 654.6000 302.8500 707.4000 ;
	    RECT 304.3500 657.6000 305.2500 887.4000 ;
	    RECT 306.7500 858.6000 307.6500 1004.4000 ;
	    RECT 316.3500 999.6000 317.2500 1391.4000 ;
	    RECT 333.1500 1317.6000 334.0500 1418.4000 ;
	    RECT 335.4000 1416.3000 336.6000 1433.7001 ;
	    RECT 337.8000 1433.4000 339.0000 1434.6000 ;
	    RECT 337.9500 1422.6000 338.8500 1433.4000 ;
	    RECT 337.8000 1421.4000 339.0000 1422.6000 ;
	    RECT 340.2000 1416.3000 341.4000 1433.7001 ;
	    RECT 342.6000 1416.3000 343.8000 1436.7001 ;
	    RECT 345.0000 1416.3000 346.2000 1436.7001 ;
	    RECT 352.2000 1436.4000 353.4000 1437.6000 ;
	    RECT 352.3500 1428.6000 353.2500 1436.4000 ;
	    RECT 347.4000 1427.4000 348.6000 1428.6000 ;
	    RECT 352.2000 1427.4000 353.4000 1428.6000 ;
	    RECT 376.2000 1427.4000 377.4000 1428.6000 ;
	    RECT 381.0000 1427.4000 382.2000 1428.6000 ;
	    RECT 347.5500 1425.6000 348.4500 1427.4000 ;
	    RECT 347.4000 1424.4000 348.6000 1425.6000 ;
	    RECT 347.5500 1407.6000 348.4500 1424.4000 ;
	    RECT 376.3500 1422.6000 377.2500 1427.4000 ;
	    RECT 376.2000 1421.4000 377.4000 1422.6000 ;
	    RECT 340.2000 1406.4000 341.4000 1407.6000 ;
	    RECT 347.4000 1406.4000 348.6000 1407.6000 ;
	    RECT 333.0000 1316.4000 334.2000 1317.6000 ;
	    RECT 328.2000 1289.4000 329.4000 1290.6000 ;
	    RECT 328.3500 1284.6000 329.2500 1289.4000 ;
	    RECT 328.2000 1283.4000 329.4000 1284.6000 ;
	    RECT 323.4000 1280.4000 324.6000 1281.6000 ;
	    RECT 325.8000 1280.4000 327.0000 1281.6000 ;
	    RECT 323.5500 1278.6000 324.4500 1280.4000 ;
	    RECT 323.4000 1277.4000 324.6000 1278.6000 ;
	    RECT 325.9500 1254.6000 326.8500 1280.4000 ;
	    RECT 337.8000 1274.4000 339.0000 1275.6000 ;
	    RECT 325.8000 1253.4000 327.0000 1254.6000 ;
	    RECT 325.8000 1250.4000 327.0000 1251.6000 ;
	    RECT 325.9500 1224.6000 326.8500 1250.4000 ;
	    RECT 335.4000 1235.4000 336.6000 1236.6000 ;
	    RECT 335.5500 1230.6000 336.4500 1235.4000 ;
	    RECT 335.4000 1229.4000 336.6000 1230.6000 ;
	    RECT 325.8000 1223.4000 327.0000 1224.6000 ;
	    RECT 330.6000 1220.4000 331.8000 1221.6000 ;
	    RECT 323.4000 1169.4000 324.6000 1170.6000 ;
	    RECT 323.5500 1164.6000 324.4500 1169.4000 ;
	    RECT 323.4000 1163.4000 324.6000 1164.6000 ;
	    RECT 328.2000 1124.4000 329.4000 1125.6000 ;
	    RECT 328.3500 1122.6000 329.2500 1124.4000 ;
	    RECT 325.8000 1121.4000 327.0000 1122.6000 ;
	    RECT 328.2000 1121.4000 329.4000 1122.6000 ;
	    RECT 325.9500 1062.6000 326.8500 1121.4000 ;
	    RECT 330.7500 1101.6000 331.6500 1220.4000 ;
	    RECT 337.9500 1218.6000 338.8500 1274.4000 ;
	    RECT 340.3500 1272.6000 341.2500 1406.4000 ;
	    RECT 376.3500 1380.6000 377.2500 1421.4000 ;
	    RECT 381.1500 1410.6000 382.0500 1427.4000 ;
	    RECT 385.9500 1422.6000 386.8500 1460.4000 ;
	    RECT 445.8000 1457.4000 447.0000 1458.6000 ;
	    RECT 441.0000 1454.4000 442.2000 1455.6000 ;
	    RECT 407.4000 1451.4000 408.6000 1452.6000 ;
	    RECT 407.5500 1422.6000 408.4500 1451.4000 ;
	    RECT 441.1500 1446.6000 442.0500 1454.4000 ;
	    RECT 441.0000 1445.4000 442.2000 1446.6000 ;
	    RECT 426.6000 1427.4000 427.8000 1428.6000 ;
	    RECT 385.8000 1421.4000 387.0000 1422.6000 ;
	    RECT 407.4000 1421.4000 408.6000 1422.6000 ;
	    RECT 414.6000 1421.4000 415.8000 1422.6000 ;
	    RECT 381.0000 1409.4000 382.2000 1410.6000 ;
	    RECT 369.0000 1379.4000 370.2000 1380.6000 ;
	    RECT 376.2000 1379.4000 377.4000 1380.6000 ;
	    RECT 354.6000 1376.4000 355.8000 1377.6000 ;
	    RECT 354.7500 1368.6000 355.6500 1376.4000 ;
	    RECT 354.6000 1367.4000 355.8000 1368.6000 ;
	    RECT 359.4000 1364.4000 360.6000 1365.6000 ;
	    RECT 359.5500 1362.6000 360.4500 1364.4000 ;
	    RECT 359.4000 1361.4000 360.6000 1362.6000 ;
	    RECT 361.8000 1356.3000 363.0000 1376.7001 ;
	    RECT 364.2000 1356.3000 365.4000 1376.7001 ;
	    RECT 366.6000 1356.3000 367.8000 1373.7001 ;
	    RECT 369.1500 1362.6000 370.0500 1379.4000 ;
	    RECT 369.0000 1361.4000 370.2000 1362.6000 ;
	    RECT 371.4000 1356.3000 372.6000 1373.7001 ;
	    RECT 373.8000 1358.4000 375.0000 1359.6000 ;
	    RECT 342.6000 1326.3000 343.8000 1346.7001 ;
	    RECT 345.0000 1326.3000 346.2000 1346.7001 ;
	    RECT 347.4000 1326.3000 348.6000 1346.7001 ;
	    RECT 349.8000 1329.3000 351.0000 1346.7001 ;
	    RECT 352.2000 1343.4000 353.4000 1344.6000 ;
	    RECT 352.3500 1320.6000 353.2500 1343.4000 ;
	    RECT 354.6000 1329.3000 355.8000 1346.7001 ;
	    RECT 357.0000 1340.4000 358.2000 1341.6000 ;
	    RECT 352.2000 1319.4000 353.4000 1320.6000 ;
	    RECT 349.8000 1316.4000 351.0000 1317.6000 ;
	    RECT 340.2000 1271.4000 341.4000 1272.6000 ;
	    RECT 340.2000 1236.3000 341.4000 1256.7001 ;
	    RECT 342.6000 1236.3000 343.8000 1256.7001 ;
	    RECT 345.0000 1236.3000 346.2000 1256.7001 ;
	    RECT 347.4000 1236.3000 348.6000 1253.7001 ;
	    RECT 349.9500 1239.6000 350.8500 1316.4000 ;
	    RECT 357.1500 1302.6000 358.0500 1340.4000 ;
	    RECT 359.4000 1329.3000 360.6000 1346.7001 ;
	    RECT 359.4000 1325.4000 360.6000 1326.6000 ;
	    RECT 361.8000 1326.3000 363.0000 1346.7001 ;
	    RECT 364.2000 1326.3000 365.4000 1346.7001 ;
	    RECT 366.6000 1337.4000 367.8000 1338.6000 ;
	    RECT 371.4000 1335.4501 372.6000 1335.6000 ;
	    RECT 369.1500 1334.5500 372.6000 1335.4501 ;
	    RECT 359.5500 1320.6000 360.4500 1325.4000 ;
	    RECT 359.4000 1319.4000 360.6000 1320.6000 ;
	    RECT 357.0000 1301.4000 358.2000 1302.6000 ;
	    RECT 354.6000 1280.4000 355.8000 1281.6000 ;
	    RECT 349.8000 1238.4000 351.0000 1239.6000 ;
	    RECT 345.0000 1220.4000 346.2000 1221.6000 ;
	    RECT 345.1500 1218.6000 346.0500 1220.4000 ;
	    RECT 337.8000 1217.4000 339.0000 1218.6000 ;
	    RECT 345.0000 1217.4000 346.2000 1218.6000 ;
	    RECT 349.9500 1212.6000 350.8500 1238.4000 ;
	    RECT 352.2000 1236.3000 353.4000 1253.7001 ;
	    RECT 354.7500 1242.6000 355.6500 1280.4000 ;
	    RECT 359.4000 1277.4000 360.6000 1278.6000 ;
	    RECT 364.2000 1271.4000 365.4000 1272.6000 ;
	    RECT 354.6000 1241.4000 355.8000 1242.6000 ;
	    RECT 357.0000 1236.3000 358.2000 1253.7001 ;
	    RECT 359.4000 1236.3000 360.6000 1256.7001 ;
	    RECT 361.8000 1236.3000 363.0000 1256.7001 ;
	    RECT 364.3500 1245.6000 365.2500 1271.4000 ;
	    RECT 369.1500 1260.6000 370.0500 1334.5500 ;
	    RECT 371.4000 1334.4000 372.6000 1334.5500 ;
	    RECT 373.9500 1317.6000 374.8500 1358.4000 ;
	    RECT 376.2000 1356.3000 377.4000 1373.7001 ;
	    RECT 378.6000 1356.3000 379.8000 1376.7001 ;
	    RECT 381.0000 1356.3000 382.2000 1376.7001 ;
	    RECT 383.4000 1356.3000 384.6000 1376.7001 ;
	    RECT 373.8000 1316.4000 375.0000 1317.6000 ;
	    RECT 373.9500 1314.6000 374.8500 1316.4000 ;
	    RECT 373.8000 1313.4000 375.0000 1314.6000 ;
	    RECT 381.0000 1310.4000 382.2000 1311.6000 ;
	    RECT 378.6000 1277.4000 379.8000 1278.6000 ;
	    RECT 369.0000 1259.4000 370.2000 1260.6000 ;
	    RECT 369.0000 1256.4000 370.2000 1257.6000 ;
	    RECT 369.1500 1248.6000 370.0500 1256.4000 ;
	    RECT 369.0000 1247.4000 370.2000 1248.6000 ;
	    RECT 364.2000 1244.4000 365.4000 1245.6000 ;
	    RECT 357.0000 1214.4000 358.2000 1215.6000 ;
	    RECT 349.8000 1211.4000 351.0000 1212.6000 ;
	    RECT 357.1500 1191.6000 358.0500 1214.4000 ;
	    RECT 361.8000 1211.4000 363.0000 1212.6000 ;
	    RECT 359.4000 1196.4000 360.6000 1197.6000 ;
	    RECT 357.0000 1190.4000 358.2000 1191.6000 ;
	    RECT 345.0000 1175.4000 346.2000 1176.6000 ;
	    RECT 333.0000 1127.4000 334.2000 1128.6000 ;
	    RECT 330.6000 1100.4000 331.8000 1101.6000 ;
	    RECT 328.2000 1067.4000 329.4000 1068.6000 ;
	    RECT 328.3500 1065.6000 329.2500 1067.4000 ;
	    RECT 333.1500 1065.6000 334.0500 1127.4000 ;
	    RECT 345.1500 1125.6000 346.0500 1175.4000 ;
	    RECT 345.0000 1124.4000 346.2000 1125.6000 ;
	    RECT 335.4000 1121.4000 336.6000 1122.6000 ;
	    RECT 357.1500 1119.6000 358.0500 1190.4000 ;
	    RECT 357.0000 1118.4000 358.2000 1119.6000 ;
	    RECT 337.8000 1109.4000 339.0000 1110.6000 ;
	    RECT 337.9500 1101.6000 338.8500 1109.4000 ;
	    RECT 357.1500 1104.6000 358.0500 1118.4000 ;
	    RECT 340.2000 1103.4000 341.4000 1104.6000 ;
	    RECT 357.0000 1103.4000 358.2000 1104.6000 ;
	    RECT 337.8000 1100.4000 339.0000 1101.6000 ;
	    RECT 340.3500 1098.6000 341.2500 1103.4000 ;
	    RECT 357.0000 1100.4000 358.2000 1101.6000 ;
	    RECT 340.2000 1097.4000 341.4000 1098.6000 ;
	    RECT 352.2000 1097.4000 353.4000 1098.6000 ;
	    RECT 335.4000 1067.4000 336.6000 1068.6000 ;
	    RECT 328.2000 1064.4000 329.4000 1065.6000 ;
	    RECT 333.0000 1064.4000 334.2000 1065.6000 ;
	    RECT 325.8000 1061.4000 327.0000 1062.6000 ;
	    RECT 335.5500 1032.6000 336.4500 1067.4000 ;
	    RECT 337.8000 1058.4000 339.0000 1059.6000 ;
	    RECT 337.9500 1044.6000 338.8500 1058.4000 ;
	    RECT 337.8000 1043.4000 339.0000 1044.6000 ;
	    RECT 340.2000 1043.4000 341.4000 1044.6000 ;
	    RECT 340.3500 1038.6000 341.2500 1043.4000 ;
	    RECT 347.4000 1040.4000 348.6000 1041.6000 ;
	    RECT 337.8000 1037.4000 339.0000 1038.6000 ;
	    RECT 340.2000 1037.4000 341.4000 1038.6000 ;
	    RECT 345.0000 1038.4501 346.2000 1038.6000 ;
	    RECT 347.5500 1038.4501 348.4500 1040.4000 ;
	    RECT 345.0000 1037.5500 348.4500 1038.4501 ;
	    RECT 345.0000 1037.4000 346.2000 1037.5500 ;
	    RECT 349.8000 1037.4000 351.0000 1038.6000 ;
	    RECT 335.4000 1031.4000 336.6000 1032.6000 ;
	    RECT 335.5500 1020.6000 336.4500 1031.4000 ;
	    RECT 335.4000 1019.4000 336.6000 1020.6000 ;
	    RECT 316.2000 998.4000 317.4000 999.6000 ;
	    RECT 316.3500 978.6000 317.2500 998.4000 ;
	    RECT 313.8000 977.4000 315.0000 978.6000 ;
	    RECT 316.2000 977.4000 317.4000 978.6000 ;
	    RECT 313.9500 972.6000 314.8500 977.4000 ;
	    RECT 313.8000 971.4000 315.0000 972.6000 ;
	    RECT 313.9500 966.6000 314.8500 971.4000 ;
	    RECT 337.9500 966.6000 338.8500 1037.4000 ;
	    RECT 349.9500 1026.6000 350.8500 1037.4000 ;
	    RECT 349.8000 1025.4000 351.0000 1026.6000 ;
	    RECT 309.0000 965.4000 310.2000 966.6000 ;
	    RECT 313.8000 965.4000 315.0000 966.6000 ;
	    RECT 337.8000 965.4000 339.0000 966.6000 ;
	    RECT 309.1500 948.6000 310.0500 965.4000 ;
	    RECT 309.0000 947.4000 310.2000 948.6000 ;
	    RECT 311.4000 947.4000 312.6000 948.6000 ;
	    RECT 309.0000 941.4000 310.2000 942.6000 ;
	    RECT 306.6000 857.4000 307.8000 858.6000 ;
	    RECT 309.1500 705.6000 310.0500 941.4000 ;
	    RECT 311.5500 906.6000 312.4500 947.4000 ;
	    RECT 313.9500 942.6000 314.8500 965.4000 ;
	    RECT 349.8000 959.4000 351.0000 960.6000 ;
	    RECT 349.9500 951.6000 350.8500 959.4000 ;
	    RECT 316.2000 950.4000 317.4000 951.6000 ;
	    RECT 318.6000 950.4000 319.8000 951.6000 ;
	    RECT 328.2000 950.4000 329.4000 951.6000 ;
	    RECT 349.8000 950.4000 351.0000 951.6000 ;
	    RECT 313.8000 941.4000 315.0000 942.6000 ;
	    RECT 313.9500 924.6000 314.8500 941.4000 ;
	    RECT 316.3500 936.6000 317.2500 950.4000 ;
	    RECT 318.7500 945.6000 319.6500 950.4000 ;
	    RECT 321.0000 947.4000 322.2000 948.6000 ;
	    RECT 318.6000 944.4000 319.8000 945.6000 ;
	    RECT 316.2000 935.4000 317.4000 936.6000 ;
	    RECT 318.7500 930.6000 319.6500 944.4000 ;
	    RECT 321.1500 942.6000 322.0500 947.4000 ;
	    RECT 321.0000 941.4000 322.2000 942.6000 ;
	    RECT 318.6000 929.4000 319.8000 930.6000 ;
	    RECT 313.8000 923.4000 315.0000 924.6000 ;
	    RECT 328.3500 921.6000 329.2500 950.4000 ;
	    RECT 342.6000 947.4000 343.8000 948.6000 ;
	    RECT 333.0000 923.4000 334.2000 924.6000 ;
	    RECT 328.2000 920.4000 329.4000 921.6000 ;
	    RECT 333.1500 918.6000 334.0500 923.4000 ;
	    RECT 342.7500 921.6000 343.6500 947.4000 ;
	    RECT 347.4000 944.4000 348.6000 945.6000 ;
	    RECT 347.5500 936.6000 348.4500 944.4000 ;
	    RECT 347.4000 935.4000 348.6000 936.6000 ;
	    RECT 342.6000 920.4000 343.8000 921.6000 ;
	    RECT 333.0000 917.4000 334.2000 918.6000 ;
	    RECT 352.3500 915.6000 353.2500 1097.4000 ;
	    RECT 357.1500 1041.6000 358.0500 1100.4000 ;
	    RECT 357.0000 1040.4000 358.2000 1041.6000 ;
	    RECT 357.0000 1025.4000 358.2000 1026.6000 ;
	    RECT 357.1500 948.6000 358.0500 1025.4000 ;
	    RECT 357.0000 947.4000 358.2000 948.6000 ;
	    RECT 354.6000 938.4000 355.8000 939.6000 ;
	    RECT 352.2000 914.4000 353.4000 915.6000 ;
	    RECT 311.4000 905.4000 312.6000 906.6000 ;
	    RECT 311.5500 849.6000 312.4500 905.4000 ;
	    RECT 323.4000 876.3000 324.6000 896.7000 ;
	    RECT 325.8000 876.3000 327.0000 896.7000 ;
	    RECT 328.2000 876.3000 329.4000 896.7000 ;
	    RECT 330.6000 876.3000 331.8000 893.7000 ;
	    RECT 333.0000 878.4000 334.2000 879.6000 ;
	    RECT 333.1500 870.6000 334.0500 878.4000 ;
	    RECT 335.4000 876.3000 336.6000 893.7000 ;
	    RECT 337.8000 881.4000 339.0000 882.6000 ;
	    RECT 333.0000 869.4000 334.2000 870.6000 ;
	    RECT 333.1500 864.6000 334.0500 869.4000 ;
	    RECT 337.9500 867.6000 338.8500 881.4000 ;
	    RECT 340.2000 876.3000 341.4000 893.7000 ;
	    RECT 342.6000 876.3000 343.8000 896.7000 ;
	    RECT 345.0000 876.3000 346.2000 896.7000 ;
	    RECT 352.2000 896.4000 353.4000 897.6000 ;
	    RECT 352.3500 888.6000 353.2500 896.4000 ;
	    RECT 347.4000 887.4000 348.6000 888.6000 ;
	    RECT 352.2000 887.4000 353.4000 888.6000 ;
	    RECT 347.5500 885.6000 348.4500 887.4000 ;
	    RECT 347.4000 884.4000 348.6000 885.6000 ;
	    RECT 352.2000 869.4000 353.4000 870.6000 ;
	    RECT 337.8000 866.4000 339.0000 867.6000 ;
	    RECT 333.0000 863.4000 334.2000 864.6000 ;
	    RECT 342.6000 851.4000 343.8000 852.6000 ;
	    RECT 311.4000 848.4000 312.6000 849.6000 ;
	    RECT 342.7500 822.6000 343.6500 851.4000 ;
	    RECT 347.4000 824.4000 348.6000 825.6000 ;
	    RECT 318.6000 821.4000 319.8000 822.6000 ;
	    RECT 323.4000 821.4000 324.6000 822.6000 ;
	    RECT 340.2000 821.4000 341.4000 822.6000 ;
	    RECT 342.6000 821.4000 343.8000 822.6000 ;
	    RECT 318.7500 810.6000 319.6500 821.4000 ;
	    RECT 318.6000 809.4000 319.8000 810.6000 ;
	    RECT 323.5500 801.6000 324.4500 821.4000 ;
	    RECT 347.5500 801.6000 348.4500 824.4000 ;
	    RECT 349.8000 821.4000 351.0000 822.6000 ;
	    RECT 349.9500 810.6000 350.8500 821.4000 ;
	    RECT 349.8000 809.4000 351.0000 810.6000 ;
	    RECT 323.4000 800.4000 324.6000 801.6000 ;
	    RECT 347.4000 800.4000 348.6000 801.6000 ;
	    RECT 316.2000 743.4000 317.4000 744.6000 ;
	    RECT 316.3500 726.6000 317.2500 743.4000 ;
	    RECT 316.2000 725.4000 317.4000 726.6000 ;
	    RECT 347.4000 713.4000 348.6000 714.6000 ;
	    RECT 347.5500 708.6000 348.4500 713.4000 ;
	    RECT 347.4000 707.4000 348.6000 708.6000 ;
	    RECT 309.0000 704.4000 310.2000 705.6000 ;
	    RECT 313.8000 704.4000 315.0000 705.6000 ;
	    RECT 309.1500 660.6000 310.0500 704.4000 ;
	    RECT 311.4000 701.4000 312.6000 702.6000 ;
	    RECT 311.5500 696.6000 312.4500 701.4000 ;
	    RECT 311.4000 695.4000 312.6000 696.6000 ;
	    RECT 313.9500 666.6000 314.8500 704.4000 ;
	    RECT 349.9500 702.6000 350.8500 809.4000 ;
	    RECT 352.3500 777.6000 353.2500 869.4000 ;
	    RECT 354.7500 798.6000 355.6500 938.4000 ;
	    RECT 357.0000 914.4000 358.2000 915.6000 ;
	    RECT 357.1500 888.6000 358.0500 914.4000 ;
	    RECT 357.0000 887.4000 358.2000 888.6000 ;
	    RECT 357.1500 840.6000 358.0500 887.4000 ;
	    RECT 357.0000 839.4000 358.2000 840.6000 ;
	    RECT 354.6000 797.4000 355.8000 798.6000 ;
	    RECT 352.2000 776.4000 353.4000 777.6000 ;
	    RECT 352.3500 738.6000 353.2500 776.4000 ;
	    RECT 354.6000 740.4000 355.8000 741.6000 ;
	    RECT 352.2000 737.4000 353.4000 738.6000 ;
	    RECT 354.7500 708.6000 355.6500 740.4000 ;
	    RECT 357.1500 738.6000 358.0500 839.4000 ;
	    RECT 359.5500 819.4500 360.4500 1196.4000 ;
	    RECT 361.9500 939.6000 362.8500 1211.4000 ;
	    RECT 364.3500 1161.6000 365.2500 1244.4000 ;
	    RECT 369.0000 1223.4000 370.2000 1224.6000 ;
	    RECT 364.2000 1161.4501 365.4000 1161.6000 ;
	    RECT 364.2000 1160.5500 367.6500 1161.4501 ;
	    RECT 364.2000 1160.4000 365.4000 1160.5500 ;
	    RECT 364.2000 1151.4000 365.4000 1152.6000 ;
	    RECT 364.3500 1119.6000 365.2500 1151.4000 ;
	    RECT 364.2000 1118.4000 365.4000 1119.6000 ;
	    RECT 364.3500 1050.6000 365.2500 1118.4000 ;
	    RECT 364.2000 1049.4000 365.4000 1050.6000 ;
	    RECT 361.8000 938.4000 363.0000 939.6000 ;
	    RECT 361.8000 935.4000 363.0000 936.6000 ;
	    RECT 361.9500 918.6000 362.8500 935.4000 ;
	    RECT 364.2000 923.4000 365.4000 924.6000 ;
	    RECT 361.8000 917.4000 363.0000 918.6000 ;
	    RECT 364.3500 915.6000 365.2500 923.4000 ;
	    RECT 364.2000 914.4000 365.4000 915.6000 ;
	    RECT 366.7500 894.6000 367.6500 1160.5500 ;
	    RECT 366.6000 893.4000 367.8000 894.6000 ;
	    RECT 369.1500 879.6000 370.0500 1223.4000 ;
	    RECT 378.7500 1221.6000 379.6500 1277.4000 ;
	    RECT 381.1500 1224.6000 382.0500 1310.4000 ;
	    RECT 385.9500 1281.6000 386.8500 1421.4000 ;
	    RECT 426.7500 1419.6000 427.6500 1427.4000 ;
	    RECT 426.6000 1418.4000 427.8000 1419.6000 ;
	    RECT 429.0000 1397.4000 430.2000 1398.6000 ;
	    RECT 397.8000 1379.4000 399.0000 1380.6000 ;
	    RECT 397.9500 1371.6000 398.8500 1379.4000 ;
	    RECT 397.8000 1370.4000 399.0000 1371.6000 ;
	    RECT 429.1500 1362.6000 430.0500 1397.4000 ;
	    RECT 445.9500 1374.6000 446.8500 1457.4000 ;
	    RECT 448.2000 1446.3000 449.4000 1466.7001 ;
	    RECT 450.6000 1446.3000 451.8000 1466.7001 ;
	    RECT 453.0000 1449.3000 454.2000 1466.7001 ;
	    RECT 455.4000 1460.4000 456.6000 1461.6000 ;
	    RECT 455.5500 1452.6000 456.4500 1460.4000 ;
	    RECT 455.4000 1451.4000 456.6000 1452.6000 ;
	    RECT 457.8000 1449.3000 459.0000 1466.7001 ;
	    RECT 460.2000 1463.4000 461.4000 1464.6000 ;
	    RECT 460.3500 1446.4501 461.2500 1463.4000 ;
	    RECT 462.6000 1449.3000 463.8000 1466.7001 ;
	    RECT 460.3500 1445.5500 463.6500 1446.4501 ;
	    RECT 465.0000 1446.3000 466.2000 1466.7001 ;
	    RECT 467.4000 1446.3000 468.6000 1466.7001 ;
	    RECT 469.8000 1446.3000 471.0000 1466.7001 ;
	    RECT 510.6000 1460.4000 511.8000 1461.6000 ;
	    RECT 537.0000 1460.4000 538.2000 1461.6000 ;
	    RECT 544.2000 1460.4000 545.4000 1461.6000 ;
	    RECT 505.8000 1454.4000 507.0000 1455.6000 ;
	    RECT 491.4000 1451.4000 492.6000 1452.6000 ;
	    RECT 457.8000 1424.4000 459.0000 1425.6000 ;
	    RECT 457.9500 1401.6000 458.8500 1424.4000 ;
	    RECT 460.2000 1421.4000 461.4000 1422.6000 ;
	    RECT 460.2000 1415.4000 461.4000 1416.6000 ;
	    RECT 457.8000 1400.4000 459.0000 1401.6000 ;
	    RECT 455.4000 1391.4000 456.6000 1392.6000 ;
	    RECT 431.4000 1373.4000 432.6000 1374.6000 ;
	    RECT 445.8000 1373.4000 447.0000 1374.6000 ;
	    RECT 400.2000 1361.4000 401.4000 1362.6000 ;
	    RECT 429.0000 1361.4000 430.2000 1362.6000 ;
	    RECT 400.3500 1296.6000 401.2500 1361.4000 ;
	    RECT 417.0000 1358.4000 418.2000 1359.6000 ;
	    RECT 417.1500 1356.6000 418.0500 1358.4000 ;
	    RECT 417.0000 1355.4000 418.2000 1356.6000 ;
	    RECT 405.0000 1301.4000 406.2000 1302.6000 ;
	    RECT 400.2000 1295.4000 401.4000 1296.6000 ;
	    RECT 405.1500 1281.6000 406.0500 1301.4000 ;
	    RECT 414.6000 1283.4000 415.8000 1284.6000 ;
	    RECT 383.4000 1280.4000 384.6000 1281.6000 ;
	    RECT 385.8000 1280.4000 387.0000 1281.6000 ;
	    RECT 405.0000 1280.4000 406.2000 1281.6000 ;
	    RECT 412.2000 1280.4000 413.4000 1281.6000 ;
	    RECT 381.0000 1223.4000 382.2000 1224.6000 ;
	    RECT 378.6000 1220.4000 379.8000 1221.6000 ;
	    RECT 383.5500 1218.6000 384.4500 1280.4000 ;
	    RECT 395.4000 1277.4000 396.6000 1278.6000 ;
	    RECT 409.8000 1277.4000 411.0000 1278.6000 ;
	    RECT 395.5500 1275.6000 396.4500 1277.4000 ;
	    RECT 395.4000 1274.4000 396.6000 1275.6000 ;
	    RECT 393.0000 1265.4000 394.2000 1266.6000 ;
	    RECT 393.1500 1245.6000 394.0500 1265.4000 ;
	    RECT 400.2000 1259.4000 401.4000 1260.6000 ;
	    RECT 393.0000 1244.4000 394.2000 1245.6000 ;
	    RECT 385.8000 1229.4000 387.0000 1230.6000 ;
	    RECT 385.9500 1218.6000 386.8500 1229.4000 ;
	    RECT 390.6000 1220.4000 391.8000 1221.6000 ;
	    RECT 390.7500 1218.6000 391.6500 1220.4000 ;
	    RECT 383.4000 1217.4000 384.6000 1218.6000 ;
	    RECT 385.8000 1217.4000 387.0000 1218.6000 ;
	    RECT 390.6000 1217.4000 391.8000 1218.6000 ;
	    RECT 378.6000 1157.4000 379.8000 1158.6000 ;
	    RECT 378.7500 1140.6000 379.6500 1157.4000 ;
	    RECT 378.6000 1139.4000 379.8000 1140.6000 ;
	    RECT 390.6000 1121.4000 391.8000 1122.6000 ;
	    RECT 376.2000 1115.4000 377.4000 1116.6000 ;
	    RECT 376.3500 1104.6000 377.2500 1115.4000 ;
	    RECT 376.2000 1103.4000 377.4000 1104.6000 ;
	    RECT 385.8000 1103.4000 387.0000 1104.6000 ;
	    RECT 385.9500 1074.6000 386.8500 1103.4000 ;
	    RECT 390.7500 1101.6000 391.6500 1121.4000 ;
	    RECT 388.2000 1100.4000 389.4000 1101.6000 ;
	    RECT 390.6000 1100.4000 391.8000 1101.6000 ;
	    RECT 388.3500 1098.6000 389.2500 1100.4000 ;
	    RECT 388.2000 1097.4000 389.4000 1098.6000 ;
	    RECT 385.8000 1073.4000 387.0000 1074.6000 ;
	    RECT 385.9500 1071.6000 386.8500 1073.4000 ;
	    RECT 385.8000 1070.4000 387.0000 1071.6000 ;
	    RECT 381.0000 1067.4000 382.2000 1068.6000 ;
	    RECT 390.7500 1062.6000 391.6500 1100.4000 ;
	    RECT 373.8000 1061.4000 375.0000 1062.6000 ;
	    RECT 390.6000 1061.4000 391.8000 1062.6000 ;
	    RECT 373.8000 977.4000 375.0000 978.6000 ;
	    RECT 371.4000 959.4000 372.6000 960.6000 ;
	    RECT 371.5500 912.6000 372.4500 959.4000 ;
	    RECT 373.9500 954.6000 374.8500 977.4000 ;
	    RECT 381.0000 969.3000 382.2000 986.7000 ;
	    RECT 390.6000 977.4000 391.8000 978.6000 ;
	    RECT 385.8000 959.4000 387.0000 960.6000 ;
	    RECT 373.8000 953.4000 375.0000 954.6000 ;
	    RECT 381.0000 953.4000 382.2000 954.6000 ;
	    RECT 378.6000 950.4000 379.8000 951.6000 ;
	    RECT 373.8000 944.4000 375.0000 945.6000 ;
	    RECT 371.4000 911.4000 372.6000 912.6000 ;
	    RECT 373.9500 900.6000 374.8500 944.4000 ;
	    RECT 378.7500 936.6000 379.6500 950.4000 ;
	    RECT 381.1500 945.6000 382.0500 953.4000 ;
	    RECT 385.9500 948.6000 386.8500 959.4000 ;
	    RECT 390.7500 948.6000 391.6500 977.4000 ;
	    RECT 393.1500 960.6000 394.0500 1244.4000 ;
	    RECT 400.3500 1242.6000 401.2500 1259.4000 ;
	    RECT 400.2000 1241.4000 401.4000 1242.6000 ;
	    RECT 400.3500 1221.4501 401.2500 1241.4000 ;
	    RECT 407.4000 1238.4000 408.6000 1239.6000 ;
	    RECT 400.3500 1220.5500 403.6500 1221.4501 ;
	    RECT 400.2000 1097.4000 401.4000 1098.6000 ;
	    RECT 395.4000 969.3000 396.6000 986.7000 ;
	    RECT 397.8000 983.4000 399.0000 984.6000 ;
	    RECT 397.9500 981.6000 398.8500 983.4000 ;
	    RECT 397.8000 980.4000 399.0000 981.6000 ;
	    RECT 400.2000 975.3000 401.4000 983.7000 ;
	    RECT 393.0000 959.4000 394.2000 960.6000 ;
	    RECT 393.0000 953.4000 394.2000 954.6000 ;
	    RECT 385.8000 947.4000 387.0000 948.6000 ;
	    RECT 388.2000 947.4000 389.4000 948.6000 ;
	    RECT 390.6000 947.4000 391.8000 948.6000 ;
	    RECT 381.0000 944.4000 382.2000 945.6000 ;
	    RECT 378.6000 935.4000 379.8000 936.6000 ;
	    RECT 378.7500 921.6000 379.6500 935.4000 ;
	    RECT 385.9500 924.6000 386.8500 947.4000 ;
	    RECT 388.3500 924.6000 389.2500 947.4000 ;
	    RECT 393.1500 924.6000 394.0500 953.4000 ;
	    RECT 402.7500 948.6000 403.6500 1220.5500 ;
	    RECT 407.5500 1170.6000 408.4500 1238.4000 ;
	    RECT 407.4000 1169.4000 408.6000 1170.6000 ;
	    RECT 407.5500 1014.6000 408.4500 1169.4000 ;
	    RECT 409.8000 1031.4000 411.0000 1032.6000 ;
	    RECT 407.4000 1013.4000 408.6000 1014.6000 ;
	    RECT 409.8000 950.4000 411.0000 951.6000 ;
	    RECT 402.6000 947.4000 403.8000 948.6000 ;
	    RECT 385.8000 923.4000 387.0000 924.6000 ;
	    RECT 388.2000 923.4000 389.4000 924.6000 ;
	    RECT 393.0000 923.4000 394.2000 924.6000 ;
	    RECT 378.6000 920.4000 379.8000 921.6000 ;
	    RECT 409.9500 915.6000 410.8500 950.4000 ;
	    RECT 409.8000 914.4000 411.0000 915.6000 ;
	    RECT 373.8000 899.4000 375.0000 900.6000 ;
	    RECT 409.8000 899.4000 411.0000 900.6000 ;
	    RECT 371.4000 893.4000 372.6000 894.6000 ;
	    RECT 364.2000 878.4000 365.4000 879.6000 ;
	    RECT 369.0000 878.4000 370.2000 879.6000 ;
	    RECT 361.8000 819.4500 363.0000 819.6000 ;
	    RECT 359.5500 818.5500 363.0000 819.4500 ;
	    RECT 361.8000 818.4000 363.0000 818.5500 ;
	    RECT 359.4000 803.4000 360.6000 804.6000 ;
	    RECT 359.5500 762.6000 360.4500 803.4000 ;
	    RECT 361.9500 774.6000 362.8500 818.4000 ;
	    RECT 361.8000 773.4000 363.0000 774.6000 ;
	    RECT 359.4000 761.4000 360.6000 762.6000 ;
	    RECT 361.9500 759.6000 362.8500 773.4000 ;
	    RECT 361.8000 758.4000 363.0000 759.6000 ;
	    RECT 361.8000 755.4000 363.0000 756.6000 ;
	    RECT 361.9500 750.6000 362.8500 755.4000 ;
	    RECT 361.8000 749.4000 363.0000 750.6000 ;
	    RECT 357.0000 737.4000 358.2000 738.6000 ;
	    RECT 354.6000 707.4000 355.8000 708.6000 ;
	    RECT 352.2000 704.4000 353.4000 705.6000 ;
	    RECT 316.2000 701.4000 317.4000 702.6000 ;
	    RECT 325.8000 701.4000 327.0000 702.6000 ;
	    RECT 340.2000 701.4000 341.4000 702.6000 ;
	    RECT 349.8000 701.4000 351.0000 702.6000 ;
	    RECT 316.3500 684.6000 317.2500 701.4000 ;
	    RECT 318.6000 698.4000 319.8000 699.6000 ;
	    RECT 318.7500 696.6000 319.6500 698.4000 ;
	    RECT 318.6000 695.4000 319.8000 696.6000 ;
	    RECT 316.2000 683.4000 317.4000 684.6000 ;
	    RECT 313.8000 665.4000 315.0000 666.6000 ;
	    RECT 309.0000 659.4000 310.2000 660.6000 ;
	    RECT 304.2000 656.4000 305.4000 657.6000 ;
	    RECT 301.8000 653.4000 303.0000 654.6000 ;
	    RECT 309.1500 642.6000 310.0500 659.4000 ;
	    RECT 311.4000 656.4000 312.6000 657.6000 ;
	    RECT 297.0000 641.4000 298.2000 642.6000 ;
	    RECT 309.0000 641.4000 310.2000 642.6000 ;
	    RECT 297.1500 621.6000 298.0500 641.4000 ;
	    RECT 306.6000 638.4000 307.8000 639.6000 ;
	    RECT 297.0000 620.4000 298.2000 621.6000 ;
	    RECT 292.2000 599.4000 293.4000 600.6000 ;
	    RECT 297.1500 582.6000 298.0500 620.4000 ;
	    RECT 304.2000 605.4000 305.4000 606.6000 ;
	    RECT 287.4000 582.4500 288.6000 582.6000 ;
	    RECT 287.4000 581.5500 290.8500 582.4500 ;
	    RECT 287.4000 581.4000 288.6000 581.5500 ;
	    RECT 289.9500 576.6000 290.8500 581.5500 ;
	    RECT 297.0000 581.4000 298.2000 582.6000 ;
	    RECT 289.8000 575.4000 291.0000 576.6000 ;
	    RECT 301.8000 569.4000 303.0000 570.6000 ;
	    RECT 285.0000 560.4000 286.2000 561.6000 ;
	    RECT 287.4000 549.3000 288.6000 566.7000 ;
	    RECT 289.8000 563.4000 291.0000 564.6000 ;
	    RECT 282.6000 503.4000 283.8000 504.6000 ;
	    RECT 268.2000 500.4000 269.4000 501.6000 ;
	    RECT 273.0000 500.4000 274.2000 501.6000 ;
	    RECT 263.4000 497.4000 264.6000 498.6000 ;
	    RECT 265.8000 497.4000 267.0000 498.6000 ;
	    RECT 270.6000 497.4000 271.8000 498.6000 ;
	    RECT 261.0000 485.4000 262.2000 486.6000 ;
	    RECT 261.1500 465.6000 262.0500 485.4000 ;
	    RECT 265.9500 468.6000 266.8500 497.4000 ;
	    RECT 265.8000 467.4000 267.0000 468.6000 ;
	    RECT 256.2000 464.4000 257.4000 465.6000 ;
	    RECT 261.0000 464.4000 262.2000 465.6000 ;
	    RECT 256.3500 438.6000 257.2500 464.4000 ;
	    RECT 258.6000 461.4000 259.8000 462.6000 ;
	    RECT 263.4000 461.4000 264.6000 462.6000 ;
	    RECT 258.7500 444.6000 259.6500 461.4000 ;
	    RECT 258.6000 443.4000 259.8000 444.6000 ;
	    RECT 263.5500 441.6000 264.4500 461.4000 ;
	    RECT 268.2000 455.4000 269.4000 456.6000 ;
	    RECT 268.3500 444.6000 269.2500 455.4000 ;
	    RECT 268.2000 443.4000 269.4000 444.6000 ;
	    RECT 263.4000 440.4000 264.6000 441.6000 ;
	    RECT 268.2000 440.4000 269.4000 441.6000 ;
	    RECT 256.2000 437.4000 257.4000 438.6000 ;
	    RECT 268.3500 432.6000 269.2500 440.4000 ;
	    RECT 270.7500 438.6000 271.6500 497.4000 ;
	    RECT 273.1500 492.6000 274.0500 500.4000 ;
	    RECT 273.0000 491.4000 274.2000 492.6000 ;
	    RECT 275.4000 467.4000 276.6000 468.6000 ;
	    RECT 273.0000 464.4000 274.2000 465.6000 ;
	    RECT 273.1500 441.6000 274.0500 464.4000 ;
	    RECT 273.0000 440.4000 274.2000 441.6000 ;
	    RECT 275.5500 438.6000 276.4500 467.4000 ;
	    RECT 270.6000 437.4000 271.8000 438.6000 ;
	    RECT 275.4000 437.4000 276.6000 438.6000 ;
	    RECT 268.2000 431.4000 269.4000 432.6000 ;
	    RECT 270.7500 417.6000 271.6500 437.4000 ;
	    RECT 280.2000 431.4000 281.4000 432.6000 ;
	    RECT 270.6000 416.4000 271.8000 417.6000 ;
	    RECT 275.4000 410.4000 276.6000 411.6000 ;
	    RECT 275.5500 396.6000 276.4500 410.4000 ;
	    RECT 275.4000 395.4000 276.6000 396.6000 ;
	    RECT 270.6000 383.4000 271.8000 384.6000 ;
	    RECT 270.7500 381.6000 271.6500 383.4000 ;
	    RECT 270.6000 380.4000 271.8000 381.6000 ;
	    RECT 273.0000 380.4000 274.2000 381.6000 ;
	    RECT 273.1500 378.6000 274.0500 380.4000 ;
	    RECT 273.0000 377.4000 274.2000 378.6000 ;
	    RECT 256.2000 365.4000 257.4000 366.6000 ;
	    RECT 256.3500 324.6000 257.2500 365.4000 ;
	    RECT 273.1500 324.6000 274.0500 377.4000 ;
	    RECT 280.3500 342.6000 281.2500 431.4000 ;
	    RECT 280.2000 341.4000 281.4000 342.6000 ;
	    RECT 256.2000 323.4000 257.4000 324.6000 ;
	    RECT 273.0000 323.4000 274.2000 324.6000 ;
	    RECT 253.8000 260.4000 255.0000 261.6000 ;
	    RECT 251.4000 257.4000 252.6000 258.6000 ;
	    RECT 244.2000 221.4000 245.4000 222.6000 ;
	    RECT 249.0000 221.4000 250.2000 222.6000 ;
	    RECT 246.6000 185.4000 247.8000 186.6000 ;
	    RECT 229.8000 98.4000 231.0000 99.6000 ;
	    RECT 165.0000 47.4000 166.2000 48.6000 ;
	    RECT 169.8000 47.4000 171.0000 48.6000 ;
	    RECT 181.8000 47.4000 183.0000 48.6000 ;
	    RECT 165.1500 45.6000 166.0500 47.4000 ;
	    RECT 165.0000 44.4000 166.2000 45.6000 ;
	    RECT 229.9500 42.6000 230.8500 98.4000 ;
	    RECT 232.2000 96.3000 233.4000 113.7000 ;
	    RECT 234.6000 113.4000 235.8000 114.6000 ;
	    RECT 234.6000 101.4000 235.8000 102.6000 ;
	    RECT 237.0000 96.3000 238.2000 113.7000 ;
	    RECT 239.4000 96.3000 240.6000 116.7000 ;
	    RECT 241.8000 96.3000 243.0000 116.7000 ;
	    RECT 244.2000 113.4000 245.4000 114.6000 ;
	    RECT 244.3500 105.6000 245.2500 113.4000 ;
	    RECT 244.2000 104.4000 245.4000 105.6000 ;
	    RECT 244.3500 78.6000 245.2500 104.4000 ;
	    RECT 246.7500 102.6000 247.6500 185.4000 ;
	    RECT 251.5500 168.6000 252.4500 257.4000 ;
	    RECT 253.9500 246.6000 254.8500 260.4000 ;
	    RECT 253.8000 245.4000 255.0000 246.6000 ;
	    RECT 253.8000 218.4000 255.0000 219.6000 ;
	    RECT 251.4000 167.4000 252.6000 168.6000 ;
	    RECT 249.0000 161.4000 250.2000 162.6000 ;
	    RECT 253.9500 156.6000 254.8500 218.4000 ;
	    RECT 256.3500 168.6000 257.2500 323.4000 ;
	    RECT 273.1500 321.6000 274.0500 323.4000 ;
	    RECT 273.0000 320.4000 274.2000 321.6000 ;
	    RECT 268.2000 263.4000 269.4000 264.6000 ;
	    RECT 268.3500 219.6000 269.2500 263.4000 ;
	    RECT 268.2000 218.4000 269.4000 219.6000 ;
	    RECT 256.2000 167.4000 257.4000 168.6000 ;
	    RECT 253.8000 155.4000 255.0000 156.6000 ;
	    RECT 249.0000 116.4000 250.2000 117.6000 ;
	    RECT 249.1500 108.6000 250.0500 116.4000 ;
	    RECT 249.0000 107.4000 250.2000 108.6000 ;
	    RECT 246.6000 101.4000 247.8000 102.6000 ;
	    RECT 244.2000 77.4000 245.4000 78.6000 ;
	    RECT 253.9500 51.6000 254.8500 155.4000 ;
	    RECT 253.8000 50.4000 255.0000 51.6000 ;
	    RECT 229.8000 41.4000 231.0000 42.6000 ;
	    RECT 150.6000 23.4000 151.8000 24.6000 ;
	    RECT 153.0000 9.3000 154.2000 26.7000 ;
	    RECT 155.4000 23.4000 156.6000 24.6000 ;
	    RECT 155.5500 21.6000 156.4500 23.4000 ;
	    RECT 155.4000 20.4000 156.6000 21.6000 ;
	    RECT 157.8000 9.3000 159.0000 26.7000 ;
	    RECT 160.2000 6.3000 161.4000 26.7000 ;
	    RECT 162.6000 6.3000 163.8000 26.7000 ;
	    RECT 165.0000 17.4000 166.2000 18.6000 ;
	    RECT 169.8000 14.4000 171.0000 15.6000 ;
	    RECT 169.9500 6.6000 170.8500 14.4000 ;
	    RECT 256.3500 12.6000 257.2500 167.4000 ;
	    RECT 270.6000 164.4000 271.8000 165.6000 ;
	    RECT 270.7500 129.6000 271.6500 164.4000 ;
	    RECT 273.1500 162.6000 274.0500 320.4000 ;
	    RECT 280.2000 317.4000 281.4000 318.6000 ;
	    RECT 280.3500 255.6000 281.2500 317.4000 ;
	    RECT 282.7500 315.6000 283.6500 503.4000 ;
	    RECT 289.9500 492.6000 290.8500 563.4000 ;
	    RECT 292.2000 549.3000 293.4000 566.7000 ;
	    RECT 294.6000 546.3000 295.8000 566.7000 ;
	    RECT 297.0000 546.3000 298.2000 566.7000 ;
	    RECT 299.4000 546.3000 300.6000 566.7000 ;
	    RECT 294.6000 539.4000 295.8000 540.6000 ;
	    RECT 289.8000 491.4000 291.0000 492.6000 ;
	    RECT 294.7500 462.6000 295.6500 539.4000 ;
	    RECT 301.9500 528.6000 302.8500 569.4000 ;
	    RECT 304.3500 558.6000 305.2500 605.4000 ;
	    RECT 306.7500 588.6000 307.6500 638.4000 ;
	    RECT 306.6000 587.4000 307.8000 588.6000 ;
	    RECT 304.2000 557.4000 305.4000 558.6000 ;
	    RECT 301.8000 527.4000 303.0000 528.6000 ;
	    RECT 306.7500 525.6000 307.6500 587.4000 ;
	    RECT 301.8000 524.4000 303.0000 525.6000 ;
	    RECT 306.6000 524.4000 307.8000 525.6000 ;
	    RECT 297.0000 500.4000 298.2000 501.6000 ;
	    RECT 297.1500 480.6000 298.0500 500.4000 ;
	    RECT 299.4000 497.4000 300.6000 498.6000 ;
	    RECT 299.4000 491.4000 300.6000 492.6000 ;
	    RECT 297.0000 479.4000 298.2000 480.6000 ;
	    RECT 294.6000 461.4000 295.8000 462.6000 ;
	    RECT 287.4000 458.4000 288.6000 459.6000 ;
	    RECT 287.5500 456.6000 288.4500 458.4000 ;
	    RECT 287.4000 455.4000 288.6000 456.6000 ;
	    RECT 285.0000 419.4000 286.2000 420.6000 ;
	    RECT 282.6000 314.4000 283.8000 315.6000 ;
	    RECT 282.6000 260.4000 283.8000 261.6000 ;
	    RECT 280.2000 254.4000 281.4000 255.6000 ;
	    RECT 273.0000 161.4000 274.2000 162.6000 ;
	    RECT 280.2000 140.4000 281.4000 141.6000 ;
	    RECT 270.6000 128.4000 271.8000 129.6000 ;
	    RECT 277.8000 125.4000 279.0000 126.6000 ;
	    RECT 277.9500 102.6000 278.8500 125.4000 ;
	    RECT 280.3500 105.6000 281.2500 140.4000 ;
	    RECT 280.2000 104.4000 281.4000 105.6000 ;
	    RECT 277.8000 101.4000 279.0000 102.6000 ;
	    RECT 282.7500 48.6000 283.6500 260.4000 ;
	    RECT 285.1500 225.6000 286.0500 419.4000 ;
	    RECT 287.4000 395.4000 288.6000 396.6000 ;
	    RECT 289.8000 396.3000 291.0000 416.7000 ;
	    RECT 292.2000 396.3000 293.4000 416.7000 ;
	    RECT 294.6000 396.3000 295.8000 416.7000 ;
	    RECT 297.0000 396.3000 298.2000 413.7000 ;
	    RECT 299.5500 408.6000 300.4500 491.4000 ;
	    RECT 301.9500 459.6000 302.8500 524.4000 ;
	    RECT 306.6000 515.4000 307.8000 516.6000 ;
	    RECT 306.7500 501.6000 307.6500 515.4000 ;
	    RECT 306.6000 500.4000 307.8000 501.6000 ;
	    RECT 309.0000 500.4000 310.2000 501.6000 ;
	    RECT 309.1500 498.6000 310.0500 500.4000 ;
	    RECT 309.0000 497.4000 310.2000 498.6000 ;
	    RECT 304.2000 494.4000 305.4000 495.6000 ;
	    RECT 304.3500 486.6000 305.2500 494.4000 ;
	    RECT 304.2000 485.4000 305.4000 486.6000 ;
	    RECT 301.8000 458.4000 303.0000 459.6000 ;
	    RECT 301.9500 420.6000 302.8500 458.4000 ;
	    RECT 309.0000 440.4000 310.2000 441.6000 ;
	    RECT 309.1500 432.6000 310.0500 440.4000 ;
	    RECT 309.0000 431.4000 310.2000 432.6000 ;
	    RECT 311.5500 426.6000 312.4500 656.4000 ;
	    RECT 313.9500 618.6000 314.8500 665.4000 ;
	    RECT 325.9500 648.6000 326.8500 701.4000 ;
	    RECT 340.2000 671.4000 341.4000 672.6000 ;
	    RECT 323.4000 647.4000 324.6000 648.6000 ;
	    RECT 325.8000 647.4000 327.0000 648.6000 ;
	    RECT 323.5500 645.6000 324.4500 647.4000 ;
	    RECT 323.4000 644.4000 324.6000 645.6000 ;
	    RECT 321.0000 641.4000 322.2000 642.6000 ;
	    RECT 337.8000 641.4000 339.0000 642.6000 ;
	    RECT 321.1500 630.6000 322.0500 641.4000 ;
	    RECT 321.0000 629.4000 322.2000 630.6000 ;
	    RECT 330.6000 629.4000 331.8000 630.6000 ;
	    RECT 316.2000 623.4000 317.4000 624.6000 ;
	    RECT 313.8000 617.4000 315.0000 618.6000 ;
	    RECT 316.3500 564.6000 317.2500 623.4000 ;
	    RECT 330.7500 618.6000 331.6500 629.4000 ;
	    RECT 330.6000 617.4000 331.8000 618.6000 ;
	    RECT 321.0000 599.4000 322.2000 600.6000 ;
	    RECT 316.2000 563.4000 317.4000 564.6000 ;
	    RECT 316.3500 552.6000 317.2500 563.4000 ;
	    RECT 316.2000 551.4000 317.4000 552.6000 ;
	    RECT 316.3500 504.6000 317.2500 551.4000 ;
	    RECT 316.2000 503.4000 317.4000 504.6000 ;
	    RECT 318.6000 479.4000 319.8000 480.6000 ;
	    RECT 316.2000 473.4000 317.4000 474.6000 ;
	    RECT 313.8000 443.4000 315.0000 444.6000 ;
	    RECT 311.4000 425.4000 312.6000 426.6000 ;
	    RECT 313.9500 420.6000 314.8500 443.4000 ;
	    RECT 316.3500 435.6000 317.2500 473.4000 ;
	    RECT 316.2000 434.4000 317.4000 435.6000 ;
	    RECT 316.2000 425.4000 317.4000 426.6000 ;
	    RECT 301.8000 419.4000 303.0000 420.6000 ;
	    RECT 313.8000 419.4000 315.0000 420.6000 ;
	    RECT 299.4000 407.4000 300.6000 408.6000 ;
	    RECT 299.5500 399.6000 300.4500 407.4000 ;
	    RECT 299.4000 398.4000 300.6000 399.6000 ;
	    RECT 301.8000 396.3000 303.0000 413.7000 ;
	    RECT 304.2000 401.4000 305.4000 402.6000 ;
	    RECT 287.5500 375.6000 288.4500 395.4000 ;
	    RECT 289.8000 389.4000 291.0000 390.6000 ;
	    RECT 287.4000 374.4000 288.6000 375.6000 ;
	    RECT 287.4000 344.4000 288.6000 345.6000 ;
	    RECT 287.5500 306.6000 288.4500 344.4000 ;
	    RECT 287.4000 305.4000 288.6000 306.6000 ;
	    RECT 285.0000 224.4000 286.2000 225.6000 ;
	    RECT 289.9500 171.6000 290.8500 389.4000 ;
	    RECT 304.3500 384.6000 305.2500 401.4000 ;
	    RECT 306.6000 396.3000 307.8000 413.7000 ;
	    RECT 309.0000 396.3000 310.2000 416.7000 ;
	    RECT 311.4000 396.3000 312.6000 416.7000 ;
	    RECT 313.8000 405.4500 315.0000 405.6000 ;
	    RECT 316.3500 405.4500 317.2500 425.4000 ;
	    RECT 318.6000 416.4000 319.8000 417.6000 ;
	    RECT 318.7500 408.6000 319.6500 416.4000 ;
	    RECT 318.6000 407.4000 319.8000 408.6000 ;
	    RECT 313.8000 404.5500 317.2500 405.4500 ;
	    RECT 313.8000 404.4000 315.0000 404.5500 ;
	    RECT 304.2000 383.4000 305.4000 384.6000 ;
	    RECT 301.8000 380.4000 303.0000 381.6000 ;
	    RECT 301.9500 378.6000 302.8500 380.4000 ;
	    RECT 301.8000 377.4000 303.0000 378.6000 ;
	    RECT 294.6000 371.4000 295.8000 372.6000 ;
	    RECT 294.7500 339.6000 295.6500 371.4000 ;
	    RECT 301.9500 342.6000 302.8500 377.4000 ;
	    RECT 301.8000 341.4000 303.0000 342.6000 ;
	    RECT 294.6000 338.4000 295.8000 339.6000 ;
	    RECT 301.9500 264.6000 302.8500 341.4000 ;
	    RECT 306.6000 338.4000 307.8000 339.6000 ;
	    RECT 306.7500 315.6000 307.6500 338.4000 ;
	    RECT 306.6000 314.4000 307.8000 315.6000 ;
	    RECT 301.8000 264.4500 303.0000 264.6000 ;
	    RECT 299.5500 263.5500 303.0000 264.4500 ;
	    RECT 299.5500 261.6000 300.4500 263.5500 ;
	    RECT 301.8000 263.4000 303.0000 263.5500 ;
	    RECT 292.2000 260.4000 293.4000 261.6000 ;
	    RECT 299.4000 260.4000 300.6000 261.6000 ;
	    RECT 289.8000 170.4000 291.0000 171.6000 ;
	    RECT 289.9500 168.6000 290.8500 170.4000 ;
	    RECT 289.8000 167.4000 291.0000 168.6000 ;
	    RECT 285.0000 164.4000 286.2000 165.6000 ;
	    RECT 285.1500 108.6000 286.0500 164.4000 ;
	    RECT 292.3500 144.6000 293.2500 260.4000 ;
	    RECT 313.9500 252.6000 314.8500 404.4000 ;
	    RECT 316.2000 389.4000 317.4000 390.6000 ;
	    RECT 316.3500 384.6000 317.2500 389.4000 ;
	    RECT 316.2000 383.4000 317.4000 384.6000 ;
	    RECT 316.2000 377.4000 317.4000 378.6000 ;
	    RECT 316.3500 366.6000 317.2500 377.4000 ;
	    RECT 316.2000 365.4000 317.4000 366.6000 ;
	    RECT 318.6000 347.4000 319.8000 348.6000 ;
	    RECT 318.7500 345.6000 319.6500 347.4000 ;
	    RECT 318.6000 344.4000 319.8000 345.6000 ;
	    RECT 313.8000 251.4000 315.0000 252.6000 ;
	    RECT 321.1500 246.6000 322.0500 599.4000 ;
	    RECT 337.9500 585.6000 338.8500 641.4000 ;
	    RECT 340.3500 639.6000 341.2500 671.4000 ;
	    RECT 345.0000 647.4000 346.2000 648.6000 ;
	    RECT 340.2000 638.4000 341.4000 639.6000 ;
	    RECT 340.2000 623.4000 341.4000 624.6000 ;
	    RECT 337.8000 584.4000 339.0000 585.6000 ;
	    RECT 340.3500 582.6000 341.2500 623.4000 ;
	    RECT 342.6000 617.4000 343.8000 618.6000 ;
	    RECT 342.7500 585.6000 343.6500 617.4000 ;
	    RECT 347.4000 587.4000 348.6000 588.6000 ;
	    RECT 342.6000 584.4000 343.8000 585.6000 ;
	    RECT 335.4000 581.4000 336.6000 582.6000 ;
	    RECT 340.2000 581.4000 341.4000 582.6000 ;
	    RECT 345.0000 581.4000 346.2000 582.6000 ;
	    RECT 330.6000 563.4000 331.8000 564.6000 ;
	    RECT 335.5500 561.6000 336.4500 581.4000 ;
	    RECT 335.4000 560.4000 336.6000 561.6000 ;
	    RECT 345.1500 558.6000 346.0500 581.4000 ;
	    RECT 347.5500 576.6000 348.4500 587.4000 ;
	    RECT 349.8000 581.4000 351.0000 582.6000 ;
	    RECT 347.4000 575.4000 348.6000 576.6000 ;
	    RECT 330.6000 557.4000 331.8000 558.6000 ;
	    RECT 340.2000 557.4000 341.4000 558.6000 ;
	    RECT 345.0000 557.4000 346.2000 558.6000 ;
	    RECT 328.2000 551.4000 329.4000 552.6000 ;
	    RECT 323.4000 533.4000 324.6000 534.6000 ;
	    RECT 323.5500 468.6000 324.4500 533.4000 ;
	    RECT 328.3500 522.6000 329.2500 551.4000 ;
	    RECT 328.2000 521.4000 329.4000 522.6000 ;
	    RECT 323.4000 467.4000 324.6000 468.6000 ;
	    RECT 323.5500 345.6000 324.4500 467.4000 ;
	    RECT 328.3500 462.6000 329.2500 521.4000 ;
	    RECT 330.7500 501.6000 331.6500 557.4000 ;
	    RECT 337.8000 545.4000 339.0000 546.6000 ;
	    RECT 335.4000 536.4000 336.6000 537.6000 ;
	    RECT 335.5500 528.6000 336.4500 536.4000 ;
	    RECT 335.4000 527.4000 336.6000 528.6000 ;
	    RECT 337.9500 507.4500 338.8500 545.4000 ;
	    RECT 340.3500 534.6000 341.2500 557.4000 ;
	    RECT 340.2000 533.4000 341.4000 534.6000 ;
	    RECT 340.2000 527.4000 341.4000 528.6000 ;
	    RECT 340.3500 525.6000 341.2500 527.4000 ;
	    RECT 340.2000 524.4000 341.4000 525.6000 ;
	    RECT 342.6000 516.3000 343.8000 536.7000 ;
	    RECT 345.0000 516.3000 346.2000 536.7000 ;
	    RECT 347.4000 516.3000 348.6000 533.7000 ;
	    RECT 349.9500 528.6000 350.8500 581.4000 ;
	    RECT 352.3500 546.6000 353.2500 704.4000 ;
	    RECT 354.6000 701.4000 355.8000 702.6000 ;
	    RECT 354.7500 561.6000 355.6500 701.4000 ;
	    RECT 364.3500 675.6000 365.2500 878.4000 ;
	    RECT 369.0000 854.4000 370.2000 855.6000 ;
	    RECT 369.1500 846.6000 370.0500 854.4000 ;
	    RECT 369.0000 845.4000 370.2000 846.6000 ;
	    RECT 366.6000 833.4000 367.8000 834.6000 ;
	    RECT 366.7500 828.6000 367.6500 833.4000 ;
	    RECT 371.5500 831.4500 372.4500 893.4000 ;
	    RECT 373.9500 870.6000 374.8500 899.4000 ;
	    RECT 385.8000 887.4000 387.0000 888.6000 ;
	    RECT 385.9500 885.6000 386.8500 887.4000 ;
	    RECT 409.9500 885.6000 410.8500 899.4000 ;
	    RECT 385.8000 884.4000 387.0000 885.6000 ;
	    RECT 409.8000 884.4000 411.0000 885.6000 ;
	    RECT 412.3500 882.6000 413.2500 1280.4000 ;
	    RECT 414.7500 1275.6000 415.6500 1283.4000 ;
	    RECT 414.6000 1274.4000 415.8000 1275.6000 ;
	    RECT 417.1500 1239.6000 418.0500 1355.4000 ;
	    RECT 429.0000 1331.4000 430.2000 1332.6000 ;
	    RECT 429.1500 1275.6000 430.0500 1331.4000 ;
	    RECT 429.0000 1274.4000 430.2000 1275.6000 ;
	    RECT 419.4000 1271.4000 420.6000 1272.6000 ;
	    RECT 419.5500 1245.6000 420.4500 1271.4000 ;
	    RECT 419.4000 1244.4000 420.6000 1245.6000 ;
	    RECT 417.0000 1238.4000 418.2000 1239.6000 ;
	    RECT 419.4000 1238.4000 420.6000 1239.6000 ;
	    RECT 419.5500 1212.6000 420.4500 1238.4000 ;
	    RECT 426.6000 1229.4000 427.8000 1230.6000 ;
	    RECT 419.4000 1211.4000 420.6000 1212.6000 ;
	    RECT 419.5500 1185.6000 420.4500 1211.4000 ;
	    RECT 419.4000 1184.4000 420.6000 1185.6000 ;
	    RECT 414.6000 1154.4000 415.8000 1155.6000 ;
	    RECT 414.7500 1122.6000 415.6500 1154.4000 ;
	    RECT 417.0000 1127.4000 418.2000 1128.6000 ;
	    RECT 414.6000 1121.4000 415.8000 1122.6000 ;
	    RECT 417.1500 1116.6000 418.0500 1127.4000 ;
	    RECT 426.7500 1125.6000 427.6500 1229.4000 ;
	    RECT 431.5500 1146.6000 432.4500 1373.4000 ;
	    RECT 460.3500 1368.6000 461.2500 1415.4000 ;
	    RECT 462.7500 1404.6000 463.6500 1445.5500 ;
	    RECT 491.5500 1428.6000 492.4500 1451.4000 ;
	    RECT 505.9500 1446.6000 506.8500 1454.4000 ;
	    RECT 505.8000 1445.4000 507.0000 1446.6000 ;
	    RECT 491.4000 1427.4000 492.6000 1428.6000 ;
	    RECT 472.2000 1421.4000 473.4000 1422.6000 ;
	    RECT 474.6000 1421.4000 475.8000 1422.6000 ;
	    RECT 479.4000 1421.4000 480.6000 1422.6000 ;
	    RECT 472.3500 1410.6000 473.2500 1421.4000 ;
	    RECT 472.2000 1409.4000 473.4000 1410.6000 ;
	    RECT 462.6000 1403.4000 463.8000 1404.6000 ;
	    RECT 457.8000 1367.4000 459.0000 1368.6000 ;
	    RECT 460.2000 1367.4000 461.4000 1368.6000 ;
	    RECT 457.9500 1362.6000 458.8500 1367.4000 ;
	    RECT 479.5500 1362.6000 480.4500 1421.4000 ;
	    RECT 505.9500 1416.6000 506.8500 1445.4000 ;
	    RECT 508.2000 1440.4501 509.4000 1440.6000 ;
	    RECT 510.7500 1440.4501 511.6500 1460.4000 ;
	    RECT 537.1500 1440.6000 538.0500 1460.4000 ;
	    RECT 508.2000 1439.5500 511.6500 1440.4501 ;
	    RECT 508.2000 1439.4000 509.4000 1439.5500 ;
	    RECT 537.0000 1439.4000 538.2000 1440.6000 ;
	    RECT 541.8000 1440.4501 543.0000 1440.6000 ;
	    RECT 544.3500 1440.4501 545.2500 1460.4000 ;
	    RECT 611.4000 1457.4000 612.6000 1458.6000 ;
	    RECT 652.2000 1457.4000 653.4000 1458.6000 ;
	    RECT 688.2000 1457.4000 689.4000 1458.6000 ;
	    RECT 541.8000 1439.5500 545.2500 1440.4501 ;
	    RECT 541.8000 1439.4000 543.0000 1439.5500 ;
	    RECT 561.0000 1424.4000 562.2000 1425.6000 ;
	    RECT 561.1500 1422.6000 562.0500 1424.4000 ;
	    RECT 561.0000 1421.4000 562.2000 1422.6000 ;
	    RECT 505.8000 1415.4000 507.0000 1416.6000 ;
	    RECT 568.2000 1416.3000 569.4000 1433.7001 ;
	    RECT 577.8000 1424.4000 579.0000 1425.6000 ;
	    RECT 577.9500 1416.6000 578.8500 1424.4000 ;
	    RECT 577.8000 1415.4000 579.0000 1416.6000 ;
	    RECT 582.6000 1416.3000 583.8000 1433.7001 ;
	    RECT 585.0000 1421.4000 586.2000 1422.6000 ;
	    RECT 496.2000 1409.4000 497.4000 1410.6000 ;
	    RECT 481.8000 1386.3000 483.0000 1406.7001 ;
	    RECT 484.2000 1386.3000 485.4000 1406.7001 ;
	    RECT 486.6000 1386.3000 487.8000 1406.7001 ;
	    RECT 489.0000 1389.3000 490.2000 1406.7001 ;
	    RECT 491.4000 1403.4000 492.6000 1404.6000 ;
	    RECT 457.8000 1361.4000 459.0000 1362.6000 ;
	    RECT 479.4000 1361.4000 480.6000 1362.6000 ;
	    RECT 489.0000 1361.4000 490.2000 1362.6000 ;
	    RECT 457.8000 1358.4000 459.0000 1359.6000 ;
	    RECT 457.9500 1332.6000 458.8500 1358.4000 ;
	    RECT 457.8000 1331.4000 459.0000 1332.6000 ;
	    RECT 460.2000 1319.4000 461.4000 1320.6000 ;
	    RECT 436.2000 1296.3000 437.4000 1316.7001 ;
	    RECT 438.6000 1296.3000 439.8000 1316.7001 ;
	    RECT 441.0000 1296.3000 442.2000 1316.7001 ;
	    RECT 443.4000 1296.3000 444.6000 1313.7001 ;
	    RECT 445.8000 1313.4000 447.0000 1314.6000 ;
	    RECT 445.9500 1299.6000 446.8500 1313.4000 ;
	    RECT 445.8000 1298.4000 447.0000 1299.6000 ;
	    RECT 448.2000 1296.3000 449.4000 1313.7001 ;
	    RECT 450.6000 1301.4000 451.8000 1302.6000 ;
	    RECT 453.0000 1296.3000 454.2000 1313.7001 ;
	    RECT 455.4000 1296.3000 456.6000 1316.7001 ;
	    RECT 457.8000 1296.3000 459.0000 1316.7001 ;
	    RECT 460.3500 1305.6000 461.2500 1319.4000 ;
	    RECT 465.0000 1316.4000 466.2000 1317.6000 ;
	    RECT 465.1500 1308.6000 466.0500 1316.4000 ;
	    RECT 465.0000 1307.4000 466.2000 1308.6000 ;
	    RECT 472.2000 1307.4000 473.4000 1308.6000 ;
	    RECT 472.3500 1305.6000 473.2500 1307.4000 ;
	    RECT 460.2000 1304.4000 461.4000 1305.6000 ;
	    RECT 472.2000 1304.4000 473.4000 1305.6000 ;
	    RECT 453.0000 1280.4000 454.2000 1281.6000 ;
	    RECT 453.1500 1248.6000 454.0500 1280.4000 ;
	    RECT 453.0000 1247.4000 454.2000 1248.6000 ;
	    RECT 453.1500 1242.6000 454.0500 1247.4000 ;
	    RECT 453.0000 1241.4000 454.2000 1242.6000 ;
	    RECT 453.1500 1221.4501 454.0500 1241.4000 ;
	    RECT 450.7500 1220.5500 454.0500 1221.4501 ;
	    RECT 431.4000 1145.4000 432.6000 1146.6000 ;
	    RECT 443.4000 1133.4000 444.6000 1134.6000 ;
	    RECT 450.7500 1134.4501 451.6500 1220.5500 ;
	    RECT 460.3500 1200.6000 461.2500 1304.4000 ;
	    RECT 479.5500 1302.6000 480.4500 1361.4000 ;
	    RECT 489.1500 1350.6000 490.0500 1361.4000 ;
	    RECT 489.0000 1349.4000 490.2000 1350.6000 ;
	    RECT 491.5500 1314.6000 492.4500 1403.4000 ;
	    RECT 493.8000 1389.3000 495.0000 1406.7001 ;
	    RECT 496.3500 1401.6000 497.2500 1409.4000 ;
	    RECT 585.1500 1407.6000 586.0500 1421.4000 ;
	    RECT 587.4000 1419.3000 588.6000 1427.7001 ;
	    RECT 611.5500 1422.6000 612.4500 1457.4000 ;
	    RECT 649.8000 1427.4000 651.0000 1428.6000 ;
	    RECT 613.8000 1424.4000 615.0000 1425.6000 ;
	    RECT 652.3500 1425.4501 653.2500 1457.4000 ;
	    RECT 683.4000 1454.4000 684.6000 1455.6000 ;
	    RECT 683.5500 1443.6000 684.4500 1454.4000 ;
	    RECT 683.4000 1442.4000 684.6000 1443.6000 ;
	    RECT 654.6000 1439.4000 655.8000 1440.6000 ;
	    RECT 649.9500 1424.5500 653.2500 1425.4501 ;
	    RECT 589.8000 1421.4000 591.0000 1422.6000 ;
	    RECT 606.6000 1421.4000 607.8000 1422.6000 ;
	    RECT 611.4000 1421.4000 612.6000 1422.6000 ;
	    RECT 589.9500 1416.6000 590.8500 1421.4000 ;
	    RECT 606.7500 1419.6000 607.6500 1421.4000 ;
	    RECT 606.6000 1418.4000 607.8000 1419.6000 ;
	    RECT 589.8000 1415.4000 591.0000 1416.6000 ;
	    RECT 496.2000 1400.4000 497.4000 1401.6000 ;
	    RECT 498.6000 1389.3000 499.8000 1406.7001 ;
	    RECT 501.0000 1386.3000 502.2000 1406.7001 ;
	    RECT 503.4000 1386.3000 504.6000 1406.7001 ;
	    RECT 585.0000 1406.4000 586.2000 1407.6000 ;
	    RECT 505.8000 1397.4000 507.0000 1398.6000 ;
	    RECT 493.8000 1367.4000 495.0000 1368.6000 ;
	    RECT 493.9500 1365.6000 494.8500 1367.4000 ;
	    RECT 493.8000 1364.4000 495.0000 1365.6000 ;
	    RECT 496.2000 1361.4000 497.4000 1362.6000 ;
	    RECT 491.4000 1313.4000 492.6000 1314.6000 ;
	    RECT 479.4000 1301.4000 480.6000 1302.6000 ;
	    RECT 465.0000 1280.4000 466.2000 1281.6000 ;
	    RECT 465.1500 1266.6000 466.0500 1280.4000 ;
	    RECT 467.4000 1277.4000 468.6000 1278.6000 ;
	    RECT 465.0000 1265.4000 466.2000 1266.6000 ;
	    RECT 467.5500 1260.6000 468.4500 1277.4000 ;
	    RECT 472.2000 1274.4000 473.4000 1275.6000 ;
	    RECT 472.3500 1272.6000 473.2500 1274.4000 ;
	    RECT 472.2000 1271.4000 473.4000 1272.6000 ;
	    RECT 467.4000 1259.4000 468.6000 1260.6000 ;
	    RECT 479.5500 1248.6000 480.4500 1301.4000 ;
	    RECT 479.4000 1247.4000 480.6000 1248.6000 ;
	    RECT 479.4000 1241.4000 480.6000 1242.6000 ;
	    RECT 479.5500 1230.6000 480.4500 1241.4000 ;
	    RECT 479.4000 1229.4000 480.6000 1230.6000 ;
	    RECT 460.2000 1199.4000 461.4000 1200.6000 ;
	    RECT 477.0000 1199.4000 478.2000 1200.6000 ;
	    RECT 453.0000 1176.3000 454.2000 1196.7001 ;
	    RECT 455.4000 1176.3000 456.6000 1196.7001 ;
	    RECT 457.8000 1176.3000 459.0000 1196.7001 ;
	    RECT 460.2000 1176.3000 461.4000 1193.7001 ;
	    RECT 462.6000 1178.4000 463.8000 1179.6000 ;
	    RECT 462.7500 1170.6000 463.6500 1178.4000 ;
	    RECT 465.0000 1176.3000 466.2000 1193.7001 ;
	    RECT 467.4000 1181.4000 468.6000 1182.6000 ;
	    RECT 467.5500 1176.6000 468.4500 1181.4000 ;
	    RECT 467.4000 1175.4000 468.6000 1176.6000 ;
	    RECT 469.8000 1176.3000 471.0000 1193.7001 ;
	    RECT 472.2000 1176.3000 473.4000 1196.7001 ;
	    RECT 474.6000 1176.3000 475.8000 1196.7001 ;
	    RECT 477.1500 1194.6000 478.0500 1199.4000 ;
	    RECT 481.8000 1196.4000 483.0000 1197.6000 ;
	    RECT 477.0000 1193.4000 478.2000 1194.6000 ;
	    RECT 477.1500 1185.6000 478.0500 1193.4000 ;
	    RECT 481.9500 1188.6000 482.8500 1196.4000 ;
	    RECT 505.9500 1188.6000 506.8500 1397.4000 ;
	    RECT 510.6000 1394.4000 511.8000 1395.6000 ;
	    RECT 510.7500 1386.6000 511.6500 1394.4000 ;
	    RECT 510.6000 1385.4000 511.8000 1386.6000 ;
	    RECT 508.2000 1367.4000 509.4000 1368.6000 ;
	    RECT 508.3500 1359.6000 509.2500 1367.4000 ;
	    RECT 575.4000 1361.4000 576.6000 1362.6000 ;
	    RECT 508.2000 1358.4000 509.4000 1359.6000 ;
	    RECT 508.3500 1356.6000 509.2500 1358.4000 ;
	    RECT 508.2000 1355.4000 509.4000 1356.6000 ;
	    RECT 541.8000 1349.4000 543.0000 1350.6000 ;
	    RECT 527.4000 1326.3000 528.6000 1346.7001 ;
	    RECT 529.8000 1326.3000 531.0000 1346.7001 ;
	    RECT 532.2000 1326.3000 533.4000 1346.7001 ;
	    RECT 534.6000 1329.3000 535.8000 1346.7001 ;
	    RECT 537.0000 1343.4000 538.2000 1344.6000 ;
	    RECT 537.1500 1314.6000 538.0500 1343.4000 ;
	    RECT 539.4000 1329.3000 540.6000 1346.7001 ;
	    RECT 541.9500 1341.6000 542.8500 1349.4000 ;
	    RECT 541.8000 1340.4000 543.0000 1341.6000 ;
	    RECT 544.2000 1329.3000 545.4000 1346.7001 ;
	    RECT 546.6000 1326.3000 547.8000 1346.7001 ;
	    RECT 549.0000 1326.3000 550.2000 1346.7001 ;
	    RECT 551.4000 1337.4000 552.6000 1338.6000 ;
	    RECT 537.0000 1313.4000 538.2000 1314.6000 ;
	    RECT 539.4000 1280.4000 540.6000 1281.6000 ;
	    RECT 539.5500 1278.6000 540.4500 1280.4000 ;
	    RECT 532.2000 1277.4000 533.4000 1278.6000 ;
	    RECT 539.4000 1277.4000 540.6000 1278.6000 ;
	    RECT 532.3500 1260.6000 533.2500 1277.4000 ;
	    RECT 549.0000 1269.3000 550.2000 1286.7001 ;
	    RECT 551.5500 1266.6000 552.4500 1337.4000 ;
	    RECT 556.2000 1334.4000 557.4000 1335.6000 ;
	    RECT 556.3500 1326.6000 557.2500 1334.4000 ;
	    RECT 556.2000 1325.4000 557.4000 1326.6000 ;
	    RECT 558.6000 1277.4000 559.8000 1278.6000 ;
	    RECT 563.4000 1269.3000 564.6000 1286.7001 ;
	    RECT 565.8000 1280.4000 567.0000 1281.6000 ;
	    RECT 565.9500 1278.6000 566.8500 1280.4000 ;
	    RECT 565.8000 1277.4000 567.0000 1278.6000 ;
	    RECT 568.2000 1275.3000 569.4000 1283.7001 ;
	    RECT 551.4000 1265.4000 552.6000 1266.6000 ;
	    RECT 563.4000 1265.4000 564.6000 1266.6000 ;
	    RECT 532.2000 1259.4000 533.4000 1260.6000 ;
	    RECT 553.8000 1229.4000 555.0000 1230.6000 ;
	    RECT 525.0000 1205.4000 526.2000 1206.6000 ;
	    RECT 539.4000 1206.3000 540.6000 1226.7001 ;
	    RECT 541.8000 1206.3000 543.0000 1226.7001 ;
	    RECT 544.2000 1206.3000 545.4000 1226.7001 ;
	    RECT 546.6000 1209.3000 547.8000 1226.7001 ;
	    RECT 549.0000 1223.4000 550.2000 1224.6000 ;
	    RECT 481.8000 1187.4000 483.0000 1188.6000 ;
	    RECT 505.8000 1187.4000 507.0000 1188.6000 ;
	    RECT 522.6000 1187.4000 523.8000 1188.6000 ;
	    RECT 477.0000 1184.4000 478.2000 1185.6000 ;
	    RECT 522.7500 1182.6000 523.6500 1187.4000 ;
	    RECT 501.0000 1181.4000 502.2000 1182.6000 ;
	    RECT 522.6000 1181.4000 523.8000 1182.6000 ;
	    RECT 501.1500 1179.6000 502.0500 1181.4000 ;
	    RECT 501.0000 1178.4000 502.2000 1179.6000 ;
	    RECT 462.6000 1169.4000 463.8000 1170.6000 ;
	    RECT 486.6000 1169.4000 487.8000 1170.6000 ;
	    RECT 460.2000 1154.4000 461.4000 1155.6000 ;
	    RECT 460.3500 1152.6000 461.2500 1154.4000 ;
	    RECT 460.2000 1151.4000 461.4000 1152.6000 ;
	    RECT 455.4000 1146.4501 456.6000 1146.6000 ;
	    RECT 455.4000 1145.5500 458.8500 1146.4501 ;
	    RECT 477.0000 1146.3000 478.2000 1166.7001 ;
	    RECT 479.4000 1146.3000 480.6000 1166.7001 ;
	    RECT 481.8000 1146.3000 483.0000 1166.7001 ;
	    RECT 484.2000 1149.3000 485.4000 1166.7001 ;
	    RECT 486.7500 1164.6000 487.6500 1169.4000 ;
	    RECT 486.6000 1163.4000 487.8000 1164.6000 ;
	    RECT 455.4000 1145.4000 456.6000 1145.5500 ;
	    RECT 453.0000 1134.4501 454.2000 1134.6000 ;
	    RECT 450.7500 1133.5500 454.2000 1134.4501 ;
	    RECT 453.0000 1133.4000 454.2000 1133.5500 ;
	    RECT 426.6000 1124.4000 427.8000 1125.6000 ;
	    RECT 443.5500 1122.6000 444.4500 1133.4000 ;
	    RECT 453.1500 1122.6000 454.0500 1133.4000 ;
	    RECT 443.4000 1121.4000 444.6000 1122.6000 ;
	    RECT 453.0000 1121.4000 454.2000 1122.6000 ;
	    RECT 417.0000 1115.4000 418.2000 1116.6000 ;
	    RECT 445.8000 1115.4000 447.0000 1116.6000 ;
	    RECT 445.9500 1104.6000 446.8500 1115.4000 ;
	    RECT 445.8000 1103.4000 447.0000 1104.6000 ;
	    RECT 438.6000 1100.4000 439.8000 1101.6000 ;
	    RECT 419.4000 1094.4000 420.6000 1095.6000 ;
	    RECT 419.5500 1092.6000 420.4500 1094.4000 ;
	    RECT 419.4000 1091.4000 420.6000 1092.6000 ;
	    RECT 438.7500 1086.6000 439.6500 1100.4000 ;
	    RECT 438.6000 1085.4000 439.8000 1086.6000 ;
	    RECT 453.0000 1016.4000 454.2000 1017.6000 ;
	    RECT 453.1500 1008.6000 454.0500 1016.4000 ;
	    RECT 453.0000 1007.4000 454.2000 1008.6000 ;
	    RECT 457.9500 1005.6000 458.8500 1145.5500 ;
	    RECT 479.4000 1133.4000 480.6000 1134.6000 ;
	    RECT 477.0000 1127.4000 478.2000 1128.6000 ;
	    RECT 460.2000 1121.4000 461.4000 1122.6000 ;
	    RECT 460.3500 1020.6000 461.2500 1121.4000 ;
	    RECT 467.4000 1061.4000 468.6000 1062.6000 ;
	    RECT 460.2000 1019.4000 461.4000 1020.6000 ;
	    RECT 457.8000 1004.4000 459.0000 1005.6000 ;
	    RECT 419.4000 980.4000 420.6000 981.6000 ;
	    RECT 419.5500 960.6000 420.4500 980.4000 ;
	    RECT 453.0000 977.4000 454.2000 978.6000 ;
	    RECT 455.4000 977.4000 456.6000 978.6000 ;
	    RECT 424.2000 974.4000 425.4000 975.6000 ;
	    RECT 419.4000 959.4000 420.6000 960.6000 ;
	    RECT 417.0000 950.4000 418.2000 951.6000 ;
	    RECT 417.1500 942.6000 418.0500 950.4000 ;
	    RECT 424.3500 948.6000 425.2500 974.4000 ;
	    RECT 453.1500 972.6000 454.0500 977.4000 ;
	    RECT 453.0000 971.4000 454.2000 972.6000 ;
	    RECT 455.5500 960.6000 456.4500 977.4000 ;
	    RECT 431.4000 959.4000 432.6000 960.6000 ;
	    RECT 455.4000 959.4000 456.6000 960.6000 ;
	    RECT 424.2000 947.4000 425.4000 948.6000 ;
	    RECT 417.0000 941.4000 418.2000 942.6000 ;
	    RECT 417.0000 920.4000 418.2000 921.6000 ;
	    RECT 429.0000 920.4000 430.2000 921.6000 ;
	    RECT 417.1500 912.4500 418.0500 920.4000 ;
	    RECT 429.1500 918.6000 430.0500 920.4000 ;
	    RECT 424.2000 917.4000 425.4000 918.6000 ;
	    RECT 429.0000 917.4000 430.2000 918.6000 ;
	    RECT 426.6000 914.4000 427.8000 915.6000 ;
	    RECT 421.8000 912.4500 423.0000 912.6000 ;
	    RECT 417.1500 911.5500 423.0000 912.4500 ;
	    RECT 421.8000 911.4000 423.0000 911.5500 ;
	    RECT 417.0000 905.4000 418.2000 906.6000 ;
	    RECT 407.4000 881.4000 408.6000 882.6000 ;
	    RECT 412.2000 881.4000 413.4000 882.6000 ;
	    RECT 373.8000 869.4000 375.0000 870.6000 ;
	    RECT 373.8000 857.4000 375.0000 858.6000 ;
	    RECT 373.9500 846.6000 374.8500 857.4000 ;
	    RECT 373.8000 845.4000 375.0000 846.6000 ;
	    RECT 376.2000 846.3000 377.4000 866.7000 ;
	    RECT 378.6000 846.3000 379.8000 866.7000 ;
	    RECT 381.0000 849.3000 382.2000 866.7000 ;
	    RECT 383.4000 860.4000 384.6000 861.6000 ;
	    RECT 383.5500 852.6000 384.4500 860.4000 ;
	    RECT 383.4000 851.4000 384.6000 852.6000 ;
	    RECT 385.8000 849.3000 387.0000 866.7000 ;
	    RECT 388.2000 863.4000 389.4000 864.6000 ;
	    RECT 390.6000 849.3000 391.8000 866.7000 ;
	    RECT 383.4000 845.4000 384.6000 846.6000 ;
	    RECT 393.0000 846.3000 394.2000 866.7000 ;
	    RECT 395.4000 846.3000 396.6000 866.7000 ;
	    RECT 397.8000 846.3000 399.0000 866.7000 ;
	    RECT 371.5500 830.5500 374.8500 831.4500 ;
	    RECT 366.6000 827.4000 367.8000 828.6000 ;
	    RECT 369.0000 809.4000 370.2000 810.6000 ;
	    RECT 369.1500 801.6000 370.0500 809.4000 ;
	    RECT 369.0000 800.4000 370.2000 801.6000 ;
	    RECT 366.6000 779.4000 367.8000 780.6000 ;
	    RECT 366.7500 708.6000 367.6500 779.4000 ;
	    RECT 369.0000 776.4000 370.2000 777.6000 ;
	    RECT 369.1500 768.6000 370.0500 776.4000 ;
	    RECT 369.0000 767.4000 370.2000 768.6000 ;
	    RECT 373.9500 765.6000 374.8500 830.5500 ;
	    RECT 381.0000 821.4000 382.2000 822.6000 ;
	    RECT 381.1500 798.6000 382.0500 821.4000 ;
	    RECT 383.5500 804.6000 384.4500 845.4000 ;
	    RECT 390.6000 839.4000 391.8000 840.6000 ;
	    RECT 390.7500 822.6000 391.6500 839.4000 ;
	    RECT 407.5500 828.6000 408.4500 881.4000 ;
	    RECT 412.2000 851.4000 413.4000 852.6000 ;
	    RECT 412.3500 846.6000 413.2500 851.4000 ;
	    RECT 412.2000 845.4000 413.4000 846.6000 ;
	    RECT 400.2000 827.4000 401.4000 828.6000 ;
	    RECT 405.0000 827.4000 406.2000 828.6000 ;
	    RECT 407.4000 827.4000 408.6000 828.6000 ;
	    RECT 390.6000 821.4000 391.8000 822.6000 ;
	    RECT 383.4000 803.4000 384.6000 804.6000 ;
	    RECT 385.8000 800.4000 387.0000 801.6000 ;
	    RECT 393.0000 800.4000 394.2000 801.6000 ;
	    RECT 381.0000 797.4000 382.2000 798.6000 ;
	    RECT 383.4000 791.4000 384.6000 792.6000 ;
	    RECT 373.8000 764.4000 375.0000 765.6000 ;
	    RECT 371.4000 725.4000 372.6000 726.6000 ;
	    RECT 366.6000 707.4000 367.8000 708.6000 ;
	    RECT 369.0000 707.4000 370.2000 708.6000 ;
	    RECT 364.2000 674.4000 365.4000 675.6000 ;
	    RECT 359.4000 647.4000 360.6000 648.6000 ;
	    RECT 359.5500 621.6000 360.4500 647.4000 ;
	    RECT 361.8000 641.4000 363.0000 642.6000 ;
	    RECT 357.0000 620.4000 358.2000 621.6000 ;
	    RECT 359.4000 620.4000 360.6000 621.6000 ;
	    RECT 357.1500 612.6000 358.0500 620.4000 ;
	    RECT 361.9500 618.4500 362.8500 641.4000 ;
	    RECT 366.6000 620.4000 367.8000 621.6000 ;
	    RECT 364.2000 618.4500 365.4000 618.6000 ;
	    RECT 361.9500 617.5500 365.4000 618.4500 ;
	    RECT 364.2000 617.4000 365.4000 617.5500 ;
	    RECT 359.4000 614.4000 360.6000 615.6000 ;
	    RECT 357.0000 611.4000 358.2000 612.6000 ;
	    RECT 359.5500 600.6000 360.4500 614.4000 ;
	    RECT 359.4000 599.4000 360.6000 600.6000 ;
	    RECT 364.2000 600.4500 365.4000 600.6000 ;
	    RECT 366.7500 600.4500 367.6500 620.4000 ;
	    RECT 364.2000 599.5500 367.6500 600.4500 ;
	    RECT 364.2000 599.4000 365.4000 599.5500 ;
	    RECT 359.4000 587.4000 360.6000 588.6000 ;
	    RECT 359.5500 582.6000 360.4500 587.4000 ;
	    RECT 359.4000 581.4000 360.6000 582.6000 ;
	    RECT 361.8000 578.4000 363.0000 579.6000 ;
	    RECT 361.9500 576.6000 362.8500 578.4000 ;
	    RECT 361.8000 575.4000 363.0000 576.6000 ;
	    RECT 354.6000 560.4000 355.8000 561.6000 ;
	    RECT 357.0000 560.4000 358.2000 561.6000 ;
	    RECT 354.6000 557.4000 355.8000 558.6000 ;
	    RECT 352.2000 545.4000 353.4000 546.6000 ;
	    RECT 354.7500 540.6000 355.6500 557.4000 ;
	    RECT 357.1500 552.6000 358.0500 560.4000 ;
	    RECT 366.6000 557.4000 367.8000 558.6000 ;
	    RECT 357.0000 551.4000 358.2000 552.6000 ;
	    RECT 354.6000 539.4000 355.8000 540.6000 ;
	    RECT 349.8000 527.4000 351.0000 528.6000 ;
	    RECT 349.8000 521.4000 351.0000 522.6000 ;
	    RECT 349.9500 516.6000 350.8500 521.4000 ;
	    RECT 349.8000 515.4000 351.0000 516.6000 ;
	    RECT 352.2000 516.3000 353.4000 533.7000 ;
	    RECT 354.6000 518.4000 355.8000 519.6000 ;
	    RECT 354.7500 507.6000 355.6500 518.4000 ;
	    RECT 357.0000 516.3000 358.2000 533.7000 ;
	    RECT 359.4000 516.3000 360.6000 536.7000 ;
	    RECT 361.8000 516.3000 363.0000 536.7000 ;
	    RECT 364.2000 516.3000 365.4000 536.7000 ;
	    RECT 335.5500 506.5500 338.8500 507.4500 ;
	    RECT 333.0000 503.4000 334.2000 504.6000 ;
	    RECT 330.6000 500.4000 331.8000 501.6000 ;
	    RECT 330.6000 497.4000 331.8000 498.6000 ;
	    RECT 330.7500 480.6000 331.6500 497.4000 ;
	    RECT 333.1500 492.6000 334.0500 503.4000 ;
	    RECT 333.0000 491.4000 334.2000 492.6000 ;
	    RECT 330.6000 479.4000 331.8000 480.6000 ;
	    RECT 328.2000 461.4000 329.4000 462.6000 ;
	    RECT 328.3500 441.6000 329.2500 461.4000 ;
	    RECT 328.2000 440.4000 329.4000 441.6000 ;
	    RECT 328.2000 437.4000 329.4000 438.6000 ;
	    RECT 325.8000 431.4000 327.0000 432.6000 ;
	    RECT 323.4000 344.4000 324.6000 345.6000 ;
	    RECT 323.4000 305.4000 324.6000 306.6000 ;
	    RECT 309.0000 245.4000 310.2000 246.6000 ;
	    RECT 321.0000 245.4000 322.2000 246.6000 ;
	    RECT 306.6000 233.4000 307.8000 234.6000 ;
	    RECT 304.2000 194.4000 305.4000 195.6000 ;
	    RECT 304.3500 186.6000 305.2500 194.4000 ;
	    RECT 304.2000 185.4000 305.4000 186.6000 ;
	    RECT 292.2000 143.4000 293.4000 144.6000 ;
	    RECT 292.2000 128.4000 293.4000 129.6000 ;
	    RECT 287.4000 119.4000 288.6000 120.6000 ;
	    RECT 287.5500 114.6000 288.4500 119.4000 ;
	    RECT 287.4000 113.4000 288.6000 114.6000 ;
	    RECT 292.3500 108.6000 293.2500 128.4000 ;
	    RECT 285.0000 107.4000 286.2000 108.6000 ;
	    RECT 292.2000 107.4000 293.4000 108.6000 ;
	    RECT 282.6000 47.4000 283.8000 48.6000 ;
	    RECT 306.7500 36.6000 307.6500 233.4000 ;
	    RECT 309.1500 198.6000 310.0500 245.4000 ;
	    RECT 318.6000 221.4000 319.8000 222.6000 ;
	    RECT 309.0000 197.4000 310.2000 198.6000 ;
	    RECT 311.4000 186.3000 312.6000 206.7000 ;
	    RECT 313.8000 186.3000 315.0000 206.7000 ;
	    RECT 316.2000 189.3000 317.4000 206.7000 ;
	    RECT 318.7500 201.6000 319.6500 221.4000 ;
	    RECT 318.6000 200.4000 319.8000 201.6000 ;
	    RECT 321.0000 189.3000 322.2000 206.7000 ;
	    RECT 323.5500 204.6000 324.4500 305.4000 ;
	    RECT 325.9500 294.6000 326.8500 431.4000 ;
	    RECT 328.3500 402.6000 329.2500 437.4000 ;
	    RECT 330.6000 419.4000 331.8000 420.6000 ;
	    RECT 328.2000 401.4000 329.4000 402.6000 ;
	    RECT 325.8000 293.4000 327.0000 294.6000 ;
	    RECT 330.7500 264.6000 331.6500 419.4000 ;
	    RECT 333.1500 342.6000 334.0500 491.4000 ;
	    RECT 335.5500 468.6000 336.4500 506.5500 ;
	    RECT 354.6000 506.4000 355.8000 507.6000 ;
	    RECT 337.8000 503.4000 339.0000 504.6000 ;
	    RECT 335.4000 467.4000 336.6000 468.6000 ;
	    RECT 335.4000 461.4000 336.6000 462.6000 ;
	    RECT 333.0000 341.4000 334.2000 342.6000 ;
	    RECT 330.6000 263.4000 331.8000 264.6000 ;
	    RECT 333.0000 263.4000 334.2000 264.6000 ;
	    RECT 333.1500 255.6000 334.0500 263.4000 ;
	    RECT 333.0000 254.4000 334.2000 255.6000 ;
	    RECT 333.1500 216.6000 334.0500 254.4000 ;
	    RECT 335.5500 222.6000 336.4500 461.4000 ;
	    RECT 337.9500 390.6000 338.8500 503.4000 ;
	    RECT 345.0000 500.4000 346.2000 501.6000 ;
	    RECT 342.6000 485.4000 343.8000 486.6000 ;
	    RECT 340.2000 479.4000 341.4000 480.6000 ;
	    RECT 340.3500 468.6000 341.2500 479.4000 ;
	    RECT 340.2000 467.4000 341.4000 468.6000 ;
	    RECT 342.7500 465.6000 343.6500 485.4000 ;
	    RECT 342.6000 464.4000 343.8000 465.6000 ;
	    RECT 345.1500 441.6000 346.0500 500.4000 ;
	    RECT 347.4000 497.4000 348.6000 498.6000 ;
	    RECT 347.5500 495.6000 348.4500 497.4000 ;
	    RECT 347.4000 494.4000 348.6000 495.6000 ;
	    RECT 359.4000 494.4000 360.6000 495.6000 ;
	    RECT 359.5500 468.6000 360.4500 494.4000 ;
	    RECT 366.7500 474.6000 367.6500 557.4000 ;
	    RECT 366.6000 473.4000 367.8000 474.6000 ;
	    RECT 359.4000 467.4000 360.6000 468.6000 ;
	    RECT 349.8000 461.4000 351.0000 462.6000 ;
	    RECT 352.2000 461.4000 353.4000 462.6000 ;
	    RECT 349.9500 444.6000 350.8500 461.4000 ;
	    RECT 352.3500 444.6000 353.2500 461.4000 ;
	    RECT 349.8000 443.4000 351.0000 444.6000 ;
	    RECT 352.2000 443.4000 353.4000 444.6000 ;
	    RECT 345.0000 440.4000 346.2000 441.6000 ;
	    RECT 337.8000 389.4000 339.0000 390.6000 ;
	    RECT 342.6000 380.4000 343.8000 381.6000 ;
	    RECT 342.7500 378.6000 343.6500 380.4000 ;
	    RECT 342.6000 377.4000 343.8000 378.6000 ;
	    RECT 342.6000 344.4000 343.8000 345.6000 ;
	    RECT 340.2000 263.4000 341.4000 264.6000 ;
	    RECT 340.3500 261.6000 341.2500 263.4000 ;
	    RECT 340.2000 260.4000 341.4000 261.6000 ;
	    RECT 335.4000 221.4000 336.6000 222.6000 ;
	    RECT 337.8000 221.4000 339.0000 222.6000 ;
	    RECT 333.0000 215.4000 334.2000 216.6000 ;
	    RECT 323.4000 203.4000 324.6000 204.6000 ;
	    RECT 323.5500 150.6000 324.4500 203.4000 ;
	    RECT 325.8000 189.3000 327.0000 206.7000 ;
	    RECT 328.2000 186.3000 329.4000 206.7000 ;
	    RECT 330.6000 186.3000 331.8000 206.7000 ;
	    RECT 333.0000 186.3000 334.2000 206.7000 ;
	    RECT 323.4000 149.4000 324.6000 150.6000 ;
	    RECT 335.4000 149.4000 336.6000 150.6000 ;
	    RECT 321.0000 137.4000 322.2000 138.6000 ;
	    RECT 309.0000 101.4000 310.2000 102.6000 ;
	    RECT 311.4000 101.4000 312.6000 102.6000 ;
	    RECT 318.6000 101.4000 319.8000 102.6000 ;
	    RECT 309.1500 54.6000 310.0500 101.4000 ;
	    RECT 311.5500 90.6000 312.4500 101.4000 ;
	    RECT 321.1500 99.6000 322.0500 137.4000 ;
	    RECT 333.0000 134.4000 334.2000 135.6000 ;
	    RECT 333.1500 126.6000 334.0500 134.4000 ;
	    RECT 333.0000 125.4000 334.2000 126.6000 ;
	    RECT 321.0000 98.4000 322.2000 99.6000 ;
	    RECT 311.4000 89.4000 312.6000 90.6000 ;
	    RECT 321.1500 72.6000 322.0500 98.4000 ;
	    RECT 311.4000 71.4000 312.6000 72.6000 ;
	    RECT 321.0000 71.4000 322.2000 72.6000 ;
	    RECT 325.8000 66.3000 327.0000 86.7000 ;
	    RECT 328.2000 66.3000 329.4000 86.7000 ;
	    RECT 330.6000 66.3000 331.8000 86.7000 ;
	    RECT 333.0000 69.3000 334.2000 86.7000 ;
	    RECT 335.5500 84.6000 336.4500 149.4000 ;
	    RECT 337.9500 138.6000 338.8500 221.4000 ;
	    RECT 342.7500 174.6000 343.6500 344.4000 ;
	    RECT 345.1500 306.6000 346.0500 440.4000 ;
	    RECT 349.8000 374.4000 351.0000 375.6000 ;
	    RECT 349.9500 366.6000 350.8500 374.4000 ;
	    RECT 352.3500 372.6000 353.2500 443.4000 ;
	    RECT 371.5500 399.6000 372.4500 725.4000 ;
	    RECT 373.9500 606.6000 374.8500 764.4000 ;
	    RECT 376.2000 756.3000 377.4000 776.7000 ;
	    RECT 378.6000 756.3000 379.8000 776.7000 ;
	    RECT 381.0000 756.3000 382.2000 773.7000 ;
	    RECT 383.5500 762.6000 384.4500 791.4000 ;
	    RECT 385.9500 786.6000 386.8500 800.4000 ;
	    RECT 388.2000 797.4000 389.4000 798.6000 ;
	    RECT 385.8000 785.4000 387.0000 786.6000 ;
	    RECT 383.4000 761.4000 384.6000 762.6000 ;
	    RECT 385.8000 756.3000 387.0000 773.7000 ;
	    RECT 388.3500 759.6000 389.2500 797.4000 ;
	    RECT 393.1500 792.6000 394.0500 800.4000 ;
	    RECT 393.0000 791.4000 394.2000 792.6000 ;
	    RECT 388.2000 758.4000 389.4000 759.6000 ;
	    RECT 390.6000 756.3000 391.8000 773.7000 ;
	    RECT 393.0000 756.3000 394.2000 776.7000 ;
	    RECT 395.4000 756.3000 396.6000 776.7000 ;
	    RECT 397.8000 756.3000 399.0000 776.7000 ;
	    RECT 381.0000 671.4000 382.2000 672.6000 ;
	    RECT 373.8000 605.4000 375.0000 606.6000 ;
	    RECT 381.1500 582.6000 382.0500 671.4000 ;
	    RECT 400.3500 630.6000 401.2500 827.4000 ;
	    RECT 402.6000 824.4000 403.8000 825.6000 ;
	    RECT 400.2000 629.4000 401.4000 630.6000 ;
	    RECT 390.6000 620.4000 391.8000 621.6000 ;
	    RECT 388.2000 617.4000 389.4000 618.6000 ;
	    RECT 385.8000 614.4000 387.0000 615.6000 ;
	    RECT 385.9500 612.6000 386.8500 614.4000 ;
	    RECT 385.8000 611.4000 387.0000 612.6000 ;
	    RECT 383.4000 599.4000 384.6000 600.6000 ;
	    RECT 381.0000 581.4000 382.2000 582.6000 ;
	    RECT 378.6000 530.4000 379.8000 531.6000 ;
	    RECT 378.7500 492.6000 379.6500 530.4000 ;
	    RECT 373.8000 491.4000 375.0000 492.6000 ;
	    RECT 378.6000 491.4000 379.8000 492.6000 ;
	    RECT 373.9500 459.6000 374.8500 491.4000 ;
	    RECT 383.5500 465.6000 384.4500 599.4000 ;
	    RECT 385.8000 581.4000 387.0000 582.6000 ;
	    RECT 390.7500 558.6000 391.6500 620.4000 ;
	    RECT 393.0000 596.4000 394.2000 597.6000 ;
	    RECT 393.1500 588.6000 394.0500 596.4000 ;
	    RECT 402.7500 594.6000 403.6500 824.4000 ;
	    RECT 405.1500 726.6000 406.0500 827.4000 ;
	    RECT 407.4000 821.4000 408.6000 822.6000 ;
	    RECT 412.2000 821.4000 413.4000 822.6000 ;
	    RECT 407.5500 810.6000 408.4500 821.4000 ;
	    RECT 407.4000 809.4000 408.6000 810.6000 ;
	    RECT 412.3500 801.6000 413.2500 821.4000 ;
	    RECT 412.2000 800.4000 413.4000 801.6000 ;
	    RECT 412.3500 786.6000 413.2500 800.4000 ;
	    RECT 412.2000 785.4000 413.4000 786.6000 ;
	    RECT 412.2000 773.4000 413.4000 774.6000 ;
	    RECT 412.3500 771.6000 413.2500 773.4000 ;
	    RECT 412.2000 770.4000 413.4000 771.6000 ;
	    RECT 405.0000 725.4000 406.2000 726.6000 ;
	    RECT 412.2000 707.4000 413.4000 708.6000 ;
	    RECT 412.3500 705.6000 413.2500 707.4000 ;
	    RECT 412.2000 704.4000 413.4000 705.6000 ;
	    RECT 414.6000 704.4000 415.8000 705.6000 ;
	    RECT 414.7500 702.6000 415.6500 704.4000 ;
	    RECT 405.0000 701.4000 406.2000 702.6000 ;
	    RECT 412.2000 701.4000 413.4000 702.6000 ;
	    RECT 414.6000 701.4000 415.8000 702.6000 ;
	    RECT 405.1500 660.6000 406.0500 701.4000 ;
	    RECT 412.3500 660.6000 413.2500 701.4000 ;
	    RECT 405.0000 659.4000 406.2000 660.6000 ;
	    RECT 412.2000 659.4000 413.4000 660.6000 ;
	    RECT 417.1500 618.6000 418.0500 905.4000 ;
	    RECT 426.7500 861.6000 427.6500 914.4000 ;
	    RECT 431.5500 864.6000 432.4500 959.4000 ;
	    RECT 433.8000 953.4000 435.0000 954.6000 ;
	    RECT 433.9500 948.6000 434.8500 953.4000 ;
	    RECT 433.8000 947.4000 435.0000 948.6000 ;
	    RECT 453.0000 947.4000 454.2000 948.6000 ;
	    RECT 453.1500 945.6000 454.0500 947.4000 ;
	    RECT 453.0000 944.4000 454.2000 945.6000 ;
	    RECT 453.1500 924.6000 454.0500 944.4000 ;
	    RECT 455.5500 942.6000 456.4500 959.4000 ;
	    RECT 455.4000 941.4000 456.6000 942.6000 ;
	    RECT 453.0000 923.4000 454.2000 924.6000 ;
	    RECT 457.9500 921.4500 458.8500 1004.4000 ;
	    RECT 460.2000 996.3000 461.4000 1016.7000 ;
	    RECT 462.6000 996.3000 463.8000 1016.7000 ;
	    RECT 465.0000 996.3000 466.2000 1013.7000 ;
	    RECT 467.5500 1002.6000 468.4500 1061.4000 ;
	    RECT 472.2000 1049.4000 473.4000 1050.6000 ;
	    RECT 467.4000 1001.4000 468.6000 1002.6000 ;
	    RECT 469.8000 996.3000 471.0000 1013.7000 ;
	    RECT 472.3500 999.6000 473.2500 1049.4000 ;
	    RECT 477.1500 1044.6000 478.0500 1127.4000 ;
	    RECT 479.5500 1122.6000 480.4500 1133.4000 ;
	    RECT 479.4000 1121.4000 480.6000 1122.6000 ;
	    RECT 486.7500 1050.6000 487.6500 1163.4000 ;
	    RECT 489.0000 1149.3000 490.2000 1166.7001 ;
	    RECT 491.4000 1160.4000 492.6000 1161.6000 ;
	    RECT 491.5500 1152.6000 492.4500 1160.4000 ;
	    RECT 491.4000 1151.4000 492.6000 1152.6000 ;
	    RECT 493.8000 1149.3000 495.0000 1166.7001 ;
	    RECT 496.2000 1146.3000 497.4000 1166.7001 ;
	    RECT 498.6000 1146.3000 499.8000 1166.7001 ;
	    RECT 501.0000 1157.4000 502.2000 1158.6000 ;
	    RECT 501.1500 1140.6000 502.0500 1157.4000 ;
	    RECT 505.8000 1154.4000 507.0000 1155.6000 ;
	    RECT 505.9500 1146.6000 506.8500 1154.4000 ;
	    RECT 505.8000 1145.4000 507.0000 1146.6000 ;
	    RECT 501.0000 1139.4000 502.2000 1140.6000 ;
	    RECT 501.0000 1127.4000 502.2000 1128.6000 ;
	    RECT 508.2000 1127.4000 509.4000 1128.6000 ;
	    RECT 501.1500 1125.6000 502.0500 1127.4000 ;
	    RECT 501.0000 1124.4000 502.2000 1125.6000 ;
	    RECT 503.4000 1124.4000 504.6000 1125.6000 ;
	    RECT 503.5500 1101.6000 504.4500 1124.4000 ;
	    RECT 503.4000 1100.4000 504.6000 1101.6000 ;
	    RECT 498.6000 1091.4000 499.8000 1092.6000 ;
	    RECT 486.6000 1049.4000 487.8000 1050.6000 ;
	    RECT 477.0000 1043.4000 478.2000 1044.6000 ;
	    RECT 496.2000 1043.4000 497.4000 1044.6000 ;
	    RECT 486.6000 1031.4000 487.8000 1032.6000 ;
	    RECT 472.2000 998.4000 473.4000 999.6000 ;
	    RECT 465.0000 986.4000 466.2000 987.6000 ;
	    RECT 460.2000 974.4000 461.4000 975.6000 ;
	    RECT 460.3500 942.6000 461.2500 974.4000 ;
	    RECT 460.2000 941.4000 461.4000 942.6000 ;
	    RECT 465.1500 924.6000 466.0500 986.4000 ;
	    RECT 465.0000 923.4000 466.2000 924.6000 ;
	    RECT 455.5500 920.5500 458.8500 921.4500 ;
	    RECT 450.6000 890.4000 451.8000 891.6000 ;
	    RECT 450.7500 864.6000 451.6500 890.4000 ;
	    RECT 431.4000 863.4000 432.6000 864.6000 ;
	    RECT 450.6000 863.4000 451.8000 864.6000 ;
	    RECT 426.6000 860.4000 427.8000 861.6000 ;
	    RECT 429.0000 860.4000 430.2000 861.6000 ;
	    RECT 429.1500 804.6000 430.0500 860.4000 ;
	    RECT 431.4000 821.4000 432.6000 822.6000 ;
	    RECT 431.5500 810.6000 432.4500 821.4000 ;
	    RECT 431.4000 809.4000 432.6000 810.6000 ;
	    RECT 424.2000 803.4000 425.4000 804.6000 ;
	    RECT 429.0000 803.4000 430.2000 804.6000 ;
	    RECT 419.4000 800.4000 420.6000 801.6000 ;
	    RECT 419.5500 741.6000 420.4500 800.4000 ;
	    RECT 419.4000 740.4000 420.6000 741.6000 ;
	    RECT 424.3500 738.6000 425.2500 803.4000 ;
	    RECT 429.1500 795.6000 430.0500 803.4000 ;
	    RECT 429.0000 794.4000 430.2000 795.6000 ;
	    RECT 431.4000 767.4000 432.6000 768.6000 ;
	    RECT 431.5500 750.6000 432.4500 767.4000 ;
	    RECT 445.8000 761.4000 447.0000 762.6000 ;
	    RECT 431.4000 749.4000 432.6000 750.6000 ;
	    RECT 445.9500 744.6000 446.8500 761.4000 ;
	    RECT 445.8000 743.4000 447.0000 744.6000 ;
	    RECT 424.2000 737.4000 425.4000 738.6000 ;
	    RECT 419.4000 707.4000 420.6000 708.6000 ;
	    RECT 419.4000 701.4000 420.6000 702.6000 ;
	    RECT 421.8000 701.4000 423.0000 702.6000 ;
	    RECT 419.5500 696.6000 420.4500 701.4000 ;
	    RECT 419.4000 695.4000 420.6000 696.6000 ;
	    RECT 448.2000 695.4000 449.4000 696.6000 ;
	    RECT 421.8000 666.3000 423.0000 686.7000 ;
	    RECT 424.2000 666.3000 425.4000 686.7000 ;
	    RECT 426.6000 666.3000 427.8000 686.7000 ;
	    RECT 429.0000 669.3000 430.2000 686.7000 ;
	    RECT 431.4000 683.4000 432.6000 684.6000 ;
	    RECT 431.5500 672.6000 432.4500 683.4000 ;
	    RECT 431.4000 671.4000 432.6000 672.6000 ;
	    RECT 433.8000 669.3000 435.0000 686.7000 ;
	    RECT 436.2000 680.4000 437.4000 681.6000 ;
	    RECT 424.2000 656.4000 425.4000 657.6000 ;
	    RECT 419.4000 653.4000 420.6000 654.6000 ;
	    RECT 417.0000 617.4000 418.2000 618.6000 ;
	    RECT 402.6000 593.4000 403.8000 594.6000 ;
	    RECT 419.5500 588.6000 420.4500 653.4000 ;
	    RECT 424.3500 621.6000 425.2500 656.4000 ;
	    RECT 436.3500 648.6000 437.2500 680.4000 ;
	    RECT 438.6000 669.3000 439.8000 686.7000 ;
	    RECT 441.0000 666.3000 442.2000 686.7000 ;
	    RECT 443.4000 666.3000 444.6000 686.7000 ;
	    RECT 448.3500 684.6000 449.2500 695.4000 ;
	    RECT 448.2000 683.4000 449.4000 684.6000 ;
	    RECT 445.8000 677.4000 447.0000 678.6000 ;
	    RECT 445.9500 657.6000 446.8500 677.4000 ;
	    RECT 450.6000 674.4000 451.8000 675.6000 ;
	    RECT 450.7500 666.6000 451.6500 674.4000 ;
	    RECT 450.6000 665.4000 451.8000 666.6000 ;
	    RECT 450.6000 662.4000 451.8000 663.6000 ;
	    RECT 445.8000 656.4000 447.0000 657.6000 ;
	    RECT 450.7500 654.6000 451.6500 662.4000 ;
	    RECT 450.6000 653.4000 451.8000 654.6000 ;
	    RECT 436.2000 647.4000 437.4000 648.6000 ;
	    RECT 429.0000 644.4000 430.2000 645.6000 ;
	    RECT 426.6000 623.4000 427.8000 624.6000 ;
	    RECT 424.2000 620.4000 425.4000 621.6000 ;
	    RECT 393.0000 587.4000 394.2000 588.6000 ;
	    RECT 419.4000 587.4000 420.6000 588.6000 ;
	    RECT 421.8000 587.4000 423.0000 588.6000 ;
	    RECT 421.9500 585.6000 422.8500 587.4000 ;
	    RECT 405.0000 584.4000 406.2000 585.6000 ;
	    RECT 421.8000 584.4000 423.0000 585.6000 ;
	    RECT 390.6000 557.4000 391.8000 558.6000 ;
	    RECT 405.1500 486.6000 406.0500 584.4000 ;
	    RECT 409.8000 581.4000 411.0000 582.6000 ;
	    RECT 409.9500 570.6000 410.8500 581.4000 ;
	    RECT 426.7500 579.6000 427.6500 623.4000 ;
	    RECT 429.1500 615.6000 430.0500 644.4000 ;
	    RECT 450.7500 642.6000 451.6500 653.4000 ;
	    RECT 431.4000 641.4000 432.6000 642.6000 ;
	    RECT 450.6000 641.4000 451.8000 642.6000 ;
	    RECT 431.5500 621.6000 432.4500 641.4000 ;
	    RECT 450.7500 621.6000 451.6500 641.4000 ;
	    RECT 431.4000 620.4000 432.6000 621.6000 ;
	    RECT 450.6000 620.4000 451.8000 621.6000 ;
	    RECT 445.8000 617.4000 447.0000 618.6000 ;
	    RECT 429.0000 614.4000 430.2000 615.6000 ;
	    RECT 426.6000 578.4000 427.8000 579.6000 ;
	    RECT 453.0000 578.4000 454.2000 579.6000 ;
	    RECT 426.7500 576.6000 427.6500 578.4000 ;
	    RECT 426.6000 575.4000 427.8000 576.6000 ;
	    RECT 409.8000 569.4000 411.0000 570.6000 ;
	    RECT 445.8000 509.4000 447.0000 510.6000 ;
	    RECT 445.9500 507.6000 446.8500 509.4000 ;
	    RECT 445.8000 506.4000 447.0000 507.6000 ;
	    RECT 450.6000 497.4000 451.8000 498.6000 ;
	    RECT 409.8000 491.4000 411.0000 492.6000 ;
	    RECT 405.0000 485.4000 406.2000 486.6000 ;
	    RECT 393.0000 467.4000 394.2000 468.6000 ;
	    RECT 400.2000 467.4000 401.4000 468.6000 ;
	    RECT 383.4000 464.4000 384.6000 465.6000 ;
	    RECT 393.1500 462.6000 394.0500 467.4000 ;
	    RECT 393.0000 461.4000 394.2000 462.6000 ;
	    RECT 395.4000 461.4000 396.6000 462.6000 ;
	    RECT 373.8000 458.4000 375.0000 459.6000 ;
	    RECT 378.6000 440.4000 379.8000 441.6000 ;
	    RECT 378.7500 420.6000 379.6500 440.4000 ;
	    RECT 378.6000 419.4000 379.8000 420.6000 ;
	    RECT 371.4000 398.4000 372.6000 399.6000 ;
	    RECT 393.0000 398.4000 394.2000 399.6000 ;
	    RECT 352.2000 371.4000 353.4000 372.6000 ;
	    RECT 349.8000 365.4000 351.0000 366.6000 ;
	    RECT 347.4000 359.4000 348.6000 360.6000 ;
	    RECT 347.5500 348.6000 348.4500 359.4000 ;
	    RECT 347.4000 347.4000 348.6000 348.6000 ;
	    RECT 383.4000 347.4000 384.6000 348.6000 ;
	    RECT 390.6000 347.4000 391.8000 348.6000 ;
	    RECT 390.7500 345.6000 391.6500 347.4000 ;
	    RECT 388.2000 344.4000 389.4000 345.6000 ;
	    RECT 390.6000 344.4000 391.8000 345.6000 ;
	    RECT 388.3500 342.6000 389.2500 344.4000 ;
	    RECT 381.0000 341.4000 382.2000 342.6000 ;
	    RECT 383.4000 341.4000 384.6000 342.6000 ;
	    RECT 388.2000 341.4000 389.4000 342.6000 ;
	    RECT 357.0000 338.4000 358.2000 339.6000 ;
	    RECT 357.1500 312.6000 358.0500 338.4000 ;
	    RECT 383.5500 330.6000 384.4500 341.4000 ;
	    RECT 383.4000 329.4000 384.6000 330.6000 ;
	    RECT 385.8000 314.4000 387.0000 315.6000 ;
	    RECT 357.0000 311.4000 358.2000 312.6000 ;
	    RECT 345.0000 305.4000 346.2000 306.6000 ;
	    RECT 364.2000 305.4000 365.4000 306.6000 ;
	    RECT 345.0000 296.4000 346.2000 297.6000 ;
	    RECT 345.1500 288.6000 346.0500 296.4000 ;
	    RECT 345.0000 287.4000 346.2000 288.6000 ;
	    RECT 349.8000 284.4000 351.0000 285.6000 ;
	    RECT 349.9500 246.6000 350.8500 284.4000 ;
	    RECT 352.2000 276.3000 353.4000 296.7000 ;
	    RECT 354.6000 276.3000 355.8000 296.7000 ;
	    RECT 357.0000 276.3000 358.2000 293.7000 ;
	    RECT 359.4000 293.4000 360.6000 294.6000 ;
	    RECT 359.5500 282.6000 360.4500 293.4000 ;
	    RECT 359.4000 281.4000 360.6000 282.6000 ;
	    RECT 361.8000 276.3000 363.0000 293.7000 ;
	    RECT 364.3500 279.6000 365.2500 305.4000 ;
	    RECT 364.2000 278.4000 365.4000 279.6000 ;
	    RECT 366.6000 276.3000 367.8000 293.7000 ;
	    RECT 369.0000 276.3000 370.2000 296.7000 ;
	    RECT 371.4000 276.3000 372.6000 296.7000 ;
	    RECT 373.8000 276.3000 375.0000 296.7000 ;
	    RECT 385.9500 264.6000 386.8500 314.4000 ;
	    RECT 393.1500 291.6000 394.0500 398.4000 ;
	    RECT 393.0000 290.4000 394.2000 291.6000 ;
	    RECT 395.5500 264.6000 396.4500 461.4000 ;
	    RECT 400.3500 420.6000 401.2500 467.4000 ;
	    RECT 402.6000 440.4000 403.8000 441.6000 ;
	    RECT 400.2000 419.4000 401.4000 420.6000 ;
	    RECT 402.7500 384.6000 403.6500 440.4000 ;
	    RECT 405.0000 434.4000 406.2000 435.6000 ;
	    RECT 405.1500 420.6000 406.0500 434.4000 ;
	    RECT 405.0000 419.4000 406.2000 420.6000 ;
	    RECT 402.6000 383.4000 403.8000 384.6000 ;
	    RECT 402.6000 380.4000 403.8000 381.6000 ;
	    RECT 385.8000 263.4000 387.0000 264.6000 ;
	    RECT 395.4000 263.4000 396.6000 264.6000 ;
	    RECT 376.2000 260.4000 377.4000 261.6000 ;
	    RECT 376.3500 258.6000 377.2500 260.4000 ;
	    RECT 366.6000 257.4000 367.8000 258.6000 ;
	    RECT 369.0000 257.4000 370.2000 258.6000 ;
	    RECT 376.2000 257.4000 377.4000 258.6000 ;
	    RECT 383.4000 257.4000 384.6000 258.6000 ;
	    RECT 366.7500 252.6000 367.6500 257.4000 ;
	    RECT 373.8000 254.4000 375.0000 255.6000 ;
	    RECT 373.9500 252.6000 374.8500 254.4000 ;
	    RECT 366.6000 251.4000 367.8000 252.6000 ;
	    RECT 373.8000 251.4000 375.0000 252.6000 ;
	    RECT 349.8000 245.4000 351.0000 246.6000 ;
	    RECT 383.5500 228.6000 384.4500 257.4000 ;
	    RECT 385.9500 231.6000 386.8500 263.4000 ;
	    RECT 385.8000 230.4000 387.0000 231.6000 ;
	    RECT 383.4000 227.4000 384.6000 228.6000 ;
	    RECT 347.4000 224.4000 348.6000 225.6000 ;
	    RECT 347.5500 192.6000 348.4500 224.4000 ;
	    RECT 364.2000 218.4000 365.4000 219.6000 ;
	    RECT 364.3500 210.6000 365.2500 218.4000 ;
	    RECT 376.2000 215.4000 377.4000 216.6000 ;
	    RECT 364.2000 209.4000 365.4000 210.6000 ;
	    RECT 364.3500 204.6000 365.2500 209.4000 ;
	    RECT 364.2000 203.4000 365.4000 204.6000 ;
	    RECT 347.4000 191.4000 348.6000 192.6000 ;
	    RECT 364.2000 179.4000 365.4000 180.6000 ;
	    RECT 342.6000 173.4000 343.8000 174.6000 ;
	    RECT 352.2000 149.4000 353.4000 150.6000 ;
	    RECT 337.8000 137.4000 339.0000 138.6000 ;
	    RECT 337.9500 96.6000 338.8500 137.4000 ;
	    RECT 340.2000 126.3000 341.4000 146.7000 ;
	    RECT 342.6000 126.3000 343.8000 146.7000 ;
	    RECT 345.0000 129.3000 346.2000 146.7000 ;
	    RECT 347.4000 143.4000 348.6000 144.6000 ;
	    RECT 347.5500 141.6000 348.4500 143.4000 ;
	    RECT 347.4000 140.4000 348.6000 141.6000 ;
	    RECT 349.8000 129.3000 351.0000 146.7000 ;
	    RECT 352.3500 144.6000 353.2500 149.4000 ;
	    RECT 352.2000 143.4000 353.4000 144.6000 ;
	    RECT 354.6000 129.3000 355.8000 146.7000 ;
	    RECT 347.4000 125.4000 348.6000 126.6000 ;
	    RECT 357.0000 126.3000 358.2000 146.7000 ;
	    RECT 359.4000 126.3000 360.6000 146.7000 ;
	    RECT 361.8000 126.3000 363.0000 146.7000 ;
	    RECT 347.5500 114.6000 348.4500 125.4000 ;
	    RECT 347.4000 113.4000 348.6000 114.6000 ;
	    RECT 337.8000 95.4000 339.0000 96.6000 ;
	    RECT 357.0000 95.4000 358.2000 96.6000 ;
	    RECT 340.2000 89.4000 341.4000 90.6000 ;
	    RECT 349.8000 89.4000 351.0000 90.6000 ;
	    RECT 335.4000 83.4000 336.6000 84.6000 ;
	    RECT 335.5500 60.6000 336.4500 83.4000 ;
	    RECT 337.8000 69.3000 339.0000 86.7000 ;
	    RECT 340.3500 81.6000 341.2500 89.4000 ;
	    RECT 340.2000 80.4000 341.4000 81.6000 ;
	    RECT 342.6000 69.3000 343.8000 86.7000 ;
	    RECT 345.0000 66.3000 346.2000 86.7000 ;
	    RECT 347.4000 66.3000 348.6000 86.7000 ;
	    RECT 349.9500 78.6000 350.8500 89.4000 ;
	    RECT 349.8000 77.4000 351.0000 78.6000 ;
	    RECT 354.6000 74.4000 355.8000 75.6000 ;
	    RECT 354.7500 66.6000 355.6500 74.4000 ;
	    RECT 354.6000 65.4000 355.8000 66.6000 ;
	    RECT 335.4000 59.4000 336.6000 60.6000 ;
	    RECT 349.8000 59.4000 351.0000 60.6000 ;
	    RECT 309.0000 53.4000 310.2000 54.6000 ;
	    RECT 306.6000 35.4000 307.8000 36.6000 ;
	    RECT 323.4000 36.3000 324.6000 56.7000 ;
	    RECT 325.8000 36.3000 327.0000 56.7000 ;
	    RECT 328.2000 36.3000 329.4000 56.7000 ;
	    RECT 330.6000 36.3000 331.8000 53.7000 ;
	    RECT 333.0000 41.4000 334.2000 42.6000 ;
	    RECT 333.1500 39.6000 334.0500 41.4000 ;
	    RECT 333.0000 38.4000 334.2000 39.6000 ;
	    RECT 335.4000 36.3000 336.6000 53.7000 ;
	    RECT 337.8000 53.4000 339.0000 54.6000 ;
	    RECT 337.9500 42.6000 338.8500 53.4000 ;
	    RECT 337.8000 41.4000 339.0000 42.6000 ;
	    RECT 337.8000 35.4000 339.0000 36.6000 ;
	    RECT 340.2000 36.3000 341.4000 53.7000 ;
	    RECT 342.6000 36.3000 343.8000 56.7000 ;
	    RECT 345.0000 36.3000 346.2000 56.7000 ;
	    RECT 347.4000 47.4000 348.6000 48.6000 ;
	    RECT 347.5500 45.6000 348.4500 47.4000 ;
	    RECT 347.4000 44.4000 348.6000 45.6000 ;
	    RECT 256.2000 11.4000 257.4000 12.6000 ;
	    RECT 169.8000 5.4000 171.0000 6.6000 ;
	    RECT 323.4000 6.3000 324.6000 26.7000 ;
	    RECT 325.8000 6.3000 327.0000 26.7000 ;
	    RECT 328.2000 6.3000 329.4000 26.7000 ;
	    RECT 330.6000 9.3000 331.8000 26.7000 ;
	    RECT 333.0000 23.4000 334.2000 24.6000 ;
	    RECT 335.4000 9.3000 336.6000 26.7000 ;
	    RECT 337.9500 21.6000 338.8500 35.4000 ;
	    RECT 347.4000 29.4000 348.6000 30.6000 ;
	    RECT 337.8000 20.4000 339.0000 21.6000 ;
	    RECT 340.2000 9.3000 341.4000 26.7000 ;
	    RECT 342.6000 6.3000 343.8000 26.7000 ;
	    RECT 345.0000 6.3000 346.2000 26.7000 ;
	    RECT 347.5500 18.6000 348.4500 29.4000 ;
	    RECT 349.9500 24.6000 350.8500 59.4000 ;
	    RECT 352.2000 56.4000 353.4000 57.6000 ;
	    RECT 352.3500 48.6000 353.2500 56.4000 ;
	    RECT 352.2000 47.4000 353.4000 48.6000 ;
	    RECT 357.1500 30.6000 358.0500 95.4000 ;
	    RECT 364.3500 90.6000 365.2500 179.4000 ;
	    RECT 376.3500 132.6000 377.2500 215.4000 ;
	    RECT 381.0000 209.4000 382.2000 210.6000 ;
	    RECT 397.8000 209.4000 399.0000 210.6000 ;
	    RECT 381.1500 204.6000 382.0500 209.4000 ;
	    RECT 397.9500 204.6000 398.8500 209.4000 ;
	    RECT 381.0000 203.4000 382.2000 204.6000 ;
	    RECT 397.8000 203.4000 399.0000 204.6000 ;
	    RECT 381.0000 200.4000 382.2000 201.6000 ;
	    RECT 395.4000 200.4000 396.6000 201.6000 ;
	    RECT 376.2000 131.4000 377.4000 132.6000 ;
	    RECT 381.1500 108.6000 382.0500 200.4000 ;
	    RECT 381.0000 107.4000 382.2000 108.6000 ;
	    RECT 364.2000 89.4000 365.4000 90.6000 ;
	    RECT 369.0000 59.4000 370.2000 60.6000 ;
	    RECT 369.1500 39.6000 370.0500 59.4000 ;
	    RECT 369.0000 38.4000 370.2000 39.6000 ;
	    RECT 357.0000 29.4000 358.2000 30.6000 ;
	    RECT 349.8000 23.4000 351.0000 24.6000 ;
	    RECT 347.4000 17.4000 348.6000 18.6000 ;
	    RECT 352.2000 14.4000 353.4000 15.6000 ;
	    RECT 352.3500 6.6000 353.2500 14.4000 ;
	    RECT 395.5500 12.6000 396.4500 200.4000 ;
	    RECT 402.7500 168.6000 403.6500 380.4000 ;
	    RECT 409.9500 342.6000 410.8500 491.4000 ;
	    RECT 431.4000 485.4000 432.6000 486.6000 ;
	    RECT 431.5500 468.6000 432.4500 485.4000 ;
	    RECT 426.6000 467.4000 427.8000 468.6000 ;
	    RECT 431.4000 467.4000 432.6000 468.6000 ;
	    RECT 426.7500 465.6000 427.6500 467.4000 ;
	    RECT 426.6000 464.4000 427.8000 465.6000 ;
	    RECT 450.7500 462.6000 451.6500 497.4000 ;
	    RECT 453.1500 462.6000 454.0500 578.4000 ;
	    RECT 455.5500 501.6000 456.4500 920.5500 ;
	    RECT 472.3500 900.6000 473.2500 998.4000 ;
	    RECT 474.6000 996.3000 475.8000 1013.7000 ;
	    RECT 477.0000 996.3000 478.2000 1016.7000 ;
	    RECT 479.4000 996.3000 480.6000 1016.7000 ;
	    RECT 481.8000 996.3000 483.0000 1016.7000 ;
	    RECT 486.7500 987.6000 487.6500 1031.4000 ;
	    RECT 491.4000 1019.4000 492.6000 1020.6000 ;
	    RECT 486.6000 986.4000 487.8000 987.6000 ;
	    RECT 479.4000 938.4000 480.6000 939.6000 ;
	    RECT 477.0000 920.4000 478.2000 921.6000 ;
	    RECT 472.2000 899.4000 473.4000 900.6000 ;
	    RECT 477.1500 861.6000 478.0500 920.4000 ;
	    RECT 477.0000 860.4000 478.2000 861.6000 ;
	    RECT 474.6000 851.4000 475.8000 852.6000 ;
	    RECT 474.7500 825.6000 475.6500 851.4000 ;
	    RECT 474.6000 824.4000 475.8000 825.6000 ;
	    RECT 460.2000 713.4000 461.4000 714.6000 ;
	    RECT 460.3500 699.6000 461.2500 713.4000 ;
	    RECT 479.5500 702.6000 480.4500 938.4000 ;
	    RECT 491.5500 924.6000 492.4500 1019.4000 ;
	    RECT 496.3500 1011.6000 497.2500 1043.4000 ;
	    RECT 496.2000 1010.4000 497.4000 1011.6000 ;
	    RECT 491.4000 923.4000 492.6000 924.6000 ;
	    RECT 491.5500 921.6000 492.4500 923.4000 ;
	    RECT 491.4000 920.4000 492.6000 921.6000 ;
	    RECT 498.7500 918.6000 499.6500 1091.4000 ;
	    RECT 517.8000 1067.4000 519.0000 1068.6000 ;
	    RECT 517.9500 1050.6000 518.8500 1067.4000 ;
	    RECT 525.1500 1062.6000 526.0500 1205.4000 ;
	    RECT 544.2000 1184.4000 545.4000 1185.6000 ;
	    RECT 527.4000 1181.4000 528.6000 1182.6000 ;
	    RECT 529.8000 1181.4000 531.0000 1182.6000 ;
	    RECT 527.5500 1164.6000 528.4500 1181.4000 ;
	    RECT 527.4000 1163.4000 528.6000 1164.6000 ;
	    RECT 544.3500 1161.6000 545.2500 1184.4000 ;
	    RECT 546.6000 1181.4000 547.8000 1182.6000 ;
	    RECT 546.7500 1179.6000 547.6500 1181.4000 ;
	    RECT 546.6000 1178.4000 547.8000 1179.6000 ;
	    RECT 544.2000 1160.4000 545.4000 1161.6000 ;
	    RECT 549.1500 1104.6000 550.0500 1223.4000 ;
	    RECT 551.4000 1209.3000 552.6000 1226.7001 ;
	    RECT 553.9500 1221.6000 554.8500 1229.4000 ;
	    RECT 553.8000 1220.4000 555.0000 1221.6000 ;
	    RECT 556.2000 1209.3000 557.4000 1226.7001 ;
	    RECT 558.6000 1206.3000 559.8000 1226.7001 ;
	    RECT 561.0000 1206.3000 562.2000 1226.7001 ;
	    RECT 563.5500 1218.6000 564.4500 1265.4000 ;
	    RECT 563.4000 1217.4000 564.6000 1218.6000 ;
	    RECT 563.5500 1206.6000 564.4500 1217.4000 ;
	    RECT 568.2000 1214.4000 569.4000 1215.6000 ;
	    RECT 568.3500 1206.6000 569.2500 1214.4000 ;
	    RECT 563.4000 1205.4000 564.6000 1206.6000 ;
	    RECT 568.2000 1205.4000 569.4000 1206.6000 ;
	    RECT 570.6000 1193.4000 571.8000 1194.6000 ;
	    RECT 551.4000 1184.4000 552.6000 1185.6000 ;
	    RECT 551.5500 1146.6000 552.4500 1184.4000 ;
	    RECT 563.4000 1181.4000 564.6000 1182.6000 ;
	    RECT 563.5500 1170.6000 564.4500 1181.4000 ;
	    RECT 563.4000 1169.4000 564.6000 1170.6000 ;
	    RECT 554.1000 1163.4000 555.3000 1163.7001 ;
	    RECT 554.1000 1162.5000 562.5000 1163.4000 ;
	    RECT 563.4000 1162.5000 564.6000 1163.7001 ;
	    RECT 554.1000 1155.3000 555.0000 1162.5000 ;
	    RECT 556.2000 1162.2001 557.4000 1162.5000 ;
	    RECT 561.3000 1162.2001 562.5000 1162.5000 ;
	    RECT 563.7000 1161.3000 564.6000 1162.5000 ;
	    RECT 556.2000 1160.4000 564.6000 1161.3000 ;
	    RECT 565.8000 1160.4000 567.0000 1161.6000 ;
	    RECT 556.2000 1158.3000 557.1000 1160.4000 ;
	    RECT 555.9000 1157.1000 557.1000 1158.3000 ;
	    RECT 563.7000 1155.3000 564.6000 1160.4000 ;
	    RECT 565.9500 1158.6000 566.8500 1160.4000 ;
	    RECT 565.8000 1157.4000 567.0000 1158.6000 ;
	    RECT 554.1000 1154.1000 555.3000 1155.3000 ;
	    RECT 563.4000 1154.1000 564.6000 1155.3000 ;
	    RECT 551.4000 1145.4000 552.6000 1146.6000 ;
	    RECT 541.8000 1103.4000 543.0000 1104.6000 ;
	    RECT 549.0000 1103.4000 550.2000 1104.6000 ;
	    RECT 525.0000 1061.4000 526.2000 1062.6000 ;
	    RECT 510.6000 1049.4000 511.8000 1050.6000 ;
	    RECT 517.8000 1049.4000 519.0000 1050.6000 ;
	    RECT 501.0000 1026.3000 502.2000 1046.7001 ;
	    RECT 503.4000 1026.3000 504.6000 1046.7001 ;
	    RECT 505.8000 1026.3000 507.0000 1046.7001 ;
	    RECT 508.2000 1029.3000 509.4000 1046.7001 ;
	    RECT 510.7500 1044.6000 511.6500 1049.4000 ;
	    RECT 510.6000 1043.4000 511.8000 1044.6000 ;
	    RECT 513.0000 1029.3000 514.2000 1046.7001 ;
	    RECT 515.4000 1040.4000 516.6000 1041.6000 ;
	    RECT 515.5500 1026.4501 516.4500 1040.4000 ;
	    RECT 517.8000 1029.3000 519.0000 1046.7001 ;
	    RECT 513.1500 1025.5500 516.4500 1026.4501 ;
	    RECT 520.2000 1026.3000 521.4000 1046.7001 ;
	    RECT 522.6000 1026.3000 523.8000 1046.7001 ;
	    RECT 525.1500 1038.6000 526.0500 1061.4000 ;
	    RECT 532.2000 1056.3000 533.4000 1076.7001 ;
	    RECT 534.6000 1056.3000 535.8000 1076.7001 ;
	    RECT 537.0000 1056.3000 538.2000 1076.7001 ;
	    RECT 539.4000 1056.3000 540.6000 1073.7001 ;
	    RECT 541.9500 1068.6000 542.8500 1103.4000 ;
	    RECT 546.6000 1085.4000 547.8000 1086.6000 ;
	    RECT 541.8000 1067.4000 543.0000 1068.6000 ;
	    RECT 541.9500 1059.6000 542.8500 1067.4000 ;
	    RECT 541.8000 1058.4000 543.0000 1059.6000 ;
	    RECT 544.2000 1056.3000 545.4000 1073.7001 ;
	    RECT 546.7500 1062.6000 547.6500 1085.4000 ;
	    RECT 546.6000 1061.4000 547.8000 1062.6000 ;
	    RECT 549.0000 1056.3000 550.2000 1073.7001 ;
	    RECT 551.4000 1056.3000 552.6000 1076.7001 ;
	    RECT 553.8000 1056.3000 555.0000 1076.7001 ;
	    RECT 561.0000 1076.4000 562.2000 1077.6000 ;
	    RECT 561.1500 1068.6000 562.0500 1076.4000 ;
	    RECT 561.0000 1067.4000 562.2000 1068.6000 ;
	    RECT 556.2000 1064.4000 557.4000 1065.6000 ;
	    RECT 556.3500 1062.6000 557.2500 1064.4000 ;
	    RECT 556.2000 1061.4000 557.4000 1062.6000 ;
	    RECT 525.0000 1037.4000 526.2000 1038.6000 ;
	    RECT 539.4000 1037.4000 540.6000 1038.6000 ;
	    RECT 510.6000 1013.4000 511.8000 1014.6000 ;
	    RECT 510.7500 999.6000 511.6500 1013.4000 ;
	    RECT 510.6000 998.4000 511.8000 999.6000 ;
	    RECT 508.2000 969.3000 509.4000 986.7000 ;
	    RECT 508.2000 965.4000 509.4000 966.6000 ;
	    RECT 498.6000 917.4000 499.8000 918.6000 ;
	    RECT 498.6000 899.4000 499.8000 900.6000 ;
	    RECT 496.2000 860.4000 497.4000 861.6000 ;
	    RECT 484.2000 854.4000 485.4000 855.6000 ;
	    RECT 484.3500 852.6000 485.2500 854.4000 ;
	    RECT 484.2000 851.4000 485.4000 852.6000 ;
	    RECT 496.3500 840.6000 497.2500 860.4000 ;
	    RECT 496.2000 839.4000 497.4000 840.6000 ;
	    RECT 498.7500 825.6000 499.6500 899.4000 ;
	    RECT 501.0000 863.4000 502.2000 864.6000 ;
	    RECT 501.1500 858.6000 502.0500 863.4000 ;
	    RECT 501.0000 857.4000 502.2000 858.6000 ;
	    RECT 498.6000 824.4000 499.8000 825.6000 ;
	    RECT 496.2000 821.4000 497.4000 822.6000 ;
	    RECT 496.3500 765.6000 497.2500 821.4000 ;
	    RECT 501.1500 810.4500 502.0500 857.4000 ;
	    RECT 508.3500 819.6000 509.2500 965.4000 ;
	    RECT 510.7500 939.6000 511.6500 998.4000 ;
	    RECT 510.6000 938.4000 511.8000 939.6000 ;
	    RECT 513.1500 921.6000 514.0500 1025.5500 ;
	    RECT 525.1500 1020.6000 526.0500 1037.4000 ;
	    RECT 529.8000 1034.4000 531.0000 1035.6000 ;
	    RECT 529.9500 1026.6000 530.8500 1034.4000 ;
	    RECT 529.8000 1025.4000 531.0000 1026.6000 ;
	    RECT 520.2000 1019.4000 521.4000 1020.6000 ;
	    RECT 525.0000 1019.4000 526.2000 1020.6000 ;
	    RECT 515.4000 1007.4000 516.6000 1008.6000 ;
	    RECT 517.8000 977.4000 519.0000 978.6000 ;
	    RECT 517.9500 972.6000 518.8500 977.4000 ;
	    RECT 517.8000 971.4000 519.0000 972.6000 ;
	    RECT 517.8000 923.4000 519.0000 924.6000 ;
	    RECT 517.9500 921.6000 518.8500 923.4000 ;
	    RECT 513.0000 920.4000 514.2000 921.6000 ;
	    RECT 517.8000 920.4000 519.0000 921.6000 ;
	    RECT 517.8000 917.4000 519.0000 918.6000 ;
	    RECT 517.9500 915.6000 518.8500 917.4000 ;
	    RECT 517.8000 914.4000 519.0000 915.6000 ;
	    RECT 517.8000 860.4000 519.0000 861.6000 ;
	    RECT 517.9500 846.6000 518.8500 860.4000 ;
	    RECT 517.8000 845.4000 519.0000 846.6000 ;
	    RECT 508.2000 818.4000 509.4000 819.6000 ;
	    RECT 498.7500 809.5500 502.0500 810.4500 ;
	    RECT 496.2000 764.4000 497.4000 765.6000 ;
	    RECT 493.8000 761.4000 495.0000 762.6000 ;
	    RECT 493.9500 726.4500 494.8500 761.4000 ;
	    RECT 496.2000 734.4000 497.4000 735.6000 ;
	    RECT 496.3500 726.6000 497.2500 734.4000 ;
	    RECT 496.2000 726.4500 497.4000 726.6000 ;
	    RECT 493.9500 725.5500 497.4000 726.4500 ;
	    RECT 496.2000 725.4000 497.4000 725.5500 ;
	    RECT 479.4000 701.4000 480.6000 702.6000 ;
	    RECT 460.2000 698.4000 461.4000 699.6000 ;
	    RECT 474.6000 623.4000 475.8000 624.6000 ;
	    RECT 491.4000 623.4000 492.6000 624.6000 ;
	    RECT 462.6000 620.4000 463.8000 621.6000 ;
	    RECT 465.0000 620.4000 466.2000 621.6000 ;
	    RECT 457.8000 587.4000 459.0000 588.6000 ;
	    RECT 462.7500 585.6000 463.6500 620.4000 ;
	    RECT 465.1500 618.6000 466.0500 620.4000 ;
	    RECT 465.0000 617.4000 466.2000 618.6000 ;
	    RECT 474.7500 606.6000 475.6500 623.4000 ;
	    RECT 498.7500 609.6000 499.6500 809.5500 ;
	    RECT 508.3500 750.6000 509.2500 818.4000 ;
	    RECT 520.3500 804.6000 521.2500 1019.4000 ;
	    RECT 532.2000 1001.4000 533.4000 1002.6000 ;
	    RECT 537.0000 1001.4000 538.2000 1002.6000 ;
	    RECT 522.6000 969.3000 523.8000 986.7000 ;
	    RECT 525.0000 983.4000 526.2000 984.6000 ;
	    RECT 525.1500 981.6000 526.0500 983.4000 ;
	    RECT 525.0000 980.4000 526.2000 981.6000 ;
	    RECT 527.4000 975.3000 528.6000 983.7000 ;
	    RECT 525.0000 959.4000 526.2000 960.6000 ;
	    RECT 532.3500 954.6000 533.2500 1001.4000 ;
	    RECT 537.1500 960.6000 538.0500 1001.4000 ;
	    RECT 539.5500 984.6000 540.4500 1037.4000 ;
	    RECT 561.0000 1025.4000 562.2000 1026.6000 ;
	    RECT 561.1500 1002.6000 562.0500 1025.4000 ;
	    RECT 568.2000 1013.4000 569.4000 1014.6000 ;
	    RECT 568.3500 1002.6000 569.2500 1013.4000 ;
	    RECT 561.0000 1001.4000 562.2000 1002.6000 ;
	    RECT 568.2000 1001.4000 569.4000 1002.6000 ;
	    RECT 539.4000 983.4000 540.6000 984.6000 ;
	    RECT 537.0000 959.4000 538.2000 960.6000 ;
	    RECT 532.2000 953.4000 533.4000 954.6000 ;
	    RECT 561.0000 935.4000 562.2000 936.6000 ;
	    RECT 534.6000 923.4000 535.8000 924.6000 ;
	    RECT 534.7500 921.6000 535.6500 923.4000 ;
	    RECT 534.6000 920.4000 535.8000 921.6000 ;
	    RECT 522.6000 917.4000 523.8000 918.6000 ;
	    RECT 541.8000 914.4000 543.0000 915.6000 ;
	    RECT 525.0000 864.4500 526.2000 864.6000 ;
	    RECT 522.7500 863.5500 526.2000 864.4500 ;
	    RECT 522.7500 819.6000 523.6500 863.5500 ;
	    RECT 525.0000 863.4000 526.2000 863.5500 ;
	    RECT 541.9500 828.6000 542.8500 914.4000 ;
	    RECT 556.2000 893.4000 557.4000 894.6000 ;
	    RECT 549.0000 863.4000 550.2000 864.6000 ;
	    RECT 549.1500 861.6000 550.0500 863.4000 ;
	    RECT 549.0000 860.4000 550.2000 861.6000 ;
	    RECT 551.4000 860.4000 552.6000 861.6000 ;
	    RECT 551.5500 858.4500 552.4500 860.4000 ;
	    RECT 556.3500 858.6000 557.2500 893.4000 ;
	    RECT 549.1500 857.5500 552.4500 858.4500 ;
	    RECT 541.8000 827.4000 543.0000 828.6000 ;
	    RECT 522.6000 818.4000 523.8000 819.6000 ;
	    RECT 520.2000 803.4000 521.4000 804.6000 ;
	    RECT 522.7500 792.6000 523.6500 818.4000 ;
	    RECT 522.6000 791.4000 523.8000 792.6000 ;
	    RECT 515.4000 773.4000 516.6000 774.6000 ;
	    RECT 508.2000 749.4000 509.4000 750.6000 ;
	    RECT 501.0000 737.4000 502.2000 738.6000 ;
	    RECT 501.1500 690.6000 502.0500 737.4000 ;
	    RECT 503.4000 726.3000 504.6000 746.7000 ;
	    RECT 505.8000 726.3000 507.0000 746.7000 ;
	    RECT 508.2000 729.3000 509.4000 746.7000 ;
	    RECT 510.6000 743.4000 511.8000 744.6000 ;
	    RECT 510.7500 741.6000 511.6500 743.4000 ;
	    RECT 510.6000 740.4000 511.8000 741.6000 ;
	    RECT 513.0000 729.3000 514.2000 746.7000 ;
	    RECT 515.5500 744.6000 516.4500 773.4000 ;
	    RECT 549.1500 762.6000 550.0500 857.5500 ;
	    RECT 556.2000 857.4000 557.4000 858.6000 ;
	    RECT 551.4000 854.4000 552.6000 855.6000 ;
	    RECT 561.1500 855.4500 562.0500 935.4000 ;
	    RECT 570.7500 930.6000 571.6500 1193.4000 ;
	    RECT 573.0000 1094.4000 574.2000 1095.6000 ;
	    RECT 573.1500 1086.6000 574.0500 1094.4000 ;
	    RECT 573.0000 1085.4000 574.2000 1086.6000 ;
	    RECT 573.0000 1067.4000 574.2000 1068.6000 ;
	    RECT 570.6000 929.4000 571.8000 930.6000 ;
	    RECT 565.8000 923.4000 567.0000 924.6000 ;
	    RECT 565.9500 915.6000 566.8500 923.4000 ;
	    RECT 565.8000 914.4000 567.0000 915.6000 ;
	    RECT 573.1500 906.6000 574.0500 1067.4000 ;
	    RECT 575.5500 936.6000 576.4500 1361.4000 ;
	    RECT 580.2000 1310.4000 581.4000 1311.6000 ;
	    RECT 580.3500 1284.6000 581.2500 1310.4000 ;
	    RECT 580.2000 1283.4000 581.4000 1284.6000 ;
	    RECT 577.8000 1187.4000 579.0000 1188.6000 ;
	    RECT 577.9500 1098.6000 578.8500 1187.4000 ;
	    RECT 580.3500 1182.6000 581.2500 1283.4000 ;
	    RECT 597.0000 1235.4000 598.2000 1236.6000 ;
	    RECT 597.1500 1221.6000 598.0500 1235.4000 ;
	    RECT 597.0000 1220.4000 598.2000 1221.6000 ;
	    RECT 604.2000 1220.4000 605.4000 1221.6000 ;
	    RECT 601.8000 1217.4000 603.0000 1218.6000 ;
	    RECT 597.0000 1214.4000 598.2000 1215.6000 ;
	    RECT 580.2000 1181.4000 581.4000 1182.6000 ;
	    RECT 580.3500 1161.6000 581.2500 1181.4000 ;
	    RECT 585.0000 1163.4000 586.2000 1164.6000 ;
	    RECT 580.2000 1160.4000 581.4000 1161.6000 ;
	    RECT 585.1500 1158.6000 586.0500 1163.4000 ;
	    RECT 589.8000 1160.4000 591.0000 1161.6000 ;
	    RECT 589.9500 1158.6000 590.8500 1160.4000 ;
	    RECT 582.6000 1157.4000 583.8000 1158.6000 ;
	    RECT 585.0000 1157.4000 586.2000 1158.6000 ;
	    RECT 589.8000 1157.4000 591.0000 1158.6000 ;
	    RECT 582.7500 1152.6000 583.6500 1157.4000 ;
	    RECT 589.8000 1154.4000 591.0000 1155.6000 ;
	    RECT 582.6000 1151.4000 583.8000 1152.6000 ;
	    RECT 589.9500 1146.6000 590.8500 1154.4000 ;
	    RECT 589.8000 1145.4000 591.0000 1146.6000 ;
	    RECT 587.4000 1121.4000 588.6000 1122.6000 ;
	    RECT 577.8000 1097.4000 579.0000 1098.6000 ;
	    RECT 580.2000 1086.3000 581.4000 1106.7001 ;
	    RECT 582.6000 1086.3000 583.8000 1106.7001 ;
	    RECT 585.0000 1089.3000 586.2000 1106.7001 ;
	    RECT 587.5500 1101.6000 588.4500 1121.4000 ;
	    RECT 597.1500 1110.6000 598.0500 1214.4000 ;
	    RECT 601.9500 1182.6000 602.8500 1217.4000 ;
	    RECT 604.3500 1197.6000 605.2500 1220.4000 ;
	    RECT 604.2000 1196.4000 605.4000 1197.6000 ;
	    RECT 601.8000 1181.4000 603.0000 1182.6000 ;
	    RECT 597.0000 1109.4000 598.2000 1110.6000 ;
	    RECT 587.4000 1100.4000 588.6000 1101.6000 ;
	    RECT 589.8000 1089.3000 591.0000 1106.7001 ;
	    RECT 592.2000 1103.4000 593.4000 1104.6000 ;
	    RECT 592.2000 1097.4000 593.4000 1098.6000 ;
	    RECT 592.3500 1065.6000 593.2500 1097.4000 ;
	    RECT 594.6000 1089.3000 595.8000 1106.7001 ;
	    RECT 597.0000 1086.3000 598.2000 1106.7001 ;
	    RECT 599.4000 1086.3000 600.6000 1106.7001 ;
	    RECT 601.8000 1086.3000 603.0000 1106.7001 ;
	    RECT 594.6000 1079.4000 595.8000 1080.6000 ;
	    RECT 592.2000 1064.4000 593.4000 1065.6000 ;
	    RECT 594.7500 1062.6000 595.6500 1079.4000 ;
	    RECT 594.6000 1061.4000 595.8000 1062.6000 ;
	    RECT 601.8000 1058.4000 603.0000 1059.6000 ;
	    RECT 601.9500 1002.6000 602.8500 1058.4000 ;
	    RECT 606.7500 1056.6000 607.6500 1418.4000 ;
	    RECT 613.9500 1368.6000 614.8500 1424.4000 ;
	    RECT 649.9500 1422.6000 650.8500 1424.5500 ;
	    RECT 647.4000 1421.4000 648.6000 1422.6000 ;
	    RECT 649.8000 1421.4000 651.0000 1422.6000 ;
	    RECT 647.5500 1419.6000 648.4500 1421.4000 ;
	    RECT 625.8000 1418.4000 627.0000 1419.6000 ;
	    RECT 647.4000 1418.4000 648.6000 1419.6000 ;
	    RECT 613.8000 1367.4000 615.0000 1368.6000 ;
	    RECT 623.4000 1367.4000 624.6000 1368.6000 ;
	    RECT 609.0000 1319.4000 610.2000 1320.6000 ;
	    RECT 609.1500 1281.6000 610.0500 1319.4000 ;
	    RECT 618.6000 1307.4000 619.8000 1308.6000 ;
	    RECT 618.7500 1296.6000 619.6500 1307.4000 ;
	    RECT 618.6000 1295.4000 619.8000 1296.6000 ;
	    RECT 609.0000 1280.4000 610.2000 1281.6000 ;
	    RECT 618.7500 1275.6000 619.6500 1295.4000 ;
	    RECT 621.0000 1283.4000 622.2000 1284.6000 ;
	    RECT 618.6000 1274.4000 619.8000 1275.6000 ;
	    RECT 611.4000 1271.4000 612.6000 1272.6000 ;
	    RECT 611.5500 1242.6000 612.4500 1271.4000 ;
	    RECT 613.8000 1250.4000 615.0000 1251.6000 ;
	    RECT 611.4000 1241.4000 612.6000 1242.6000 ;
	    RECT 609.0000 1196.4000 610.2000 1197.6000 ;
	    RECT 606.6000 1055.4000 607.8000 1056.6000 ;
	    RECT 609.1500 1053.4501 610.0500 1196.4000 ;
	    RECT 613.9500 1179.6000 614.8500 1250.4000 ;
	    RECT 613.8000 1178.4000 615.0000 1179.6000 ;
	    RECT 616.2000 1169.4000 617.4000 1170.6000 ;
	    RECT 613.8000 1160.4000 615.0000 1161.6000 ;
	    RECT 611.4000 1157.4000 612.6000 1158.6000 ;
	    RECT 606.7500 1052.5500 610.0500 1053.4501 ;
	    RECT 601.8000 1001.4000 603.0000 1002.6000 ;
	    RECT 589.8000 983.4000 591.0000 984.6000 ;
	    RECT 575.4000 935.4000 576.6000 936.6000 ;
	    RECT 587.4000 929.4000 588.6000 930.6000 ;
	    RECT 573.0000 905.4000 574.2000 906.6000 ;
	    RECT 573.0000 899.4000 574.2000 900.6000 ;
	    RECT 563.4000 876.3000 564.6000 896.7000 ;
	    RECT 565.8000 876.3000 567.0000 896.7000 ;
	    RECT 568.2000 876.3000 569.4000 896.7000 ;
	    RECT 570.6000 876.3000 571.8000 893.7000 ;
	    RECT 573.1500 879.6000 574.0500 899.4000 ;
	    RECT 573.0000 878.4000 574.2000 879.6000 ;
	    RECT 575.4000 876.3000 576.6000 893.7000 ;
	    RECT 577.8000 881.4000 579.0000 882.6000 ;
	    RECT 577.9500 873.4500 578.8500 881.4000 ;
	    RECT 580.2000 876.3000 581.4000 893.7000 ;
	    RECT 582.6000 876.3000 583.8000 896.7000 ;
	    RECT 585.0000 876.3000 586.2000 896.7000 ;
	    RECT 587.5500 885.6000 588.4500 929.4000 ;
	    RECT 587.4000 884.4000 588.6000 885.6000 ;
	    RECT 575.5500 872.5500 578.8500 873.4500 ;
	    RECT 573.0000 863.4000 574.2000 864.6000 ;
	    RECT 563.4000 860.4000 564.6000 861.6000 ;
	    RECT 558.7500 854.5500 562.0500 855.4500 ;
	    RECT 551.5500 852.4500 552.4500 854.4000 ;
	    RECT 551.5500 851.5500 554.8500 852.4500 ;
	    RECT 553.9500 834.6000 554.8500 851.5500 ;
	    RECT 553.8000 833.4000 555.0000 834.6000 ;
	    RECT 551.4000 821.4000 552.6000 822.6000 ;
	    RECT 549.0000 761.4000 550.2000 762.6000 ;
	    RECT 539.4000 749.4000 540.6000 750.6000 ;
	    RECT 515.4000 743.4000 516.6000 744.6000 ;
	    RECT 515.5500 690.6000 516.4500 743.4000 ;
	    RECT 517.8000 729.3000 519.0000 746.7000 ;
	    RECT 520.2000 726.3000 521.4000 746.7000 ;
	    RECT 522.6000 726.3000 523.8000 746.7000 ;
	    RECT 525.0000 726.3000 526.2000 746.7000 ;
	    RECT 539.5500 732.6000 540.4500 749.4000 ;
	    RECT 546.6000 743.4000 547.8000 744.6000 ;
	    RECT 546.7500 738.6000 547.6500 743.4000 ;
	    RECT 546.6000 737.4000 547.8000 738.6000 ;
	    RECT 539.4000 731.4000 540.6000 732.6000 ;
	    RECT 501.0000 689.4000 502.2000 690.6000 ;
	    RECT 508.2000 689.4000 509.4000 690.6000 ;
	    RECT 515.4000 689.4000 516.6000 690.6000 ;
	    RECT 508.3500 678.6000 509.2500 689.4000 ;
	    RECT 508.2000 677.4000 509.4000 678.6000 ;
	    RECT 503.4000 656.4000 504.6000 657.6000 ;
	    RECT 503.5500 648.6000 504.4500 656.4000 ;
	    RECT 503.4000 647.4000 504.6000 648.6000 ;
	    RECT 508.3500 645.6000 509.2500 677.4000 ;
	    RECT 515.5500 672.6000 516.4500 689.4000 ;
	    RECT 515.4000 671.4000 516.6000 672.6000 ;
	    RECT 515.5500 660.6000 516.4500 671.4000 ;
	    RECT 515.4000 659.4000 516.6000 660.6000 ;
	    RECT 522.6000 659.4000 523.8000 660.6000 ;
	    RECT 508.2000 644.4000 509.4000 645.6000 ;
	    RECT 508.3500 621.6000 509.2500 644.4000 ;
	    RECT 510.6000 636.3000 511.8000 656.7000 ;
	    RECT 513.0000 636.3000 514.2000 656.7000 ;
	    RECT 515.4000 636.3000 516.6000 653.7000 ;
	    RECT 517.8000 641.4000 519.0000 642.6000 ;
	    RECT 520.2000 636.3000 521.4000 653.7000 ;
	    RECT 522.7500 639.6000 523.6500 659.4000 ;
	    RECT 522.6000 638.4000 523.8000 639.6000 ;
	    RECT 522.7500 624.4500 523.6500 638.4000 ;
	    RECT 525.0000 636.3000 526.2000 653.7000 ;
	    RECT 527.4000 636.3000 528.6000 656.7000 ;
	    RECT 529.8000 636.3000 531.0000 656.7000 ;
	    RECT 532.2000 636.3000 533.4000 656.7000 ;
	    RECT 546.7500 651.6000 547.6500 737.4000 ;
	    RECT 551.4000 653.4000 552.6000 654.6000 ;
	    RECT 546.6000 650.4000 547.8000 651.6000 ;
	    RECT 546.7500 624.6000 547.6500 650.4000 ;
	    RECT 522.7500 623.5500 526.0500 624.4500 ;
	    RECT 508.2000 620.4000 509.4000 621.6000 ;
	    RECT 522.6000 620.4000 523.8000 621.6000 ;
	    RECT 498.6000 608.4000 499.8000 609.6000 ;
	    RECT 520.2000 608.4000 521.4000 609.6000 ;
	    RECT 474.6000 605.4000 475.8000 606.6000 ;
	    RECT 489.0000 593.4000 490.2000 594.6000 ;
	    RECT 489.1500 588.6000 490.0500 593.4000 ;
	    RECT 489.0000 587.4000 490.2000 588.6000 ;
	    RECT 462.6000 584.4000 463.8000 585.6000 ;
	    RECT 457.8000 581.4000 459.0000 582.6000 ;
	    RECT 484.2000 581.4000 485.4000 582.6000 ;
	    RECT 486.6000 581.4000 487.8000 582.6000 ;
	    RECT 489.0000 581.4000 490.2000 582.6000 ;
	    RECT 503.4000 581.4000 504.6000 582.6000 ;
	    RECT 515.4000 581.4000 516.6000 582.6000 ;
	    RECT 457.9500 522.6000 458.8500 581.4000 ;
	    RECT 457.8000 521.4000 459.0000 522.6000 ;
	    RECT 455.4000 500.4000 456.6000 501.6000 ;
	    RECT 467.4000 491.4000 468.6000 492.6000 ;
	    RECT 467.5500 462.6000 468.4500 491.4000 ;
	    RECT 469.8000 479.4000 471.0000 480.6000 ;
	    RECT 469.9500 462.6000 470.8500 479.4000 ;
	    RECT 421.8000 461.4000 423.0000 462.6000 ;
	    RECT 450.6000 461.4000 451.8000 462.6000 ;
	    RECT 453.0000 461.4000 454.2000 462.6000 ;
	    RECT 467.4000 461.4000 468.6000 462.6000 ;
	    RECT 469.8000 461.4000 471.0000 462.6000 ;
	    RECT 421.9500 417.6000 422.8500 461.4000 ;
	    RECT 453.1500 459.6000 454.0500 461.4000 ;
	    RECT 453.0000 458.4000 454.2000 459.6000 ;
	    RECT 467.4000 458.4000 468.6000 459.6000 ;
	    RECT 453.1500 444.6000 454.0500 458.4000 ;
	    RECT 424.2000 443.4000 425.4000 444.6000 ;
	    RECT 453.0000 443.4000 454.2000 444.6000 ;
	    RECT 421.8000 416.4000 423.0000 417.6000 ;
	    RECT 424.3500 411.6000 425.2500 443.4000 ;
	    RECT 429.0000 440.4000 430.2000 441.6000 ;
	    RECT 462.6000 440.4000 463.8000 441.6000 ;
	    RECT 424.2000 410.4000 425.4000 411.6000 ;
	    RECT 429.1500 348.6000 430.0500 440.4000 ;
	    RECT 448.2000 419.4000 449.4000 420.6000 ;
	    RECT 431.4000 353.4000 432.6000 354.6000 ;
	    RECT 417.0000 347.4000 418.2000 348.6000 ;
	    RECT 429.0000 347.4000 430.2000 348.6000 ;
	    RECT 405.0000 341.4000 406.2000 342.6000 ;
	    RECT 409.8000 341.4000 411.0000 342.6000 ;
	    RECT 405.1500 300.6000 406.0500 341.4000 ;
	    RECT 407.4000 335.4000 408.6000 336.6000 ;
	    RECT 407.5500 312.6000 408.4500 335.4000 ;
	    RECT 407.4000 311.4000 408.6000 312.6000 ;
	    RECT 417.1500 300.6000 418.0500 347.4000 ;
	    RECT 421.8000 341.4000 423.0000 342.6000 ;
	    RECT 421.9500 330.6000 422.8500 341.4000 ;
	    RECT 421.8000 329.4000 423.0000 330.6000 ;
	    RECT 419.4000 305.4000 420.6000 306.6000 ;
	    RECT 421.8000 306.3000 423.0000 326.7000 ;
	    RECT 424.2000 306.3000 425.4000 326.7000 ;
	    RECT 426.6000 306.3000 427.8000 326.7000 ;
	    RECT 429.0000 309.3000 430.2000 326.7000 ;
	    RECT 431.5500 324.6000 432.4500 353.4000 ;
	    RECT 448.3500 348.6000 449.2500 419.4000 ;
	    RECT 462.7500 408.6000 463.6500 440.4000 ;
	    RECT 467.5500 420.6000 468.4500 458.4000 ;
	    RECT 467.4000 419.4000 468.6000 420.6000 ;
	    RECT 462.6000 407.4000 463.8000 408.6000 ;
	    RECT 469.8000 401.4000 471.0000 402.6000 ;
	    RECT 448.2000 347.4000 449.4000 348.6000 ;
	    RECT 469.9500 342.6000 470.8500 401.4000 ;
	    RECT 474.6000 347.4000 475.8000 348.6000 ;
	    RECT 474.7500 345.6000 475.6500 347.4000 ;
	    RECT 474.6000 344.4000 475.8000 345.6000 ;
	    RECT 441.0000 341.4000 442.2000 342.6000 ;
	    RECT 445.8000 341.4000 447.0000 342.6000 ;
	    RECT 469.8000 341.4000 471.0000 342.6000 ;
	    RECT 441.1500 336.6000 442.0500 341.4000 ;
	    RECT 441.0000 335.4000 442.2000 336.6000 ;
	    RECT 431.4000 323.4000 432.6000 324.6000 ;
	    RECT 433.8000 309.3000 435.0000 326.7000 ;
	    RECT 436.2000 323.4000 437.4000 324.6000 ;
	    RECT 436.3500 321.6000 437.2500 323.4000 ;
	    RECT 436.2000 320.4000 437.4000 321.6000 ;
	    RECT 438.6000 309.3000 439.8000 326.7000 ;
	    RECT 441.0000 306.3000 442.2000 326.7000 ;
	    RECT 443.4000 306.3000 444.6000 326.7000 ;
	    RECT 445.9500 324.6000 446.8500 341.4000 ;
	    RECT 445.8000 323.4000 447.0000 324.6000 ;
	    RECT 457.8000 320.4000 459.0000 321.6000 ;
	    RECT 479.4000 320.4000 480.6000 321.6000 ;
	    RECT 457.9500 318.6000 458.8500 320.4000 ;
	    RECT 445.8000 317.4000 447.0000 318.6000 ;
	    RECT 457.8000 317.4000 459.0000 318.6000 ;
	    RECT 450.6000 314.4000 451.8000 315.6000 ;
	    RECT 450.7500 306.6000 451.6500 314.4000 ;
	    RECT 450.6000 305.4000 451.8000 306.6000 ;
	    RECT 405.0000 299.4000 406.2000 300.6000 ;
	    RECT 417.0000 299.4000 418.2000 300.6000 ;
	    RECT 405.0000 263.4000 406.2000 264.6000 ;
	    RECT 405.1500 210.6000 406.0500 263.4000 ;
	    RECT 419.5500 246.6000 420.4500 305.4000 ;
	    RECT 450.6000 302.4000 451.8000 303.6000 ;
	    RECT 450.7500 300.6000 451.6500 302.4000 ;
	    RECT 450.6000 299.4000 451.8000 300.6000 ;
	    RECT 453.0000 284.4000 454.2000 285.6000 ;
	    RECT 445.8000 260.4000 447.0000 261.6000 ;
	    RECT 419.4000 245.4000 420.6000 246.6000 ;
	    RECT 431.4000 245.4000 432.6000 246.6000 ;
	    RECT 443.4000 245.4000 444.6000 246.6000 ;
	    RECT 407.4000 216.3000 408.6000 236.7000 ;
	    RECT 409.8000 216.3000 411.0000 236.7000 ;
	    RECT 412.2000 216.3000 413.4000 236.7000 ;
	    RECT 414.6000 216.3000 415.8000 233.7000 ;
	    RECT 417.0000 218.4000 418.2000 219.6000 ;
	    RECT 405.0000 209.4000 406.2000 210.6000 ;
	    RECT 402.6000 167.4000 403.8000 168.6000 ;
	    RECT 417.1500 150.6000 418.0500 218.4000 ;
	    RECT 419.4000 216.3000 420.6000 233.7000 ;
	    RECT 421.8000 227.4000 423.0000 228.6000 ;
	    RECT 421.9500 222.6000 422.8500 227.4000 ;
	    RECT 421.8000 221.4000 423.0000 222.6000 ;
	    RECT 424.2000 216.3000 425.4000 233.7000 ;
	    RECT 426.6000 216.3000 427.8000 236.7000 ;
	    RECT 429.0000 216.3000 430.2000 236.7000 ;
	    RECT 431.5500 225.6000 432.4500 245.4000 ;
	    RECT 436.2000 236.4000 437.4000 237.6000 ;
	    RECT 436.3500 228.6000 437.2500 236.4000 ;
	    RECT 436.2000 227.4000 437.4000 228.6000 ;
	    RECT 431.4000 224.4000 432.6000 225.6000 ;
	    RECT 431.5500 180.6000 432.4500 224.4000 ;
	    RECT 443.5500 222.6000 444.4500 245.4000 ;
	    RECT 443.4000 221.4000 444.6000 222.6000 ;
	    RECT 431.4000 179.4000 432.6000 180.6000 ;
	    RECT 421.8000 156.3000 423.0000 176.7000 ;
	    RECT 424.2000 156.3000 425.4000 176.7000 ;
	    RECT 426.6000 156.3000 427.8000 176.7000 ;
	    RECT 429.0000 156.3000 430.2000 173.7000 ;
	    RECT 431.4000 158.4000 432.6000 159.6000 ;
	    RECT 431.5500 150.6000 432.4500 158.4000 ;
	    RECT 433.8000 156.3000 435.0000 173.7000 ;
	    RECT 436.2000 167.4000 437.4000 168.6000 ;
	    RECT 436.3500 162.6000 437.2500 167.4000 ;
	    RECT 436.2000 161.4000 437.4000 162.6000 ;
	    RECT 438.6000 156.3000 439.8000 173.7000 ;
	    RECT 441.0000 156.3000 442.2000 176.7000 ;
	    RECT 443.4000 156.3000 444.6000 176.7000 ;
	    RECT 445.9500 165.6000 446.8500 260.4000 ;
	    RECT 450.6000 176.4000 451.8000 177.6000 ;
	    RECT 450.7500 168.6000 451.6500 176.4000 ;
	    RECT 450.6000 167.4000 451.8000 168.6000 ;
	    RECT 445.8000 164.4000 447.0000 165.6000 ;
	    RECT 417.0000 149.4000 418.2000 150.6000 ;
	    RECT 431.4000 149.4000 432.6000 150.6000 ;
	    RECT 424.2000 143.4000 425.4000 144.6000 ;
	    RECT 397.8000 116.4000 399.0000 117.6000 ;
	    RECT 397.9500 42.6000 398.8500 116.4000 ;
	    RECT 421.8000 101.4000 423.0000 102.6000 ;
	    RECT 421.9500 42.6000 422.8500 101.4000 ;
	    RECT 424.3500 42.6000 425.2500 143.4000 ;
	    RECT 445.9500 120.6000 446.8500 164.4000 ;
	    RECT 453.1500 120.6000 454.0500 284.4000 ;
	    RECT 479.5500 264.6000 480.4500 320.4000 ;
	    RECT 484.3500 279.6000 485.2500 581.4000 ;
	    RECT 486.7500 576.6000 487.6500 581.4000 ;
	    RECT 486.6000 575.4000 487.8000 576.6000 ;
	    RECT 489.1500 564.6000 490.0500 581.4000 ;
	    RECT 503.5500 576.6000 504.4500 581.4000 ;
	    RECT 515.5500 576.6000 516.4500 581.4000 ;
	    RECT 520.3500 579.6000 521.2500 608.4000 ;
	    RECT 520.2000 578.4000 521.4000 579.6000 ;
	    RECT 503.4000 575.4000 504.6000 576.6000 ;
	    RECT 515.4000 575.4000 516.6000 576.6000 ;
	    RECT 510.6000 569.4000 511.8000 570.6000 ;
	    RECT 489.0000 563.4000 490.2000 564.6000 ;
	    RECT 510.7500 555.6000 511.6500 569.4000 ;
	    RECT 515.5500 555.6000 516.4500 575.4000 ;
	    RECT 510.6000 554.4000 511.8000 555.6000 ;
	    RECT 515.4000 554.4000 516.6000 555.6000 ;
	    RECT 515.5500 546.4500 516.4500 554.4000 ;
	    RECT 520.3500 552.6000 521.2500 578.4000 ;
	    RECT 522.7500 558.6000 523.6500 620.4000 ;
	    RECT 525.1500 576.6000 526.0500 623.5500 ;
	    RECT 546.6000 623.4000 547.8000 624.6000 ;
	    RECT 537.0000 587.4000 538.2000 588.6000 ;
	    RECT 537.1500 582.6000 538.0500 587.4000 ;
	    RECT 537.0000 581.4000 538.2000 582.6000 ;
	    RECT 525.0000 575.4000 526.2000 576.6000 ;
	    RECT 537.0000 575.4000 538.2000 576.6000 ;
	    RECT 522.6000 557.4000 523.8000 558.6000 ;
	    RECT 520.2000 551.4000 521.4000 552.6000 ;
	    RECT 517.8000 546.4500 519.0000 546.6000 ;
	    RECT 515.5500 545.5500 519.0000 546.4500 ;
	    RECT 517.8000 545.4000 519.0000 545.5500 ;
	    RECT 517.9500 528.6000 518.8500 545.4000 ;
	    RECT 517.8000 527.4000 519.0000 528.6000 ;
	    RECT 522.7500 525.6000 523.6500 557.4000 ;
	    RECT 525.0000 546.3000 526.2000 566.7000 ;
	    RECT 527.4000 546.3000 528.6000 566.7000 ;
	    RECT 529.8000 549.3000 531.0000 566.7000 ;
	    RECT 532.2000 563.4000 533.4000 564.6000 ;
	    RECT 532.3500 561.6000 533.2500 563.4000 ;
	    RECT 532.2000 560.4000 533.4000 561.6000 ;
	    RECT 534.6000 549.3000 535.8000 566.7000 ;
	    RECT 537.1500 564.6000 538.0500 575.4000 ;
	    RECT 537.0000 563.4000 538.2000 564.6000 ;
	    RECT 539.4000 549.3000 540.6000 566.7000 ;
	    RECT 541.8000 546.3000 543.0000 566.7000 ;
	    RECT 544.2000 546.3000 545.4000 566.7000 ;
	    RECT 546.6000 546.3000 547.8000 566.7000 ;
	    RECT 522.6000 524.4000 523.8000 525.6000 ;
	    RECT 525.0000 516.3000 526.2000 536.7000 ;
	    RECT 527.4000 516.3000 528.6000 536.7000 ;
	    RECT 529.8000 516.3000 531.0000 533.7000 ;
	    RECT 532.2000 521.4000 533.4000 522.6000 ;
	    RECT 534.6000 516.3000 535.8000 533.7000 ;
	    RECT 537.0000 521.4000 538.2000 522.6000 ;
	    RECT 537.1500 519.6000 538.0500 521.4000 ;
	    RECT 537.0000 518.4000 538.2000 519.6000 ;
	    RECT 496.2000 509.4000 497.4000 510.6000 ;
	    RECT 486.6000 486.3000 487.8000 506.7000 ;
	    RECT 489.0000 486.3000 490.2000 506.7000 ;
	    RECT 491.4000 486.3000 492.6000 506.7000 ;
	    RECT 493.8000 489.3000 495.0000 506.7000 ;
	    RECT 496.3500 504.6000 497.2500 509.4000 ;
	    RECT 496.2000 503.4000 497.4000 504.6000 ;
	    RECT 486.6000 443.4000 487.8000 444.6000 ;
	    RECT 491.4000 443.4000 492.6000 444.6000 ;
	    RECT 486.7500 441.6000 487.6500 443.4000 ;
	    RECT 486.6000 440.4000 487.8000 441.6000 ;
	    RECT 496.3500 417.4500 497.2500 503.4000 ;
	    RECT 498.6000 489.3000 499.8000 506.7000 ;
	    RECT 501.0000 500.4000 502.2000 501.6000 ;
	    RECT 501.1500 498.6000 502.0500 500.4000 ;
	    RECT 501.0000 497.4000 502.2000 498.6000 ;
	    RECT 503.4000 489.3000 504.6000 506.7000 ;
	    RECT 505.8000 486.3000 507.0000 506.7000 ;
	    RECT 508.2000 486.3000 509.4000 506.7000 ;
	    RECT 537.1500 504.6000 538.0500 518.4000 ;
	    RECT 539.4000 516.3000 540.6000 533.7000 ;
	    RECT 541.8000 516.3000 543.0000 536.7000 ;
	    RECT 544.2000 516.3000 545.4000 536.7000 ;
	    RECT 546.6000 516.3000 547.8000 536.7000 ;
	    RECT 539.4000 509.4000 540.6000 510.6000 ;
	    RECT 537.0000 503.4000 538.2000 504.6000 ;
	    RECT 539.5500 501.6000 540.4500 509.4000 ;
	    RECT 539.4000 500.4000 540.6000 501.6000 ;
	    RECT 510.6000 497.4000 511.8000 498.6000 ;
	    RECT 510.7500 492.6000 511.6500 497.4000 ;
	    RECT 515.4000 494.4000 516.6000 495.6000 ;
	    RECT 515.5500 492.6000 516.4500 494.4000 ;
	    RECT 510.6000 491.4000 511.8000 492.6000 ;
	    RECT 515.4000 491.4000 516.6000 492.6000 ;
	    RECT 515.5500 486.6000 516.4500 491.4000 ;
	    RECT 515.4000 485.4000 516.6000 486.6000 ;
	    RECT 549.0000 455.4000 550.2000 456.6000 ;
	    RECT 522.6000 440.4000 523.8000 441.6000 ;
	    RECT 489.0000 396.3000 490.2000 416.7000 ;
	    RECT 491.4000 396.3000 492.6000 416.7000 ;
	    RECT 493.8000 396.3000 495.0000 416.7000 ;
	    RECT 496.3500 416.5500 499.6500 417.4500 ;
	    RECT 496.2000 396.3000 497.4000 413.7000 ;
	    RECT 498.7500 399.6000 499.6500 416.5500 ;
	    RECT 498.6000 398.4000 499.8000 399.6000 ;
	    RECT 498.7500 390.6000 499.6500 398.4000 ;
	    RECT 501.0000 396.3000 502.2000 413.7000 ;
	    RECT 503.4000 401.4000 504.6000 402.6000 ;
	    RECT 505.8000 396.3000 507.0000 413.7000 ;
	    RECT 508.2000 396.3000 509.4000 416.7000 ;
	    RECT 510.6000 396.3000 511.8000 416.7000 ;
	    RECT 517.8000 416.4000 519.0000 417.6000 ;
	    RECT 517.9500 408.6000 518.8500 416.4000 ;
	    RECT 513.0000 407.4000 514.2000 408.6000 ;
	    RECT 517.8000 407.4000 519.0000 408.6000 ;
	    RECT 513.1500 405.6000 514.0500 407.4000 ;
	    RECT 513.0000 404.4000 514.2000 405.6000 ;
	    RECT 498.6000 389.4000 499.8000 390.6000 ;
	    RECT 508.2000 389.4000 509.4000 390.6000 ;
	    RECT 498.6000 366.3000 499.8000 386.7000 ;
	    RECT 501.0000 366.3000 502.2000 386.7000 ;
	    RECT 503.4000 366.3000 504.6000 386.7000 ;
	    RECT 505.8000 369.3000 507.0000 386.7000 ;
	    RECT 508.3500 384.6000 509.2500 389.4000 ;
	    RECT 508.2000 383.4000 509.4000 384.6000 ;
	    RECT 508.3500 354.6000 509.2500 383.4000 ;
	    RECT 510.6000 369.3000 511.8000 386.7000 ;
	    RECT 513.0000 383.4000 514.2000 384.6000 ;
	    RECT 513.1500 381.6000 514.0500 383.4000 ;
	    RECT 513.0000 380.4000 514.2000 381.6000 ;
	    RECT 515.4000 369.3000 516.6000 386.7000 ;
	    RECT 517.8000 366.3000 519.0000 386.7000 ;
	    RECT 520.2000 366.3000 521.4000 386.7000 ;
	    RECT 522.7500 378.6000 523.6500 440.4000 ;
	    RECT 537.0000 398.4000 538.2000 399.6000 ;
	    RECT 522.6000 377.4000 523.8000 378.6000 ;
	    RECT 534.6000 377.4000 535.8000 378.6000 ;
	    RECT 527.4000 374.4000 528.6000 375.6000 ;
	    RECT 527.5500 366.6000 528.4500 374.4000 ;
	    RECT 527.4000 365.4000 528.6000 366.6000 ;
	    RECT 508.2000 353.4000 509.4000 354.6000 ;
	    RECT 501.0000 341.4000 502.2000 342.6000 ;
	    RECT 501.1500 300.6000 502.0500 341.4000 ;
	    RECT 534.7500 324.6000 535.6500 377.4000 ;
	    RECT 537.1500 351.6000 538.0500 398.4000 ;
	    RECT 537.0000 350.4000 538.2000 351.6000 ;
	    RECT 544.2000 350.4000 545.4000 351.6000 ;
	    RECT 527.4000 323.4000 528.6000 324.6000 ;
	    RECT 534.6000 323.4000 535.8000 324.6000 ;
	    RECT 527.5500 315.6000 528.4500 323.4000 ;
	    RECT 529.8000 320.4000 531.0000 321.6000 ;
	    RECT 537.0000 320.4000 538.2000 321.6000 ;
	    RECT 527.4000 314.4000 528.6000 315.6000 ;
	    RECT 501.0000 299.4000 502.2000 300.6000 ;
	    RECT 501.1500 282.6000 502.0500 299.4000 ;
	    RECT 501.0000 281.4000 502.2000 282.6000 ;
	    RECT 527.4000 281.4000 528.6000 282.6000 ;
	    RECT 484.2000 278.4000 485.4000 279.6000 ;
	    RECT 479.4000 263.4000 480.6000 264.6000 ;
	    RECT 479.5500 219.6000 480.4500 263.4000 ;
	    RECT 479.4000 218.4000 480.6000 219.6000 ;
	    RECT 484.3500 192.6000 485.2500 278.4000 ;
	    RECT 501.1500 249.6000 502.0500 281.4000 ;
	    RECT 510.6000 263.4000 511.8000 264.6000 ;
	    RECT 489.0000 248.4000 490.2000 249.6000 ;
	    RECT 501.0000 248.4000 502.2000 249.6000 ;
	    RECT 489.1500 222.6000 490.0500 248.4000 ;
	    RECT 496.2000 227.4000 497.4000 228.6000 ;
	    RECT 491.4000 224.4000 492.6000 225.6000 ;
	    RECT 491.5500 222.6000 492.4500 224.4000 ;
	    RECT 489.0000 221.4000 490.2000 222.6000 ;
	    RECT 491.4000 221.4000 492.6000 222.6000 ;
	    RECT 496.2000 221.4000 497.4000 222.6000 ;
	    RECT 498.6000 221.4000 499.8000 222.6000 ;
	    RECT 484.2000 191.4000 485.4000 192.6000 ;
	    RECT 457.8000 173.4000 459.0000 174.6000 ;
	    RECT 457.9500 168.6000 458.8500 173.4000 ;
	    RECT 457.8000 167.4000 459.0000 168.6000 ;
	    RECT 486.6000 161.4000 487.8000 162.6000 ;
	    RECT 493.8000 161.4000 495.0000 162.6000 ;
	    RECT 460.2000 140.4000 461.4000 141.6000 ;
	    RECT 457.8000 125.4000 459.0000 126.6000 ;
	    RECT 445.8000 119.4000 447.0000 120.6000 ;
	    RECT 453.0000 119.4000 454.2000 120.6000 ;
	    RECT 429.0000 116.4000 430.2000 117.6000 ;
	    RECT 429.1500 48.6000 430.0500 116.4000 ;
	    RECT 429.0000 47.4000 430.2000 48.6000 ;
	    RECT 457.9500 42.6000 458.8500 125.4000 ;
	    RECT 460.3500 45.6000 461.2500 140.4000 ;
	    RECT 486.7500 126.6000 487.6500 161.4000 ;
	    RECT 493.9500 132.6000 494.8500 161.4000 ;
	    RECT 496.3500 144.6000 497.2500 221.4000 ;
	    RECT 510.7500 165.6000 511.6500 263.4000 ;
	    RECT 513.0000 227.4000 514.2000 228.6000 ;
	    RECT 513.1500 225.6000 514.0500 227.4000 ;
	    RECT 513.0000 224.4000 514.2000 225.6000 ;
	    RECT 527.5500 216.6000 528.4500 281.4000 ;
	    RECT 529.9500 264.6000 530.8500 320.4000 ;
	    RECT 537.1500 279.4500 538.0500 320.4000 ;
	    RECT 544.3500 288.6000 545.2500 350.4000 ;
	    RECT 544.2000 287.4000 545.4000 288.6000 ;
	    RECT 539.4000 281.4000 540.6000 282.6000 ;
	    RECT 539.5500 279.4500 540.4500 281.4000 ;
	    RECT 537.1500 278.5500 540.4500 279.4500 ;
	    RECT 534.6000 269.4000 535.8000 270.6000 ;
	    RECT 529.8000 263.4000 531.0000 264.6000 ;
	    RECT 529.8000 221.4000 531.0000 222.6000 ;
	    RECT 532.2000 221.4000 533.4000 222.6000 ;
	    RECT 529.9500 219.6000 530.8500 221.4000 ;
	    RECT 529.8000 218.4000 531.0000 219.6000 ;
	    RECT 527.4000 215.4000 528.6000 216.6000 ;
	    RECT 529.8000 200.4000 531.0000 201.6000 ;
	    RECT 510.6000 164.4000 511.8000 165.6000 ;
	    RECT 517.8000 161.4000 519.0000 162.6000 ;
	    RECT 496.2000 143.4000 497.4000 144.6000 ;
	    RECT 493.8000 131.4000 495.0000 132.6000 ;
	    RECT 469.8000 125.4000 471.0000 126.6000 ;
	    RECT 486.6000 125.4000 487.8000 126.6000 ;
	    RECT 469.9500 120.6000 470.8500 125.4000 ;
	    RECT 469.8000 119.4000 471.0000 120.6000 ;
	    RECT 489.0000 119.4000 490.2000 120.6000 ;
	    RECT 469.8000 116.4000 471.0000 117.6000 ;
	    RECT 469.9500 108.6000 470.8500 116.4000 ;
	    RECT 469.8000 107.4000 471.0000 108.6000 ;
	    RECT 474.6000 107.4000 475.8000 108.6000 ;
	    RECT 474.7500 105.6000 475.6500 107.4000 ;
	    RECT 474.6000 104.4000 475.8000 105.6000 ;
	    RECT 477.0000 96.3000 478.2000 116.7000 ;
	    RECT 479.4000 96.3000 480.6000 116.7000 ;
	    RECT 481.8000 96.3000 483.0000 113.7000 ;
	    RECT 484.2000 101.4000 485.4000 102.6000 ;
	    RECT 486.6000 96.3000 487.8000 113.7000 ;
	    RECT 489.1500 99.6000 490.0500 119.4000 ;
	    RECT 489.0000 98.4000 490.2000 99.6000 ;
	    RECT 469.8000 47.4000 471.0000 48.6000 ;
	    RECT 460.2000 44.4000 461.4000 45.6000 ;
	    RECT 397.8000 41.4000 399.0000 42.6000 ;
	    RECT 421.8000 41.4000 423.0000 42.6000 ;
	    RECT 424.2000 41.4000 425.4000 42.6000 ;
	    RECT 457.8000 41.4000 459.0000 42.6000 ;
	    RECT 424.3500 12.6000 425.2500 41.4000 ;
	    RECT 469.9500 36.6000 470.8500 47.4000 ;
	    RECT 486.6000 41.4000 487.8000 42.6000 ;
	    RECT 469.8000 35.4000 471.0000 36.6000 ;
	    RECT 486.7500 24.6000 487.6500 41.4000 ;
	    RECT 489.1500 30.6000 490.0500 98.4000 ;
	    RECT 491.4000 96.3000 492.6000 113.7000 ;
	    RECT 493.8000 96.3000 495.0000 116.7000 ;
	    RECT 496.2000 96.3000 497.4000 116.7000 ;
	    RECT 498.6000 96.3000 499.8000 116.7000 ;
	    RECT 513.0000 113.4000 514.2000 114.6000 ;
	    RECT 513.1500 111.6000 514.0500 113.4000 ;
	    RECT 513.0000 110.4000 514.2000 111.6000 ;
	    RECT 491.4000 77.4000 492.6000 78.6000 ;
	    RECT 491.5500 42.6000 492.4500 77.4000 ;
	    RECT 493.8000 71.4000 495.0000 72.6000 ;
	    RECT 493.9500 60.6000 494.8500 71.4000 ;
	    RECT 508.2000 66.3000 509.4000 86.7000 ;
	    RECT 510.6000 66.3000 511.8000 86.7000 ;
	    RECT 513.0000 66.3000 514.2000 86.7000 ;
	    RECT 515.4000 69.3000 516.6000 86.7000 ;
	    RECT 517.9500 84.6000 518.8500 161.4000 ;
	    RECT 529.9500 138.6000 530.8500 200.4000 ;
	    RECT 532.3500 159.6000 533.2500 221.4000 ;
	    RECT 532.2000 158.4000 533.4000 159.6000 ;
	    RECT 529.8000 137.4000 531.0000 138.6000 ;
	    RECT 532.2000 134.4000 533.4000 135.6000 ;
	    RECT 532.3500 132.6000 533.2500 134.4000 ;
	    RECT 532.2000 131.4000 533.4000 132.6000 ;
	    RECT 532.3500 126.6000 533.2500 131.4000 ;
	    RECT 532.2000 125.4000 533.4000 126.6000 ;
	    RECT 517.8000 83.4000 519.0000 84.6000 ;
	    RECT 520.2000 69.3000 521.4000 86.7000 ;
	    RECT 522.6000 80.4000 523.8000 81.6000 ;
	    RECT 522.7500 78.6000 523.6500 80.4000 ;
	    RECT 522.6000 77.4000 523.8000 78.6000 ;
	    RECT 525.0000 69.3000 526.2000 86.7000 ;
	    RECT 527.4000 66.3000 528.6000 86.7000 ;
	    RECT 529.8000 66.3000 531.0000 86.7000 ;
	    RECT 532.2000 78.4500 533.4000 78.6000 ;
	    RECT 534.7500 78.4500 535.6500 269.4000 ;
	    RECT 539.5500 246.6000 540.4500 278.5500 ;
	    RECT 549.1500 258.6000 550.0500 455.4000 ;
	    RECT 551.5500 375.6000 552.4500 653.4000 ;
	    RECT 551.4000 374.4000 552.6000 375.6000 ;
	    RECT 558.7500 270.6000 559.6500 854.5500 ;
	    RECT 563.5500 822.6000 564.4500 860.4000 ;
	    RECT 575.5500 840.6000 576.4500 872.5500 ;
	    RECT 577.8000 863.4000 579.0000 864.6000 ;
	    RECT 577.8000 857.4000 579.0000 858.6000 ;
	    RECT 577.9500 846.6000 578.8500 857.4000 ;
	    RECT 577.8000 845.4000 579.0000 846.6000 ;
	    RECT 575.4000 839.4000 576.6000 840.6000 ;
	    RECT 582.6000 833.4000 583.8000 834.6000 ;
	    RECT 577.8000 827.4000 579.0000 828.6000 ;
	    RECT 577.9500 822.6000 578.8500 827.4000 ;
	    RECT 582.7500 825.6000 583.6500 833.4000 ;
	    RECT 582.6000 824.4000 583.8000 825.6000 ;
	    RECT 563.4000 821.4000 564.6000 822.6000 ;
	    RECT 570.6000 821.4000 571.8000 822.6000 ;
	    RECT 577.8000 821.4000 579.0000 822.6000 ;
	    RECT 563.5500 780.6000 564.4500 821.4000 ;
	    RECT 570.7500 804.6000 571.6500 821.4000 ;
	    RECT 573.0000 815.4000 574.2000 816.6000 ;
	    RECT 570.6000 803.4000 571.8000 804.6000 ;
	    RECT 573.1500 798.6000 574.0500 815.4000 ;
	    RECT 589.9500 810.4500 590.8500 983.4000 ;
	    RECT 592.2000 959.4000 593.4000 960.6000 ;
	    RECT 601.8000 959.4000 603.0000 960.6000 ;
	    RECT 592.3500 921.6000 593.2500 959.4000 ;
	    RECT 601.8000 957.4500 603.0000 957.6000 ;
	    RECT 601.8000 956.5500 605.2500 957.4500 ;
	    RECT 601.8000 956.4000 603.0000 956.5500 ;
	    RECT 594.6000 953.4000 595.8000 954.6000 ;
	    RECT 592.2000 920.4000 593.4000 921.6000 ;
	    RECT 592.2000 896.4000 593.4000 897.6000 ;
	    RECT 592.3500 888.6000 593.2500 896.4000 ;
	    RECT 592.2000 887.4000 593.4000 888.6000 ;
	    RECT 592.2000 869.4000 593.4000 870.6000 ;
	    RECT 592.3500 864.6000 593.2500 869.4000 ;
	    RECT 592.2000 863.4000 593.4000 864.6000 ;
	    RECT 594.7500 816.6000 595.6500 953.4000 ;
	    RECT 601.9500 948.6000 602.8500 956.4000 ;
	    RECT 601.8000 947.4000 603.0000 948.6000 ;
	    RECT 597.0000 941.4000 598.2000 942.6000 ;
	    RECT 597.1500 921.6000 598.0500 941.4000 ;
	    RECT 604.3500 921.6000 605.2500 956.5500 ;
	    RECT 606.7500 954.6000 607.6500 1052.5500 ;
	    RECT 613.9500 987.6000 614.8500 1160.4000 ;
	    RECT 616.3500 1158.6000 617.2500 1169.4000 ;
	    RECT 616.2000 1157.4000 617.4000 1158.6000 ;
	    RECT 616.2000 1115.4000 617.4000 1116.6000 ;
	    RECT 616.3500 1092.6000 617.2500 1115.4000 ;
	    RECT 618.6000 1094.4000 619.8000 1095.6000 ;
	    RECT 616.2000 1091.4000 617.4000 1092.6000 ;
	    RECT 618.7500 1080.6000 619.6500 1094.4000 ;
	    RECT 618.6000 1079.4000 619.8000 1080.6000 ;
	    RECT 618.6000 1001.4000 619.8000 1002.6000 ;
	    RECT 613.8000 986.4000 615.0000 987.6000 ;
	    RECT 618.7500 966.6000 619.6500 1001.4000 ;
	    RECT 621.1500 987.4500 622.0500 1283.4000 ;
	    RECT 623.5500 1230.6000 624.4500 1367.4000 ;
	    RECT 623.4000 1229.4000 624.6000 1230.6000 ;
	    RECT 625.9500 1221.6000 626.8500 1418.4000 ;
	    RECT 649.8000 1415.4000 651.0000 1416.6000 ;
	    RECT 645.0000 1406.4000 646.2000 1407.6000 ;
	    RECT 645.1500 1386.6000 646.0500 1406.4000 ;
	    RECT 649.9500 1395.6000 650.8500 1415.4000 ;
	    RECT 654.7500 1410.6000 655.6500 1439.4000 ;
	    RECT 659.4000 1427.4000 660.6000 1428.6000 ;
	    RECT 676.2000 1427.4000 677.4000 1428.6000 ;
	    RECT 681.0000 1427.4000 682.2000 1428.6000 ;
	    RECT 681.1500 1425.6000 682.0500 1427.4000 ;
	    RECT 681.0000 1424.4000 682.2000 1425.6000 ;
	    RECT 683.5500 1422.6000 684.4500 1442.4000 ;
	    RECT 657.0000 1421.4000 658.2000 1422.6000 ;
	    RECT 676.2000 1421.4000 677.4000 1422.6000 ;
	    RECT 683.4000 1421.4000 684.6000 1422.6000 ;
	    RECT 657.1500 1416.6000 658.0500 1421.4000 ;
	    RECT 676.3500 1416.6000 677.2500 1421.4000 ;
	    RECT 657.0000 1415.4000 658.2000 1416.6000 ;
	    RECT 676.2000 1415.4000 677.4000 1416.6000 ;
	    RECT 654.6000 1409.4000 655.8000 1410.6000 ;
	    RECT 666.6000 1409.4000 667.8000 1410.6000 ;
	    RECT 657.0000 1397.4000 658.2000 1398.6000 ;
	    RECT 649.8000 1394.4000 651.0000 1395.6000 ;
	    RECT 645.0000 1385.4000 646.2000 1386.6000 ;
	    RECT 633.0000 1370.4000 634.2000 1371.6000 ;
	    RECT 633.1500 1284.6000 634.0500 1370.4000 ;
	    RECT 637.8000 1367.4000 639.0000 1368.6000 ;
	    RECT 637.9500 1362.6000 638.8500 1367.4000 ;
	    RECT 637.8000 1361.4000 639.0000 1362.6000 ;
	    RECT 645.1500 1326.6000 646.0500 1385.4000 ;
	    RECT 649.9500 1356.6000 650.8500 1394.4000 ;
	    RECT 657.1500 1380.6000 658.0500 1397.4000 ;
	    RECT 659.4000 1386.3000 660.6000 1406.7001 ;
	    RECT 661.8000 1386.3000 663.0000 1406.7001 ;
	    RECT 664.2000 1389.3000 665.4000 1406.7001 ;
	    RECT 666.7500 1401.6000 667.6500 1409.4000 ;
	    RECT 666.6000 1400.4000 667.8000 1401.6000 ;
	    RECT 669.0000 1389.3000 670.2000 1406.7001 ;
	    RECT 671.4000 1403.4000 672.6000 1404.6000 ;
	    RECT 671.5500 1386.6000 672.4500 1403.4000 ;
	    RECT 673.8000 1389.3000 675.0000 1406.7001 ;
	    RECT 671.4000 1385.4000 672.6000 1386.6000 ;
	    RECT 676.2000 1386.3000 677.4000 1406.7001 ;
	    RECT 678.6000 1386.3000 679.8000 1406.7001 ;
	    RECT 681.0000 1386.3000 682.2000 1406.7001 ;
	    RECT 688.3500 1380.6000 689.2500 1457.4000 ;
	    RECT 690.6000 1446.3000 691.8000 1466.7001 ;
	    RECT 693.0000 1446.3000 694.2000 1466.7001 ;
	    RECT 695.4000 1449.3000 696.6000 1466.7001 ;
	    RECT 697.8000 1460.4000 699.0000 1461.6000 ;
	    RECT 697.9500 1458.6000 698.8500 1460.4000 ;
	    RECT 697.8000 1457.4000 699.0000 1458.6000 ;
	    RECT 700.2000 1449.3000 701.4000 1466.7001 ;
	    RECT 702.6000 1463.4000 703.8000 1464.6000 ;
	    RECT 705.0000 1449.3000 706.2000 1466.7001 ;
	    RECT 707.4000 1446.3000 708.6000 1466.7001 ;
	    RECT 709.8000 1446.3000 711.0000 1466.7001 ;
	    RECT 712.2000 1446.3000 713.4000 1466.7001 ;
	    RECT 726.6000 1451.4000 727.8000 1452.6000 ;
	    RECT 757.8000 1451.4000 759.0000 1452.6000 ;
	    RECT 856.2000 1451.4000 857.4000 1452.6000 ;
	    RECT 726.7500 1428.6000 727.6500 1451.4000 ;
	    RECT 748.2000 1445.4000 749.4000 1446.6000 ;
	    RECT 697.8000 1427.4000 699.0000 1428.6000 ;
	    RECT 726.6000 1427.4000 727.8000 1428.6000 ;
	    RECT 697.9500 1419.6000 698.8500 1427.4000 ;
	    RECT 697.8000 1418.4000 699.0000 1419.6000 ;
	    RECT 695.4000 1415.4000 696.6000 1416.6000 ;
	    RECT 695.5500 1392.6000 696.4500 1415.4000 ;
	    RECT 695.4000 1391.4000 696.6000 1392.6000 ;
	    RECT 652.2000 1379.4000 653.4000 1380.6000 ;
	    RECT 657.0000 1379.4000 658.2000 1380.6000 ;
	    RECT 688.2000 1379.4000 689.4000 1380.6000 ;
	    RECT 649.8000 1355.4000 651.0000 1356.6000 ;
	    RECT 645.0000 1325.4000 646.2000 1326.6000 ;
	    RECT 635.4000 1296.3000 636.6000 1316.7001 ;
	    RECT 637.8000 1296.3000 639.0000 1316.7001 ;
	    RECT 640.2000 1296.3000 641.4000 1316.7001 ;
	    RECT 642.6000 1296.3000 643.8000 1313.7001 ;
	    RECT 645.1500 1299.6000 646.0500 1325.4000 ;
	    RECT 649.9500 1320.6000 650.8500 1355.4000 ;
	    RECT 652.3500 1347.6000 653.2500 1379.4000 ;
	    RECT 654.6000 1356.3000 655.8000 1376.7001 ;
	    RECT 657.0000 1356.3000 658.2000 1376.7001 ;
	    RECT 659.4000 1356.3000 660.6000 1376.7001 ;
	    RECT 661.8000 1356.3000 663.0000 1373.7001 ;
	    RECT 664.2000 1358.4000 665.4000 1359.6000 ;
	    RECT 652.2000 1346.4000 653.4000 1347.6000 ;
	    RECT 659.4000 1346.4000 660.6000 1347.6000 ;
	    RECT 649.8000 1319.4000 651.0000 1320.6000 ;
	    RECT 649.9500 1314.6000 650.8500 1319.4000 ;
	    RECT 645.0000 1298.4000 646.2000 1299.6000 ;
	    RECT 635.4000 1289.4000 636.6000 1290.6000 ;
	    RECT 633.0000 1283.4000 634.2000 1284.6000 ;
	    RECT 635.5500 1281.6000 636.4500 1289.4000 ;
	    RECT 642.6000 1283.4000 643.8000 1284.6000 ;
	    RECT 635.4000 1280.4000 636.6000 1281.6000 ;
	    RECT 645.1500 1278.6000 646.0500 1298.4000 ;
	    RECT 647.4000 1296.3000 648.6000 1313.7001 ;
	    RECT 649.8000 1313.4000 651.0000 1314.6000 ;
	    RECT 649.8000 1301.4000 651.0000 1302.6000 ;
	    RECT 649.9500 1290.6000 650.8500 1301.4000 ;
	    RECT 652.2000 1296.3000 653.4000 1313.7001 ;
	    RECT 654.6000 1296.3000 655.8000 1316.7001 ;
	    RECT 657.0000 1296.3000 658.2000 1316.7001 ;
	    RECT 659.5500 1305.6000 660.4500 1346.4000 ;
	    RECT 664.3500 1344.6000 665.2500 1358.4000 ;
	    RECT 666.6000 1356.3000 667.8000 1373.7001 ;
	    RECT 669.0000 1361.4000 670.2000 1362.6000 ;
	    RECT 671.4000 1356.3000 672.6000 1373.7001 ;
	    RECT 673.8000 1356.3000 675.0000 1376.7001 ;
	    RECT 676.2000 1356.3000 677.4000 1376.7001 ;
	    RECT 683.4000 1376.4000 684.6000 1377.6000 ;
	    RECT 683.5500 1368.6000 684.4500 1376.4000 ;
	    RECT 697.9500 1368.6000 698.8500 1418.4000 ;
	    RECT 724.2000 1415.4000 725.4000 1416.6000 ;
	    RECT 724.3500 1401.6000 725.2500 1415.4000 ;
	    RECT 724.2000 1400.4000 725.4000 1401.6000 ;
	    RECT 741.0000 1400.4000 742.2000 1401.6000 ;
	    RECT 743.4000 1400.4000 744.6000 1401.6000 ;
	    RECT 729.0000 1397.4000 730.2000 1398.6000 ;
	    RECT 724.2000 1394.4000 725.4000 1395.6000 ;
	    RECT 683.4000 1367.4000 684.6000 1368.6000 ;
	    RECT 697.8000 1367.4000 699.0000 1368.6000 ;
	    RECT 714.6000 1367.4000 715.8000 1368.6000 ;
	    RECT 678.6000 1364.4000 679.8000 1365.6000 ;
	    RECT 678.7500 1347.6000 679.6500 1364.4000 ;
	    RECT 714.7500 1362.6000 715.6500 1367.4000 ;
	    RECT 724.3500 1365.6000 725.2500 1394.4000 ;
	    RECT 741.1500 1377.6000 742.0500 1400.4000 ;
	    RECT 743.5500 1398.6000 744.4500 1400.4000 ;
	    RECT 743.4000 1397.4000 744.6000 1398.6000 ;
	    RECT 741.0000 1376.4000 742.2000 1377.6000 ;
	    RECT 724.2000 1364.4000 725.4000 1365.6000 ;
	    RECT 695.4000 1361.4000 696.6000 1362.6000 ;
	    RECT 714.6000 1361.4000 715.8000 1362.6000 ;
	    RECT 719.4000 1361.4000 720.6000 1362.6000 ;
	    RECT 678.6000 1346.4000 679.8000 1347.6000 ;
	    RECT 664.2000 1343.4000 665.4000 1344.6000 ;
	    RECT 664.3500 1326.6000 665.2500 1343.4000 ;
	    RECT 678.7500 1338.6000 679.6500 1346.4000 ;
	    RECT 678.6000 1337.4000 679.8000 1338.6000 ;
	    RECT 664.2000 1325.4000 665.4000 1326.6000 ;
	    RECT 688.2000 1319.4000 689.4000 1320.6000 ;
	    RECT 664.2000 1316.4000 665.4000 1317.6000 ;
	    RECT 664.3500 1314.6000 665.2500 1316.4000 ;
	    RECT 664.2000 1313.4000 665.4000 1314.6000 ;
	    RECT 664.3500 1308.6000 665.2500 1313.4000 ;
	    RECT 664.2000 1307.4000 665.4000 1308.6000 ;
	    RECT 659.4000 1304.4000 660.6000 1305.6000 ;
	    RECT 649.8000 1289.4000 651.0000 1290.6000 ;
	    RECT 652.2000 1280.4000 653.4000 1281.6000 ;
	    RECT 645.0000 1277.4000 646.2000 1278.6000 ;
	    RECT 645.1500 1260.6000 646.0500 1277.4000 ;
	    RECT 652.3500 1260.6000 653.2500 1280.4000 ;
	    RECT 637.8000 1259.4000 639.0000 1260.6000 ;
	    RECT 645.0000 1259.4000 646.2000 1260.6000 ;
	    RECT 652.2000 1259.4000 653.4000 1260.6000 ;
	    RECT 657.0000 1259.4000 658.2000 1260.6000 ;
	    RECT 628.2000 1236.3000 629.4000 1256.7001 ;
	    RECT 630.6000 1236.3000 631.8000 1256.7001 ;
	    RECT 633.0000 1236.3000 634.2000 1256.7001 ;
	    RECT 635.4000 1236.3000 636.6000 1253.7001 ;
	    RECT 637.9500 1239.6000 638.8500 1259.4000 ;
	    RECT 657.1500 1257.6000 658.0500 1259.4000 ;
	    RECT 637.8000 1238.4000 639.0000 1239.6000 ;
	    RECT 640.2000 1236.3000 641.4000 1253.7001 ;
	    RECT 642.6000 1241.4000 643.8000 1242.6000 ;
	    RECT 642.7500 1236.6000 643.6500 1241.4000 ;
	    RECT 642.6000 1235.4000 643.8000 1236.6000 ;
	    RECT 645.0000 1236.3000 646.2000 1253.7001 ;
	    RECT 647.4000 1236.3000 648.6000 1256.7001 ;
	    RECT 649.8000 1236.3000 651.0000 1256.7001 ;
	    RECT 657.0000 1256.4000 658.2000 1257.6000 ;
	    RECT 657.1500 1251.6000 658.0500 1256.4000 ;
	    RECT 657.0000 1250.4000 658.2000 1251.6000 ;
	    RECT 657.1500 1248.6000 658.0500 1250.4000 ;
	    RECT 657.0000 1247.4000 658.2000 1248.6000 ;
	    RECT 652.2000 1244.4000 653.4000 1245.6000 ;
	    RECT 649.8000 1229.4000 651.0000 1230.6000 ;
	    RECT 649.9500 1224.6000 650.8500 1229.4000 ;
	    RECT 649.8000 1223.4000 651.0000 1224.6000 ;
	    RECT 625.8000 1220.4000 627.0000 1221.6000 ;
	    RECT 623.4000 1157.4000 624.6000 1158.6000 ;
	    RECT 623.5500 1155.6000 624.4500 1157.4000 ;
	    RECT 623.4000 1154.4000 624.6000 1155.6000 ;
	    RECT 625.9500 1146.6000 626.8500 1220.4000 ;
	    RECT 633.0000 1217.4000 634.2000 1218.6000 ;
	    RECT 640.2000 1217.4000 641.4000 1218.6000 ;
	    RECT 633.1500 1179.6000 634.0500 1217.4000 ;
	    RECT 633.0000 1178.4000 634.2000 1179.6000 ;
	    RECT 628.2000 1160.4000 629.4000 1161.6000 ;
	    RECT 625.8000 1145.4000 627.0000 1146.6000 ;
	    RECT 628.3500 1080.6000 629.2500 1160.4000 ;
	    RECT 633.1500 1110.6000 634.0500 1178.4000 ;
	    RECT 637.8000 1137.4501 639.0000 1137.6000 ;
	    RECT 635.5500 1136.5500 639.0000 1137.4501 ;
	    RECT 633.0000 1109.4000 634.2000 1110.6000 ;
	    RECT 635.5500 1104.6000 636.4500 1136.5500 ;
	    RECT 637.8000 1136.4000 639.0000 1136.5500 ;
	    RECT 637.9500 1128.6000 638.8500 1136.4000 ;
	    RECT 637.8000 1127.4000 639.0000 1128.6000 ;
	    RECT 635.4000 1103.4000 636.6000 1104.6000 ;
	    RECT 628.2000 1079.4000 629.4000 1080.6000 ;
	    RECT 625.8000 1068.4501 627.0000 1068.6000 ;
	    RECT 623.5500 1067.5500 627.0000 1068.4501 ;
	    RECT 623.5500 1065.6000 624.4500 1067.5500 ;
	    RECT 625.8000 1067.4000 627.0000 1067.5500 ;
	    RECT 635.4000 1067.4000 636.6000 1068.6000 ;
	    RECT 623.4000 1064.4000 624.6000 1065.6000 ;
	    RECT 637.8000 1064.4000 639.0000 1065.6000 ;
	    RECT 625.8000 1061.4000 627.0000 1062.6000 ;
	    RECT 628.2000 1061.4000 629.4000 1062.6000 ;
	    RECT 625.9500 1044.6000 626.8500 1061.4000 ;
	    RECT 628.3500 1059.6000 629.2500 1061.4000 ;
	    RECT 628.2000 1058.4000 629.4000 1059.6000 ;
	    RECT 625.8000 1043.4000 627.0000 1044.6000 ;
	    RECT 637.9500 1041.6000 638.8500 1064.4000 ;
	    RECT 640.3500 1044.6000 641.2500 1217.4000 ;
	    RECT 652.3500 1200.6000 653.2500 1244.4000 ;
	    RECT 657.0000 1220.4000 658.2000 1221.6000 ;
	    RECT 642.6000 1199.4000 643.8000 1200.6000 ;
	    RECT 652.2000 1199.4000 653.4000 1200.6000 ;
	    RECT 642.7500 1125.6000 643.6500 1199.4000 ;
	    RECT 642.6000 1124.4000 643.8000 1125.6000 ;
	    RECT 642.7500 1113.4501 643.6500 1124.4000 ;
	    RECT 645.0000 1116.3000 646.2000 1136.7001 ;
	    RECT 647.4000 1116.3000 648.6000 1136.7001 ;
	    RECT 657.1500 1134.6000 658.0500 1220.4000 ;
	    RECT 659.5500 1197.6000 660.4500 1304.4000 ;
	    RECT 688.3500 1299.6000 689.2500 1319.4000 ;
	    RECT 676.2000 1298.4000 677.4000 1299.6000 ;
	    RECT 688.2000 1298.4000 689.4000 1299.6000 ;
	    RECT 661.8000 1247.4000 663.0000 1248.6000 ;
	    RECT 661.9500 1221.6000 662.8500 1247.4000 ;
	    RECT 661.8000 1220.4000 663.0000 1221.6000 ;
	    RECT 659.4000 1196.4000 660.6000 1197.6000 ;
	    RECT 649.8000 1116.3000 651.0000 1133.7001 ;
	    RECT 652.2000 1121.4000 653.4000 1122.6000 ;
	    RECT 642.7500 1112.5500 646.0500 1113.4501 ;
	    RECT 642.6000 1103.4000 643.8000 1104.6000 ;
	    RECT 642.7500 1101.6000 643.6500 1103.4000 ;
	    RECT 642.6000 1100.4000 643.8000 1101.6000 ;
	    RECT 642.6000 1079.4000 643.8000 1080.6000 ;
	    RECT 640.2000 1043.4000 641.4000 1044.6000 ;
	    RECT 637.8000 1040.4000 639.0000 1041.6000 ;
	    RECT 640.3500 1038.6000 641.2500 1043.4000 ;
	    RECT 642.7500 1038.6000 643.6500 1079.4000 ;
	    RECT 633.0000 1037.4000 634.2000 1038.6000 ;
	    RECT 640.2000 1037.4000 641.4000 1038.6000 ;
	    RECT 642.6000 1037.4000 643.8000 1038.6000 ;
	    RECT 630.6000 1019.4000 631.8000 1020.6000 ;
	    RECT 625.8000 1013.4000 627.0000 1014.6000 ;
	    RECT 625.9500 1002.6000 626.8500 1013.4000 ;
	    RECT 628.2000 1007.7000 629.4000 1008.9000 ;
	    RECT 628.2000 1002.6000 629.1000 1007.7000 ;
	    RECT 630.7500 1005.6000 631.6500 1019.4000 ;
	    RECT 633.1500 1014.6000 634.0500 1037.4000 ;
	    RECT 633.0000 1013.4000 634.2000 1014.6000 ;
	    RECT 640.2000 1013.4000 641.4000 1014.6000 ;
	    RECT 637.5000 1007.7000 638.7000 1008.9000 ;
	    RECT 630.6000 1004.4000 631.8000 1005.6000 ;
	    RECT 635.7000 1004.7000 636.9000 1005.9000 ;
	    RECT 635.7000 1002.6000 636.6000 1004.7000 ;
	    RECT 625.8000 1001.4000 627.0000 1002.6000 ;
	    RECT 628.2000 1001.7000 636.6000 1002.6000 ;
	    RECT 628.2000 1000.5000 629.1000 1001.7000 ;
	    RECT 630.3000 1000.5000 631.5000 1000.8000 ;
	    RECT 635.4000 1000.5000 636.6000 1000.8000 ;
	    RECT 637.8000 1000.5000 638.7000 1007.7000 ;
	    RECT 623.4000 998.4000 624.6000 999.6000 ;
	    RECT 628.2000 999.3000 629.4000 1000.5000 ;
	    RECT 630.3000 999.6000 638.7000 1000.5000 ;
	    RECT 637.5000 999.3000 638.7000 999.6000 ;
	    RECT 623.5500 990.6000 624.4500 998.4000 ;
	    RECT 635.4000 995.4000 636.6000 996.6000 ;
	    RECT 623.4000 989.4000 624.6000 990.6000 ;
	    RECT 621.1500 986.5500 624.4500 987.4500 ;
	    RECT 623.5500 984.6000 624.4500 986.5500 ;
	    RECT 633.0000 986.4000 634.2000 987.6000 ;
	    RECT 621.0000 983.4000 622.2000 984.6000 ;
	    RECT 623.4000 983.4000 624.6000 984.6000 ;
	    RECT 618.6000 965.4000 619.8000 966.6000 ;
	    RECT 606.6000 953.4000 607.8000 954.6000 ;
	    RECT 606.7500 945.6000 607.6500 953.4000 ;
	    RECT 606.6000 944.4000 607.8000 945.6000 ;
	    RECT 609.0000 936.3000 610.2000 956.7000 ;
	    RECT 611.4000 936.3000 612.6000 956.7000 ;
	    RECT 621.1500 954.6000 622.0500 983.4000 ;
	    RECT 613.8000 936.3000 615.0000 953.7000 ;
	    RECT 616.2000 941.4000 617.4000 942.6000 ;
	    RECT 618.6000 936.3000 619.8000 953.7000 ;
	    RECT 621.0000 953.4000 622.2000 954.6000 ;
	    RECT 621.1500 939.6000 622.0500 953.4000 ;
	    RECT 621.0000 938.4000 622.2000 939.6000 ;
	    RECT 623.4000 936.3000 624.6000 953.7000 ;
	    RECT 625.8000 936.3000 627.0000 956.7000 ;
	    RECT 628.2000 936.3000 629.4000 956.7000 ;
	    RECT 630.6000 936.3000 631.8000 956.7000 ;
	    RECT 616.2000 929.4000 617.4000 930.6000 ;
	    RECT 597.0000 920.4000 598.2000 921.6000 ;
	    RECT 604.2000 920.4000 605.4000 921.6000 ;
	    RECT 599.4000 881.4000 600.6000 882.6000 ;
	    RECT 599.5500 864.6000 600.4500 881.4000 ;
	    RECT 611.4000 878.4000 612.6000 879.6000 ;
	    RECT 606.6000 869.4000 607.8000 870.6000 ;
	    RECT 606.7500 864.6000 607.6500 869.4000 ;
	    RECT 599.4000 863.4000 600.6000 864.6000 ;
	    RECT 606.6000 863.4000 607.8000 864.6000 ;
	    RECT 601.8000 857.4000 603.0000 858.6000 ;
	    RECT 606.6000 827.4000 607.8000 828.6000 ;
	    RECT 599.4000 821.4000 600.6000 822.6000 ;
	    RECT 594.6000 815.4000 595.8000 816.6000 ;
	    RECT 587.5500 809.5500 590.8500 810.4500 ;
	    RECT 573.0000 797.4000 574.2000 798.6000 ;
	    RECT 568.2000 794.4000 569.4000 795.6000 ;
	    RECT 568.3500 786.6000 569.2500 794.4000 ;
	    RECT 568.2000 785.4000 569.4000 786.6000 ;
	    RECT 563.4000 779.4000 564.6000 780.6000 ;
	    RECT 568.2000 737.4000 569.4000 738.6000 ;
	    RECT 568.3500 735.6000 569.2500 737.4000 ;
	    RECT 568.2000 734.4000 569.4000 735.6000 ;
	    RECT 563.4000 638.4000 564.6000 639.6000 ;
	    RECT 563.5500 588.6000 564.4500 638.4000 ;
	    RECT 563.4000 587.4000 564.6000 588.6000 ;
	    RECT 563.4000 581.4000 564.6000 582.6000 ;
	    RECT 561.0000 551.4000 562.2000 552.6000 ;
	    RECT 563.5500 531.6000 564.4500 581.4000 ;
	    RECT 570.6000 557.4000 571.8000 558.6000 ;
	    RECT 565.8000 533.4000 567.0000 534.6000 ;
	    RECT 563.4000 530.4000 564.6000 531.6000 ;
	    RECT 563.4000 383.4000 564.6000 384.6000 ;
	    RECT 563.5500 381.6000 564.4500 383.4000 ;
	    RECT 563.4000 380.4000 564.6000 381.6000 ;
	    RECT 563.4000 353.4000 564.6000 354.6000 ;
	    RECT 563.5500 330.6000 564.4500 353.4000 ;
	    RECT 563.4000 329.4000 564.6000 330.6000 ;
	    RECT 558.6000 269.4000 559.8000 270.6000 ;
	    RECT 549.0000 257.4000 550.2000 258.6000 ;
	    RECT 544.2000 254.4000 545.4000 255.6000 ;
	    RECT 544.3500 246.6000 545.2500 254.4000 ;
	    RECT 539.4000 245.4000 540.6000 246.6000 ;
	    RECT 544.2000 245.4000 545.4000 246.6000 ;
	    RECT 551.4000 246.3000 552.6000 266.7000 ;
	    RECT 553.8000 246.3000 555.0000 266.7000 ;
	    RECT 556.2000 249.3000 557.4000 266.7000 ;
	    RECT 558.6000 263.4000 559.8000 264.6000 ;
	    RECT 558.7500 261.6000 559.6500 263.4000 ;
	    RECT 558.6000 260.4000 559.8000 261.6000 ;
	    RECT 561.0000 249.3000 562.2000 266.7000 ;
	    RECT 563.5500 264.6000 564.4500 329.4000 ;
	    RECT 565.9500 324.6000 566.8500 533.4000 ;
	    RECT 568.2000 500.4000 569.4000 501.6000 ;
	    RECT 568.3500 480.6000 569.2500 500.4000 ;
	    RECT 570.7500 495.6000 571.6500 557.4000 ;
	    RECT 570.6000 494.4000 571.8000 495.6000 ;
	    RECT 568.2000 479.4000 569.4000 480.6000 ;
	    RECT 573.1500 456.6000 574.0500 797.4000 ;
	    RECT 575.4000 786.3000 576.6000 806.7000 ;
	    RECT 577.8000 786.3000 579.0000 806.7000 ;
	    RECT 580.2000 789.3000 581.4000 806.7000 ;
	    RECT 582.6000 803.4000 583.8000 804.6000 ;
	    RECT 582.7500 801.6000 583.6500 803.4000 ;
	    RECT 582.6000 800.4000 583.8000 801.6000 ;
	    RECT 585.0000 789.3000 586.2000 806.7000 ;
	    RECT 587.5500 804.6000 588.4500 809.5500 ;
	    RECT 587.4000 803.4000 588.6000 804.6000 ;
	    RECT 582.6000 785.4000 583.8000 786.6000 ;
	    RECT 582.7500 780.6000 583.6500 785.4000 ;
	    RECT 582.6000 779.4000 583.8000 780.6000 ;
	    RECT 582.7500 768.6000 583.6500 779.4000 ;
	    RECT 587.5500 774.6000 588.4500 803.4000 ;
	    RECT 589.8000 789.3000 591.0000 806.7000 ;
	    RECT 592.2000 786.3000 593.4000 806.7000 ;
	    RECT 594.6000 786.3000 595.8000 806.7000 ;
	    RECT 597.0000 786.3000 598.2000 806.7000 ;
	    RECT 599.5500 786.6000 600.4500 821.4000 ;
	    RECT 606.7500 804.6000 607.6500 827.4000 ;
	    RECT 606.6000 803.4000 607.8000 804.6000 ;
	    RECT 611.5500 792.6000 612.4500 878.4000 ;
	    RECT 613.8000 860.4000 615.0000 861.6000 ;
	    RECT 613.9500 852.6000 614.8500 860.4000 ;
	    RECT 613.8000 851.4000 615.0000 852.6000 ;
	    RECT 611.4000 791.4000 612.6000 792.6000 ;
	    RECT 599.4000 785.4000 600.6000 786.6000 ;
	    RECT 587.4000 773.4000 588.6000 774.6000 ;
	    RECT 582.6000 767.4000 583.8000 768.6000 ;
	    RECT 587.4000 767.4000 588.6000 768.6000 ;
	    RECT 587.5500 765.6000 588.4500 767.4000 ;
	    RECT 587.4000 765.4500 588.6000 765.6000 ;
	    RECT 585.1500 764.5500 588.6000 765.4500 ;
	    RECT 577.8000 740.4000 579.0000 741.6000 ;
	    RECT 577.9500 732.6000 578.8500 740.4000 ;
	    RECT 577.8000 731.4000 579.0000 732.6000 ;
	    RECT 575.4000 719.4000 576.6000 720.6000 ;
	    RECT 575.5500 606.6000 576.4500 719.4000 ;
	    RECT 582.6000 677.4000 583.8000 678.6000 ;
	    RECT 582.6000 653.4000 583.8000 654.6000 ;
	    RECT 577.8000 647.4000 579.0000 648.6000 ;
	    RECT 575.4000 605.4000 576.6000 606.6000 ;
	    RECT 575.5500 582.6000 576.4500 605.4000 ;
	    RECT 577.9500 585.6000 578.8500 647.4000 ;
	    RECT 582.7500 642.6000 583.6500 653.4000 ;
	    RECT 582.6000 641.4000 583.8000 642.6000 ;
	    RECT 580.2000 587.7000 581.4000 588.9000 ;
	    RECT 585.1500 588.6000 586.0500 764.5500 ;
	    RECT 587.4000 764.4000 588.6000 764.5500 ;
	    RECT 589.8000 756.3000 591.0000 776.7000 ;
	    RECT 592.2000 756.3000 593.4000 776.7000 ;
	    RECT 594.6000 756.3000 595.8000 773.7000 ;
	    RECT 597.0000 761.4000 598.2000 762.6000 ;
	    RECT 597.0000 755.4000 598.2000 756.6000 ;
	    RECT 599.4000 756.3000 600.6000 773.7000 ;
	    RECT 601.8000 758.4000 603.0000 759.6000 ;
	    RECT 592.2000 743.4000 593.4000 744.6000 ;
	    RECT 592.3500 741.6000 593.2500 743.4000 ;
	    RECT 592.2000 740.4000 593.4000 741.6000 ;
	    RECT 587.4000 701.4000 588.6000 702.6000 ;
	    RECT 587.5500 654.6000 588.4500 701.4000 ;
	    RECT 589.8000 695.4000 591.0000 696.6000 ;
	    RECT 589.9500 675.6000 590.8500 695.4000 ;
	    RECT 592.3500 687.4500 593.2500 740.4000 ;
	    RECT 594.6000 737.4000 595.8000 738.6000 ;
	    RECT 592.3500 686.5500 595.6500 687.4500 ;
	    RECT 589.8000 674.4000 591.0000 675.6000 ;
	    RECT 589.8000 671.4000 591.0000 672.6000 ;
	    RECT 587.4000 653.4000 588.6000 654.6000 ;
	    RECT 589.9500 642.6000 590.8500 671.4000 ;
	    RECT 592.2000 665.4000 593.4000 666.6000 ;
	    RECT 592.3500 648.6000 593.2500 665.4000 ;
	    RECT 592.2000 647.4000 593.4000 648.6000 ;
	    RECT 589.8000 641.4000 591.0000 642.6000 ;
	    RECT 592.2000 641.4000 593.4000 642.6000 ;
	    RECT 592.3500 624.6000 593.2500 641.4000 ;
	    RECT 592.2000 623.4000 593.4000 624.6000 ;
	    RECT 577.8000 584.4000 579.0000 585.6000 ;
	    RECT 580.2000 582.6000 581.1000 587.7000 ;
	    RECT 585.0000 587.4000 586.2000 588.6000 ;
	    RECT 589.5000 587.7000 590.7000 588.9000 ;
	    RECT 585.0000 584.4000 586.2000 585.6000 ;
	    RECT 587.7000 584.7000 588.9000 585.9000 ;
	    RECT 587.7000 582.6000 588.6000 584.7000 ;
	    RECT 575.4000 581.4000 576.6000 582.6000 ;
	    RECT 580.2000 581.7000 588.6000 582.6000 ;
	    RECT 580.2000 580.5000 581.1000 581.7000 ;
	    RECT 582.3000 580.5000 583.5000 580.8000 ;
	    RECT 587.4000 580.5000 588.6000 580.8000 ;
	    RECT 589.8000 580.5000 590.7000 587.7000 ;
	    RECT 580.2000 579.3000 581.4000 580.5000 ;
	    RECT 582.3000 579.6000 590.7000 580.5000 ;
	    RECT 589.5000 579.3000 590.7000 579.6000 ;
	    RECT 589.8000 575.4000 591.0000 576.6000 ;
	    RECT 582.6000 569.4000 583.8000 570.6000 ;
	    RECT 582.7500 555.6000 583.6500 569.4000 ;
	    RECT 587.4000 560.4000 588.6000 561.6000 ;
	    RECT 582.6000 554.4000 583.8000 555.6000 ;
	    RECT 587.5500 546.6000 588.4500 560.4000 ;
	    RECT 587.4000 545.4000 588.6000 546.6000 ;
	    RECT 575.4000 521.4000 576.6000 522.6000 ;
	    RECT 575.5500 498.6000 576.4500 521.4000 ;
	    RECT 577.8000 500.4000 579.0000 501.6000 ;
	    RECT 575.4000 497.4000 576.6000 498.6000 ;
	    RECT 577.9500 492.6000 578.8500 500.4000 ;
	    RECT 577.8000 491.4000 579.0000 492.6000 ;
	    RECT 582.6000 491.4000 583.8000 492.6000 ;
	    RECT 573.0000 455.4000 574.2000 456.6000 ;
	    RECT 580.2000 380.4000 581.4000 381.6000 ;
	    RECT 577.8000 374.4000 579.0000 375.6000 ;
	    RECT 577.9500 339.4500 578.8500 374.4000 ;
	    RECT 580.3500 342.6000 581.2500 380.4000 ;
	    RECT 580.2000 341.4000 581.4000 342.6000 ;
	    RECT 577.9500 338.5500 581.2500 339.4500 ;
	    RECT 565.8000 323.4000 567.0000 324.6000 ;
	    RECT 575.4000 323.4000 576.6000 324.6000 ;
	    RECT 568.2000 284.4000 569.4000 285.6000 ;
	    RECT 568.3500 282.6000 569.2500 284.4000 ;
	    RECT 568.2000 281.4000 569.4000 282.6000 ;
	    RECT 570.6000 281.4000 571.8000 282.6000 ;
	    RECT 570.7500 276.6000 571.6500 281.4000 ;
	    RECT 570.6000 275.4000 571.8000 276.6000 ;
	    RECT 563.4000 263.4000 564.6000 264.6000 ;
	    RECT 565.8000 249.3000 567.0000 266.7000 ;
	    RECT 568.2000 246.3000 569.4000 266.7000 ;
	    RECT 570.6000 246.3000 571.8000 266.7000 ;
	    RECT 573.0000 246.3000 574.2000 266.7000 ;
	    RECT 575.5500 258.6000 576.4500 323.4000 ;
	    RECT 577.8000 317.4000 579.0000 318.6000 ;
	    RECT 575.4000 257.4000 576.6000 258.6000 ;
	    RECT 575.4000 245.4000 576.6000 246.6000 ;
	    RECT 539.5500 228.6000 540.4500 245.4000 ;
	    RECT 565.8000 239.4000 567.0000 240.6000 ;
	    RECT 565.9500 228.6000 566.8500 239.4000 ;
	    RECT 539.4000 227.4000 540.6000 228.6000 ;
	    RECT 565.8000 227.4000 567.0000 228.6000 ;
	    RECT 575.5500 225.6000 576.4500 245.4000 ;
	    RECT 575.4000 224.4000 576.6000 225.6000 ;
	    RECT 546.6000 221.4000 547.8000 222.6000 ;
	    RECT 546.7500 156.6000 547.6500 221.4000 ;
	    RECT 575.4000 218.4000 576.6000 219.6000 ;
	    RECT 563.4000 215.4000 564.6000 216.6000 ;
	    RECT 573.0000 215.4000 574.2000 216.6000 ;
	    RECT 549.0000 186.3000 550.2000 206.7000 ;
	    RECT 551.4000 186.3000 552.6000 206.7000 ;
	    RECT 553.8000 186.3000 555.0000 206.7000 ;
	    RECT 556.2000 189.3000 557.4000 206.7000 ;
	    RECT 558.6000 203.4000 559.8000 204.6000 ;
	    RECT 558.7500 162.6000 559.6500 203.4000 ;
	    RECT 561.0000 189.3000 562.2000 206.7000 ;
	    RECT 563.5500 201.6000 564.4500 215.4000 ;
	    RECT 563.4000 200.4000 564.6000 201.6000 ;
	    RECT 565.8000 189.3000 567.0000 206.7000 ;
	    RECT 568.2000 186.3000 569.4000 206.7000 ;
	    RECT 570.6000 186.3000 571.8000 206.7000 ;
	    RECT 573.1500 198.6000 574.0500 215.4000 ;
	    RECT 573.0000 197.4000 574.2000 198.6000 ;
	    RECT 573.0000 191.4000 574.2000 192.6000 ;
	    RECT 558.6000 161.4000 559.8000 162.6000 ;
	    RECT 546.6000 155.4000 547.8000 156.6000 ;
	    RECT 551.4000 155.4000 552.6000 156.6000 ;
	    RECT 537.0000 137.4000 538.2000 138.6000 ;
	    RECT 539.4000 126.3000 540.6000 146.7000 ;
	    RECT 541.8000 126.3000 543.0000 146.7000 ;
	    RECT 544.2000 129.3000 545.4000 146.7000 ;
	    RECT 546.6000 143.4000 547.8000 144.6000 ;
	    RECT 546.7500 141.6000 547.6500 143.4000 ;
	    RECT 546.6000 140.4000 547.8000 141.6000 ;
	    RECT 549.0000 129.3000 550.2000 146.7000 ;
	    RECT 551.5500 144.6000 552.4500 155.4000 ;
	    RECT 551.4000 143.4000 552.6000 144.6000 ;
	    RECT 551.5500 120.6000 552.4500 143.4000 ;
	    RECT 553.8000 129.3000 555.0000 146.7000 ;
	    RECT 556.2000 126.3000 557.4000 146.7000 ;
	    RECT 558.6000 126.3000 559.8000 146.7000 ;
	    RECT 561.0000 126.3000 562.2000 146.7000 ;
	    RECT 551.4000 119.4000 552.6000 120.6000 ;
	    RECT 565.8000 80.4000 567.0000 81.6000 ;
	    RECT 532.2000 77.5500 535.6500 78.4500 ;
	    RECT 532.2000 77.4000 533.4000 77.5500 ;
	    RECT 534.7500 72.6000 535.6500 77.5500 ;
	    RECT 537.0000 74.4000 538.2000 75.6000 ;
	    RECT 544.2000 74.4000 545.4000 75.6000 ;
	    RECT 534.6000 71.4000 535.8000 72.6000 ;
	    RECT 537.1500 66.6000 538.0500 74.4000 ;
	    RECT 537.0000 66.4500 538.2000 66.6000 ;
	    RECT 537.0000 65.5500 540.4500 66.4500 ;
	    RECT 537.0000 65.4000 538.2000 65.5500 ;
	    RECT 493.8000 59.4000 495.0000 60.6000 ;
	    RECT 503.4000 59.4000 504.6000 60.6000 ;
	    RECT 493.8000 47.4000 495.0000 48.6000 ;
	    RECT 501.0000 47.4000 502.2000 48.6000 ;
	    RECT 501.1500 45.6000 502.0500 47.4000 ;
	    RECT 498.6000 44.4000 499.8000 45.6000 ;
	    RECT 501.0000 44.4000 502.2000 45.6000 ;
	    RECT 498.7500 42.6000 499.6500 44.4000 ;
	    RECT 503.5500 42.6000 504.4500 59.4000 ;
	    RECT 539.5500 54.6000 540.4500 65.5500 ;
	    RECT 544.3500 60.6000 545.2500 74.4000 ;
	    RECT 565.9500 66.6000 566.8500 80.4000 ;
	    RECT 573.1500 78.6000 574.0500 191.4000 ;
	    RECT 575.5500 186.6000 576.4500 218.4000 ;
	    RECT 577.9500 198.6000 578.8500 317.4000 ;
	    RECT 577.8000 197.4000 579.0000 198.6000 ;
	    RECT 577.8000 194.4000 579.0000 195.6000 ;
	    RECT 577.9500 186.6000 578.8500 194.4000 ;
	    RECT 580.3500 192.6000 581.2500 338.5500 ;
	    RECT 582.7500 318.6000 583.6500 491.4000 ;
	    RECT 585.0000 401.4000 586.2000 402.6000 ;
	    RECT 585.1500 378.6000 586.0500 401.4000 ;
	    RECT 585.0000 377.4000 586.2000 378.6000 ;
	    RECT 589.9500 336.6000 590.8500 575.4000 ;
	    RECT 594.7500 519.6000 595.6500 686.5500 ;
	    RECT 597.1500 678.6000 598.0500 755.4000 ;
	    RECT 599.4000 716.4000 600.6000 717.6000 ;
	    RECT 599.5500 708.6000 600.4500 716.4000 ;
	    RECT 601.9500 708.6000 602.8500 758.4000 ;
	    RECT 604.2000 756.3000 605.4000 773.7000 ;
	    RECT 606.6000 756.3000 607.8000 776.7000 ;
	    RECT 609.0000 756.3000 610.2000 776.7000 ;
	    RECT 611.4000 756.3000 612.6000 776.7000 ;
	    RECT 616.3500 750.6000 617.2500 929.4000 ;
	    RECT 621.0000 926.4000 622.2000 927.6000 ;
	    RECT 618.6000 863.4000 619.8000 864.6000 ;
	    RECT 618.7500 828.6000 619.6500 863.4000 ;
	    RECT 618.6000 827.4000 619.8000 828.6000 ;
	    RECT 621.1500 780.6000 622.0500 926.4000 ;
	    RECT 623.4000 887.4000 624.6000 888.6000 ;
	    RECT 621.0000 779.4000 622.2000 780.6000 ;
	    RECT 604.2000 749.4000 605.4000 750.6000 ;
	    RECT 616.2000 749.4000 617.4000 750.6000 ;
	    RECT 599.4000 707.4000 600.6000 708.6000 ;
	    RECT 601.8000 707.4000 603.0000 708.6000 ;
	    RECT 599.5500 696.6000 600.4500 707.4000 ;
	    RECT 604.3500 705.6000 605.2500 749.4000 ;
	    RECT 621.0000 734.4000 622.2000 735.6000 ;
	    RECT 621.1500 732.6000 622.0500 734.4000 ;
	    RECT 621.0000 731.4000 622.2000 732.6000 ;
	    RECT 623.5500 720.6000 624.4500 887.4000 ;
	    RECT 633.1500 885.6000 634.0500 986.4000 ;
	    RECT 635.5500 984.6000 636.4500 995.4000 ;
	    RECT 635.4000 983.4000 636.6000 984.6000 ;
	    RECT 637.8000 983.4000 639.0000 984.6000 ;
	    RECT 633.0000 884.4000 634.2000 885.6000 ;
	    RECT 637.9500 882.6000 638.8500 983.4000 ;
	    RECT 640.3500 948.6000 641.2500 1013.4000 ;
	    RECT 642.6000 1001.4000 643.8000 1002.6000 ;
	    RECT 642.6000 978.4500 643.8000 978.6000 ;
	    RECT 645.1500 978.4500 646.0500 1112.5500 ;
	    RECT 652.3500 1101.6000 653.2500 1121.4000 ;
	    RECT 654.6000 1116.3000 655.8000 1133.7001 ;
	    RECT 657.0000 1133.4000 658.2000 1134.6000 ;
	    RECT 657.0000 1127.4000 658.2000 1128.6000 ;
	    RECT 657.1500 1119.6000 658.0500 1127.4000 ;
	    RECT 657.0000 1118.4000 658.2000 1119.6000 ;
	    RECT 659.4000 1116.3000 660.6000 1133.7001 ;
	    RECT 661.8000 1116.3000 663.0000 1136.7001 ;
	    RECT 664.2000 1116.3000 665.4000 1136.7001 ;
	    RECT 666.6000 1116.3000 667.8000 1136.7001 ;
	    RECT 669.0000 1133.4000 670.2000 1134.6000 ;
	    RECT 652.2000 1100.4000 653.4000 1101.6000 ;
	    RECT 669.1500 1086.6000 670.0500 1133.4000 ;
	    RECT 647.4000 1085.4000 648.6000 1086.6000 ;
	    RECT 669.0000 1085.4000 670.2000 1086.6000 ;
	    RECT 642.6000 977.5500 646.0500 978.4500 ;
	    RECT 642.6000 977.4000 643.8000 977.5500 ;
	    RECT 640.2000 947.4000 641.4000 948.6000 ;
	    RECT 642.7500 945.4500 643.6500 977.4000 ;
	    RECT 645.0000 950.4000 646.2000 951.6000 ;
	    RECT 640.3500 944.5500 643.6500 945.4500 ;
	    RECT 637.8000 881.4000 639.0000 882.6000 ;
	    RECT 625.8000 875.4000 627.0000 876.6000 ;
	    RECT 625.9500 771.6000 626.8500 875.4000 ;
	    RECT 628.2000 827.4000 629.4000 828.6000 ;
	    RECT 628.3500 801.6000 629.2500 827.4000 ;
	    RECT 630.6000 821.4000 631.8000 822.6000 ;
	    RECT 630.7500 816.6000 631.6500 821.4000 ;
	    RECT 630.6000 815.4000 631.8000 816.6000 ;
	    RECT 637.9500 810.6000 638.8500 881.4000 ;
	    RECT 633.0000 809.4000 634.2000 810.6000 ;
	    RECT 637.8000 809.4000 639.0000 810.6000 ;
	    RECT 628.2000 800.4000 629.4000 801.6000 ;
	    RECT 628.3500 798.6000 629.2500 800.4000 ;
	    RECT 628.2000 797.4000 629.4000 798.6000 ;
	    RECT 625.8000 770.4000 627.0000 771.6000 ;
	    RECT 628.3500 738.6000 629.2500 797.4000 ;
	    RECT 628.2000 737.4000 629.4000 738.6000 ;
	    RECT 623.4000 719.4000 624.6000 720.6000 ;
	    RECT 604.2000 704.4000 605.4000 705.6000 ;
	    RECT 604.3500 702.6000 605.2500 704.4000 ;
	    RECT 604.2000 701.4000 605.4000 702.6000 ;
	    RECT 599.4000 695.4000 600.6000 696.6000 ;
	    RECT 606.6000 696.3000 607.8000 716.7000 ;
	    RECT 609.0000 696.3000 610.2000 716.7000 ;
	    RECT 611.4000 696.3000 612.6000 713.7000 ;
	    RECT 613.8000 701.4000 615.0000 702.6000 ;
	    RECT 616.2000 696.3000 617.4000 713.7000 ;
	    RECT 618.6000 707.4000 619.8000 708.6000 ;
	    RECT 618.7500 699.6000 619.6500 707.4000 ;
	    RECT 618.6000 698.4000 619.8000 699.6000 ;
	    RECT 621.0000 696.3000 622.2000 713.7000 ;
	    RECT 623.4000 696.3000 624.6000 716.7000 ;
	    RECT 625.8000 696.3000 627.0000 716.7000 ;
	    RECT 628.2000 696.3000 629.4000 716.7000 ;
	    RECT 609.0000 690.4500 610.2000 690.6000 ;
	    RECT 609.0000 689.5500 612.4500 690.4500 ;
	    RECT 609.0000 689.4000 610.2000 689.5500 ;
	    RECT 597.0000 677.4000 598.2000 678.6000 ;
	    RECT 599.4000 666.3000 600.6000 686.7000 ;
	    RECT 601.8000 666.3000 603.0000 686.7000 ;
	    RECT 604.2000 669.3000 605.4000 686.7000 ;
	    RECT 606.6000 683.4000 607.8000 684.6000 ;
	    RECT 606.7500 681.6000 607.6500 683.4000 ;
	    RECT 606.6000 680.4000 607.8000 681.6000 ;
	    RECT 609.0000 669.3000 610.2000 686.7000 ;
	    RECT 611.5500 684.6000 612.4500 689.5500 ;
	    RECT 611.4000 683.4000 612.6000 684.6000 ;
	    RECT 611.4000 671.4000 612.6000 672.6000 ;
	    RECT 601.8000 660.4500 603.0000 660.6000 ;
	    RECT 599.5500 659.5500 603.0000 660.4500 ;
	    RECT 597.0000 653.4000 598.2000 654.6000 ;
	    RECT 597.1500 561.6000 598.0500 653.4000 ;
	    RECT 599.5500 642.6000 600.4500 659.5500 ;
	    RECT 601.8000 659.4000 603.0000 659.5500 ;
	    RECT 611.5500 654.6000 612.4500 671.4000 ;
	    RECT 613.8000 669.3000 615.0000 686.7000 ;
	    RECT 613.8000 665.4000 615.0000 666.6000 ;
	    RECT 616.2000 666.3000 617.4000 686.7000 ;
	    RECT 618.6000 666.3000 619.8000 686.7000 ;
	    RECT 621.0000 666.3000 622.2000 686.7000 ;
	    RECT 630.6000 677.4000 631.8000 678.6000 ;
	    RECT 613.9500 660.6000 614.8500 665.4000 ;
	    RECT 630.7500 660.6000 631.6500 677.4000 ;
	    RECT 613.8000 659.4000 615.0000 660.6000 ;
	    RECT 630.6000 659.4000 631.8000 660.6000 ;
	    RECT 611.4000 653.4000 612.6000 654.6000 ;
	    RECT 599.4000 641.4000 600.6000 642.6000 ;
	    RECT 628.2000 638.4000 629.4000 639.6000 ;
	    RECT 628.3500 636.6000 629.2500 638.4000 ;
	    RECT 628.2000 635.4000 629.4000 636.6000 ;
	    RECT 618.6000 623.4000 619.8000 624.6000 ;
	    RECT 618.7500 612.6000 619.6500 623.4000 ;
	    RECT 633.1500 621.4500 634.0500 809.4000 ;
	    RECT 637.8000 800.4000 639.0000 801.6000 ;
	    RECT 637.9500 795.6000 638.8500 800.4000 ;
	    RECT 637.8000 794.4000 639.0000 795.6000 ;
	    RECT 635.4000 791.4000 636.6000 792.6000 ;
	    RECT 635.5500 714.6000 636.4500 791.4000 ;
	    RECT 637.9500 738.6000 638.8500 794.4000 ;
	    RECT 640.3500 756.6000 641.2500 944.5500 ;
	    RECT 645.1500 936.6000 646.0500 950.4000 ;
	    RECT 645.0000 935.4000 646.2000 936.6000 ;
	    RECT 645.1500 924.6000 646.0500 935.4000 ;
	    RECT 645.0000 923.4000 646.2000 924.6000 ;
	    RECT 642.6000 893.4000 643.8000 894.6000 ;
	    RECT 642.7500 882.6000 643.6500 893.4000 ;
	    RECT 642.6000 881.4000 643.8000 882.6000 ;
	    RECT 647.5500 861.4500 648.4500 1085.4000 ;
	    RECT 652.2000 1061.4000 653.4000 1062.6000 ;
	    RECT 676.3500 1059.6000 677.2500 1298.4000 ;
	    RECT 688.2000 1283.4000 689.4000 1284.6000 ;
	    RECT 688.3500 1281.6000 689.2500 1283.4000 ;
	    RECT 695.5500 1281.6000 696.4500 1361.4000 ;
	    RECT 719.5500 1356.6000 720.4500 1361.4000 ;
	    RECT 719.4000 1355.4000 720.6000 1356.6000 ;
	    RECT 705.0000 1337.4000 706.2000 1338.6000 ;
	    RECT 700.2000 1334.4000 701.4000 1335.6000 ;
	    RECT 700.3500 1323.6000 701.2500 1334.4000 ;
	    RECT 707.4000 1326.3000 708.6000 1346.7001 ;
	    RECT 709.8000 1326.3000 711.0000 1346.7001 ;
	    RECT 712.2000 1329.3000 713.4000 1346.7001 ;
	    RECT 714.6000 1340.4000 715.8000 1341.6000 ;
	    RECT 700.2000 1322.4000 701.4000 1323.6000 ;
	    RECT 700.3500 1284.6000 701.2500 1322.4000 ;
	    RECT 714.7500 1317.6000 715.6500 1340.4000 ;
	    RECT 717.0000 1329.3000 718.2000 1346.7001 ;
	    RECT 719.4000 1343.4000 720.6000 1344.6000 ;
	    RECT 714.6000 1316.4000 715.8000 1317.6000 ;
	    RECT 719.5500 1305.6000 720.4500 1343.4000 ;
	    RECT 721.8000 1329.3000 723.0000 1346.7001 ;
	    RECT 724.2000 1326.3000 725.4000 1346.7001 ;
	    RECT 726.6000 1326.3000 727.8000 1346.7001 ;
	    RECT 729.0000 1326.3000 730.2000 1346.7001 ;
	    RECT 729.0000 1316.4000 730.2000 1317.6000 ;
	    RECT 702.6000 1304.4000 703.8000 1305.6000 ;
	    RECT 719.4000 1304.4000 720.6000 1305.6000 ;
	    RECT 700.2000 1283.4000 701.4000 1284.6000 ;
	    RECT 700.3500 1281.6000 701.2500 1283.4000 ;
	    RECT 688.2000 1280.4000 689.4000 1281.6000 ;
	    RECT 695.4000 1280.4000 696.6000 1281.6000 ;
	    RECT 700.2000 1280.4000 701.4000 1281.6000 ;
	    RECT 695.4000 1277.4000 696.6000 1278.6000 ;
	    RECT 695.5500 1275.6000 696.4500 1277.4000 ;
	    RECT 695.4000 1274.4000 696.6000 1275.6000 ;
	    RECT 693.0000 1253.4000 694.2000 1254.6000 ;
	    RECT 690.6000 1247.4000 691.8000 1248.6000 ;
	    RECT 690.7500 1218.6000 691.6500 1247.4000 ;
	    RECT 693.1500 1242.6000 694.0500 1253.4000 ;
	    RECT 700.3500 1245.6000 701.2500 1280.4000 ;
	    RECT 697.8000 1244.4000 699.0000 1245.6000 ;
	    RECT 700.2000 1244.4000 701.4000 1245.6000 ;
	    RECT 693.0000 1241.4000 694.2000 1242.6000 ;
	    RECT 697.9500 1221.6000 698.8500 1244.4000 ;
	    RECT 700.3500 1242.6000 701.2500 1244.4000 ;
	    RECT 700.2000 1241.4000 701.4000 1242.6000 ;
	    RECT 697.8000 1220.4000 699.0000 1221.6000 ;
	    RECT 690.6000 1217.4000 691.8000 1218.6000 ;
	    RECT 693.0000 1214.4000 694.2000 1215.6000 ;
	    RECT 693.1500 1206.6000 694.0500 1214.4000 ;
	    RECT 693.0000 1205.4000 694.2000 1206.6000 ;
	    RECT 695.4000 1181.4000 696.6000 1182.6000 ;
	    RECT 683.4000 1145.4000 684.6000 1146.6000 ;
	    RECT 693.0000 1145.4000 694.2000 1146.6000 ;
	    RECT 683.5500 1131.6000 684.4500 1145.4000 ;
	    RECT 683.4000 1130.4000 684.6000 1131.6000 ;
	    RECT 681.0000 1121.4000 682.2000 1122.6000 ;
	    RECT 681.1500 1101.6000 682.0500 1121.4000 ;
	    RECT 683.5500 1104.6000 684.4500 1130.4000 ;
	    RECT 693.1500 1104.6000 694.0500 1145.4000 ;
	    RECT 683.4000 1103.4000 684.6000 1104.6000 ;
	    RECT 693.0000 1103.4000 694.2000 1104.6000 ;
	    RECT 681.0000 1100.4000 682.2000 1101.6000 ;
	    RECT 676.2000 1058.4000 677.4000 1059.6000 ;
	    RECT 652.2000 1055.4000 653.4000 1056.6000 ;
	    RECT 673.8000 1055.4000 675.0000 1056.6000 ;
	    RECT 645.1500 860.5500 648.4500 861.4500 ;
	    RECT 642.6000 833.4000 643.8000 834.6000 ;
	    RECT 642.7500 822.6000 643.6500 833.4000 ;
	    RECT 642.6000 821.4000 643.8000 822.6000 ;
	    RECT 642.7500 798.6000 643.6500 821.4000 ;
	    RECT 642.6000 797.4000 643.8000 798.6000 ;
	    RECT 645.1500 768.6000 646.0500 860.5500 ;
	    RECT 647.4000 857.4000 648.6000 858.6000 ;
	    RECT 647.5500 852.6000 648.4500 857.4000 ;
	    RECT 647.4000 851.4000 648.6000 852.6000 ;
	    RECT 645.0000 767.4000 646.2000 768.6000 ;
	    RECT 645.0000 764.4000 646.2000 765.6000 ;
	    RECT 640.2000 755.4000 641.4000 756.6000 ;
	    RECT 637.8000 737.4000 639.0000 738.6000 ;
	    RECT 645.1500 735.6000 646.0500 764.4000 ;
	    RECT 649.8000 737.4000 651.0000 738.6000 ;
	    RECT 652.3500 735.6000 653.2500 1055.4000 ;
	    RECT 673.9500 1041.6000 674.8500 1055.4000 ;
	    RECT 673.8000 1040.4000 675.0000 1041.6000 ;
	    RECT 657.0000 1037.4000 658.2000 1038.6000 ;
	    RECT 671.4000 1037.4000 672.6000 1038.6000 ;
	    RECT 657.1500 1011.6000 658.0500 1037.4000 ;
	    RECT 659.4000 1019.4000 660.6000 1020.6000 ;
	    RECT 657.0000 1010.4000 658.2000 1011.6000 ;
	    RECT 659.5500 1008.6000 660.4500 1019.4000 ;
	    RECT 673.9500 1008.6000 674.8500 1040.4000 ;
	    RECT 659.4000 1007.4000 660.6000 1008.6000 ;
	    RECT 671.4000 1007.4000 672.6000 1008.6000 ;
	    RECT 673.8000 1007.4000 675.0000 1008.6000 ;
	    RECT 671.5500 1005.4500 672.4500 1007.4000 ;
	    RECT 673.8000 1005.4500 675.0000 1005.6000 ;
	    RECT 671.5500 1004.5500 675.0000 1005.4500 ;
	    RECT 673.8000 1004.4000 675.0000 1004.5500 ;
	    RECT 676.3500 1002.6000 677.2500 1058.4000 ;
	    RECT 678.6000 1043.4000 679.8000 1044.6000 ;
	    RECT 678.6000 1025.4000 679.8000 1026.6000 ;
	    RECT 676.2000 1001.4000 677.4000 1002.6000 ;
	    RECT 676.2000 995.4000 677.4000 996.6000 ;
	    RECT 676.3500 990.6000 677.2500 995.4000 ;
	    RECT 676.2000 989.4000 677.4000 990.6000 ;
	    RECT 661.8000 983.4000 663.0000 984.6000 ;
	    RECT 661.9500 969.4500 662.8500 983.4000 ;
	    RECT 669.0000 977.4000 670.2000 978.6000 ;
	    RECT 664.2000 974.4000 665.4000 975.6000 ;
	    RECT 664.3500 969.4500 665.2500 974.4000 ;
	    RECT 661.9500 968.5500 665.2500 969.4500 ;
	    RECT 664.3500 966.6000 665.2500 968.5500 ;
	    RECT 664.2000 965.4000 665.4000 966.6000 ;
	    RECT 671.4000 966.3000 672.6000 986.7000 ;
	    RECT 673.8000 966.3000 675.0000 986.7000 ;
	    RECT 676.2000 969.3000 677.4000 986.7000 ;
	    RECT 678.7500 981.6000 679.6500 1025.4000 ;
	    RECT 678.6000 980.4000 679.8000 981.6000 ;
	    RECT 681.0000 969.3000 682.2000 986.7000 ;
	    RECT 683.4000 983.4000 684.6000 984.6000 ;
	    RECT 683.5500 966.6000 684.4500 983.4000 ;
	    RECT 685.8000 969.3000 687.0000 986.7000 ;
	    RECT 676.2000 965.4000 677.4000 966.6000 ;
	    RECT 683.4000 965.4000 684.6000 966.6000 ;
	    RECT 688.2000 966.3000 689.4000 986.7000 ;
	    RECT 690.6000 966.3000 691.8000 986.7000 ;
	    RECT 693.0000 966.3000 694.2000 986.7000 ;
	    RECT 676.3500 954.6000 677.2500 965.4000 ;
	    RECT 676.2000 953.4000 677.4000 954.6000 ;
	    RECT 683.4000 953.4000 684.6000 954.6000 ;
	    RECT 681.0000 947.4000 682.2000 948.6000 ;
	    RECT 681.1500 945.6000 682.0500 947.4000 ;
	    RECT 681.0000 944.4000 682.2000 945.6000 ;
	    RECT 683.5500 942.6000 684.4500 953.4000 ;
	    RECT 688.2000 944.4000 689.4000 945.6000 ;
	    RECT 678.6000 941.4000 679.8000 942.6000 ;
	    RECT 683.4000 941.4000 684.6000 942.6000 ;
	    RECT 654.6000 911.4000 655.8000 912.6000 ;
	    RECT 654.7500 879.6000 655.6500 911.4000 ;
	    RECT 678.6000 887.4000 679.8000 888.6000 ;
	    RECT 654.6000 878.4000 655.8000 879.6000 ;
	    RECT 654.7500 876.6000 655.6500 878.4000 ;
	    RECT 654.6000 875.4000 655.8000 876.6000 ;
	    RECT 657.0000 863.4000 658.2000 864.6000 ;
	    RECT 657.1500 858.6000 658.0500 863.4000 ;
	    RECT 657.0000 857.4000 658.2000 858.6000 ;
	    RECT 671.4000 857.4000 672.6000 858.6000 ;
	    RECT 673.8000 857.4000 675.0000 858.6000 ;
	    RECT 671.5500 846.6000 672.4500 857.4000 ;
	    RECT 671.4000 845.4000 672.6000 846.6000 ;
	    RECT 673.9500 825.6000 674.8500 857.4000 ;
	    RECT 678.7500 852.6000 679.6500 887.4000 ;
	    RECT 685.8000 884.4000 687.0000 885.6000 ;
	    RECT 681.0000 881.4000 682.2000 882.6000 ;
	    RECT 683.4000 881.4000 684.6000 882.6000 ;
	    RECT 678.6000 851.4000 679.8000 852.6000 ;
	    RECT 673.8000 824.4000 675.0000 825.6000 ;
	    RECT 681.1500 804.6000 682.0500 881.4000 ;
	    RECT 683.5500 864.6000 684.4500 881.4000 ;
	    RECT 683.4000 863.4000 684.6000 864.6000 ;
	    RECT 678.6000 803.4000 679.8000 804.6000 ;
	    RECT 681.0000 803.4000 682.2000 804.6000 ;
	    RECT 671.4000 797.4000 672.6000 798.6000 ;
	    RECT 678.7500 792.6000 679.6500 803.4000 ;
	    RECT 678.6000 791.4000 679.8000 792.6000 ;
	    RECT 661.8000 767.4000 663.0000 768.6000 ;
	    RECT 661.9500 765.6000 662.8500 767.4000 ;
	    RECT 661.8000 764.4000 663.0000 765.6000 ;
	    RECT 664.2000 764.4000 665.4000 765.6000 ;
	    RECT 664.3500 762.6000 665.2500 764.4000 ;
	    RECT 657.0000 761.4000 658.2000 762.6000 ;
	    RECT 664.2000 761.4000 665.4000 762.6000 ;
	    RECT 661.8000 758.4000 663.0000 759.6000 ;
	    RECT 661.9500 750.6000 662.8500 758.4000 ;
	    RECT 661.8000 749.4000 663.0000 750.6000 ;
	    RECT 673.8000 743.4000 675.0000 744.6000 ;
	    RECT 654.6000 740.4000 655.8000 741.6000 ;
	    RECT 645.0000 734.4000 646.2000 735.6000 ;
	    RECT 652.2000 734.4000 653.4000 735.6000 ;
	    RECT 652.3500 732.6000 653.2500 734.4000 ;
	    RECT 654.7500 732.6000 655.6500 740.4000 ;
	    RECT 652.2000 731.4000 653.4000 732.6000 ;
	    RECT 654.6000 731.4000 655.8000 732.6000 ;
	    RECT 659.4000 731.4000 660.6000 732.6000 ;
	    RECT 635.4000 713.4000 636.6000 714.6000 ;
	    RECT 635.5500 672.6000 636.4500 713.4000 ;
	    RECT 642.6000 710.4000 643.8000 711.6000 ;
	    RECT 637.8000 701.4000 639.0000 702.6000 ;
	    RECT 637.9500 681.6000 638.8500 701.4000 ;
	    RECT 642.7500 684.6000 643.6500 710.4000 ;
	    RECT 647.4000 707.4000 648.6000 708.6000 ;
	    RECT 642.6000 683.4000 643.8000 684.6000 ;
	    RECT 637.8000 680.4000 639.0000 681.6000 ;
	    RECT 642.6000 674.4000 643.8000 675.6000 ;
	    RECT 635.4000 671.4000 636.6000 672.6000 ;
	    RECT 642.7500 648.6000 643.6500 674.4000 ;
	    RECT 647.5500 651.6000 648.4500 707.4000 ;
	    RECT 654.6000 704.4000 655.8000 705.6000 ;
	    RECT 649.8000 689.4000 651.0000 690.6000 ;
	    RECT 647.4000 650.4000 648.6000 651.6000 ;
	    RECT 642.6000 647.4000 643.8000 648.6000 ;
	    RECT 630.7500 620.5500 634.0500 621.4500 ;
	    RECT 628.2000 614.4000 629.4000 615.6000 ;
	    RECT 618.6000 611.4000 619.8000 612.6000 ;
	    RECT 609.0000 596.4000 610.2000 597.6000 ;
	    RECT 599.4000 587.4000 600.6000 588.6000 ;
	    RECT 597.0000 560.4000 598.2000 561.6000 ;
	    RECT 594.6000 518.4000 595.8000 519.6000 ;
	    RECT 599.5500 471.4500 600.4500 587.4000 ;
	    RECT 609.1500 570.6000 610.0500 596.4000 ;
	    RECT 609.0000 569.4000 610.2000 570.6000 ;
	    RECT 618.7500 564.6000 619.6500 611.4000 ;
	    RECT 628.3500 606.6000 629.2500 614.4000 ;
	    RECT 628.2000 605.4000 629.4000 606.6000 ;
	    RECT 628.2000 602.4000 629.4000 603.6000 ;
	    RECT 628.3500 600.6000 629.2500 602.4000 ;
	    RECT 628.2000 599.4000 629.4000 600.6000 ;
	    RECT 630.7500 582.6000 631.6500 620.5500 ;
	    RECT 633.0000 617.4000 634.2000 618.6000 ;
	    RECT 633.1500 588.6000 634.0500 617.4000 ;
	    RECT 635.4000 606.3000 636.6000 626.7000 ;
	    RECT 637.8000 606.3000 639.0000 626.7000 ;
	    RECT 640.2000 609.3000 641.4000 626.7000 ;
	    RECT 642.6000 623.4000 643.8000 624.6000 ;
	    RECT 642.7500 621.6000 643.6500 623.4000 ;
	    RECT 642.6000 620.4000 643.8000 621.6000 ;
	    RECT 645.0000 609.3000 646.2000 626.7000 ;
	    RECT 647.5500 624.6000 648.4500 650.4000 ;
	    RECT 649.9500 642.6000 650.8500 689.4000 ;
	    RECT 652.2000 671.4000 653.4000 672.6000 ;
	    RECT 652.3500 654.6000 653.2500 671.4000 ;
	    RECT 652.2000 653.4000 653.4000 654.6000 ;
	    RECT 654.7500 642.6000 655.6500 704.4000 ;
	    RECT 657.0000 650.4000 658.2000 651.6000 ;
	    RECT 657.1500 648.6000 658.0500 650.4000 ;
	    RECT 659.5500 648.6000 660.4500 731.4000 ;
	    RECT 678.6000 713.4000 679.8000 714.6000 ;
	    RECT 676.2000 707.4000 677.4000 708.6000 ;
	    RECT 676.3500 702.6000 677.2500 707.4000 ;
	    RECT 678.7500 702.6000 679.6500 713.4000 ;
	    RECT 671.4000 701.4000 672.6000 702.6000 ;
	    RECT 676.2000 701.4000 677.4000 702.6000 ;
	    RECT 678.6000 701.4000 679.8000 702.6000 ;
	    RECT 676.2000 680.4000 677.4000 681.6000 ;
	    RECT 673.8000 660.4500 675.0000 660.6000 ;
	    RECT 676.3500 660.4500 677.2500 680.4000 ;
	    RECT 673.8000 659.5500 677.2500 660.4500 ;
	    RECT 673.8000 659.4000 675.0000 659.5500 ;
	    RECT 676.3500 657.6000 677.2500 659.5500 ;
	    RECT 676.2000 656.4000 677.4000 657.6000 ;
	    RECT 661.8000 650.4000 663.0000 651.6000 ;
	    RECT 657.0000 647.4000 658.2000 648.6000 ;
	    RECT 659.4000 647.4000 660.6000 648.6000 ;
	    RECT 659.4000 644.4000 660.6000 645.6000 ;
	    RECT 659.5500 642.6000 660.4500 644.4000 ;
	    RECT 649.8000 641.4000 651.0000 642.6000 ;
	    RECT 654.6000 641.4000 655.8000 642.6000 ;
	    RECT 659.4000 641.4000 660.6000 642.6000 ;
	    RECT 647.4000 623.4000 648.6000 624.6000 ;
	    RECT 647.4000 617.4000 648.6000 618.6000 ;
	    RECT 642.6000 599.4000 643.8000 600.6000 ;
	    RECT 633.0000 587.4000 634.2000 588.6000 ;
	    RECT 630.6000 581.4000 631.8000 582.6000 ;
	    RECT 601.8000 563.4000 603.0000 564.6000 ;
	    RECT 618.6000 563.4000 619.8000 564.6000 ;
	    RECT 601.8000 560.4000 603.0000 561.6000 ;
	    RECT 597.1500 470.5500 600.4500 471.4500 ;
	    RECT 589.8000 335.4000 591.0000 336.6000 ;
	    RECT 582.6000 317.4000 583.8000 318.6000 ;
	    RECT 589.8000 278.4000 591.0000 279.6000 ;
	    RECT 589.9500 261.6000 590.8500 278.4000 ;
	    RECT 589.8000 260.4000 591.0000 261.6000 ;
	    RECT 587.4000 257.4000 588.6000 258.6000 ;
	    RECT 587.5500 252.6000 588.4500 257.4000 ;
	    RECT 587.4000 251.4000 588.6000 252.6000 ;
	    RECT 597.1500 234.6000 598.0500 470.5500 ;
	    RECT 599.4000 467.4000 600.6000 468.6000 ;
	    RECT 599.5500 402.6000 600.4500 467.4000 ;
	    RECT 599.4000 401.4000 600.6000 402.6000 ;
	    RECT 599.5500 384.6000 600.4500 401.4000 ;
	    RECT 599.4000 383.4000 600.6000 384.6000 ;
	    RECT 599.5500 381.6000 600.4500 383.4000 ;
	    RECT 599.4000 380.4000 600.6000 381.6000 ;
	    RECT 601.9500 366.6000 602.8500 560.4000 ;
	    RECT 604.2000 518.4000 605.4000 519.6000 ;
	    RECT 604.3500 474.6000 605.2500 518.4000 ;
	    RECT 616.2000 510.4500 617.4000 510.6000 ;
	    RECT 618.7500 510.4500 619.6500 563.4000 ;
	    RECT 633.1500 561.6000 634.0500 587.4000 ;
	    RECT 642.7500 561.6000 643.6500 599.4000 ;
	    RECT 633.0000 560.4000 634.2000 561.6000 ;
	    RECT 642.6000 560.4000 643.8000 561.6000 ;
	    RECT 616.2000 509.5500 619.6500 510.4500 ;
	    RECT 616.2000 509.4000 617.4000 509.5500 ;
	    RECT 616.3500 504.6000 617.2500 509.4000 ;
	    RECT 616.2000 503.4000 617.4000 504.6000 ;
	    RECT 611.4000 500.4000 612.6000 501.6000 ;
	    RECT 611.5500 498.6000 612.4500 500.4000 ;
	    RECT 611.4000 497.4000 612.6000 498.6000 ;
	    RECT 613.8000 479.4000 615.0000 480.6000 ;
	    RECT 604.2000 473.4000 605.4000 474.6000 ;
	    RECT 604.2000 464.4000 605.4000 465.6000 ;
	    RECT 604.3500 456.6000 605.2500 464.4000 ;
	    RECT 604.2000 455.4000 605.4000 456.6000 ;
	    RECT 606.6000 456.3000 607.8000 476.7000 ;
	    RECT 609.0000 456.3000 610.2000 476.7000 ;
	    RECT 611.4000 456.3000 612.6000 473.7000 ;
	    RECT 613.9500 462.6000 614.8500 479.4000 ;
	    RECT 613.8000 461.4000 615.0000 462.6000 ;
	    RECT 616.2000 456.3000 617.4000 473.7000 ;
	    RECT 618.6000 461.4000 619.8000 462.6000 ;
	    RECT 618.7500 459.6000 619.6500 461.4000 ;
	    RECT 618.6000 458.4000 619.8000 459.6000 ;
	    RECT 621.0000 456.3000 622.2000 473.7000 ;
	    RECT 623.4000 456.3000 624.6000 476.7000 ;
	    RECT 625.8000 456.3000 627.0000 476.7000 ;
	    RECT 628.2000 456.3000 629.4000 476.7000 ;
	    RECT 633.1500 450.6000 634.0500 560.4000 ;
	    RECT 637.8000 554.4000 639.0000 555.6000 ;
	    RECT 637.9500 552.6000 638.8500 554.4000 ;
	    RECT 637.8000 551.4000 639.0000 552.6000 ;
	    RECT 647.5500 516.6000 648.4500 617.4000 ;
	    RECT 649.8000 609.3000 651.0000 626.7000 ;
	    RECT 652.2000 606.3000 653.4000 626.7000 ;
	    RECT 654.6000 606.3000 655.8000 626.7000 ;
	    RECT 657.0000 606.3000 658.2000 626.7000 ;
	    RECT 652.2000 551.4000 653.4000 552.6000 ;
	    RECT 649.8000 524.4000 651.0000 525.6000 ;
	    RECT 649.9500 522.6000 650.8500 524.4000 ;
	    RECT 649.8000 521.4000 651.0000 522.6000 ;
	    RECT 647.4000 515.4000 648.6000 516.6000 ;
	    RECT 647.5500 504.6000 648.4500 515.4000 ;
	    RECT 635.4000 503.4000 636.6000 504.6000 ;
	    RECT 647.4000 503.4000 648.6000 504.6000 ;
	    RECT 635.5500 501.6000 636.4500 503.4000 ;
	    RECT 635.4000 500.4000 636.6000 501.6000 ;
	    RECT 637.8000 500.4000 639.0000 501.6000 ;
	    RECT 635.4000 497.4000 636.6000 498.6000 ;
	    RECT 635.5500 456.6000 636.4500 497.4000 ;
	    RECT 637.9500 492.6000 638.8500 500.4000 ;
	    RECT 637.8000 491.4000 639.0000 492.6000 ;
	    RECT 642.6000 473.4000 643.8000 474.6000 ;
	    RECT 642.7500 471.6000 643.6500 473.4000 ;
	    RECT 642.6000 470.4000 643.8000 471.6000 ;
	    RECT 649.9500 462.6000 650.8500 521.4000 ;
	    RECT 652.3500 519.6000 653.2500 551.4000 ;
	    RECT 652.2000 518.4000 653.4000 519.6000 ;
	    RECT 649.8000 461.4000 651.0000 462.6000 ;
	    RECT 657.0000 458.4000 658.2000 459.6000 ;
	    RECT 635.4000 455.4000 636.6000 456.6000 ;
	    RECT 657.1500 450.6000 658.0500 458.4000 ;
	    RECT 628.2000 449.4000 629.4000 450.6000 ;
	    RECT 633.0000 449.4000 634.2000 450.6000 ;
	    RECT 657.0000 449.4000 658.2000 450.6000 ;
	    RECT 628.3500 438.6000 629.2500 449.4000 ;
	    RECT 628.2000 437.4000 629.4000 438.6000 ;
	    RECT 623.4000 434.4000 624.6000 435.6000 ;
	    RECT 606.6000 425.4000 607.8000 426.6000 ;
	    RECT 606.7500 378.6000 607.6500 425.4000 ;
	    RECT 623.5500 423.6000 624.4500 434.4000 ;
	    RECT 628.2000 431.4000 629.4000 432.6000 ;
	    RECT 623.4000 422.4000 624.6000 423.6000 ;
	    RECT 621.0000 410.4000 622.2000 411.6000 ;
	    RECT 616.2000 407.4000 617.4000 408.6000 ;
	    RECT 616.3500 384.6000 617.2500 407.4000 ;
	    RECT 621.1500 384.6000 622.0500 410.4000 ;
	    RECT 623.5500 402.6000 624.4500 422.4000 ;
	    RECT 628.3500 420.6000 629.2500 431.4000 ;
	    RECT 630.6000 426.3000 631.8000 446.7000 ;
	    RECT 633.0000 426.3000 634.2000 446.7000 ;
	    RECT 635.4000 429.3000 636.6000 446.7000 ;
	    RECT 637.8000 443.4000 639.0000 444.6000 ;
	    RECT 637.9500 441.6000 638.8500 443.4000 ;
	    RECT 637.8000 440.4000 639.0000 441.6000 ;
	    RECT 640.2000 429.3000 641.4000 446.7000 ;
	    RECT 642.6000 443.4000 643.8000 444.6000 ;
	    RECT 642.7500 432.6000 643.6500 443.4000 ;
	    RECT 642.6000 431.4000 643.8000 432.6000 ;
	    RECT 645.0000 429.3000 646.2000 446.7000 ;
	    RECT 647.4000 426.3000 648.6000 446.7000 ;
	    RECT 649.8000 426.3000 651.0000 446.7000 ;
	    RECT 652.2000 426.3000 653.4000 446.7000 ;
	    RECT 628.2000 419.4000 629.4000 420.6000 ;
	    RECT 623.4000 401.4000 624.6000 402.6000 ;
	    RECT 616.2000 383.4000 617.4000 384.6000 ;
	    RECT 621.0000 383.4000 622.2000 384.6000 ;
	    RECT 609.0000 380.4000 610.2000 381.6000 ;
	    RECT 606.6000 377.4000 607.8000 378.6000 ;
	    RECT 604.2000 371.4000 605.4000 372.6000 ;
	    RECT 601.8000 365.4000 603.0000 366.6000 ;
	    RECT 604.3500 351.6000 605.2500 371.4000 ;
	    RECT 604.2000 350.4000 605.4000 351.6000 ;
	    RECT 606.7500 282.6000 607.6500 377.4000 ;
	    RECT 609.1500 321.6000 610.0500 380.4000 ;
	    RECT 609.0000 320.4000 610.2000 321.6000 ;
	    RECT 606.6000 281.4000 607.8000 282.6000 ;
	    RECT 606.7500 276.6000 607.6500 281.4000 ;
	    RECT 616.3500 276.6000 617.2500 383.4000 ;
	    RECT 618.6000 336.3000 619.8000 356.7000 ;
	    RECT 621.0000 336.3000 622.2000 356.7000 ;
	    RECT 623.4000 336.3000 624.6000 356.7000 ;
	    RECT 625.8000 336.3000 627.0000 353.7000 ;
	    RECT 628.3500 339.6000 629.2500 419.4000 ;
	    RECT 659.5500 408.6000 660.4500 641.4000 ;
	    RECT 661.9500 618.6000 662.8500 650.4000 ;
	    RECT 671.4000 635.4000 672.6000 636.6000 ;
	    RECT 661.8000 617.4000 663.0000 618.6000 ;
	    RECT 671.5500 612.6000 672.4500 635.4000 ;
	    RECT 671.4000 611.4000 672.6000 612.6000 ;
	    RECT 676.3500 609.6000 677.2500 656.4000 ;
	    RECT 676.2000 608.4000 677.4000 609.6000 ;
	    RECT 676.2000 575.4000 677.4000 576.6000 ;
	    RECT 676.3500 561.6000 677.2500 575.4000 ;
	    RECT 676.2000 560.4000 677.4000 561.6000 ;
	    RECT 681.1500 501.6000 682.0500 803.4000 ;
	    RECT 683.5500 798.6000 684.4500 863.4000 ;
	    RECT 685.9500 861.6000 686.8500 884.4000 ;
	    RECT 685.8000 860.4000 687.0000 861.6000 ;
	    RECT 688.3500 858.6000 689.2500 944.4000 ;
	    RECT 695.5500 930.6000 696.4500 1181.4000 ;
	    RECT 700.2000 1155.3000 701.4000 1163.7001 ;
	    RECT 702.7500 1161.6000 703.6500 1304.4000 ;
	    RECT 724.2000 1301.4000 725.4000 1302.6000 ;
	    RECT 709.8000 1289.4000 711.0000 1290.6000 ;
	    RECT 705.0000 1196.4000 706.2000 1197.6000 ;
	    RECT 705.1500 1188.6000 706.0500 1196.4000 ;
	    RECT 705.0000 1187.4000 706.2000 1188.6000 ;
	    RECT 709.9500 1185.6000 710.8500 1289.4000 ;
	    RECT 724.3500 1278.6000 725.2500 1301.4000 ;
	    RECT 729.1500 1281.6000 730.0500 1316.4000 ;
	    RECT 731.4000 1313.4000 732.6000 1314.6000 ;
	    RECT 729.0000 1280.4000 730.2000 1281.6000 ;
	    RECT 724.2000 1277.4000 725.4000 1278.6000 ;
	    RECT 729.0000 1277.4000 730.2000 1278.6000 ;
	    RECT 731.5500 1248.6000 732.4500 1313.4000 ;
	    RECT 741.1500 1275.6000 742.0500 1376.4000 ;
	    RECT 748.3500 1374.6000 749.2500 1445.4000 ;
	    RECT 755.4000 1409.4000 756.6000 1410.6000 ;
	    RECT 755.5500 1404.6000 756.4500 1409.4000 ;
	    RECT 755.4000 1403.4000 756.6000 1404.6000 ;
	    RECT 748.2000 1373.4000 749.4000 1374.6000 ;
	    RECT 750.6000 1361.4000 751.8000 1362.6000 ;
	    RECT 750.7500 1344.6000 751.6500 1361.4000 ;
	    RECT 750.6000 1343.4000 751.8000 1344.6000 ;
	    RECT 743.4000 1331.4000 744.6000 1332.6000 ;
	    RECT 743.5500 1320.6000 744.4500 1331.4000 ;
	    RECT 743.4000 1319.4000 744.6000 1320.6000 ;
	    RECT 755.5500 1314.6000 756.4500 1403.4000 ;
	    RECT 755.4000 1313.4000 756.6000 1314.6000 ;
	    RECT 757.9500 1290.6000 758.8500 1451.4000 ;
	    RECT 856.3500 1446.6000 857.2500 1451.4000 ;
	    RECT 856.2000 1445.4000 857.4000 1446.6000 ;
	    RECT 870.6000 1446.3000 871.8000 1466.7001 ;
	    RECT 873.0000 1446.3000 874.2000 1466.7001 ;
	    RECT 875.4000 1446.3000 876.6000 1466.7001 ;
	    RECT 877.8000 1449.3000 879.0000 1466.7001 ;
	    RECT 880.2000 1463.4000 881.4000 1464.6000 ;
	    RECT 834.6000 1436.4000 835.8000 1437.6000 ;
	    RECT 834.7500 1428.6000 835.6500 1436.4000 ;
	    RECT 762.6000 1427.4000 763.8000 1428.6000 ;
	    RECT 834.6000 1427.4000 835.8000 1428.6000 ;
	    RECT 762.7500 1404.6000 763.6500 1427.4000 ;
	    RECT 839.4000 1424.4000 840.6000 1425.6000 ;
	    RECT 762.6000 1403.4000 763.8000 1404.6000 ;
	    RECT 803.4000 1400.4000 804.6000 1401.6000 ;
	    RECT 767.4000 1355.4000 768.6000 1356.6000 ;
	    RECT 765.0000 1313.4000 766.2000 1314.6000 ;
	    RECT 765.1500 1299.6000 766.0500 1313.4000 ;
	    RECT 765.0000 1298.4000 766.2000 1299.6000 ;
	    RECT 757.8000 1289.4000 759.0000 1290.6000 ;
	    RECT 753.0000 1280.4000 754.2000 1281.6000 ;
	    RECT 738.6000 1274.4000 739.8000 1275.6000 ;
	    RECT 741.0000 1274.4000 742.2000 1275.6000 ;
	    RECT 731.4000 1247.4000 732.6000 1248.6000 ;
	    RECT 721.8000 1205.4000 723.0000 1206.6000 ;
	    RECT 721.9500 1200.6000 722.8500 1205.4000 ;
	    RECT 721.8000 1199.4000 723.0000 1200.6000 ;
	    RECT 709.8000 1184.4000 711.0000 1185.6000 ;
	    RECT 709.9500 1182.6000 710.8500 1184.4000 ;
	    RECT 709.8000 1181.4000 711.0000 1182.6000 ;
	    RECT 712.2000 1176.3000 713.4000 1196.7001 ;
	    RECT 714.6000 1176.3000 715.8000 1196.7001 ;
	    RECT 717.0000 1176.3000 718.2000 1193.7001 ;
	    RECT 719.4000 1181.4000 720.6000 1182.6000 ;
	    RECT 719.5500 1173.4501 720.4500 1181.4000 ;
	    RECT 721.8000 1176.3000 723.0000 1193.7001 ;
	    RECT 724.2000 1181.4000 725.4000 1182.6000 ;
	    RECT 724.3500 1179.6000 725.2500 1181.4000 ;
	    RECT 724.2000 1178.4000 725.4000 1179.6000 ;
	    RECT 726.6000 1176.3000 727.8000 1193.7001 ;
	    RECT 729.0000 1176.3000 730.2000 1196.7001 ;
	    RECT 731.4000 1176.3000 732.6000 1196.7001 ;
	    RECT 733.8000 1176.3000 735.0000 1196.7001 ;
	    RECT 719.5500 1172.5500 722.8500 1173.4501 ;
	    RECT 702.6000 1160.4000 703.8000 1161.6000 ;
	    RECT 702.7500 1128.6000 703.6500 1160.4000 ;
	    RECT 705.0000 1149.3000 706.2000 1166.7001 ;
	    RECT 709.8000 1157.4000 711.0000 1158.6000 ;
	    RECT 709.9500 1152.6000 710.8500 1157.4000 ;
	    RECT 709.8000 1151.4000 711.0000 1152.6000 ;
	    RECT 719.4000 1149.3000 720.6000 1166.7001 ;
	    RECT 712.2000 1139.4000 713.4000 1140.6000 ;
	    RECT 702.6000 1127.4000 703.8000 1128.6000 ;
	    RECT 702.7500 1068.6000 703.6500 1127.4000 ;
	    RECT 712.3500 1122.6000 713.2500 1139.4000 ;
	    RECT 717.0000 1124.4000 718.2000 1125.6000 ;
	    RECT 717.1500 1122.6000 718.0500 1124.4000 ;
	    RECT 721.9500 1122.6000 722.8500 1172.5500 ;
	    RECT 726.6000 1127.4000 727.8000 1128.6000 ;
	    RECT 712.2000 1121.4000 713.4000 1122.6000 ;
	    RECT 717.0000 1121.4000 718.2000 1122.6000 ;
	    RECT 721.8000 1121.4000 723.0000 1122.6000 ;
	    RECT 724.2000 1121.4000 725.4000 1122.6000 ;
	    RECT 707.4000 1109.4000 708.6000 1110.6000 ;
	    RECT 707.5500 1101.6000 708.4500 1109.4000 ;
	    RECT 707.4000 1100.4000 708.6000 1101.6000 ;
	    RECT 726.7500 1098.6000 727.6500 1127.4000 ;
	    RECT 726.6000 1097.4000 727.8000 1098.6000 ;
	    RECT 733.8000 1097.4000 735.0000 1098.6000 ;
	    RECT 702.6000 1067.4000 703.8000 1068.6000 ;
	    RECT 733.9500 1056.6000 734.8500 1097.4000 ;
	    RECT 733.8000 1055.4000 735.0000 1056.6000 ;
	    RECT 722.1000 1043.4000 723.3000 1043.7001 ;
	    RECT 722.1000 1042.5000 730.5000 1043.4000 ;
	    RECT 731.4000 1042.5000 732.6000 1043.7001 ;
	    RECT 700.2000 1040.4000 701.4000 1041.6000 ;
	    RECT 700.3500 1038.6000 701.2500 1040.4000 ;
	    RECT 700.2000 1037.4000 701.4000 1038.6000 ;
	    RECT 719.4000 1037.4000 720.6000 1038.6000 ;
	    RECT 714.6000 1031.4000 715.8000 1032.6000 ;
	    RECT 702.6000 1025.4000 703.8000 1026.6000 ;
	    RECT 695.4000 929.4000 696.6000 930.6000 ;
	    RECT 688.2000 857.4000 689.4000 858.6000 ;
	    RECT 693.0000 854.4000 694.2000 855.6000 ;
	    RECT 693.1500 846.6000 694.0500 854.4000 ;
	    RECT 700.2000 851.4000 701.4000 852.6000 ;
	    RECT 693.0000 845.4000 694.2000 846.6000 ;
	    RECT 688.5000 827.7000 689.7000 828.9000 ;
	    RECT 697.8000 827.7000 699.0000 828.9000 ;
	    RECT 685.8000 821.4000 687.0000 822.6000 ;
	    RECT 685.9500 816.6000 686.8500 821.4000 ;
	    RECT 688.5000 820.5000 689.4000 827.7000 ;
	    RECT 690.3000 824.7000 691.5000 825.9000 ;
	    RECT 690.6000 822.6000 691.5000 824.7000 ;
	    RECT 698.1000 822.6000 699.0000 827.7000 ;
	    RECT 700.3500 822.6000 701.2500 851.4000 ;
	    RECT 690.6000 821.7000 699.0000 822.6000 ;
	    RECT 690.6000 820.5000 691.8000 820.8000 ;
	    RECT 695.7000 820.5000 696.9000 820.8000 ;
	    RECT 698.1000 820.5000 699.0000 821.7000 ;
	    RECT 700.2000 821.4000 701.4000 822.6000 ;
	    RECT 688.5000 819.6000 696.9000 820.5000 ;
	    RECT 688.5000 819.3000 689.7000 819.6000 ;
	    RECT 697.8000 819.3000 699.0000 820.5000 ;
	    RECT 685.8000 815.4000 687.0000 816.6000 ;
	    RECT 690.6000 803.4000 691.8000 804.6000 ;
	    RECT 683.4000 797.4000 684.6000 798.6000 ;
	    RECT 702.7500 768.6000 703.6500 1025.4000 ;
	    RECT 709.8000 1007.4000 711.0000 1008.6000 ;
	    RECT 707.4000 995.4000 708.6000 996.6000 ;
	    RECT 707.5500 972.6000 708.4500 995.4000 ;
	    RECT 707.4000 971.4000 708.6000 972.6000 ;
	    RECT 707.5500 960.6000 708.4500 971.4000 ;
	    RECT 707.4000 959.4000 708.6000 960.6000 ;
	    RECT 709.9500 954.6000 710.8500 1007.4000 ;
	    RECT 709.8000 953.4000 711.0000 954.6000 ;
	    RECT 709.9500 945.6000 710.8500 953.4000 ;
	    RECT 712.2000 947.4000 713.4000 948.6000 ;
	    RECT 709.8000 944.4000 711.0000 945.6000 ;
	    RECT 712.3500 942.6000 713.2500 947.4000 ;
	    RECT 712.2000 941.4000 713.4000 942.6000 ;
	    RECT 714.7500 924.6000 715.6500 1031.4000 ;
	    RECT 719.5500 1002.6000 720.4500 1037.4000 ;
	    RECT 722.1000 1035.3000 723.0000 1042.5000 ;
	    RECT 724.2000 1042.2001 725.4000 1042.5000 ;
	    RECT 729.3000 1042.2001 730.5000 1042.5000 ;
	    RECT 731.7000 1041.3000 732.6000 1042.5000 ;
	    RECT 733.9500 1041.6000 734.8500 1055.4000 ;
	    RECT 724.2000 1040.4000 732.6000 1041.3000 ;
	    RECT 733.8000 1040.4000 735.0000 1041.6000 ;
	    RECT 724.2000 1038.3000 725.1000 1040.4000 ;
	    RECT 723.9000 1037.1000 725.1000 1038.3000 ;
	    RECT 731.7000 1035.3000 732.6000 1040.4000 ;
	    RECT 722.1000 1034.1000 723.3000 1035.3000 ;
	    RECT 731.4000 1034.1000 732.6000 1035.3000 ;
	    RECT 723.9000 1007.7000 725.1000 1008.9000 ;
	    RECT 733.8000 1007.7000 735.0000 1008.9000 ;
	    RECT 719.4000 1001.4000 720.6000 1002.6000 ;
	    RECT 723.9000 1000.5000 724.8000 1007.7000 ;
	    RECT 727.8000 1002.6000 729.0000 1002.9000 ;
	    RECT 734.1000 1002.6000 735.0000 1007.7000 ;
	    RECT 736.2000 1007.4000 737.4000 1008.6000 ;
	    RECT 736.3500 1002.6000 737.2500 1007.4000 ;
	    RECT 727.8000 1001.7000 735.0000 1002.6000 ;
	    RECT 726.6000 1000.5000 727.8000 1000.8000 ;
	    RECT 731.7000 1000.5000 732.9000 1000.8000 ;
	    RECT 734.1000 1000.5000 735.0000 1001.7000 ;
	    RECT 736.2000 1001.4000 737.4000 1002.6000 ;
	    RECT 723.9000 999.3000 725.1000 1000.5000 ;
	    RECT 726.6000 999.6000 732.9000 1000.5000 ;
	    RECT 733.8000 999.3000 735.0000 1000.5000 ;
	    RECT 738.7500 978.6000 739.6500 1274.4000 ;
	    RECT 741.1500 1242.6000 742.0500 1274.4000 ;
	    RECT 753.1500 1272.6000 754.0500 1280.4000 ;
	    RECT 753.0000 1271.4000 754.2000 1272.6000 ;
	    RECT 767.5500 1254.6000 768.4500 1355.4000 ;
	    RECT 767.4000 1253.4000 768.6000 1254.6000 ;
	    RECT 777.0000 1253.4000 778.2000 1254.6000 ;
	    RECT 755.4000 1248.4501 756.6000 1248.6000 ;
	    RECT 753.1500 1247.5500 756.6000 1248.4501 ;
	    RECT 745.8000 1244.4000 747.0000 1245.6000 ;
	    RECT 750.6000 1244.4000 751.8000 1245.6000 ;
	    RECT 741.0000 1241.4000 742.2000 1242.6000 ;
	    RECT 745.9500 1188.6000 746.8500 1244.4000 ;
	    RECT 750.7500 1242.6000 751.6500 1244.4000 ;
	    RECT 750.6000 1241.4000 751.8000 1242.6000 ;
	    RECT 748.2000 1199.4000 749.4000 1200.6000 ;
	    RECT 748.3500 1191.6000 749.2500 1199.4000 ;
	    RECT 748.2000 1190.4000 749.4000 1191.6000 ;
	    RECT 745.8000 1187.4000 747.0000 1188.6000 ;
	    RECT 745.8000 1160.4000 747.0000 1161.6000 ;
	    RECT 743.4000 1157.4000 744.6000 1158.6000 ;
	    RECT 743.5500 1152.6000 744.4500 1157.4000 ;
	    RECT 743.4000 1151.4000 744.6000 1152.6000 ;
	    RECT 745.9500 1146.6000 746.8500 1160.4000 ;
	    RECT 745.8000 1145.4000 747.0000 1146.6000 ;
	    RECT 748.3500 1119.6000 749.2500 1190.4000 ;
	    RECT 753.1500 1158.6000 754.0500 1247.5500 ;
	    RECT 755.4000 1247.4000 756.6000 1247.5500 ;
	    RECT 755.4000 1241.4000 756.6000 1242.6000 ;
	    RECT 757.8000 1241.4000 759.0000 1242.6000 ;
	    RECT 755.5500 1236.6000 756.4500 1241.4000 ;
	    RECT 777.1500 1239.6000 778.0500 1253.4000 ;
	    RECT 803.5500 1242.6000 804.4500 1400.4000 ;
	    RECT 825.0000 1370.4000 826.2000 1371.6000 ;
	    RECT 817.8000 1340.4000 819.0000 1341.6000 ;
	    RECT 813.0000 1307.4000 814.2000 1308.6000 ;
	    RECT 810.6000 1304.4000 811.8000 1305.6000 ;
	    RECT 810.7500 1284.6000 811.6500 1304.4000 ;
	    RECT 813.1500 1302.6000 814.0500 1307.4000 ;
	    RECT 817.9500 1302.6000 818.8500 1340.4000 ;
	    RECT 820.2000 1307.4000 821.4000 1308.6000 ;
	    RECT 813.0000 1301.4000 814.2000 1302.6000 ;
	    RECT 817.8000 1301.4000 819.0000 1302.6000 ;
	    RECT 810.6000 1283.4000 811.8000 1284.6000 ;
	    RECT 808.2000 1247.4000 809.4000 1248.6000 ;
	    RECT 805.8000 1244.4000 807.0000 1245.6000 ;
	    RECT 805.9500 1242.6000 806.8500 1244.4000 ;
	    RECT 808.3500 1242.6000 809.2500 1247.4000 ;
	    RECT 803.4000 1241.4000 804.6000 1242.6000 ;
	    RECT 805.8000 1241.4000 807.0000 1242.6000 ;
	    RECT 808.2000 1241.4000 809.4000 1242.6000 ;
	    RECT 777.0000 1238.4000 778.2000 1239.6000 ;
	    RECT 755.4000 1235.4000 756.6000 1236.6000 ;
	    RECT 757.8000 1223.4000 759.0000 1224.6000 ;
	    RECT 753.0000 1157.4000 754.2000 1158.6000 ;
	    RECT 755.4000 1154.4000 756.6000 1155.6000 ;
	    RECT 748.2000 1118.4000 749.4000 1119.6000 ;
	    RECT 748.3500 1110.6000 749.2500 1118.4000 ;
	    RECT 748.2000 1109.4000 749.4000 1110.6000 ;
	    RECT 741.0000 1102.5000 742.2000 1103.7001 ;
	    RECT 750.3000 1103.4000 751.5000 1103.7001 ;
	    RECT 753.0000 1103.4000 754.2000 1104.6000 ;
	    RECT 743.1000 1102.5000 751.5000 1103.4000 ;
	    RECT 741.0000 1101.3000 741.9000 1102.5000 ;
	    RECT 743.1000 1102.2001 744.3000 1102.5000 ;
	    RECT 748.2000 1102.2001 749.4000 1102.5000 ;
	    RECT 741.0000 1100.4000 749.4000 1101.3000 ;
	    RECT 741.0000 1095.3000 741.9000 1100.4000 ;
	    RECT 748.5000 1098.3000 749.4000 1100.4000 ;
	    RECT 748.5000 1097.1000 749.7000 1098.3000 ;
	    RECT 750.6000 1095.3000 751.5000 1102.5000 ;
	    RECT 753.1500 1101.6000 754.0500 1103.4000 ;
	    RECT 753.0000 1100.4000 754.2000 1101.6000 ;
	    RECT 753.0000 1097.4000 754.2000 1098.6000 ;
	    RECT 755.5500 1095.4501 756.4500 1154.4000 ;
	    RECT 757.9500 1128.6000 758.8500 1223.4000 ;
	    RECT 772.2000 1217.4000 773.4000 1218.6000 ;
	    RECT 772.3500 1182.6000 773.2500 1217.4000 ;
	    RECT 774.6000 1187.4000 775.8000 1188.6000 ;
	    RECT 772.2000 1181.4000 773.4000 1182.6000 ;
	    RECT 777.1500 1164.6000 778.0500 1238.4000 ;
	    RECT 810.7500 1227.6000 811.6500 1283.4000 ;
	    RECT 813.0000 1265.4000 814.2000 1266.6000 ;
	    RECT 813.1500 1245.6000 814.0500 1265.4000 ;
	    RECT 813.0000 1244.4000 814.2000 1245.6000 ;
	    RECT 803.4000 1226.4000 804.6000 1227.6000 ;
	    RECT 810.6000 1226.4000 811.8000 1227.6000 ;
	    RECT 781.8000 1181.4000 783.0000 1182.6000 ;
	    RECT 777.0000 1163.4000 778.2000 1164.6000 ;
	    RECT 767.4000 1145.4000 768.6000 1146.6000 ;
	    RECT 767.5500 1140.6000 768.4500 1145.4000 ;
	    RECT 781.9500 1140.6000 782.8500 1181.4000 ;
	    RECT 798.6000 1175.4000 799.8000 1176.6000 ;
	    RECT 798.7500 1158.6000 799.6500 1175.4000 ;
	    RECT 801.0000 1160.4000 802.2000 1161.6000 ;
	    RECT 798.6000 1157.4000 799.8000 1158.6000 ;
	    RECT 767.4000 1139.4000 768.6000 1140.6000 ;
	    RECT 781.8000 1139.4000 783.0000 1140.6000 ;
	    RECT 767.5500 1137.6000 768.4500 1139.4000 ;
	    RECT 767.4000 1136.4000 768.6000 1137.6000 ;
	    RECT 757.8000 1127.4000 759.0000 1128.6000 ;
	    RECT 741.0000 1094.1000 742.2000 1095.3000 ;
	    RECT 750.3000 1094.1000 751.5000 1095.3000 ;
	    RECT 753.1500 1094.5500 756.4500 1095.4501 ;
	    RECT 745.8000 1059.3000 747.0000 1067.7001 ;
	    RECT 748.2000 1067.4000 749.4000 1068.6000 ;
	    RECT 748.3500 1062.6000 749.2500 1067.4000 ;
	    RECT 748.2000 1061.4000 749.4000 1062.6000 ;
	    RECT 745.8000 1055.4000 747.0000 1056.6000 ;
	    RECT 750.6000 1056.3000 751.8000 1073.7001 ;
	    RECT 753.1500 1056.6000 754.0500 1094.5500 ;
	    RECT 755.4000 1064.4000 756.6000 1065.6000 ;
	    RECT 753.0000 1055.4000 754.2000 1056.6000 ;
	    RECT 745.9500 1044.6000 746.8500 1055.4000 ;
	    RECT 745.8000 1043.4000 747.0000 1044.6000 ;
	    RECT 750.6000 1043.4000 751.8000 1044.6000 ;
	    RECT 743.4000 989.4000 744.6000 990.6000 ;
	    RECT 743.5500 981.6000 744.4500 989.4000 ;
	    RECT 745.9500 984.6000 746.8500 1043.4000 ;
	    RECT 748.2000 1037.4000 749.4000 1038.6000 ;
	    RECT 748.3500 1014.6000 749.2500 1037.4000 ;
	    RECT 748.2000 1013.4000 749.4000 1014.6000 ;
	    RECT 748.2000 1004.4000 749.4000 1005.6000 ;
	    RECT 745.8000 983.4000 747.0000 984.6000 ;
	    RECT 743.4000 980.4000 744.6000 981.6000 ;
	    RECT 738.6000 977.4000 739.8000 978.6000 ;
	    RECT 729.0000 974.4000 730.2000 975.6000 ;
	    RECT 724.2000 941.4000 725.4000 942.6000 ;
	    RECT 717.0000 938.4000 718.2000 939.6000 ;
	    RECT 714.6000 923.4000 715.8000 924.6000 ;
	    RECT 717.1500 885.6000 718.0500 938.4000 ;
	    RECT 719.4000 887.4000 720.6000 888.6000 ;
	    RECT 717.0000 884.4000 718.2000 885.6000 ;
	    RECT 707.4000 863.4000 708.6000 864.6000 ;
	    RECT 705.0000 860.4000 706.2000 861.6000 ;
	    RECT 705.1500 840.6000 706.0500 860.4000 ;
	    RECT 707.5500 855.6000 708.4500 863.4000 ;
	    RECT 707.4000 854.4000 708.6000 855.6000 ;
	    RECT 705.0000 839.4000 706.2000 840.6000 ;
	    RECT 705.0000 824.4000 706.2000 825.6000 ;
	    RECT 693.0000 767.4000 694.2000 768.6000 ;
	    RECT 702.6000 767.4000 703.8000 768.6000 ;
	    RECT 688.2000 761.4000 689.4000 762.6000 ;
	    RECT 688.3500 744.6000 689.2500 761.4000 ;
	    RECT 688.2000 743.4000 689.4000 744.6000 ;
	    RECT 685.8000 641.4000 687.0000 642.6000 ;
	    RECT 683.4000 608.4000 684.6000 609.6000 ;
	    RECT 683.5500 561.6000 684.4500 608.4000 ;
	    RECT 683.4000 560.4000 684.6000 561.6000 ;
	    RECT 676.2000 500.4000 677.4000 501.6000 ;
	    RECT 681.0000 500.4000 682.2000 501.6000 ;
	    RECT 666.6000 449.4000 667.8000 450.6000 ;
	    RECT 666.7500 432.6000 667.6500 449.4000 ;
	    RECT 666.6000 431.4000 667.8000 432.6000 ;
	    RECT 676.3500 411.6000 677.2500 500.4000 ;
	    RECT 676.2000 410.4000 677.4000 411.6000 ;
	    RECT 659.4000 407.4000 660.6000 408.6000 ;
	    RECT 681.0000 389.4000 682.2000 390.6000 ;
	    RECT 671.4000 383.4000 672.6000 384.6000 ;
	    RECT 647.4000 380.4000 648.6000 381.6000 ;
	    RECT 647.5500 357.6000 648.4500 380.4000 ;
	    RECT 659.4000 374.4000 660.6000 375.6000 ;
	    RECT 628.2000 338.4000 629.4000 339.6000 ;
	    RECT 606.6000 275.4000 607.8000 276.6000 ;
	    RECT 616.2000 275.4000 617.4000 276.6000 ;
	    RECT 621.0000 275.4000 622.2000 276.6000 ;
	    RECT 616.3500 258.4500 617.2500 275.4000 ;
	    RECT 621.1500 261.6000 622.0500 275.4000 ;
	    RECT 621.0000 260.4000 622.2000 261.6000 ;
	    RECT 618.6000 258.4500 619.8000 258.6000 ;
	    RECT 616.3500 257.5500 619.8000 258.4500 ;
	    RECT 618.6000 257.4000 619.8000 257.5500 ;
	    RECT 601.8000 254.4000 603.0000 255.6000 ;
	    RECT 597.0000 233.4000 598.2000 234.6000 ;
	    RECT 597.1500 216.6000 598.0500 233.4000 ;
	    RECT 601.9500 222.6000 602.8500 254.4000 ;
	    RECT 628.3500 240.6000 629.2500 338.4000 ;
	    RECT 630.6000 336.3000 631.8000 353.7000 ;
	    RECT 633.0000 341.4000 634.2000 342.6000 ;
	    RECT 635.4000 336.3000 636.6000 353.7000 ;
	    RECT 637.8000 336.3000 639.0000 356.7000 ;
	    RECT 640.2000 336.3000 641.4000 356.7000 ;
	    RECT 647.4000 356.4000 648.6000 357.6000 ;
	    RECT 647.5500 354.6000 648.4500 356.4000 ;
	    RECT 647.4000 353.4000 648.6000 354.6000 ;
	    RECT 654.6000 353.4000 655.8000 354.6000 ;
	    RECT 647.5500 348.6000 648.4500 353.4000 ;
	    RECT 642.6000 347.4000 643.8000 348.6000 ;
	    RECT 647.4000 347.4000 648.6000 348.6000 ;
	    RECT 642.7500 345.6000 643.6500 347.4000 ;
	    RECT 642.6000 344.4000 643.8000 345.6000 ;
	    RECT 654.7500 342.6000 655.6500 353.4000 ;
	    RECT 659.5500 345.6000 660.4500 374.4000 ;
	    RECT 671.5500 372.6000 672.4500 383.4000 ;
	    RECT 681.1500 381.6000 682.0500 389.4000 ;
	    RECT 685.9500 381.6000 686.8500 641.4000 ;
	    RECT 688.3500 618.6000 689.2500 743.4000 ;
	    RECT 693.1500 738.6000 694.0500 767.4000 ;
	    RECT 700.2000 758.4000 701.4000 759.6000 ;
	    RECT 700.3500 750.6000 701.2500 758.4000 ;
	    RECT 700.2000 749.4000 701.4000 750.6000 ;
	    RECT 690.6000 737.4000 691.8000 738.6000 ;
	    RECT 693.0000 737.4000 694.2000 738.6000 ;
	    RECT 690.7500 735.6000 691.6500 737.4000 ;
	    RECT 690.6000 734.4000 691.8000 735.6000 ;
	    RECT 690.7500 642.6000 691.6500 734.4000 ;
	    RECT 695.4000 725.4000 696.6000 726.6000 ;
	    RECT 695.5500 705.6000 696.4500 725.4000 ;
	    RECT 695.4000 704.4000 696.6000 705.6000 ;
	    RECT 695.4000 680.4000 696.6000 681.6000 ;
	    RECT 693.0000 677.4000 694.2000 678.6000 ;
	    RECT 695.5500 657.6000 696.4500 680.4000 ;
	    RECT 695.4000 656.4000 696.6000 657.6000 ;
	    RECT 697.8000 653.4000 699.0000 654.6000 ;
	    RECT 697.9500 648.6000 698.8500 653.4000 ;
	    RECT 697.8000 647.4000 699.0000 648.6000 ;
	    RECT 700.3500 642.6000 701.2500 749.4000 ;
	    RECT 705.1500 720.6000 706.0500 824.4000 ;
	    RECT 707.5500 822.6000 708.4500 854.4000 ;
	    RECT 707.4000 821.4000 708.6000 822.6000 ;
	    RECT 709.8000 809.4000 711.0000 810.6000 ;
	    RECT 717.0000 809.4000 718.2000 810.6000 ;
	    RECT 709.9500 801.6000 710.8500 809.4000 ;
	    RECT 709.8000 800.4000 711.0000 801.6000 ;
	    RECT 712.2000 800.4000 713.4000 801.6000 ;
	    RECT 712.3500 759.6000 713.2500 800.4000 ;
	    RECT 717.1500 795.6000 718.0500 809.4000 ;
	    RECT 717.0000 794.4000 718.2000 795.6000 ;
	    RECT 719.5500 768.6000 720.4500 887.4000 ;
	    RECT 724.3500 861.6000 725.2500 941.4000 ;
	    RECT 729.1500 927.6000 730.0500 974.4000 ;
	    RECT 745.9500 966.6000 746.8500 983.4000 ;
	    RECT 745.8000 965.4000 747.0000 966.6000 ;
	    RECT 729.0000 926.4000 730.2000 927.6000 ;
	    RECT 741.0000 926.4000 742.2000 927.6000 ;
	    RECT 738.6000 884.4000 739.8000 885.6000 ;
	    RECT 736.2000 881.4000 737.4000 882.6000 ;
	    RECT 733.8000 878.4000 735.0000 879.6000 ;
	    RECT 726.6000 875.4000 727.8000 876.6000 ;
	    RECT 724.2000 860.4000 725.4000 861.6000 ;
	    RECT 726.7500 825.6000 727.6500 875.4000 ;
	    RECT 729.0000 861.4500 730.2000 861.6000 ;
	    RECT 729.0000 860.5500 732.4500 861.4500 ;
	    RECT 729.0000 860.4000 730.2000 860.5500 ;
	    RECT 731.5500 828.6000 732.4500 860.5500 ;
	    RECT 733.9500 858.6000 734.8500 878.4000 ;
	    RECT 736.3500 870.6000 737.2500 881.4000 ;
	    RECT 736.2000 869.4000 737.4000 870.6000 ;
	    RECT 733.8000 857.4000 735.0000 858.6000 ;
	    RECT 733.8000 854.4000 735.0000 855.6000 ;
	    RECT 731.4000 827.4000 732.6000 828.6000 ;
	    RECT 726.6000 824.4000 727.8000 825.6000 ;
	    RECT 733.9500 816.6000 734.8500 854.4000 ;
	    RECT 736.2000 845.4000 737.4000 846.6000 ;
	    RECT 736.3500 825.6000 737.2500 845.4000 ;
	    RECT 738.7500 834.6000 739.6500 884.4000 ;
	    RECT 741.1500 846.6000 742.0500 926.4000 ;
	    RECT 745.8000 884.4000 747.0000 885.6000 ;
	    RECT 745.9500 876.6000 746.8500 884.4000 ;
	    RECT 745.8000 875.4000 747.0000 876.6000 ;
	    RECT 743.4000 851.4000 744.6000 852.6000 ;
	    RECT 741.0000 845.4000 742.2000 846.6000 ;
	    RECT 738.6000 833.4000 739.8000 834.6000 ;
	    RECT 738.6000 827.4000 739.8000 828.6000 ;
	    RECT 736.2000 824.4000 737.4000 825.6000 ;
	    RECT 738.7500 825.4500 739.6500 827.4000 ;
	    RECT 741.0000 825.4500 742.2000 825.6000 ;
	    RECT 738.7500 824.5500 742.2000 825.4500 ;
	    RECT 733.8000 815.4000 735.0000 816.6000 ;
	    RECT 731.4000 809.4000 732.6000 810.6000 ;
	    RECT 729.0000 803.4000 730.2000 804.6000 ;
	    RECT 729.1500 801.6000 730.0500 803.4000 ;
	    RECT 729.0000 800.4000 730.2000 801.6000 ;
	    RECT 724.2000 779.4000 725.4000 780.6000 ;
	    RECT 719.4000 767.4000 720.6000 768.6000 ;
	    RECT 719.5500 762.6000 720.4500 767.4000 ;
	    RECT 719.4000 761.4000 720.6000 762.6000 ;
	    RECT 712.2000 758.4000 713.4000 759.6000 ;
	    RECT 719.4000 758.4000 720.6000 759.6000 ;
	    RECT 712.2000 743.4000 713.4000 744.6000 ;
	    RECT 712.3500 738.6000 713.2500 743.4000 ;
	    RECT 714.6000 740.4000 715.8000 741.6000 ;
	    RECT 712.2000 737.4000 713.4000 738.6000 ;
	    RECT 714.7500 732.6000 715.6500 740.4000 ;
	    RECT 714.6000 731.4000 715.8000 732.6000 ;
	    RECT 705.0000 719.4000 706.2000 720.6000 ;
	    RECT 714.7500 708.6000 715.6500 731.4000 ;
	    RECT 714.6000 707.4000 715.8000 708.6000 ;
	    RECT 714.7500 699.6000 715.6500 707.4000 ;
	    RECT 709.8000 698.4000 711.0000 699.6000 ;
	    RECT 714.6000 698.4000 715.8000 699.6000 ;
	    RECT 707.4000 683.4000 708.6000 684.6000 ;
	    RECT 702.6000 665.4000 703.8000 666.6000 ;
	    RECT 702.7500 645.6000 703.6500 665.4000 ;
	    RECT 707.4000 653.4000 708.6000 654.6000 ;
	    RECT 707.5500 645.6000 708.4500 653.4000 ;
	    RECT 709.9500 645.6000 710.8500 698.4000 ;
	    RECT 717.0000 695.4000 718.2000 696.6000 ;
	    RECT 717.1500 690.6000 718.0500 695.4000 ;
	    RECT 717.0000 689.4000 718.2000 690.6000 ;
	    RECT 717.0000 677.4000 718.2000 678.6000 ;
	    RECT 717.1500 675.6000 718.0500 677.4000 ;
	    RECT 717.0000 674.4000 718.2000 675.6000 ;
	    RECT 717.0000 665.4000 718.2000 666.6000 ;
	    RECT 717.1500 660.6000 718.0500 665.4000 ;
	    RECT 717.0000 659.4000 718.2000 660.6000 ;
	    RECT 717.0000 653.4000 718.2000 654.6000 ;
	    RECT 714.6000 647.4000 715.8000 648.6000 ;
	    RECT 702.6000 644.4000 703.8000 645.6000 ;
	    RECT 707.4000 644.4000 708.6000 645.6000 ;
	    RECT 709.8000 644.4000 711.0000 645.6000 ;
	    RECT 714.7500 642.6000 715.6500 647.4000 ;
	    RECT 690.6000 641.4000 691.8000 642.6000 ;
	    RECT 695.4000 641.4000 696.6000 642.6000 ;
	    RECT 700.2000 641.4000 701.4000 642.6000 ;
	    RECT 705.0000 641.4000 706.2000 642.6000 ;
	    RECT 712.2000 641.4000 713.4000 642.6000 ;
	    RECT 714.6000 641.4000 715.8000 642.6000 ;
	    RECT 695.5500 624.6000 696.4500 641.4000 ;
	    RECT 695.4000 623.4000 696.6000 624.6000 ;
	    RECT 688.2000 617.4000 689.4000 618.6000 ;
	    RECT 695.5500 612.6000 696.4500 623.4000 ;
	    RECT 712.3500 621.6000 713.2500 641.4000 ;
	    RECT 714.6000 623.4000 715.8000 624.6000 ;
	    RECT 709.8000 620.4000 711.0000 621.6000 ;
	    RECT 712.2000 620.4000 713.4000 621.6000 ;
	    RECT 695.4000 611.4000 696.6000 612.6000 ;
	    RECT 707.4000 605.4000 708.6000 606.6000 ;
	    RECT 707.5500 564.6000 708.4500 605.4000 ;
	    RECT 707.4000 563.4000 708.6000 564.6000 ;
	    RECT 709.9500 558.6000 710.8500 620.4000 ;
	    RECT 714.7500 606.6000 715.6500 623.4000 ;
	    RECT 714.6000 605.4000 715.8000 606.6000 ;
	    RECT 712.2000 599.4000 713.4000 600.6000 ;
	    RECT 712.3500 570.6000 713.2500 599.4000 ;
	    RECT 712.2000 569.4000 713.4000 570.6000 ;
	    RECT 712.2000 563.4000 713.4000 564.6000 ;
	    RECT 709.8000 557.4000 711.0000 558.6000 ;
	    RECT 712.3500 552.6000 713.2500 563.4000 ;
	    RECT 712.2000 551.4000 713.4000 552.6000 ;
	    RECT 695.4000 539.4000 696.6000 540.6000 ;
	    RECT 695.5500 522.6000 696.4500 539.4000 ;
	    RECT 695.4000 521.4000 696.6000 522.6000 ;
	    RECT 712.3500 492.6000 713.2500 551.4000 ;
	    RECT 719.5500 534.6000 720.4500 758.4000 ;
	    RECT 721.8000 737.4000 723.0000 738.6000 ;
	    RECT 721.9500 708.6000 722.8500 737.4000 ;
	    RECT 724.3500 714.6000 725.2500 779.4000 ;
	    RECT 729.0000 719.4000 730.2000 720.6000 ;
	    RECT 724.2000 713.4000 725.4000 714.6000 ;
	    RECT 721.8000 707.4000 723.0000 708.6000 ;
	    RECT 724.2000 695.4000 725.4000 696.6000 ;
	    RECT 724.3500 690.6000 725.2500 695.4000 ;
	    RECT 724.2000 689.4000 725.4000 690.6000 ;
	    RECT 721.8000 653.4000 723.0000 654.6000 ;
	    RECT 721.9500 642.6000 722.8500 653.4000 ;
	    RECT 721.8000 641.4000 723.0000 642.6000 ;
	    RECT 721.8000 629.4000 723.0000 630.6000 ;
	    RECT 721.9500 597.6000 722.8500 629.4000 ;
	    RECT 724.2000 623.4000 725.4000 624.6000 ;
	    RECT 721.8000 596.4000 723.0000 597.6000 ;
	    RECT 724.3500 561.6000 725.2500 623.4000 ;
	    RECT 729.1500 594.6000 730.0500 719.4000 ;
	    RECT 731.5500 684.6000 732.4500 809.4000 ;
	    RECT 733.9500 798.6000 734.8500 815.4000 ;
	    RECT 738.7500 798.6000 739.6500 824.5500 ;
	    RECT 741.0000 824.4000 742.2000 824.5500 ;
	    RECT 741.0000 821.4000 742.2000 822.6000 ;
	    RECT 741.1500 816.6000 742.0500 821.4000 ;
	    RECT 741.0000 815.4000 742.2000 816.6000 ;
	    RECT 733.8000 797.4000 735.0000 798.6000 ;
	    RECT 736.2000 797.4000 737.4000 798.6000 ;
	    RECT 738.6000 797.4000 739.8000 798.6000 ;
	    RECT 736.3500 795.6000 737.2500 797.4000 ;
	    RECT 736.2000 794.4000 737.4000 795.6000 ;
	    RECT 741.0000 794.4000 742.2000 795.6000 ;
	    RECT 741.1500 786.6000 742.0500 794.4000 ;
	    RECT 741.0000 785.4000 742.2000 786.6000 ;
	    RECT 736.2000 767.4000 737.4000 768.6000 ;
	    RECT 738.6000 767.4000 739.8000 768.6000 ;
	    RECT 733.8000 740.4000 735.0000 741.6000 ;
	    RECT 733.9500 738.6000 734.8500 740.4000 ;
	    RECT 733.8000 737.4000 735.0000 738.6000 ;
	    RECT 733.8000 734.4000 735.0000 735.6000 ;
	    RECT 733.9500 711.6000 734.8500 734.4000 ;
	    RECT 733.8000 710.4000 735.0000 711.6000 ;
	    RECT 733.9500 702.6000 734.8500 710.4000 ;
	    RECT 733.8000 701.4000 735.0000 702.6000 ;
	    RECT 731.4000 683.4000 732.6000 684.6000 ;
	    RECT 736.3500 642.6000 737.2500 767.4000 ;
	    RECT 738.7500 708.6000 739.6500 767.4000 ;
	    RECT 741.1500 762.6000 742.0500 785.4000 ;
	    RECT 741.0000 761.4000 742.2000 762.6000 ;
	    RECT 743.5500 741.4500 744.4500 851.4000 ;
	    RECT 748.3500 786.6000 749.2500 1004.4000 ;
	    RECT 750.7500 912.6000 751.6500 1043.4000 ;
	    RECT 755.5500 1026.6000 756.4500 1064.4000 ;
	    RECT 757.9500 1050.6000 758.8500 1127.4000 ;
	    RECT 760.2000 1124.4000 761.4000 1125.6000 ;
	    RECT 757.8000 1049.4000 759.0000 1050.6000 ;
	    RECT 755.4000 1025.4000 756.6000 1026.6000 ;
	    RECT 760.3500 1008.6000 761.2500 1124.4000 ;
	    RECT 767.5500 1122.6000 768.4500 1136.4000 ;
	    RECT 801.1500 1122.6000 802.0500 1160.4000 ;
	    RECT 767.4000 1121.4000 768.6000 1122.6000 ;
	    RECT 781.8000 1121.4000 783.0000 1122.6000 ;
	    RECT 789.0000 1121.4000 790.2000 1122.6000 ;
	    RECT 801.0000 1121.4000 802.2000 1122.6000 ;
	    RECT 781.9500 1119.6000 782.8500 1121.4000 ;
	    RECT 781.8000 1118.4000 783.0000 1119.6000 ;
	    RECT 777.0000 1100.4000 778.2000 1101.6000 ;
	    RECT 767.4000 1094.4000 768.6000 1095.6000 ;
	    RECT 765.0000 1056.3000 766.2000 1073.7001 ;
	    RECT 767.5500 1044.6000 768.4500 1094.4000 ;
	    RECT 774.6000 1080.4501 775.8000 1080.6000 ;
	    RECT 777.1500 1080.4501 778.0500 1100.4000 ;
	    RECT 779.4000 1085.4000 780.6000 1086.6000 ;
	    RECT 774.6000 1079.5500 778.0500 1080.4501 ;
	    RECT 774.6000 1079.4000 775.8000 1079.5500 ;
	    RECT 772.2000 1064.4000 773.4000 1065.6000 ;
	    RECT 767.4000 1043.4000 768.6000 1044.6000 ;
	    RECT 762.6000 1040.4000 763.8000 1041.6000 ;
	    RECT 762.7500 1038.6000 763.6500 1040.4000 ;
	    RECT 762.6000 1037.4000 763.8000 1038.6000 ;
	    RECT 760.2000 1007.4000 761.4000 1008.6000 ;
	    RECT 767.4000 1004.4000 768.6000 1005.6000 ;
	    RECT 762.6000 1001.4000 763.8000 1002.6000 ;
	    RECT 757.8000 995.4000 759.0000 996.6000 ;
	    RECT 753.0000 947.4000 754.2000 948.6000 ;
	    RECT 750.6000 911.4000 751.8000 912.6000 ;
	    RECT 753.1500 864.6000 754.0500 947.4000 ;
	    RECT 755.4000 914.4000 756.6000 915.6000 ;
	    RECT 755.5500 903.6000 756.4500 914.4000 ;
	    RECT 755.4000 902.4000 756.6000 903.6000 ;
	    RECT 755.5500 894.6000 756.4500 902.4000 ;
	    RECT 755.4000 893.4000 756.6000 894.6000 ;
	    RECT 757.9500 882.6000 758.8500 995.4000 ;
	    RECT 762.7500 966.6000 763.6500 1001.4000 ;
	    RECT 767.5500 981.6000 768.4500 1004.4000 ;
	    RECT 767.4000 980.4000 768.6000 981.6000 ;
	    RECT 765.0000 968.4000 766.2000 969.6000 ;
	    RECT 760.2000 965.4000 761.4000 966.6000 ;
	    RECT 762.6000 965.4000 763.8000 966.6000 ;
	    RECT 760.3500 942.6000 761.2500 965.4000 ;
	    RECT 765.1500 942.6000 766.0500 968.4000 ;
	    RECT 769.8000 965.4000 771.0000 966.6000 ;
	    RECT 767.4000 953.4000 768.6000 954.6000 ;
	    RECT 767.5500 948.6000 768.4500 953.4000 ;
	    RECT 767.4000 947.4000 768.6000 948.6000 ;
	    RECT 760.2000 941.4000 761.4000 942.6000 ;
	    RECT 765.0000 941.4000 766.2000 942.6000 ;
	    RECT 760.2000 917.4000 761.4000 918.6000 ;
	    RECT 760.3500 888.6000 761.2500 917.4000 ;
	    RECT 762.6000 906.3000 763.8000 926.7000 ;
	    RECT 765.0000 906.3000 766.2000 926.7000 ;
	    RECT 767.4000 909.3000 768.6000 926.7000 ;
	    RECT 769.9500 921.6000 770.8500 965.4000 ;
	    RECT 772.3500 954.6000 773.2500 1064.4000 ;
	    RECT 779.5500 1041.6000 780.4500 1085.4000 ;
	    RECT 789.1500 1062.6000 790.0500 1121.4000 ;
	    RECT 791.4000 1109.4000 792.6000 1110.6000 ;
	    RECT 791.5500 1104.6000 792.4500 1109.4000 ;
	    RECT 791.4000 1103.4000 792.6000 1104.6000 ;
	    RECT 796.2000 1067.4000 797.4000 1068.6000 ;
	    RECT 793.8000 1064.4000 795.0000 1065.6000 ;
	    RECT 789.0000 1061.4000 790.2000 1062.6000 ;
	    RECT 781.8000 1049.4000 783.0000 1050.6000 ;
	    RECT 781.9500 1044.6000 782.8500 1049.4000 ;
	    RECT 781.8000 1043.4000 783.0000 1044.6000 ;
	    RECT 779.4000 1040.4000 780.6000 1041.6000 ;
	    RECT 793.9500 1032.6000 794.8500 1064.4000 ;
	    RECT 796.3500 1062.6000 797.2500 1067.4000 ;
	    RECT 796.2000 1061.4000 797.4000 1062.6000 ;
	    RECT 793.8000 1031.4000 795.0000 1032.6000 ;
	    RECT 803.5500 1026.6000 804.4500 1226.4000 ;
	    RECT 805.8000 1181.4000 807.0000 1182.6000 ;
	    RECT 805.9500 1161.6000 806.8500 1181.4000 ;
	    RECT 808.2000 1178.4000 809.4000 1179.6000 ;
	    RECT 808.3500 1164.6000 809.2500 1178.4000 ;
	    RECT 813.1500 1176.6000 814.0500 1244.4000 ;
	    RECT 815.4000 1241.4000 816.6000 1242.6000 ;
	    RECT 813.0000 1175.4000 814.2000 1176.6000 ;
	    RECT 808.2000 1163.4000 809.4000 1164.6000 ;
	    RECT 815.5500 1161.6000 816.4500 1241.4000 ;
	    RECT 825.1500 1224.6000 826.0500 1370.4000 ;
	    RECT 839.5500 1344.6000 840.4500 1424.4000 ;
	    RECT 841.8000 1416.3000 843.0000 1436.7001 ;
	    RECT 844.2000 1416.3000 845.4000 1436.7001 ;
	    RECT 846.6000 1416.3000 847.8000 1433.7001 ;
	    RECT 849.0000 1421.4000 850.2000 1422.6000 ;
	    RECT 849.1500 1416.6000 850.0500 1421.4000 ;
	    RECT 849.0000 1415.4000 850.2000 1416.6000 ;
	    RECT 851.4000 1416.3000 852.6000 1433.7001 ;
	    RECT 853.8000 1418.4000 855.0000 1419.6000 ;
	    RECT 853.9500 1416.6000 854.8500 1418.4000 ;
	    RECT 853.8000 1415.4000 855.0000 1416.6000 ;
	    RECT 856.2000 1416.3000 857.4000 1433.7001 ;
	    RECT 858.6000 1416.3000 859.8000 1436.7001 ;
	    RECT 861.0000 1416.3000 862.2000 1436.7001 ;
	    RECT 863.4000 1416.3000 864.6000 1436.7001 ;
	    RECT 877.8000 1430.4000 879.0000 1431.6000 ;
	    RECT 873.0000 1415.4000 874.2000 1416.6000 ;
	    RECT 863.4000 1356.3000 864.6000 1376.7001 ;
	    RECT 865.8000 1356.3000 867.0000 1376.7001 ;
	    RECT 868.2000 1356.3000 869.4000 1376.7001 ;
	    RECT 870.6000 1356.3000 871.8000 1373.7001 ;
	    RECT 873.1500 1359.6000 874.0500 1415.4000 ;
	    RECT 877.9500 1410.6000 878.8500 1430.4000 ;
	    RECT 880.3500 1416.6000 881.2500 1463.4000 ;
	    RECT 882.6000 1449.3000 883.8000 1466.7001 ;
	    RECT 885.0000 1463.4000 886.2000 1464.6000 ;
	    RECT 885.1500 1461.6000 886.0500 1463.4000 ;
	    RECT 885.0000 1460.4000 886.2000 1461.6000 ;
	    RECT 887.4000 1449.3000 888.6000 1466.7001 ;
	    RECT 882.6000 1445.4000 883.8000 1446.6000 ;
	    RECT 889.8000 1446.3000 891.0000 1466.7001 ;
	    RECT 892.2000 1446.3000 893.4000 1466.7001 ;
	    RECT 906.6000 1463.4000 907.8000 1464.6000 ;
	    RECT 906.7500 1461.6000 907.6500 1463.4000 ;
	    RECT 906.6000 1460.4000 907.8000 1461.6000 ;
	    RECT 942.6000 1460.4000 943.8000 1461.6000 ;
	    RECT 894.6000 1457.4000 895.8000 1458.6000 ;
	    RECT 940.2000 1458.4501 941.4000 1458.6000 ;
	    RECT 937.9500 1457.5500 941.4000 1458.4501 ;
	    RECT 894.7500 1452.6000 895.6500 1457.4000 ;
	    RECT 899.4000 1454.4000 900.6000 1455.6000 ;
	    RECT 935.4000 1454.4000 936.6000 1455.6000 ;
	    RECT 894.6000 1451.4000 895.8000 1452.6000 ;
	    RECT 882.7500 1419.6000 883.6500 1445.4000 ;
	    RECT 899.5500 1443.6000 900.4500 1454.4000 ;
	    RECT 899.4000 1442.4000 900.6000 1443.6000 ;
	    RECT 899.5500 1440.6000 900.4500 1442.4000 ;
	    RECT 899.4000 1439.4000 900.6000 1440.6000 ;
	    RECT 906.6000 1439.4000 907.8000 1440.6000 ;
	    RECT 904.2000 1427.4000 905.4000 1428.6000 ;
	    RECT 904.3500 1422.6000 905.2500 1427.4000 ;
	    RECT 906.7500 1422.6000 907.6500 1439.4000 ;
	    RECT 935.5500 1425.6000 936.4500 1454.4000 ;
	    RECT 937.9500 1428.6000 938.8500 1457.5500 ;
	    RECT 940.2000 1457.4000 941.4000 1457.5500 ;
	    RECT 940.2000 1440.4501 941.4000 1440.6000 ;
	    RECT 942.7500 1440.4501 943.6500 1460.4000 ;
	    RECT 1043.4000 1457.4000 1044.6000 1458.6000 ;
	    RECT 945.0000 1451.4000 946.2000 1452.6000 ;
	    RECT 945.1500 1446.6000 946.0500 1451.4000 ;
	    RECT 945.0000 1445.4000 946.2000 1446.6000 ;
	    RECT 940.2000 1439.5500 943.6500 1440.4501 ;
	    RECT 940.2000 1439.4000 941.4000 1439.5500 ;
	    RECT 1031.4000 1430.4000 1032.6000 1431.6000 ;
	    RECT 937.8000 1427.4000 939.0000 1428.6000 ;
	    RECT 966.6000 1427.4000 967.8000 1428.6000 ;
	    RECT 935.4000 1424.4000 936.6000 1425.6000 ;
	    RECT 904.2000 1421.4000 905.4000 1422.6000 ;
	    RECT 906.6000 1421.4000 907.8000 1422.6000 ;
	    RECT 882.6000 1418.4000 883.8000 1419.6000 ;
	    RECT 880.2000 1415.4000 881.4000 1416.6000 ;
	    RECT 877.8000 1409.4000 879.0000 1410.6000 ;
	    RECT 882.7500 1404.6000 883.6500 1418.4000 ;
	    RECT 882.6000 1403.4000 883.8000 1404.6000 ;
	    RECT 904.2000 1397.4000 905.4000 1398.6000 ;
	    RECT 899.4000 1394.4000 900.6000 1395.6000 ;
	    RECT 899.5500 1386.6000 900.4500 1394.4000 ;
	    RECT 899.4000 1385.4000 900.6000 1386.6000 ;
	    RECT 887.4000 1379.4000 888.6000 1380.6000 ;
	    RECT 873.0000 1358.4000 874.2000 1359.6000 ;
	    RECT 873.1500 1344.6000 874.0500 1358.4000 ;
	    RECT 875.4000 1356.3000 876.6000 1373.7001 ;
	    RECT 877.8000 1361.4000 879.0000 1362.6000 ;
	    RECT 877.9500 1356.6000 878.8500 1361.4000 ;
	    RECT 877.8000 1355.4000 879.0000 1356.6000 ;
	    RECT 880.2000 1356.3000 881.4000 1373.7001 ;
	    RECT 882.6000 1356.3000 883.8000 1376.7001 ;
	    RECT 885.0000 1356.3000 886.2000 1376.7001 ;
	    RECT 887.5500 1365.6000 888.4500 1379.4000 ;
	    RECT 892.2000 1376.4000 893.4000 1377.6000 ;
	    RECT 892.3500 1368.6000 893.2500 1376.4000 ;
	    RECT 892.2000 1367.4000 893.4000 1368.6000 ;
	    RECT 887.4000 1364.4000 888.6000 1365.6000 ;
	    RECT 839.4000 1343.4000 840.6000 1344.6000 ;
	    RECT 873.0000 1343.4000 874.2000 1344.6000 ;
	    RECT 880.2000 1343.4000 881.4000 1344.6000 ;
	    RECT 827.4000 1325.4000 828.6000 1326.6000 ;
	    RECT 825.0000 1223.4000 826.2000 1224.6000 ;
	    RECT 827.5500 1188.6000 828.4500 1325.4000 ;
	    RECT 829.8000 1313.4000 831.0000 1314.6000 ;
	    RECT 829.9500 1305.6000 830.8500 1313.4000 ;
	    RECT 832.2000 1307.4000 833.4000 1308.6000 ;
	    RECT 834.6000 1307.4000 835.8000 1308.6000 ;
	    RECT 861.0000 1307.4000 862.2000 1308.6000 ;
	    RECT 829.8000 1304.4000 831.0000 1305.6000 ;
	    RECT 827.4000 1187.4000 828.6000 1188.6000 ;
	    RECT 827.5500 1179.6000 828.4500 1187.4000 ;
	    RECT 827.4000 1178.4000 828.6000 1179.6000 ;
	    RECT 820.2000 1163.4000 821.4000 1164.6000 ;
	    RECT 805.8000 1160.4000 807.0000 1161.6000 ;
	    RECT 815.4000 1160.4000 816.6000 1161.6000 ;
	    RECT 808.2000 1157.4000 809.4000 1158.6000 ;
	    RECT 808.3500 1137.6000 809.2500 1157.4000 ;
	    RECT 808.2000 1136.4000 809.4000 1137.6000 ;
	    RECT 805.8000 1058.4000 807.0000 1059.6000 ;
	    RECT 805.9500 1032.6000 806.8500 1058.4000 ;
	    RECT 808.3500 1041.4501 809.2500 1136.4000 ;
	    RECT 827.4000 1124.4000 828.6000 1125.6000 ;
	    RECT 820.2000 1109.4000 821.4000 1110.6000 ;
	    RECT 820.3500 1101.6000 821.2500 1109.4000 ;
	    RECT 827.5500 1101.6000 828.4500 1124.4000 ;
	    RECT 820.2000 1100.4000 821.4000 1101.6000 ;
	    RECT 822.6000 1100.4000 823.8000 1101.6000 ;
	    RECT 827.4000 1100.4000 828.6000 1101.6000 ;
	    RECT 822.7500 1086.6000 823.6500 1100.4000 ;
	    RECT 825.0000 1097.4000 826.2000 1098.6000 ;
	    RECT 822.6000 1085.4000 823.8000 1086.6000 ;
	    RECT 813.1500 1043.5500 821.2500 1044.4501 ;
	    RECT 808.3500 1040.5500 811.6500 1041.4501 ;
	    RECT 808.2000 1037.4000 809.4000 1038.6000 ;
	    RECT 805.8000 1031.4000 807.0000 1032.6000 ;
	    RECT 803.4000 1025.4000 804.6000 1026.6000 ;
	    RECT 808.2000 1025.4000 809.4000 1026.6000 ;
	    RECT 781.8000 1019.4000 783.0000 1020.6000 ;
	    RECT 781.9500 1002.6000 782.8500 1019.4000 ;
	    RECT 781.8000 1001.4000 783.0000 1002.6000 ;
	    RECT 781.9500 990.6000 782.8500 1001.4000 ;
	    RECT 786.6000 998.4000 787.8000 999.6000 ;
	    RECT 786.7500 996.6000 787.6500 998.4000 ;
	    RECT 786.6000 995.4000 787.8000 996.6000 ;
	    RECT 781.8000 989.4000 783.0000 990.6000 ;
	    RECT 791.7000 983.4000 792.9000 983.7000 ;
	    RECT 791.7000 982.5000 800.1000 983.4000 ;
	    RECT 801.0000 982.5000 802.2000 983.7000 ;
	    RECT 789.0000 980.4000 790.2000 981.6000 ;
	    RECT 786.6000 968.4000 787.8000 969.6000 ;
	    RECT 786.7500 966.6000 787.6500 968.4000 ;
	    RECT 786.6000 965.4000 787.8000 966.6000 ;
	    RECT 772.2000 953.4000 773.4000 954.6000 ;
	    RECT 772.2000 947.4000 773.4000 948.6000 ;
	    RECT 772.3500 942.6000 773.2500 947.4000 ;
	    RECT 786.6000 944.4000 787.8000 945.6000 ;
	    RECT 772.2000 941.4000 773.4000 942.6000 ;
	    RECT 769.8000 920.4000 771.0000 921.6000 ;
	    RECT 772.2000 909.3000 773.4000 926.7000 ;
	    RECT 774.6000 923.4000 775.8000 924.6000 ;
	    RECT 774.6000 911.4000 775.8000 912.6000 ;
	    RECT 765.0000 893.4000 766.2000 894.6000 ;
	    RECT 760.2000 887.4000 761.4000 888.6000 ;
	    RECT 757.8000 881.4000 759.0000 882.6000 ;
	    RECT 753.0000 863.4000 754.2000 864.6000 ;
	    RECT 753.1500 858.6000 754.0500 863.4000 ;
	    RECT 753.0000 857.4000 754.2000 858.6000 ;
	    RECT 757.8000 858.4500 759.0000 858.6000 ;
	    RECT 755.5500 857.5500 759.0000 858.4500 ;
	    RECT 750.6000 845.4000 751.8000 846.6000 ;
	    RECT 750.7500 816.6000 751.6500 845.4000 ;
	    RECT 755.5500 840.6000 756.4500 857.5500 ;
	    RECT 757.8000 857.4000 759.0000 857.5500 ;
	    RECT 755.4000 839.4000 756.6000 840.6000 ;
	    RECT 760.2000 827.4000 761.4000 828.6000 ;
	    RECT 750.6000 815.4000 751.8000 816.6000 ;
	    RECT 760.3500 810.6000 761.2500 827.4000 ;
	    RECT 765.1500 822.6000 766.0500 893.4000 ;
	    RECT 767.4000 887.4000 768.6000 888.6000 ;
	    RECT 767.5500 882.6000 768.4500 887.4000 ;
	    RECT 767.4000 881.4000 768.6000 882.6000 ;
	    RECT 765.0000 821.4000 766.2000 822.6000 ;
	    RECT 760.2000 809.4000 761.4000 810.6000 ;
	    RECT 765.0000 803.4000 766.2000 804.6000 ;
	    RECT 750.6000 797.4000 751.8000 798.6000 ;
	    RECT 757.8000 791.4000 759.0000 792.6000 ;
	    RECT 748.2000 785.4000 749.4000 786.6000 ;
	    RECT 753.0000 785.4000 754.2000 786.6000 ;
	    RECT 750.6000 770.4000 751.8000 771.6000 ;
	    RECT 748.2000 764.4000 749.4000 765.6000 ;
	    RECT 748.3500 756.6000 749.2500 764.4000 ;
	    RECT 748.2000 755.4000 749.4000 756.6000 ;
	    RECT 741.1500 740.5500 744.4500 741.4500 ;
	    RECT 741.1500 726.6000 742.0500 740.5500 ;
	    RECT 748.3500 738.6000 749.2500 755.4000 ;
	    RECT 750.7500 741.6000 751.6500 770.4000 ;
	    RECT 750.6000 740.4000 751.8000 741.6000 ;
	    RECT 743.4000 737.4000 744.6000 738.6000 ;
	    RECT 748.2000 737.4000 749.4000 738.6000 ;
	    RECT 748.2000 734.4000 749.4000 735.6000 ;
	    RECT 745.8000 731.4000 747.0000 732.6000 ;
	    RECT 741.0000 725.4000 742.2000 726.6000 ;
	    RECT 743.4000 719.4000 744.6000 720.6000 ;
	    RECT 743.5500 711.6000 744.4500 719.4000 ;
	    RECT 745.9500 711.6000 746.8500 731.4000 ;
	    RECT 743.4000 710.4000 744.6000 711.6000 ;
	    RECT 745.8000 710.4000 747.0000 711.6000 ;
	    RECT 738.6000 707.4000 739.8000 708.6000 ;
	    RECT 741.0000 707.4000 742.2000 708.6000 ;
	    RECT 741.1500 702.6000 742.0500 707.4000 ;
	    RECT 743.5500 705.6000 744.4500 710.4000 ;
	    RECT 743.4000 704.4000 744.6000 705.6000 ;
	    RECT 741.0000 701.4000 742.2000 702.6000 ;
	    RECT 748.3500 660.6000 749.2500 734.4000 ;
	    RECT 750.7500 732.6000 751.6500 740.4000 ;
	    RECT 750.6000 731.4000 751.8000 732.6000 ;
	    RECT 750.7500 711.6000 751.6500 731.4000 ;
	    RECT 750.6000 710.4000 751.8000 711.6000 ;
	    RECT 748.2000 659.4000 749.4000 660.6000 ;
	    RECT 748.3500 648.6000 749.2500 659.4000 ;
	    RECT 748.2000 647.4000 749.4000 648.6000 ;
	    RECT 736.2000 641.4000 737.4000 642.6000 ;
	    RECT 753.1500 636.6000 754.0500 785.4000 ;
	    RECT 757.9500 654.6000 758.8500 791.4000 ;
	    RECT 765.1500 786.6000 766.0500 803.4000 ;
	    RECT 774.7500 801.6000 775.6500 911.4000 ;
	    RECT 777.0000 909.3000 778.2000 926.7000 ;
	    RECT 779.4000 906.3000 780.6000 926.7000 ;
	    RECT 781.8000 906.3000 783.0000 926.7000 ;
	    RECT 784.2000 906.3000 785.4000 926.7000 ;
	    RECT 786.7500 888.6000 787.6500 944.4000 ;
	    RECT 789.1500 936.6000 790.0500 980.4000 ;
	    RECT 791.7000 975.3000 792.6000 982.5000 ;
	    RECT 793.8000 982.2000 795.0000 982.5000 ;
	    RECT 798.9000 982.2000 800.1000 982.5000 ;
	    RECT 801.3000 981.3000 802.2000 982.5000 ;
	    RECT 793.8000 980.4000 802.2000 981.3000 ;
	    RECT 803.4000 980.4000 804.6000 981.6000 ;
	    RECT 793.8000 978.3000 794.7000 980.4000 ;
	    RECT 793.5000 977.1000 794.7000 978.3000 ;
	    RECT 801.3000 975.3000 802.2000 980.4000 ;
	    RECT 791.7000 974.1000 792.9000 975.3000 ;
	    RECT 801.0000 974.1000 802.2000 975.3000 ;
	    RECT 803.5500 960.6000 804.4500 980.4000 ;
	    RECT 803.4000 959.4000 804.6000 960.6000 ;
	    RECT 793.8000 953.4000 795.0000 954.6000 ;
	    RECT 791.4000 944.4000 792.6000 945.6000 ;
	    RECT 789.0000 935.4000 790.2000 936.6000 ;
	    RECT 786.6000 887.4000 787.8000 888.6000 ;
	    RECT 784.2000 860.4000 785.4000 861.6000 ;
	    RECT 781.8000 845.4000 783.0000 846.6000 ;
	    RECT 781.9500 825.6000 782.8500 845.4000 ;
	    RECT 784.3500 825.6000 785.2500 860.4000 ;
	    RECT 781.8000 824.4000 783.0000 825.6000 ;
	    RECT 784.2000 824.4000 785.4000 825.6000 ;
	    RECT 784.2000 821.4000 785.4000 822.6000 ;
	    RECT 774.6000 800.4000 775.8000 801.6000 ;
	    RECT 784.3500 798.6000 785.2500 821.4000 ;
	    RECT 789.0000 819.4500 790.2000 819.6000 ;
	    RECT 791.5500 819.4500 792.4500 944.4000 ;
	    RECT 789.0000 818.5500 792.4500 819.4500 ;
	    RECT 789.0000 818.4000 790.2000 818.5500 ;
	    RECT 789.1500 816.6000 790.0500 818.4000 ;
	    RECT 789.0000 815.4000 790.2000 816.6000 ;
	    RECT 786.6000 803.4000 787.8000 804.6000 ;
	    RECT 791.4000 803.4000 792.6000 804.6000 ;
	    RECT 784.2000 797.4000 785.4000 798.6000 ;
	    RECT 784.2000 795.4500 785.4000 795.6000 ;
	    RECT 786.7500 795.4500 787.6500 803.4000 ;
	    RECT 791.5500 801.6000 792.4500 803.4000 ;
	    RECT 789.0000 800.4000 790.2000 801.6000 ;
	    RECT 791.4000 800.4000 792.6000 801.6000 ;
	    RECT 784.2000 794.5500 787.6500 795.4500 ;
	    RECT 784.2000 794.4000 785.4000 794.5500 ;
	    RECT 765.0000 785.4000 766.2000 786.6000 ;
	    RECT 786.6000 779.4000 787.8000 780.6000 ;
	    RECT 781.8000 770.4000 783.0000 771.6000 ;
	    RECT 760.2000 767.4000 761.4000 768.6000 ;
	    RECT 765.0000 767.4000 766.2000 768.6000 ;
	    RECT 760.3500 762.6000 761.2500 767.4000 ;
	    RECT 760.2000 761.4000 761.4000 762.6000 ;
	    RECT 760.2000 755.4000 761.4000 756.6000 ;
	    RECT 760.3500 690.6000 761.2500 755.4000 ;
	    RECT 765.1500 744.6000 766.0500 767.4000 ;
	    RECT 769.8000 764.4000 771.0000 765.6000 ;
	    RECT 779.4000 764.4000 780.6000 765.6000 ;
	    RECT 765.0000 743.4000 766.2000 744.6000 ;
	    RECT 762.6000 713.4000 763.8000 714.6000 ;
	    RECT 760.2000 689.4000 761.4000 690.6000 ;
	    RECT 762.7500 678.6000 763.6500 713.4000 ;
	    RECT 765.0000 707.4000 766.2000 708.6000 ;
	    RECT 765.1500 678.6000 766.0500 707.4000 ;
	    RECT 767.4000 683.4000 768.6000 684.6000 ;
	    RECT 767.5500 681.6000 768.4500 683.4000 ;
	    RECT 767.4000 680.4000 768.6000 681.6000 ;
	    RECT 769.9500 678.6000 770.8500 764.4000 ;
	    RECT 774.6000 755.4000 775.8000 756.6000 ;
	    RECT 774.7500 744.6000 775.6500 755.4000 ;
	    RECT 774.6000 743.4000 775.8000 744.6000 ;
	    RECT 774.6000 731.4000 775.8000 732.6000 ;
	    RECT 772.2000 707.4000 773.4000 708.6000 ;
	    RECT 772.3500 696.6000 773.2500 707.4000 ;
	    RECT 774.7500 705.6000 775.6500 731.4000 ;
	    RECT 779.5500 720.6000 780.4500 764.4000 ;
	    RECT 781.9500 756.6000 782.8500 770.4000 ;
	    RECT 784.2000 767.4000 785.4000 768.6000 ;
	    RECT 781.8000 755.4000 783.0000 756.6000 ;
	    RECT 779.4000 719.4000 780.6000 720.6000 ;
	    RECT 781.8000 713.4000 783.0000 714.6000 ;
	    RECT 781.9500 711.6000 782.8500 713.4000 ;
	    RECT 781.8000 710.4000 783.0000 711.6000 ;
	    RECT 784.3500 708.6000 785.2500 767.4000 ;
	    RECT 786.7500 762.6000 787.6500 779.4000 ;
	    RECT 786.6000 761.4000 787.8000 762.6000 ;
	    RECT 786.6000 743.4000 787.8000 744.6000 ;
	    RECT 786.7500 738.6000 787.6500 743.4000 ;
	    RECT 786.6000 737.4000 787.8000 738.6000 ;
	    RECT 784.2000 707.4000 785.4000 708.6000 ;
	    RECT 774.6000 704.4000 775.8000 705.6000 ;
	    RECT 774.7500 702.6000 775.6500 704.4000 ;
	    RECT 774.6000 701.4000 775.8000 702.6000 ;
	    RECT 772.2000 695.4000 773.4000 696.6000 ;
	    RECT 781.8000 683.4000 783.0000 684.6000 ;
	    RECT 772.2000 680.4000 773.4000 681.6000 ;
	    RECT 762.6000 677.4000 763.8000 678.6000 ;
	    RECT 765.0000 677.4000 766.2000 678.6000 ;
	    RECT 769.8000 677.4000 771.0000 678.6000 ;
	    RECT 765.1500 666.6000 766.0500 677.4000 ;
	    RECT 772.3500 672.6000 773.2500 680.4000 ;
	    RECT 772.2000 671.4000 773.4000 672.6000 ;
	    RECT 765.0000 665.4000 766.2000 666.6000 ;
	    RECT 757.8000 653.4000 759.0000 654.6000 ;
	    RECT 762.6000 654.4500 763.8000 654.6000 ;
	    RECT 765.0000 654.4500 766.2000 654.6000 ;
	    RECT 762.6000 653.5500 766.2000 654.4500 ;
	    RECT 762.6000 653.4000 763.8000 653.5500 ;
	    RECT 765.0000 653.4000 766.2000 653.5500 ;
	    RECT 755.4000 644.4000 756.6000 645.6000 ;
	    RECT 760.2000 644.4000 761.4000 645.6000 ;
	    RECT 750.6000 636.4500 751.8000 636.6000 ;
	    RECT 748.3500 635.5500 751.8000 636.4500 ;
	    RECT 748.3500 621.6000 749.2500 635.5500 ;
	    RECT 750.6000 635.4000 751.8000 635.5500 ;
	    RECT 753.0000 635.4000 754.2000 636.6000 ;
	    RECT 755.5500 627.6000 756.4500 644.4000 ;
	    RECT 760.3500 642.6000 761.2500 644.4000 ;
	    RECT 760.2000 641.4000 761.4000 642.6000 ;
	    RECT 779.4000 641.4000 780.6000 642.6000 ;
	    RECT 755.4000 626.4000 756.6000 627.6000 ;
	    RECT 753.0000 623.4000 754.2000 624.6000 ;
	    RECT 753.1500 621.6000 754.0500 623.4000 ;
	    RECT 731.4000 620.4000 732.6000 621.6000 ;
	    RECT 748.2000 620.4000 749.4000 621.6000 ;
	    RECT 753.0000 620.4000 754.2000 621.6000 ;
	    RECT 729.0000 593.4000 730.2000 594.6000 ;
	    RECT 726.6000 587.4000 727.8000 588.6000 ;
	    RECT 726.7500 570.6000 727.6500 587.4000 ;
	    RECT 726.6000 569.4000 727.8000 570.6000 ;
	    RECT 724.2000 560.4000 725.4000 561.6000 ;
	    RECT 719.4000 533.4000 720.6000 534.6000 ;
	    RECT 731.5500 522.6000 732.4500 620.4000 ;
	    RECT 745.8000 617.4000 747.0000 618.6000 ;
	    RECT 745.9500 612.6000 746.8500 617.4000 ;
	    RECT 745.8000 611.4000 747.0000 612.6000 ;
	    RECT 733.8000 587.4000 735.0000 588.6000 ;
	    RECT 733.9500 585.6000 734.8500 587.4000 ;
	    RECT 733.8000 584.4000 735.0000 585.6000 ;
	    RECT 733.9500 564.6000 734.8500 584.4000 ;
	    RECT 736.2000 576.3000 737.4000 596.7000 ;
	    RECT 738.6000 576.3000 739.8000 596.7000 ;
	    RECT 741.0000 576.3000 742.2000 593.7000 ;
	    RECT 743.4000 581.4000 744.6000 582.6000 ;
	    RECT 743.5500 576.6000 744.4500 581.4000 ;
	    RECT 743.4000 575.4000 744.6000 576.6000 ;
	    RECT 745.8000 576.3000 747.0000 593.7000 ;
	    RECT 748.2000 581.4000 749.4000 582.6000 ;
	    RECT 748.3500 579.6000 749.2500 581.4000 ;
	    RECT 748.2000 578.4000 749.4000 579.6000 ;
	    RECT 750.6000 576.3000 751.8000 593.7000 ;
	    RECT 753.0000 576.3000 754.2000 596.7000 ;
	    RECT 755.4000 576.3000 756.6000 596.7000 ;
	    RECT 757.8000 576.3000 759.0000 596.7000 ;
	    RECT 760.3500 582.6000 761.2500 641.4000 ;
	    RECT 762.6000 635.4000 763.8000 636.6000 ;
	    RECT 760.2000 581.4000 761.4000 582.6000 ;
	    RECT 760.3500 576.6000 761.2500 581.4000 ;
	    RECT 760.2000 575.4000 761.4000 576.6000 ;
	    RECT 733.8000 563.4000 735.0000 564.6000 ;
	    RECT 721.8000 521.4000 723.0000 522.6000 ;
	    RECT 724.2000 521.4000 725.4000 522.6000 ;
	    RECT 731.4000 521.4000 732.6000 522.6000 ;
	    RECT 721.9500 504.6000 722.8500 521.4000 ;
	    RECT 714.6000 503.4000 715.8000 504.6000 ;
	    RECT 721.8000 503.4000 723.0000 504.6000 ;
	    RECT 714.7500 492.6000 715.6500 503.4000 ;
	    RECT 712.2000 491.4000 713.4000 492.6000 ;
	    RECT 714.6000 491.4000 715.8000 492.6000 ;
	    RECT 700.2000 485.4000 701.4000 486.6000 ;
	    RECT 700.3500 468.6000 701.2500 485.4000 ;
	    RECT 700.2000 467.4000 701.4000 468.6000 ;
	    RECT 693.0000 461.4000 694.2000 462.6000 ;
	    RECT 700.2000 461.4000 701.4000 462.6000 ;
	    RECT 688.2000 455.4000 689.4000 456.6000 ;
	    RECT 688.3500 420.6000 689.2500 455.4000 ;
	    RECT 693.1500 426.6000 694.0500 461.4000 ;
	    RECT 700.3500 444.6000 701.2500 461.4000 ;
	    RECT 700.2000 443.4000 701.4000 444.6000 ;
	    RECT 700.2000 431.4000 701.4000 432.6000 ;
	    RECT 693.0000 425.4000 694.2000 426.6000 ;
	    RECT 688.2000 419.4000 689.4000 420.6000 ;
	    RECT 690.6000 396.3000 691.8000 416.7000 ;
	    RECT 693.0000 396.3000 694.2000 416.7000 ;
	    RECT 695.4000 396.3000 696.6000 416.7000 ;
	    RECT 697.8000 396.3000 699.0000 413.7000 ;
	    RECT 700.3500 399.6000 701.2500 431.4000 ;
	    RECT 700.2000 398.4000 701.4000 399.6000 ;
	    RECT 700.3500 387.6000 701.2500 398.4000 ;
	    RECT 702.6000 396.3000 703.8000 413.7000 ;
	    RECT 705.0000 401.4000 706.2000 402.6000 ;
	    RECT 705.1500 390.6000 706.0500 401.4000 ;
	    RECT 707.4000 396.3000 708.6000 413.7000 ;
	    RECT 709.8000 396.3000 711.0000 416.7000 ;
	    RECT 712.2000 396.3000 713.4000 416.7000 ;
	    RECT 714.7500 405.6000 715.6500 491.4000 ;
	    RECT 719.4000 464.4000 720.6000 465.6000 ;
	    RECT 724.3500 465.4500 725.2500 521.4000 ;
	    RECT 721.9500 464.5500 725.2500 465.4500 ;
	    RECT 719.5500 450.6000 720.4500 464.4000 ;
	    RECT 719.4000 449.4000 720.6000 450.6000 ;
	    RECT 719.4000 425.4000 720.6000 426.6000 ;
	    RECT 717.0000 419.4000 718.2000 420.6000 ;
	    RECT 714.6000 404.4000 715.8000 405.6000 ;
	    RECT 705.0000 389.4000 706.2000 390.6000 ;
	    RECT 700.2000 386.4000 701.4000 387.6000 ;
	    RECT 681.0000 380.4000 682.2000 381.6000 ;
	    RECT 685.8000 380.4000 687.0000 381.6000 ;
	    RECT 671.4000 371.4000 672.6000 372.6000 ;
	    RECT 714.7500 348.6000 715.6500 404.4000 ;
	    RECT 690.6000 347.4000 691.8000 348.6000 ;
	    RECT 714.6000 347.4000 715.8000 348.6000 ;
	    RECT 659.4000 344.4000 660.6000 345.6000 ;
	    RECT 654.6000 341.4000 655.8000 342.6000 ;
	    RECT 671.4000 335.4000 672.6000 336.6000 ;
	    RECT 664.2000 329.4000 665.4000 330.6000 ;
	    RECT 661.8000 315.3000 663.0000 323.7000 ;
	    RECT 664.3500 321.6000 665.2500 329.4000 ;
	    RECT 664.2000 320.4000 665.4000 321.6000 ;
	    RECT 666.6000 309.3000 667.8000 326.7000 ;
	    RECT 671.5500 318.6000 672.4500 335.4000 ;
	    RECT 671.4000 317.4000 672.6000 318.6000 ;
	    RECT 681.0000 309.3000 682.2000 326.7000 ;
	    RECT 688.2000 317.4000 689.4000 318.6000 ;
	    RECT 688.3500 306.6000 689.2500 317.4000 ;
	    RECT 688.2000 305.4000 689.4000 306.6000 ;
	    RECT 606.6000 239.4000 607.8000 240.6000 ;
	    RECT 628.2000 239.4000 629.4000 240.6000 ;
	    RECT 604.2000 224.4000 605.4000 225.6000 ;
	    RECT 601.8000 221.4000 603.0000 222.6000 ;
	    RECT 604.3500 216.6000 605.2500 224.4000 ;
	    RECT 597.0000 215.4000 598.2000 216.6000 ;
	    RECT 604.2000 215.4000 605.4000 216.6000 ;
	    RECT 597.0000 197.4000 598.2000 198.6000 ;
	    RECT 580.2000 191.4000 581.4000 192.6000 ;
	    RECT 575.4000 185.4000 576.6000 186.6000 ;
	    RECT 577.8000 185.4000 579.0000 186.6000 ;
	    RECT 577.9500 162.6000 578.8500 185.4000 ;
	    RECT 580.2000 164.4000 581.4000 165.6000 ;
	    RECT 577.8000 161.4000 579.0000 162.6000 ;
	    RECT 577.8000 158.4000 579.0000 159.6000 ;
	    RECT 575.4000 155.4000 576.6000 156.6000 ;
	    RECT 575.5500 132.6000 576.4500 155.4000 ;
	    RECT 575.4000 131.4000 576.6000 132.6000 ;
	    RECT 577.9500 111.6000 578.8500 158.4000 ;
	    RECT 580.3500 141.6000 581.2500 164.4000 ;
	    RECT 587.4000 156.3000 588.6000 173.7000 ;
	    RECT 597.1500 165.6000 598.0500 197.4000 ;
	    RECT 604.3500 192.6000 605.2500 215.4000 ;
	    RECT 606.7500 204.6000 607.6500 239.4000 ;
	    RECT 609.0000 227.4000 610.2000 228.6000 ;
	    RECT 633.0000 227.4000 634.2000 228.6000 ;
	    RECT 645.0000 227.4000 646.2000 228.6000 ;
	    RECT 654.6000 227.4000 655.8000 228.6000 ;
	    RECT 609.1500 225.6000 610.0500 227.4000 ;
	    RECT 633.1500 225.6000 634.0500 227.4000 ;
	    RECT 609.0000 224.4000 610.2000 225.6000 ;
	    RECT 633.0000 224.4000 634.2000 225.6000 ;
	    RECT 613.8000 221.4000 615.0000 222.6000 ;
	    RECT 606.6000 203.4000 607.8000 204.6000 ;
	    RECT 606.7500 195.6000 607.6500 203.4000 ;
	    RECT 609.0000 197.4000 610.2000 198.6000 ;
	    RECT 606.6000 194.4000 607.8000 195.6000 ;
	    RECT 604.2000 191.4000 605.4000 192.6000 ;
	    RECT 597.0000 164.4000 598.2000 165.6000 ;
	    RECT 601.8000 156.3000 603.0000 173.7000 ;
	    RECT 604.2000 161.4000 605.4000 162.6000 ;
	    RECT 604.3500 156.6000 605.2500 161.4000 ;
	    RECT 606.6000 159.3000 607.8000 167.7000 ;
	    RECT 609.0000 161.4000 610.2000 162.6000 ;
	    RECT 604.2000 155.4000 605.4000 156.6000 ;
	    RECT 580.2000 140.4000 581.4000 141.6000 ;
	    RECT 609.1500 135.6000 610.0500 161.4000 ;
	    RECT 613.9500 144.6000 614.8500 221.4000 ;
	    RECT 628.2000 215.4000 629.4000 216.6000 ;
	    RECT 628.3500 204.6000 629.2500 215.4000 ;
	    RECT 633.1500 204.6000 634.0500 224.4000 ;
	    RECT 637.8000 221.4000 639.0000 222.6000 ;
	    RECT 645.0000 221.4000 646.2000 222.6000 ;
	    RECT 628.2000 203.4000 629.4000 204.6000 ;
	    RECT 633.0000 203.4000 634.2000 204.6000 ;
	    RECT 637.8000 203.4000 639.0000 204.6000 ;
	    RECT 637.9500 198.6000 638.8500 203.4000 ;
	    RECT 645.1500 198.6000 646.0500 221.4000 ;
	    RECT 649.8000 215.4000 651.0000 216.6000 ;
	    RECT 649.9500 204.6000 650.8500 215.4000 ;
	    RECT 654.7500 204.6000 655.6500 227.4000 ;
	    RECT 685.8000 224.4000 687.0000 225.6000 ;
	    RECT 676.2000 221.4000 677.4000 222.6000 ;
	    RECT 683.4000 221.4000 684.6000 222.6000 ;
	    RECT 649.8000 203.4000 651.0000 204.6000 ;
	    RECT 654.6000 203.4000 655.8000 204.6000 ;
	    RECT 649.8000 200.4000 651.0000 201.6000 ;
	    RECT 637.8000 197.4000 639.0000 198.6000 ;
	    RECT 645.0000 197.4000 646.2000 198.6000 ;
	    RECT 628.2000 194.4000 629.4000 195.6000 ;
	    RECT 625.8000 191.4000 627.0000 192.6000 ;
	    RECT 625.9500 186.6000 626.8500 191.4000 ;
	    RECT 625.8000 185.4000 627.0000 186.6000 ;
	    RECT 625.9500 162.6000 626.8500 185.4000 ;
	    RECT 625.8000 161.4000 627.0000 162.6000 ;
	    RECT 613.8000 143.4000 615.0000 144.6000 ;
	    RECT 625.9500 138.6000 626.8500 161.4000 ;
	    RECT 621.0000 137.4000 622.2000 138.6000 ;
	    RECT 625.8000 137.4000 627.0000 138.6000 ;
	    RECT 609.0000 134.4000 610.2000 135.6000 ;
	    RECT 577.8000 110.4000 579.0000 111.6000 ;
	    RECT 621.1500 108.6000 622.0500 137.4000 ;
	    RECT 621.0000 107.4000 622.2000 108.6000 ;
	    RECT 594.6000 95.4000 595.8000 96.6000 ;
	    RECT 582.6000 83.4000 583.8000 84.6000 ;
	    RECT 573.0000 77.4000 574.2000 78.6000 ;
	    RECT 558.6000 65.4000 559.8000 66.6000 ;
	    RECT 565.8000 65.4000 567.0000 66.6000 ;
	    RECT 544.2000 59.4000 545.4000 60.6000 ;
	    RECT 520.2000 53.4000 521.4000 54.6000 ;
	    RECT 539.4000 53.4000 540.6000 54.6000 ;
	    RECT 520.3500 42.6000 521.2500 53.4000 ;
	    RECT 491.4000 41.4000 492.6000 42.6000 ;
	    RECT 498.6000 41.4000 499.8000 42.6000 ;
	    RECT 503.4000 41.4000 504.6000 42.6000 ;
	    RECT 520.2000 41.4000 521.4000 42.6000 ;
	    RECT 525.0000 41.4000 526.2000 42.6000 ;
	    RECT 544.3500 39.6000 545.2500 59.4000 ;
	    RECT 544.2000 38.4000 545.4000 39.6000 ;
	    RECT 541.8000 35.4000 543.0000 36.6000 ;
	    RECT 489.0000 29.4000 490.2000 30.6000 ;
	    RECT 515.4000 29.4000 516.6000 30.6000 ;
	    RECT 486.6000 23.4000 487.8000 24.6000 ;
	    RECT 395.4000 11.4000 396.6000 12.6000 ;
	    RECT 424.2000 11.4000 425.4000 12.6000 ;
	    RECT 352.2000 5.4000 353.4000 6.6000 ;
	    RECT 505.8000 6.3000 507.0000 26.7000 ;
	    RECT 508.2000 6.3000 509.4000 26.7000 ;
	    RECT 510.6000 6.3000 511.8000 26.7000 ;
	    RECT 513.0000 9.3000 514.2000 26.7000 ;
	    RECT 515.5500 24.6000 516.4500 29.4000 ;
	    RECT 515.4000 23.4000 516.6000 24.6000 ;
	    RECT 517.8000 9.3000 519.0000 26.7000 ;
	    RECT 520.2000 23.4000 521.4000 24.6000 ;
	    RECT 520.3500 21.6000 521.2500 23.4000 ;
	    RECT 520.2000 20.4000 521.4000 21.6000 ;
	    RECT 522.6000 9.3000 523.8000 26.7000 ;
	    RECT 525.0000 6.3000 526.2000 26.7000 ;
	    RECT 527.4000 6.3000 528.6000 26.7000 ;
	    RECT 541.9500 18.6000 542.8500 35.4000 ;
	    RECT 529.8000 17.4000 531.0000 18.6000 ;
	    RECT 541.8000 17.4000 543.0000 18.6000 ;
	    RECT 529.9500 12.6000 530.8500 17.4000 ;
	    RECT 558.7500 15.6000 559.6500 65.4000 ;
	    RECT 563.4000 29.4000 564.6000 30.6000 ;
	    RECT 563.5500 21.6000 564.4500 29.4000 ;
	    RECT 582.7500 24.6000 583.6500 83.4000 ;
	    RECT 594.7500 81.6000 595.6500 95.4000 ;
	    RECT 625.9500 84.6000 626.8500 137.4000 ;
	    RECT 628.3500 132.6000 629.2500 194.4000 ;
	    RECT 649.9500 168.6000 650.8500 200.4000 ;
	    RECT 649.8000 167.4000 651.0000 168.6000 ;
	    RECT 654.7500 165.6000 655.6500 203.4000 ;
	    RECT 654.6000 164.4000 655.8000 165.6000 ;
	    RECT 673.8000 155.4000 675.0000 156.6000 ;
	    RECT 628.2000 131.4000 629.4000 132.6000 ;
	    RECT 664.2000 96.3000 665.4000 116.7000 ;
	    RECT 666.6000 96.3000 667.8000 116.7000 ;
	    RECT 669.0000 96.3000 670.2000 116.7000 ;
	    RECT 671.4000 96.3000 672.6000 113.7000 ;
	    RECT 673.9500 99.6000 674.8500 155.4000 ;
	    RECT 676.3500 138.6000 677.2500 221.4000 ;
	    RECT 683.5500 201.6000 684.4500 221.4000 ;
	    RECT 685.9500 210.6000 686.8500 224.4000 ;
	    RECT 688.2000 218.4000 689.4000 219.6000 ;
	    RECT 685.8000 209.4000 687.0000 210.6000 ;
	    RECT 685.9500 201.6000 686.8500 209.4000 ;
	    RECT 683.4000 200.4000 684.6000 201.6000 ;
	    RECT 685.8000 200.4000 687.0000 201.6000 ;
	    RECT 688.3500 192.6000 689.2500 218.4000 ;
	    RECT 688.2000 191.4000 689.4000 192.6000 ;
	    RECT 676.2000 137.4000 677.4000 138.6000 ;
	    RECT 678.6000 125.4000 679.8000 126.6000 ;
	    RECT 673.8000 98.4000 675.0000 99.6000 ;
	    RECT 676.2000 96.3000 677.4000 113.7000 ;
	    RECT 678.7500 102.6000 679.6500 125.4000 ;
	    RECT 678.6000 101.4000 679.8000 102.6000 ;
	    RECT 681.0000 96.3000 682.2000 113.7000 ;
	    RECT 683.4000 96.3000 684.6000 116.7000 ;
	    RECT 685.8000 96.3000 687.0000 116.7000 ;
	    RECT 688.2000 104.4000 689.4000 105.6000 ;
	    RECT 688.3500 96.6000 689.2500 104.4000 ;
	    RECT 688.2000 95.4000 689.4000 96.6000 ;
	    RECT 597.0000 83.4000 598.2000 84.6000 ;
	    RECT 625.8000 83.4000 627.0000 84.6000 ;
	    RECT 594.6000 80.4000 595.8000 81.6000 ;
	    RECT 625.9500 54.6000 626.8500 83.4000 ;
	    RECT 690.7500 60.6000 691.6500 347.4000 ;
	    RECT 700.2000 329.4000 701.4000 330.6000 ;
	    RECT 697.8000 255.3000 699.0000 263.7000 ;
	    RECT 700.3500 261.6000 701.2500 329.4000 ;
	    RECT 717.1500 324.6000 718.0500 419.4000 ;
	    RECT 719.5500 417.6000 720.4500 425.4000 ;
	    RECT 719.4000 417.4500 720.6000 417.6000 ;
	    RECT 721.9500 417.4500 722.8500 464.5500 ;
	    RECT 719.4000 416.5500 722.8500 417.4500 ;
	    RECT 719.4000 416.4000 720.6000 416.5500 ;
	    RECT 719.5500 408.6000 720.4500 416.4000 ;
	    RECT 733.9500 414.6000 734.8500 563.4000 ;
	    RECT 743.4000 527.4000 744.6000 528.6000 ;
	    RECT 743.5500 519.6000 744.4500 527.4000 ;
	    RECT 743.4000 518.4000 744.6000 519.6000 ;
	    RECT 753.0000 518.4000 754.2000 519.6000 ;
	    RECT 743.5500 510.6000 744.4500 518.4000 ;
	    RECT 743.4000 509.4000 744.6000 510.6000 ;
	    RECT 750.6000 509.4000 751.8000 510.6000 ;
	    RECT 741.0000 464.4000 742.2000 465.6000 ;
	    RECT 738.6000 419.4000 739.8000 420.6000 ;
	    RECT 733.8000 413.4000 735.0000 414.6000 ;
	    RECT 719.4000 407.4000 720.6000 408.6000 ;
	    RECT 738.7500 399.6000 739.6500 419.4000 ;
	    RECT 738.6000 398.4000 739.8000 399.6000 ;
	    RECT 738.6000 390.4500 739.8000 390.6000 ;
	    RECT 741.1500 390.4500 742.0500 464.4000 ;
	    RECT 750.7500 459.6000 751.6500 509.4000 ;
	    RECT 750.6000 458.4000 751.8000 459.6000 ;
	    RECT 745.8000 437.4000 747.0000 438.6000 ;
	    RECT 745.9500 408.6000 746.8500 437.4000 ;
	    RECT 745.8000 407.4000 747.0000 408.6000 ;
	    RECT 738.6000 389.5500 742.0500 390.4500 ;
	    RECT 738.6000 389.4000 739.8000 389.5500 ;
	    RECT 717.0000 323.4000 718.2000 324.6000 ;
	    RECT 721.8000 320.4000 723.0000 321.6000 ;
	    RECT 709.8000 290.4000 711.0000 291.6000 ;
	    RECT 707.4000 284.4000 708.6000 285.6000 ;
	    RECT 700.2000 260.4000 701.4000 261.6000 ;
	    RECT 702.6000 249.3000 703.8000 266.7000 ;
	    RECT 707.5500 258.6000 708.4500 284.4000 ;
	    RECT 709.9500 264.6000 710.8500 290.4000 ;
	    RECT 721.9500 288.6000 722.8500 320.4000 ;
	    RECT 738.7500 318.6000 739.6500 389.4000 ;
	    RECT 750.7500 372.6000 751.6500 458.4000 ;
	    RECT 753.1500 450.6000 754.0500 518.4000 ;
	    RECT 762.7500 474.6000 763.6500 635.4000 ;
	    RECT 777.0000 623.4000 778.2000 624.6000 ;
	    RECT 772.2000 605.4000 773.4000 606.6000 ;
	    RECT 772.3500 591.6000 773.2500 605.4000 ;
	    RECT 772.2000 590.4000 773.4000 591.6000 ;
	    RECT 774.6000 584.4000 775.8000 585.6000 ;
	    RECT 762.6000 473.4000 763.8000 474.6000 ;
	    RECT 753.0000 449.4000 754.2000 450.6000 ;
	    RECT 753.0000 429.3000 754.2000 446.7000 ;
	    RECT 762.6000 443.4000 763.8000 444.6000 ;
	    RECT 762.7500 438.6000 763.6500 443.4000 ;
	    RECT 762.6000 437.4000 763.8000 438.6000 ;
	    RECT 767.4000 429.3000 768.6000 446.7000 ;
	    RECT 774.7500 444.6000 775.6500 584.4000 ;
	    RECT 777.1500 522.6000 778.0500 623.4000 ;
	    RECT 779.5500 621.6000 780.4500 641.4000 ;
	    RECT 781.9500 636.6000 782.8500 683.4000 ;
	    RECT 789.1500 681.6000 790.0500 800.4000 ;
	    RECT 793.9500 798.4500 794.8500 953.4000 ;
	    RECT 796.2000 947.4000 797.4000 948.6000 ;
	    RECT 796.3500 942.6000 797.2500 947.4000 ;
	    RECT 796.2000 941.4000 797.4000 942.6000 ;
	    RECT 798.6000 941.4000 799.8000 942.6000 ;
	    RECT 796.3500 912.6000 797.2500 941.4000 ;
	    RECT 798.7500 912.6000 799.6500 941.4000 ;
	    RECT 808.3500 924.6000 809.2500 1025.4000 ;
	    RECT 808.2000 923.4000 809.4000 924.6000 ;
	    RECT 796.2000 911.4000 797.4000 912.6000 ;
	    RECT 798.6000 911.4000 799.8000 912.6000 ;
	    RECT 798.6000 845.4000 799.8000 846.6000 ;
	    RECT 796.2000 798.4500 797.4000 798.6000 ;
	    RECT 793.9500 797.5500 797.4000 798.4500 ;
	    RECT 796.2000 797.4000 797.4000 797.5500 ;
	    RECT 796.3500 738.6000 797.2500 797.4000 ;
	    RECT 798.7500 759.4500 799.6500 845.4000 ;
	    RECT 808.3500 822.6000 809.2500 923.4000 ;
	    RECT 801.0000 821.4000 802.2000 822.6000 ;
	    RECT 808.2000 821.4000 809.4000 822.6000 ;
	    RECT 801.1500 768.6000 802.0500 821.4000 ;
	    RECT 808.2000 797.4000 809.4000 798.6000 ;
	    RECT 808.3500 792.6000 809.2500 797.4000 ;
	    RECT 808.2000 791.4000 809.4000 792.6000 ;
	    RECT 801.0000 767.4000 802.2000 768.6000 ;
	    RECT 801.1500 762.6000 802.0500 767.4000 ;
	    RECT 803.4000 765.4500 804.6000 765.6000 ;
	    RECT 808.2000 765.4500 809.4000 765.6000 ;
	    RECT 803.4000 764.5500 809.4000 765.4500 ;
	    RECT 803.4000 764.4000 804.6000 764.5500 ;
	    RECT 808.2000 764.4000 809.4000 764.5500 ;
	    RECT 801.0000 761.4000 802.2000 762.6000 ;
	    RECT 798.7500 758.5500 802.0500 759.4500 ;
	    RECT 796.2000 737.4000 797.4000 738.6000 ;
	    RECT 791.4000 734.4000 792.6000 735.6000 ;
	    RECT 798.6000 734.4000 799.8000 735.6000 ;
	    RECT 791.5500 714.6000 792.4500 734.4000 ;
	    RECT 798.7500 732.6000 799.6500 734.4000 ;
	    RECT 793.8000 731.4000 795.0000 732.6000 ;
	    RECT 798.6000 731.4000 799.8000 732.6000 ;
	    RECT 793.9500 720.6000 794.8500 731.4000 ;
	    RECT 793.8000 719.4000 795.0000 720.6000 ;
	    RECT 791.4000 713.4000 792.6000 714.6000 ;
	    RECT 798.6000 710.4000 799.8000 711.6000 ;
	    RECT 798.7500 708.6000 799.6500 710.4000 ;
	    RECT 798.6000 707.4000 799.8000 708.6000 ;
	    RECT 801.1500 705.6000 802.0500 758.5500 ;
	    RECT 808.2000 758.4000 809.4000 759.6000 ;
	    RECT 808.3500 750.6000 809.2500 758.4000 ;
	    RECT 808.2000 749.4000 809.4000 750.6000 ;
	    RECT 805.8000 734.4000 807.0000 735.6000 ;
	    RECT 801.0000 704.4000 802.2000 705.6000 ;
	    RECT 798.6000 701.4000 799.8000 702.6000 ;
	    RECT 803.4000 701.4000 804.6000 702.6000 ;
	    RECT 796.2000 683.4000 797.4000 684.6000 ;
	    RECT 789.0000 680.4000 790.2000 681.6000 ;
	    RECT 796.3500 678.6000 797.2500 683.4000 ;
	    RECT 796.2000 677.4000 797.4000 678.6000 ;
	    RECT 784.2000 641.4000 785.4000 642.6000 ;
	    RECT 786.6000 641.4000 787.8000 642.6000 ;
	    RECT 786.7500 639.4500 787.6500 641.4000 ;
	    RECT 784.3500 638.5500 787.6500 639.4500 ;
	    RECT 781.8000 635.4000 783.0000 636.6000 ;
	    RECT 779.4000 620.4000 780.6000 621.6000 ;
	    RECT 779.4000 593.4000 780.6000 594.6000 ;
	    RECT 777.0000 521.4000 778.2000 522.6000 ;
	    RECT 779.5500 456.6000 780.4500 593.4000 ;
	    RECT 781.8000 527.4000 783.0000 528.6000 ;
	    RECT 781.9500 522.6000 782.8500 527.4000 ;
	    RECT 781.8000 521.4000 783.0000 522.6000 ;
	    RECT 779.4000 455.4000 780.6000 456.6000 ;
	    RECT 769.8000 440.4000 771.0000 441.6000 ;
	    RECT 769.9500 438.6000 770.8500 440.4000 ;
	    RECT 769.8000 437.4000 771.0000 438.6000 ;
	    RECT 772.2000 435.3000 773.4000 443.7000 ;
	    RECT 774.6000 443.4000 775.8000 444.6000 ;
	    RECT 774.6000 431.4000 775.8000 432.6000 ;
	    RECT 774.7500 408.6000 775.6500 431.4000 ;
	    RECT 781.9500 426.6000 782.8500 521.4000 ;
	    RECT 784.3500 441.6000 785.2500 638.5500 ;
	    RECT 789.0000 587.4000 790.2000 588.6000 ;
	    RECT 786.6000 581.4000 787.8000 582.6000 ;
	    RECT 786.7500 528.6000 787.6500 581.4000 ;
	    RECT 786.6000 527.4000 787.8000 528.6000 ;
	    RECT 786.7500 522.6000 787.6500 527.4000 ;
	    RECT 786.6000 521.4000 787.8000 522.6000 ;
	    RECT 789.1500 510.4500 790.0500 587.4000 ;
	    RECT 805.9500 582.6000 806.8500 734.4000 ;
	    RECT 810.7500 714.6000 811.6500 1040.5500 ;
	    RECT 813.1500 1038.6000 814.0500 1043.5500 ;
	    RECT 817.8000 1040.4000 819.0000 1041.6000 ;
	    RECT 820.3500 1041.4501 821.2500 1043.5500 ;
	    RECT 822.6000 1041.4501 823.8000 1041.6000 ;
	    RECT 820.3500 1040.5500 823.8000 1041.4501 ;
	    RECT 822.6000 1040.4000 823.8000 1040.5500 ;
	    RECT 813.0000 1037.4000 814.2000 1038.6000 ;
	    RECT 815.4000 1037.4000 816.6000 1038.6000 ;
	    RECT 815.4000 1032.4501 816.6000 1032.6000 ;
	    RECT 817.9500 1032.4501 818.8500 1040.4000 ;
	    RECT 820.2000 1037.4000 821.4000 1038.6000 ;
	    RECT 815.4000 1031.5500 818.8500 1032.4501 ;
	    RECT 815.4000 1031.4000 816.6000 1031.5500 ;
	    RECT 820.3500 1026.6000 821.2500 1037.4000 ;
	    RECT 820.2000 1025.4000 821.4000 1026.6000 ;
	    RECT 825.1500 1008.6000 826.0500 1097.4000 ;
	    RECT 829.9500 1038.6000 830.8500 1304.4000 ;
	    RECT 832.2000 1247.4000 833.4000 1248.6000 ;
	    RECT 832.3500 1239.6000 833.2500 1247.4000 ;
	    RECT 834.7500 1242.6000 835.6500 1307.4000 ;
	    RECT 861.1500 1305.6000 862.0500 1307.4000 ;
	    RECT 839.4000 1304.4000 840.6000 1305.6000 ;
	    RECT 861.0000 1304.4000 862.2000 1305.6000 ;
	    RECT 839.5500 1296.6000 840.4500 1304.4000 ;
	    RECT 865.8000 1298.4000 867.0000 1299.6000 ;
	    RECT 839.4000 1295.4000 840.6000 1296.6000 ;
	    RECT 837.0000 1277.4000 838.2000 1278.6000 ;
	    RECT 865.9500 1278.4501 866.8500 1298.4000 ;
	    RECT 863.5500 1277.5500 866.8500 1278.4501 ;
	    RECT 834.6000 1241.4000 835.8000 1242.6000 ;
	    RECT 832.2000 1238.4000 833.4000 1239.6000 ;
	    RECT 837.1500 1218.6000 838.0500 1277.4000 ;
	    RECT 851.4000 1265.4000 852.6000 1266.6000 ;
	    RECT 837.0000 1217.4000 838.2000 1218.6000 ;
	    RECT 832.2000 1214.4000 833.4000 1215.6000 ;
	    RECT 832.3500 1206.6000 833.2500 1214.4000 ;
	    RECT 832.2000 1205.4000 833.4000 1206.6000 ;
	    RECT 832.2000 1181.4000 833.4000 1182.6000 ;
	    RECT 832.3500 1140.6000 833.2500 1181.4000 ;
	    RECT 832.2000 1139.4000 833.4000 1140.6000 ;
	    RECT 832.2000 1109.4000 833.4000 1110.6000 ;
	    RECT 832.3500 1101.6000 833.2500 1109.4000 ;
	    RECT 832.2000 1100.4000 833.4000 1101.6000 ;
	    RECT 832.2000 1097.4000 833.4000 1098.6000 ;
	    RECT 829.8000 1037.4000 831.0000 1038.6000 ;
	    RECT 827.4000 1013.4000 828.6000 1014.6000 ;
	    RECT 825.0000 1007.4000 826.2000 1008.6000 ;
	    RECT 820.2000 995.4000 821.4000 996.6000 ;
	    RECT 815.4000 983.4000 816.6000 984.6000 ;
	    RECT 815.5500 948.6000 816.4500 983.4000 ;
	    RECT 820.3500 981.6000 821.2500 995.4000 ;
	    RECT 820.2000 980.4000 821.4000 981.6000 ;
	    RECT 822.6000 980.4000 823.8000 981.6000 ;
	    RECT 817.8000 977.4000 819.0000 978.6000 ;
	    RECT 817.8000 959.4000 819.0000 960.6000 ;
	    RECT 822.7500 948.6000 823.6500 980.4000 ;
	    RECT 825.0000 953.4000 826.2000 954.6000 ;
	    RECT 815.4000 947.4000 816.6000 948.6000 ;
	    RECT 822.6000 947.4000 823.8000 948.6000 ;
	    RECT 825.1500 942.6000 826.0500 953.4000 ;
	    RECT 827.5500 942.6000 828.4500 1013.4000 ;
	    RECT 829.8000 947.4000 831.0000 948.6000 ;
	    RECT 825.0000 941.4000 826.2000 942.6000 ;
	    RECT 827.4000 941.4000 828.6000 942.6000 ;
	    RECT 817.8000 887.7000 819.0000 888.9000 ;
	    RECT 827.1000 887.7000 828.3000 888.9000 ;
	    RECT 813.0000 884.4000 814.2000 885.6000 ;
	    RECT 813.1500 849.6000 814.0500 884.4000 ;
	    RECT 817.8000 882.6000 818.7000 887.7000 ;
	    RECT 825.3000 884.7000 826.5000 885.9000 ;
	    RECT 825.3000 882.6000 826.2000 884.7000 ;
	    RECT 815.4000 881.4000 816.6000 882.6000 ;
	    RECT 817.8000 881.7000 826.2000 882.6000 ;
	    RECT 815.5500 864.6000 816.4500 881.4000 ;
	    RECT 817.8000 880.5000 818.7000 881.7000 ;
	    RECT 819.9000 880.5000 821.1000 880.8000 ;
	    RECT 825.0000 880.5000 826.2000 880.8000 ;
	    RECT 827.4000 880.5000 828.3000 887.7000 ;
	    RECT 829.8000 887.4000 831.0000 888.6000 ;
	    RECT 829.9500 882.6000 830.8500 887.4000 ;
	    RECT 829.8000 881.4000 831.0000 882.6000 ;
	    RECT 817.8000 879.3000 819.0000 880.5000 ;
	    RECT 819.9000 879.6000 828.3000 880.5000 ;
	    RECT 827.1000 879.3000 828.3000 879.6000 ;
	    RECT 815.4000 863.4000 816.6000 864.6000 ;
	    RECT 815.4000 851.4000 816.6000 852.6000 ;
	    RECT 813.0000 848.4000 814.2000 849.6000 ;
	    RECT 815.5500 825.4500 816.4500 851.4000 ;
	    RECT 813.1500 824.5500 816.4500 825.4500 ;
	    RECT 810.6000 713.4000 811.8000 714.6000 ;
	    RECT 813.1500 708.6000 814.0500 824.5500 ;
	    RECT 820.2000 824.4000 821.4000 825.6000 ;
	    RECT 825.0000 824.4000 826.2000 825.6000 ;
	    RECT 820.3500 822.6000 821.2500 824.4000 ;
	    RECT 815.4000 821.4000 816.6000 822.6000 ;
	    RECT 817.8000 821.4000 819.0000 822.6000 ;
	    RECT 820.2000 821.4000 821.4000 822.6000 ;
	    RECT 822.6000 821.4000 823.8000 822.6000 ;
	    RECT 815.5500 780.6000 816.4500 821.4000 ;
	    RECT 817.9500 816.6000 818.8500 821.4000 ;
	    RECT 817.8000 815.4000 819.0000 816.6000 ;
	    RECT 822.7500 804.6000 823.6500 821.4000 ;
	    RECT 820.2000 803.4000 821.4000 804.6000 ;
	    RECT 822.6000 803.4000 823.8000 804.6000 ;
	    RECT 815.4000 779.4000 816.6000 780.6000 ;
	    RECT 820.3500 738.6000 821.2500 803.4000 ;
	    RECT 825.1500 768.6000 826.0500 824.4000 ;
	    RECT 827.4000 821.4000 828.6000 822.6000 ;
	    RECT 829.8000 821.4000 831.0000 822.6000 ;
	    RECT 829.9500 816.6000 830.8500 821.4000 ;
	    RECT 829.8000 815.4000 831.0000 816.6000 ;
	    RECT 825.0000 767.4000 826.2000 768.6000 ;
	    RECT 822.6000 765.4500 823.8000 765.6000 ;
	    RECT 827.4000 765.4500 828.6000 765.6000 ;
	    RECT 822.6000 764.5500 828.6000 765.4500 ;
	    RECT 822.6000 764.4000 823.8000 764.5500 ;
	    RECT 827.4000 764.4000 828.6000 764.5500 ;
	    RECT 822.6000 758.4000 823.8000 759.6000 ;
	    RECT 820.2000 737.4000 821.4000 738.6000 ;
	    RECT 817.8000 713.4000 819.0000 714.6000 ;
	    RECT 817.9500 708.6000 818.8500 713.4000 ;
	    RECT 808.2000 707.4000 809.4000 708.6000 ;
	    RECT 813.0000 707.4000 814.2000 708.6000 ;
	    RECT 817.8000 707.4000 819.0000 708.6000 ;
	    RECT 808.3500 702.6000 809.2500 707.4000 ;
	    RECT 808.2000 701.4000 809.4000 702.6000 ;
	    RECT 810.6000 684.4500 811.8000 684.6000 ;
	    RECT 813.1500 684.4500 814.0500 707.4000 ;
	    RECT 810.6000 683.5500 814.0500 684.4500 ;
	    RECT 810.6000 683.4000 811.8000 683.5500 ;
	    RECT 815.4000 665.4000 816.6000 666.6000 ;
	    RECT 815.5500 645.6000 816.4500 665.4000 ;
	    RECT 815.4000 644.4000 816.6000 645.6000 ;
	    RECT 817.9500 645.4500 818.8500 707.4000 ;
	    RECT 820.3500 654.6000 821.2500 737.4000 ;
	    RECT 822.7500 726.6000 823.6500 758.4000 ;
	    RECT 832.3500 750.6000 833.2500 1097.4000 ;
	    RECT 837.1500 1017.6000 838.0500 1217.4000 ;
	    RECT 839.4000 1206.3000 840.6000 1226.7001 ;
	    RECT 841.8000 1206.3000 843.0000 1226.7001 ;
	    RECT 844.2000 1209.3000 845.4000 1226.7001 ;
	    RECT 846.6000 1220.4000 847.8000 1221.6000 ;
	    RECT 846.7500 1218.6000 847.6500 1220.4000 ;
	    RECT 846.6000 1217.4000 847.8000 1218.6000 ;
	    RECT 849.0000 1209.3000 850.2000 1226.7001 ;
	    RECT 851.5500 1224.6000 852.4500 1265.4000 ;
	    RECT 863.5500 1230.6000 864.4500 1277.5500 ;
	    RECT 868.3500 1250.5500 878.8500 1251.4501 ;
	    RECT 865.8000 1244.4000 867.0000 1245.6000 ;
	    RECT 863.4000 1229.4000 864.6000 1230.6000 ;
	    RECT 851.4000 1223.4000 852.6000 1224.6000 ;
	    RECT 839.4000 1187.4000 840.6000 1188.6000 ;
	    RECT 844.2000 1187.4000 845.4000 1188.6000 ;
	    RECT 844.3500 1185.6000 845.2500 1187.4000 ;
	    RECT 844.2000 1184.4000 845.4000 1185.6000 ;
	    RECT 846.6000 1184.4000 847.8000 1185.6000 ;
	    RECT 839.4000 1163.4000 840.6000 1164.6000 ;
	    RECT 839.5500 1035.6000 840.4500 1163.4000 ;
	    RECT 846.7500 1161.6000 847.6500 1184.4000 ;
	    RECT 851.5500 1182.6000 852.4500 1223.4000 ;
	    RECT 853.8000 1209.3000 855.0000 1226.7001 ;
	    RECT 856.2000 1206.3000 857.4000 1226.7001 ;
	    RECT 858.6000 1206.3000 859.8000 1226.7001 ;
	    RECT 861.0000 1206.3000 862.2000 1226.7001 ;
	    RECT 865.9500 1218.6000 866.8500 1244.4000 ;
	    RECT 868.3500 1242.6000 869.2500 1250.5500 ;
	    RECT 870.6000 1247.4000 871.8000 1248.6000 ;
	    RECT 870.7500 1245.6000 871.6500 1247.4000 ;
	    RECT 877.9500 1245.6000 878.8500 1250.5500 ;
	    RECT 870.6000 1244.4000 871.8000 1245.6000 ;
	    RECT 875.4000 1244.4000 876.6000 1245.6000 ;
	    RECT 877.8000 1244.4000 879.0000 1245.6000 ;
	    RECT 868.2000 1241.4000 869.4000 1242.6000 ;
	    RECT 873.0000 1241.4000 874.2000 1242.6000 ;
	    RECT 873.1500 1230.6000 874.0500 1241.4000 ;
	    RECT 873.0000 1229.4000 874.2000 1230.6000 ;
	    RECT 875.5500 1224.6000 876.4500 1244.4000 ;
	    RECT 877.8000 1241.4000 879.0000 1242.6000 ;
	    RECT 877.9500 1230.6000 878.8500 1241.4000 ;
	    RECT 877.8000 1229.4000 879.0000 1230.6000 ;
	    RECT 868.2000 1223.4000 869.4000 1224.6000 ;
	    RECT 875.4000 1223.4000 876.6000 1224.6000 ;
	    RECT 865.8000 1217.4000 867.0000 1218.6000 ;
	    RECT 863.4000 1199.4000 864.6000 1200.6000 ;
	    RECT 863.5500 1182.6000 864.4500 1199.4000 ;
	    RECT 851.4000 1181.4000 852.6000 1182.6000 ;
	    RECT 863.4000 1181.4000 864.6000 1182.6000 ;
	    RECT 849.0000 1169.4000 850.2000 1170.6000 ;
	    RECT 849.1500 1164.6000 850.0500 1169.4000 ;
	    RECT 849.0000 1163.4000 850.2000 1164.6000 ;
	    RECT 846.6000 1160.4000 847.8000 1161.6000 ;
	    RECT 849.0000 1160.4000 850.2000 1161.6000 ;
	    RECT 846.6000 1073.4000 847.8000 1074.6000 ;
	    RECT 846.7500 1065.6000 847.6500 1073.4000 ;
	    RECT 846.6000 1064.4000 847.8000 1065.6000 ;
	    RECT 849.1500 1062.6000 850.0500 1160.4000 ;
	    RECT 868.3500 1140.6000 869.2500 1223.4000 ;
	    RECT 875.4000 1211.4000 876.6000 1212.6000 ;
	    RECT 873.0000 1187.4000 874.2000 1188.6000 ;
	    RECT 870.6000 1175.4000 871.8000 1176.6000 ;
	    RECT 870.7500 1164.6000 871.6500 1175.4000 ;
	    RECT 875.5500 1164.6000 876.4500 1211.4000 ;
	    RECT 870.6000 1163.4000 871.8000 1164.6000 ;
	    RECT 875.4000 1163.4000 876.6000 1164.6000 ;
	    RECT 875.4000 1160.4000 876.6000 1161.6000 ;
	    RECT 851.4000 1139.4000 852.6000 1140.6000 ;
	    RECT 868.2000 1139.4000 869.4000 1140.6000 ;
	    RECT 851.5500 1092.6000 852.4500 1139.4000 ;
	    RECT 863.4000 1133.4000 864.6000 1134.6000 ;
	    RECT 851.4000 1091.4000 852.6000 1092.6000 ;
	    RECT 851.5500 1065.6000 852.4500 1091.4000 ;
	    RECT 863.5500 1086.6000 864.4500 1133.4000 ;
	    RECT 873.0000 1097.4000 874.2000 1098.6000 ;
	    RECT 863.4000 1085.4000 864.6000 1086.6000 ;
	    RECT 853.8000 1073.4000 855.0000 1074.6000 ;
	    RECT 851.4000 1064.4000 852.6000 1065.6000 ;
	    RECT 849.0000 1061.4000 850.2000 1062.6000 ;
	    RECT 841.8000 1037.4000 843.0000 1038.6000 ;
	    RECT 839.4000 1034.4000 840.6000 1035.6000 ;
	    RECT 837.0000 1016.4000 838.2000 1017.6000 ;
	    RECT 839.4000 995.4000 840.6000 996.6000 ;
	    RECT 837.0000 983.4000 838.2000 984.6000 ;
	    RECT 837.1500 978.6000 838.0500 983.4000 ;
	    RECT 837.0000 977.4000 838.2000 978.6000 ;
	    RECT 839.5500 975.6000 840.4500 995.4000 ;
	    RECT 839.4000 974.4000 840.6000 975.6000 ;
	    RECT 837.0000 959.4000 838.2000 960.6000 ;
	    RECT 834.6000 944.4000 835.8000 945.6000 ;
	    RECT 834.7500 942.6000 835.6500 944.4000 ;
	    RECT 837.1500 942.6000 838.0500 959.4000 ;
	    RECT 839.4000 947.4000 840.6000 948.6000 ;
	    RECT 839.5500 945.6000 840.4500 947.4000 ;
	    RECT 839.4000 944.4000 840.6000 945.6000 ;
	    RECT 834.6000 941.4000 835.8000 942.6000 ;
	    RECT 837.0000 941.4000 838.2000 942.6000 ;
	    RECT 841.9500 918.6000 842.8500 1037.4000 ;
	    RECT 849.0000 1013.4000 850.2000 1014.6000 ;
	    RECT 844.2000 983.4000 845.4000 984.6000 ;
	    RECT 841.8000 917.4000 843.0000 918.6000 ;
	    RECT 837.0000 881.4000 838.2000 882.6000 ;
	    RECT 834.6000 794.4000 835.8000 795.6000 ;
	    RECT 827.4000 750.4500 828.6000 750.6000 ;
	    RECT 827.4000 749.5500 830.8500 750.4500 ;
	    RECT 827.4000 749.4000 828.6000 749.5500 ;
	    RECT 829.9500 747.4500 830.8500 749.5500 ;
	    RECT 832.2000 749.4000 833.4000 750.6000 ;
	    RECT 829.9500 746.5500 833.2500 747.4500 ;
	    RECT 827.4000 743.4000 828.6000 744.6000 ;
	    RECT 827.5500 741.6000 828.4500 743.4000 ;
	    RECT 832.3500 741.6000 833.2500 746.5500 ;
	    RECT 834.7500 744.6000 835.6500 794.4000 ;
	    RECT 834.6000 743.4000 835.8000 744.6000 ;
	    RECT 827.4000 740.4000 828.6000 741.6000 ;
	    RECT 832.2000 740.4000 833.4000 741.6000 ;
	    RECT 834.7500 738.6000 835.6500 743.4000 ;
	    RECT 837.1500 741.6000 838.0500 881.4000 ;
	    RECT 844.3500 852.6000 845.2500 983.4000 ;
	    RECT 846.6000 953.4000 847.8000 954.6000 ;
	    RECT 846.7500 948.6000 847.6500 953.4000 ;
	    RECT 846.6000 947.4000 847.8000 948.6000 ;
	    RECT 846.6000 911.4000 847.8000 912.6000 ;
	    RECT 846.7500 879.6000 847.6500 911.4000 ;
	    RECT 846.6000 878.4000 847.8000 879.6000 ;
	    RECT 844.2000 851.4000 845.4000 852.6000 ;
	    RECT 841.8000 822.4500 843.0000 822.6000 ;
	    RECT 844.2000 822.4500 845.4000 822.6000 ;
	    RECT 841.8000 821.5500 845.4000 822.4500 ;
	    RECT 841.8000 821.4000 843.0000 821.5500 ;
	    RECT 844.2000 821.4000 845.4000 821.5500 ;
	    RECT 846.6000 821.4000 847.8000 822.6000 ;
	    RECT 846.7500 819.6000 847.6500 821.4000 ;
	    RECT 846.6000 818.4000 847.8000 819.6000 ;
	    RECT 841.8000 797.4000 843.0000 798.6000 ;
	    RECT 844.2000 794.4000 845.4000 795.6000 ;
	    RECT 839.4000 791.4000 840.6000 792.6000 ;
	    RECT 841.8000 791.4000 843.0000 792.6000 ;
	    RECT 839.5500 756.6000 840.4500 791.4000 ;
	    RECT 839.4000 755.4000 840.6000 756.6000 ;
	    RECT 839.4000 749.4000 840.6000 750.6000 ;
	    RECT 837.0000 740.4000 838.2000 741.6000 ;
	    RECT 834.6000 737.4000 835.8000 738.6000 ;
	    RECT 822.6000 725.4000 823.8000 726.6000 ;
	    RECT 827.4000 719.4000 828.6000 720.6000 ;
	    RECT 822.6000 713.4000 823.8000 714.6000 ;
	    RECT 822.7500 705.6000 823.6500 713.4000 ;
	    RECT 822.6000 704.4000 823.8000 705.6000 ;
	    RECT 827.5500 699.6000 828.4500 719.4000 ;
	    RECT 832.2000 704.4000 833.4000 705.6000 ;
	    RECT 829.8000 701.4000 831.0000 702.6000 ;
	    RECT 827.4000 698.4000 828.6000 699.6000 ;
	    RECT 822.6000 680.4000 823.8000 681.6000 ;
	    RECT 820.2000 653.4000 821.4000 654.6000 ;
	    RECT 820.2000 645.4500 821.4000 645.6000 ;
	    RECT 817.9500 644.5500 821.4000 645.4500 ;
	    RECT 820.2000 644.4000 821.4000 644.5500 ;
	    RECT 815.4000 641.4000 816.6000 642.6000 ;
	    RECT 817.8000 641.4000 819.0000 642.6000 ;
	    RECT 805.8000 581.4000 807.0000 582.6000 ;
	    RECT 810.6000 530.4000 811.8000 531.6000 ;
	    RECT 810.7500 522.6000 811.6500 530.4000 ;
	    RECT 810.6000 521.4000 811.8000 522.6000 ;
	    RECT 810.7500 516.6000 811.6500 521.4000 ;
	    RECT 810.6000 515.4000 811.8000 516.6000 ;
	    RECT 786.7500 509.5500 790.0500 510.4500 ;
	    RECT 786.7500 468.6000 787.6500 509.5500 ;
	    RECT 813.0000 509.4000 814.2000 510.6000 ;
	    RECT 789.0000 486.3000 790.2000 506.7000 ;
	    RECT 791.4000 486.3000 792.6000 506.7000 ;
	    RECT 793.8000 486.3000 795.0000 506.7000 ;
	    RECT 796.2000 489.3000 797.4000 506.7000 ;
	    RECT 798.6000 503.4000 799.8000 504.6000 ;
	    RECT 786.6000 467.4000 787.8000 468.6000 ;
	    RECT 793.8000 464.4000 795.0000 465.6000 ;
	    RECT 793.9500 462.6000 794.8500 464.4000 ;
	    RECT 786.6000 461.4000 787.8000 462.6000 ;
	    RECT 789.0000 461.4000 790.2000 462.6000 ;
	    RECT 793.8000 461.4000 795.0000 462.6000 ;
	    RECT 786.6000 443.4000 787.8000 444.6000 ;
	    RECT 784.2000 440.4000 785.4000 441.6000 ;
	    RECT 781.8000 425.4000 783.0000 426.6000 ;
	    RECT 774.6000 407.4000 775.8000 408.6000 ;
	    RECT 769.8000 405.4500 771.0000 405.6000 ;
	    RECT 769.8000 404.5500 778.0500 405.4500 ;
	    RECT 769.8000 404.4000 771.0000 404.5500 ;
	    RECT 777.1500 402.6000 778.0500 404.5500 ;
	    RECT 765.0000 401.4000 766.2000 402.6000 ;
	    RECT 767.4000 401.4000 768.6000 402.6000 ;
	    RECT 774.6000 401.4000 775.8000 402.6000 ;
	    RECT 777.0000 401.4000 778.2000 402.6000 ;
	    RECT 750.6000 371.4000 751.8000 372.6000 ;
	    RECT 767.5500 321.6000 768.4500 401.4000 ;
	    RECT 774.7500 354.6000 775.6500 401.4000 ;
	    RECT 774.6000 353.4000 775.8000 354.6000 ;
	    RECT 755.4000 320.4000 756.6000 321.6000 ;
	    RECT 767.4000 320.4000 768.6000 321.6000 ;
	    RECT 738.6000 317.4000 739.8000 318.6000 ;
	    RECT 753.0000 317.4000 754.2000 318.6000 ;
	    RECT 753.1500 303.4500 754.0500 317.4000 ;
	    RECT 750.7500 302.5500 754.0500 303.4500 ;
	    RECT 721.8000 287.4000 723.0000 288.6000 ;
	    RECT 724.2000 276.3000 725.4000 296.7000 ;
	    RECT 726.6000 276.3000 727.8000 296.7000 ;
	    RECT 729.0000 276.3000 730.2000 296.7000 ;
	    RECT 731.4000 276.3000 732.6000 293.7000 ;
	    RECT 733.8000 281.4000 735.0000 282.6000 ;
	    RECT 733.9500 279.6000 734.8500 281.4000 ;
	    RECT 733.8000 278.4000 735.0000 279.6000 ;
	    RECT 736.2000 276.3000 737.4000 293.7000 ;
	    RECT 738.6000 281.4000 739.8000 282.6000 ;
	    RECT 709.8000 263.4000 711.0000 264.6000 ;
	    RECT 707.4000 257.4000 708.6000 258.6000 ;
	    RECT 717.0000 249.3000 718.2000 266.7000 ;
	    RECT 738.7500 261.6000 739.6500 281.4000 ;
	    RECT 741.0000 276.3000 742.2000 293.7000 ;
	    RECT 743.4000 276.3000 744.6000 296.7000 ;
	    RECT 745.8000 276.3000 747.0000 296.7000 ;
	    RECT 748.2000 287.4000 749.4000 288.6000 ;
	    RECT 748.3500 285.6000 749.2500 287.4000 ;
	    RECT 748.2000 284.4000 749.4000 285.6000 ;
	    RECT 750.7500 273.6000 751.6500 302.5500 ;
	    RECT 753.0000 300.4500 754.2000 300.6000 ;
	    RECT 755.5500 300.4500 756.4500 320.4000 ;
	    RECT 779.4000 317.4000 780.6000 318.6000 ;
	    RECT 753.0000 299.5500 756.4500 300.4500 ;
	    RECT 753.0000 299.4000 754.2000 299.5500 ;
	    RECT 753.1500 288.6000 754.0500 299.4000 ;
	    RECT 753.0000 287.4000 754.2000 288.6000 ;
	    RECT 750.6000 272.4000 751.8000 273.6000 ;
	    RECT 738.6000 260.4000 739.8000 261.6000 ;
	    RECT 724.2000 257.4000 725.4000 258.6000 ;
	    RECT 748.2000 254.4000 749.4000 255.6000 ;
	    RECT 748.3500 246.6000 749.2500 254.4000 ;
	    RECT 748.2000 245.4000 749.4000 246.6000 ;
	    RECT 693.0000 227.4000 694.2000 228.6000 ;
	    RECT 693.1500 222.6000 694.0500 227.4000 ;
	    RECT 750.7500 225.6000 751.6500 272.4000 ;
	    RECT 755.5500 261.6000 756.4500 299.5500 ;
	    RECT 779.5500 282.6000 780.4500 317.4000 ;
	    RECT 786.7500 312.6000 787.6500 443.4000 ;
	    RECT 789.1500 390.6000 790.0500 461.4000 ;
	    RECT 796.2000 443.4000 797.4000 444.6000 ;
	    RECT 796.3500 426.6000 797.2500 443.4000 ;
	    RECT 796.2000 425.4000 797.4000 426.6000 ;
	    RECT 789.0000 389.4000 790.2000 390.6000 ;
	    RECT 798.7500 387.6000 799.6500 503.4000 ;
	    RECT 801.0000 489.3000 802.2000 506.7000 ;
	    RECT 803.4000 503.4000 804.6000 504.6000 ;
	    RECT 803.5500 501.6000 804.4500 503.4000 ;
	    RECT 803.4000 500.4000 804.6000 501.6000 ;
	    RECT 805.8000 489.3000 807.0000 506.7000 ;
	    RECT 808.2000 486.3000 809.4000 506.7000 ;
	    RECT 810.6000 486.3000 811.8000 506.7000 ;
	    RECT 813.1500 498.6000 814.0500 509.4000 ;
	    RECT 815.5500 504.6000 816.4500 641.4000 ;
	    RECT 817.9500 627.6000 818.8500 641.4000 ;
	    RECT 817.8000 626.4000 819.0000 627.6000 ;
	    RECT 820.3500 618.6000 821.2500 644.4000 ;
	    RECT 822.7500 642.6000 823.6500 680.4000 ;
	    RECT 825.0000 677.4000 826.2000 678.6000 ;
	    RECT 822.6000 641.4000 823.8000 642.6000 ;
	    RECT 820.2000 617.4000 821.4000 618.6000 ;
	    RECT 820.2000 587.7000 821.4000 588.9000 ;
	    RECT 825.1500 588.6000 826.0500 677.4000 ;
	    RECT 832.3500 675.6000 833.2500 704.4000 ;
	    RECT 832.2000 674.4000 833.4000 675.6000 ;
	    RECT 832.2000 638.4000 833.4000 639.6000 ;
	    RECT 820.2000 582.6000 821.1000 587.7000 ;
	    RECT 825.0000 587.4000 826.2000 588.6000 ;
	    RECT 829.5000 587.7000 830.7000 588.9000 ;
	    RECT 827.7000 584.7000 828.9000 585.9000 ;
	    RECT 827.7000 582.6000 828.6000 584.7000 ;
	    RECT 817.8000 581.4000 819.0000 582.6000 ;
	    RECT 820.2000 581.7000 828.6000 582.6000 ;
	    RECT 820.2000 580.5000 821.1000 581.7000 ;
	    RECT 822.3000 580.5000 823.5000 580.8000 ;
	    RECT 827.4000 580.5000 828.6000 580.8000 ;
	    RECT 829.8000 580.5000 830.7000 587.7000 ;
	    RECT 820.2000 579.3000 821.4000 580.5000 ;
	    RECT 822.3000 579.6000 830.7000 580.5000 ;
	    RECT 829.5000 579.3000 830.7000 579.6000 ;
	    RECT 817.8000 527.4000 819.0000 528.6000 ;
	    RECT 817.8000 515.4000 819.0000 516.6000 ;
	    RECT 815.4000 503.4000 816.6000 504.6000 ;
	    RECT 813.0000 497.4000 814.2000 498.6000 ;
	    RECT 817.9500 495.6000 818.8500 515.4000 ;
	    RECT 825.0000 509.4000 826.2000 510.6000 ;
	    RECT 820.2000 503.4000 821.4000 504.6000 ;
	    RECT 817.8000 494.4000 819.0000 495.6000 ;
	    RECT 801.0000 479.4000 802.2000 480.6000 ;
	    RECT 801.1500 462.6000 802.0500 479.4000 ;
	    RECT 810.6000 473.4000 811.8000 474.6000 ;
	    RECT 803.4000 467.4000 804.6000 468.6000 ;
	    RECT 801.0000 461.4000 802.2000 462.6000 ;
	    RECT 801.0000 419.4000 802.2000 420.6000 ;
	    RECT 801.1500 402.6000 802.0500 419.4000 ;
	    RECT 801.0000 401.4000 802.2000 402.6000 ;
	    RECT 798.6000 386.4000 799.8000 387.6000 ;
	    RECT 798.7500 384.6000 799.6500 386.4000 ;
	    RECT 798.6000 383.4000 799.8000 384.6000 ;
	    RECT 786.6000 311.4000 787.8000 312.6000 ;
	    RECT 781.8000 299.4000 783.0000 300.6000 ;
	    RECT 779.4000 281.4000 780.6000 282.6000 ;
	    RECT 781.9500 261.6000 782.8500 299.4000 ;
	    RECT 784.2000 281.4000 785.4000 282.6000 ;
	    RECT 755.4000 260.4000 756.6000 261.6000 ;
	    RECT 781.8000 260.4000 783.0000 261.6000 ;
	    RECT 781.9500 258.6000 782.8500 260.4000 ;
	    RECT 781.8000 257.4000 783.0000 258.6000 ;
	    RECT 769.8000 239.4000 771.0000 240.6000 ;
	    RECT 762.6000 227.4000 763.8000 228.6000 ;
	    RECT 721.8000 224.4000 723.0000 225.6000 ;
	    RECT 750.6000 224.4000 751.8000 225.6000 ;
	    RECT 693.0000 221.4000 694.2000 222.6000 ;
	    RECT 695.4000 221.4000 696.6000 222.6000 ;
	    RECT 695.5500 204.6000 696.4500 221.4000 ;
	    RECT 721.9500 210.6000 722.8500 224.4000 ;
	    RECT 724.2000 221.4000 725.4000 222.6000 ;
	    RECT 753.0000 221.4000 754.2000 222.6000 ;
	    RECT 721.8000 209.4000 723.0000 210.6000 ;
	    RECT 695.4000 203.4000 696.6000 204.6000 ;
	    RECT 721.9500 174.6000 722.8500 209.4000 ;
	    RECT 714.6000 156.3000 715.8000 173.7000 ;
	    RECT 721.8000 173.4000 723.0000 174.6000 ;
	    RECT 724.2000 167.4000 725.4000 168.6000 ;
	    RECT 724.3500 165.6000 725.2500 167.4000 ;
	    RECT 724.2000 164.4000 725.4000 165.6000 ;
	    RECT 726.6000 155.4000 727.8000 156.6000 ;
	    RECT 729.0000 156.3000 730.2000 173.7000 ;
	    RECT 743.4000 173.4000 744.6000 174.6000 ;
	    RECT 731.4000 161.4000 732.6000 162.6000 ;
	    RECT 731.5500 156.6000 732.4500 161.4000 ;
	    RECT 733.8000 159.3000 735.0000 167.7000 ;
	    RECT 743.5500 165.6000 744.4500 173.4000 ;
	    RECT 743.4000 164.4000 744.6000 165.6000 ;
	    RECT 753.1500 162.6000 754.0500 221.4000 ;
	    RECT 762.7500 219.6000 763.6500 227.4000 ;
	    RECT 769.9500 222.6000 770.8500 239.4000 ;
	    RECT 769.8000 221.4000 771.0000 222.6000 ;
	    RECT 762.6000 218.4000 763.8000 219.6000 ;
	    RECT 760.2000 215.4000 761.4000 216.6000 ;
	    RECT 760.3500 198.6000 761.2500 215.4000 ;
	    RECT 757.8000 197.4000 759.0000 198.6000 ;
	    RECT 760.2000 197.4000 761.4000 198.6000 ;
	    RECT 767.4000 189.3000 768.6000 206.7000 ;
	    RECT 777.0000 197.4000 778.2000 198.6000 ;
	    RECT 781.8000 189.3000 783.0000 206.7000 ;
	    RECT 784.3500 201.6000 785.2500 281.4000 ;
	    RECT 786.7500 279.6000 787.6500 311.4000 ;
	    RECT 786.6000 278.4000 787.8000 279.6000 ;
	    RECT 796.2000 278.4000 797.4000 279.6000 ;
	    RECT 789.0000 263.4000 790.2000 264.6000 ;
	    RECT 793.8000 257.4000 795.0000 258.6000 ;
	    RECT 793.9500 228.4500 794.8500 257.4000 ;
	    RECT 796.3500 255.6000 797.2500 278.4000 ;
	    RECT 796.2000 254.4000 797.4000 255.6000 ;
	    RECT 796.2000 228.4500 797.4000 228.6000 ;
	    RECT 793.9500 227.5500 797.4000 228.4500 ;
	    RECT 796.2000 227.4000 797.4000 227.5500 ;
	    RECT 793.8000 209.4000 795.0000 210.6000 ;
	    RECT 793.9500 204.6000 794.8500 209.4000 ;
	    RECT 784.2000 200.4000 785.4000 201.6000 ;
	    RECT 779.4000 167.4000 780.6000 168.6000 ;
	    RECT 753.0000 161.4000 754.2000 162.6000 ;
	    RECT 774.6000 161.4000 775.8000 162.6000 ;
	    RECT 731.4000 155.4000 732.6000 156.6000 ;
	    RECT 755.4000 155.4000 756.6000 156.6000 ;
	    RECT 700.2000 140.4000 701.4000 141.6000 ;
	    RECT 700.3500 138.6000 701.2500 140.4000 ;
	    RECT 700.2000 137.4000 701.4000 138.6000 ;
	    RECT 709.8000 129.3000 711.0000 146.7000 ;
	    RECT 719.4000 137.4000 720.6000 138.6000 ;
	    RECT 724.2000 129.3000 725.4000 146.7000 ;
	    RECT 726.7500 141.6000 727.6500 155.4000 ;
	    RECT 726.6000 140.4000 727.8000 141.6000 ;
	    RECT 729.0000 135.3000 730.2000 143.7000 ;
	    RECT 693.0000 116.4000 694.2000 117.6000 ;
	    RECT 693.1500 108.6000 694.0500 116.4000 ;
	    RECT 693.0000 107.4000 694.2000 108.6000 ;
	    RECT 721.8000 107.4000 723.0000 108.6000 ;
	    RECT 721.8000 101.4000 723.0000 102.6000 ;
	    RECT 729.0000 101.4000 730.2000 102.6000 ;
	    RECT 721.9500 84.6000 722.8500 101.4000 ;
	    RECT 729.1500 84.6000 730.0500 101.4000 ;
	    RECT 731.4000 89.4000 732.6000 90.6000 ;
	    RECT 717.0000 83.4000 718.2000 84.6000 ;
	    RECT 721.8000 83.4000 723.0000 84.6000 ;
	    RECT 729.0000 83.4000 730.2000 84.6000 ;
	    RECT 717.1500 60.6000 718.0500 83.4000 ;
	    RECT 729.0000 80.4000 730.2000 81.6000 ;
	    RECT 729.1500 78.6000 730.0500 80.4000 ;
	    RECT 729.0000 77.4000 730.2000 78.6000 ;
	    RECT 724.2000 71.4000 725.4000 72.6000 ;
	    RECT 724.3500 66.6000 725.2500 71.4000 ;
	    RECT 724.2000 65.4000 725.4000 66.6000 ;
	    RECT 690.6000 59.4000 691.8000 60.6000 ;
	    RECT 717.0000 59.4000 718.2000 60.6000 ;
	    RECT 625.8000 53.4000 627.0000 54.6000 ;
	    RECT 585.0000 50.4000 586.2000 51.6000 ;
	    RECT 585.1500 30.6000 586.0500 50.4000 ;
	    RECT 688.2000 36.3000 689.4000 56.7000 ;
	    RECT 690.6000 36.3000 691.8000 56.7000 ;
	    RECT 693.0000 36.3000 694.2000 56.7000 ;
	    RECT 695.4000 36.3000 696.6000 53.7000 ;
	    RECT 697.8000 38.4000 699.0000 39.6000 ;
	    RECT 697.9500 36.6000 698.8500 38.4000 ;
	    RECT 697.8000 35.4000 699.0000 36.6000 ;
	    RECT 700.2000 36.3000 701.4000 53.7000 ;
	    RECT 702.6000 47.4000 703.8000 48.6000 ;
	    RECT 702.7500 42.6000 703.6500 47.4000 ;
	    RECT 702.6000 41.4000 703.8000 42.6000 ;
	    RECT 705.0000 36.3000 706.2000 53.7000 ;
	    RECT 707.4000 36.3000 708.6000 56.7000 ;
	    RECT 709.8000 36.3000 711.0000 56.7000 ;
	    RECT 717.0000 56.4000 718.2000 57.6000 ;
	    RECT 717.1500 48.6000 718.0500 56.4000 ;
	    RECT 731.5500 54.6000 732.4500 89.4000 ;
	    RECT 741.0000 77.4000 742.2000 78.6000 ;
	    RECT 736.2000 74.4000 737.4000 75.6000 ;
	    RECT 736.3500 66.6000 737.2500 74.4000 ;
	    RECT 736.2000 65.4000 737.4000 66.6000 ;
	    RECT 743.4000 66.3000 744.6000 86.7000 ;
	    RECT 745.8000 66.3000 747.0000 86.7000 ;
	    RECT 748.2000 69.3000 749.4000 86.7000 ;
	    RECT 750.6000 83.4000 751.8000 84.6000 ;
	    RECT 750.7500 81.6000 751.6500 83.4000 ;
	    RECT 750.6000 80.4000 751.8000 81.6000 ;
	    RECT 753.0000 69.3000 754.2000 86.7000 ;
	    RECT 755.5500 84.6000 756.4500 155.4000 ;
	    RECT 772.2000 131.4000 773.4000 132.6000 ;
	    RECT 772.3500 105.6000 773.2500 131.4000 ;
	    RECT 772.2000 104.4000 773.4000 105.6000 ;
	    RECT 774.7500 102.6000 775.6500 161.4000 ;
	    RECT 779.5500 159.6000 780.4500 167.4000 ;
	    RECT 779.4000 158.4000 780.6000 159.6000 ;
	    RECT 779.5500 138.6000 780.4500 158.4000 ;
	    RECT 784.3500 150.6000 785.2500 200.4000 ;
	    RECT 786.6000 195.3000 787.8000 203.7000 ;
	    RECT 793.8000 203.4000 795.0000 204.6000 ;
	    RECT 803.5500 162.6000 804.4500 467.4000 ;
	    RECT 805.8000 398.4000 807.0000 399.6000 ;
	    RECT 805.9500 396.6000 806.8500 398.4000 ;
	    RECT 805.8000 395.4000 807.0000 396.6000 ;
	    RECT 808.2000 383.4000 809.4000 384.6000 ;
	    RECT 805.8000 353.4000 807.0000 354.6000 ;
	    RECT 803.4000 161.4000 804.6000 162.6000 ;
	    RECT 784.2000 149.4000 785.4000 150.6000 ;
	    RECT 779.4000 137.4000 780.6000 138.6000 ;
	    RECT 791.4000 119.4000 792.6000 120.6000 ;
	    RECT 791.5500 105.6000 792.4500 119.4000 ;
	    RECT 803.5500 114.6000 804.4500 161.4000 ;
	    RECT 805.8000 129.3000 807.0000 146.7000 ;
	    RECT 805.8000 119.4000 807.0000 120.6000 ;
	    RECT 803.4000 113.4000 804.6000 114.6000 ;
	    RECT 805.9500 108.6000 806.8500 119.4000 ;
	    RECT 805.8000 107.4000 807.0000 108.6000 ;
	    RECT 791.4000 104.4000 792.6000 105.6000 ;
	    RECT 793.8000 104.4000 795.0000 105.6000 ;
	    RECT 769.8000 101.4000 771.0000 102.6000 ;
	    RECT 774.6000 101.4000 775.8000 102.6000 ;
	    RECT 779.4000 101.4000 780.6000 102.6000 ;
	    RECT 769.9500 99.6000 770.8500 101.4000 ;
	    RECT 769.8000 98.4000 771.0000 99.6000 ;
	    RECT 755.4000 83.4000 756.6000 84.6000 ;
	    RECT 731.4000 53.4000 732.6000 54.6000 ;
	    RECT 717.0000 47.4000 718.2000 48.6000 ;
	    RECT 712.2000 44.4000 713.4000 45.6000 ;
	    RECT 712.3500 42.6000 713.2500 44.4000 ;
	    RECT 712.2000 41.4000 713.4000 42.6000 ;
	    RECT 724.2000 41.4000 725.4000 42.6000 ;
	    RECT 731.5500 39.6000 732.4500 53.4000 ;
	    RECT 731.4000 38.4000 732.6000 39.6000 ;
	    RECT 755.5500 36.6000 756.4500 83.4000 ;
	    RECT 757.8000 69.3000 759.0000 86.7000 ;
	    RECT 760.2000 66.3000 761.4000 86.7000 ;
	    RECT 762.6000 66.3000 763.8000 86.7000 ;
	    RECT 765.0000 66.3000 766.2000 86.7000 ;
	    RECT 779.5500 72.6000 780.4500 101.4000 ;
	    RECT 781.8000 98.4000 783.0000 99.6000 ;
	    RECT 781.9500 90.6000 782.8500 98.4000 ;
	    RECT 781.8000 89.4000 783.0000 90.6000 ;
	    RECT 779.4000 71.4000 780.6000 72.6000 ;
	    RECT 760.2000 59.4000 761.4000 60.6000 ;
	    RECT 760.3500 42.6000 761.2500 59.4000 ;
	    RECT 793.9500 48.6000 794.8500 104.4000 ;
	    RECT 798.6000 101.4000 799.8000 102.6000 ;
	    RECT 808.3500 78.6000 809.2500 383.4000 ;
	    RECT 810.7500 300.6000 811.6500 473.4000 ;
	    RECT 820.3500 468.6000 821.2500 503.4000 ;
	    RECT 825.1500 501.6000 826.0500 509.4000 ;
	    RECT 825.0000 500.4000 826.2000 501.6000 ;
	    RECT 832.3500 480.6000 833.2500 638.4000 ;
	    RECT 834.7500 612.6000 835.6500 737.4000 ;
	    RECT 839.5500 666.6000 840.4500 749.4000 ;
	    RECT 839.4000 665.4000 840.6000 666.6000 ;
	    RECT 841.9500 648.6000 842.8500 791.4000 ;
	    RECT 844.3500 696.6000 845.2500 794.4000 ;
	    RECT 846.7500 705.6000 847.6500 818.4000 ;
	    RECT 846.6000 704.4000 847.8000 705.6000 ;
	    RECT 846.6000 701.4000 847.8000 702.6000 ;
	    RECT 846.7500 699.6000 847.6500 701.4000 ;
	    RECT 846.6000 698.4000 847.8000 699.6000 ;
	    RECT 844.2000 695.4000 845.4000 696.6000 ;
	    RECT 841.8000 647.4000 843.0000 648.6000 ;
	    RECT 834.6000 611.4000 835.8000 612.6000 ;
	    RECT 844.3500 588.6000 845.2500 695.4000 ;
	    RECT 849.1500 639.6000 850.0500 1013.4000 ;
	    RECT 851.5500 804.6000 852.4500 1064.4000 ;
	    RECT 853.9500 1062.6000 854.8500 1073.4000 ;
	    RECT 856.2000 1064.4000 857.4000 1065.6000 ;
	    RECT 853.8000 1061.4000 855.0000 1062.6000 ;
	    RECT 856.3500 1059.4501 857.2500 1064.4000 ;
	    RECT 858.6000 1061.4000 859.8000 1062.6000 ;
	    RECT 853.9500 1058.5500 857.2500 1059.4501 ;
	    RECT 853.9500 954.6000 854.8500 1058.5500 ;
	    RECT 856.2000 1040.4000 857.4000 1041.6000 ;
	    RECT 856.3500 960.6000 857.2500 1040.4000 ;
	    RECT 858.7500 1002.6000 859.6500 1061.4000 ;
	    RECT 873.1500 1041.6000 874.0500 1097.4000 ;
	    RECT 873.0000 1040.4000 874.2000 1041.6000 ;
	    RECT 873.0000 1019.4000 874.2000 1020.6000 ;
	    RECT 858.6000 1001.4000 859.8000 1002.6000 ;
	    RECT 865.8000 977.4000 867.0000 978.6000 ;
	    RECT 868.2000 971.4000 869.4000 972.6000 ;
	    RECT 868.3500 966.6000 869.2500 971.4000 ;
	    RECT 868.2000 965.4000 869.4000 966.6000 ;
	    RECT 856.2000 959.4000 857.4000 960.6000 ;
	    RECT 863.4000 959.4000 864.6000 960.6000 ;
	    RECT 853.8000 953.4000 855.0000 954.6000 ;
	    RECT 851.4000 803.4000 852.6000 804.6000 ;
	    RECT 853.9500 792.6000 854.8500 953.4000 ;
	    RECT 856.3500 942.6000 857.2500 959.4000 ;
	    RECT 861.0000 947.4000 862.2000 948.6000 ;
	    RECT 856.2000 942.4500 857.4000 942.6000 ;
	    RECT 856.2000 941.5500 859.6500 942.4500 ;
	    RECT 856.2000 941.4000 857.4000 941.5500 ;
	    RECT 858.7500 915.6000 859.6500 941.5500 ;
	    RECT 861.1500 927.6000 862.0500 947.4000 ;
	    RECT 863.4000 941.4000 864.6000 942.6000 ;
	    RECT 873.1500 939.6000 874.0500 1019.4000 ;
	    RECT 865.8000 938.4000 867.0000 939.6000 ;
	    RECT 873.0000 938.4000 874.2000 939.6000 ;
	    RECT 861.0000 926.4000 862.2000 927.6000 ;
	    RECT 863.4000 926.4000 864.6000 927.6000 ;
	    RECT 858.6000 914.4000 859.8000 915.6000 ;
	    RECT 861.0000 878.4000 862.2000 879.6000 ;
	    RECT 861.1500 852.6000 862.0500 878.4000 ;
	    RECT 861.0000 851.4000 862.2000 852.6000 ;
	    RECT 863.5500 819.6000 864.4500 926.4000 ;
	    RECT 865.9500 822.6000 866.8500 938.4000 ;
	    RECT 870.6000 917.4000 871.8000 918.6000 ;
	    RECT 868.2000 824.4000 869.4000 825.6000 ;
	    RECT 865.8000 821.4000 867.0000 822.6000 ;
	    RECT 863.4000 818.4000 864.6000 819.6000 ;
	    RECT 868.3500 819.4500 869.2500 824.4000 ;
	    RECT 865.9500 818.5500 869.2500 819.4500 ;
	    RECT 858.6000 803.4000 859.8000 804.6000 ;
	    RECT 863.4000 800.4000 864.6000 801.6000 ;
	    RECT 853.8000 791.4000 855.0000 792.6000 ;
	    RECT 856.2000 767.4000 857.4000 768.6000 ;
	    RECT 856.3500 765.6000 857.2500 767.4000 ;
	    RECT 853.8000 764.4000 855.0000 765.6000 ;
	    RECT 856.2000 764.4000 857.4000 765.6000 ;
	    RECT 861.0000 764.4000 862.2000 765.6000 ;
	    RECT 853.9500 762.4500 854.8500 764.4000 ;
	    RECT 861.1500 762.6000 862.0500 764.4000 ;
	    RECT 863.5500 762.6000 864.4500 800.4000 ;
	    RECT 858.6000 762.4500 859.8000 762.6000 ;
	    RECT 853.9500 761.5500 859.8000 762.4500 ;
	    RECT 858.6000 761.4000 859.8000 761.5500 ;
	    RECT 861.0000 761.4000 862.2000 762.6000 ;
	    RECT 863.4000 761.4000 864.6000 762.6000 ;
	    RECT 861.0000 740.4000 862.2000 741.6000 ;
	    RECT 856.2000 734.4000 857.4000 735.6000 ;
	    RECT 856.3500 726.6000 857.2500 734.4000 ;
	    RECT 856.2000 725.4000 857.4000 726.6000 ;
	    RECT 853.8000 707.4000 855.0000 708.6000 ;
	    RECT 851.4000 680.4000 852.6000 681.6000 ;
	    RECT 849.0000 638.4000 850.2000 639.6000 ;
	    RECT 849.0000 635.4000 850.2000 636.6000 ;
	    RECT 837.0000 587.4000 838.2000 588.6000 ;
	    RECT 844.2000 587.4000 845.4000 588.6000 ;
	    RECT 837.1500 582.6000 838.0500 587.4000 ;
	    RECT 837.0000 581.4000 838.2000 582.6000 ;
	    RECT 834.6000 533.4000 835.8000 534.6000 ;
	    RECT 834.7500 525.6000 835.6500 533.4000 ;
	    RECT 837.1500 528.6000 838.0500 581.4000 ;
	    RECT 841.8000 578.4000 843.0000 579.6000 ;
	    RECT 841.9500 531.6000 842.8500 578.4000 ;
	    RECT 849.1500 558.6000 850.0500 635.4000 ;
	    RECT 851.5500 624.6000 852.4500 680.4000 ;
	    RECT 853.8000 665.4000 855.0000 666.6000 ;
	    RECT 853.9500 660.6000 854.8500 665.4000 ;
	    RECT 853.8000 659.4000 855.0000 660.6000 ;
	    RECT 851.4000 623.4000 852.6000 624.6000 ;
	    RECT 856.3500 600.6000 857.2500 725.4000 ;
	    RECT 858.6000 720.4500 859.8000 720.6000 ;
	    RECT 861.1500 720.4500 862.0500 740.4000 ;
	    RECT 858.6000 719.5500 862.0500 720.4500 ;
	    RECT 858.6000 719.4000 859.8000 719.5500 ;
	    RECT 858.7500 702.6000 859.6500 719.4000 ;
	    RECT 858.6000 701.4000 859.8000 702.6000 ;
	    RECT 858.7500 684.6000 859.6500 701.4000 ;
	    RECT 858.6000 683.4000 859.8000 684.6000 ;
	    RECT 863.4000 677.4000 864.6000 678.6000 ;
	    RECT 863.5500 672.6000 864.4500 677.4000 ;
	    RECT 863.4000 671.4000 864.6000 672.6000 ;
	    RECT 865.9500 630.6000 866.8500 818.5500 ;
	    RECT 870.7500 768.6000 871.6500 917.4000 ;
	    RECT 875.5500 828.6000 876.4500 1160.4000 ;
	    RECT 877.8000 1157.4000 879.0000 1158.6000 ;
	    RECT 877.9500 1116.6000 878.8500 1157.4000 ;
	    RECT 877.8000 1115.4000 879.0000 1116.6000 ;
	    RECT 880.3500 1095.6000 881.2500 1343.4000 ;
	    RECT 887.5500 1332.6000 888.4500 1364.4000 ;
	    RECT 904.3500 1332.6000 905.2500 1397.4000 ;
	    RECT 906.6000 1386.3000 907.8000 1406.7001 ;
	    RECT 909.0000 1386.3000 910.2000 1406.7001 ;
	    RECT 911.4000 1389.3000 912.6000 1406.7001 ;
	    RECT 913.8000 1400.4000 915.0000 1401.6000 ;
	    RECT 913.9500 1398.6000 914.8500 1400.4000 ;
	    RECT 913.8000 1397.4000 915.0000 1398.6000 ;
	    RECT 916.2000 1389.3000 917.4000 1406.7001 ;
	    RECT 918.6000 1403.4000 919.8000 1404.6000 ;
	    RECT 918.7500 1380.6000 919.6500 1403.4000 ;
	    RECT 921.0000 1389.3000 922.2000 1406.7001 ;
	    RECT 923.4000 1386.3000 924.6000 1406.7001 ;
	    RECT 925.8000 1386.3000 927.0000 1406.7001 ;
	    RECT 928.2000 1386.3000 929.4000 1406.7001 ;
	    RECT 930.6000 1403.4000 931.8000 1404.6000 ;
	    RECT 930.7500 1398.6000 931.6500 1403.4000 ;
	    RECT 930.6000 1397.4000 931.8000 1398.6000 ;
	    RECT 954.6000 1397.4000 955.8000 1398.6000 ;
	    RECT 942.6000 1392.4501 943.8000 1392.6000 ;
	    RECT 940.3500 1391.5500 943.8000 1392.4501 ;
	    RECT 918.6000 1379.4000 919.8000 1380.6000 ;
	    RECT 923.4000 1379.4000 924.6000 1380.6000 ;
	    RECT 921.0000 1373.4000 922.2000 1374.6000 ;
	    RECT 921.1500 1365.6000 922.0500 1373.4000 ;
	    RECT 921.0000 1364.4000 922.2000 1365.6000 ;
	    RECT 909.0000 1361.4000 910.2000 1362.6000 ;
	    RECT 911.4000 1361.4000 912.6000 1362.6000 ;
	    RECT 887.4000 1331.4000 888.6000 1332.6000 ;
	    RECT 899.4000 1331.4000 900.6000 1332.6000 ;
	    RECT 904.2000 1331.4000 905.4000 1332.6000 ;
	    RECT 899.5500 1326.6000 900.4500 1331.4000 ;
	    RECT 899.4000 1325.4000 900.6000 1326.6000 ;
	    RECT 909.1500 1296.6000 910.0500 1361.4000 ;
	    RECT 911.5500 1338.6000 912.4500 1361.4000 ;
	    RECT 911.4000 1337.4000 912.6000 1338.6000 ;
	    RECT 913.8000 1326.3000 915.0000 1346.7001 ;
	    RECT 916.2000 1326.3000 917.4000 1346.7001 ;
	    RECT 918.6000 1326.3000 919.8000 1346.7001 ;
	    RECT 921.0000 1329.3000 922.2000 1346.7001 ;
	    RECT 923.5500 1344.6000 924.4500 1379.4000 ;
	    RECT 925.8000 1367.4000 927.0000 1368.6000 ;
	    RECT 925.9500 1362.6000 926.8500 1367.4000 ;
	    RECT 925.8000 1361.4000 927.0000 1362.6000 ;
	    RECT 940.3500 1359.6000 941.2500 1391.5500 ;
	    RECT 942.6000 1391.4000 943.8000 1391.5500 ;
	    RECT 945.0000 1391.4000 946.2000 1392.6000 ;
	    RECT 940.2000 1358.4000 941.4000 1359.6000 ;
	    RECT 940.3500 1350.6000 941.2500 1358.4000 ;
	    RECT 940.2000 1349.4000 941.4000 1350.6000 ;
	    RECT 923.4000 1343.4000 924.6000 1344.6000 ;
	    RECT 923.5500 1305.6000 924.4500 1343.4000 ;
	    RECT 925.8000 1329.3000 927.0000 1346.7001 ;
	    RECT 928.2000 1343.4000 929.4000 1344.6000 ;
	    RECT 928.3500 1341.6000 929.2500 1343.4000 ;
	    RECT 928.2000 1340.4000 929.4000 1341.6000 ;
	    RECT 928.2000 1337.4000 929.4000 1338.6000 ;
	    RECT 911.4000 1304.4000 912.6000 1305.6000 ;
	    RECT 923.4000 1304.4000 924.6000 1305.6000 ;
	    RECT 909.0000 1295.4000 910.2000 1296.6000 ;
	    RECT 885.0000 1283.4000 886.2000 1284.6000 ;
	    RECT 882.6000 1277.4000 883.8000 1278.6000 ;
	    RECT 897.0000 1277.4000 898.2000 1278.6000 ;
	    RECT 892.2000 1274.4000 893.4000 1275.6000 ;
	    RECT 882.6000 1271.4000 883.8000 1272.6000 ;
	    RECT 885.0000 1271.4000 886.2000 1272.6000 ;
	    RECT 882.7500 1185.6000 883.6500 1271.4000 ;
	    RECT 885.1500 1266.6000 886.0500 1271.4000 ;
	    RECT 892.3500 1266.6000 893.2500 1274.4000 ;
	    RECT 885.0000 1265.4000 886.2000 1266.6000 ;
	    RECT 892.2000 1265.4000 893.4000 1266.6000 ;
	    RECT 899.4000 1266.3000 900.6000 1286.7001 ;
	    RECT 901.8000 1266.3000 903.0000 1286.7001 ;
	    RECT 904.2000 1269.3000 905.4000 1286.7001 ;
	    RECT 906.6000 1280.4000 907.8000 1281.6000 ;
	    RECT 892.2000 1241.4000 893.4000 1242.6000 ;
	    RECT 892.3500 1236.4501 893.2500 1241.4000 ;
	    RECT 906.7500 1236.6000 907.6500 1280.4000 ;
	    RECT 909.0000 1269.3000 910.2000 1286.7001 ;
	    RECT 911.5500 1284.6000 912.4500 1304.4000 ;
	    RECT 911.4000 1283.4000 912.6000 1284.6000 ;
	    RECT 911.5500 1266.6000 912.4500 1283.4000 ;
	    RECT 913.8000 1269.3000 915.0000 1286.7001 ;
	    RECT 911.4000 1265.4000 912.6000 1266.6000 ;
	    RECT 916.2000 1266.3000 917.4000 1286.7001 ;
	    RECT 918.6000 1266.3000 919.8000 1286.7001 ;
	    RECT 921.0000 1266.3000 922.2000 1286.7001 ;
	    RECT 913.8000 1241.4000 915.0000 1242.6000 ;
	    RECT 909.0000 1238.4000 910.2000 1239.6000 ;
	    RECT 889.9500 1235.5500 893.2500 1236.4501 ;
	    RECT 889.9500 1230.6000 890.8500 1235.5500 ;
	    RECT 906.6000 1235.4000 907.8000 1236.6000 ;
	    RECT 889.8000 1229.4000 891.0000 1230.6000 ;
	    RECT 904.2000 1220.4000 905.4000 1221.6000 ;
	    RECT 904.3500 1200.6000 905.2500 1220.4000 ;
	    RECT 906.6000 1217.4000 907.8000 1218.6000 ;
	    RECT 904.2000 1199.4000 905.4000 1200.6000 ;
	    RECT 889.8000 1193.4000 891.0000 1194.6000 ;
	    RECT 882.6000 1184.4000 883.8000 1185.6000 ;
	    RECT 889.9500 1182.6000 890.8500 1193.4000 ;
	    RECT 892.2000 1187.4000 893.4000 1188.6000 ;
	    RECT 892.3500 1182.6000 893.2500 1187.4000 ;
	    RECT 904.2000 1184.4000 905.4000 1185.6000 ;
	    RECT 889.8000 1181.4000 891.0000 1182.6000 ;
	    RECT 892.2000 1181.4000 893.4000 1182.6000 ;
	    RECT 899.4000 1181.4000 900.6000 1182.6000 ;
	    RECT 899.4000 1175.4000 900.6000 1176.6000 ;
	    RECT 889.8000 1169.4000 891.0000 1170.6000 ;
	    RECT 889.9500 1164.4501 890.8500 1169.4000 ;
	    RECT 892.2000 1164.4501 893.4000 1164.6000 ;
	    RECT 889.9500 1163.5500 893.4000 1164.4501 ;
	    RECT 892.2000 1163.4000 893.4000 1163.5500 ;
	    RECT 904.3500 1107.6000 905.2500 1184.4000 ;
	    RECT 904.2000 1106.4000 905.4000 1107.6000 ;
	    RECT 901.8000 1103.4000 903.0000 1104.6000 ;
	    RECT 880.2000 1094.4000 881.4000 1095.6000 ;
	    RECT 885.0000 1091.4000 886.2000 1092.6000 ;
	    RECT 887.4000 1091.4000 888.6000 1092.6000 ;
	    RECT 877.8000 1061.4000 879.0000 1062.6000 ;
	    RECT 877.9500 1038.6000 878.8500 1061.4000 ;
	    RECT 877.8000 1037.4000 879.0000 1038.6000 ;
	    RECT 887.5500 1020.6000 888.4500 1091.4000 ;
	    RECT 901.9500 1059.6000 902.8500 1103.4000 ;
	    RECT 906.7500 1101.4501 907.6500 1217.4000 ;
	    RECT 909.1500 1215.6000 910.0500 1238.4000 ;
	    RECT 909.0000 1214.4000 910.2000 1215.6000 ;
	    RECT 909.1500 1146.6000 910.0500 1214.4000 ;
	    RECT 911.4000 1169.4000 912.6000 1170.6000 ;
	    RECT 911.5500 1161.6000 912.4500 1169.4000 ;
	    RECT 911.4000 1160.4000 912.6000 1161.6000 ;
	    RECT 913.9500 1158.6000 914.8500 1241.4000 ;
	    RECT 928.3500 1221.6000 929.2500 1337.4000 ;
	    RECT 930.6000 1329.3000 931.8000 1346.7001 ;
	    RECT 933.0000 1326.3000 934.2000 1346.7001 ;
	    RECT 935.4000 1326.3000 936.6000 1346.7001 ;
	    RECT 937.8000 1337.4000 939.0000 1338.6000 ;
	    RECT 937.9500 1278.6000 938.8500 1337.4000 ;
	    RECT 945.1500 1335.6000 946.0500 1391.4000 ;
	    RECT 954.7500 1362.6000 955.6500 1397.4000 ;
	    RECT 957.0000 1385.4000 958.2000 1386.6000 ;
	    RECT 954.6000 1361.4000 955.8000 1362.6000 ;
	    RECT 957.1500 1359.6000 958.0500 1385.4000 ;
	    RECT 961.8000 1361.4000 963.0000 1362.6000 ;
	    RECT 957.0000 1358.4000 958.2000 1359.6000 ;
	    RECT 949.8000 1343.4000 951.0000 1344.6000 ;
	    RECT 949.9500 1341.6000 950.8500 1343.4000 ;
	    RECT 949.8000 1340.4000 951.0000 1341.6000 ;
	    RECT 945.0000 1334.4000 946.2000 1335.6000 ;
	    RECT 942.6000 1325.4000 943.8000 1326.6000 ;
	    RECT 947.4000 1325.4000 948.6000 1326.6000 ;
	    RECT 942.7500 1320.6000 943.6500 1325.4000 ;
	    RECT 942.6000 1319.4000 943.8000 1320.6000 ;
	    RECT 947.5500 1302.6000 948.4500 1325.4000 ;
	    RECT 952.2000 1319.4000 953.4000 1320.6000 ;
	    RECT 952.3500 1308.6000 953.2500 1319.4000 ;
	    RECT 952.2000 1307.4000 953.4000 1308.6000 ;
	    RECT 947.4000 1301.4000 948.6000 1302.6000 ;
	    RECT 930.6000 1277.4000 931.8000 1278.6000 ;
	    RECT 937.8000 1277.4000 939.0000 1278.6000 ;
	    RECT 928.2000 1220.4000 929.4000 1221.6000 ;
	    RECT 925.8000 1217.4000 927.0000 1218.6000 ;
	    RECT 928.2000 1217.4000 929.4000 1218.6000 ;
	    RECT 925.9500 1206.6000 926.8500 1217.4000 ;
	    RECT 925.8000 1205.4000 927.0000 1206.6000 ;
	    RECT 923.4000 1184.4000 924.6000 1185.6000 ;
	    RECT 923.5500 1182.6000 924.4500 1184.4000 ;
	    RECT 923.4000 1181.4000 924.6000 1182.6000 ;
	    RECT 916.2000 1175.4000 917.4000 1176.6000 ;
	    RECT 916.3500 1161.6000 917.2500 1175.4000 ;
	    RECT 916.2000 1160.4000 917.4000 1161.6000 ;
	    RECT 921.0000 1160.4000 922.2000 1161.6000 ;
	    RECT 913.8000 1157.4000 915.0000 1158.6000 ;
	    RECT 918.6000 1157.4000 919.8000 1158.6000 ;
	    RECT 909.0000 1145.4000 910.2000 1146.6000 ;
	    RECT 909.1500 1104.6000 910.0500 1145.4000 ;
	    RECT 913.9500 1134.6000 914.8500 1157.4000 ;
	    RECT 918.7500 1137.6000 919.6500 1157.4000 ;
	    RECT 918.6000 1136.4000 919.8000 1137.6000 ;
	    RECT 913.8000 1133.4000 915.0000 1134.6000 ;
	    RECT 909.0000 1103.4000 910.2000 1104.6000 ;
	    RECT 906.7500 1100.5500 910.0500 1101.4501 ;
	    RECT 906.6000 1067.4000 907.8000 1068.6000 ;
	    RECT 904.2000 1061.4000 905.4000 1062.6000 ;
	    RECT 901.8000 1058.4000 903.0000 1059.6000 ;
	    RECT 901.8000 1046.4000 903.0000 1047.6000 ;
	    RECT 892.2000 1043.4000 893.4000 1044.6000 ;
	    RECT 889.8000 1040.4000 891.0000 1041.6000 ;
	    RECT 889.9500 1032.6000 890.8500 1040.4000 ;
	    RECT 889.8000 1031.4000 891.0000 1032.6000 ;
	    RECT 887.4000 1019.4000 888.6000 1020.6000 ;
	    RECT 892.3500 996.6000 893.2500 1043.4000 ;
	    RECT 901.9500 1014.6000 902.8500 1046.4000 ;
	    RECT 904.3500 1038.6000 905.2500 1061.4000 ;
	    RECT 906.7500 1038.6000 907.6500 1067.4000 ;
	    RECT 904.2000 1037.4000 905.4000 1038.6000 ;
	    RECT 906.6000 1037.4000 907.8000 1038.6000 ;
	    RECT 906.6000 1016.4000 907.8000 1017.6000 ;
	    RECT 901.8000 1013.4000 903.0000 1014.6000 ;
	    RECT 892.2000 995.4000 893.4000 996.6000 ;
	    RECT 904.2000 995.4000 905.4000 996.6000 ;
	    RECT 889.8000 980.4000 891.0000 981.6000 ;
	    RECT 889.9500 975.6000 890.8500 980.4000 ;
	    RECT 889.8000 974.4000 891.0000 975.6000 ;
	    RECT 894.6000 974.4000 895.8000 975.6000 ;
	    RECT 894.7500 948.6000 895.6500 974.4000 ;
	    RECT 899.4000 965.4000 900.6000 966.6000 ;
	    RECT 899.5500 954.6000 900.4500 965.4000 ;
	    RECT 899.4000 953.4000 900.6000 954.6000 ;
	    RECT 894.6000 947.4000 895.8000 948.6000 ;
	    RECT 889.8000 941.4000 891.0000 942.6000 ;
	    RECT 889.9500 939.6000 890.8500 941.4000 ;
	    RECT 889.8000 938.4000 891.0000 939.6000 ;
	    RECT 897.0000 926.4000 898.2000 927.6000 ;
	    RECT 877.8000 911.4000 879.0000 912.6000 ;
	    RECT 875.4000 827.4000 876.6000 828.6000 ;
	    RECT 870.6000 767.4000 871.8000 768.6000 ;
	    RECT 873.0000 764.4000 874.2000 765.6000 ;
	    RECT 873.1500 738.6000 874.0500 764.4000 ;
	    RECT 875.4000 755.4000 876.6000 756.6000 ;
	    RECT 875.5500 744.6000 876.4500 755.4000 ;
	    RECT 875.4000 743.4000 876.6000 744.6000 ;
	    RECT 873.0000 737.4000 874.2000 738.6000 ;
	    RECT 870.6000 707.4000 871.8000 708.6000 ;
	    RECT 868.2000 704.4000 869.4000 705.6000 ;
	    RECT 875.5500 705.4500 876.4500 743.4000 ;
	    RECT 877.9500 708.6000 878.8500 911.4000 ;
	    RECT 887.4000 899.4000 888.6000 900.6000 ;
	    RECT 894.6000 899.4000 895.8000 900.6000 ;
	    RECT 887.5500 888.6000 888.4500 899.4000 ;
	    RECT 887.4000 887.4000 888.6000 888.6000 ;
	    RECT 889.8000 887.4000 891.0000 888.6000 ;
	    RECT 889.9500 885.4500 890.8500 887.4000 ;
	    RECT 894.7500 885.6000 895.6500 899.4000 ;
	    RECT 887.5500 884.5500 890.8500 885.4500 ;
	    RECT 887.5500 882.6000 888.4500 884.5500 ;
	    RECT 892.2000 884.4000 893.4000 885.6000 ;
	    RECT 894.6000 884.4000 895.8000 885.6000 ;
	    RECT 892.3500 882.6000 893.2500 884.4000 ;
	    RECT 885.0000 881.4000 886.2000 882.6000 ;
	    RECT 887.4000 881.4000 888.6000 882.6000 ;
	    RECT 892.2000 881.4000 893.4000 882.6000 ;
	    RECT 897.1500 876.6000 898.0500 926.4000 ;
	    RECT 899.4000 914.4000 900.6000 915.6000 ;
	    RECT 899.5500 882.6000 900.4500 914.4000 ;
	    RECT 899.4000 881.4000 900.6000 882.6000 ;
	    RECT 897.0000 875.4000 898.2000 876.6000 ;
	    RECT 882.6000 848.4000 883.8000 849.6000 ;
	    RECT 880.2000 803.4000 881.4000 804.6000 ;
	    RECT 880.3500 795.6000 881.2500 803.4000 ;
	    RECT 880.2000 794.4000 881.4000 795.6000 ;
	    RECT 882.7500 735.6000 883.6500 848.4000 ;
	    RECT 887.4000 845.4000 888.6000 846.6000 ;
	    RECT 887.5500 840.6000 888.4500 845.4000 ;
	    RECT 887.4000 839.4000 888.6000 840.6000 ;
	    RECT 904.3500 828.6000 905.2500 995.4000 ;
	    RECT 906.7500 960.6000 907.6500 1016.4000 ;
	    RECT 909.1500 990.6000 910.0500 1100.5500 ;
	    RECT 913.9500 1098.6000 914.8500 1133.4000 ;
	    RECT 918.6000 1109.4000 919.8000 1110.6000 ;
	    RECT 913.8000 1097.4000 915.0000 1098.6000 ;
	    RECT 916.2000 1067.4000 917.4000 1068.6000 ;
	    RECT 911.4000 1064.4000 912.6000 1065.6000 ;
	    RECT 911.5500 1041.6000 912.4500 1064.4000 ;
	    RECT 916.3500 1047.6000 917.2500 1067.4000 ;
	    RECT 916.2000 1046.4000 917.4000 1047.6000 ;
	    RECT 911.4000 1040.4000 912.6000 1041.6000 ;
	    RECT 916.2000 1031.4000 917.4000 1032.6000 ;
	    RECT 913.8000 1025.4000 915.0000 1026.6000 ;
	    RECT 909.0000 989.4000 910.2000 990.6000 ;
	    RECT 913.9500 978.6000 914.8500 1025.4000 ;
	    RECT 916.2000 1013.4000 917.4000 1014.6000 ;
	    RECT 916.3500 996.6000 917.2500 1013.4000 ;
	    RECT 916.2000 995.4000 917.4000 996.6000 ;
	    RECT 916.3500 984.6000 917.2500 995.4000 ;
	    RECT 916.2000 983.4000 917.4000 984.6000 ;
	    RECT 918.7500 978.6000 919.6500 1109.4000 ;
	    RECT 921.1500 1059.6000 922.0500 1160.4000 ;
	    RECT 923.4000 1145.4000 924.6000 1146.6000 ;
	    RECT 923.5500 1116.6000 924.4500 1145.4000 ;
	    RECT 925.8000 1136.4000 927.0000 1137.6000 ;
	    RECT 925.9500 1128.6000 926.8500 1136.4000 ;
	    RECT 925.8000 1127.4000 927.0000 1128.6000 ;
	    RECT 930.7500 1125.6000 931.6500 1277.4000 ;
	    RECT 935.4000 1271.4000 936.6000 1272.6000 ;
	    RECT 935.5500 1254.6000 936.4500 1271.4000 ;
	    RECT 945.0000 1265.4000 946.2000 1266.6000 ;
	    RECT 935.4000 1253.4000 936.6000 1254.6000 ;
	    RECT 945.1500 1242.6000 946.0500 1265.4000 ;
	    RECT 945.0000 1241.4000 946.2000 1242.6000 ;
	    RECT 935.4000 1238.4000 936.6000 1239.6000 ;
	    RECT 935.5500 1230.6000 936.4500 1238.4000 ;
	    RECT 935.4000 1229.4000 936.6000 1230.6000 ;
	    RECT 935.5500 1224.6000 936.4500 1229.4000 ;
	    RECT 933.0000 1223.4000 934.2000 1224.6000 ;
	    RECT 935.4000 1223.4000 936.6000 1224.6000 ;
	    RECT 933.1500 1212.6000 934.0500 1223.4000 ;
	    RECT 933.0000 1211.4000 934.2000 1212.6000 ;
	    RECT 947.5500 1200.6000 948.4500 1301.4000 ;
	    RECT 959.4000 1295.4000 960.6000 1296.6000 ;
	    RECT 959.5500 1290.6000 960.4500 1295.4000 ;
	    RECT 959.4000 1289.4000 960.6000 1290.6000 ;
	    RECT 957.0000 1280.4000 958.2000 1281.6000 ;
	    RECT 954.6000 1247.4000 955.8000 1248.6000 ;
	    RECT 954.7500 1245.6000 955.6500 1247.4000 ;
	    RECT 949.8000 1244.4000 951.0000 1245.6000 ;
	    RECT 954.6000 1244.4000 955.8000 1245.6000 ;
	    RECT 949.9500 1242.6000 950.8500 1244.4000 ;
	    RECT 949.8000 1241.4000 951.0000 1242.6000 ;
	    RECT 952.2000 1241.4000 953.4000 1242.6000 ;
	    RECT 949.8000 1217.4000 951.0000 1218.6000 ;
	    RECT 952.3500 1212.6000 953.2500 1241.4000 ;
	    RECT 952.2000 1211.4000 953.4000 1212.6000 ;
	    RECT 947.4000 1199.4000 948.6000 1200.6000 ;
	    RECT 933.0000 1178.4000 934.2000 1179.6000 ;
	    RECT 933.1500 1140.6000 934.0500 1178.4000 ;
	    RECT 954.7500 1158.6000 955.6500 1244.4000 ;
	    RECT 957.1500 1242.6000 958.0500 1280.4000 ;
	    RECT 959.4000 1271.4000 960.6000 1272.6000 ;
	    RECT 959.5500 1257.6000 960.4500 1271.4000 ;
	    RECT 959.4000 1256.4000 960.6000 1257.6000 ;
	    RECT 957.0000 1241.4000 958.2000 1242.6000 ;
	    RECT 959.4000 1235.4000 960.6000 1236.6000 ;
	    RECT 959.5500 1218.6000 960.4500 1235.4000 ;
	    RECT 959.4000 1217.4000 960.6000 1218.6000 ;
	    RECT 957.0000 1199.4000 958.2000 1200.6000 ;
	    RECT 954.6000 1157.4000 955.8000 1158.6000 ;
	    RECT 933.0000 1139.4000 934.2000 1140.6000 ;
	    RECT 930.6000 1124.4000 931.8000 1125.6000 ;
	    RECT 923.4000 1115.4000 924.6000 1116.6000 ;
	    RECT 930.7500 1110.6000 931.6500 1124.4000 ;
	    RECT 933.0000 1116.3000 934.2000 1136.7001 ;
	    RECT 935.4000 1116.3000 936.6000 1136.7001 ;
	    RECT 937.8000 1116.3000 939.0000 1133.7001 ;
	    RECT 940.2000 1121.4000 941.4000 1122.6000 ;
	    RECT 930.6000 1109.4000 931.8000 1110.6000 ;
	    RECT 928.2000 1106.4000 929.4000 1107.6000 ;
	    RECT 923.4000 1064.4000 924.6000 1065.6000 ;
	    RECT 921.0000 1058.4000 922.2000 1059.6000 ;
	    RECT 921.0000 1040.4000 922.2000 1041.6000 ;
	    RECT 921.1500 1032.6000 922.0500 1040.4000 ;
	    RECT 921.0000 1031.4000 922.2000 1032.6000 ;
	    RECT 921.1500 1020.6000 922.0500 1031.4000 ;
	    RECT 921.0000 1019.4000 922.2000 1020.6000 ;
	    RECT 921.0000 1007.4000 922.2000 1008.6000 ;
	    RECT 921.1500 978.6000 922.0500 1007.4000 ;
	    RECT 923.5500 987.6000 924.4500 1064.4000 ;
	    RECT 928.3500 1062.6000 929.2500 1106.4000 ;
	    RECT 930.6000 1103.4000 931.8000 1104.6000 ;
	    RECT 930.7500 1086.6000 931.6500 1103.4000 ;
	    RECT 940.3500 1098.6000 941.2500 1121.4000 ;
	    RECT 942.6000 1116.3000 943.8000 1133.7001 ;
	    RECT 945.0000 1118.4000 946.2000 1119.6000 ;
	    RECT 945.1500 1116.6000 946.0500 1118.4000 ;
	    RECT 945.0000 1115.4000 946.2000 1116.6000 ;
	    RECT 947.4000 1116.3000 948.6000 1133.7001 ;
	    RECT 949.8000 1116.3000 951.0000 1136.7001 ;
	    RECT 952.2000 1116.3000 953.4000 1136.7001 ;
	    RECT 954.6000 1116.3000 955.8000 1136.7001 ;
	    RECT 940.2000 1097.4000 941.4000 1098.6000 ;
	    RECT 940.2000 1094.4000 941.4000 1095.6000 ;
	    RECT 930.6000 1085.4000 931.8000 1086.6000 ;
	    RECT 925.8000 1061.4000 927.0000 1062.6000 ;
	    RECT 928.2000 1061.4000 929.4000 1062.6000 ;
	    RECT 925.9500 1020.6000 926.8500 1061.4000 ;
	    RECT 928.2000 1058.4000 929.4000 1059.6000 ;
	    RECT 925.8000 1019.4000 927.0000 1020.6000 ;
	    RECT 925.9500 1008.6000 926.8500 1019.4000 ;
	    RECT 925.8000 1007.4000 927.0000 1008.6000 ;
	    RECT 923.4000 986.4000 924.6000 987.6000 ;
	    RECT 913.8000 977.4000 915.0000 978.6000 ;
	    RECT 918.6000 977.4000 919.8000 978.6000 ;
	    RECT 921.0000 977.4000 922.2000 978.6000 ;
	    RECT 906.6000 959.4000 907.8000 960.6000 ;
	    RECT 913.8000 941.4000 915.0000 942.6000 ;
	    RECT 913.9500 936.6000 914.8500 941.4000 ;
	    RECT 913.8000 935.4000 915.0000 936.6000 ;
	    RECT 916.2000 923.4000 917.4000 924.6000 ;
	    RECT 906.6000 846.3000 907.8000 866.7000 ;
	    RECT 909.0000 846.3000 910.2000 866.7000 ;
	    RECT 911.4000 846.3000 912.6000 866.7000 ;
	    RECT 913.8000 849.3000 915.0000 866.7000 ;
	    RECT 916.3500 864.6000 917.2500 923.4000 ;
	    RECT 921.0000 911.4000 922.2000 912.6000 ;
	    RECT 921.1500 888.6000 922.0500 911.4000 ;
	    RECT 918.6000 887.4000 919.8000 888.6000 ;
	    RECT 921.0000 887.4000 922.2000 888.6000 ;
	    RECT 918.7500 870.4500 919.6500 887.4000 ;
	    RECT 928.3500 885.6000 929.2500 1058.4000 ;
	    RECT 930.7500 1005.6000 931.6500 1085.4000 ;
	    RECT 940.3500 1077.6000 941.2500 1094.4000 ;
	    RECT 940.2000 1076.4000 941.4000 1077.6000 ;
	    RECT 940.2000 1037.4000 941.4000 1038.6000 ;
	    RECT 930.6000 1004.4000 931.8000 1005.6000 ;
	    RECT 933.0000 996.3000 934.2000 1016.7000 ;
	    RECT 935.4000 996.3000 936.6000 1016.7000 ;
	    RECT 937.8000 996.3000 939.0000 1013.7000 ;
	    RECT 940.3500 1002.6000 941.2500 1037.4000 ;
	    RECT 940.2000 1001.4000 941.4000 1002.6000 ;
	    RECT 942.6000 996.3000 943.8000 1013.7000 ;
	    RECT 945.1500 999.6000 946.0500 1115.4000 ;
	    RECT 957.1500 1041.6000 958.0500 1199.4000 ;
	    RECT 961.9500 1188.4501 962.8500 1361.4000 ;
	    RECT 964.2000 1307.4000 965.4000 1308.6000 ;
	    RECT 964.3500 1254.6000 965.2500 1307.4000 ;
	    RECT 964.2000 1253.4000 965.4000 1254.6000 ;
	    RECT 966.7500 1215.6000 967.6500 1427.4000 ;
	    RECT 1031.5500 1404.6000 1032.4501 1430.4000 ;
	    RECT 976.2000 1403.4000 977.4000 1404.6000 ;
	    RECT 993.0000 1403.4000 994.2000 1404.6000 ;
	    RECT 1012.2000 1403.4000 1013.4000 1404.6000 ;
	    RECT 1031.4000 1403.4000 1032.6000 1404.6000 ;
	    RECT 976.3500 1401.6000 977.2500 1403.4000 ;
	    RECT 969.0000 1400.4000 970.2000 1401.6000 ;
	    RECT 976.2000 1400.4000 977.4000 1401.6000 ;
	    RECT 981.0000 1400.4000 982.2000 1401.6000 ;
	    RECT 969.1500 1392.6000 970.0500 1400.4000 ;
	    RECT 976.2000 1397.4000 977.4000 1398.6000 ;
	    RECT 976.3500 1395.6000 977.2500 1397.4000 ;
	    RECT 976.2000 1394.4000 977.4000 1395.6000 ;
	    RECT 969.0000 1391.4000 970.2000 1392.6000 ;
	    RECT 969.1500 1380.6000 970.0500 1391.4000 ;
	    RECT 969.0000 1379.4000 970.2000 1380.6000 ;
	    RECT 978.6000 1379.4000 979.8000 1380.6000 ;
	    RECT 969.1500 1302.6000 970.0500 1379.4000 ;
	    RECT 973.8000 1367.4000 975.0000 1368.6000 ;
	    RECT 973.9500 1356.6000 974.8500 1367.4000 ;
	    RECT 973.8000 1355.4000 975.0000 1356.6000 ;
	    RECT 971.4000 1334.4000 972.6000 1335.6000 ;
	    RECT 971.5500 1305.6000 972.4500 1334.4000 ;
	    RECT 971.4000 1304.4000 972.6000 1305.6000 ;
	    RECT 969.0000 1301.4000 970.2000 1302.6000 ;
	    RECT 973.9500 1284.6000 974.8500 1355.4000 ;
	    RECT 978.7500 1341.6000 979.6500 1379.4000 ;
	    RECT 978.6000 1340.4000 979.8000 1341.6000 ;
	    RECT 976.2000 1331.4000 977.4000 1332.6000 ;
	    RECT 969.0000 1283.4000 970.2000 1284.6000 ;
	    RECT 973.8000 1283.4000 975.0000 1284.6000 ;
	    RECT 969.1500 1254.6000 970.0500 1283.4000 ;
	    RECT 976.3500 1278.6000 977.2500 1331.4000 ;
	    RECT 978.6000 1280.4000 979.8000 1281.6000 ;
	    RECT 976.2000 1277.4000 977.4000 1278.6000 ;
	    RECT 978.7500 1260.6000 979.6500 1280.4000 ;
	    RECT 981.1500 1266.6000 982.0500 1400.4000 ;
	    RECT 993.0000 1397.4000 994.2000 1398.6000 ;
	    RECT 1012.3500 1395.6000 1013.2500 1403.4000 ;
	    RECT 1019.4000 1400.4000 1020.6000 1401.6000 ;
	    RECT 1031.4000 1400.4000 1032.6000 1401.6000 ;
	    RECT 1012.2000 1394.4000 1013.4000 1395.6000 ;
	    RECT 983.4000 1379.4000 984.6000 1380.6000 ;
	    RECT 983.5500 1362.6000 984.4500 1379.4000 ;
	    RECT 1017.0000 1367.4000 1018.2000 1368.6000 ;
	    RECT 1012.2000 1364.4000 1013.4000 1365.6000 ;
	    RECT 983.4000 1361.4000 984.6000 1362.6000 ;
	    RECT 985.8000 1349.4000 987.0000 1350.6000 ;
	    RECT 983.4000 1343.4000 984.6000 1344.6000 ;
	    RECT 983.5500 1308.6000 984.4500 1343.4000 ;
	    RECT 983.4000 1307.4000 984.6000 1308.6000 ;
	    RECT 985.9500 1299.6000 986.8500 1349.4000 ;
	    RECT 997.8000 1313.4000 999.0000 1314.6000 ;
	    RECT 993.0000 1301.4000 994.2000 1302.6000 ;
	    RECT 985.8000 1298.4000 987.0000 1299.6000 ;
	    RECT 983.4000 1283.4000 984.6000 1284.6000 ;
	    RECT 988.2000 1283.4000 989.4000 1284.6000 ;
	    RECT 983.5500 1278.4501 984.4500 1283.4000 ;
	    RECT 988.3500 1281.6000 989.2500 1283.4000 ;
	    RECT 993.1500 1281.6000 994.0500 1301.4000 ;
	    RECT 995.4000 1289.4000 996.6000 1290.6000 ;
	    RECT 995.5500 1281.6000 996.4500 1289.4000 ;
	    RECT 988.2000 1280.4000 989.4000 1281.6000 ;
	    RECT 993.0000 1280.4000 994.2000 1281.6000 ;
	    RECT 995.4000 1280.4000 996.6000 1281.6000 ;
	    RECT 997.9500 1278.6000 998.8500 1313.4000 ;
	    RECT 1012.3500 1308.6000 1013.2500 1364.4000 ;
	    RECT 1017.1500 1362.6000 1018.0500 1367.4000 ;
	    RECT 1017.0000 1361.4000 1018.2000 1362.6000 ;
	    RECT 1019.5500 1341.6000 1020.4500 1400.4000 ;
	    RECT 1031.5500 1380.6000 1032.4501 1400.4000 ;
	    RECT 1031.4000 1379.4000 1032.6000 1380.6000 ;
	    RECT 1031.5500 1344.6000 1032.4501 1379.4000 ;
	    RECT 1031.4000 1343.4000 1032.6000 1344.6000 ;
	    RECT 1041.0000 1343.4000 1042.2001 1344.6000 ;
	    RECT 1041.1500 1341.6000 1042.0500 1343.4000 ;
	    RECT 1019.4000 1340.4000 1020.6000 1341.6000 ;
	    RECT 1041.0000 1340.4000 1042.2001 1341.6000 ;
	    RECT 1021.8000 1337.4000 1023.0000 1338.6000 ;
	    RECT 1012.2000 1307.4000 1013.4000 1308.6000 ;
	    RECT 1012.2000 1301.4000 1013.4000 1302.6000 ;
	    RECT 1019.4000 1301.4000 1020.6000 1302.6000 ;
	    RECT 1005.0000 1298.4000 1006.2000 1299.6000 ;
	    RECT 985.8000 1278.4501 987.0000 1278.6000 ;
	    RECT 983.5500 1277.5500 987.0000 1278.4501 ;
	    RECT 985.8000 1277.4000 987.0000 1277.5500 ;
	    RECT 997.8000 1277.4000 999.0000 1278.6000 ;
	    RECT 981.0000 1265.4000 982.2000 1266.6000 ;
	    RECT 978.6000 1259.4000 979.8000 1260.6000 ;
	    RECT 983.4000 1259.4000 984.6000 1260.6000 ;
	    RECT 985.8000 1259.4000 987.0000 1260.6000 ;
	    RECT 969.0000 1253.4000 970.2000 1254.6000 ;
	    RECT 973.8000 1247.4000 975.0000 1248.6000 ;
	    RECT 973.9500 1221.6000 974.8500 1247.4000 ;
	    RECT 971.4000 1220.4000 972.6000 1221.6000 ;
	    RECT 973.8000 1220.4000 975.0000 1221.6000 ;
	    RECT 971.5500 1218.6000 972.4500 1220.4000 ;
	    RECT 971.4000 1217.4000 972.6000 1218.6000 ;
	    RECT 978.6000 1217.4000 979.8000 1218.6000 ;
	    RECT 983.5500 1218.4501 984.4500 1259.4000 ;
	    RECT 985.9500 1221.6000 986.8500 1259.4000 ;
	    RECT 997.8000 1253.4000 999.0000 1254.6000 ;
	    RECT 1000.2000 1253.4000 1001.4000 1254.6000 ;
	    RECT 985.8000 1220.4000 987.0000 1221.6000 ;
	    RECT 981.1500 1217.5500 984.4500 1218.4501 ;
	    RECT 966.6000 1214.4000 967.8000 1215.6000 ;
	    RECT 971.4000 1214.4000 972.6000 1215.6000 ;
	    RECT 973.8000 1214.4000 975.0000 1215.6000 ;
	    RECT 959.5500 1187.5500 962.8500 1188.4501 ;
	    RECT 959.5500 1182.6000 960.4500 1187.5500 ;
	    RECT 966.6000 1187.4000 967.8000 1188.6000 ;
	    RECT 966.7500 1185.6000 967.6500 1187.4000 ;
	    RECT 961.8000 1184.4000 963.0000 1185.6000 ;
	    RECT 966.6000 1184.4000 967.8000 1185.6000 ;
	    RECT 959.4000 1181.4000 960.6000 1182.6000 ;
	    RECT 961.9500 1164.6000 962.8500 1184.4000 ;
	    RECT 964.2000 1181.4000 965.4000 1182.6000 ;
	    RECT 964.2000 1166.4000 965.4000 1167.6000 ;
	    RECT 961.8000 1163.4000 963.0000 1164.6000 ;
	    RECT 964.3500 1104.6000 965.2500 1166.4000 ;
	    RECT 969.0000 1145.4000 970.2000 1146.6000 ;
	    RECT 969.1500 1131.6000 970.0500 1145.4000 ;
	    RECT 969.0000 1130.4000 970.2000 1131.6000 ;
	    RECT 964.2000 1103.4000 965.4000 1104.6000 ;
	    RECT 971.5500 1074.6000 972.4500 1214.4000 ;
	    RECT 973.9500 1206.6000 974.8500 1214.4000 ;
	    RECT 973.8000 1205.4000 975.0000 1206.6000 ;
	    RECT 981.1500 1182.6000 982.0500 1217.5500 ;
	    RECT 976.2000 1181.4000 977.4000 1182.6000 ;
	    RECT 981.0000 1181.4000 982.2000 1182.6000 ;
	    RECT 983.4000 1181.4000 984.6000 1182.6000 ;
	    RECT 997.9500 1179.6000 998.8500 1253.4000 ;
	    RECT 1000.3500 1179.6000 1001.2500 1253.4000 ;
	    RECT 983.4000 1178.4000 984.6000 1179.6000 ;
	    RECT 997.8000 1178.4000 999.0000 1179.6000 ;
	    RECT 1000.2000 1178.4000 1001.4000 1179.6000 ;
	    RECT 983.5500 1176.6000 984.4500 1178.4000 ;
	    RECT 983.4000 1175.4000 984.6000 1176.6000 ;
	    RECT 973.8000 1163.4000 975.0000 1164.6000 ;
	    RECT 973.9500 1152.6000 974.8500 1163.4000 ;
	    RECT 973.8000 1151.4000 975.0000 1152.6000 ;
	    RECT 997.9500 1146.6000 998.8500 1178.4000 ;
	    RECT 1005.1500 1149.6000 1006.0500 1298.4000 ;
	    RECT 1012.3500 1296.6000 1013.2500 1301.4000 ;
	    RECT 1012.2000 1295.4000 1013.4000 1296.6000 ;
	    RECT 1012.2000 1283.4000 1013.4000 1284.6000 ;
	    RECT 1012.3500 1278.6000 1013.2500 1283.4000 ;
	    RECT 1012.2000 1277.4000 1013.4000 1278.6000 ;
	    RECT 1019.4000 1250.4000 1020.6000 1251.6000 ;
	    RECT 1017.0000 1235.4000 1018.2000 1236.6000 ;
	    RECT 1012.2000 1223.4000 1013.4000 1224.6000 ;
	    RECT 1012.3500 1221.6000 1013.2500 1223.4000 ;
	    RECT 1017.1500 1221.6000 1018.0500 1235.4000 ;
	    RECT 1019.5500 1230.6000 1020.4500 1250.4000 ;
	    RECT 1019.4000 1229.4000 1020.6000 1230.6000 ;
	    RECT 1012.2000 1220.4000 1013.4000 1221.6000 ;
	    RECT 1017.0000 1220.4000 1018.2000 1221.6000 ;
	    RECT 1014.6000 1217.4000 1015.8000 1218.6000 ;
	    RECT 1009.8000 1175.4000 1011.0000 1176.6000 ;
	    RECT 1007.4000 1157.4000 1008.6000 1158.6000 ;
	    RECT 1005.0000 1148.4000 1006.2000 1149.6000 ;
	    RECT 997.8000 1145.4000 999.0000 1146.6000 ;
	    RECT 1005.0000 1139.4000 1006.2000 1140.6000 ;
	    RECT 1002.6000 1133.4000 1003.8000 1134.6000 ;
	    RECT 1002.7500 1125.6000 1003.6500 1133.4000 ;
	    RECT 1002.6000 1124.4000 1003.8000 1125.6000 ;
	    RECT 1005.1500 1122.6000 1006.0500 1139.4000 ;
	    RECT 1007.5500 1125.6000 1008.4500 1157.4000 ;
	    RECT 1007.4000 1124.4000 1008.6000 1125.6000 ;
	    RECT 1000.2000 1121.4000 1001.4000 1122.6000 ;
	    RECT 1005.0000 1121.4000 1006.2000 1122.6000 ;
	    RECT 1007.4000 1121.4000 1008.6000 1122.6000 ;
	    RECT 990.6000 1115.4000 991.8000 1116.6000 ;
	    RECT 981.0000 1086.3000 982.2000 1106.7001 ;
	    RECT 983.4000 1086.3000 984.6000 1106.7001 ;
	    RECT 985.8000 1086.3000 987.0000 1106.7001 ;
	    RECT 988.2000 1089.3000 989.4000 1106.7001 ;
	    RECT 990.7500 1104.6000 991.6500 1115.4000 ;
	    RECT 1000.3500 1110.6000 1001.2500 1121.4000 ;
	    RECT 1000.2000 1109.4000 1001.4000 1110.6000 ;
	    RECT 990.6000 1103.4000 991.8000 1104.6000 ;
	    RECT 990.7500 1086.6000 991.6500 1103.4000 ;
	    RECT 993.0000 1089.3000 994.2000 1106.7001 ;
	    RECT 995.4000 1100.4000 996.6000 1101.6000 ;
	    RECT 990.6000 1085.4000 991.8000 1086.6000 ;
	    RECT 971.4000 1073.4000 972.6000 1074.6000 ;
	    RECT 988.2000 1073.4000 989.4000 1074.6000 ;
	    RECT 957.0000 1040.4000 958.2000 1041.6000 ;
	    RECT 978.6000 1040.4000 979.8000 1041.6000 ;
	    RECT 973.8000 1034.4000 975.0000 1035.6000 ;
	    RECT 945.0000 998.4000 946.2000 999.6000 ;
	    RECT 947.4000 996.3000 948.6000 1013.7000 ;
	    RECT 949.8000 996.3000 951.0000 1016.7000 ;
	    RECT 952.2000 996.3000 953.4000 1016.7000 ;
	    RECT 954.6000 996.3000 955.8000 1016.7000 ;
	    RECT 969.0000 1013.4000 970.2000 1014.6000 ;
	    RECT 969.1500 1011.6000 970.0500 1013.4000 ;
	    RECT 969.0000 1010.4000 970.2000 1011.6000 ;
	    RECT 973.9500 1002.6000 974.8500 1034.4000 ;
	    RECT 973.8000 1001.4000 975.0000 1002.6000 ;
	    RECT 935.4000 986.4000 936.6000 987.6000 ;
	    RECT 930.6000 977.4000 931.8000 978.6000 ;
	    RECT 928.2000 884.4000 929.4000 885.6000 ;
	    RECT 928.2000 881.4000 929.4000 882.6000 ;
	    RECT 928.3500 870.6000 929.2500 881.4000 ;
	    RECT 918.7500 869.5500 922.0500 870.4500 ;
	    RECT 916.2000 863.4000 917.4000 864.6000 ;
	    RECT 904.2000 827.4000 905.4000 828.6000 ;
	    RECT 887.4000 821.4000 888.6000 822.6000 ;
	    RECT 913.8000 821.4000 915.0000 822.6000 ;
	    RECT 887.4000 818.4000 888.6000 819.6000 ;
	    RECT 904.2000 818.4000 905.4000 819.6000 ;
	    RECT 887.5500 804.6000 888.4500 818.4000 ;
	    RECT 887.4000 803.4000 888.6000 804.6000 ;
	    RECT 885.0000 800.4000 886.2000 801.6000 ;
	    RECT 887.4000 800.4000 888.6000 801.6000 ;
	    RECT 885.1500 795.6000 886.0500 800.4000 ;
	    RECT 885.0000 794.4000 886.2000 795.6000 ;
	    RECT 885.0000 761.4000 886.2000 762.6000 ;
	    RECT 885.1500 741.6000 886.0500 761.4000 ;
	    RECT 887.5500 744.6000 888.4500 800.4000 ;
	    RECT 904.3500 792.6000 905.2500 818.4000 ;
	    RECT 904.2000 791.4000 905.4000 792.6000 ;
	    RECT 899.4000 773.4000 900.6000 774.6000 ;
	    RECT 899.5500 765.6000 900.4500 773.4000 ;
	    RECT 901.8000 767.4000 903.0000 768.6000 ;
	    RECT 901.9500 765.6000 902.8500 767.4000 ;
	    RECT 913.9500 765.6000 914.8500 821.4000 ;
	    RECT 899.4000 764.4000 900.6000 765.6000 ;
	    RECT 901.8000 764.4000 903.0000 765.6000 ;
	    RECT 906.6000 764.4000 907.8000 765.6000 ;
	    RECT 913.8000 764.4000 915.0000 765.6000 ;
	    RECT 906.7500 762.6000 907.6500 764.4000 ;
	    RECT 904.2000 761.4000 905.4000 762.6000 ;
	    RECT 906.6000 761.4000 907.8000 762.6000 ;
	    RECT 911.4000 761.4000 912.6000 762.6000 ;
	    RECT 889.8000 755.4000 891.0000 756.6000 ;
	    RECT 889.9500 747.6000 890.8500 755.4000 ;
	    RECT 889.8000 746.4000 891.0000 747.6000 ;
	    RECT 887.4000 743.4000 888.6000 744.6000 ;
	    RECT 885.0000 740.4000 886.2000 741.6000 ;
	    RECT 882.6000 734.4000 883.8000 735.6000 ;
	    RECT 880.2000 725.4000 881.4000 726.6000 ;
	    RECT 880.3500 714.6000 881.2500 725.4000 ;
	    RECT 887.5500 714.6000 888.4500 743.4000 ;
	    RECT 889.8000 728.4000 891.0000 729.6000 ;
	    RECT 880.2000 713.4000 881.4000 714.6000 ;
	    RECT 887.4000 713.4000 888.6000 714.6000 ;
	    RECT 877.8000 707.4000 879.0000 708.6000 ;
	    RECT 875.5500 704.5500 878.8500 705.4500 ;
	    RECT 868.3500 699.4500 869.2500 704.4000 ;
	    RECT 875.4000 701.4000 876.6000 702.6000 ;
	    RECT 868.3500 698.5500 871.6500 699.4500 ;
	    RECT 870.7500 681.6000 871.6500 698.5500 ;
	    RECT 870.6000 680.4000 871.8000 681.6000 ;
	    RECT 868.2000 677.4000 869.4000 678.6000 ;
	    RECT 873.0000 677.4000 874.2000 678.6000 ;
	    RECT 868.3500 654.6000 869.2500 677.4000 ;
	    RECT 868.2000 653.4000 869.4000 654.6000 ;
	    RECT 873.1500 648.6000 874.0500 677.4000 ;
	    RECT 873.0000 647.4000 874.2000 648.6000 ;
	    RECT 865.8000 629.4000 867.0000 630.6000 ;
	    RECT 863.4000 623.4000 864.6000 624.6000 ;
	    RECT 856.2000 599.4000 857.4000 600.6000 ;
	    RECT 861.0000 587.4000 862.2000 588.6000 ;
	    RECT 863.5500 576.6000 864.4500 623.4000 ;
	    RECT 870.6000 590.4000 871.8000 591.6000 ;
	    RECT 870.7500 582.6000 871.6500 590.4000 ;
	    RECT 875.4000 584.4000 876.6000 585.6000 ;
	    RECT 875.5500 582.6000 876.4500 584.4000 ;
	    RECT 870.6000 581.4000 871.8000 582.6000 ;
	    RECT 875.4000 581.4000 876.6000 582.6000 ;
	    RECT 863.4000 575.4000 864.6000 576.6000 ;
	    RECT 849.0000 557.4000 850.2000 558.6000 ;
	    RECT 844.2000 554.4000 845.4000 555.6000 ;
	    RECT 844.3500 543.6000 845.2500 554.4000 ;
	    RECT 851.4000 546.3000 852.6000 566.7000 ;
	    RECT 853.8000 546.3000 855.0000 566.7000 ;
	    RECT 856.2000 549.3000 857.4000 566.7000 ;
	    RECT 858.6000 560.4000 859.8000 561.6000 ;
	    RECT 858.7500 558.6000 859.6500 560.4000 ;
	    RECT 858.6000 557.4000 859.8000 558.6000 ;
	    RECT 858.6000 551.4000 859.8000 552.6000 ;
	    RECT 844.2000 542.4000 845.4000 543.6000 ;
	    RECT 844.3500 540.6000 845.2500 542.4000 ;
	    RECT 844.2000 539.4000 845.4000 540.6000 ;
	    RECT 841.8000 530.4000 843.0000 531.6000 ;
	    RECT 837.0000 527.4000 838.2000 528.6000 ;
	    RECT 834.6000 524.4000 835.8000 525.6000 ;
	    RECT 839.4000 524.4000 840.6000 525.6000 ;
	    RECT 839.5500 522.6000 840.4500 524.4000 ;
	    RECT 839.4000 521.4000 840.6000 522.6000 ;
	    RECT 844.3500 516.6000 845.2500 539.4000 ;
	    RECT 851.4000 533.4000 852.6000 534.6000 ;
	    RECT 851.5500 528.6000 852.4500 533.4000 ;
	    RECT 851.4000 527.4000 852.6000 528.6000 ;
	    RECT 856.2000 527.4000 857.4000 528.6000 ;
	    RECT 856.3500 522.6000 857.2500 527.4000 ;
	    RECT 856.2000 521.4000 857.4000 522.6000 ;
	    RECT 858.7500 519.6000 859.6500 551.4000 ;
	    RECT 861.0000 549.3000 862.2000 566.7000 ;
	    RECT 863.5500 564.6000 864.4500 575.4000 ;
	    RECT 863.4000 563.4000 864.6000 564.6000 ;
	    RECT 863.4000 557.4000 864.6000 558.6000 ;
	    RECT 861.0000 533.4000 862.2000 534.6000 ;
	    RECT 858.6000 518.4000 859.8000 519.6000 ;
	    RECT 844.2000 515.4000 845.4000 516.6000 ;
	    RECT 841.8000 503.4000 843.0000 504.6000 ;
	    RECT 822.6000 479.4000 823.8000 480.6000 ;
	    RECT 832.2000 479.4000 833.4000 480.6000 ;
	    RECT 839.4000 479.4000 840.6000 480.6000 ;
	    RECT 820.2000 467.4000 821.4000 468.6000 ;
	    RECT 815.4000 464.4000 816.6000 465.6000 ;
	    RECT 815.5500 450.6000 816.4500 464.4000 ;
	    RECT 815.4000 449.4000 816.6000 450.6000 ;
	    RECT 817.8000 413.4000 819.0000 414.6000 ;
	    RECT 813.0000 407.4000 814.2000 408.6000 ;
	    RECT 813.0000 356.4000 814.2000 357.6000 ;
	    RECT 813.1500 348.6000 814.0500 356.4000 ;
	    RECT 813.0000 347.4000 814.2000 348.6000 ;
	    RECT 817.9500 345.6000 818.8500 413.4000 ;
	    RECT 822.7500 396.6000 823.6500 479.4000 ;
	    RECT 825.0000 464.4000 826.2000 465.6000 ;
	    RECT 825.1500 432.6000 826.0500 464.4000 ;
	    RECT 839.5500 462.6000 840.4500 479.4000 ;
	    RECT 839.4000 461.4000 840.6000 462.6000 ;
	    RECT 825.0000 431.4000 826.2000 432.6000 ;
	    RECT 841.9500 420.6000 842.8500 503.4000 ;
	    RECT 861.1500 501.6000 862.0500 533.4000 ;
	    RECT 863.5500 501.6000 864.4500 557.4000 ;
	    RECT 865.8000 549.3000 867.0000 566.7000 ;
	    RECT 868.2000 546.3000 869.4000 566.7000 ;
	    RECT 870.6000 546.3000 871.8000 566.7000 ;
	    RECT 873.0000 546.3000 874.2000 566.7000 ;
	    RECT 877.9500 552.6000 878.8500 704.5500 ;
	    RECT 880.2000 704.4000 881.4000 705.6000 ;
	    RECT 877.8000 551.4000 879.0000 552.6000 ;
	    RECT 870.6000 539.4000 871.8000 540.6000 ;
	    RECT 870.7500 522.6000 871.6500 539.4000 ;
	    RECT 873.0000 524.4000 874.2000 525.6000 ;
	    RECT 880.3500 525.4500 881.2500 704.4000 ;
	    RECT 885.0000 665.4000 886.2000 666.6000 ;
	    RECT 882.6000 656.4000 883.8000 657.6000 ;
	    RECT 882.7500 621.6000 883.6500 656.4000 ;
	    RECT 882.6000 620.4000 883.8000 621.6000 ;
	    RECT 882.7500 618.6000 883.6500 620.4000 ;
	    RECT 882.6000 617.4000 883.8000 618.6000 ;
	    RECT 885.1500 528.6000 886.0500 665.4000 ;
	    RECT 889.9500 564.6000 890.8500 728.4000 ;
	    RECT 904.3500 711.4500 905.2500 761.4000 ;
	    RECT 916.3500 732.6000 917.2500 863.4000 ;
	    RECT 918.6000 849.3000 919.8000 866.7000 ;
	    RECT 921.1500 861.6000 922.0500 869.5500 ;
	    RECT 928.2000 869.4000 929.4000 870.6000 ;
	    RECT 921.0000 860.4000 922.2000 861.6000 ;
	    RECT 923.4000 849.3000 924.6000 866.7000 ;
	    RECT 921.0000 845.4000 922.2000 846.6000 ;
	    RECT 925.8000 846.3000 927.0000 866.7000 ;
	    RECT 928.2000 846.3000 929.4000 866.7000 ;
	    RECT 930.7500 858.6000 931.6500 977.4000 ;
	    RECT 933.0000 944.4000 934.2000 945.6000 ;
	    RECT 933.1500 924.6000 934.0500 944.4000 ;
	    RECT 935.5500 942.6000 936.4500 986.4000 ;
	    RECT 973.9500 984.6000 974.8500 1001.4000 ;
	    RECT 952.2000 983.4000 953.4000 984.6000 ;
	    RECT 973.8000 983.4000 975.0000 984.6000 ;
	    RECT 952.3500 981.6000 953.2500 983.4000 ;
	    RECT 952.2000 980.4000 953.4000 981.6000 ;
	    RECT 949.8000 977.4000 951.0000 978.6000 ;
	    RECT 954.6000 977.4000 955.8000 978.6000 ;
	    RECT 954.7500 972.6000 955.6500 977.4000 ;
	    RECT 954.6000 971.4000 955.8000 972.6000 ;
	    RECT 954.7500 966.6000 955.6500 971.4000 ;
	    RECT 954.6000 965.4000 955.8000 966.6000 ;
	    RECT 973.8000 959.4000 975.0000 960.6000 ;
	    RECT 937.8000 944.4000 939.0000 945.6000 ;
	    RECT 935.4000 941.4000 936.6000 942.6000 ;
	    RECT 933.0000 923.4000 934.2000 924.6000 ;
	    RECT 933.1500 888.6000 934.0500 923.4000 ;
	    RECT 937.9500 918.6000 938.8500 944.4000 ;
	    RECT 973.9500 942.6000 974.8500 959.4000 ;
	    RECT 976.2000 947.4000 977.4000 948.6000 ;
	    RECT 940.2000 941.4000 941.4000 942.6000 ;
	    RECT 942.6000 941.4000 943.8000 942.6000 ;
	    RECT 959.4000 941.4000 960.6000 942.6000 ;
	    RECT 973.8000 941.4000 975.0000 942.6000 ;
	    RECT 940.3500 936.6000 941.2500 941.4000 ;
	    RECT 940.2000 935.4000 941.4000 936.6000 ;
	    RECT 937.8000 917.4000 939.0000 918.6000 ;
	    RECT 935.4000 911.4000 936.6000 912.6000 ;
	    RECT 933.0000 887.4000 934.2000 888.6000 ;
	    RECT 935.5500 882.6000 936.4500 911.4000 ;
	    RECT 937.9500 894.6000 938.8500 917.4000 ;
	    RECT 937.8000 893.4000 939.0000 894.6000 ;
	    RECT 940.3500 891.4500 941.2500 935.4000 ;
	    RECT 937.9500 890.5500 941.2500 891.4500 ;
	    RECT 935.4000 881.4000 936.6000 882.6000 ;
	    RECT 933.0000 869.4000 934.2000 870.6000 ;
	    RECT 930.6000 857.4000 931.8000 858.6000 ;
	    RECT 921.1500 825.6000 922.0500 845.4000 ;
	    RECT 923.4000 827.4000 924.6000 828.6000 ;
	    RECT 921.0000 824.4000 922.2000 825.6000 ;
	    RECT 918.6000 821.4000 919.8000 822.6000 ;
	    RECT 906.6000 731.4000 907.8000 732.6000 ;
	    RECT 916.2000 731.4000 917.4000 732.6000 ;
	    RECT 901.9500 710.5500 905.2500 711.4500 ;
	    RECT 901.9500 702.6000 902.8500 710.5500 ;
	    RECT 904.2000 707.4000 905.4000 708.6000 ;
	    RECT 901.8000 701.4000 903.0000 702.6000 ;
	    RECT 904.3500 684.6000 905.2500 707.4000 ;
	    RECT 904.2000 683.4000 905.4000 684.6000 ;
	    RECT 897.0000 617.4000 898.2000 618.6000 ;
	    RECT 892.2000 614.4000 893.4000 615.6000 ;
	    RECT 892.3500 606.6000 893.2500 614.4000 ;
	    RECT 892.2000 605.4000 893.4000 606.6000 ;
	    RECT 899.4000 606.3000 900.6000 626.7000 ;
	    RECT 901.8000 606.3000 903.0000 626.7000 ;
	    RECT 904.2000 609.3000 905.4000 626.7000 ;
	    RECT 906.7500 624.6000 907.6500 731.4000 ;
	    RECT 916.2000 719.4000 917.4000 720.6000 ;
	    RECT 913.8000 713.4000 915.0000 714.6000 ;
	    RECT 913.9500 705.6000 914.8500 713.4000 ;
	    RECT 913.8000 704.4000 915.0000 705.6000 ;
	    RECT 916.3500 702.6000 917.2500 719.4000 ;
	    RECT 918.6000 707.4000 919.8000 708.6000 ;
	    RECT 918.7500 705.6000 919.6500 707.4000 ;
	    RECT 918.6000 704.4000 919.8000 705.6000 ;
	    RECT 911.4000 702.4500 912.6000 702.6000 ;
	    RECT 911.4000 701.5500 914.8500 702.4500 ;
	    RECT 911.4000 701.4000 912.6000 701.5500 ;
	    RECT 913.9500 699.4500 914.8500 701.5500 ;
	    RECT 916.2000 701.4000 917.4000 702.6000 ;
	    RECT 918.6000 701.4000 919.8000 702.6000 ;
	    RECT 921.0000 701.4000 922.2000 702.6000 ;
	    RECT 918.7500 699.4500 919.6500 701.4000 ;
	    RECT 913.9500 698.5500 919.6500 699.4500 ;
	    RECT 913.8000 683.4000 915.0000 684.6000 ;
	    RECT 913.9500 666.6000 914.8500 683.4000 ;
	    RECT 921.1500 681.6000 922.0500 701.4000 ;
	    RECT 921.0000 680.4000 922.2000 681.6000 ;
	    RECT 913.8000 665.4000 915.0000 666.6000 ;
	    RECT 906.6000 623.4000 907.8000 624.6000 ;
	    RECT 906.6000 620.4000 907.8000 621.6000 ;
	    RECT 906.7500 612.6000 907.6500 620.4000 ;
	    RECT 906.6000 611.4000 907.8000 612.6000 ;
	    RECT 909.0000 609.3000 910.2000 626.7000 ;
	    RECT 911.4000 623.4000 912.6000 624.6000 ;
	    RECT 913.8000 609.3000 915.0000 626.7000 ;
	    RECT 913.8000 605.4000 915.0000 606.6000 ;
	    RECT 916.2000 606.3000 917.4000 626.7000 ;
	    RECT 918.6000 606.3000 919.8000 626.7000 ;
	    RECT 921.0000 606.3000 922.2000 626.7000 ;
	    RECT 909.0000 599.4000 910.2000 600.6000 ;
	    RECT 889.8000 563.4000 891.0000 564.6000 ;
	    RECT 887.4000 551.4000 888.6000 552.6000 ;
	    RECT 885.0000 527.4000 886.2000 528.6000 ;
	    RECT 880.3500 524.5500 883.6500 525.4500 ;
	    RECT 868.2000 521.4000 869.4000 522.6000 ;
	    RECT 870.6000 521.4000 871.8000 522.6000 ;
	    RECT 861.0000 500.4000 862.2000 501.6000 ;
	    RECT 863.4000 500.4000 864.6000 501.6000 ;
	    RECT 868.3500 498.6000 869.2500 521.4000 ;
	    RECT 870.7500 501.6000 871.6500 521.4000 ;
	    RECT 870.6000 500.4000 871.8000 501.6000 ;
	    RECT 868.2000 497.4000 869.4000 498.6000 ;
	    RECT 870.6000 497.4000 871.8000 498.6000 ;
	    RECT 863.4000 495.4500 864.6000 495.6000 ;
	    RECT 870.7500 495.4500 871.6500 497.4000 ;
	    RECT 863.4000 494.5500 871.6500 495.4500 ;
	    RECT 863.4000 494.4000 864.6000 494.5500 ;
	    RECT 873.1500 486.6000 874.0500 524.4000 ;
	    RECT 873.0000 485.4000 874.2000 486.6000 ;
	    RECT 844.2000 473.4000 845.4000 474.6000 ;
	    RECT 844.3500 468.6000 845.2500 473.4000 ;
	    RECT 844.2000 467.4000 845.4000 468.6000 ;
	    RECT 863.4000 464.4000 864.6000 465.6000 ;
	    RECT 863.5500 450.6000 864.4500 464.4000 ;
	    RECT 882.7500 453.4500 883.6500 524.5500 ;
	    RECT 904.2000 521.4000 905.4000 522.6000 ;
	    RECT 904.3500 519.6000 905.2500 521.4000 ;
	    RECT 904.2000 518.4000 905.4000 519.6000 ;
	    RECT 889.8000 500.4000 891.0000 501.6000 ;
	    RECT 889.9500 480.6000 890.8500 500.4000 ;
	    RECT 906.6000 494.4000 907.8000 495.6000 ;
	    RECT 889.8000 479.4000 891.0000 480.6000 ;
	    RECT 882.7500 452.5500 886.0500 453.4500 ;
	    RECT 863.4000 449.4000 864.6000 450.6000 ;
	    RECT 870.6000 449.4000 871.8000 450.6000 ;
	    RECT 882.6000 449.4000 883.8000 450.6000 ;
	    RECT 870.7500 441.6000 871.6500 449.4000 ;
	    RECT 870.6000 440.4000 871.8000 441.6000 ;
	    RECT 873.0000 435.3000 874.2000 443.7000 ;
	    RECT 875.4000 440.4000 876.6000 441.6000 ;
	    RECT 875.5500 438.6000 876.4500 440.4000 ;
	    RECT 875.4000 437.4000 876.6000 438.6000 ;
	    RECT 877.8000 429.3000 879.0000 446.7000 ;
	    RECT 882.7500 438.6000 883.6500 449.4000 ;
	    RECT 882.6000 437.4000 883.8000 438.6000 ;
	    RECT 877.8000 425.4000 879.0000 426.6000 ;
	    RECT 841.8000 419.4000 843.0000 420.6000 ;
	    RECT 849.0000 401.4000 850.2000 402.6000 ;
	    RECT 822.6000 395.4000 823.8000 396.6000 ;
	    RECT 822.7500 378.6000 823.6500 395.4000 ;
	    RECT 839.4000 389.4000 840.6000 390.6000 ;
	    RECT 822.6000 377.4000 823.8000 378.6000 ;
	    RECT 825.0000 366.3000 826.2000 386.7000 ;
	    RECT 827.4000 366.3000 828.6000 386.7000 ;
	    RECT 829.8000 366.3000 831.0000 386.7000 ;
	    RECT 832.2000 369.3000 833.4000 386.7000 ;
	    RECT 834.6000 383.4000 835.8000 384.6000 ;
	    RECT 837.0000 369.3000 838.2000 386.7000 ;
	    RECT 839.5500 381.6000 840.4500 389.4000 ;
	    RECT 839.4000 380.4000 840.6000 381.6000 ;
	    RECT 841.8000 369.3000 843.0000 386.7000 ;
	    RECT 844.2000 366.3000 845.4000 386.7000 ;
	    RECT 846.6000 366.3000 847.8000 386.7000 ;
	    RECT 849.1500 378.6000 850.0500 401.4000 ;
	    RECT 877.9500 381.6000 878.8500 425.4000 ;
	    RECT 877.8000 380.4000 879.0000 381.6000 ;
	    RECT 849.0000 377.4000 850.2000 378.6000 ;
	    RECT 856.2000 377.4000 857.4000 378.6000 ;
	    RECT 853.8000 374.4000 855.0000 375.6000 ;
	    RECT 853.9500 363.6000 854.8500 374.4000 ;
	    RECT 853.8000 362.4000 855.0000 363.6000 ;
	    RECT 853.9500 360.6000 854.8500 362.4000 ;
	    RECT 853.8000 359.4000 855.0000 360.6000 ;
	    RECT 817.8000 344.4000 819.0000 345.6000 ;
	    RECT 820.2000 336.3000 821.4000 356.7000 ;
	    RECT 822.6000 336.3000 823.8000 356.7000 ;
	    RECT 825.0000 336.3000 826.2000 353.7000 ;
	    RECT 827.4000 353.4000 828.6000 354.6000 ;
	    RECT 827.5500 342.6000 828.4500 353.4000 ;
	    RECT 827.4000 341.4000 828.6000 342.6000 ;
	    RECT 829.8000 336.3000 831.0000 353.7000 ;
	    RECT 832.2000 338.4000 833.4000 339.6000 ;
	    RECT 832.3500 324.6000 833.2500 338.4000 ;
	    RECT 834.6000 336.3000 835.8000 353.7000 ;
	    RECT 837.0000 336.3000 838.2000 356.7000 ;
	    RECT 839.4000 336.3000 840.6000 356.7000 ;
	    RECT 841.8000 336.3000 843.0000 356.7000 ;
	    RECT 856.3500 351.6000 857.2500 377.4000 ;
	    RECT 882.6000 374.4000 883.8000 375.6000 ;
	    RECT 858.6000 359.4000 859.8000 360.6000 ;
	    RECT 856.2000 350.4000 857.4000 351.6000 ;
	    RECT 858.7500 342.6000 859.6500 359.4000 ;
	    RECT 861.0000 344.4000 862.2000 345.6000 ;
	    RECT 858.6000 341.4000 859.8000 342.6000 ;
	    RECT 832.2000 323.4000 833.4000 324.6000 ;
	    RECT 810.6000 299.4000 811.8000 300.6000 ;
	    RECT 844.2000 284.4000 845.4000 285.6000 ;
	    RECT 844.3500 282.6000 845.2500 284.4000 ;
	    RECT 858.7500 282.6000 859.6500 341.4000 ;
	    RECT 861.1500 315.6000 862.0500 344.4000 ;
	    RECT 882.7500 342.6000 883.6500 374.4000 ;
	    RECT 875.4000 341.4000 876.6000 342.6000 ;
	    RECT 882.6000 341.4000 883.8000 342.6000 ;
	    RECT 861.0000 314.4000 862.2000 315.6000 ;
	    RECT 877.8000 288.4500 879.0000 288.6000 ;
	    RECT 875.5500 287.5500 879.0000 288.4500 ;
	    RECT 873.0000 284.4000 874.2000 285.6000 ;
	    RECT 873.1500 282.6000 874.0500 284.4000 ;
	    RECT 844.2000 281.4000 845.4000 282.6000 ;
	    RECT 858.6000 281.4000 859.8000 282.6000 ;
	    RECT 873.0000 281.4000 874.2000 282.6000 ;
	    RECT 815.4000 263.4000 816.6000 264.6000 ;
	    RECT 815.5500 261.6000 816.4500 263.4000 ;
	    RECT 858.7500 261.6000 859.6500 281.4000 ;
	    RECT 870.6000 269.4000 871.8000 270.6000 ;
	    RECT 815.4000 260.4000 816.6000 261.6000 ;
	    RECT 858.6000 260.4000 859.8000 261.6000 ;
	    RECT 820.2000 257.4000 821.4000 258.6000 ;
	    RECT 837.0000 257.4000 838.2000 258.6000 ;
	    RECT 839.4000 257.4000 840.6000 258.6000 ;
	    RECT 820.3500 255.6000 821.2500 257.4000 ;
	    RECT 820.2000 254.4000 821.4000 255.6000 ;
	    RECT 837.1500 252.6000 838.0500 257.4000 ;
	    RECT 837.0000 251.4000 838.2000 252.6000 ;
	    RECT 839.5500 204.6000 840.4500 257.4000 ;
	    RECT 870.7500 255.6000 871.6500 269.4000 ;
	    RECT 875.5500 258.6000 876.4500 287.5500 ;
	    RECT 877.8000 287.4000 879.0000 287.5500 ;
	    RECT 877.8000 281.4000 879.0000 282.6000 ;
	    RECT 880.2000 281.4000 881.4000 282.6000 ;
	    RECT 877.9500 264.6000 878.8500 281.4000 ;
	    RECT 877.8000 263.4000 879.0000 264.6000 ;
	    RECT 875.4000 257.4000 876.6000 258.6000 ;
	    RECT 870.6000 254.4000 871.8000 255.6000 ;
	    RECT 810.6000 203.4000 811.8000 204.6000 ;
	    RECT 829.8000 203.4000 831.0000 204.6000 ;
	    RECT 839.4000 203.4000 840.6000 204.6000 ;
	    RECT 858.6000 203.4000 859.8000 204.6000 ;
	    RECT 810.7500 198.6000 811.6500 203.4000 ;
	    RECT 829.9500 198.6000 830.8500 203.4000 ;
	    RECT 853.8000 200.4000 855.0000 201.6000 ;
	    RECT 810.6000 197.4000 811.8000 198.6000 ;
	    RECT 829.8000 197.4000 831.0000 198.6000 ;
	    RECT 853.9500 186.6000 854.8500 200.4000 ;
	    RECT 856.2000 197.4000 857.4000 198.6000 ;
	    RECT 853.8000 185.4000 855.0000 186.6000 ;
	    RECT 832.2000 179.4000 833.4000 180.6000 ;
	    RECT 822.6000 149.4000 823.8000 150.6000 ;
	    RECT 815.4000 137.4000 816.6000 138.6000 ;
	    RECT 815.5500 120.6000 816.4500 137.4000 ;
	    RECT 820.2000 129.3000 821.4000 146.7000 ;
	    RECT 822.7500 141.6000 823.6500 149.4000 ;
	    RECT 822.6000 140.4000 823.8000 141.6000 ;
	    RECT 822.7500 120.6000 823.6500 140.4000 ;
	    RECT 825.0000 135.3000 826.2000 143.7000 ;
	    RECT 832.3500 141.6000 833.2500 179.4000 ;
	    RECT 832.2000 140.4000 833.4000 141.6000 ;
	    RECT 853.8000 137.4000 855.0000 138.6000 ;
	    RECT 856.3500 135.4500 857.2500 197.4000 ;
	    RECT 858.7500 195.6000 859.6500 203.4000 ;
	    RECT 882.6000 200.4000 883.8000 201.6000 ;
	    RECT 858.6000 194.4000 859.8000 195.6000 ;
	    RECT 882.7500 156.6000 883.6500 200.4000 ;
	    RECT 885.1500 195.6000 886.0500 452.5500 ;
	    RECT 892.2000 429.3000 893.4000 446.7000 ;
	    RECT 904.2000 443.4000 905.4000 444.6000 ;
	    RECT 899.4000 437.4000 900.6000 438.6000 ;
	    RECT 899.5500 426.6000 900.4500 437.4000 ;
	    RECT 899.4000 425.4000 900.6000 426.6000 ;
	    RECT 904.3500 420.6000 905.2500 443.4000 ;
	    RECT 904.2000 419.4000 905.4000 420.6000 ;
	    RECT 889.8000 197.4000 891.0000 198.6000 ;
	    RECT 885.0000 194.4000 886.2000 195.6000 ;
	    RECT 882.6000 155.4000 883.8000 156.6000 ;
	    RECT 906.7500 150.6000 907.6500 494.4000 ;
	    RECT 909.1500 228.6000 910.0500 599.4000 ;
	    RECT 913.9500 585.6000 914.8500 605.4000 ;
	    RECT 913.8000 584.4000 915.0000 585.6000 ;
	    RECT 911.4000 581.4000 912.6000 582.6000 ;
	    RECT 911.5500 528.6000 912.4500 581.4000 ;
	    RECT 911.4000 527.4000 912.6000 528.6000 ;
	    RECT 918.6000 449.4000 919.8000 450.6000 ;
	    RECT 918.7500 444.6000 919.6500 449.4000 ;
	    RECT 918.6000 443.4000 919.8000 444.6000 ;
	    RECT 916.2000 395.4000 917.4000 396.6000 ;
	    RECT 916.3500 381.6000 917.2500 395.4000 ;
	    RECT 923.5500 384.4500 924.4500 827.4000 ;
	    RECT 930.7500 738.6000 931.6500 857.4000 ;
	    RECT 933.1500 846.4500 934.0500 869.4000 ;
	    RECT 935.4000 854.4000 936.6000 855.6000 ;
	    RECT 935.5500 846.4500 936.4500 854.4000 ;
	    RECT 933.1500 845.5500 936.4500 846.4500 ;
	    RECT 935.5500 843.6000 936.4500 845.5500 ;
	    RECT 935.4000 842.4000 936.6000 843.6000 ;
	    RECT 935.5500 795.6000 936.4500 842.4000 ;
	    RECT 935.4000 794.4000 936.6000 795.6000 ;
	    RECT 935.5500 762.6000 936.4500 794.4000 ;
	    RECT 935.4000 761.4000 936.6000 762.6000 ;
	    RECT 930.6000 737.4000 931.8000 738.6000 ;
	    RECT 925.8000 731.4000 927.0000 732.6000 ;
	    RECT 925.9500 474.6000 926.8500 731.4000 ;
	    RECT 928.2000 578.4000 929.4000 579.6000 ;
	    RECT 928.3500 495.6000 929.2500 578.4000 ;
	    RECT 930.7500 534.6000 931.6500 737.4000 ;
	    RECT 933.0000 680.4000 934.2000 681.6000 ;
	    RECT 933.1500 582.6000 934.0500 680.4000 ;
	    RECT 937.9500 624.6000 938.8500 890.5500 ;
	    RECT 940.2000 887.4000 941.4000 888.6000 ;
	    RECT 940.3500 798.6000 941.2500 887.4000 ;
	    RECT 942.7500 858.6000 943.6500 941.4000 ;
	    RECT 947.4000 917.4000 948.6000 918.6000 ;
	    RECT 947.5500 882.6000 948.4500 917.4000 ;
	    RECT 949.8000 906.3000 951.0000 926.7000 ;
	    RECT 952.2000 906.3000 953.4000 926.7000 ;
	    RECT 954.6000 906.3000 955.8000 926.7000 ;
	    RECT 957.0000 909.3000 958.2000 926.7000 ;
	    RECT 959.4000 923.4000 960.6000 924.6000 ;
	    RECT 961.8000 909.3000 963.0000 926.7000 ;
	    RECT 964.2000 920.4000 965.4000 921.6000 ;
	    RECT 964.3500 918.6000 965.2500 920.4000 ;
	    RECT 964.2000 917.4000 965.4000 918.6000 ;
	    RECT 966.6000 909.3000 967.8000 926.7000 ;
	    RECT 957.0000 905.4000 958.2000 906.6000 ;
	    RECT 966.6000 905.4000 967.8000 906.6000 ;
	    RECT 969.0000 906.3000 970.2000 926.7000 ;
	    RECT 971.4000 906.3000 972.6000 926.7000 ;
	    RECT 973.9500 918.6000 974.8500 941.4000 ;
	    RECT 973.8000 917.4000 975.0000 918.6000 ;
	    RECT 949.8000 884.4000 951.0000 885.6000 ;
	    RECT 945.0000 881.4000 946.2000 882.6000 ;
	    RECT 947.4000 881.4000 948.6000 882.6000 ;
	    RECT 949.9500 861.6000 950.8500 884.4000 ;
	    RECT 957.1500 882.6000 958.0500 905.4000 ;
	    RECT 966.7500 900.6000 967.6500 905.4000 ;
	    RECT 966.6000 899.4000 967.8000 900.6000 ;
	    RECT 957.0000 881.4000 958.2000 882.6000 ;
	    RECT 959.4000 881.4000 960.6000 882.6000 ;
	    RECT 959.5500 879.6000 960.4500 881.4000 ;
	    RECT 959.4000 878.4000 960.6000 879.6000 ;
	    RECT 969.0000 863.4000 970.2000 864.6000 ;
	    RECT 949.8000 860.4000 951.0000 861.6000 ;
	    RECT 942.6000 857.4000 943.8000 858.6000 ;
	    RECT 966.6000 827.4000 967.8000 828.6000 ;
	    RECT 966.7500 825.6000 967.6500 827.4000 ;
	    RECT 961.8000 824.4000 963.0000 825.6000 ;
	    RECT 966.6000 824.4000 967.8000 825.6000 ;
	    RECT 945.0000 821.4000 946.2000 822.6000 ;
	    RECT 942.6000 818.4000 943.8000 819.6000 ;
	    RECT 942.7500 816.6000 943.6500 818.4000 ;
	    RECT 942.6000 815.4000 943.8000 816.6000 ;
	    RECT 940.2000 797.4000 941.4000 798.6000 ;
	    RECT 942.6000 773.4000 943.8000 774.6000 ;
	    RECT 942.7500 768.6000 943.6500 773.4000 ;
	    RECT 942.6000 767.4000 943.8000 768.6000 ;
	    RECT 945.1500 765.4500 946.0500 821.4000 ;
	    RECT 947.4000 809.4000 948.6000 810.6000 ;
	    RECT 942.7500 764.5500 946.0500 765.4500 ;
	    RECT 942.7500 642.6000 943.6500 764.5500 ;
	    RECT 947.5500 762.6000 948.4500 809.4000 ;
	    RECT 959.4000 791.4000 960.6000 792.6000 ;
	    RECT 947.4000 761.4000 948.6000 762.6000 ;
	    RECT 949.8000 761.4000 951.0000 762.6000 ;
	    RECT 959.5500 759.6000 960.4500 791.4000 ;
	    RECT 959.4000 758.4000 960.6000 759.6000 ;
	    RECT 949.8000 725.4000 951.0000 726.6000 ;
	    RECT 945.0000 707.4000 946.2000 708.6000 ;
	    RECT 945.0000 701.4000 946.2000 702.6000 ;
	    RECT 945.1500 684.6000 946.0500 701.4000 ;
	    RECT 945.0000 683.4000 946.2000 684.6000 ;
	    RECT 949.9500 681.6000 950.8500 725.4000 ;
	    RECT 954.6000 701.4000 955.8000 702.6000 ;
	    RECT 952.2000 689.4000 953.4000 690.6000 ;
	    RECT 949.8000 680.4000 951.0000 681.6000 ;
	    RECT 952.3500 678.6000 953.2500 689.4000 ;
	    RECT 945.0000 677.4000 946.2000 678.6000 ;
	    RECT 947.4000 677.4000 948.6000 678.6000 ;
	    RECT 952.2000 677.4000 953.4000 678.6000 ;
	    RECT 945.1500 672.6000 946.0500 677.4000 ;
	    RECT 945.0000 671.4000 946.2000 672.6000 ;
	    RECT 947.5500 660.6000 948.4500 677.4000 ;
	    RECT 954.7500 672.6000 955.6500 701.4000 ;
	    RECT 954.6000 671.4000 955.8000 672.6000 ;
	    RECT 947.4000 659.4000 948.6000 660.6000 ;
	    RECT 961.9500 654.6000 962.8500 824.4000 ;
	    RECT 964.2000 821.4000 965.4000 822.6000 ;
	    RECT 964.3500 816.6000 965.2500 821.4000 ;
	    RECT 964.2000 815.4000 965.4000 816.6000 ;
	    RECT 966.7500 801.6000 967.6500 824.4000 ;
	    RECT 966.6000 800.4000 967.8000 801.6000 ;
	    RECT 966.6000 773.4000 967.8000 774.6000 ;
	    RECT 966.7500 657.6000 967.6500 773.4000 ;
	    RECT 969.1500 759.6000 970.0500 863.4000 ;
	    RECT 973.9500 837.6000 974.8500 917.4000 ;
	    RECT 976.3500 903.4500 977.2500 947.4000 ;
	    RECT 978.7500 930.6000 979.6500 1040.4000 ;
	    RECT 988.3500 984.6000 989.2500 1073.4000 ;
	    RECT 995.5500 1068.6000 996.4500 1100.4000 ;
	    RECT 997.8000 1089.3000 999.0000 1106.7001 ;
	    RECT 997.8000 1085.4000 999.0000 1086.6000 ;
	    RECT 1000.2000 1086.3000 1001.4000 1106.7001 ;
	    RECT 1002.6000 1086.3000 1003.8000 1106.7001 ;
	    RECT 1005.0000 1097.4000 1006.2000 1098.6000 ;
	    RECT 995.4000 1067.4000 996.6000 1068.6000 ;
	    RECT 997.9500 1038.6000 998.8500 1085.4000 ;
	    RECT 1005.1500 1077.6000 1006.0500 1097.4000 ;
	    RECT 1005.0000 1076.4000 1006.2000 1077.6000 ;
	    RECT 997.8000 1037.4000 999.0000 1038.6000 ;
	    RECT 1000.2000 1007.4000 1001.4000 1008.6000 ;
	    RECT 990.6000 998.4000 991.8000 999.6000 ;
	    RECT 988.2000 983.4000 989.4000 984.6000 ;
	    RECT 988.3500 960.6000 989.2500 983.4000 ;
	    RECT 988.2000 959.4000 989.4000 960.6000 ;
	    RECT 990.7500 951.6000 991.6500 998.4000 ;
	    RECT 993.0000 977.4000 994.2000 978.6000 ;
	    RECT 990.6000 950.4000 991.8000 951.6000 ;
	    RECT 1000.3500 945.6000 1001.2500 1007.4000 ;
	    RECT 1002.6000 977.4000 1003.8000 978.6000 ;
	    RECT 1000.2000 944.4000 1001.4000 945.6000 ;
	    RECT 1000.2000 941.4000 1001.4000 942.6000 ;
	    RECT 978.6000 929.4000 979.8000 930.6000 ;
	    RECT 978.6000 914.4000 979.8000 915.6000 ;
	    RECT 978.7500 903.6000 979.6500 914.4000 ;
	    RECT 997.8000 911.4000 999.0000 912.6000 ;
	    RECT 978.6000 903.4500 979.8000 903.6000 ;
	    RECT 976.3500 902.5500 979.8000 903.4500 ;
	    RECT 976.3500 900.6000 977.2500 902.5500 ;
	    RECT 978.6000 902.4000 979.8000 902.5500 ;
	    RECT 976.2000 899.4000 977.4000 900.6000 ;
	    RECT 978.7500 894.6000 979.6500 902.4000 ;
	    RECT 978.6000 893.4000 979.8000 894.6000 ;
	    RECT 988.2000 893.4000 989.4000 894.6000 ;
	    RECT 976.2000 884.4000 977.4000 885.6000 ;
	    RECT 973.8000 836.4000 975.0000 837.6000 ;
	    RECT 973.8000 821.4000 975.0000 822.6000 ;
	    RECT 969.0000 758.4000 970.2000 759.6000 ;
	    RECT 973.8000 758.4000 975.0000 759.6000 ;
	    RECT 971.4000 734.4000 972.6000 735.6000 ;
	    RECT 969.0000 701.4000 970.2000 702.6000 ;
	    RECT 966.6000 656.4000 967.8000 657.6000 ;
	    RECT 961.8000 653.4000 963.0000 654.6000 ;
	    RECT 942.6000 641.4000 943.8000 642.6000 ;
	    RECT 942.6000 638.4000 943.8000 639.6000 ;
	    RECT 940.2000 629.4000 941.4000 630.6000 ;
	    RECT 937.8000 623.4000 939.0000 624.6000 ;
	    RECT 937.9500 612.6000 938.8500 623.4000 ;
	    RECT 935.4000 611.4000 936.6000 612.6000 ;
	    RECT 937.8000 611.4000 939.0000 612.6000 ;
	    RECT 935.5500 582.6000 936.4500 611.4000 ;
	    RECT 933.0000 581.4000 934.2000 582.6000 ;
	    RECT 935.4000 581.4000 936.6000 582.6000 ;
	    RECT 930.6000 533.4000 931.8000 534.6000 ;
	    RECT 928.2000 494.4000 929.4000 495.6000 ;
	    RECT 925.8000 473.4000 927.0000 474.6000 ;
	    RECT 940.3500 402.6000 941.2500 629.4000 ;
	    RECT 940.2000 401.4000 941.4000 402.6000 ;
	    RECT 921.1500 383.5500 924.4500 384.4500 ;
	    RECT 916.2000 380.4000 917.4000 381.6000 ;
	    RECT 921.1500 348.6000 922.0500 383.5500 ;
	    RECT 923.4000 380.4000 924.6000 381.6000 ;
	    RECT 921.0000 347.4000 922.2000 348.6000 ;
	    RECT 916.2000 320.4000 917.4000 321.6000 ;
	    RECT 916.3500 318.6000 917.2500 320.4000 ;
	    RECT 916.2000 317.4000 917.4000 318.6000 ;
	    RECT 923.5500 312.6000 924.4500 380.4000 ;
	    RECT 942.7500 330.6000 943.6500 638.4000 ;
	    RECT 959.4000 620.4000 960.6000 621.6000 ;
	    RECT 949.8000 599.4000 951.0000 600.6000 ;
	    RECT 954.6000 588.4500 955.8000 588.6000 ;
	    RECT 954.6000 587.5500 958.0500 588.4500 ;
	    RECT 954.6000 587.4000 955.8000 587.5500 ;
	    RECT 957.1500 582.6000 958.0500 587.5500 ;
	    RECT 959.5500 585.6000 960.4500 620.4000 ;
	    RECT 961.8000 599.4000 963.0000 600.6000 ;
	    RECT 959.4000 584.4000 960.6000 585.6000 ;
	    RECT 961.9500 582.6000 962.8500 599.4000 ;
	    RECT 964.2000 584.4000 965.4000 585.6000 ;
	    RECT 964.3500 582.6000 965.2500 584.4000 ;
	    RECT 957.0000 581.4000 958.2000 582.6000 ;
	    RECT 961.8000 581.4000 963.0000 582.6000 ;
	    RECT 964.2000 581.4000 965.4000 582.6000 ;
	    RECT 971.5500 570.6000 972.4500 734.4000 ;
	    RECT 973.9500 732.6000 974.8500 758.4000 ;
	    RECT 973.8000 731.4000 975.0000 732.6000 ;
	    RECT 976.3500 708.6000 977.2500 884.4000 ;
	    RECT 988.3500 882.6000 989.2500 893.4000 ;
	    RECT 997.9500 888.6000 998.8500 911.4000 ;
	    RECT 997.8000 887.4000 999.0000 888.6000 ;
	    RECT 988.2000 881.4000 989.4000 882.6000 ;
	    RECT 988.3500 861.6000 989.2500 881.4000 ;
	    RECT 981.0000 860.4000 982.2000 861.6000 ;
	    RECT 988.2000 860.4000 989.4000 861.6000 ;
	    RECT 978.6000 854.4000 979.8000 855.6000 ;
	    RECT 978.7500 840.6000 979.6500 854.4000 ;
	    RECT 981.1500 852.6000 982.0500 860.4000 ;
	    RECT 983.4000 857.4000 984.6000 858.6000 ;
	    RECT 981.0000 851.4000 982.2000 852.6000 ;
	    RECT 978.6000 839.4000 979.8000 840.6000 ;
	    RECT 981.0000 836.4000 982.2000 837.6000 ;
	    RECT 981.1500 708.6000 982.0500 836.4000 ;
	    RECT 983.5500 822.6000 984.4500 857.4000 ;
	    RECT 983.4000 821.4000 984.6000 822.6000 ;
	    RECT 985.8000 821.4000 987.0000 822.6000 ;
	    RECT 988.2000 818.4000 989.4000 819.6000 ;
	    RECT 985.8000 713.4000 987.0000 714.6000 ;
	    RECT 976.2000 707.4000 977.4000 708.6000 ;
	    RECT 981.0000 707.4000 982.2000 708.6000 ;
	    RECT 978.6000 698.4000 979.8000 699.6000 ;
	    RECT 976.2000 671.4000 977.4000 672.6000 ;
	    RECT 973.8000 659.4000 975.0000 660.6000 ;
	    RECT 973.9500 636.6000 974.8500 659.4000 ;
	    RECT 976.3500 657.6000 977.2500 671.4000 ;
	    RECT 976.2000 656.4000 977.4000 657.6000 ;
	    RECT 976.3500 651.4500 977.2500 656.4000 ;
	    RECT 978.7500 654.6000 979.6500 698.4000 ;
	    RECT 978.6000 653.4000 979.8000 654.6000 ;
	    RECT 976.3500 650.5500 979.6500 651.4500 ;
	    RECT 976.3500 648.6000 977.2500 650.5500 ;
	    RECT 976.2000 647.4000 977.4000 648.6000 ;
	    RECT 973.8000 635.4000 975.0000 636.6000 ;
	    RECT 971.4000 569.4000 972.6000 570.6000 ;
	    RECT 959.4000 563.4000 960.6000 564.6000 ;
	    RECT 959.5500 492.6000 960.4500 563.4000 ;
	    RECT 966.6000 555.3000 967.8000 563.7000 ;
	    RECT 969.0000 560.4000 970.2000 561.6000 ;
	    RECT 969.1500 552.6000 970.0500 560.4000 ;
	    RECT 969.0000 551.4000 970.2000 552.6000 ;
	    RECT 971.4000 549.3000 972.6000 566.7000 ;
	    RECT 973.9500 534.6000 974.8500 635.4000 ;
	    RECT 978.7500 588.6000 979.6500 650.5500 ;
	    RECT 981.1500 645.6000 982.0500 707.4000 ;
	    RECT 985.9500 699.6000 986.8500 713.4000 ;
	    RECT 988.3500 699.6000 989.2500 818.4000 ;
	    RECT 995.4000 779.4000 996.6000 780.6000 ;
	    RECT 995.5500 768.6000 996.4500 779.4000 ;
	    RECT 1000.3500 774.6000 1001.2500 941.4000 ;
	    RECT 1000.2000 773.4000 1001.4000 774.6000 ;
	    RECT 995.4000 767.4000 996.6000 768.6000 ;
	    RECT 1000.2000 761.4000 1001.4000 762.6000 ;
	    RECT 1000.3500 744.6000 1001.2500 761.4000 ;
	    RECT 1000.2000 743.4000 1001.4000 744.6000 ;
	    RECT 995.4000 731.4000 996.6000 732.6000 ;
	    RECT 985.8000 698.4000 987.0000 699.6000 ;
	    RECT 988.2000 698.4000 989.4000 699.6000 ;
	    RECT 990.6000 683.4000 991.8000 684.6000 ;
	    RECT 981.0000 644.4000 982.2000 645.6000 ;
	    RECT 981.1500 630.6000 982.0500 644.4000 ;
	    RECT 983.4000 636.3000 984.6000 656.7000 ;
	    RECT 985.8000 636.3000 987.0000 656.7000 ;
	    RECT 988.2000 636.3000 989.4000 653.7000 ;
	    RECT 990.7500 642.6000 991.6500 683.4000 ;
	    RECT 990.6000 641.4000 991.8000 642.6000 ;
	    RECT 993.0000 636.3000 994.2000 653.7000 ;
	    RECT 995.5500 639.6000 996.4500 731.4000 ;
	    RECT 1000.2000 698.4000 1001.4000 699.6000 ;
	    RECT 1000.3500 672.6000 1001.2500 698.4000 ;
	    RECT 1002.7500 690.6000 1003.6500 977.4000 ;
	    RECT 1005.1500 942.6000 1006.0500 1076.4000 ;
	    RECT 1005.0000 941.4000 1006.2000 942.6000 ;
	    RECT 1005.0000 875.4000 1006.2000 876.6000 ;
	    RECT 1005.1500 864.6000 1006.0500 875.4000 ;
	    RECT 1005.0000 863.4000 1006.2000 864.6000 ;
	    RECT 1005.0000 755.4000 1006.2000 756.6000 ;
	    RECT 1005.1500 747.6000 1006.0500 755.4000 ;
	    RECT 1005.0000 746.4000 1006.2000 747.6000 ;
	    RECT 1007.5500 729.6000 1008.4500 1121.4000 ;
	    RECT 1009.9500 1104.6000 1010.8500 1175.4000 ;
	    RECT 1014.7500 1164.6000 1015.6500 1217.4000 ;
	    RECT 1021.9500 1182.6000 1022.8500 1337.4000 ;
	    RECT 1024.2001 1319.4000 1025.4000 1320.6000 ;
	    RECT 1024.3500 1302.6000 1025.2500 1319.4000 ;
	    RECT 1024.2001 1301.4000 1025.4000 1302.6000 ;
	    RECT 1041.0000 1301.4000 1042.2001 1302.6000 ;
	    RECT 1041.1500 1299.6000 1042.0500 1301.4000 ;
	    RECT 1041.0000 1298.4000 1042.2001 1299.6000 ;
	    RECT 1033.8000 1283.4000 1035.0000 1284.6000 ;
	    RECT 1036.2001 1229.4000 1037.4000 1230.6000 ;
	    RECT 1024.2001 1217.4000 1025.4000 1218.6000 ;
	    RECT 1024.3500 1188.6000 1025.2500 1217.4000 ;
	    RECT 1033.8000 1205.4000 1035.0000 1206.6000 ;
	    RECT 1024.2001 1187.4000 1025.4000 1188.6000 ;
	    RECT 1021.8000 1181.4000 1023.0000 1182.6000 ;
	    RECT 1014.6000 1163.4000 1015.8000 1164.6000 ;
	    RECT 1014.7500 1134.6000 1015.6500 1163.4000 ;
	    RECT 1017.0000 1148.4000 1018.2000 1149.6000 ;
	    RECT 1014.6000 1133.4000 1015.8000 1134.6000 ;
	    RECT 1012.2000 1109.4000 1013.4000 1110.6000 ;
	    RECT 1009.8000 1103.4000 1011.0000 1104.6000 ;
	    RECT 1009.8000 1094.4000 1011.0000 1095.6000 ;
	    RECT 1009.9500 1083.6000 1010.8500 1094.4000 ;
	    RECT 1009.8000 1082.4000 1011.0000 1083.6000 ;
	    RECT 1009.9500 1080.6000 1010.8500 1082.4000 ;
	    RECT 1009.8000 1079.4000 1011.0000 1080.6000 ;
	    RECT 1012.3500 1077.4501 1013.2500 1109.4000 ;
	    RECT 1009.9500 1076.5500 1013.2500 1077.4501 ;
	    RECT 1009.9500 1002.6000 1010.8500 1076.5500 ;
	    RECT 1012.2000 1049.4000 1013.4000 1050.6000 ;
	    RECT 1012.3500 1002.6000 1013.2500 1049.4000 ;
	    RECT 1017.1500 1035.6000 1018.0500 1148.4000 ;
	    RECT 1024.3500 1128.6000 1025.2500 1187.4000 ;
	    RECT 1029.0000 1133.4000 1030.2001 1134.6000 ;
	    RECT 1024.2001 1127.4000 1025.4000 1128.6000 ;
	    RECT 1019.4000 1121.4000 1020.6000 1122.6000 ;
	    RECT 1019.5500 1110.6000 1020.4500 1121.4000 ;
	    RECT 1019.4000 1109.4000 1020.6000 1110.6000 ;
	    RECT 1021.8000 1097.4000 1023.0000 1098.6000 ;
	    RECT 1021.9500 1092.6000 1022.8500 1097.4000 ;
	    RECT 1021.8000 1091.4000 1023.0000 1092.6000 ;
	    RECT 1021.8000 1079.4000 1023.0000 1080.6000 ;
	    RECT 1021.9500 1044.4501 1022.8500 1079.4000 ;
	    RECT 1019.5500 1043.5500 1022.8500 1044.4501 ;
	    RECT 1017.0000 1034.4000 1018.2000 1035.6000 ;
	    RECT 1019.5500 1002.6000 1020.4500 1043.5500 ;
	    RECT 1021.9500 1041.6000 1022.8500 1043.5500 ;
	    RECT 1021.8000 1040.4000 1023.0000 1041.6000 ;
	    RECT 1009.8000 1001.4000 1011.0000 1002.6000 ;
	    RECT 1012.2000 1001.4000 1013.4000 1002.6000 ;
	    RECT 1019.4000 1001.4000 1020.6000 1002.6000 ;
	    RECT 1024.3500 978.6000 1025.2500 1127.4000 ;
	    RECT 1026.6000 1040.4000 1027.8000 1041.6000 ;
	    RECT 1026.7500 1005.6000 1027.6500 1040.4000 ;
	    RECT 1026.6000 1004.4000 1027.8000 1005.6000 ;
	    RECT 1026.6000 989.4000 1027.8000 990.6000 ;
	    RECT 1026.7500 981.6000 1027.6500 989.4000 ;
	    RECT 1026.6000 980.4000 1027.8000 981.6000 ;
	    RECT 1029.1500 978.6000 1030.0500 1133.4000 ;
	    RECT 1031.4000 983.4000 1032.6000 984.6000 ;
	    RECT 1031.5500 981.6000 1032.4501 983.4000 ;
	    RECT 1031.4000 980.4000 1032.6000 981.6000 ;
	    RECT 1024.2001 977.4000 1025.4000 978.6000 ;
	    RECT 1029.0000 977.4000 1030.2001 978.6000 ;
	    RECT 1029.1500 972.6000 1030.0500 977.4000 ;
	    RECT 1029.0000 971.4000 1030.2001 972.6000 ;
	    RECT 1024.2001 959.4000 1025.4000 960.6000 ;
	    RECT 1019.4000 956.4000 1020.6000 957.6000 ;
	    RECT 1009.8000 893.4000 1011.0000 894.6000 ;
	    RECT 1009.9500 882.6000 1010.8500 893.4000 ;
	    RECT 1009.8000 881.4000 1011.0000 882.6000 ;
	    RECT 1012.2000 737.4000 1013.4000 738.6000 ;
	    RECT 1007.4000 728.4000 1008.6000 729.6000 ;
	    RECT 1002.6000 689.4000 1003.8000 690.6000 ;
	    RECT 1009.8000 680.4000 1011.0000 681.6000 ;
	    RECT 1000.2000 671.4000 1001.4000 672.6000 ;
	    RECT 1007.4000 671.4000 1008.6000 672.6000 ;
	    RECT 995.4000 638.4000 996.6000 639.6000 ;
	    RECT 997.8000 636.3000 999.0000 653.7000 ;
	    RECT 1000.2000 636.3000 1001.4000 656.7000 ;
	    RECT 1002.6000 636.3000 1003.8000 656.7000 ;
	    RECT 1005.0000 636.3000 1006.2000 656.7000 ;
	    RECT 981.0000 629.4000 982.2000 630.6000 ;
	    RECT 1000.2000 629.4000 1001.4000 630.6000 ;
	    RECT 978.6000 587.4000 979.8000 588.6000 ;
	    RECT 978.7500 576.6000 979.6500 587.4000 ;
	    RECT 978.6000 575.4000 979.8000 576.6000 ;
	    RECT 976.2000 569.4000 977.4000 570.6000 ;
	    RECT 976.3500 558.6000 977.2500 569.4000 ;
	    RECT 976.2000 557.4000 977.4000 558.6000 ;
	    RECT 978.6000 551.4000 979.8000 552.6000 ;
	    RECT 973.8000 533.4000 975.0000 534.6000 ;
	    RECT 973.8000 527.4000 975.0000 528.6000 ;
	    RECT 973.9500 522.6000 974.8500 527.4000 ;
	    RECT 973.8000 521.4000 975.0000 522.6000 ;
	    RECT 976.2000 519.3000 977.4000 527.7000 ;
	    RECT 978.7500 522.6000 979.6500 551.4000 ;
	    RECT 985.8000 549.3000 987.0000 566.7000 ;
	    RECT 993.0000 557.4000 994.2000 558.6000 ;
	    RECT 978.6000 521.4000 979.8000 522.6000 ;
	    RECT 978.7500 492.6000 979.6500 521.4000 ;
	    RECT 981.0000 516.3000 982.2000 533.7000 ;
	    RECT 988.2000 533.4000 989.4000 534.6000 ;
	    RECT 985.8000 527.4000 987.0000 528.6000 ;
	    RECT 985.9500 525.6000 986.8500 527.4000 ;
	    RECT 985.8000 524.4000 987.0000 525.6000 ;
	    RECT 959.4000 491.4000 960.6000 492.6000 ;
	    RECT 978.6000 491.4000 979.8000 492.6000 ;
	    RECT 945.0000 459.3000 946.2000 467.7000 ;
	    RECT 947.4000 461.4000 948.6000 462.6000 ;
	    RECT 947.5500 438.6000 948.4500 461.4000 ;
	    RECT 949.8000 456.3000 951.0000 473.7000 ;
	    RECT 954.6000 464.4000 955.8000 465.6000 ;
	    RECT 954.7500 456.6000 955.6500 464.4000 ;
	    RECT 954.6000 455.4000 955.8000 456.6000 ;
	    RECT 964.2000 456.3000 965.4000 473.7000 ;
	    RECT 971.4000 464.4000 972.6000 465.6000 ;
	    RECT 971.5500 441.6000 972.4500 464.4000 ;
	    RECT 957.0000 440.4000 958.2000 441.6000 ;
	    RECT 971.4000 440.4000 972.6000 441.6000 ;
	    RECT 957.1500 438.6000 958.0500 440.4000 ;
	    RECT 947.4000 437.4000 948.6000 438.6000 ;
	    RECT 957.0000 437.4000 958.2000 438.6000 ;
	    RECT 947.5500 426.6000 948.4500 437.4000 ;
	    RECT 947.4000 425.4000 948.6000 426.6000 ;
	    RECT 952.2000 416.4000 953.4000 417.6000 ;
	    RECT 952.3500 408.6000 953.2500 416.4000 ;
	    RECT 945.0000 407.4000 946.2000 408.6000 ;
	    RECT 952.2000 407.4000 953.4000 408.6000 ;
	    RECT 945.1500 405.6000 946.0500 407.4000 ;
	    RECT 957.1500 405.6000 958.0500 437.4000 ;
	    RECT 978.7500 426.6000 979.6500 491.4000 ;
	    RECT 971.4000 425.4000 972.6000 426.6000 ;
	    RECT 978.6000 425.4000 979.8000 426.6000 ;
	    RECT 945.0000 404.4000 946.2000 405.6000 ;
	    RECT 957.0000 404.4000 958.2000 405.6000 ;
	    RECT 959.4000 396.3000 960.6000 416.7000 ;
	    RECT 961.8000 396.3000 963.0000 416.7000 ;
	    RECT 964.2000 396.3000 965.4000 413.7000 ;
	    RECT 966.6000 401.4000 967.8000 402.6000 ;
	    RECT 966.7500 396.6000 967.6500 401.4000 ;
	    RECT 966.6000 395.4000 967.8000 396.6000 ;
	    RECT 969.0000 396.3000 970.2000 413.7000 ;
	    RECT 971.5500 399.6000 972.4500 425.4000 ;
	    RECT 971.4000 398.4000 972.6000 399.6000 ;
	    RECT 969.0000 383.4000 970.2000 384.6000 ;
	    RECT 957.0000 365.4000 958.2000 366.6000 ;
	    RECT 942.6000 329.4000 943.8000 330.6000 ;
	    RECT 923.4000 311.4000 924.6000 312.6000 ;
	    RECT 933.0000 306.3000 934.2000 326.7000 ;
	    RECT 935.4000 306.3000 936.6000 326.7000 ;
	    RECT 937.8000 306.3000 939.0000 326.7000 ;
	    RECT 940.2000 309.3000 941.4000 326.7000 ;
	    RECT 942.6000 323.4000 943.8000 324.6000 ;
	    RECT 916.2000 278.4000 917.4000 279.6000 ;
	    RECT 909.0000 227.4000 910.2000 228.6000 ;
	    RECT 909.0000 200.4000 910.2000 201.6000 ;
	    RECT 911.4000 200.4000 912.6000 201.6000 ;
	    RECT 909.1500 186.6000 910.0500 200.4000 ;
	    RECT 911.5500 198.6000 912.4500 200.4000 ;
	    RECT 911.4000 197.4000 912.6000 198.6000 ;
	    RECT 916.3500 192.6000 917.2500 278.4000 ;
	    RECT 925.8000 233.4000 927.0000 234.6000 ;
	    RECT 921.0000 200.4000 922.2000 201.6000 ;
	    RECT 916.2000 191.4000 917.4000 192.6000 ;
	    RECT 909.0000 185.4000 910.2000 186.6000 ;
	    RECT 909.1500 180.6000 910.0500 185.4000 ;
	    RECT 921.1500 180.6000 922.0500 200.4000 ;
	    RECT 909.0000 179.4000 910.2000 180.6000 ;
	    RECT 921.0000 179.4000 922.2000 180.6000 ;
	    RECT 921.1500 168.6000 922.0500 179.4000 ;
	    RECT 921.0000 167.4000 922.2000 168.6000 ;
	    RECT 925.9500 165.6000 926.8500 233.4000 ;
	    RECT 930.6000 230.4000 931.8000 231.6000 ;
	    RECT 930.7500 228.6000 931.6500 230.4000 ;
	    RECT 930.6000 227.4000 931.8000 228.6000 ;
	    RECT 928.2000 221.4000 929.4000 222.6000 ;
	    RECT 928.3500 216.6000 929.2500 221.4000 ;
	    RECT 928.2000 215.4000 929.4000 216.6000 ;
	    RECT 940.2000 209.4000 941.4000 210.6000 ;
	    RECT 930.6000 203.4000 931.8000 204.6000 ;
	    RECT 930.7500 180.6000 931.6500 203.4000 ;
	    RECT 940.3500 195.6000 941.2500 209.4000 ;
	    RECT 940.2000 194.4000 941.4000 195.6000 ;
	    RECT 942.7500 192.6000 943.6500 323.4000 ;
	    RECT 945.0000 309.3000 946.2000 326.7000 ;
	    RECT 947.4000 320.4000 948.6000 321.6000 ;
	    RECT 947.5500 318.6000 948.4500 320.4000 ;
	    RECT 947.4000 317.4000 948.6000 318.6000 ;
	    RECT 949.8000 309.3000 951.0000 326.7000 ;
	    RECT 952.2000 306.3000 953.4000 326.7000 ;
	    RECT 954.6000 306.3000 955.8000 326.7000 ;
	    RECT 957.1500 318.6000 958.0500 365.4000 ;
	    RECT 969.1500 318.6000 970.0500 383.4000 ;
	    RECT 971.5500 378.6000 972.4500 398.4000 ;
	    RECT 973.8000 396.3000 975.0000 413.7000 ;
	    RECT 976.2000 396.3000 977.4000 416.7000 ;
	    RECT 978.6000 396.3000 979.8000 416.7000 ;
	    RECT 981.0000 396.3000 982.2000 416.7000 ;
	    RECT 983.4000 389.4000 984.6000 390.6000 ;
	    RECT 971.4000 377.4000 972.6000 378.6000 ;
	    RECT 981.0000 329.4000 982.2000 330.6000 ;
	    RECT 957.0000 317.4000 958.2000 318.6000 ;
	    RECT 969.0000 317.4000 970.2000 318.6000 ;
	    RECT 957.1500 246.6000 958.0500 317.4000 ;
	    RECT 961.8000 314.4000 963.0000 315.6000 ;
	    RECT 961.9500 312.6000 962.8500 314.4000 ;
	    RECT 961.8000 311.4000 963.0000 312.6000 ;
	    RECT 961.9500 306.6000 962.8500 311.4000 ;
	    RECT 961.8000 305.4000 963.0000 306.6000 ;
	    RECT 971.4000 305.4000 972.6000 306.6000 ;
	    RECT 969.0000 287.4000 970.2000 288.6000 ;
	    RECT 969.1500 285.6000 970.0500 287.4000 ;
	    RECT 969.0000 284.4000 970.2000 285.6000 ;
	    RECT 969.0000 248.4000 970.2000 249.6000 ;
	    RECT 957.0000 245.4000 958.2000 246.6000 ;
	    RECT 945.0000 216.3000 946.2000 236.7000 ;
	    RECT 947.4000 216.3000 948.6000 236.7000 ;
	    RECT 949.8000 216.3000 951.0000 236.7000 ;
	    RECT 952.2000 216.3000 953.4000 233.7000 ;
	    RECT 954.6000 218.4000 955.8000 219.6000 ;
	    RECT 954.7500 192.6000 955.6500 218.4000 ;
	    RECT 957.0000 216.3000 958.2000 233.7000 ;
	    RECT 959.4000 221.4000 960.6000 222.6000 ;
	    RECT 959.5500 216.6000 960.4500 221.4000 ;
	    RECT 959.4000 215.4000 960.6000 216.6000 ;
	    RECT 961.8000 216.3000 963.0000 233.7000 ;
	    RECT 964.2000 216.3000 965.4000 236.7000 ;
	    RECT 966.6000 216.3000 967.8000 236.7000 ;
	    RECT 969.1500 225.6000 970.0500 248.4000 ;
	    RECT 969.0000 224.4000 970.2000 225.6000 ;
	    RECT 969.0000 201.4500 970.2000 201.6000 ;
	    RECT 971.5500 201.4500 972.4500 305.4000 ;
	    RECT 976.2000 276.3000 977.4000 293.7000 ;
	    RECT 973.8000 236.4000 975.0000 237.6000 ;
	    RECT 973.9500 228.6000 974.8500 236.4000 ;
	    RECT 973.8000 227.4000 975.0000 228.6000 ;
	    RECT 969.0000 200.5500 972.4500 201.4500 ;
	    RECT 969.0000 200.4000 970.2000 200.5500 ;
	    RECT 959.4000 197.4000 960.6000 198.6000 ;
	    RECT 961.8000 197.4000 963.0000 198.6000 ;
	    RECT 966.6000 197.4000 967.8000 198.6000 ;
	    RECT 940.2000 191.4000 941.4000 192.6000 ;
	    RECT 942.6000 191.4000 943.8000 192.6000 ;
	    RECT 954.6000 191.4000 955.8000 192.6000 ;
	    RECT 930.6000 179.4000 931.8000 180.6000 ;
	    RECT 925.8000 164.4000 927.0000 165.6000 ;
	    RECT 928.2000 156.3000 929.4000 176.7000 ;
	    RECT 930.6000 156.3000 931.8000 176.7000 ;
	    RECT 933.0000 156.3000 934.2000 173.7000 ;
	    RECT 935.4000 161.4000 936.6000 162.6000 ;
	    RECT 935.5500 156.6000 936.4500 161.4000 ;
	    RECT 935.4000 155.4000 936.6000 156.6000 ;
	    RECT 937.8000 156.3000 939.0000 173.7000 ;
	    RECT 940.3500 159.6000 941.2500 191.4000 ;
	    RECT 940.2000 158.4000 941.4000 159.6000 ;
	    RECT 906.6000 149.4000 907.8000 150.6000 ;
	    RECT 935.4000 143.4000 936.6000 144.6000 ;
	    RECT 861.0000 140.4000 862.2000 141.6000 ;
	    RECT 861.1500 138.6000 862.0500 140.4000 ;
	    RECT 861.0000 137.4000 862.2000 138.6000 ;
	    RECT 868.2000 137.4000 869.4000 138.6000 ;
	    RECT 858.6000 135.4500 859.8000 135.6000 ;
	    RECT 856.3500 134.5500 859.8000 135.4500 ;
	    RECT 858.6000 134.4000 859.8000 134.5500 ;
	    RECT 868.3500 126.6000 869.2500 137.4000 ;
	    RECT 868.2000 125.4000 869.4000 126.6000 ;
	    RECT 815.4000 119.4000 816.6000 120.6000 ;
	    RECT 822.6000 119.4000 823.8000 120.6000 ;
	    RECT 935.5500 114.6000 936.4500 143.4000 ;
	    RECT 940.3500 129.4500 941.2500 158.4000 ;
	    RECT 942.6000 156.3000 943.8000 173.7000 ;
	    RECT 945.0000 156.3000 946.2000 176.7000 ;
	    RECT 947.4000 156.3000 948.6000 176.7000 ;
	    RECT 949.8000 156.3000 951.0000 176.7000 ;
	    RECT 959.5500 174.6000 960.4500 197.4000 ;
	    RECT 966.7500 192.6000 967.6500 197.4000 ;
	    RECT 966.6000 191.4000 967.8000 192.6000 ;
	    RECT 964.2000 179.4000 965.4000 180.6000 ;
	    RECT 959.4000 173.4000 960.6000 174.6000 ;
	    RECT 964.3500 171.6000 965.2500 179.4000 ;
	    RECT 964.2000 170.4000 965.4000 171.6000 ;
	    RECT 969.1500 156.6000 970.0500 200.4000 ;
	    RECT 978.6000 170.4000 979.8000 171.6000 ;
	    RECT 969.0000 156.4500 970.2000 156.6000 ;
	    RECT 969.0000 155.5500 972.4500 156.4500 ;
	    RECT 969.0000 155.4000 970.2000 155.5500 ;
	    RECT 959.4000 137.4000 960.6000 138.6000 ;
	    RECT 940.3500 128.5500 943.6500 129.4500 ;
	    RECT 940.2000 116.4000 941.4000 117.6000 ;
	    RECT 851.4000 113.4000 852.6000 114.6000 ;
	    RECT 935.4000 113.4000 936.6000 114.6000 ;
	    RECT 851.5500 81.6000 852.4500 113.4000 ;
	    RECT 851.4000 80.4000 852.6000 81.6000 ;
	    RECT 808.2000 77.4000 809.4000 78.6000 ;
	    RECT 935.5500 75.6000 936.4500 113.4000 ;
	    RECT 940.3500 108.6000 941.2500 116.4000 ;
	    RECT 940.2000 107.4000 941.4000 108.6000 ;
	    RECT 942.7500 78.6000 943.6500 128.5500 ;
	    RECT 954.6000 125.4000 955.8000 126.6000 ;
	    RECT 945.0000 107.4000 946.2000 108.6000 ;
	    RECT 945.1500 105.6000 946.0500 107.4000 ;
	    RECT 945.0000 104.4000 946.2000 105.6000 ;
	    RECT 947.4000 96.3000 948.6000 116.7000 ;
	    RECT 949.8000 96.3000 951.0000 116.7000 ;
	    RECT 952.2000 96.3000 953.4000 113.7000 ;
	    RECT 954.7500 102.6000 955.6500 125.4000 ;
	    RECT 959.5500 120.6000 960.4500 137.4000 ;
	    RECT 959.4000 119.4000 960.6000 120.6000 ;
	    RECT 954.6000 101.4000 955.8000 102.6000 ;
	    RECT 957.0000 96.3000 958.2000 113.7000 ;
	    RECT 959.5500 99.6000 960.4500 119.4000 ;
	    RECT 959.4000 98.4000 960.6000 99.6000 ;
	    RECT 961.8000 96.3000 963.0000 113.7000 ;
	    RECT 964.2000 96.3000 965.4000 116.7000 ;
	    RECT 966.6000 96.3000 967.8000 116.7000 ;
	    RECT 969.0000 96.3000 970.2000 116.7000 ;
	    RECT 971.5500 81.6000 972.4500 155.5500 ;
	    RECT 973.8000 125.4000 975.0000 126.6000 ;
	    RECT 973.9500 81.6000 974.8500 125.4000 ;
	    RECT 971.4000 80.4000 972.6000 81.6000 ;
	    RECT 973.8000 80.4000 975.0000 81.6000 ;
	    RECT 942.6000 77.4000 943.8000 78.6000 ;
	    RECT 947.4000 77.4000 948.6000 78.6000 ;
	    RECT 964.2000 77.4000 965.4000 78.6000 ;
	    RECT 935.4000 74.4000 936.6000 75.6000 ;
	    RECT 832.2000 59.4000 833.4000 60.6000 ;
	    RECT 839.4000 59.4000 840.6000 60.6000 ;
	    RECT 856.2000 59.4000 857.4000 60.6000 ;
	    RECT 769.8000 47.4000 771.0000 48.6000 ;
	    RECT 774.6000 47.4000 775.8000 48.6000 ;
	    RECT 793.8000 47.4000 795.0000 48.6000 ;
	    RECT 765.0000 44.4000 766.2000 45.6000 ;
	    RECT 760.2000 41.4000 761.4000 42.6000 ;
	    RECT 755.4000 35.4000 756.6000 36.6000 ;
	    RECT 585.0000 29.4000 586.2000 30.6000 ;
	    RECT 726.6000 29.4000 727.8000 30.6000 ;
	    RECT 755.5500 30.4500 756.4500 35.4000 ;
	    RECT 765.1500 30.6000 766.0500 44.4000 ;
	    RECT 769.9500 42.6000 770.8500 47.4000 ;
	    RECT 769.8000 41.4000 771.0000 42.6000 ;
	    RECT 772.2000 41.4000 773.4000 42.6000 ;
	    RECT 753.1500 29.5500 756.4500 30.4500 ;
	    RECT 585.1500 24.6000 586.0500 29.4000 ;
	    RECT 577.8000 23.4000 579.0000 24.6000 ;
	    RECT 582.6000 23.4000 583.8000 24.6000 ;
	    RECT 585.0000 23.4000 586.2000 24.6000 ;
	    RECT 726.7500 21.6000 727.6500 29.4000 ;
	    RECT 563.4000 20.4000 564.6000 21.6000 ;
	    RECT 594.6000 20.4000 595.8000 21.6000 ;
	    RECT 726.6000 20.4000 727.8000 21.6000 ;
	    RECT 594.7500 18.6000 595.6500 20.4000 ;
	    RECT 594.6000 17.4000 595.8000 18.6000 ;
	    RECT 738.6000 17.4000 739.8000 18.6000 ;
	    RECT 534.6000 14.4000 535.8000 15.6000 ;
	    RECT 558.6000 14.4000 559.8000 15.6000 ;
	    RECT 733.8000 14.4000 735.0000 15.6000 ;
	    RECT 529.8000 11.4000 531.0000 12.6000 ;
	    RECT 534.7500 6.6000 535.6500 14.4000 ;
	    RECT 733.9500 6.6000 734.8500 14.4000 ;
	    RECT 534.6000 5.4000 535.8000 6.6000 ;
	    RECT 733.8000 5.4000 735.0000 6.6000 ;
	    RECT 741.0000 6.3000 742.2000 26.7000 ;
	    RECT 743.4000 6.3000 744.6000 26.7000 ;
	    RECT 745.8000 9.3000 747.0000 26.7000 ;
	    RECT 748.2000 23.4000 749.4000 24.6000 ;
	    RECT 748.3500 21.6000 749.2500 23.4000 ;
	    RECT 748.2000 20.4000 749.4000 21.6000 ;
	    RECT 750.6000 9.3000 751.8000 26.7000 ;
	    RECT 753.1500 24.6000 754.0500 29.5500 ;
	    RECT 765.0000 29.4000 766.2000 30.6000 ;
	    RECT 753.0000 23.4000 754.2000 24.6000 ;
	    RECT 755.4000 9.3000 756.6000 26.7000 ;
	    RECT 757.8000 6.3000 759.0000 26.7000 ;
	    RECT 760.2000 6.3000 761.4000 26.7000 ;
	    RECT 762.6000 6.3000 763.8000 26.7000 ;
	    RECT 772.3500 24.6000 773.2500 41.4000 ;
	    RECT 774.7500 30.6000 775.6500 47.4000 ;
	    RECT 798.6000 44.4000 799.8000 45.6000 ;
	    RECT 774.6000 29.4000 775.8000 30.6000 ;
	    RECT 772.2000 23.4000 773.4000 24.6000 ;
	    RECT 796.2000 23.4000 797.4000 24.6000 ;
	    RECT 796.3500 12.6000 797.2500 23.4000 ;
	    RECT 798.7500 21.6000 799.6500 44.4000 ;
	    RECT 832.3500 42.6000 833.2500 59.4000 ;
	    RECT 832.2000 41.4000 833.4000 42.6000 ;
	    RECT 801.0000 29.4000 802.2000 30.6000 ;
	    RECT 798.6000 20.4000 799.8000 21.6000 ;
	    RECT 801.1500 18.6000 802.0500 29.4000 ;
	    RECT 839.5500 21.6000 840.4500 59.4000 ;
	    RECT 856.3500 51.6000 857.2500 59.4000 ;
	    RECT 885.0000 56.4000 886.2000 57.6000 ;
	    RECT 856.2000 50.4000 857.4000 51.6000 ;
	    RECT 856.3500 24.6000 857.2500 50.4000 ;
	    RECT 856.2000 23.4000 857.4000 24.6000 ;
	    RECT 885.1500 21.6000 886.0500 56.4000 ;
	    RECT 947.5500 42.6000 948.4500 77.4000 ;
	    RECT 947.4000 41.4000 948.6000 42.6000 ;
	    RECT 949.8000 36.3000 951.0000 56.7000 ;
	    RECT 952.2000 36.3000 953.4000 56.7000 ;
	    RECT 954.6000 36.3000 955.8000 56.7000 ;
	    RECT 964.3500 54.6000 965.2500 77.4000 ;
	    RECT 978.7500 75.6000 979.6500 170.4000 ;
	    RECT 981.1500 120.6000 982.0500 329.4000 ;
	    RECT 983.5500 171.6000 984.4500 389.4000 ;
	    RECT 985.8000 299.4000 987.0000 300.6000 ;
	    RECT 985.9500 285.6000 986.8500 299.4000 ;
	    RECT 985.8000 284.4000 987.0000 285.6000 ;
	    RECT 988.3500 249.6000 989.2500 533.4000 ;
	    RECT 990.6000 467.4000 991.8000 468.6000 ;
	    RECT 990.7500 465.6000 991.6500 467.4000 ;
	    RECT 990.6000 464.4000 991.8000 465.6000 ;
	    RECT 993.1500 444.6000 994.0500 557.4000 ;
	    RECT 995.4000 516.3000 996.6000 533.7000 ;
	    RECT 995.4000 467.4000 996.6000 468.6000 ;
	    RECT 993.0000 443.4000 994.2000 444.6000 ;
	    RECT 995.5500 411.6000 996.4500 467.4000 ;
	    RECT 995.4000 410.4000 996.6000 411.6000 ;
	    RECT 990.6000 377.4000 991.8000 378.6000 ;
	    RECT 990.7500 366.6000 991.6500 377.4000 ;
	    RECT 990.6000 365.4000 991.8000 366.6000 ;
	    RECT 990.7500 309.4500 991.6500 365.4000 ;
	    RECT 997.8000 323.4000 999.0000 324.6000 ;
	    RECT 997.9500 318.6000 998.8500 323.4000 ;
	    RECT 1000.3500 321.6000 1001.2500 629.4000 ;
	    RECT 1007.5500 582.6000 1008.4500 671.4000 ;
	    RECT 1007.4000 581.4000 1008.6000 582.6000 ;
	    RECT 1002.6000 554.4000 1003.8000 555.6000 ;
	    RECT 1002.7500 525.6000 1003.6500 554.4000 ;
	    RECT 1002.6000 524.4000 1003.8000 525.6000 ;
	    RECT 1005.0000 440.4000 1006.2000 441.6000 ;
	    RECT 1005.1500 321.6000 1006.0500 440.4000 ;
	    RECT 1009.9500 402.6000 1010.8500 680.4000 ;
	    RECT 1019.5500 654.6000 1020.4500 956.4000 ;
	    RECT 1024.3500 834.6000 1025.2500 959.4000 ;
	    RECT 1033.9501 957.6000 1034.8500 1205.4000 ;
	    RECT 1036.3500 1089.4501 1037.2500 1229.4000 ;
	    RECT 1038.6000 1223.4000 1039.8000 1224.6000 ;
	    RECT 1038.7500 1200.6000 1039.6500 1223.4000 ;
	    RECT 1038.6000 1199.4000 1039.8000 1200.6000 ;
	    RECT 1043.5500 1188.6000 1044.4501 1457.4000 ;
	    RECT 1069.8000 1451.4000 1071.0000 1452.6000 ;
	    RECT 1067.4000 1439.4000 1068.6000 1440.6000 ;
	    RECT 1057.8000 1427.4000 1059.0000 1428.6000 ;
	    RECT 1057.9501 1401.6000 1058.8500 1427.4000 ;
	    RECT 1067.5500 1401.6000 1068.4501 1439.4000 ;
	    RECT 1069.9501 1404.6000 1070.8500 1451.4000 ;
	    RECT 1086.6000 1446.3000 1087.8000 1466.7001 ;
	    RECT 1089.0000 1446.3000 1090.2001 1466.7001 ;
	    RECT 1091.4000 1446.3000 1092.6000 1466.7001 ;
	    RECT 1093.8000 1449.3000 1095.0000 1466.7001 ;
	    RECT 1096.2001 1463.4000 1097.4000 1464.6000 ;
	    RECT 1098.6000 1449.3000 1099.8000 1466.7001 ;
	    RECT 1101.0000 1460.4000 1102.2001 1461.6000 ;
	    RECT 1101.1500 1452.6000 1102.0500 1460.4000 ;
	    RECT 1101.0000 1451.4000 1102.2001 1452.6000 ;
	    RECT 1103.4000 1449.3000 1104.6000 1466.7001 ;
	    RECT 1096.2001 1445.4000 1097.4000 1446.6000 ;
	    RECT 1105.8000 1446.3000 1107.0000 1466.7001 ;
	    RECT 1108.2001 1446.3000 1109.4000 1466.7001 ;
	    RECT 1139.4000 1463.4000 1140.6000 1464.6000 ;
	    RECT 1199.4000 1463.4000 1200.6000 1464.6000 ;
	    RECT 1312.2001 1463.4000 1313.4000 1464.6000 ;
	    RECT 1333.8000 1463.4000 1335.0000 1464.6000 ;
	    RECT 1446.6000 1463.4000 1447.8000 1464.6000 ;
	    RECT 1110.6000 1457.4000 1111.8000 1458.6000 ;
	    RECT 1115.4000 1454.4000 1116.6000 1455.6000 ;
	    RECT 1110.6000 1451.4000 1111.8000 1452.6000 ;
	    RECT 1072.2001 1416.3000 1073.4000 1436.7001 ;
	    RECT 1074.6000 1416.3000 1075.8000 1436.7001 ;
	    RECT 1077.0000 1416.3000 1078.2001 1436.7001 ;
	    RECT 1079.4000 1416.3000 1080.6000 1433.7001 ;
	    RECT 1081.8000 1418.4000 1083.0000 1419.6000 ;
	    RECT 1069.8000 1403.4000 1071.0000 1404.6000 ;
	    RECT 1055.4000 1400.4000 1056.6000 1401.6000 ;
	    RECT 1057.8000 1400.4000 1059.0000 1401.6000 ;
	    RECT 1067.4000 1400.4000 1068.6000 1401.6000 ;
	    RECT 1055.5500 1398.6000 1056.4501 1400.4000 ;
	    RECT 1055.4000 1397.4000 1056.6000 1398.6000 ;
	    RECT 1062.6000 1397.4000 1063.8000 1398.6000 ;
	    RECT 1065.0000 1397.4000 1066.2001 1398.6000 ;
	    RECT 1057.8000 1394.4000 1059.0000 1395.6000 ;
	    RECT 1057.9501 1392.6000 1058.8500 1394.4000 ;
	    RECT 1065.1500 1392.6000 1066.0500 1397.4000 ;
	    RECT 1057.8000 1391.4000 1059.0000 1392.6000 ;
	    RECT 1065.0000 1391.4000 1066.2001 1392.6000 ;
	    RECT 1048.2001 1310.4000 1049.4000 1311.6000 ;
	    RECT 1048.3500 1302.6000 1049.2500 1310.4000 ;
	    RECT 1045.8000 1301.4000 1047.0000 1302.6000 ;
	    RECT 1048.2001 1301.4000 1049.4000 1302.6000 ;
	    RECT 1045.9501 1281.6000 1046.8500 1301.4000 ;
	    RECT 1048.3500 1299.6000 1049.2500 1301.4000 ;
	    RECT 1048.2001 1298.4000 1049.4000 1299.6000 ;
	    RECT 1053.0000 1283.4000 1054.2001 1284.6000 ;
	    RECT 1053.1500 1281.6000 1054.0500 1283.4000 ;
	    RECT 1045.8000 1280.4000 1047.0000 1281.6000 ;
	    RECT 1053.0000 1280.4000 1054.2001 1281.6000 ;
	    RECT 1050.6000 1277.4000 1051.8000 1278.6000 ;
	    RECT 1055.4000 1277.4000 1056.6000 1278.6000 ;
	    RECT 1043.4000 1187.4000 1044.6000 1188.6000 ;
	    RECT 1043.5500 1167.6000 1044.4501 1187.4000 ;
	    RECT 1043.4000 1166.4000 1044.6000 1167.6000 ;
	    RECT 1043.4000 1145.4000 1044.6000 1146.6000 ;
	    RECT 1041.0000 1133.4000 1042.2001 1134.6000 ;
	    RECT 1041.1500 1125.6000 1042.0500 1133.4000 ;
	    RECT 1041.0000 1124.4000 1042.2001 1125.6000 ;
	    RECT 1043.5500 1122.6000 1044.4501 1145.4000 ;
	    RECT 1045.8000 1127.4000 1047.0000 1128.6000 ;
	    RECT 1045.9501 1125.6000 1046.8500 1127.4000 ;
	    RECT 1045.8000 1124.4000 1047.0000 1125.6000 ;
	    RECT 1048.2001 1124.4000 1049.4000 1125.6000 ;
	    RECT 1038.6000 1122.4501 1039.8000 1122.6000 ;
	    RECT 1038.6000 1121.5500 1042.0500 1122.4501 ;
	    RECT 1038.6000 1121.4000 1039.8000 1121.5500 ;
	    RECT 1041.1500 1119.4501 1042.0500 1121.5500 ;
	    RECT 1043.4000 1121.4000 1044.6000 1122.6000 ;
	    RECT 1048.3500 1122.4501 1049.2500 1124.4000 ;
	    RECT 1045.9501 1121.5500 1049.2500 1122.4501 ;
	    RECT 1045.9501 1119.4501 1046.8500 1121.5500 ;
	    RECT 1050.7500 1119.4501 1051.6500 1277.4000 ;
	    RECT 1055.5500 1257.6000 1056.4501 1277.4000 ;
	    RECT 1055.4000 1256.4000 1056.6000 1257.6000 ;
	    RECT 1053.0000 1220.4000 1054.2001 1221.6000 ;
	    RECT 1053.1500 1131.6000 1054.0500 1220.4000 ;
	    RECT 1053.0000 1130.4000 1054.2001 1131.6000 ;
	    RECT 1053.0000 1127.4000 1054.2001 1128.6000 ;
	    RECT 1053.1500 1125.6000 1054.0500 1127.4000 ;
	    RECT 1053.0000 1124.4000 1054.2001 1125.6000 ;
	    RECT 1055.5500 1122.4501 1056.4501 1256.4000 ;
	    RECT 1069.9501 1254.6000 1070.8500 1403.4000 ;
	    RECT 1074.6000 1334.4000 1075.8000 1335.6000 ;
	    RECT 1072.2001 1295.4000 1073.4000 1296.6000 ;
	    RECT 1074.7500 1284.6000 1075.6500 1334.4000 ;
	    RECT 1081.9501 1287.6000 1082.8500 1418.4000 ;
	    RECT 1084.2001 1416.3000 1085.4000 1433.7001 ;
	    RECT 1086.6000 1427.4000 1087.8000 1428.6000 ;
	    RECT 1086.7500 1422.6000 1087.6500 1427.4000 ;
	    RECT 1086.6000 1421.4000 1087.8000 1422.6000 ;
	    RECT 1089.0000 1416.3000 1090.2001 1433.7001 ;
	    RECT 1091.4000 1416.3000 1092.6000 1436.7001 ;
	    RECT 1093.8000 1416.3000 1095.0000 1436.7001 ;
	    RECT 1096.3500 1425.6000 1097.2500 1445.4000 ;
	    RECT 1101.0000 1439.4000 1102.2001 1440.6000 ;
	    RECT 1101.1500 1428.6000 1102.0500 1439.4000 ;
	    RECT 1101.0000 1427.4000 1102.2001 1428.6000 ;
	    RECT 1096.2001 1424.4000 1097.4000 1425.6000 ;
	    RECT 1091.4000 1403.4000 1092.6000 1404.6000 ;
	    RECT 1084.2001 1400.4000 1085.4000 1401.6000 ;
	    RECT 1084.3500 1380.6000 1085.2500 1400.4000 ;
	    RECT 1089.0000 1394.4000 1090.2001 1395.6000 ;
	    RECT 1084.2001 1379.4000 1085.4000 1380.6000 ;
	    RECT 1081.8000 1286.4000 1083.0000 1287.6000 ;
	    RECT 1074.6000 1283.4000 1075.8000 1284.6000 ;
	    RECT 1069.8000 1253.4000 1071.0000 1254.6000 ;
	    RECT 1057.8000 1223.4000 1059.0000 1224.6000 ;
	    RECT 1060.2001 1223.4000 1061.4000 1224.6000 ;
	    RECT 1069.8000 1223.4000 1071.0000 1224.6000 ;
	    RECT 1057.9501 1212.6000 1058.8500 1223.4000 ;
	    RECT 1060.3500 1221.6000 1061.2500 1223.4000 ;
	    RECT 1060.2001 1220.4000 1061.4000 1221.6000 ;
	    RECT 1057.8000 1211.4000 1059.0000 1212.6000 ;
	    RECT 1074.7500 1206.6000 1075.6500 1283.4000 ;
	    RECT 1084.2001 1271.4000 1085.4000 1272.6000 ;
	    RECT 1084.3500 1230.6000 1085.2500 1271.4000 ;
	    RECT 1084.2001 1229.4000 1085.4000 1230.6000 ;
	    RECT 1084.3500 1224.6000 1085.2500 1229.4000 ;
	    RECT 1084.2001 1223.4000 1085.4000 1224.6000 ;
	    RECT 1074.6000 1205.4000 1075.8000 1206.6000 ;
	    RECT 1079.4000 1199.4000 1080.6000 1200.6000 ;
	    RECT 1079.5500 1194.6000 1080.4501 1199.4000 ;
	    RECT 1089.1500 1194.6000 1090.0500 1394.4000 ;
	    RECT 1096.3500 1368.6000 1097.2500 1424.4000 ;
	    RECT 1110.7500 1422.6000 1111.6500 1451.4000 ;
	    RECT 1115.5500 1446.6000 1116.4501 1454.4000 ;
	    RECT 1115.4000 1445.4000 1116.6000 1446.6000 ;
	    RECT 1137.0000 1427.4000 1138.2001 1428.6000 ;
	    RECT 1110.6000 1421.4000 1111.8000 1422.6000 ;
	    RECT 1122.6000 1421.4000 1123.8000 1422.6000 ;
	    RECT 1122.7500 1401.6000 1123.6500 1421.4000 ;
	    RECT 1122.6000 1400.4000 1123.8000 1401.6000 ;
	    RECT 1127.4000 1400.4000 1128.6000 1401.6000 ;
	    RECT 1120.2001 1394.4000 1121.4000 1395.6000 ;
	    RECT 1120.3500 1380.6000 1121.2500 1394.4000 ;
	    RECT 1127.5500 1392.6000 1128.4501 1400.4000 ;
	    RECT 1137.1500 1398.6000 1138.0500 1427.4000 ;
	    RECT 1139.5500 1404.6000 1140.4501 1463.4000 ;
	    RECT 1146.6000 1460.4000 1147.8000 1461.6000 ;
	    RECT 1177.8000 1460.4000 1179.0000 1461.6000 ;
	    RECT 1185.0000 1460.4000 1186.2001 1461.6000 ;
	    RECT 1146.7500 1440.4501 1147.6500 1460.4000 ;
	    RECT 1149.0000 1440.4501 1150.2001 1440.6000 ;
	    RECT 1146.7500 1439.5500 1150.2001 1440.4501 ;
	    RECT 1149.0000 1439.4000 1150.2001 1439.5500 ;
	    RECT 1149.1500 1437.6000 1150.0500 1439.4000 ;
	    RECT 1149.0000 1436.4000 1150.2001 1437.6000 ;
	    RECT 1144.2001 1424.4000 1145.4000 1425.6000 ;
	    RECT 1144.3500 1422.6000 1145.2500 1424.4000 ;
	    RECT 1149.1500 1422.6000 1150.0500 1436.4000 ;
	    RECT 1177.9501 1428.6000 1178.8500 1460.4000 ;
	    RECT 1185.1500 1437.6000 1186.0500 1460.4000 ;
	    RECT 1185.0000 1436.4000 1186.2001 1437.6000 ;
	    RECT 1199.5500 1431.6000 1200.4501 1463.4000 ;
	    RECT 1252.2001 1460.4000 1253.4000 1461.6000 ;
	    RECT 1199.4000 1430.4000 1200.6000 1431.6000 ;
	    RECT 1177.8000 1427.4000 1179.0000 1428.6000 ;
	    RECT 1144.2001 1421.4000 1145.4000 1422.6000 ;
	    RECT 1149.0000 1421.4000 1150.2001 1422.6000 ;
	    RECT 1139.4000 1403.4000 1140.6000 1404.6000 ;
	    RECT 1137.0000 1397.4000 1138.2001 1398.6000 ;
	    RECT 1127.4000 1391.4000 1128.6000 1392.6000 ;
	    RECT 1127.5500 1386.6000 1128.4501 1391.4000 ;
	    RECT 1127.4000 1385.4000 1128.6000 1386.6000 ;
	    RECT 1120.2001 1379.4000 1121.4000 1380.6000 ;
	    RECT 1120.3500 1368.6000 1121.2500 1379.4000 ;
	    RECT 1096.2001 1367.4000 1097.4000 1368.6000 ;
	    RECT 1120.2001 1367.4000 1121.4000 1368.6000 ;
	    RECT 1125.0000 1367.4000 1126.2001 1368.6000 ;
	    RECT 1074.6000 1193.4000 1075.8000 1194.6000 ;
	    RECT 1079.4000 1193.4000 1080.6000 1194.6000 ;
	    RECT 1072.2001 1181.4000 1073.4000 1182.6000 ;
	    RECT 1057.8000 1145.4000 1059.0000 1146.6000 ;
	    RECT 1062.6000 1146.3000 1063.8000 1166.7001 ;
	    RECT 1065.0000 1146.3000 1066.2001 1166.7001 ;
	    RECT 1067.4000 1146.3000 1068.6000 1166.7001 ;
	    RECT 1069.8000 1149.3000 1071.0000 1166.7001 ;
	    RECT 1072.3500 1164.6000 1073.2500 1181.4000 ;
	    RECT 1074.7500 1170.4501 1075.6500 1193.4000 ;
	    RECT 1079.4000 1187.4000 1080.6000 1188.6000 ;
	    RECT 1081.8000 1179.3000 1083.0000 1187.7001 ;
	    RECT 1084.2001 1181.4000 1085.4000 1182.6000 ;
	    RECT 1084.3500 1176.6000 1085.2500 1181.4000 ;
	    RECT 1084.2001 1175.4000 1085.4000 1176.6000 ;
	    RECT 1086.6000 1176.3000 1087.8000 1193.7001 ;
	    RECT 1089.0000 1193.4000 1090.2001 1194.6000 ;
	    RECT 1093.8000 1184.4000 1095.0000 1185.6000 ;
	    RECT 1074.7500 1169.5500 1078.0500 1170.4501 ;
	    RECT 1072.2001 1163.4000 1073.4000 1164.6000 ;
	    RECT 1069.8000 1145.4000 1071.0000 1146.6000 ;
	    RECT 1041.1500 1118.5500 1046.8500 1119.4501 ;
	    RECT 1048.3500 1118.5500 1051.6500 1119.4501 ;
	    RECT 1053.1500 1121.5500 1056.4501 1122.4501 ;
	    RECT 1043.4000 1103.4000 1044.6000 1104.6000 ;
	    RECT 1036.3500 1088.5500 1039.6500 1089.4501 ;
	    RECT 1036.2001 1085.4000 1037.4000 1086.6000 ;
	    RECT 1036.3500 1044.6000 1037.2500 1085.4000 ;
	    RECT 1036.2001 1043.4000 1037.4000 1044.6000 ;
	    RECT 1036.2001 1037.4000 1037.4000 1038.6000 ;
	    RECT 1036.3500 1020.6000 1037.2500 1037.4000 ;
	    RECT 1036.2001 1019.4000 1037.4000 1020.6000 ;
	    RECT 1038.7500 1008.6000 1039.6500 1088.5500 ;
	    RECT 1038.6000 1007.4000 1039.8000 1008.6000 ;
	    RECT 1036.2001 1001.4000 1037.4000 1002.6000 ;
	    RECT 1033.8000 956.4000 1035.0000 957.6000 ;
	    RECT 1029.0000 887.4000 1030.2001 888.6000 ;
	    RECT 1029.1500 885.6000 1030.0500 887.4000 ;
	    RECT 1029.0000 884.4000 1030.2001 885.6000 ;
	    RECT 1033.8000 884.4000 1035.0000 885.6000 ;
	    RECT 1033.9501 882.6000 1034.8500 884.4000 ;
	    RECT 1036.3500 882.6000 1037.2500 1001.4000 ;
	    RECT 1038.7500 999.6000 1039.6500 1007.4000 ;
	    RECT 1038.6000 998.4000 1039.8000 999.6000 ;
	    RECT 1043.5500 984.6000 1044.4501 1103.4000 ;
	    RECT 1045.8000 1100.4000 1047.0000 1101.6000 ;
	    RECT 1045.9501 1098.6000 1046.8500 1100.4000 ;
	    RECT 1048.3500 1098.6000 1049.2500 1118.5500 ;
	    RECT 1050.6000 1100.4000 1051.8000 1101.6000 ;
	    RECT 1045.8000 1097.4000 1047.0000 1098.6000 ;
	    RECT 1048.2001 1097.4000 1049.4000 1098.6000 ;
	    RECT 1050.7500 1059.6000 1051.6500 1100.4000 ;
	    RECT 1053.1500 1098.6000 1054.0500 1121.5500 ;
	    RECT 1053.0000 1097.4000 1054.2001 1098.6000 ;
	    RECT 1050.6000 1058.4000 1051.8000 1059.6000 ;
	    RECT 1043.4000 983.4000 1044.6000 984.6000 ;
	    RECT 1043.5500 912.6000 1044.4501 983.4000 ;
	    RECT 1043.4000 911.4000 1044.6000 912.6000 ;
	    RECT 1053.1500 900.4500 1054.0500 1097.4000 ;
	    RECT 1055.4000 1073.4000 1056.6000 1074.6000 ;
	    RECT 1055.5500 1008.6000 1056.4501 1073.4000 ;
	    RECT 1055.4000 1007.4000 1056.6000 1008.6000 ;
	    RECT 1057.9501 1002.4500 1058.8500 1145.4000 ;
	    RECT 1060.2001 1121.4000 1061.4000 1122.6000 ;
	    RECT 1060.3500 1101.6000 1061.2500 1121.4000 ;
	    RECT 1062.6000 1118.4000 1063.8000 1119.6000 ;
	    RECT 1060.2001 1100.4000 1061.4000 1101.6000 ;
	    RECT 1062.7500 1086.6000 1063.6500 1118.4000 ;
	    RECT 1062.6000 1085.4000 1063.8000 1086.6000 ;
	    RECT 1067.4000 1076.4000 1068.6000 1077.6000 ;
	    RECT 1067.5500 1074.6000 1068.4501 1076.4000 ;
	    RECT 1067.4000 1073.4000 1068.6000 1074.6000 ;
	    RECT 1067.5500 1068.6000 1068.4501 1073.4000 ;
	    RECT 1067.4000 1067.4000 1068.6000 1068.6000 ;
	    RECT 1069.9501 1065.4501 1070.8500 1145.4000 ;
	    RECT 1072.3500 1116.6000 1073.2500 1163.4000 ;
	    RECT 1074.6000 1149.3000 1075.8000 1166.7001 ;
	    RECT 1077.1500 1161.6000 1078.0500 1169.5500 ;
	    RECT 1077.0000 1160.4000 1078.2001 1161.6000 ;
	    RECT 1079.4000 1149.3000 1080.6000 1166.7001 ;
	    RECT 1081.8000 1146.3000 1083.0000 1166.7001 ;
	    RECT 1084.2001 1146.3000 1085.4000 1166.7001 ;
	    RECT 1086.6000 1163.4000 1087.8000 1164.6000 ;
	    RECT 1086.7500 1158.6000 1087.6500 1163.4000 ;
	    RECT 1086.6000 1157.4000 1087.8000 1158.6000 ;
	    RECT 1086.7500 1143.4501 1087.6500 1157.4000 ;
	    RECT 1091.4000 1154.4000 1092.6000 1155.6000 ;
	    RECT 1091.5500 1143.6000 1092.4501 1154.4000 ;
	    RECT 1093.9501 1146.6000 1094.8500 1184.4000 ;
	    RECT 1093.8000 1145.4000 1095.0000 1146.6000 ;
	    RECT 1084.3500 1142.5500 1087.6500 1143.4501 ;
	    RECT 1084.3500 1122.6000 1085.2500 1142.5500 ;
	    RECT 1091.4000 1142.4000 1092.6000 1143.6000 ;
	    RECT 1091.5500 1140.6000 1092.4501 1142.4000 ;
	    RECT 1091.4000 1139.4000 1092.6000 1140.6000 ;
	    RECT 1091.5500 1128.6000 1092.4501 1139.4000 ;
	    RECT 1091.4000 1127.4000 1092.6000 1128.6000 ;
	    RECT 1093.8000 1127.4000 1095.0000 1128.6000 ;
	    RECT 1084.2001 1121.4000 1085.4000 1122.6000 ;
	    RECT 1093.9501 1116.6000 1094.8500 1127.4000 ;
	    RECT 1072.2001 1115.4000 1073.4000 1116.6000 ;
	    RECT 1093.8000 1115.4000 1095.0000 1116.6000 ;
	    RECT 1096.3500 1080.6000 1097.2500 1367.4000 ;
	    RECT 1125.1500 1365.6000 1126.0500 1367.4000 ;
	    RECT 1125.0000 1364.4000 1126.2001 1365.6000 ;
	    RECT 1125.0000 1355.4000 1126.2001 1356.6000 ;
	    RECT 1127.4000 1356.3000 1128.6000 1376.7001 ;
	    RECT 1129.8000 1356.3000 1131.0000 1376.7001 ;
	    RECT 1132.2001 1356.3000 1133.4000 1373.7001 ;
	    RECT 1134.6000 1361.4000 1135.8000 1362.6000 ;
	    RECT 1134.7500 1356.6000 1135.6500 1361.4000 ;
	    RECT 1134.6000 1355.4000 1135.8000 1356.6000 ;
	    RECT 1137.0000 1356.3000 1138.2001 1373.7001 ;
	    RECT 1139.5500 1359.6000 1140.4501 1403.4000 ;
	    RECT 1139.4000 1358.4000 1140.6000 1359.6000 ;
	    RECT 1141.8000 1356.3000 1143.0000 1373.7001 ;
	    RECT 1144.2001 1356.3000 1145.4000 1376.7001 ;
	    RECT 1146.6000 1356.3000 1147.8000 1376.7001 ;
	    RECT 1149.0000 1356.3000 1150.2001 1376.7001 ;
	    RECT 1163.4000 1370.4000 1164.6000 1371.6000 ;
	    RECT 1235.4000 1370.4000 1236.6000 1371.6000 ;
	    RECT 1125.1500 1332.6000 1126.0500 1355.4000 ;
	    RECT 1125.0000 1331.4000 1126.2001 1332.6000 ;
	    RECT 1134.6000 1301.4000 1135.8000 1302.6000 ;
	    RECT 1108.2001 1286.4000 1109.4000 1287.6000 ;
	    RECT 1098.6000 1236.3000 1099.8000 1256.7001 ;
	    RECT 1101.0000 1236.3000 1102.2001 1256.7001 ;
	    RECT 1103.4000 1236.3000 1104.6000 1256.7001 ;
	    RECT 1105.8000 1236.3000 1107.0000 1253.7001 ;
	    RECT 1108.3500 1239.6000 1109.2500 1286.4000 ;
	    RECT 1108.2001 1238.4000 1109.4000 1239.6000 ;
	    RECT 1108.3500 1224.4501 1109.2500 1238.4000 ;
	    RECT 1110.6000 1236.3000 1111.8000 1253.7001 ;
	    RECT 1113.0000 1247.4000 1114.2001 1248.6000 ;
	    RECT 1113.1500 1242.6000 1114.0500 1247.4000 ;
	    RECT 1113.0000 1241.4000 1114.2001 1242.6000 ;
	    RECT 1115.4000 1236.3000 1116.6000 1253.7001 ;
	    RECT 1117.8000 1236.3000 1119.0000 1256.7001 ;
	    RECT 1120.2001 1236.3000 1121.4000 1256.7001 ;
	    RECT 1127.4000 1256.4000 1128.6000 1257.6000 ;
	    RECT 1127.5500 1248.6000 1128.4501 1256.4000 ;
	    RECT 1134.7500 1248.6000 1135.6500 1301.4000 ;
	    RECT 1163.5500 1248.6000 1164.4501 1370.4000 ;
	    RECT 1170.6000 1343.4000 1171.8000 1344.6000 ;
	    RECT 1170.7500 1332.6000 1171.6500 1343.4000 ;
	    RECT 1170.6000 1331.4000 1171.8000 1332.6000 ;
	    RECT 1199.4000 1326.3000 1200.6000 1346.7001 ;
	    RECT 1201.8000 1326.3000 1203.0000 1346.7001 ;
	    RECT 1204.2001 1326.3000 1205.4000 1346.7001 ;
	    RECT 1206.6000 1329.3000 1207.8000 1346.7001 ;
	    RECT 1209.0000 1343.4000 1210.2001 1344.6000 ;
	    RECT 1209.1500 1326.4501 1210.0500 1343.4000 ;
	    RECT 1211.4000 1329.3000 1212.6000 1346.7001 ;
	    RECT 1213.8000 1340.4000 1215.0000 1341.6000 ;
	    RECT 1213.9501 1332.6000 1214.8500 1340.4000 ;
	    RECT 1213.8000 1331.4000 1215.0000 1332.6000 ;
	    RECT 1216.2001 1329.3000 1217.4000 1346.7001 ;
	    RECT 1206.7500 1325.5500 1210.0500 1326.4501 ;
	    RECT 1218.6000 1326.3000 1219.8000 1346.7001 ;
	    RECT 1221.0000 1326.3000 1222.2001 1346.7001 ;
	    RECT 1235.5500 1344.6000 1236.4501 1370.4000 ;
	    RECT 1235.4000 1343.4000 1236.6000 1344.6000 ;
	    RECT 1223.4000 1337.4000 1224.6000 1338.6000 ;
	    RECT 1192.2001 1307.4000 1193.4000 1308.6000 ;
	    RECT 1192.3500 1296.6000 1193.2500 1307.4000 ;
	    RECT 1177.8000 1295.4000 1179.0000 1296.6000 ;
	    RECT 1192.2001 1295.4000 1193.4000 1296.6000 ;
	    RECT 1197.0000 1296.3000 1198.2001 1316.7001 ;
	    RECT 1199.4000 1296.3000 1200.6000 1316.7001 ;
	    RECT 1201.8000 1296.3000 1203.0000 1316.7001 ;
	    RECT 1204.2001 1296.3000 1205.4000 1313.7001 ;
	    RECT 1206.7500 1299.6000 1207.6500 1325.5500 ;
	    RECT 1206.6000 1298.4000 1207.8000 1299.6000 ;
	    RECT 1206.7500 1287.6000 1207.6500 1298.4000 ;
	    RECT 1209.0000 1296.3000 1210.2001 1313.7001 ;
	    RECT 1211.4000 1307.4000 1212.6000 1308.6000 ;
	    RECT 1211.5500 1302.6000 1212.4501 1307.4000 ;
	    RECT 1211.4000 1301.4000 1212.6000 1302.6000 ;
	    RECT 1213.8000 1296.3000 1215.0000 1313.7001 ;
	    RECT 1216.2001 1296.3000 1217.4000 1316.7001 ;
	    RECT 1218.6000 1296.3000 1219.8000 1316.7001 ;
	    RECT 1221.0000 1304.4000 1222.2001 1305.6000 ;
	    RECT 1221.1500 1302.6000 1222.0500 1304.4000 ;
	    RECT 1221.0000 1301.4000 1222.2001 1302.6000 ;
	    RECT 1223.5500 1290.6000 1224.4501 1337.4000 ;
	    RECT 1228.2001 1334.4000 1229.4000 1335.6000 ;
	    RECT 1228.3500 1326.6000 1229.2500 1334.4000 ;
	    RECT 1252.3500 1326.6000 1253.2500 1460.4000 ;
	    RECT 1312.3500 1458.6000 1313.2500 1463.4000 ;
	    RECT 1314.6000 1460.4000 1315.8000 1461.6000 ;
	    RECT 1285.8000 1457.4000 1287.0000 1458.6000 ;
	    RECT 1312.2001 1457.4000 1313.4000 1458.6000 ;
	    RECT 1269.0000 1430.4000 1270.2001 1431.6000 ;
	    RECT 1264.2001 1391.4000 1265.4000 1392.6000 ;
	    RECT 1264.3500 1380.6000 1265.2500 1391.4000 ;
	    RECT 1264.2001 1379.4000 1265.4000 1380.6000 ;
	    RECT 1228.2001 1325.4000 1229.4000 1326.6000 ;
	    RECT 1252.2001 1325.4000 1253.4000 1326.6000 ;
	    RECT 1225.8000 1316.4000 1227.0000 1317.6000 ;
	    RECT 1225.9501 1314.6000 1226.8500 1316.4000 ;
	    RECT 1225.8000 1313.4000 1227.0000 1314.6000 ;
	    RECT 1233.0000 1313.4000 1234.2001 1314.6000 ;
	    RECT 1225.9501 1308.6000 1226.8500 1313.4000 ;
	    RECT 1225.8000 1307.4000 1227.0000 1308.6000 ;
	    RECT 1233.1500 1302.6000 1234.0500 1313.4000 ;
	    RECT 1269.1500 1308.6000 1270.0500 1430.4000 ;
	    RECT 1285.9501 1422.6000 1286.8500 1457.4000 ;
	    RECT 1314.7500 1440.4501 1315.6500 1460.4000 ;
	    RECT 1331.4000 1457.4000 1332.6000 1458.6000 ;
	    RECT 1317.0000 1440.4501 1318.2001 1440.6000 ;
	    RECT 1314.7500 1439.5500 1318.2001 1440.4501 ;
	    RECT 1317.0000 1439.4000 1318.2001 1439.5500 ;
	    RECT 1285.8000 1421.4000 1287.0000 1422.6000 ;
	    RECT 1285.9501 1410.4501 1286.8500 1421.4000 ;
	    RECT 1288.2001 1416.3000 1289.4000 1436.7001 ;
	    RECT 1290.6000 1416.3000 1291.8000 1436.7001 ;
	    RECT 1293.0000 1416.3000 1294.2001 1436.7001 ;
	    RECT 1295.4000 1416.3000 1296.6000 1433.7001 ;
	    RECT 1297.8000 1421.4000 1299.0000 1422.6000 ;
	    RECT 1297.9501 1419.6000 1298.8500 1421.4000 ;
	    RECT 1297.8000 1418.4000 1299.0000 1419.6000 ;
	    RECT 1300.2001 1416.3000 1301.4000 1433.7001 ;
	    RECT 1302.6000 1427.4000 1303.8000 1428.6000 ;
	    RECT 1302.7500 1422.6000 1303.6500 1427.4000 ;
	    RECT 1302.6000 1421.4000 1303.8000 1422.6000 ;
	    RECT 1305.0000 1416.3000 1306.2001 1433.7001 ;
	    RECT 1307.4000 1416.3000 1308.6000 1436.7001 ;
	    RECT 1309.8000 1416.3000 1311.0000 1436.7001 ;
	    RECT 1317.0000 1436.4000 1318.2001 1437.6000 ;
	    RECT 1317.1500 1428.6000 1318.0500 1436.4000 ;
	    RECT 1317.0000 1427.4000 1318.2001 1428.6000 ;
	    RECT 1312.2001 1424.4000 1313.4000 1425.6000 ;
	    RECT 1285.9501 1409.5500 1289.2500 1410.4501 ;
	    RECT 1278.6000 1386.3000 1279.8000 1406.7001 ;
	    RECT 1281.0000 1386.3000 1282.2001 1406.7001 ;
	    RECT 1283.4000 1386.3000 1284.6000 1406.7001 ;
	    RECT 1285.8000 1389.3000 1287.0000 1406.7001 ;
	    RECT 1288.3500 1404.6000 1289.2500 1409.5500 ;
	    RECT 1288.2001 1403.4000 1289.4000 1404.6000 ;
	    RECT 1290.6000 1389.3000 1291.8000 1406.7001 ;
	    RECT 1293.0000 1400.4000 1294.2001 1401.6000 ;
	    RECT 1293.1500 1356.6000 1294.0500 1400.4000 ;
	    RECT 1295.4000 1389.3000 1296.6000 1406.7001 ;
	    RECT 1297.8000 1386.3000 1299.0000 1406.7001 ;
	    RECT 1300.2001 1386.3000 1301.4000 1406.7001 ;
	    RECT 1302.6000 1397.4000 1303.8000 1398.6000 ;
	    RECT 1300.2001 1379.4000 1301.4000 1380.6000 ;
	    RECT 1297.8000 1376.4000 1299.0000 1377.6000 ;
	    RECT 1295.4000 1373.4000 1296.6000 1374.6000 ;
	    RECT 1295.5500 1362.6000 1296.4501 1373.4000 ;
	    RECT 1297.9501 1368.6000 1298.8500 1376.4000 ;
	    RECT 1297.8000 1367.4000 1299.0000 1368.6000 ;
	    RECT 1295.4000 1361.4000 1296.6000 1362.6000 ;
	    RECT 1281.0000 1355.4000 1282.2001 1356.6000 ;
	    RECT 1293.0000 1355.4000 1294.2001 1356.6000 ;
	    RECT 1281.1500 1341.6000 1282.0500 1355.4000 ;
	    RECT 1300.3500 1344.6000 1301.2500 1379.4000 ;
	    RECT 1302.7500 1368.6000 1303.6500 1397.4000 ;
	    RECT 1307.4000 1394.4000 1308.6000 1395.6000 ;
	    RECT 1307.5500 1386.6000 1308.4501 1394.4000 ;
	    RECT 1307.4000 1385.4000 1308.6000 1386.6000 ;
	    RECT 1302.6000 1367.4000 1303.8000 1368.6000 ;
	    RECT 1302.6000 1364.4000 1303.8000 1365.6000 ;
	    RECT 1302.7500 1362.6000 1303.6500 1364.4000 ;
	    RECT 1302.6000 1361.4000 1303.8000 1362.6000 ;
	    RECT 1295.4000 1343.4000 1296.6000 1344.6000 ;
	    RECT 1300.2001 1343.4000 1301.4000 1344.6000 ;
	    RECT 1273.8000 1340.4000 1275.0000 1341.6000 ;
	    RECT 1281.0000 1340.4000 1282.2001 1341.6000 ;
	    RECT 1273.9501 1320.4501 1274.8500 1340.4000 ;
	    RECT 1295.5500 1338.6000 1296.4501 1343.4000 ;
	    RECT 1295.4000 1337.4000 1296.6000 1338.6000 ;
	    RECT 1283.4000 1334.4000 1284.6000 1335.6000 ;
	    RECT 1276.2001 1320.4501 1277.4000 1320.6000 ;
	    RECT 1273.9501 1319.5500 1277.4000 1320.4501 ;
	    RECT 1276.2001 1319.4000 1277.4000 1319.5500 ;
	    RECT 1269.0000 1307.4000 1270.2001 1308.6000 ;
	    RECT 1276.3500 1302.6000 1277.2500 1319.4000 ;
	    RECT 1278.6000 1307.4000 1279.8000 1308.6000 ;
	    RECT 1278.7500 1305.6000 1279.6500 1307.4000 ;
	    RECT 1278.6000 1304.4000 1279.8000 1305.6000 ;
	    RECT 1281.0000 1304.4000 1282.2001 1305.6000 ;
	    RECT 1233.0000 1301.4000 1234.2001 1302.6000 ;
	    RECT 1276.2001 1301.4000 1277.4000 1302.6000 ;
	    RECT 1216.2001 1289.4000 1217.4000 1290.6000 ;
	    RECT 1223.4000 1289.4000 1224.6000 1290.6000 ;
	    RECT 1206.6000 1286.4000 1207.8000 1287.6000 ;
	    RECT 1206.7500 1284.6000 1207.6500 1286.4000 ;
	    RECT 1206.6000 1283.4000 1207.8000 1284.6000 ;
	    RECT 1177.8000 1277.4000 1179.0000 1278.6000 ;
	    RECT 1168.2001 1271.4000 1169.4000 1272.6000 ;
	    RECT 1168.2001 1253.4000 1169.4000 1254.6000 ;
	    RECT 1165.8000 1250.4000 1167.0000 1251.6000 ;
	    RECT 1122.6000 1247.4000 1123.8000 1248.6000 ;
	    RECT 1127.4000 1247.4000 1128.6000 1248.6000 ;
	    RECT 1134.6000 1247.4000 1135.8000 1248.6000 ;
	    RECT 1144.2001 1247.4000 1145.4000 1248.6000 ;
	    RECT 1158.6000 1247.4000 1159.8000 1248.6000 ;
	    RECT 1163.4000 1247.4000 1164.6000 1248.6000 ;
	    RECT 1122.7500 1245.6000 1123.6500 1247.4000 ;
	    RECT 1122.6000 1244.4000 1123.8000 1245.6000 ;
	    RECT 1134.6000 1244.4000 1135.8000 1245.6000 ;
	    RECT 1122.7500 1233.4501 1123.6500 1244.4000 ;
	    RECT 1105.9501 1223.5500 1109.2500 1224.4501 ;
	    RECT 1120.3500 1232.5500 1123.6500 1233.4501 ;
	    RECT 1101.0000 1176.3000 1102.2001 1193.7001 ;
	    RECT 1105.9501 1182.6000 1106.8500 1223.5500 ;
	    RECT 1110.6000 1220.4000 1111.8000 1221.6000 ;
	    RECT 1110.7500 1200.6000 1111.6500 1220.4000 ;
	    RECT 1110.6000 1199.4000 1111.8000 1200.6000 ;
	    RECT 1117.8000 1184.4000 1119.0000 1185.6000 ;
	    RECT 1105.8000 1181.4000 1107.0000 1182.6000 ;
	    RECT 1110.6000 1181.4000 1111.8000 1182.6000 ;
	    RECT 1110.7500 1161.6000 1111.6500 1181.4000 ;
	    RECT 1110.6000 1160.4000 1111.8000 1161.6000 ;
	    RECT 1117.9501 1161.4501 1118.8500 1184.4000 ;
	    RECT 1120.3500 1164.6000 1121.2500 1232.5500 ;
	    RECT 1134.7500 1215.6000 1135.6500 1244.4000 ;
	    RECT 1134.6000 1214.4000 1135.8000 1215.6000 ;
	    RECT 1134.6000 1175.4000 1135.8000 1176.6000 ;
	    RECT 1122.6000 1169.4000 1123.8000 1170.6000 ;
	    RECT 1120.2001 1163.4000 1121.4000 1164.6000 ;
	    RECT 1122.7500 1161.6000 1123.6500 1169.4000 ;
	    RECT 1117.9501 1160.5500 1121.2500 1161.4501 ;
	    RECT 1101.0000 1157.4000 1102.2001 1158.6000 ;
	    RECT 1098.6000 1151.4000 1099.8000 1152.6000 ;
	    RECT 1096.2001 1079.4000 1097.4000 1080.6000 ;
	    RECT 1067.5500 1064.5500 1070.8500 1065.4501 ;
	    RECT 1060.2001 1002.4500 1061.4000 1002.6000 ;
	    RECT 1057.9501 1001.5500 1061.4000 1002.4500 ;
	    RECT 1060.2001 1001.4000 1061.4000 1001.5500 ;
	    RECT 1062.6000 995.4000 1063.8000 996.6000 ;
	    RECT 1062.7500 984.6000 1063.6500 995.4000 ;
	    RECT 1062.6000 983.4000 1063.8000 984.6000 ;
	    RECT 1050.7500 899.5500 1054.0500 900.4500 ;
	    RECT 1026.6000 881.4000 1027.8000 882.6000 ;
	    RECT 1031.4000 881.4000 1032.6000 882.6000 ;
	    RECT 1033.8000 881.4000 1035.0000 882.6000 ;
	    RECT 1036.2001 881.4000 1037.4000 882.6000 ;
	    RECT 1038.6000 881.4000 1039.8000 882.6000 ;
	    RECT 1026.7500 876.6000 1027.6500 881.4000 ;
	    RECT 1026.6000 875.4000 1027.8000 876.6000 ;
	    RECT 1031.5500 846.6000 1032.4501 881.4000 ;
	    RECT 1038.7500 876.6000 1039.6500 881.4000 ;
	    RECT 1038.6000 875.4000 1039.8000 876.6000 ;
	    RECT 1031.4000 845.4000 1032.6000 846.6000 ;
	    RECT 1024.2001 833.4000 1025.4000 834.6000 ;
	    RECT 1050.7500 828.6000 1051.6500 899.5500 ;
	    RECT 1053.0000 878.4000 1054.2001 879.6000 ;
	    RECT 1053.1500 864.6000 1054.0500 878.4000 ;
	    RECT 1053.0000 863.4000 1054.2001 864.6000 ;
	    RECT 1050.6000 827.4000 1051.8000 828.6000 ;
	    RECT 1050.6000 809.4000 1051.8000 810.6000 ;
	    RECT 1060.2001 809.4000 1061.4000 810.6000 ;
	    RECT 1036.2001 786.3000 1037.4000 806.7000 ;
	    RECT 1038.6000 786.3000 1039.8000 806.7000 ;
	    RECT 1041.0000 786.3000 1042.2001 806.7000 ;
	    RECT 1043.4000 789.3000 1044.6000 806.7000 ;
	    RECT 1045.8000 803.4000 1047.0000 804.6000 ;
	    RECT 1045.9501 780.6000 1046.8500 803.4000 ;
	    RECT 1048.2001 789.3000 1049.4000 806.7000 ;
	    RECT 1050.7500 801.6000 1051.6500 809.4000 ;
	    RECT 1050.6000 800.4000 1051.8000 801.6000 ;
	    RECT 1053.0000 789.3000 1054.2001 806.7000 ;
	    RECT 1055.4000 786.3000 1056.6000 806.7000 ;
	    RECT 1057.8000 786.3000 1059.0000 806.7000 ;
	    RECT 1060.3500 798.6000 1061.2500 809.4000 ;
	    RECT 1060.2001 797.4000 1061.4000 798.6000 ;
	    RECT 1038.6000 779.4000 1039.8000 780.6000 ;
	    RECT 1045.8000 779.4000 1047.0000 780.6000 ;
	    RECT 1026.6000 743.4000 1027.8000 744.6000 ;
	    RECT 1026.7500 720.6000 1027.6500 743.4000 ;
	    RECT 1029.0000 726.3000 1030.2001 746.7000 ;
	    RECT 1031.4000 726.3000 1032.6000 746.7000 ;
	    RECT 1033.8000 726.3000 1035.0000 746.7000 ;
	    RECT 1036.2001 729.3000 1037.4000 746.7000 ;
	    RECT 1038.7500 744.6000 1039.6500 779.4000 ;
	    RECT 1060.3500 774.6000 1061.2500 797.4000 ;
	    RECT 1065.0000 794.4000 1066.2001 795.6000 ;
	    RECT 1065.1500 786.6000 1066.0500 794.4000 ;
	    RECT 1065.0000 785.4000 1066.2001 786.6000 ;
	    RECT 1060.2001 773.4000 1061.4000 774.6000 ;
	    RECT 1065.0000 773.4000 1066.2001 774.6000 ;
	    RECT 1065.1500 768.6000 1066.0500 773.4000 ;
	    RECT 1065.0000 767.4000 1066.2001 768.6000 ;
	    RECT 1055.4000 764.4000 1056.6000 765.6000 ;
	    RECT 1043.4000 761.4000 1044.6000 762.6000 ;
	    RECT 1038.6000 743.4000 1039.8000 744.6000 ;
	    RECT 1038.7500 732.6000 1039.6500 743.4000 ;
	    RECT 1038.6000 731.4000 1039.8000 732.6000 ;
	    RECT 1041.0000 729.3000 1042.2001 746.7000 ;
	    RECT 1043.5500 741.6000 1044.4501 761.4000 ;
	    RECT 1043.4000 740.4000 1044.6000 741.6000 ;
	    RECT 1045.8000 729.3000 1047.0000 746.7000 ;
	    RECT 1048.2001 726.3000 1049.4000 746.7000 ;
	    RECT 1050.6000 726.3000 1051.8000 746.7000 ;
	    RECT 1053.0000 737.4000 1054.2001 738.6000 ;
	    RECT 1026.6000 719.4000 1027.8000 720.6000 ;
	    RECT 1026.7500 702.6000 1027.6500 719.4000 ;
	    RECT 1026.6000 701.4000 1027.8000 702.6000 ;
	    RECT 1036.2001 665.4000 1037.4000 666.6000 ;
	    RECT 1019.4000 653.4000 1020.6000 654.6000 ;
	    RECT 1019.5500 651.6000 1020.4500 653.4000 ;
	    RECT 1019.4000 650.4000 1020.6000 651.6000 ;
	    RECT 1036.3500 639.6000 1037.2500 665.4000 ;
	    RECT 1036.2001 638.4000 1037.4000 639.6000 ;
	    RECT 1036.3500 612.6000 1037.2500 638.4000 ;
	    RECT 1055.5500 630.6000 1056.4501 764.4000 ;
	    RECT 1060.2001 737.4000 1061.4000 738.6000 ;
	    RECT 1057.8000 734.4000 1059.0000 735.6000 ;
	    RECT 1057.9501 723.6000 1058.8500 734.4000 ;
	    RECT 1057.8000 722.4000 1059.0000 723.6000 ;
	    RECT 1057.9501 720.6000 1058.8500 722.4000 ;
	    RECT 1057.8000 719.4000 1059.0000 720.6000 ;
	    RECT 1057.9501 642.6000 1058.8500 719.4000 ;
	    RECT 1057.8000 641.4000 1059.0000 642.6000 ;
	    RECT 1055.4000 629.4000 1056.6000 630.6000 ;
	    RECT 1060.3500 618.6000 1061.2500 737.4000 ;
	    RECT 1065.0000 629.4000 1066.2001 630.6000 ;
	    RECT 1060.2001 617.4000 1061.4000 618.6000 ;
	    RECT 1036.2001 611.4000 1037.4000 612.6000 ;
	    RECT 1036.2001 581.4000 1037.4000 582.6000 ;
	    RECT 1017.0000 575.4000 1018.2000 576.6000 ;
	    RECT 1017.1500 561.6000 1018.0500 575.4000 ;
	    RECT 1017.0000 560.4000 1018.2000 561.6000 ;
	    RECT 1021.8000 527.4000 1023.0000 528.6000 ;
	    RECT 1021.9500 525.6000 1022.8500 527.4000 ;
	    RECT 1021.8000 524.4000 1023.0000 525.6000 ;
	    RECT 1021.9500 486.6000 1022.8500 524.4000 ;
	    RECT 1033.8000 515.4000 1035.0000 516.6000 ;
	    RECT 1031.4000 494.4000 1032.6000 495.6000 ;
	    RECT 1031.5500 486.6000 1032.4501 494.4000 ;
	    RECT 1021.8000 485.4000 1023.0000 486.6000 ;
	    RECT 1031.4000 485.4000 1032.6000 486.6000 ;
	    RECT 1019.4000 473.4000 1020.6000 474.6000 ;
	    RECT 1019.5500 462.6000 1020.4500 473.4000 ;
	    RECT 1021.9500 468.6000 1022.8500 485.4000 ;
	    RECT 1026.6000 479.4000 1027.8000 480.6000 ;
	    RECT 1031.4000 479.4000 1032.6000 480.6000 ;
	    RECT 1026.7500 474.6000 1027.6500 479.4000 ;
	    RECT 1031.5500 474.6000 1032.4501 479.4000 ;
	    RECT 1026.6000 473.4000 1027.8000 474.6000 ;
	    RECT 1031.4000 474.4500 1032.6000 474.6000 ;
	    RECT 1033.9501 474.4500 1034.8500 515.4000 ;
	    RECT 1036.3500 498.6000 1037.2500 581.4000 ;
	    RECT 1043.4000 575.4000 1044.6000 576.6000 ;
	    RECT 1043.5500 561.6000 1044.4501 575.4000 ;
	    RECT 1043.4000 560.4000 1044.6000 561.6000 ;
	    RECT 1050.6000 560.4000 1051.8000 561.6000 ;
	    RECT 1050.7500 540.6000 1051.6500 560.4000 ;
	    RECT 1043.4000 539.4000 1044.6000 540.6000 ;
	    RECT 1050.6000 539.4000 1051.8000 540.6000 ;
	    RECT 1060.2001 539.4000 1061.4000 540.6000 ;
	    RECT 1045.8000 527.4000 1047.0000 528.6000 ;
	    RECT 1045.9501 525.6000 1046.8500 527.4000 ;
	    RECT 1045.8000 524.4000 1047.0000 525.6000 ;
	    RECT 1060.3500 522.6000 1061.2500 539.4000 ;
	    RECT 1043.4000 521.4000 1044.6000 522.6000 ;
	    RECT 1060.2001 521.4000 1061.4000 522.6000 ;
	    RECT 1062.6000 521.4000 1063.8000 522.6000 ;
	    RECT 1036.2001 497.4000 1037.4000 498.6000 ;
	    RECT 1036.3500 480.6000 1037.2500 497.4000 ;
	    RECT 1038.6000 486.3000 1039.8000 506.7000 ;
	    RECT 1041.0000 486.3000 1042.2001 506.7000 ;
	    RECT 1043.4000 489.3000 1044.6000 506.7000 ;
	    RECT 1045.8000 503.4000 1047.0000 504.6000 ;
	    RECT 1045.9501 501.6000 1046.8500 503.4000 ;
	    RECT 1045.8000 500.4000 1047.0000 501.6000 ;
	    RECT 1048.2001 489.3000 1049.4000 506.7000 ;
	    RECT 1050.6000 503.4000 1051.8000 504.6000 ;
	    RECT 1050.7500 492.6000 1051.6500 503.4000 ;
	    RECT 1050.6000 491.4000 1051.8000 492.6000 ;
	    RECT 1053.0000 489.3000 1054.2001 506.7000 ;
	    RECT 1048.2001 485.4000 1049.4000 486.6000 ;
	    RECT 1055.4000 486.3000 1056.6000 506.7000 ;
	    RECT 1057.8000 486.3000 1059.0000 506.7000 ;
	    RECT 1060.2001 486.3000 1061.4000 506.7000 ;
	    RECT 1065.1500 504.6000 1066.0500 629.4000 ;
	    RECT 1067.5500 606.6000 1068.4501 1064.5500 ;
	    RECT 1072.2001 1064.4000 1073.4000 1065.6000 ;
	    RECT 1072.3500 1062.4501 1073.2500 1064.4000 ;
	    RECT 1069.9501 1061.5500 1073.2500 1062.4501 ;
	    RECT 1069.9501 942.6000 1070.8500 1061.5500 ;
	    RECT 1074.6000 1056.3000 1075.8000 1076.7001 ;
	    RECT 1077.0000 1056.3000 1078.2001 1076.7001 ;
	    RECT 1079.4000 1056.3000 1080.6000 1073.7001 ;
	    RECT 1081.8000 1061.4000 1083.0000 1062.6000 ;
	    RECT 1081.9501 1050.6000 1082.8500 1061.4000 ;
	    RECT 1084.2001 1056.3000 1085.4000 1073.7001 ;
	    RECT 1086.6000 1058.4000 1087.8000 1059.6000 ;
	    RECT 1081.8000 1049.4000 1083.0000 1050.6000 ;
	    RECT 1079.4000 1019.4000 1080.6000 1020.6000 ;
	    RECT 1072.2001 980.4000 1073.4000 981.6000 ;
	    RECT 1072.3500 960.6000 1073.2500 980.4000 ;
	    RECT 1079.5500 975.6000 1080.4501 1019.4000 ;
	    RECT 1084.2001 980.4000 1085.4000 981.6000 ;
	    RECT 1079.4000 974.4000 1080.6000 975.6000 ;
	    RECT 1072.2001 959.4000 1073.4000 960.6000 ;
	    RECT 1069.8000 941.4000 1071.0000 942.6000 ;
	    RECT 1084.3500 924.6000 1085.2500 980.4000 ;
	    RECT 1086.7500 966.6000 1087.6500 1058.4000 ;
	    RECT 1089.0000 1056.3000 1090.2001 1073.7001 ;
	    RECT 1091.4000 1056.3000 1092.6000 1076.7001 ;
	    RECT 1093.8000 1056.3000 1095.0000 1076.7001 ;
	    RECT 1096.2001 1056.3000 1097.4000 1076.7001 ;
	    RECT 1093.8000 1004.4000 1095.0000 1005.6000 ;
	    RECT 1091.4000 995.4000 1092.6000 996.6000 ;
	    RECT 1089.0000 983.4000 1090.2001 984.6000 ;
	    RECT 1086.6000 965.4000 1087.8000 966.6000 ;
	    RECT 1089.1500 951.6000 1090.0500 983.4000 ;
	    RECT 1089.0000 950.4000 1090.2001 951.6000 ;
	    RECT 1084.2001 923.4000 1085.4000 924.6000 ;
	    RECT 1089.1500 801.6000 1090.0500 950.4000 ;
	    RECT 1089.0000 800.4000 1090.2001 801.6000 ;
	    RECT 1072.2001 797.4000 1073.4000 798.6000 ;
	    RECT 1069.8000 737.4000 1071.0000 738.6000 ;
	    RECT 1069.9501 648.6000 1070.8500 737.4000 ;
	    RECT 1072.3500 708.6000 1073.2500 797.4000 ;
	    RECT 1086.6000 785.4000 1087.8000 786.6000 ;
	    RECT 1077.0000 755.4000 1078.2001 756.6000 ;
	    RECT 1084.2001 756.3000 1085.4000 773.7000 ;
	    RECT 1077.1500 750.6000 1078.0500 755.4000 ;
	    RECT 1077.0000 749.4000 1078.2001 750.6000 ;
	    RECT 1086.7500 741.6000 1087.6500 785.4000 ;
	    RECT 1086.6000 740.4000 1087.8000 741.6000 ;
	    RECT 1081.8000 734.4000 1083.0000 735.6000 ;
	    RECT 1081.9501 714.6000 1082.8500 734.4000 ;
	    RECT 1081.8000 713.4000 1083.0000 714.6000 ;
	    RECT 1081.9501 711.6000 1082.8500 713.4000 ;
	    RECT 1081.8000 710.4000 1083.0000 711.6000 ;
	    RECT 1072.2001 707.4000 1073.4000 708.6000 ;
	    RECT 1069.8000 647.4000 1071.0000 648.6000 ;
	    RECT 1081.8000 641.4000 1083.0000 642.6000 ;
	    RECT 1074.6000 638.4000 1075.8000 639.6000 ;
	    RECT 1067.4000 605.4000 1068.6000 606.6000 ;
	    RECT 1069.8000 509.4000 1071.0000 510.6000 ;
	    RECT 1065.0000 503.4000 1066.2001 504.6000 ;
	    RECT 1036.2001 479.4000 1037.4000 480.6000 ;
	    RECT 1041.0000 479.4000 1042.2001 480.6000 ;
	    RECT 1045.8000 479.4000 1047.0000 480.6000 ;
	    RECT 1031.4000 473.5500 1034.8500 474.4500 ;
	    RECT 1031.4000 473.4000 1032.6000 473.5500 ;
	    RECT 1036.2001 473.4000 1037.4000 474.6000 ;
	    RECT 1021.8000 467.4000 1023.0000 468.6000 ;
	    RECT 1026.6000 467.4000 1027.8000 468.6000 ;
	    RECT 1026.7500 465.6000 1027.6500 467.4000 ;
	    RECT 1036.3500 465.6000 1037.2500 473.4000 ;
	    RECT 1026.6000 464.4000 1027.8000 465.6000 ;
	    RECT 1031.4000 464.4000 1032.6000 465.6000 ;
	    RECT 1036.2001 464.4000 1037.4000 465.6000 ;
	    RECT 1019.4000 461.4000 1020.6000 462.6000 ;
	    RECT 1029.0000 461.4000 1030.2001 462.6000 ;
	    RECT 1031.5500 444.6000 1032.4501 464.4000 ;
	    RECT 1033.8000 461.4000 1035.0000 462.6000 ;
	    RECT 1033.9501 444.6000 1034.8500 461.4000 ;
	    RECT 1031.4000 443.4000 1032.6000 444.6000 ;
	    RECT 1033.8000 443.4000 1035.0000 444.6000 ;
	    RECT 1021.8000 437.4000 1023.0000 438.6000 ;
	    RECT 1009.8000 401.4000 1011.0000 402.6000 ;
	    RECT 1014.6000 398.4000 1015.8000 399.6000 ;
	    RECT 1014.7500 390.6000 1015.6500 398.4000 ;
	    RECT 1012.2000 389.4000 1013.4000 390.6000 ;
	    RECT 1014.6000 389.4000 1015.8000 390.6000 ;
	    RECT 1012.3500 375.6000 1013.2500 389.4000 ;
	    RECT 1012.2000 374.4000 1013.4000 375.6000 ;
	    RECT 1019.4000 359.4000 1020.6000 360.6000 ;
	    RECT 1019.4000 356.4000 1020.6000 357.6000 ;
	    RECT 1019.5500 348.6000 1020.4500 356.4000 ;
	    RECT 1019.4000 347.4000 1020.6000 348.6000 ;
	    RECT 1021.9500 345.4500 1022.8500 437.4000 ;
	    RECT 1033.9501 396.6000 1034.8500 443.4000 ;
	    RECT 1041.1500 438.6000 1042.0500 479.4000 ;
	    RECT 1045.9501 462.6000 1046.8500 479.4000 ;
	    RECT 1048.3500 465.6000 1049.2500 485.4000 ;
	    RECT 1048.2001 464.4000 1049.4000 465.6000 ;
	    RECT 1045.8000 461.4000 1047.0000 462.6000 ;
	    RECT 1053.0000 443.4000 1054.2001 444.6000 ;
	    RECT 1041.0000 437.4000 1042.2001 438.6000 ;
	    RECT 1050.6000 434.4000 1051.8000 435.6000 ;
	    RECT 1050.7500 426.6000 1051.6500 434.4000 ;
	    RECT 1050.6000 425.4000 1051.8000 426.6000 ;
	    RECT 1050.6000 423.4500 1051.8000 423.6000 ;
	    RECT 1048.3500 422.5500 1051.8000 423.4500 ;
	    RECT 1041.0000 407.4000 1042.2001 408.6000 ;
	    RECT 1048.3500 402.6000 1049.2500 422.5500 ;
	    RECT 1050.6000 422.4000 1051.8000 422.5500 ;
	    RECT 1053.1500 414.6000 1054.0500 443.4000 ;
	    RECT 1055.4000 437.4000 1056.6000 438.6000 ;
	    RECT 1057.8000 426.3000 1059.0000 446.7000 ;
	    RECT 1060.2001 426.3000 1061.4000 446.7000 ;
	    RECT 1062.6000 429.3000 1063.8000 446.7000 ;
	    RECT 1065.0000 440.4000 1066.2001 441.6000 ;
	    RECT 1065.1500 420.6000 1066.0500 440.4000 ;
	    RECT 1067.4000 429.3000 1068.6000 446.7000 ;
	    RECT 1069.9501 444.6000 1070.8500 509.4000 ;
	    RECT 1074.7500 492.6000 1075.6500 638.4000 ;
	    RECT 1081.9501 624.6000 1082.8500 641.4000 ;
	    RECT 1081.8000 623.4000 1083.0000 624.6000 ;
	    RECT 1091.5500 564.6000 1092.4501 995.4000 ;
	    RECT 1093.9501 975.6000 1094.8500 1004.4000 ;
	    RECT 1096.2001 989.4000 1097.4000 990.6000 ;
	    RECT 1093.8000 974.4000 1095.0000 975.6000 ;
	    RECT 1093.8000 794.4000 1095.0000 795.6000 ;
	    RECT 1093.9501 786.6000 1094.8500 794.4000 ;
	    RECT 1093.8000 785.4000 1095.0000 786.6000 ;
	    RECT 1093.9501 780.6000 1094.8500 785.4000 ;
	    RECT 1093.8000 779.4000 1095.0000 780.6000 ;
	    RECT 1093.8000 767.4000 1095.0000 768.6000 ;
	    RECT 1093.9501 765.6000 1094.8500 767.4000 ;
	    RECT 1093.8000 764.4000 1095.0000 765.6000 ;
	    RECT 1096.3500 756.6000 1097.2500 989.4000 ;
	    RECT 1098.7500 804.6000 1099.6500 1151.4000 ;
	    RECT 1098.6000 803.4000 1099.8000 804.6000 ;
	    RECT 1098.6000 800.4000 1099.8000 801.6000 ;
	    RECT 1098.7500 780.6000 1099.6500 800.4000 ;
	    RECT 1098.6000 779.4000 1099.8000 780.6000 ;
	    RECT 1096.2001 755.4000 1097.4000 756.6000 ;
	    RECT 1098.6000 756.3000 1099.8000 773.7000 ;
	    RECT 1101.1500 768.6000 1102.0500 1157.4000 ;
	    RECT 1110.7500 1140.6000 1111.6500 1160.4000 ;
	    RECT 1120.3500 1155.6000 1121.2500 1160.5500 ;
	    RECT 1122.6000 1160.4000 1123.8000 1161.6000 ;
	    RECT 1120.2001 1154.4000 1121.4000 1155.6000 ;
	    RECT 1110.6000 1139.4000 1111.8000 1140.6000 ;
	    RECT 1113.0000 1109.4000 1114.2001 1110.6000 ;
	    RECT 1110.6000 1085.4000 1111.8000 1086.6000 ;
	    RECT 1110.7500 1071.6000 1111.6500 1085.4000 ;
	    RECT 1110.6000 1070.4000 1111.8000 1071.6000 ;
	    RECT 1113.1500 1062.6000 1114.0500 1109.4000 ;
	    RECT 1129.8000 1100.4000 1131.0000 1101.6000 ;
	    RECT 1129.9501 1098.6000 1130.8500 1100.4000 ;
	    RECT 1134.7500 1098.6000 1135.6500 1175.4000 ;
	    RECT 1144.3500 1164.6000 1145.2500 1247.4000 ;
	    RECT 1165.9501 1224.6000 1166.8500 1250.4000 ;
	    RECT 1165.8000 1223.4000 1167.0000 1224.6000 ;
	    RECT 1156.2001 1193.4000 1157.4000 1194.6000 ;
	    RECT 1156.3500 1170.6000 1157.2500 1193.4000 ;
	    RECT 1165.9501 1188.6000 1166.8500 1223.4000 ;
	    RECT 1165.8000 1187.4000 1167.0000 1188.6000 ;
	    RECT 1156.2001 1169.4000 1157.4000 1170.6000 ;
	    RECT 1156.3500 1164.6000 1157.2500 1169.4000 ;
	    RECT 1144.2001 1163.4000 1145.4000 1164.6000 ;
	    RECT 1156.2001 1163.4000 1157.4000 1164.6000 ;
	    RECT 1115.4000 1098.4501 1116.6000 1098.6000 ;
	    RECT 1120.2001 1098.4501 1121.4000 1098.6000 ;
	    RECT 1115.4000 1097.5500 1121.4000 1098.4501 ;
	    RECT 1115.4000 1097.4000 1116.6000 1097.5500 ;
	    RECT 1120.2001 1097.4000 1121.4000 1097.5500 ;
	    RECT 1129.8000 1097.4000 1131.0000 1098.6000 ;
	    RECT 1134.6000 1097.4000 1135.8000 1098.6000 ;
	    RECT 1146.6000 1097.4000 1147.8000 1098.6000 ;
	    RECT 1120.2001 1079.4000 1121.4000 1080.6000 ;
	    RECT 1113.0000 1061.4000 1114.2001 1062.6000 ;
	    RECT 1110.6000 1037.4000 1111.8000 1038.6000 ;
	    RECT 1110.7500 990.6000 1111.6500 1037.4000 ;
	    RECT 1110.6000 989.4000 1111.8000 990.6000 ;
	    RECT 1103.4000 980.4000 1104.6000 981.6000 ;
	    RECT 1103.5500 942.6000 1104.4501 980.4000 ;
	    RECT 1115.4000 965.4000 1116.6000 966.6000 ;
	    RECT 1103.4000 941.4000 1104.6000 942.6000 ;
	    RECT 1105.8000 936.3000 1107.0000 956.7000 ;
	    RECT 1108.2001 936.3000 1109.4000 956.7000 ;
	    RECT 1110.6000 936.3000 1111.8000 956.7000 ;
	    RECT 1113.0000 936.3000 1114.2001 953.7000 ;
	    RECT 1115.5500 939.6000 1116.4501 965.4000 ;
	    RECT 1115.4000 938.4000 1116.6000 939.6000 ;
	    RECT 1115.5500 936.6000 1116.4501 938.4000 ;
	    RECT 1115.4000 935.4000 1116.6000 936.6000 ;
	    RECT 1117.8000 936.3000 1119.0000 953.7000 ;
	    RECT 1120.3500 948.6000 1121.2500 1079.4000 ;
	    RECT 1146.7500 1044.6000 1147.6500 1097.4000 ;
	    RECT 1153.8000 1079.4000 1155.0000 1080.6000 ;
	    RECT 1153.9501 1062.6000 1154.8500 1079.4000 ;
	    RECT 1158.6000 1067.4000 1159.8000 1068.6000 ;
	    RECT 1153.8000 1061.4000 1155.0000 1062.6000 ;
	    RECT 1146.6000 1043.4000 1147.8000 1044.6000 ;
	    RECT 1137.0000 995.4000 1138.2001 996.6000 ;
	    RECT 1129.8000 989.4000 1131.0000 990.6000 ;
	    RECT 1129.9501 981.6000 1130.8500 989.4000 ;
	    RECT 1134.6000 983.4000 1135.8000 984.6000 ;
	    RECT 1137.1500 981.6000 1138.0500 995.4000 ;
	    RECT 1158.7500 990.6000 1159.6500 1067.4000 ;
	    RECT 1163.4000 1010.4000 1164.6000 1011.6000 ;
	    RECT 1163.5500 1002.6000 1164.4501 1010.4000 ;
	    RECT 1163.4000 1001.4000 1164.6000 1002.6000 ;
	    RECT 1158.6000 989.4000 1159.8000 990.6000 ;
	    RECT 1163.5500 984.6000 1164.4501 1001.4000 ;
	    RECT 1149.0000 983.4000 1150.2001 984.6000 ;
	    RECT 1163.4000 983.4000 1164.6000 984.6000 ;
	    RECT 1129.8000 980.4000 1131.0000 981.6000 ;
	    RECT 1132.2001 980.4000 1133.4000 981.6000 ;
	    RECT 1137.0000 980.4000 1138.2001 981.6000 ;
	    RECT 1122.6000 977.4000 1123.8000 978.6000 ;
	    RECT 1129.9501 966.6000 1130.8500 980.4000 ;
	    RECT 1132.3500 978.6000 1133.2500 980.4000 ;
	    RECT 1132.2001 977.4000 1133.4000 978.6000 ;
	    RECT 1129.8000 965.4000 1131.0000 966.6000 ;
	    RECT 1134.6000 965.4000 1135.8000 966.6000 ;
	    RECT 1134.7500 960.6000 1135.6500 965.4000 ;
	    RECT 1134.6000 959.4000 1135.8000 960.6000 ;
	    RECT 1120.2001 947.4000 1121.4000 948.6000 ;
	    RECT 1120.2001 941.4000 1121.4000 942.6000 ;
	    RECT 1122.6000 936.3000 1123.8000 953.7000 ;
	    RECT 1125.0000 936.3000 1126.2001 956.7000 ;
	    RECT 1127.4000 936.3000 1128.6000 956.7000 ;
	    RECT 1134.7500 948.6000 1135.6500 959.4000 ;
	    RECT 1149.1500 948.6000 1150.0500 983.4000 ;
	    RECT 1129.8000 947.4000 1131.0000 948.6000 ;
	    RECT 1134.6000 947.4000 1135.8000 948.6000 ;
	    RECT 1149.0000 947.4000 1150.2001 948.6000 ;
	    RECT 1165.8000 947.4000 1167.0000 948.6000 ;
	    RECT 1129.9501 945.6000 1130.8500 947.4000 ;
	    RECT 1129.8000 944.4000 1131.0000 945.6000 ;
	    RECT 1141.8000 935.4000 1143.0000 936.6000 ;
	    RECT 1132.2001 906.3000 1133.4000 926.7000 ;
	    RECT 1134.6000 906.3000 1135.8000 926.7000 ;
	    RECT 1137.0000 906.3000 1138.2001 926.7000 ;
	    RECT 1139.4000 909.3000 1140.6000 926.7000 ;
	    RECT 1141.9501 924.6000 1142.8500 935.4000 ;
	    RECT 1141.8000 923.4000 1143.0000 924.6000 ;
	    RECT 1141.9501 906.6000 1142.8500 923.4000 ;
	    RECT 1144.2001 909.3000 1145.4000 926.7000 ;
	    RECT 1146.6000 923.4000 1147.8000 924.6000 ;
	    RECT 1146.7500 921.6000 1147.6500 923.4000 ;
	    RECT 1146.6000 920.4000 1147.8000 921.6000 ;
	    RECT 1149.0000 909.3000 1150.2001 926.7000 ;
	    RECT 1141.8000 905.4000 1143.0000 906.6000 ;
	    RECT 1151.4000 906.3000 1152.6000 926.7000 ;
	    RECT 1153.8000 906.3000 1155.0000 926.7000 ;
	    RECT 1156.2001 917.4000 1157.4000 918.6000 ;
	    RECT 1156.3500 900.6000 1157.2500 917.4000 ;
	    RECT 1161.0000 914.4000 1162.2001 915.6000 ;
	    RECT 1161.1500 906.6000 1162.0500 914.4000 ;
	    RECT 1168.3500 912.6000 1169.2500 1253.4000 ;
	    RECT 1168.2001 911.4000 1169.4000 912.6000 ;
	    RECT 1161.0000 905.4000 1162.2001 906.6000 ;
	    RECT 1156.2001 899.4000 1157.4000 900.6000 ;
	    RECT 1137.0000 863.4000 1138.2001 864.6000 ;
	    RECT 1120.2001 857.4000 1121.4000 858.6000 ;
	    RECT 1117.8000 818.4000 1119.0000 819.6000 ;
	    RECT 1117.9501 816.6000 1118.8500 818.4000 ;
	    RECT 1117.8000 815.4000 1119.0000 816.6000 ;
	    RECT 1103.4000 797.4000 1104.6000 798.6000 ;
	    RECT 1103.5500 774.6000 1104.4501 797.4000 ;
	    RECT 1117.9501 795.6000 1118.8500 815.4000 ;
	    RECT 1117.8000 794.4000 1119.0000 795.6000 ;
	    RECT 1103.4000 773.4000 1104.6000 774.6000 ;
	    RECT 1101.0000 767.4000 1102.2001 768.6000 ;
	    RECT 1101.0000 761.4000 1102.2001 762.6000 ;
	    RECT 1101.1500 756.6000 1102.0500 761.4000 ;
	    RECT 1103.4000 759.3000 1104.6000 767.7000 ;
	    RECT 1117.8000 767.4000 1119.0000 768.6000 ;
	    RECT 1101.0000 755.4000 1102.2001 756.6000 ;
	    RECT 1117.9501 750.6000 1118.8500 767.4000 ;
	    RECT 1117.8000 749.4000 1119.0000 750.6000 ;
	    RECT 1105.8000 737.4000 1107.0000 738.6000 ;
	    RECT 1105.9501 732.6000 1106.8500 737.4000 ;
	    RECT 1105.8000 731.4000 1107.0000 732.6000 ;
	    RECT 1096.2001 666.3000 1097.4000 686.7000 ;
	    RECT 1098.6000 666.3000 1099.8000 686.7000 ;
	    RECT 1101.0000 666.3000 1102.2001 686.7000 ;
	    RECT 1103.4000 669.3000 1104.6000 686.7000 ;
	    RECT 1105.9501 684.6000 1106.8500 731.4000 ;
	    RECT 1110.6000 701.4000 1111.8000 702.6000 ;
	    RECT 1105.8000 683.4000 1107.0000 684.6000 ;
	    RECT 1105.9501 630.4500 1106.8500 683.4000 ;
	    RECT 1108.2001 669.3000 1109.4000 686.7000 ;
	    RECT 1110.7500 681.6000 1111.6500 701.4000 ;
	    RECT 1110.6000 680.4000 1111.8000 681.6000 ;
	    RECT 1110.6000 671.4000 1111.8000 672.6000 ;
	    RECT 1110.7500 642.6000 1111.6500 671.4000 ;
	    RECT 1113.0000 669.3000 1114.2001 686.7000 ;
	    RECT 1115.4000 666.3000 1116.6000 686.7000 ;
	    RECT 1117.8000 666.3000 1119.0000 686.7000 ;
	    RECT 1120.3500 678.6000 1121.2500 857.4000 ;
	    RECT 1137.1500 852.6000 1138.0500 863.4000 ;
	    RECT 1137.0000 851.4000 1138.2001 852.6000 ;
	    RECT 1153.8000 846.3000 1155.0000 866.7000 ;
	    RECT 1156.2001 846.3000 1157.4000 866.7000 ;
	    RECT 1158.6000 846.3000 1159.8000 866.7000 ;
	    RECT 1161.0000 849.3000 1162.2001 866.7000 ;
	    RECT 1163.4000 863.4000 1164.6000 864.6000 ;
	    RECT 1139.4000 830.4000 1140.6000 831.6000 ;
	    RECT 1139.5500 798.6000 1140.4501 830.4000 ;
	    RECT 1151.4000 827.4000 1152.6000 828.6000 ;
	    RECT 1151.5500 801.6000 1152.4501 827.4000 ;
	    RECT 1153.8000 816.3000 1155.0000 836.7000 ;
	    RECT 1156.2001 816.3000 1157.4000 836.7000 ;
	    RECT 1158.6000 816.3000 1159.8000 836.7000 ;
	    RECT 1161.0000 816.3000 1162.2001 833.7000 ;
	    RECT 1163.5500 819.6000 1164.4501 863.4000 ;
	    RECT 1165.8000 849.3000 1167.0000 866.7000 ;
	    RECT 1168.2001 860.4000 1169.4000 861.6000 ;
	    RECT 1168.3500 852.6000 1169.2500 860.4000 ;
	    RECT 1168.2001 851.4000 1169.4000 852.6000 ;
	    RECT 1170.6000 849.3000 1171.8000 866.7000 ;
	    RECT 1173.0000 846.3000 1174.2001 866.7000 ;
	    RECT 1175.4000 846.3000 1176.6000 866.7000 ;
	    RECT 1177.9501 858.6000 1178.8500 1277.4000 ;
	    RECT 1213.8000 1274.4000 1215.0000 1275.6000 ;
	    RECT 1192.2001 1265.4000 1193.4000 1266.6000 ;
	    RECT 1192.3500 1221.6000 1193.2500 1265.4000 ;
	    RECT 1213.9501 1263.6000 1214.8500 1274.4000 ;
	    RECT 1213.8000 1262.4000 1215.0000 1263.6000 ;
	    RECT 1213.9501 1242.6000 1214.8500 1262.4000 ;
	    RECT 1213.8000 1241.4000 1215.0000 1242.6000 ;
	    RECT 1192.2001 1220.4000 1193.4000 1221.6000 ;
	    RECT 1194.6000 1215.3000 1195.8000 1223.7001 ;
	    RECT 1197.0000 1220.4000 1198.2001 1221.6000 ;
	    RECT 1197.1500 1218.6000 1198.0500 1220.4000 ;
	    RECT 1197.0000 1217.4000 1198.2001 1218.6000 ;
	    RECT 1180.2001 1184.4000 1181.4000 1185.6000 ;
	    RECT 1180.3500 1155.6000 1181.2500 1184.4000 ;
	    RECT 1197.1500 1176.6000 1198.0500 1217.4000 ;
	    RECT 1199.4000 1209.3000 1200.6000 1226.7001 ;
	    RECT 1204.2001 1218.4501 1205.4000 1218.6000 ;
	    RECT 1201.9501 1217.5500 1205.4000 1218.4501 ;
	    RECT 1197.0000 1175.4000 1198.2001 1176.6000 ;
	    RECT 1182.6000 1160.4000 1183.8000 1161.6000 ;
	    RECT 1185.0000 1160.4000 1186.2001 1161.6000 ;
	    RECT 1182.7500 1158.6000 1183.6500 1160.4000 ;
	    RECT 1182.6000 1157.4000 1183.8000 1158.6000 ;
	    RECT 1180.2001 1154.4000 1181.4000 1155.6000 ;
	    RECT 1185.1500 1152.6000 1186.0500 1160.4000 ;
	    RECT 1189.8000 1157.4000 1191.0000 1158.6000 ;
	    RECT 1185.0000 1151.4000 1186.2001 1152.6000 ;
	    RECT 1180.2001 1085.4000 1181.4000 1086.6000 ;
	    RECT 1180.3500 1065.6000 1181.2500 1085.4000 ;
	    RECT 1182.6000 1073.4000 1183.8000 1074.6000 ;
	    RECT 1182.7500 1065.6000 1183.6500 1073.4000 ;
	    RECT 1192.2001 1067.4000 1193.4000 1068.6000 ;
	    RECT 1180.2001 1064.4000 1181.4000 1065.6000 ;
	    RECT 1182.6000 1064.4000 1183.8000 1065.6000 ;
	    RECT 1187.4000 1064.4000 1188.6000 1065.6000 ;
	    RECT 1187.5500 1062.6000 1188.4501 1064.4000 ;
	    RECT 1192.3500 1062.6000 1193.2500 1067.4000 ;
	    RECT 1187.4000 1061.4000 1188.6000 1062.6000 ;
	    RECT 1192.2001 1061.4000 1193.4000 1062.6000 ;
	    RECT 1187.4000 1035.3000 1188.6000 1043.7001 ;
	    RECT 1189.8000 1043.4000 1191.0000 1044.6000 ;
	    RECT 1189.9501 1041.6000 1190.8500 1043.4000 ;
	    RECT 1189.8000 1040.4000 1191.0000 1041.6000 ;
	    RECT 1192.2001 1029.3000 1193.4000 1046.7001 ;
	    RECT 1197.0000 1043.4000 1198.2001 1044.6000 ;
	    RECT 1197.1500 1038.6000 1198.0500 1043.4000 ;
	    RECT 1197.0000 1037.4000 1198.2001 1038.6000 ;
	    RECT 1201.9501 1026.6000 1202.8500 1217.5500 ;
	    RECT 1204.2001 1217.4000 1205.4000 1217.5500 ;
	    RECT 1213.8000 1209.3000 1215.0000 1226.7001 ;
	    RECT 1216.3500 1146.6000 1217.2500 1289.4000 ;
	    RECT 1218.6000 1277.4000 1219.8000 1278.6000 ;
	    RECT 1221.0000 1266.3000 1222.2001 1286.7001 ;
	    RECT 1223.4000 1266.3000 1224.6000 1286.7001 ;
	    RECT 1225.8000 1269.3000 1227.0000 1286.7001 ;
	    RECT 1228.2001 1280.4000 1229.4000 1281.6000 ;
	    RECT 1228.3500 1266.6000 1229.2500 1280.4000 ;
	    RECT 1230.6000 1269.3000 1231.8000 1286.7001 ;
	    RECT 1233.0000 1283.4000 1234.2001 1284.6000 ;
	    RECT 1235.4000 1269.3000 1236.6000 1286.7001 ;
	    RECT 1228.2001 1265.4000 1229.4000 1266.6000 ;
	    RECT 1237.8000 1266.3000 1239.0000 1286.7001 ;
	    RECT 1240.2001 1266.3000 1241.4000 1286.7001 ;
	    RECT 1242.6000 1266.3000 1243.8000 1286.7001 ;
	    RECT 1273.8000 1283.4000 1275.0000 1284.6000 ;
	    RECT 1257.0000 1271.4000 1258.2001 1272.6000 ;
	    RECT 1273.9501 1251.6000 1274.8500 1283.4000 ;
	    RECT 1281.1500 1281.6000 1282.0500 1304.4000 ;
	    RECT 1281.0000 1280.4000 1282.2001 1281.6000 ;
	    RECT 1283.5500 1278.6000 1284.4501 1334.4000 ;
	    RECT 1302.7500 1326.6000 1303.6500 1361.4000 ;
	    RECT 1305.0000 1356.3000 1306.2001 1376.7001 ;
	    RECT 1307.4000 1356.3000 1308.6000 1376.7001 ;
	    RECT 1312.3500 1374.6000 1313.2500 1424.4000 ;
	    RECT 1317.0000 1403.4000 1318.2001 1404.6000 ;
	    RECT 1314.6000 1400.4000 1315.8000 1401.6000 ;
	    RECT 1314.7500 1386.6000 1315.6500 1400.4000 ;
	    RECT 1314.6000 1385.4000 1315.8000 1386.6000 ;
	    RECT 1309.8000 1356.3000 1311.0000 1373.7001 ;
	    RECT 1312.2001 1373.4000 1313.4000 1374.6000 ;
	    RECT 1312.2001 1361.4000 1313.4000 1362.6000 ;
	    RECT 1314.6000 1356.3000 1315.8000 1373.7001 ;
	    RECT 1317.1500 1359.6000 1318.0500 1403.4000 ;
	    RECT 1331.5500 1398.6000 1332.4501 1457.4000 ;
	    RECT 1333.9501 1431.6000 1334.8500 1463.4000 ;
	    RECT 1374.6000 1460.4000 1375.8000 1461.6000 ;
	    RECT 1333.8000 1430.4000 1335.0000 1431.6000 ;
	    RECT 1348.2001 1400.4000 1349.4000 1401.6000 ;
	    RECT 1331.4000 1397.4000 1332.6000 1398.6000 ;
	    RECT 1341.0000 1397.4000 1342.2001 1398.6000 ;
	    RECT 1345.8000 1397.4000 1347.0000 1398.6000 ;
	    RECT 1317.0000 1358.4000 1318.2001 1359.6000 ;
	    RECT 1319.4000 1356.3000 1320.6000 1373.7001 ;
	    RECT 1321.8000 1356.3000 1323.0000 1376.7001 ;
	    RECT 1324.2001 1356.3000 1325.4000 1376.7001 ;
	    RECT 1326.6000 1356.3000 1327.8000 1376.7001 ;
	    RECT 1329.0000 1367.4000 1330.2001 1368.6000 ;
	    RECT 1309.8000 1349.4000 1311.0000 1350.6000 ;
	    RECT 1309.9501 1341.6000 1310.8500 1349.4000 ;
	    RECT 1309.8000 1340.4000 1311.0000 1341.6000 ;
	    RECT 1302.6000 1325.4000 1303.8000 1326.6000 ;
	    RECT 1285.8000 1307.4000 1287.0000 1308.6000 ;
	    RECT 1297.8000 1301.4000 1299.0000 1302.6000 ;
	    RECT 1326.6000 1301.4000 1327.8000 1302.6000 ;
	    RECT 1283.4000 1277.4000 1284.6000 1278.6000 ;
	    RECT 1295.4000 1274.4000 1296.6000 1275.6000 ;
	    RECT 1273.8000 1250.4000 1275.0000 1251.6000 ;
	    RECT 1295.5500 1230.6000 1296.4501 1274.4000 ;
	    RECT 1297.9501 1242.6000 1298.8500 1301.4000 ;
	    RECT 1300.2001 1298.4000 1301.4000 1299.6000 ;
	    RECT 1300.3500 1284.4501 1301.2500 1298.4000 ;
	    RECT 1300.3500 1283.5500 1303.6500 1284.4501 ;
	    RECT 1302.7500 1272.6000 1303.6500 1283.5500 ;
	    RECT 1326.7500 1281.6000 1327.6500 1301.4000 ;
	    RECT 1326.6000 1280.4000 1327.8000 1281.6000 ;
	    RECT 1302.6000 1271.4000 1303.8000 1272.6000 ;
	    RECT 1302.7500 1254.6000 1303.6500 1271.4000 ;
	    RECT 1326.7500 1260.6000 1327.6500 1280.4000 ;
	    RECT 1326.6000 1259.4000 1327.8000 1260.6000 ;
	    RECT 1302.6000 1253.4000 1303.8000 1254.6000 ;
	    RECT 1297.8000 1241.4000 1299.0000 1242.6000 ;
	    RECT 1305.0000 1236.3000 1306.2001 1256.7001 ;
	    RECT 1307.4000 1236.3000 1308.6000 1256.7001 ;
	    RECT 1309.8000 1236.3000 1311.0000 1256.7001 ;
	    RECT 1312.2001 1236.3000 1313.4000 1253.7001 ;
	    RECT 1314.6000 1238.4000 1315.8000 1239.6000 ;
	    RECT 1233.0000 1229.4000 1234.2001 1230.6000 ;
	    RECT 1295.4000 1229.4000 1296.6000 1230.6000 ;
	    RECT 1233.1500 1224.6000 1234.0500 1229.4000 ;
	    RECT 1233.0000 1223.4000 1234.2001 1224.6000 ;
	    RECT 1221.0000 1217.4000 1222.2001 1218.6000 ;
	    RECT 1216.2001 1145.4000 1217.4000 1146.6000 ;
	    RECT 1216.2001 1127.4000 1217.4000 1128.6000 ;
	    RECT 1216.3500 1125.6000 1217.2500 1127.4000 ;
	    RECT 1216.2001 1124.4000 1217.4000 1125.6000 ;
	    RECT 1218.6000 1109.4000 1219.8000 1110.6000 ;
	    RECT 1213.8000 1067.4000 1215.0000 1068.6000 ;
	    RECT 1213.9501 1065.6000 1214.8500 1067.4000 ;
	    RECT 1213.8000 1064.4000 1215.0000 1065.6000 ;
	    RECT 1213.9501 1062.6000 1214.8500 1064.4000 ;
	    RECT 1209.0000 1061.4000 1210.2001 1062.6000 ;
	    RECT 1213.8000 1061.4000 1215.0000 1062.6000 ;
	    RECT 1209.1500 1059.6000 1210.0500 1061.4000 ;
	    RECT 1209.0000 1058.4000 1210.2001 1059.6000 ;
	    RECT 1206.6000 1029.3000 1207.8000 1046.7001 ;
	    RECT 1209.1500 1038.6000 1210.0500 1058.4000 ;
	    RECT 1216.2001 1043.4000 1217.4000 1044.6000 ;
	    RECT 1216.3500 1041.6000 1217.2500 1043.4000 ;
	    RECT 1216.2001 1040.4000 1217.4000 1041.6000 ;
	    RECT 1209.0000 1037.4000 1210.2001 1038.6000 ;
	    RECT 1201.8000 1025.4000 1203.0000 1026.6000 ;
	    RECT 1206.6000 1025.4000 1207.8000 1026.6000 ;
	    RECT 1204.2001 1007.4000 1205.4000 1008.6000 ;
	    RECT 1201.8000 1001.4000 1203.0000 1002.6000 ;
	    RECT 1201.9501 981.6000 1202.8500 1001.4000 ;
	    RECT 1189.8000 980.4000 1191.0000 981.6000 ;
	    RECT 1201.8000 980.4000 1203.0000 981.6000 ;
	    RECT 1189.9501 942.6000 1190.8500 980.4000 ;
	    RECT 1204.3500 975.6000 1205.2500 1007.4000 ;
	    RECT 1206.7500 990.6000 1207.6500 1025.4000 ;
	    RECT 1209.0000 996.3000 1210.2001 1016.7000 ;
	    RECT 1211.4000 996.3000 1212.6000 1016.7000 ;
	    RECT 1213.8000 996.3000 1215.0000 1016.7000 ;
	    RECT 1216.2001 996.3000 1217.4000 1013.7000 ;
	    RECT 1218.7500 999.6000 1219.6500 1109.4000 ;
	    RECT 1221.1500 1026.6000 1222.0500 1217.4000 ;
	    RECT 1233.1500 1212.6000 1234.0500 1223.4000 ;
	    RECT 1233.0000 1211.4000 1234.2001 1212.6000 ;
	    RECT 1233.1500 1191.6000 1234.0500 1211.4000 ;
	    RECT 1309.8000 1199.4000 1311.0000 1200.6000 ;
	    RECT 1233.0000 1190.4000 1234.2001 1191.6000 ;
	    RECT 1257.0000 1187.4000 1258.2001 1188.6000 ;
	    RECT 1223.4000 1160.4000 1224.6000 1161.6000 ;
	    RECT 1223.5500 1140.6000 1224.4501 1160.4000 ;
	    RECT 1228.2001 1145.4000 1229.4000 1146.6000 ;
	    RECT 1223.4000 1139.4000 1224.6000 1140.6000 ;
	    RECT 1223.5500 1128.6000 1224.4501 1139.4000 ;
	    RECT 1223.4000 1127.4000 1224.6000 1128.6000 ;
	    RECT 1228.3500 1125.6000 1229.2500 1145.4000 ;
	    RECT 1228.2001 1124.4000 1229.4000 1125.6000 ;
	    RECT 1228.2001 1121.4000 1229.4000 1122.6000 ;
	    RECT 1223.4000 1103.4000 1224.6000 1104.6000 ;
	    RECT 1223.5500 1092.6000 1224.4501 1103.4000 ;
	    RECT 1228.3500 1098.6000 1229.2500 1121.4000 ;
	    RECT 1230.6000 1116.3000 1231.8000 1136.7001 ;
	    RECT 1233.0000 1116.3000 1234.2001 1136.7001 ;
	    RECT 1235.4000 1116.3000 1236.6000 1133.7001 ;
	    RECT 1237.8000 1121.4000 1239.0000 1122.6000 ;
	    RECT 1240.2001 1116.3000 1241.4000 1133.7001 ;
	    RECT 1242.6000 1118.4000 1243.8000 1119.6000 ;
	    RECT 1242.7500 1110.6000 1243.6500 1118.4000 ;
	    RECT 1245.0000 1116.3000 1246.2001 1133.7001 ;
	    RECT 1247.4000 1116.3000 1248.6000 1136.7001 ;
	    RECT 1249.8000 1116.3000 1251.0000 1136.7001 ;
	    RECT 1252.2001 1116.3000 1253.4000 1136.7001 ;
	    RECT 1242.6000 1109.4000 1243.8000 1110.6000 ;
	    RECT 1242.7500 1104.6000 1243.6500 1109.4000 ;
	    RECT 1242.6000 1103.4000 1243.8000 1104.6000 ;
	    RECT 1228.2001 1097.4000 1229.4000 1098.6000 ;
	    RECT 1223.4000 1091.4000 1224.6000 1092.6000 ;
	    RECT 1242.6000 1073.4000 1243.8000 1074.6000 ;
	    RECT 1247.4000 1073.4000 1248.6000 1074.6000 ;
	    RECT 1242.7500 1065.6000 1243.6500 1073.4000 ;
	    RECT 1247.5500 1068.6000 1248.4501 1073.4000 ;
	    RECT 1247.4000 1068.4501 1248.6000 1068.6000 ;
	    RECT 1245.1500 1067.5500 1248.6000 1068.4501 ;
	    RECT 1242.6000 1064.4000 1243.8000 1065.6000 ;
	    RECT 1237.8000 1043.4000 1239.0000 1044.6000 ;
	    RECT 1223.4000 1037.4000 1224.6000 1038.6000 ;
	    RECT 1221.0000 1025.4000 1222.2001 1026.6000 ;
	    RECT 1223.5500 1014.6000 1224.4501 1037.4000 ;
	    RECT 1237.9501 1035.6000 1238.8500 1043.4000 ;
	    RECT 1245.1500 1041.6000 1246.0500 1067.5500 ;
	    RECT 1247.4000 1067.4000 1248.6000 1067.5500 ;
	    RECT 1247.4000 1061.4000 1248.6000 1062.6000 ;
	    RECT 1249.8000 1061.4000 1251.0000 1062.6000 ;
	    RECT 1247.5500 1044.6000 1248.4501 1061.4000 ;
	    RECT 1247.4000 1043.4000 1248.6000 1044.6000 ;
	    RECT 1245.0000 1040.4000 1246.2001 1041.6000 ;
	    RECT 1245.0000 1037.4000 1246.2001 1038.6000 ;
	    RECT 1237.8000 1034.4000 1239.0000 1035.6000 ;
	    RECT 1218.6000 998.4000 1219.8000 999.6000 ;
	    RECT 1206.6000 989.4000 1207.8000 990.6000 ;
	    RECT 1199.4000 974.4000 1200.6000 975.6000 ;
	    RECT 1204.2001 974.4000 1205.4000 975.6000 ;
	    RECT 1199.5500 966.6000 1200.4501 974.4000 ;
	    RECT 1199.4000 965.4000 1200.6000 966.6000 ;
	    RECT 1189.8000 941.4000 1191.0000 942.6000 ;
	    RECT 1189.9501 900.6000 1190.8500 941.4000 ;
	    RECT 1218.7500 906.6000 1219.6500 998.4000 ;
	    RECT 1221.0000 996.3000 1222.2001 1013.7000 ;
	    RECT 1223.4000 1013.4000 1224.6000 1014.6000 ;
	    RECT 1223.4000 1001.4000 1224.6000 1002.6000 ;
	    RECT 1225.8000 996.3000 1227.0000 1013.7000 ;
	    RECT 1228.2001 996.3000 1229.4000 1016.7000 ;
	    RECT 1230.6000 996.3000 1231.8000 1016.7000 ;
	    RECT 1237.8000 1016.4000 1239.0000 1017.6000 ;
	    RECT 1237.9501 1011.4500 1238.8500 1016.4000 ;
	    RECT 1235.5500 1010.5500 1238.8500 1011.4500 ;
	    RECT 1233.0000 1004.4000 1234.2001 1005.6000 ;
	    RECT 1233.1500 996.6000 1234.0500 1004.4000 ;
	    RECT 1233.0000 995.4000 1234.2001 996.6000 ;
	    RECT 1221.0000 989.4000 1222.2001 990.6000 ;
	    RECT 1209.0000 905.4000 1210.2001 906.6000 ;
	    RECT 1218.6000 905.4000 1219.8000 906.6000 ;
	    RECT 1189.8000 899.4000 1191.0000 900.6000 ;
	    RECT 1194.6000 899.4000 1195.8000 900.6000 ;
	    RECT 1189.9501 888.6000 1190.8500 899.4000 ;
	    RECT 1189.8000 887.4000 1191.0000 888.6000 ;
	    RECT 1194.7500 885.6000 1195.6500 899.4000 ;
	    RECT 1194.6000 884.4000 1195.8000 885.6000 ;
	    RECT 1177.8000 857.4000 1179.0000 858.6000 ;
	    RECT 1182.6000 854.4000 1183.8000 855.6000 ;
	    RECT 1182.7500 846.6000 1183.6500 854.4000 ;
	    RECT 1182.6000 845.4000 1183.8000 846.6000 ;
	    RECT 1177.8000 839.4000 1179.0000 840.6000 ;
	    RECT 1163.4000 818.4000 1164.6000 819.6000 ;
	    RECT 1151.4000 800.4000 1152.6000 801.6000 ;
	    RECT 1158.6000 800.4000 1159.8000 801.6000 ;
	    RECT 1139.4000 797.4000 1140.6000 798.6000 ;
	    RECT 1139.5500 792.6000 1140.4501 797.4000 ;
	    RECT 1144.2001 794.4000 1145.4000 795.6000 ;
	    RECT 1139.4000 791.4000 1140.6000 792.6000 ;
	    RECT 1134.6000 767.4000 1135.8000 768.6000 ;
	    RECT 1120.2001 677.4000 1121.4000 678.6000 ;
	    RECT 1120.3500 660.6000 1121.2500 677.4000 ;
	    RECT 1125.0000 674.4000 1126.2001 675.6000 ;
	    RECT 1125.1500 672.6000 1126.0500 674.4000 ;
	    RECT 1125.0000 671.4000 1126.2001 672.6000 ;
	    RECT 1125.1500 666.6000 1126.0500 671.4000 ;
	    RECT 1125.0000 665.4000 1126.2001 666.6000 ;
	    RECT 1120.2001 659.4000 1121.4000 660.6000 ;
	    RECT 1134.7500 648.6000 1135.6500 767.4000 ;
	    RECT 1144.3500 765.6000 1145.2500 794.4000 ;
	    RECT 1158.7500 780.6000 1159.6500 800.4000 ;
	    RECT 1151.4000 779.4000 1152.6000 780.6000 ;
	    RECT 1158.6000 779.4000 1159.8000 780.6000 ;
	    RECT 1144.2001 764.4000 1145.4000 765.6000 ;
	    RECT 1151.5500 762.6000 1152.4501 779.4000 ;
	    RECT 1161.0000 764.4000 1162.2001 765.6000 ;
	    RECT 1144.2001 761.4000 1145.4000 762.6000 ;
	    RECT 1151.4000 761.4000 1152.6000 762.6000 ;
	    RECT 1144.3500 756.6000 1145.2500 761.4000 ;
	    RECT 1144.2001 755.4000 1145.4000 756.6000 ;
	    RECT 1134.6000 647.4000 1135.8000 648.6000 ;
	    RECT 1110.6000 641.4000 1111.8000 642.6000 ;
	    RECT 1117.8000 641.4000 1119.0000 642.6000 ;
	    RECT 1117.9501 630.6000 1118.8500 641.4000 ;
	    RECT 1103.5500 629.5500 1106.8500 630.4500 ;
	    RECT 1093.8000 606.3000 1095.0000 626.7000 ;
	    RECT 1096.2001 606.3000 1097.4000 626.7000 ;
	    RECT 1098.6000 606.3000 1099.8000 626.7000 ;
	    RECT 1101.0000 609.3000 1102.2001 626.7000 ;
	    RECT 1103.5500 624.6000 1104.4501 629.5500 ;
	    RECT 1117.8000 629.4000 1119.0000 630.6000 ;
	    RECT 1103.4000 623.4000 1104.6000 624.6000 ;
	    RECT 1105.8000 609.3000 1107.0000 626.7000 ;
	    RECT 1108.2001 623.4000 1109.4000 624.6000 ;
	    RECT 1108.3500 621.6000 1109.2500 623.4000 ;
	    RECT 1108.2001 620.4000 1109.4000 621.6000 ;
	    RECT 1108.2001 611.4000 1109.4000 612.6000 ;
	    RECT 1101.0000 605.4000 1102.2001 606.6000 ;
	    RECT 1096.2001 593.4000 1097.4000 594.6000 ;
	    RECT 1093.8000 569.4000 1095.0000 570.6000 ;
	    RECT 1093.9501 564.6000 1094.8500 569.4000 ;
	    RECT 1091.4000 563.4000 1092.6000 564.6000 ;
	    RECT 1093.8000 563.4000 1095.0000 564.6000 ;
	    RECT 1079.4000 560.4000 1080.6000 561.6000 ;
	    RECT 1079.5500 525.6000 1080.4501 560.4000 ;
	    RECT 1096.3500 558.6000 1097.2500 593.4000 ;
	    RECT 1098.6000 563.4000 1099.8000 564.6000 ;
	    RECT 1098.7500 561.6000 1099.6500 563.4000 ;
	    RECT 1098.6000 560.4000 1099.8000 561.6000 ;
	    RECT 1101.1500 558.6000 1102.0500 605.4000 ;
	    RECT 1103.4000 560.4000 1104.6000 561.6000 ;
	    RECT 1103.5500 558.6000 1104.4501 560.4000 ;
	    RECT 1084.2001 557.4000 1085.4000 558.6000 ;
	    RECT 1096.2001 557.4000 1097.4000 558.6000 ;
	    RECT 1101.0000 557.4000 1102.2001 558.6000 ;
	    RECT 1103.4000 557.4000 1104.6000 558.6000 ;
	    RECT 1079.4000 524.4000 1080.6000 525.6000 ;
	    RECT 1077.0000 521.4000 1078.2001 522.6000 ;
	    RECT 1077.1500 504.6000 1078.0500 521.4000 ;
	    RECT 1077.0000 503.4000 1078.2001 504.6000 ;
	    RECT 1074.6000 491.4000 1075.8000 492.6000 ;
	    RECT 1074.7500 486.6000 1075.6500 491.4000 ;
	    RECT 1074.6000 485.4000 1075.8000 486.6000 ;
	    RECT 1079.5500 465.6000 1080.4501 524.4000 ;
	    RECT 1079.4000 464.4000 1080.6000 465.6000 ;
	    RECT 1084.3500 462.6000 1085.2500 557.4000 ;
	    RECT 1089.0000 539.4000 1090.2001 540.6000 ;
	    RECT 1086.6000 485.4000 1087.8000 486.6000 ;
	    RECT 1084.2001 461.4000 1085.4000 462.6000 ;
	    RECT 1084.3500 456.6000 1085.2500 461.4000 ;
	    RECT 1084.2001 455.4000 1085.4000 456.6000 ;
	    RECT 1084.2001 449.4000 1085.4000 450.6000 ;
	    RECT 1069.8000 443.4000 1071.0000 444.6000 ;
	    RECT 1072.2001 429.3000 1073.4000 446.7000 ;
	    RECT 1074.6000 426.3000 1075.8000 446.7000 ;
	    RECT 1077.0000 426.3000 1078.2001 446.7000 ;
	    RECT 1079.4000 426.3000 1080.6000 446.7000 ;
	    RECT 1084.3500 444.6000 1085.2500 449.4000 ;
	    RECT 1084.2001 443.4000 1085.4000 444.6000 ;
	    RECT 1057.8000 419.4000 1059.0000 420.6000 ;
	    RECT 1065.0000 419.4000 1066.2001 420.6000 ;
	    RECT 1067.4000 419.4000 1068.6000 420.6000 ;
	    RECT 1053.0000 413.4000 1054.2001 414.6000 ;
	    RECT 1036.2001 401.4000 1037.4000 402.6000 ;
	    RECT 1048.2001 401.4000 1049.4000 402.6000 ;
	    RECT 1033.8000 395.4000 1035.0000 396.6000 ;
	    RECT 1033.8000 380.4000 1035.0000 381.6000 ;
	    RECT 1033.9501 360.6000 1034.8500 380.4000 ;
	    RECT 1033.8000 359.4000 1035.0000 360.6000 ;
	    RECT 1036.3500 357.4500 1037.2500 401.4000 ;
	    RECT 1050.6000 389.4000 1051.8000 390.6000 ;
	    RECT 1038.6000 365.4000 1039.8000 366.6000 ;
	    RECT 1024.2001 345.4500 1025.4000 345.6000 ;
	    RECT 1021.9500 344.5500 1025.4000 345.4500 ;
	    RECT 1000.2000 320.4000 1001.4000 321.6000 ;
	    RECT 1005.0000 320.4000 1006.2000 321.6000 ;
	    RECT 997.8000 317.4000 999.0000 318.6000 ;
	    RECT 990.7500 308.5500 994.0500 309.4500 ;
	    RECT 990.6000 276.3000 991.8000 293.7000 ;
	    RECT 993.1500 282.6000 994.0500 308.5500 ;
	    RECT 1000.3500 306.6000 1001.2500 320.4000 ;
	    RECT 1005.1500 318.6000 1006.0500 320.4000 ;
	    RECT 1002.6000 317.4000 1003.8000 318.6000 ;
	    RECT 1005.0000 317.4000 1006.2000 318.6000 ;
	    RECT 1014.6000 317.4000 1015.8000 318.6000 ;
	    RECT 1000.2000 305.4000 1001.4000 306.6000 ;
	    RECT 993.0000 281.4000 994.2000 282.6000 ;
	    RECT 995.4000 279.3000 996.6000 287.7000 ;
	    RECT 988.2000 248.4000 989.4000 249.6000 ;
	    RECT 988.2000 245.4000 989.4000 246.6000 ;
	    RECT 983.4000 170.4000 984.6000 171.6000 ;
	    RECT 981.0000 119.4000 982.2000 120.6000 ;
	    RECT 983.4000 113.4000 984.6000 114.6000 ;
	    RECT 983.5500 111.6000 984.4500 113.4000 ;
	    RECT 983.4000 110.4000 984.6000 111.6000 ;
	    RECT 978.6000 74.4000 979.8000 75.6000 ;
	    RECT 973.8000 65.4000 975.0000 66.6000 ;
	    RECT 957.0000 36.3000 958.2000 53.7000 ;
	    RECT 959.4000 41.4000 960.6000 42.6000 ;
	    RECT 959.5500 39.6000 960.4500 41.4000 ;
	    RECT 959.4000 38.4000 960.6000 39.6000 ;
	    RECT 959.5500 30.6000 960.4500 38.4000 ;
	    RECT 961.8000 36.3000 963.0000 53.7000 ;
	    RECT 964.2000 53.4000 965.4000 54.6000 ;
	    RECT 964.2000 41.4000 965.4000 42.6000 ;
	    RECT 959.4000 29.4000 960.6000 30.6000 ;
	    RECT 964.3500 21.6000 965.2500 41.4000 ;
	    RECT 966.6000 36.3000 967.8000 53.7000 ;
	    RECT 969.0000 36.3000 970.2000 56.7000 ;
	    RECT 971.4000 36.3000 972.6000 56.7000 ;
	    RECT 973.9500 45.6000 974.8500 65.4000 ;
	    RECT 978.6000 56.4000 979.8000 57.6000 ;
	    RECT 978.7500 48.6000 979.6500 56.4000 ;
	    RECT 978.6000 47.4000 979.8000 48.6000 ;
	    RECT 973.8000 44.4000 975.0000 45.6000 ;
	    RECT 839.4000 20.4000 840.6000 21.6000 ;
	    RECT 885.0000 20.4000 886.2000 21.6000 ;
	    RECT 964.2000 20.4000 965.4000 21.6000 ;
	    RECT 988.3500 18.6000 989.2500 245.4000 ;
	    RECT 997.8000 224.4000 999.0000 225.6000 ;
	    RECT 995.4000 221.4000 996.6000 222.6000 ;
	    RECT 995.5500 204.6000 996.4500 221.4000 ;
	    RECT 995.4000 203.4000 996.6000 204.6000 ;
	    RECT 995.5500 201.6000 996.4500 203.4000 ;
	    RECT 995.4000 200.4000 996.6000 201.6000 ;
	    RECT 997.9500 198.6000 998.8500 224.4000 ;
	    RECT 1002.7500 222.6000 1003.6500 317.4000 ;
	    RECT 1014.7500 282.6000 1015.6500 317.4000 ;
	    RECT 1019.4000 305.4000 1020.6000 306.6000 ;
	    RECT 1019.5500 288.6000 1020.4500 305.4000 ;
	    RECT 1019.4000 287.4000 1020.6000 288.6000 ;
	    RECT 1014.6000 281.4000 1015.8000 282.6000 ;
	    RECT 1021.9500 270.6000 1022.8500 344.5500 ;
	    RECT 1024.2001 344.4000 1025.4000 344.5500 ;
	    RECT 1026.6000 336.3000 1027.8000 356.7000 ;
	    RECT 1029.0000 336.3000 1030.2001 356.7000 ;
	    RECT 1033.9501 356.5500 1037.2500 357.4500 ;
	    RECT 1031.4000 336.3000 1032.6000 353.7000 ;
	    RECT 1033.9501 342.6000 1034.8500 356.5500 ;
	    RECT 1033.8000 341.4000 1035.0000 342.6000 ;
	    RECT 1036.2001 336.3000 1037.4000 353.7000 ;
	    RECT 1038.7500 339.6000 1039.6500 365.4000 ;
	    RECT 1038.6000 338.4000 1039.8000 339.6000 ;
	    RECT 1041.0000 336.3000 1042.2001 353.7000 ;
	    RECT 1043.4000 336.3000 1044.6000 356.7000 ;
	    RECT 1045.8000 336.3000 1047.0000 356.7000 ;
	    RECT 1048.2001 336.3000 1049.4000 356.7000 ;
	    RECT 1038.6000 329.4000 1039.8000 330.6000 ;
	    RECT 1038.7500 318.6000 1039.6500 329.4000 ;
	    RECT 1041.0000 323.4000 1042.2001 324.6000 ;
	    RECT 1041.1500 321.6000 1042.0500 323.4000 ;
	    RECT 1050.7500 321.6000 1051.6500 389.4000 ;
	    RECT 1057.9501 381.6000 1058.8500 419.4000 ;
	    RECT 1060.2001 398.4000 1061.4000 399.6000 ;
	    RECT 1057.8000 380.4000 1059.0000 381.6000 ;
	    RECT 1060.3500 360.6000 1061.2500 398.4000 ;
	    RECT 1067.5500 381.6000 1068.4501 419.4000 ;
	    RECT 1079.4000 401.4000 1080.6000 402.6000 ;
	    RECT 1067.4000 380.4000 1068.6000 381.6000 ;
	    RECT 1060.2001 359.4000 1061.4000 360.6000 ;
	    RECT 1060.3500 351.4500 1061.2500 359.4000 ;
	    RECT 1062.6000 351.4500 1063.8000 351.6000 ;
	    RECT 1060.3500 350.5500 1063.8000 351.4500 ;
	    RECT 1062.6000 350.4000 1063.8000 350.5500 ;
	    RECT 1041.0000 320.4000 1042.2001 321.6000 ;
	    RECT 1050.6000 320.4000 1051.8000 321.6000 ;
	    RECT 1033.8000 317.4000 1035.0000 318.6000 ;
	    RECT 1038.6000 317.4000 1039.8000 318.6000 ;
	    RECT 1033.9501 294.6000 1034.8500 317.4000 ;
	    RECT 1062.7500 315.6000 1063.6500 350.4000 ;
	    RECT 1077.0000 329.4000 1078.2001 330.6000 ;
	    RECT 1077.1500 327.6000 1078.0500 329.4000 ;
	    RECT 1077.0000 326.4000 1078.2001 327.6000 ;
	    RECT 1069.8000 317.4000 1071.0000 318.6000 ;
	    RECT 1043.4000 314.4000 1044.6000 315.6000 ;
	    RECT 1062.6000 314.4000 1063.8000 315.6000 ;
	    RECT 1033.8000 293.4000 1035.0000 294.6000 ;
	    RECT 1043.5500 288.6000 1044.4501 314.4000 ;
	    RECT 1072.2001 311.4000 1073.4000 312.6000 ;
	    RECT 1048.2001 305.4000 1049.4000 306.6000 ;
	    RECT 1048.3500 294.6000 1049.2500 305.4000 ;
	    RECT 1072.3500 300.6000 1073.2500 311.4000 ;
	    RECT 1072.2001 299.4000 1073.4000 300.6000 ;
	    RECT 1048.2001 293.4000 1049.4000 294.6000 ;
	    RECT 1048.3500 291.6000 1049.2500 293.4000 ;
	    RECT 1045.8000 290.4000 1047.0000 291.6000 ;
	    RECT 1048.2001 290.4000 1049.4000 291.6000 ;
	    RECT 1043.4000 287.4000 1044.6000 288.6000 ;
	    RECT 1041.0000 284.4000 1042.2001 285.6000 ;
	    RECT 1012.2000 269.4000 1013.4000 270.6000 ;
	    RECT 1021.8000 269.4000 1023.0000 270.6000 ;
	    RECT 1012.3500 258.6000 1013.2500 269.4000 ;
	    RECT 1012.2000 257.4000 1013.4000 258.6000 ;
	    RECT 1007.4000 254.4000 1008.6000 255.6000 ;
	    RECT 1007.5500 246.6000 1008.4500 254.4000 ;
	    RECT 1007.4000 245.4000 1008.6000 246.6000 ;
	    RECT 1005.0000 233.4000 1006.2000 234.6000 ;
	    RECT 1005.1500 225.6000 1006.0500 233.4000 ;
	    RECT 1005.0000 224.4000 1006.2000 225.6000 ;
	    RECT 1002.6000 221.4000 1003.8000 222.6000 ;
	    RECT 997.8000 197.4000 999.0000 198.6000 ;
	    RECT 1002.6000 194.4000 1003.8000 195.6000 ;
	    RECT 1002.7500 186.6000 1003.6500 194.4000 ;
	    RECT 1002.6000 185.4000 1003.8000 186.6000 ;
	    RECT 993.0000 173.4000 994.2000 174.6000 ;
	    RECT 993.1500 168.6000 994.0500 173.4000 ;
	    RECT 993.0000 167.4000 994.2000 168.6000 ;
	    RECT 997.8000 164.4000 999.0000 165.6000 ;
	    RECT 993.0000 161.4000 994.2000 162.6000 ;
	    RECT 993.1500 144.6000 994.0500 161.4000 ;
	    RECT 993.0000 143.4000 994.2000 144.6000 ;
	    RECT 990.6000 131.4000 991.8000 132.6000 ;
	    RECT 990.7500 84.6000 991.6500 131.4000 ;
	    RECT 990.6000 83.4000 991.8000 84.6000 ;
	    RECT 997.9500 81.6000 998.8500 164.4000 ;
	    RECT 1002.7500 162.6000 1003.6500 185.4000 ;
	    RECT 1000.2000 161.4000 1001.4000 162.6000 ;
	    RECT 1002.6000 161.4000 1003.8000 162.6000 ;
	    RECT 1000.3500 126.6000 1001.2500 161.4000 ;
	    RECT 1002.6000 149.4000 1003.8000 150.6000 ;
	    RECT 1000.2000 125.4000 1001.4000 126.6000 ;
	    RECT 1002.7500 99.6000 1003.6500 149.4000 ;
	    RECT 1012.3500 138.4500 1013.2500 257.4000 ;
	    RECT 1014.6000 246.3000 1015.8000 266.7000 ;
	    RECT 1017.0000 246.3000 1018.2000 266.7000 ;
	    RECT 1019.4000 249.3000 1020.6000 266.7000 ;
	    RECT 1021.8000 263.4000 1023.0000 264.6000 ;
	    RECT 1021.9500 261.6000 1022.8500 263.4000 ;
	    RECT 1021.8000 260.4000 1023.0000 261.6000 ;
	    RECT 1024.2001 249.3000 1025.4000 266.7000 ;
	    RECT 1026.6000 263.4000 1027.8000 264.6000 ;
	    RECT 1017.0000 224.4000 1018.2000 225.6000 ;
	    RECT 1014.6000 215.4000 1015.8000 216.6000 ;
	    RECT 1014.7500 204.6000 1015.6500 215.4000 ;
	    RECT 1014.6000 203.4000 1015.8000 204.6000 ;
	    RECT 1014.6000 200.4000 1015.8000 201.6000 ;
	    RECT 1014.7500 180.6000 1015.6500 200.4000 ;
	    RECT 1014.6000 179.4000 1015.8000 180.6000 ;
	    RECT 1017.1500 159.6000 1018.0500 224.4000 ;
	    RECT 1024.2001 221.4000 1025.4000 222.6000 ;
	    RECT 1026.7500 222.4500 1027.6500 263.4000 ;
	    RECT 1029.0000 249.3000 1030.2001 266.7000 ;
	    RECT 1031.4000 246.3000 1032.6000 266.7000 ;
	    RECT 1033.8000 246.3000 1035.0000 266.7000 ;
	    RECT 1036.2001 246.3000 1037.4000 266.7000 ;
	    RECT 1041.1500 264.6000 1042.0500 284.4000 ;
	    RECT 1043.5500 282.6000 1044.4501 287.4000 ;
	    RECT 1045.9501 285.6000 1046.8500 290.4000 ;
	    RECT 1067.4000 287.4000 1068.6000 288.6000 ;
	    RECT 1045.8000 284.4000 1047.0000 285.6000 ;
	    RECT 1043.4000 281.4000 1044.6000 282.6000 ;
	    RECT 1041.0000 263.4000 1042.2001 264.6000 ;
	    RECT 1053.0000 260.4000 1054.2001 261.6000 ;
	    RECT 1050.6000 251.4000 1051.8000 252.6000 ;
	    RECT 1029.0000 227.4000 1030.2001 228.6000 ;
	    RECT 1026.7500 221.5500 1030.0500 222.4500 ;
	    RECT 1024.3500 204.6000 1025.2500 221.4000 ;
	    RECT 1024.2001 203.4000 1025.4000 204.6000 ;
	    RECT 1017.0000 158.4000 1018.2000 159.6000 ;
	    RECT 1014.6000 138.4500 1015.8000 138.6000 ;
	    RECT 1012.3500 137.5500 1015.8000 138.4500 ;
	    RECT 1009.8000 134.4000 1011.0000 135.6000 ;
	    RECT 1009.9500 126.6000 1010.8500 134.4000 ;
	    RECT 1009.8000 125.4000 1011.0000 126.6000 ;
	    RECT 1012.3500 108.6000 1013.2500 137.5500 ;
	    RECT 1014.6000 137.4000 1015.8000 137.5500 ;
	    RECT 1017.0000 126.3000 1018.2000 146.7000 ;
	    RECT 1019.4000 126.3000 1020.6000 146.7000 ;
	    RECT 1021.8000 129.3000 1023.0000 146.7000 ;
	    RECT 1024.2001 143.4000 1025.4000 144.6000 ;
	    RECT 1024.3500 141.6000 1025.2500 143.4000 ;
	    RECT 1024.2001 140.4000 1025.4000 141.6000 ;
	    RECT 1026.6000 129.3000 1027.8000 146.7000 ;
	    RECT 1029.1500 144.6000 1030.0500 221.5500 ;
	    RECT 1033.8000 221.4000 1035.0000 222.6000 ;
	    RECT 1041.0000 200.4000 1042.2001 201.6000 ;
	    RECT 1041.1500 195.6000 1042.0500 200.4000 ;
	    RECT 1045.8000 197.4000 1047.0000 198.6000 ;
	    RECT 1041.0000 194.4000 1042.2001 195.6000 ;
	    RECT 1033.8000 191.4000 1035.0000 192.6000 ;
	    RECT 1033.9501 168.6000 1034.8500 191.4000 ;
	    RECT 1041.1500 174.6000 1042.0500 194.4000 ;
	    RECT 1045.9501 186.6000 1046.8500 197.4000 ;
	    RECT 1050.7500 192.6000 1051.6500 251.4000 ;
	    RECT 1053.1500 234.6000 1054.0500 260.4000 ;
	    RECT 1053.0000 233.4000 1054.2001 234.6000 ;
	    RECT 1067.5500 228.6000 1068.4501 287.4000 ;
	    RECT 1069.8000 281.4000 1071.0000 282.6000 ;
	    RECT 1069.9501 279.6000 1070.8500 281.4000 ;
	    RECT 1069.8000 278.4000 1071.0000 279.6000 ;
	    RECT 1079.5500 264.6000 1080.4501 401.4000 ;
	    RECT 1081.8000 395.4000 1083.0000 396.6000 ;
	    RECT 1081.9501 348.6000 1082.8500 395.4000 ;
	    RECT 1081.8000 347.4000 1083.0000 348.6000 ;
	    RECT 1084.2001 347.4000 1085.4000 348.6000 ;
	    RECT 1081.9501 318.6000 1082.8500 347.4000 ;
	    RECT 1084.3500 324.6000 1085.2500 347.4000 ;
	    RECT 1084.2001 323.4000 1085.4000 324.6000 ;
	    RECT 1081.8000 317.4000 1083.0000 318.6000 ;
	    RECT 1072.2001 263.4000 1073.4000 264.6000 ;
	    RECT 1079.4000 263.4000 1080.6000 264.6000 ;
	    RECT 1072.3500 258.6000 1073.2500 263.4000 ;
	    RECT 1072.2001 257.4000 1073.4000 258.6000 ;
	    RECT 1079.4000 245.4000 1080.6000 246.6000 ;
	    RECT 1067.4000 228.4500 1068.6000 228.6000 ;
	    RECT 1067.4000 227.5500 1070.8500 228.4500 ;
	    RECT 1067.4000 227.4000 1068.6000 227.5500 ;
	    RECT 1060.2001 224.4000 1061.4000 225.6000 ;
	    RECT 1057.8000 221.4000 1059.0000 222.6000 ;
	    RECT 1048.2001 191.4000 1049.4000 192.6000 ;
	    RECT 1050.6000 191.4000 1051.8000 192.6000 ;
	    RECT 1045.8000 185.4000 1047.0000 186.6000 ;
	    RECT 1041.0000 173.4000 1042.2001 174.6000 ;
	    RECT 1048.3500 171.6000 1049.2500 191.4000 ;
	    RECT 1048.2001 170.4000 1049.4000 171.6000 ;
	    RECT 1057.9501 168.6000 1058.8500 221.4000 ;
	    RECT 1060.3500 216.6000 1061.2500 224.4000 ;
	    RECT 1060.2001 215.4000 1061.4000 216.6000 ;
	    RECT 1067.4000 173.4000 1068.6000 174.6000 ;
	    RECT 1033.8000 167.4000 1035.0000 168.6000 ;
	    RECT 1057.8000 167.4000 1059.0000 168.6000 ;
	    RECT 1067.5500 165.6000 1068.4501 173.4000 ;
	    RECT 1069.9501 171.6000 1070.8500 227.5500 ;
	    RECT 1079.5500 222.6000 1080.4501 245.4000 ;
	    RECT 1081.9501 228.6000 1082.8500 317.4000 ;
	    RECT 1084.2001 299.4000 1085.4000 300.6000 ;
	    RECT 1084.3500 294.6000 1085.2500 299.4000 ;
	    RECT 1084.2001 293.4000 1085.4000 294.6000 ;
	    RECT 1084.3500 285.6000 1085.2500 293.4000 ;
	    RECT 1084.2001 284.4000 1085.4000 285.6000 ;
	    RECT 1084.3500 264.6000 1085.2500 284.4000 ;
	    RECT 1084.2001 263.4000 1085.4000 264.6000 ;
	    RECT 1081.8000 227.4000 1083.0000 228.6000 ;
	    RECT 1079.4000 221.4000 1080.6000 222.6000 ;
	    RECT 1077.0000 203.4000 1078.2001 204.6000 ;
	    RECT 1077.1500 198.6000 1078.0500 203.4000 ;
	    RECT 1077.0000 197.4000 1078.2001 198.6000 ;
	    RECT 1077.0000 194.4000 1078.2001 195.6000 ;
	    RECT 1077.1500 192.6000 1078.0500 194.4000 ;
	    RECT 1077.0000 191.4000 1078.2001 192.6000 ;
	    RECT 1079.4000 191.4000 1080.6000 192.6000 ;
	    RECT 1079.5500 171.6000 1080.4501 191.4000 ;
	    RECT 1069.8000 170.4000 1071.0000 171.6000 ;
	    RECT 1079.4000 170.4000 1080.6000 171.6000 ;
	    RECT 1050.6000 164.4000 1051.8000 165.6000 ;
	    RECT 1067.4000 164.4000 1068.6000 165.6000 ;
	    RECT 1041.0000 161.4000 1042.2001 162.6000 ;
	    RECT 1029.0000 143.4000 1030.2001 144.6000 ;
	    RECT 1029.1500 138.6000 1030.0500 143.4000 ;
	    RECT 1029.0000 137.4000 1030.2001 138.6000 ;
	    RECT 1031.4000 129.3000 1032.6000 146.7000 ;
	    RECT 1033.8000 126.3000 1035.0000 146.7000 ;
	    RECT 1036.2001 126.3000 1037.4000 146.7000 ;
	    RECT 1038.6000 126.3000 1039.8000 146.7000 ;
	    RECT 1012.2000 107.4000 1013.4000 108.6000 ;
	    RECT 1012.2000 101.4000 1013.4000 102.6000 ;
	    RECT 1002.6000 98.4000 1003.8000 99.6000 ;
	    RECT 997.8000 80.4000 999.0000 81.6000 ;
	    RECT 990.6000 77.4000 991.8000 78.6000 ;
	    RECT 990.7500 48.6000 991.6500 77.4000 ;
	    RECT 990.6000 47.4000 991.8000 48.6000 ;
	    RECT 1012.3500 45.6000 1013.2500 101.4000 ;
	    RECT 1048.2001 71.4000 1049.4000 72.6000 ;
	    RECT 1012.2000 44.4000 1013.4000 45.6000 ;
	    RECT 1007.4000 41.4000 1008.6000 42.6000 ;
	    RECT 1026.6000 41.4000 1027.8000 42.6000 ;
	    RECT 1007.5500 24.6000 1008.4500 41.4000 ;
	    RECT 1007.4000 23.4000 1008.6000 24.6000 ;
	    RECT 801.0000 17.4000 802.2000 18.6000 ;
	    RECT 856.2000 17.4000 857.4000 18.6000 ;
	    RECT 892.2000 17.4000 893.4000 18.6000 ;
	    RECT 988.2000 17.4000 989.4000 18.6000 ;
	    RECT 892.3500 15.6000 893.2500 17.4000 ;
	    RECT 1026.7500 15.6000 1027.6500 41.4000 ;
	    RECT 1048.3500 30.6000 1049.2500 71.4000 ;
	    RECT 1050.7500 42.6000 1051.6500 164.4000 ;
	    RECT 1074.6000 143.4000 1075.8000 144.6000 ;
	    RECT 1074.7500 141.6000 1075.6500 143.4000 ;
	    RECT 1074.6000 140.4000 1075.8000 141.6000 ;
	    RECT 1074.6000 137.4000 1075.8000 138.6000 ;
	    RECT 1079.4000 137.4000 1080.6000 138.6000 ;
	    RECT 1053.0000 131.4000 1054.2001 132.6000 ;
	    RECT 1053.1500 96.6000 1054.0500 131.4000 ;
	    RECT 1069.8000 98.4000 1071.0000 99.6000 ;
	    RECT 1072.2001 99.3000 1073.4000 107.7000 ;
	    RECT 1074.7500 102.6000 1075.6500 137.4000 ;
	    RECT 1079.5500 135.6000 1080.4501 137.4000 ;
	    RECT 1081.9501 135.6000 1082.8500 227.4000 ;
	    RECT 1084.2001 222.4500 1085.4000 222.6000 ;
	    RECT 1086.7500 222.4500 1087.6500 485.4000 ;
	    RECT 1089.1500 381.6000 1090.0500 539.4000 ;
	    RECT 1103.5500 522.6000 1104.4501 557.4000 ;
	    RECT 1105.8000 533.4000 1107.0000 534.6000 ;
	    RECT 1105.9501 525.6000 1106.8500 533.4000 ;
	    RECT 1105.8000 524.4000 1107.0000 525.6000 ;
	    RECT 1091.4000 521.4000 1092.6000 522.6000 ;
	    RECT 1103.4000 521.4000 1104.6000 522.6000 ;
	    RECT 1091.5500 501.6000 1092.4501 521.4000 ;
	    RECT 1108.3500 510.6000 1109.2500 611.4000 ;
	    RECT 1110.6000 609.3000 1111.8000 626.7000 ;
	    RECT 1113.0000 606.3000 1114.2001 626.7000 ;
	    RECT 1115.4000 606.3000 1116.6000 626.7000 ;
	    RECT 1117.8000 617.4000 1119.0000 618.6000 ;
	    RECT 1122.6000 614.4000 1123.8000 615.6000 ;
	    RECT 1122.7500 606.6000 1123.6500 614.4000 ;
	    RECT 1144.3500 612.6000 1145.2500 755.4000 ;
	    RECT 1151.4000 710.4000 1152.6000 711.6000 ;
	    RECT 1151.5500 684.6000 1152.4501 710.4000 ;
	    RECT 1151.4000 683.4000 1152.6000 684.6000 ;
	    RECT 1161.1500 681.6000 1162.0500 764.4000 ;
	    RECT 1163.5500 738.6000 1164.4501 818.4000 ;
	    RECT 1165.8000 816.3000 1167.0000 833.7000 ;
	    RECT 1168.2001 827.4000 1169.4000 828.6000 ;
	    RECT 1168.3500 822.6000 1169.2500 827.4000 ;
	    RECT 1168.2001 821.4000 1169.4000 822.6000 ;
	    RECT 1170.6000 816.3000 1171.8000 833.7000 ;
	    RECT 1173.0000 816.3000 1174.2001 836.7000 ;
	    RECT 1175.4000 816.3000 1176.6000 836.7000 ;
	    RECT 1177.9501 825.6000 1178.8500 839.4000 ;
	    RECT 1182.7500 828.6000 1183.6500 845.4000 ;
	    RECT 1194.7500 840.6000 1195.6500 884.4000 ;
	    RECT 1197.0000 876.3000 1198.2001 896.7000 ;
	    RECT 1199.4000 876.3000 1200.6000 896.7000 ;
	    RECT 1201.8000 876.3000 1203.0000 893.7000 ;
	    RECT 1204.2001 881.4000 1205.4000 882.6000 ;
	    RECT 1206.6000 876.3000 1207.8000 893.7000 ;
	    RECT 1209.1500 879.6000 1210.0500 905.4000 ;
	    RECT 1209.0000 878.4000 1210.2001 879.6000 ;
	    RECT 1209.1500 876.6000 1210.0500 878.4000 ;
	    RECT 1209.0000 875.4000 1210.2001 876.6000 ;
	    RECT 1211.4000 876.3000 1212.6000 893.7000 ;
	    RECT 1213.8000 876.3000 1215.0000 896.7000 ;
	    RECT 1216.2001 876.3000 1217.4000 896.7000 ;
	    RECT 1218.6000 876.3000 1219.8000 896.7000 ;
	    RECT 1206.6000 860.4000 1207.8000 861.6000 ;
	    RECT 1213.8000 860.4000 1215.0000 861.6000 ;
	    RECT 1218.6000 860.4000 1219.8000 861.6000 ;
	    RECT 1206.7500 846.6000 1207.6500 860.4000 ;
	    RECT 1211.4000 857.4000 1212.6000 858.6000 ;
	    RECT 1206.6000 845.4000 1207.8000 846.6000 ;
	    RECT 1194.6000 839.4000 1195.8000 840.6000 ;
	    RECT 1201.8000 833.4000 1203.0000 834.6000 ;
	    RECT 1182.6000 827.4000 1183.8000 828.6000 ;
	    RECT 1177.8000 824.4000 1179.0000 825.6000 ;
	    RECT 1177.9501 810.6000 1178.8500 824.4000 ;
	    RECT 1177.8000 809.4000 1179.0000 810.6000 ;
	    RECT 1170.6000 803.4000 1171.8000 804.6000 ;
	    RECT 1177.8000 803.4000 1179.0000 804.6000 ;
	    RECT 1170.7500 798.6000 1171.6500 803.4000 ;
	    RECT 1170.6000 797.4000 1171.8000 798.6000 ;
	    RECT 1170.7500 768.6000 1171.6500 797.4000 ;
	    RECT 1170.6000 767.4000 1171.8000 768.6000 ;
	    RECT 1163.4000 737.4000 1164.6000 738.6000 ;
	    RECT 1163.4000 731.4000 1164.6000 732.6000 ;
	    RECT 1161.0000 680.4000 1162.2001 681.6000 ;
	    RECT 1146.6000 623.4000 1147.8000 624.6000 ;
	    RECT 1144.2001 611.4000 1145.4000 612.6000 ;
	    RECT 1122.6000 605.4000 1123.8000 606.6000 ;
	    RECT 1125.0000 596.4000 1126.2001 597.6000 ;
	    RECT 1125.1500 588.6000 1126.0500 596.4000 ;
	    RECT 1125.0000 587.4000 1126.2001 588.6000 ;
	    RECT 1129.8000 584.4000 1131.0000 585.6000 ;
	    RECT 1129.9501 582.6000 1130.8500 584.4000 ;
	    RECT 1129.8000 581.4000 1131.0000 582.6000 ;
	    RECT 1127.4000 575.4000 1128.6000 576.6000 ;
	    RECT 1132.2001 576.3000 1133.4000 596.7000 ;
	    RECT 1134.6000 576.3000 1135.8000 596.7000 ;
	    RECT 1137.0000 576.3000 1138.2001 593.7000 ;
	    RECT 1139.4000 581.4000 1140.6000 582.6000 ;
	    RECT 1127.5500 567.6000 1128.4501 575.4000 ;
	    RECT 1127.4000 566.4000 1128.6000 567.6000 ;
	    RECT 1134.6000 567.4500 1135.8000 567.6000 ;
	    RECT 1139.5500 567.4500 1140.4501 581.4000 ;
	    RECT 1141.8000 576.3000 1143.0000 593.7000 ;
	    RECT 1144.3500 579.6000 1145.2500 611.4000 ;
	    RECT 1146.7500 606.6000 1147.6500 623.4000 ;
	    RECT 1146.6000 605.4000 1147.8000 606.6000 ;
	    RECT 1144.2001 578.4000 1145.4000 579.6000 ;
	    RECT 1146.6000 576.3000 1147.8000 593.7000 ;
	    RECT 1149.0000 576.3000 1150.2001 596.7000 ;
	    RECT 1151.4000 576.3000 1152.6000 596.7000 ;
	    RECT 1153.8000 576.3000 1155.0000 596.7000 ;
	    RECT 1156.2001 587.4000 1157.4000 588.6000 ;
	    RECT 1156.3500 570.6000 1157.2500 587.4000 ;
	    RECT 1156.2001 569.4000 1157.4000 570.6000 ;
	    RECT 1134.6000 566.5500 1140.4501 567.4500 ;
	    RECT 1134.6000 566.4000 1135.8000 566.5500 ;
	    RECT 1141.8000 563.4000 1143.0000 564.6000 ;
	    RECT 1141.9501 558.6000 1142.8500 563.4000 ;
	    RECT 1144.2001 560.4000 1145.4000 561.6000 ;
	    RECT 1144.3500 558.6000 1145.2500 560.4000 ;
	    RECT 1134.6000 557.4000 1135.8000 558.6000 ;
	    RECT 1137.0000 557.4000 1138.2001 558.6000 ;
	    RECT 1141.8000 557.4000 1143.0000 558.6000 ;
	    RECT 1144.2001 557.4000 1145.4000 558.6000 ;
	    RECT 1134.7500 552.6000 1135.6500 557.4000 ;
	    RECT 1134.6000 551.4000 1135.8000 552.6000 ;
	    RECT 1117.8000 539.4000 1119.0000 540.6000 ;
	    RECT 1110.6000 524.4000 1111.8000 525.6000 ;
	    RECT 1108.2001 509.4000 1109.4000 510.6000 ;
	    RECT 1091.4000 500.4000 1092.6000 501.6000 ;
	    RECT 1091.5500 468.6000 1092.4501 500.4000 ;
	    RECT 1110.7500 495.6000 1111.6500 524.4000 ;
	    RECT 1117.9501 522.6000 1118.8500 539.4000 ;
	    RECT 1137.1500 531.4500 1138.0500 557.4000 ;
	    RECT 1141.9501 546.6000 1142.8500 557.4000 ;
	    RECT 1141.8000 545.4000 1143.0000 546.6000 ;
	    RECT 1139.4000 539.4000 1140.6000 540.6000 ;
	    RECT 1134.7500 530.5500 1138.0500 531.4500 ;
	    RECT 1117.8000 521.4000 1119.0000 522.6000 ;
	    RECT 1127.4000 515.4000 1128.6000 516.6000 ;
	    RECT 1117.8000 503.4000 1119.0000 504.6000 ;
	    RECT 1103.4000 494.4000 1104.6000 495.6000 ;
	    RECT 1110.6000 494.4000 1111.8000 495.6000 ;
	    RECT 1098.6000 479.4000 1099.8000 480.6000 ;
	    RECT 1091.4000 467.4000 1092.6000 468.6000 ;
	    RECT 1091.5500 465.6000 1092.4501 467.4000 ;
	    RECT 1091.4000 464.4000 1092.6000 465.6000 ;
	    RECT 1096.2001 464.4000 1097.4000 465.6000 ;
	    RECT 1089.0000 380.4000 1090.2001 381.6000 ;
	    RECT 1091.5500 360.6000 1092.4501 464.4000 ;
	    RECT 1096.3500 432.6000 1097.2500 464.4000 ;
	    RECT 1098.7500 462.6000 1099.6500 479.4000 ;
	    RECT 1101.0000 464.4000 1102.2001 465.6000 ;
	    RECT 1098.6000 461.4000 1099.8000 462.6000 ;
	    RECT 1101.1500 456.6000 1102.0500 464.4000 ;
	    RECT 1103.5500 462.6000 1104.4501 494.4000 ;
	    RECT 1117.9501 489.4500 1118.8500 503.4000 ;
	    RECT 1127.5500 495.6000 1128.4501 515.4000 ;
	    RECT 1134.7500 510.6000 1135.6500 530.5500 ;
	    RECT 1137.0000 527.4000 1138.2001 528.6000 ;
	    RECT 1134.6000 509.4000 1135.8000 510.6000 ;
	    RECT 1132.2001 503.4000 1133.4000 504.6000 ;
	    RECT 1132.3500 498.6000 1133.2500 503.4000 ;
	    RECT 1137.1500 498.6000 1138.0500 527.4000 ;
	    RECT 1139.5500 522.6000 1140.4501 539.4000 ;
	    RECT 1146.6000 527.4000 1147.8000 528.6000 ;
	    RECT 1141.8000 524.4000 1143.0000 525.6000 ;
	    RECT 1141.9501 522.6000 1142.8500 524.4000 ;
	    RECT 1139.4000 521.4000 1140.6000 522.6000 ;
	    RECT 1141.8000 521.4000 1143.0000 522.6000 ;
	    RECT 1132.2001 497.4000 1133.4000 498.6000 ;
	    RECT 1137.0000 497.4000 1138.2001 498.6000 ;
	    RECT 1149.0000 497.4000 1150.2001 498.6000 ;
	    RECT 1127.4000 494.4000 1128.6000 495.6000 ;
	    RECT 1132.3500 492.6000 1133.2500 497.4000 ;
	    RECT 1134.6000 494.4000 1135.8000 495.6000 ;
	    RECT 1132.2001 491.4000 1133.4000 492.6000 ;
	    RECT 1117.9501 488.5500 1121.2500 489.4500 ;
	    RECT 1110.6000 485.4000 1111.8000 486.6000 ;
	    RECT 1103.4000 461.4000 1104.6000 462.6000 ;
	    RECT 1110.7500 456.6000 1111.6500 485.4000 ;
	    RECT 1115.4000 461.4000 1116.6000 462.6000 ;
	    RECT 1101.0000 455.4000 1102.2001 456.6000 ;
	    RECT 1110.6000 455.4000 1111.8000 456.6000 ;
	    RECT 1093.8000 431.4000 1095.0000 432.6000 ;
	    RECT 1096.2001 431.4000 1097.4000 432.6000 ;
	    RECT 1093.9501 384.6000 1094.8500 431.4000 ;
	    RECT 1093.8000 383.4000 1095.0000 384.6000 ;
	    RECT 1093.8000 371.4000 1095.0000 372.6000 ;
	    RECT 1091.4000 359.4000 1092.6000 360.6000 ;
	    RECT 1093.9501 345.6000 1094.8500 371.4000 ;
	    RECT 1098.6000 350.4000 1099.8000 351.6000 ;
	    RECT 1098.7500 345.6000 1099.6500 350.4000 ;
	    RECT 1101.1500 348.6000 1102.0500 455.4000 ;
	    RECT 1115.5500 435.6000 1116.4501 461.4000 ;
	    RECT 1120.3500 441.6000 1121.2500 488.5500 ;
	    RECT 1134.7500 468.4500 1135.6500 494.4000 ;
	    RECT 1132.3500 467.5500 1135.6500 468.4500 ;
	    RECT 1132.3500 462.6000 1133.2500 467.5500 ;
	    RECT 1134.6000 464.4000 1135.8000 465.6000 ;
	    RECT 1134.7500 462.6000 1135.6500 464.4000 ;
	    RECT 1132.2001 461.4000 1133.4000 462.6000 ;
	    RECT 1134.6000 461.4000 1135.8000 462.6000 ;
	    RECT 1122.6000 443.4000 1123.8000 444.6000 ;
	    RECT 1120.2001 440.4000 1121.4000 441.6000 ;
	    RECT 1115.4000 434.4000 1116.6000 435.6000 ;
	    RECT 1105.5000 407.7000 1106.7001 408.9000 ;
	    RECT 1115.4000 407.7000 1116.6000 408.9000 ;
	    RECT 1105.5000 400.5000 1106.4000 407.7000 ;
	    RECT 1109.4000 402.6000 1110.6000 402.9000 ;
	    RECT 1115.7001 402.6000 1116.6000 407.7000 ;
	    RECT 1117.8000 407.4000 1119.0000 408.6000 ;
	    RECT 1117.9501 402.6000 1118.8500 407.4000 ;
	    RECT 1109.4000 401.7000 1116.6000 402.6000 ;
	    RECT 1108.2001 400.5000 1109.4000 400.8000 ;
	    RECT 1113.3000 400.5000 1114.5000 400.8000 ;
	    RECT 1115.7001 400.5000 1116.6000 401.7000 ;
	    RECT 1117.8000 401.4000 1119.0000 402.6000 ;
	    RECT 1105.5000 399.3000 1106.7001 400.5000 ;
	    RECT 1108.2001 399.6000 1114.5000 400.5000 ;
	    RECT 1115.4000 399.3000 1116.6000 400.5000 ;
	    RECT 1120.3500 390.6000 1121.2500 440.4000 ;
	    RECT 1120.2001 389.4000 1121.4000 390.6000 ;
	    RECT 1113.0000 383.4000 1114.2001 384.6000 ;
	    RECT 1117.8000 383.4000 1119.0000 384.6000 ;
	    RECT 1108.2001 377.4000 1109.4000 378.6000 ;
	    RECT 1105.8000 374.4000 1107.0000 375.6000 ;
	    RECT 1105.9501 372.6000 1106.8500 374.4000 ;
	    RECT 1105.8000 371.4000 1107.0000 372.6000 ;
	    RECT 1101.0000 347.4000 1102.2001 348.6000 ;
	    RECT 1093.8000 344.4000 1095.0000 345.6000 ;
	    RECT 1098.6000 344.4000 1099.8000 345.6000 ;
	    RECT 1089.0000 335.4000 1090.2001 336.6000 ;
	    RECT 1089.1500 288.6000 1090.0500 335.4000 ;
	    RECT 1093.9501 327.6000 1094.8500 344.4000 ;
	    RECT 1093.8000 326.4000 1095.0000 327.6000 ;
	    RECT 1101.0000 324.4500 1102.2001 324.6000 ;
	    RECT 1101.0000 323.5500 1104.4501 324.4500 ;
	    RECT 1101.0000 323.4000 1102.2001 323.5500 ;
	    RECT 1101.1500 318.6000 1102.0500 323.4000 ;
	    RECT 1101.0000 317.4000 1102.2001 318.6000 ;
	    RECT 1096.2001 314.4000 1097.4000 315.6000 ;
	    RECT 1089.0000 287.4000 1090.2001 288.6000 ;
	    RECT 1093.8000 287.4000 1095.0000 288.6000 ;
	    RECT 1089.1500 228.6000 1090.0500 287.4000 ;
	    RECT 1093.9501 282.6000 1094.8500 287.4000 ;
	    RECT 1093.8000 281.4000 1095.0000 282.6000 ;
	    RECT 1096.3500 270.6000 1097.2500 314.4000 ;
	    RECT 1101.0000 311.4000 1102.2001 312.6000 ;
	    RECT 1101.1500 291.6000 1102.0500 311.4000 ;
	    RECT 1101.0000 290.4000 1102.2001 291.6000 ;
	    RECT 1098.6000 287.4000 1099.8000 288.6000 ;
	    RECT 1096.2001 269.4000 1097.4000 270.6000 ;
	    RECT 1098.7500 252.6000 1099.6500 287.4000 ;
	    RECT 1103.5500 285.6000 1104.4501 323.5500 ;
	    RECT 1108.3500 294.6000 1109.2500 377.4000 ;
	    RECT 1110.6000 344.4000 1111.8000 345.6000 ;
	    RECT 1108.2001 293.4000 1109.4000 294.6000 ;
	    RECT 1105.8000 287.4000 1107.0000 288.6000 ;
	    RECT 1103.4000 284.4000 1104.6000 285.6000 ;
	    RECT 1105.9501 264.6000 1106.8500 287.4000 ;
	    RECT 1101.0000 263.4000 1102.2001 264.6000 ;
	    RECT 1105.8000 263.4000 1107.0000 264.6000 ;
	    RECT 1093.8000 251.4000 1095.0000 252.6000 ;
	    RECT 1098.6000 251.4000 1099.8000 252.6000 ;
	    RECT 1093.9501 234.6000 1094.8500 251.4000 ;
	    RECT 1093.8000 233.4000 1095.0000 234.6000 ;
	    RECT 1089.0000 227.4000 1090.2001 228.6000 ;
	    RECT 1089.1500 222.6000 1090.0500 227.4000 ;
	    RECT 1101.1500 225.6000 1102.0500 263.4000 ;
	    RECT 1108.3500 258.6000 1109.2500 293.4000 ;
	    RECT 1110.7500 282.6000 1111.6500 344.4000 ;
	    RECT 1113.1500 312.6000 1114.0500 383.4000 ;
	    RECT 1117.9501 375.6000 1118.8500 383.4000 ;
	    RECT 1117.8000 374.4000 1119.0000 375.6000 ;
	    RECT 1120.2001 359.4000 1121.4000 360.6000 ;
	    RECT 1115.4000 347.4000 1116.6000 348.6000 ;
	    RECT 1120.3500 342.6000 1121.2500 359.4000 ;
	    RECT 1120.2001 341.4000 1121.4000 342.6000 ;
	    RECT 1134.7500 336.6000 1135.6500 461.4000 ;
	    RECT 1137.1500 348.6000 1138.0500 497.4000 ;
	    RECT 1141.8000 458.4000 1143.0000 459.6000 ;
	    RECT 1141.9501 444.6000 1142.8500 458.4000 ;
	    RECT 1146.6000 455.4000 1147.8000 456.6000 ;
	    RECT 1139.4000 443.4000 1140.6000 444.6000 ;
	    RECT 1141.8000 443.4000 1143.0000 444.6000 ;
	    RECT 1139.5500 432.6000 1140.4501 443.4000 ;
	    RECT 1144.2001 440.4000 1145.4000 441.6000 ;
	    RECT 1141.8000 437.4000 1143.0000 438.6000 ;
	    RECT 1139.4000 431.4000 1140.6000 432.6000 ;
	    RECT 1141.9501 402.6000 1142.8500 437.4000 ;
	    RECT 1141.8000 401.4000 1143.0000 402.6000 ;
	    RECT 1137.0000 347.4000 1138.2001 348.6000 ;
	    RECT 1134.6000 335.4000 1135.8000 336.6000 ;
	    RECT 1129.8000 329.4000 1131.0000 330.6000 ;
	    RECT 1129.9501 315.6000 1130.8500 329.4000 ;
	    RECT 1129.8000 314.4000 1131.0000 315.6000 ;
	    RECT 1132.2001 314.4000 1133.4000 315.6000 ;
	    RECT 1113.0000 311.4000 1114.2001 312.6000 ;
	    RECT 1110.6000 281.4000 1111.8000 282.6000 ;
	    RECT 1110.7500 261.6000 1111.6500 281.4000 ;
	    RECT 1110.6000 260.4000 1111.8000 261.6000 ;
	    RECT 1103.4000 257.4000 1104.6000 258.6000 ;
	    RECT 1108.2001 257.4000 1109.4000 258.6000 ;
	    RECT 1103.5500 255.4500 1104.4501 257.4000 ;
	    RECT 1110.6000 255.4500 1111.8000 255.6000 ;
	    RECT 1103.5500 254.5500 1111.8000 255.4500 ;
	    RECT 1110.6000 254.4000 1111.8000 254.5500 ;
	    RECT 1113.1500 228.6000 1114.0500 311.4000 ;
	    RECT 1132.3500 306.6000 1133.2500 314.4000 ;
	    RECT 1132.2001 305.4000 1133.4000 306.6000 ;
	    RECT 1120.2001 287.4000 1121.4000 288.6000 ;
	    RECT 1132.2001 287.4000 1133.4000 288.6000 ;
	    RECT 1115.4000 281.4000 1116.6000 282.6000 ;
	    RECT 1115.5500 270.6000 1116.4501 281.4000 ;
	    RECT 1120.3500 279.6000 1121.2500 287.4000 ;
	    RECT 1120.2001 278.4000 1121.4000 279.6000 ;
	    RECT 1115.4000 269.4000 1116.6000 270.6000 ;
	    RECT 1120.3500 264.6000 1121.2500 278.4000 ;
	    RECT 1132.3500 276.4500 1133.2500 287.4000 ;
	    RECT 1134.6000 276.4500 1135.8000 276.6000 ;
	    RECT 1132.3500 275.5500 1135.8000 276.4500 ;
	    RECT 1134.6000 275.4000 1135.8000 275.5500 ;
	    RECT 1120.2001 263.4000 1121.4000 264.6000 ;
	    RECT 1120.3500 261.6000 1121.2500 263.4000 ;
	    RECT 1120.2001 260.4000 1121.4000 261.6000 ;
	    RECT 1134.6000 239.4000 1135.8000 240.6000 ;
	    RECT 1134.7500 234.6000 1135.6500 239.4000 ;
	    RECT 1134.6000 233.4000 1135.8000 234.6000 ;
	    RECT 1113.0000 227.4000 1114.2001 228.6000 ;
	    RECT 1101.0000 224.4000 1102.2001 225.6000 ;
	    RECT 1137.0000 224.4000 1138.2001 225.6000 ;
	    RECT 1084.2001 221.5500 1087.6500 222.4500 ;
	    RECT 1084.2001 221.4000 1085.4000 221.5500 ;
	    RECT 1089.0000 221.4000 1090.2001 222.6000 ;
	    RECT 1134.6000 221.4000 1135.8000 222.6000 ;
	    RECT 1089.1500 144.6000 1090.0500 221.4000 ;
	    RECT 1101.0000 215.4000 1102.2001 216.6000 ;
	    RECT 1093.8000 194.4000 1095.0000 195.6000 ;
	    RECT 1089.0000 143.4000 1090.2001 144.6000 ;
	    RECT 1079.4000 134.4000 1080.6000 135.6000 ;
	    RECT 1081.8000 134.4000 1083.0000 135.6000 ;
	    RECT 1093.9501 126.6000 1094.8500 194.4000 ;
	    RECT 1098.6000 179.4000 1099.8000 180.6000 ;
	    RECT 1096.2001 167.4000 1097.4000 168.6000 ;
	    RECT 1098.7500 165.6000 1099.6500 179.4000 ;
	    RECT 1101.1500 171.6000 1102.0500 215.4000 ;
	    RECT 1134.7500 204.6000 1135.6500 221.4000 ;
	    RECT 1108.2001 203.4000 1109.4000 204.6000 ;
	    RECT 1134.6000 203.4000 1135.8000 204.6000 ;
	    RECT 1108.3500 198.6000 1109.2500 203.4000 ;
	    RECT 1108.2001 197.4000 1109.4000 198.6000 ;
	    RECT 1105.8000 194.4000 1107.0000 195.6000 ;
	    RECT 1134.6000 194.4000 1135.8000 195.6000 ;
	    RECT 1105.9501 192.6000 1106.8500 194.4000 ;
	    RECT 1105.8000 191.4000 1107.0000 192.6000 ;
	    RECT 1110.6000 191.4000 1111.8000 192.6000 ;
	    RECT 1113.0000 185.4000 1114.2001 186.6000 ;
	    RECT 1110.6000 173.4000 1111.8000 174.6000 ;
	    RECT 1101.0000 170.4000 1102.2001 171.6000 ;
	    RECT 1103.4000 167.4000 1104.6000 168.6000 ;
	    RECT 1108.2001 167.4000 1109.4000 168.6000 ;
	    RECT 1098.6000 164.4000 1099.8000 165.6000 ;
	    RECT 1103.5500 144.6000 1104.4501 167.4000 ;
	    RECT 1105.8000 155.4000 1107.0000 156.6000 ;
	    RECT 1103.4000 143.4000 1104.6000 144.6000 ;
	    RECT 1103.4000 140.4000 1104.6000 141.6000 ;
	    RECT 1103.5500 138.6000 1104.4501 140.4000 ;
	    RECT 1098.6000 137.4000 1099.8000 138.6000 ;
	    RECT 1103.4000 137.4000 1104.6000 138.6000 ;
	    RECT 1093.8000 125.4000 1095.0000 126.6000 ;
	    RECT 1081.8000 119.4000 1083.0000 120.6000 ;
	    RECT 1074.6000 101.4000 1075.8000 102.6000 ;
	    RECT 1053.0000 95.4000 1054.2001 96.6000 ;
	    RECT 1055.4000 53.4000 1056.6000 54.6000 ;
	    RECT 1055.5500 42.6000 1056.4501 53.4000 ;
	    RECT 1058.1000 47.7000 1059.3000 48.9000 ;
	    RECT 1067.4000 47.7000 1068.6000 48.9000 ;
	    RECT 1050.6000 41.4000 1051.8000 42.6000 ;
	    RECT 1055.4000 41.4000 1056.6000 42.6000 ;
	    RECT 1058.1000 40.5000 1059.0000 47.7000 ;
	    RECT 1059.9000 44.7000 1061.1000 45.9000 ;
	    RECT 1060.2001 42.6000 1061.1000 44.7000 ;
	    RECT 1067.7001 42.6000 1068.6000 47.7000 ;
	    RECT 1069.9501 45.4500 1070.8500 98.4000 ;
	    RECT 1069.9501 44.5500 1073.2500 45.4500 ;
	    RECT 1060.2001 41.7000 1068.6000 42.6000 ;
	    RECT 1060.2001 40.5000 1061.4000 40.8000 ;
	    RECT 1065.3000 40.5000 1066.5000 40.8000 ;
	    RECT 1067.7001 40.5000 1068.6000 41.7000 ;
	    RECT 1069.8000 41.4000 1071.0000 42.6000 ;
	    RECT 1058.1000 39.6000 1066.5000 40.5000 ;
	    RECT 1058.1000 39.3000 1059.3000 39.6000 ;
	    RECT 1067.4000 39.3000 1068.6000 40.5000 ;
	    RECT 1048.2001 29.4000 1049.4000 30.6000 ;
	    RECT 1033.8000 17.4000 1035.0000 18.6000 ;
	    RECT 829.8000 14.4000 831.0000 15.6000 ;
	    RECT 892.2000 14.4000 893.4000 15.6000 ;
	    RECT 1026.6000 14.4000 1027.8000 15.6000 ;
	    RECT 777.0000 11.4000 778.2000 12.6000 ;
	    RECT 796.2000 11.4000 797.4000 12.6000 ;
	    RECT 829.9500 6.6000 830.8500 14.4000 ;
	    RECT 1026.7500 6.6000 1027.6500 14.4000 ;
	    RECT 829.8000 5.4000 831.0000 6.6000 ;
	    RECT 1026.6000 6.4500 1027.8000 6.6000 ;
	    RECT 1029.0000 6.4500 1030.2001 6.6000 ;
	    RECT 1026.6000 5.5500 1030.2001 6.4500 ;
	    RECT 1036.2001 6.3000 1037.4000 26.7000 ;
	    RECT 1038.6000 6.3000 1039.8000 26.7000 ;
	    RECT 1041.0000 9.3000 1042.2001 26.7000 ;
	    RECT 1043.4000 23.4000 1044.6000 24.6000 ;
	    RECT 1043.5500 21.6000 1044.4501 23.4000 ;
	    RECT 1043.4000 20.4000 1044.6000 21.6000 ;
	    RECT 1045.8000 9.3000 1047.0000 26.7000 ;
	    RECT 1048.3500 24.6000 1049.2500 29.4000 ;
	    RECT 1048.2001 23.4000 1049.4000 24.6000 ;
	    RECT 1050.6000 9.3000 1051.8000 26.7000 ;
	    RECT 1053.0000 6.3000 1054.2001 26.7000 ;
	    RECT 1055.4000 6.3000 1056.6000 26.7000 ;
	    RECT 1057.8000 6.3000 1059.0000 26.7000 ;
	    RECT 1072.3500 12.6000 1073.2500 44.5500 ;
	    RECT 1074.7500 30.6000 1075.6500 101.4000 ;
	    RECT 1077.0000 96.3000 1078.2001 113.7000 ;
	    RECT 1081.9501 105.6000 1082.8500 119.4000 ;
	    RECT 1081.8000 104.4000 1083.0000 105.6000 ;
	    RECT 1091.4000 96.3000 1092.6000 113.7000 ;
	    RECT 1089.0000 71.4000 1090.2001 72.6000 ;
	    RECT 1086.6000 47.4000 1087.8000 48.6000 ;
	    RECT 1086.7500 45.6000 1087.6500 47.4000 ;
	    RECT 1089.1500 45.6000 1090.0500 71.4000 ;
	    RECT 1098.7500 66.6000 1099.6500 137.4000 ;
	    RECT 1110.7500 105.6000 1111.6500 173.4000 ;
	    RECT 1113.1500 162.6000 1114.0500 185.4000 ;
	    RECT 1120.2001 179.4000 1121.4000 180.6000 ;
	    RECT 1120.3500 171.6000 1121.2500 179.4000 ;
	    RECT 1120.2001 170.4000 1121.4000 171.6000 ;
	    RECT 1134.7500 168.6000 1135.6500 194.4000 ;
	    RECT 1134.6000 167.4000 1135.8000 168.6000 ;
	    RECT 1113.0000 161.4000 1114.2001 162.6000 ;
	    RECT 1132.2001 155.4000 1133.4000 156.6000 ;
	    RECT 1137.1500 120.6000 1138.0500 224.4000 ;
	    RECT 1141.8000 203.4000 1143.0000 204.6000 ;
	    RECT 1141.9501 192.6000 1142.8500 203.4000 ;
	    RECT 1141.8000 191.4000 1143.0000 192.6000 ;
	    RECT 1141.9501 171.6000 1142.8500 191.4000 ;
	    RECT 1139.4000 170.4000 1140.6000 171.6000 ;
	    RECT 1141.8000 170.4000 1143.0000 171.6000 ;
	    RECT 1139.5500 165.6000 1140.4501 170.4000 ;
	    RECT 1139.4000 164.4000 1140.6000 165.6000 ;
	    RECT 1141.8000 161.4000 1143.0000 162.6000 ;
	    RECT 1137.0000 119.4000 1138.2001 120.6000 ;
	    RECT 1139.4000 107.4000 1140.6000 108.6000 ;
	    RECT 1110.6000 104.4000 1111.8000 105.6000 ;
	    RECT 1113.0000 98.4000 1114.2001 99.6000 ;
	    RECT 1113.1500 72.6000 1114.0500 98.4000 ;
	    RECT 1113.0000 71.4000 1114.2001 72.6000 ;
	    RECT 1098.6000 65.4000 1099.8000 66.6000 ;
	    RECT 1139.5500 60.6000 1140.4501 107.4000 ;
	    RECT 1139.4000 59.4000 1140.6000 60.6000 ;
	    RECT 1086.6000 44.4000 1087.8000 45.6000 ;
	    RECT 1089.0000 44.4000 1090.2001 45.6000 ;
	    RECT 1141.9501 42.6000 1142.8500 161.4000 ;
	    RECT 1144.3500 132.6000 1145.2500 440.4000 ;
	    RECT 1146.7500 435.6000 1147.6500 455.4000 ;
	    RECT 1146.6000 434.4000 1147.8000 435.6000 ;
	    RECT 1149.1500 408.6000 1150.0500 497.4000 ;
	    RECT 1153.8000 467.4000 1155.0000 468.6000 ;
	    RECT 1153.9501 465.6000 1154.8500 467.4000 ;
	    RECT 1153.8000 464.4000 1155.0000 465.6000 ;
	    RECT 1153.8000 458.4000 1155.0000 459.6000 ;
	    RECT 1151.4000 425.4000 1152.6000 426.6000 ;
	    RECT 1151.5500 414.6000 1152.4501 425.4000 ;
	    RECT 1151.4000 413.4000 1152.6000 414.6000 ;
	    RECT 1149.0000 407.4000 1150.2001 408.6000 ;
	    RECT 1146.6000 404.4000 1147.8000 405.6000 ;
	    RECT 1149.0000 404.4000 1150.2001 405.6000 ;
	    RECT 1146.7500 402.6000 1147.6500 404.4000 ;
	    RECT 1146.6000 401.4000 1147.8000 402.6000 ;
	    RECT 1149.1500 375.6000 1150.0500 404.4000 ;
	    RECT 1153.9501 396.6000 1154.8500 458.4000 ;
	    RECT 1156.3500 432.6000 1157.2500 569.4000 ;
	    RECT 1161.0000 503.4000 1162.2001 504.6000 ;
	    RECT 1161.1500 501.6000 1162.0500 503.4000 ;
	    RECT 1161.0000 500.4000 1162.2001 501.6000 ;
	    RECT 1161.0000 494.4000 1162.2001 495.6000 ;
	    RECT 1161.1500 471.6000 1162.0500 494.4000 ;
	    RECT 1161.0000 470.4000 1162.2001 471.6000 ;
	    RECT 1163.5500 441.6000 1164.4501 731.4000 ;
	    RECT 1177.9501 681.6000 1178.8500 803.4000 ;
	    RECT 1180.2001 761.4000 1181.4000 762.6000 ;
	    RECT 1199.4000 761.4000 1200.6000 762.6000 ;
	    RECT 1180.3500 714.6000 1181.2500 761.4000 ;
	    RECT 1199.5500 750.6000 1200.4501 761.4000 ;
	    RECT 1201.9501 759.6000 1202.8500 833.4000 ;
	    RECT 1211.5500 828.6000 1212.4501 857.4000 ;
	    RECT 1213.9501 846.6000 1214.8500 860.4000 ;
	    RECT 1213.8000 845.4000 1215.0000 846.6000 ;
	    RECT 1211.4000 827.4000 1212.6000 828.6000 ;
	    RECT 1218.7500 822.6000 1219.6500 860.4000 ;
	    RECT 1211.4000 821.4000 1212.6000 822.6000 ;
	    RECT 1218.6000 821.4000 1219.8000 822.6000 ;
	    RECT 1211.5500 804.6000 1212.4501 821.4000 ;
	    RECT 1211.4000 803.4000 1212.6000 804.6000 ;
	    RECT 1206.6000 797.4000 1207.8000 798.6000 ;
	    RECT 1201.8000 758.4000 1203.0000 759.6000 ;
	    RECT 1199.4000 749.4000 1200.6000 750.6000 ;
	    RECT 1192.2001 737.4000 1193.4000 738.6000 ;
	    RECT 1180.2001 713.4000 1181.4000 714.6000 ;
	    RECT 1182.6000 696.3000 1183.8000 716.7000 ;
	    RECT 1185.0000 696.3000 1186.2001 716.7000 ;
	    RECT 1187.4000 696.3000 1188.6000 716.7000 ;
	    RECT 1189.8000 696.3000 1191.0000 713.7000 ;
	    RECT 1192.3500 699.6000 1193.2500 737.4000 ;
	    RECT 1201.9501 732.6000 1202.8500 758.4000 ;
	    RECT 1201.8000 731.4000 1203.0000 732.6000 ;
	    RECT 1192.2001 698.4000 1193.4000 699.6000 ;
	    RECT 1192.3500 687.6000 1193.2500 698.4000 ;
	    RECT 1194.6000 696.3000 1195.8000 713.7000 ;
	    RECT 1197.0000 713.4000 1198.2001 714.6000 ;
	    RECT 1197.1500 702.6000 1198.0500 713.4000 ;
	    RECT 1197.0000 701.4000 1198.2001 702.6000 ;
	    RECT 1199.4000 696.3000 1200.6000 713.7000 ;
	    RECT 1201.8000 696.3000 1203.0000 716.7000 ;
	    RECT 1204.2001 696.3000 1205.4000 716.7000 ;
	    RECT 1206.7500 708.6000 1207.6500 797.4000 ;
	    RECT 1211.4000 761.4000 1212.6000 762.6000 ;
	    RECT 1211.5500 750.6000 1212.4501 761.4000 ;
	    RECT 1211.4000 749.4000 1212.6000 750.6000 ;
	    RECT 1211.5500 720.6000 1212.4501 749.4000 ;
	    RECT 1211.4000 719.4000 1212.6000 720.6000 ;
	    RECT 1211.5500 708.6000 1212.4501 719.4000 ;
	    RECT 1206.6000 707.4000 1207.8000 708.6000 ;
	    RECT 1211.4000 707.4000 1212.6000 708.6000 ;
	    RECT 1206.7500 705.6000 1207.6500 707.4000 ;
	    RECT 1206.6000 704.4000 1207.8000 705.6000 ;
	    RECT 1221.1500 690.6000 1222.0500 989.4000 ;
	    RECT 1235.5500 981.6000 1236.4501 1010.5500 ;
	    RECT 1237.9501 1008.6000 1238.8500 1010.5500 ;
	    RECT 1237.8000 1007.4000 1239.0000 1008.6000 ;
	    RECT 1245.1500 1005.6000 1246.0500 1037.4000 ;
	    RECT 1245.0000 1004.4000 1246.2001 1005.6000 ;
	    RECT 1235.4000 980.4000 1236.6000 981.6000 ;
	    RECT 1235.4000 977.4000 1236.6000 978.6000 ;
	    RECT 1228.2001 965.4000 1229.4000 966.6000 ;
	    RECT 1225.8000 929.4000 1227.0000 930.6000 ;
	    RECT 1223.4000 887.4000 1224.6000 888.6000 ;
	    RECT 1223.5500 882.6000 1224.4501 887.4000 ;
	    RECT 1223.4000 881.4000 1224.6000 882.6000 ;
	    RECT 1225.9501 870.6000 1226.8500 929.4000 ;
	    RECT 1225.8000 869.4000 1227.0000 870.6000 ;
	    RECT 1223.4000 863.4000 1224.6000 864.6000 ;
	    RECT 1223.5500 858.6000 1224.4501 863.4000 ;
	    RECT 1223.4000 857.4000 1224.6000 858.6000 ;
	    RECT 1223.5500 855.6000 1224.4501 857.4000 ;
	    RECT 1223.4000 854.4000 1224.6000 855.6000 ;
	    RECT 1199.4000 689.4000 1200.6000 690.6000 ;
	    RECT 1221.0000 689.4000 1222.2001 690.6000 ;
	    RECT 1192.2001 686.4000 1193.4000 687.6000 ;
	    RECT 1197.0000 686.4000 1198.2001 687.6000 ;
	    RECT 1177.8000 680.4000 1179.0000 681.6000 ;
	    RECT 1180.2001 680.4000 1181.4000 681.6000 ;
	    RECT 1175.4000 677.4000 1176.6000 678.6000 ;
	    RECT 1177.8000 677.4000 1179.0000 678.6000 ;
	    RECT 1165.8000 674.4000 1167.0000 675.6000 ;
	    RECT 1165.9501 558.6000 1166.8500 674.4000 ;
	    RECT 1175.5500 648.6000 1176.4501 677.4000 ;
	    RECT 1175.4000 647.4000 1176.6000 648.6000 ;
	    RECT 1177.9501 642.6000 1178.8500 677.4000 ;
	    RECT 1177.8000 641.4000 1179.0000 642.6000 ;
	    RECT 1173.0000 620.4000 1174.2001 621.6000 ;
	    RECT 1173.1500 615.4500 1174.0500 620.4000 ;
	    RECT 1177.8000 617.4000 1179.0000 618.6000 ;
	    RECT 1175.4000 615.4500 1176.6000 615.6000 ;
	    RECT 1173.1500 614.5500 1176.6000 615.4500 ;
	    RECT 1175.4000 614.4000 1176.6000 614.5500 ;
	    RECT 1175.5500 612.6000 1176.4501 614.4000 ;
	    RECT 1175.4000 611.4000 1176.6000 612.6000 ;
	    RECT 1177.8000 611.4000 1179.0000 612.6000 ;
	    RECT 1170.6000 599.4000 1171.8000 600.6000 ;
	    RECT 1168.2001 590.4000 1169.4000 591.6000 ;
	    RECT 1168.3500 588.6000 1169.2500 590.4000 ;
	    RECT 1168.2001 587.4000 1169.4000 588.6000 ;
	    RECT 1170.7500 582.6000 1171.6500 599.4000 ;
	    RECT 1168.2001 581.4000 1169.4000 582.6000 ;
	    RECT 1170.6000 581.4000 1171.8000 582.6000 ;
	    RECT 1165.8000 557.4000 1167.0000 558.6000 ;
	    RECT 1168.3500 555.6000 1169.2500 581.4000 ;
	    RECT 1177.9501 570.6000 1178.8500 611.4000 ;
	    RECT 1180.3500 582.6000 1181.2500 680.4000 ;
	    RECT 1197.1500 645.6000 1198.0500 686.4000 ;
	    RECT 1197.0000 644.4000 1198.2001 645.6000 ;
	    RECT 1189.8000 641.4000 1191.0000 642.6000 ;
	    RECT 1182.6000 584.4000 1183.8000 585.6000 ;
	    RECT 1180.2001 581.4000 1181.4000 582.6000 ;
	    RECT 1177.8000 569.4000 1179.0000 570.6000 ;
	    RECT 1170.6000 557.4000 1171.8000 558.6000 ;
	    RECT 1177.9501 555.6000 1178.8500 569.4000 ;
	    RECT 1168.2001 554.4000 1169.4000 555.6000 ;
	    RECT 1177.8000 554.4000 1179.0000 555.6000 ;
	    RECT 1168.3500 552.6000 1169.2500 554.4000 ;
	    RECT 1168.2001 551.4000 1169.4000 552.6000 ;
	    RECT 1173.0000 551.4000 1174.2001 552.6000 ;
	    RECT 1173.1500 534.6000 1174.0500 551.4000 ;
	    RECT 1175.4000 545.4000 1176.6000 546.6000 ;
	    RECT 1173.0000 533.4000 1174.2001 534.6000 ;
	    RECT 1170.6000 527.4000 1171.8000 528.6000 ;
	    RECT 1170.7500 522.6000 1171.6500 527.4000 ;
	    RECT 1165.8000 521.4000 1167.0000 522.6000 ;
	    RECT 1170.6000 521.4000 1171.8000 522.6000 ;
	    RECT 1165.9501 495.6000 1166.8500 521.4000 ;
	    RECT 1165.8000 494.4000 1167.0000 495.6000 ;
	    RECT 1165.8000 467.4000 1167.0000 468.6000 ;
	    RECT 1163.4000 440.4000 1164.6000 441.6000 ;
	    RECT 1165.9501 438.6000 1166.8500 467.4000 ;
	    RECT 1168.2001 449.4000 1169.4000 450.6000 ;
	    RECT 1168.3500 444.6000 1169.2500 449.4000 ;
	    RECT 1168.2001 443.4000 1169.4000 444.6000 ;
	    RECT 1175.5500 441.6000 1176.4501 545.4000 ;
	    RECT 1182.7500 498.6000 1183.6500 584.4000 ;
	    RECT 1189.9501 582.6000 1190.8500 641.4000 ;
	    RECT 1199.5500 588.6000 1200.4501 689.4000 ;
	    RECT 1221.0000 683.4000 1222.2001 684.6000 ;
	    RECT 1204.2001 677.4000 1205.4000 678.6000 ;
	    RECT 1204.3500 615.6000 1205.2500 677.4000 ;
	    RECT 1221.1500 648.6000 1222.0500 683.4000 ;
	    RECT 1225.9501 678.6000 1226.8500 869.4000 ;
	    RECT 1228.3500 858.6000 1229.2500 965.4000 ;
	    RECT 1235.5500 888.6000 1236.4501 977.4000 ;
	    RECT 1240.2001 944.4000 1241.4000 945.6000 ;
	    RECT 1235.4000 887.4000 1236.6000 888.6000 ;
	    RECT 1237.8000 887.4000 1239.0000 888.6000 ;
	    RECT 1237.9501 882.6000 1238.8500 887.4000 ;
	    RECT 1237.8000 881.4000 1239.0000 882.6000 ;
	    RECT 1228.2001 857.4000 1229.4000 858.6000 ;
	    RECT 1235.4000 818.4000 1236.6000 819.6000 ;
	    RECT 1235.5500 816.6000 1236.4501 818.4000 ;
	    RECT 1235.4000 815.4000 1236.6000 816.6000 ;
	    RECT 1240.3500 768.6000 1241.2500 944.4000 ;
	    RECT 1242.6000 890.4000 1243.8000 891.6000 ;
	    RECT 1242.7500 864.6000 1243.6500 890.4000 ;
	    RECT 1242.6000 863.4000 1243.8000 864.6000 ;
	    RECT 1242.7500 858.6000 1243.6500 863.4000 ;
	    RECT 1242.6000 857.4000 1243.8000 858.6000 ;
	    RECT 1247.4000 854.4000 1248.6000 855.6000 ;
	    RECT 1247.5500 840.6000 1248.4501 854.4000 ;
	    RECT 1247.4000 839.4000 1248.6000 840.6000 ;
	    RECT 1245.0000 785.4000 1246.2001 786.6000 ;
	    RECT 1240.2001 767.4000 1241.4000 768.6000 ;
	    RECT 1235.4000 726.3000 1236.6000 746.7000 ;
	    RECT 1237.8000 726.3000 1239.0000 746.7000 ;
	    RECT 1240.2001 726.3000 1241.4000 746.7000 ;
	    RECT 1242.6000 729.3000 1243.8000 746.7000 ;
	    RECT 1245.1500 744.6000 1246.0500 785.4000 ;
	    RECT 1249.8000 761.4000 1251.0000 762.6000 ;
	    RECT 1245.0000 743.4000 1246.2001 744.6000 ;
	    RECT 1245.1500 738.6000 1246.0500 743.4000 ;
	    RECT 1245.0000 737.4000 1246.2001 738.6000 ;
	    RECT 1247.4000 729.3000 1248.6000 746.7000 ;
	    RECT 1249.9501 741.6000 1250.8500 761.4000 ;
	    RECT 1257.1500 750.4500 1258.0500 1187.4000 ;
	    RECT 1281.0000 1176.3000 1282.2001 1196.7001 ;
	    RECT 1283.4000 1176.3000 1284.6000 1196.7001 ;
	    RECT 1285.8000 1176.3000 1287.0000 1196.7001 ;
	    RECT 1288.2001 1176.3000 1289.4000 1193.7001 ;
	    RECT 1290.6000 1178.4000 1291.8000 1179.6000 ;
	    RECT 1290.7500 1176.6000 1291.6500 1178.4000 ;
	    RECT 1290.6000 1175.4000 1291.8000 1176.6000 ;
	    RECT 1293.0000 1176.3000 1294.2001 1193.7001 ;
	    RECT 1295.4000 1181.4000 1296.6000 1182.6000 ;
	    RECT 1295.5500 1170.6000 1296.4501 1181.4000 ;
	    RECT 1297.8000 1176.3000 1299.0000 1193.7001 ;
	    RECT 1300.2001 1176.3000 1301.4000 1196.7001 ;
	    RECT 1302.6000 1176.3000 1303.8000 1196.7001 ;
	    RECT 1309.9501 1188.6000 1310.8500 1199.4000 ;
	    RECT 1305.0000 1187.4000 1306.2001 1188.6000 ;
	    RECT 1309.8000 1187.4000 1311.0000 1188.6000 ;
	    RECT 1305.1500 1185.6000 1306.0500 1187.4000 ;
	    RECT 1305.0000 1184.4000 1306.2001 1185.6000 ;
	    RECT 1288.2001 1169.4000 1289.4000 1170.6000 ;
	    RECT 1295.4000 1169.4000 1296.6000 1170.6000 ;
	    RECT 1288.3500 1152.6000 1289.2500 1169.4000 ;
	    RECT 1305.1500 1158.6000 1306.0500 1184.4000 ;
	    RECT 1314.7500 1176.6000 1315.6500 1238.4000 ;
	    RECT 1317.0000 1236.3000 1318.2001 1253.7001 ;
	    RECT 1319.4000 1241.4000 1320.6000 1242.6000 ;
	    RECT 1321.8000 1236.3000 1323.0000 1253.7001 ;
	    RECT 1324.2001 1236.3000 1325.4000 1256.7001 ;
	    RECT 1326.6000 1236.3000 1327.8000 1256.7001 ;
	    RECT 1329.1500 1254.6000 1330.0500 1367.4000 ;
	    RECT 1341.1500 1350.6000 1342.0500 1397.4000 ;
	    RECT 1345.9501 1395.6000 1346.8500 1397.4000 ;
	    RECT 1345.8000 1394.4000 1347.0000 1395.6000 ;
	    RECT 1345.8000 1370.4000 1347.0000 1371.6000 ;
	    RECT 1343.4000 1355.4000 1344.6000 1356.6000 ;
	    RECT 1341.0000 1349.4000 1342.2001 1350.6000 ;
	    RECT 1343.5500 1341.6000 1344.4501 1355.4000 ;
	    RECT 1336.2001 1340.4000 1337.4000 1341.6000 ;
	    RECT 1343.4000 1340.4000 1344.6000 1341.6000 ;
	    RECT 1336.3500 1320.6000 1337.2500 1340.4000 ;
	    RECT 1345.9501 1338.6000 1346.8500 1370.4000 ;
	    RECT 1348.3500 1362.6000 1349.2500 1400.4000 ;
	    RECT 1374.7500 1398.6000 1375.6500 1460.4000 ;
	    RECT 1377.0000 1400.4000 1378.2001 1401.6000 ;
	    RECT 1374.6000 1397.4000 1375.8000 1398.6000 ;
	    RECT 1377.1500 1380.6000 1378.0500 1400.4000 ;
	    RECT 1384.2001 1394.4000 1385.4000 1395.6000 ;
	    RECT 1377.0000 1379.4000 1378.2001 1380.6000 ;
	    RECT 1348.2001 1361.4000 1349.4000 1362.6000 ;
	    RECT 1348.2001 1343.4000 1349.4000 1344.6000 ;
	    RECT 1348.3500 1338.6000 1349.2500 1343.4000 ;
	    RECT 1377.1500 1341.6000 1378.0500 1379.4000 ;
	    RECT 1377.0000 1340.4000 1378.2001 1341.6000 ;
	    RECT 1345.8000 1337.4000 1347.0000 1338.6000 ;
	    RECT 1348.2001 1337.4000 1349.4000 1338.6000 ;
	    RECT 1350.6000 1337.4000 1351.8000 1338.6000 ;
	    RECT 1345.9501 1335.6000 1346.8500 1337.4000 ;
	    RECT 1345.8000 1334.4000 1347.0000 1335.6000 ;
	    RECT 1336.2001 1319.4000 1337.4000 1320.6000 ;
	    RECT 1350.7500 1308.6000 1351.6500 1337.4000 ;
	    RECT 1377.1500 1335.6000 1378.0500 1340.4000 ;
	    RECT 1384.3500 1338.6000 1385.2500 1394.4000 ;
	    RECT 1398.6000 1343.4000 1399.8000 1344.6000 ;
	    RECT 1398.7500 1338.6000 1399.6500 1343.4000 ;
	    RECT 1446.7500 1341.6000 1447.6500 1463.4000 ;
	    RECT 1477.8000 1457.4000 1479.0000 1458.6000 ;
	    RECT 1473.0000 1454.4000 1474.2001 1455.6000 ;
	    RECT 1473.1500 1446.6000 1474.0500 1454.4000 ;
	    RECT 1473.0000 1445.4000 1474.2001 1446.6000 ;
	    RECT 1477.9501 1443.4501 1478.8500 1457.4000 ;
	    RECT 1480.2001 1446.3000 1481.4000 1466.7001 ;
	    RECT 1482.6000 1446.3000 1483.8000 1466.7001 ;
	    RECT 1485.0000 1449.3000 1486.2001 1466.7001 ;
	    RECT 1487.4000 1463.4000 1488.6000 1464.6000 ;
	    RECT 1487.5500 1461.6000 1488.4501 1463.4000 ;
	    RECT 1487.4000 1460.4000 1488.6000 1461.6000 ;
	    RECT 1489.8000 1449.3000 1491.0000 1466.7001 ;
	    RECT 1492.2001 1463.4000 1493.4000 1464.6000 ;
	    RECT 1477.9501 1442.5500 1481.2500 1443.4501 ;
	    RECT 1470.6000 1416.3000 1471.8000 1436.7001 ;
	    RECT 1473.0000 1416.3000 1474.2001 1436.7001 ;
	    RECT 1475.4000 1416.3000 1476.6000 1436.7001 ;
	    RECT 1480.3500 1434.6000 1481.2500 1442.5500 ;
	    RECT 1492.3500 1440.6000 1493.2500 1463.4000 ;
	    RECT 1494.6000 1449.3000 1495.8000 1466.7001 ;
	    RECT 1497.0000 1446.3000 1498.2001 1466.7001 ;
	    RECT 1499.4000 1446.3000 1500.6000 1466.7001 ;
	    RECT 1501.8000 1446.3000 1503.0000 1466.7001 ;
	    RECT 1566.6000 1460.4000 1567.8000 1461.6000 ;
	    RECT 1523.4000 1457.4000 1524.6000 1458.6000 ;
	    RECT 1564.2001 1457.4000 1565.4000 1458.6000 ;
	    RECT 1523.5500 1452.6000 1524.4501 1457.4000 ;
	    RECT 1557.0000 1454.4000 1558.2001 1455.6000 ;
	    RECT 1523.4000 1451.4000 1524.6000 1452.6000 ;
	    RECT 1492.2001 1439.4000 1493.4000 1440.6000 ;
	    RECT 1497.0000 1439.4000 1498.2001 1440.6000 ;
	    RECT 1477.8000 1416.3000 1479.0000 1433.7001 ;
	    RECT 1480.2001 1433.4000 1481.4000 1434.6000 ;
	    RECT 1480.2001 1418.4000 1481.4000 1419.6000 ;
	    RECT 1480.3500 1404.6000 1481.2500 1418.4000 ;
	    RECT 1482.6000 1416.3000 1483.8000 1433.7001 ;
	    RECT 1485.0000 1421.4000 1486.2001 1422.6000 ;
	    RECT 1480.2001 1403.4000 1481.4000 1404.6000 ;
	    RECT 1485.1500 1401.6000 1486.0500 1421.4000 ;
	    RECT 1487.4000 1416.3000 1488.6000 1433.7001 ;
	    RECT 1489.8000 1416.3000 1491.0000 1436.7001 ;
	    RECT 1492.2001 1416.3000 1493.4000 1436.7001 ;
	    RECT 1494.6000 1433.4000 1495.8000 1434.6000 ;
	    RECT 1494.7500 1425.6000 1495.6500 1433.4000 ;
	    RECT 1494.6000 1424.4000 1495.8000 1425.6000 ;
	    RECT 1485.0000 1400.4000 1486.2001 1401.6000 ;
	    RECT 1451.4000 1385.4000 1452.6000 1386.6000 ;
	    RECT 1408.2001 1340.4000 1409.4000 1341.6000 ;
	    RECT 1417.8000 1340.4000 1419.0000 1341.6000 ;
	    RECT 1446.6000 1340.4000 1447.8000 1341.6000 ;
	    RECT 1384.2001 1337.4000 1385.4000 1338.6000 ;
	    RECT 1398.6000 1337.4000 1399.8000 1338.6000 ;
	    RECT 1377.0000 1334.4000 1378.2001 1335.6000 ;
	    RECT 1350.6000 1307.4000 1351.8000 1308.6000 ;
	    RECT 1379.4000 1301.4000 1380.6000 1302.6000 ;
	    RECT 1333.8000 1259.4000 1335.0000 1260.6000 ;
	    RECT 1329.0000 1253.4000 1330.2001 1254.6000 ;
	    RECT 1329.1500 1245.6000 1330.0500 1253.4000 ;
	    RECT 1333.9501 1248.6000 1334.8500 1259.4000 ;
	    RECT 1333.8000 1247.4000 1335.0000 1248.6000 ;
	    RECT 1367.4000 1247.4000 1368.6000 1248.6000 ;
	    RECT 1329.0000 1244.4000 1330.2001 1245.6000 ;
	    RECT 1319.4000 1217.4000 1320.6000 1218.6000 ;
	    RECT 1319.5500 1212.6000 1320.4501 1217.4000 ;
	    RECT 1319.4000 1211.4000 1320.6000 1212.6000 ;
	    RECT 1317.0000 1199.4000 1318.2001 1200.6000 ;
	    RECT 1317.1500 1182.6000 1318.0500 1199.4000 ;
	    RECT 1317.0000 1181.4000 1318.2001 1182.6000 ;
	    RECT 1314.6000 1175.4000 1315.8000 1176.6000 ;
	    RECT 1305.0000 1157.4000 1306.2001 1158.6000 ;
	    RECT 1288.2001 1151.4000 1289.4000 1152.6000 ;
	    RECT 1269.0000 1130.4000 1270.2001 1131.6000 ;
	    RECT 1269.1500 1119.6000 1270.0500 1130.4000 ;
	    RECT 1309.8000 1127.4000 1311.0000 1128.6000 ;
	    RECT 1285.8000 1124.4000 1287.0000 1125.6000 ;
	    RECT 1314.6000 1124.4000 1315.8000 1125.6000 ;
	    RECT 1285.9501 1122.6000 1286.8500 1124.4000 ;
	    RECT 1314.7500 1122.6000 1315.6500 1124.4000 ;
	    RECT 1317.1500 1122.6000 1318.0500 1181.4000 ;
	    RECT 1285.8000 1121.4000 1287.0000 1122.6000 ;
	    RECT 1307.4000 1121.4000 1308.6000 1122.6000 ;
	    RECT 1314.6000 1121.4000 1315.8000 1122.6000 ;
	    RECT 1317.0000 1121.4000 1318.2001 1122.6000 ;
	    RECT 1319.4000 1121.4000 1320.6000 1122.6000 ;
	    RECT 1269.0000 1118.4000 1270.2001 1119.6000 ;
	    RECT 1269.1500 1080.6000 1270.0500 1118.4000 ;
	    RECT 1319.5500 1110.6000 1320.4501 1121.4000 ;
	    RECT 1297.8000 1109.4000 1299.0000 1110.6000 ;
	    RECT 1319.4000 1109.4000 1320.6000 1110.6000 ;
	    RECT 1288.2001 1097.4000 1289.4000 1098.6000 ;
	    RECT 1283.4000 1094.4000 1284.6000 1095.6000 ;
	    RECT 1283.5500 1086.6000 1284.4501 1094.4000 ;
	    RECT 1283.4000 1085.4000 1284.6000 1086.6000 ;
	    RECT 1290.6000 1086.3000 1291.8000 1106.7001 ;
	    RECT 1293.0000 1086.3000 1294.2001 1106.7001 ;
	    RECT 1295.4000 1089.3000 1296.6000 1106.7001 ;
	    RECT 1297.9501 1101.6000 1298.8500 1109.4000 ;
	    RECT 1297.8000 1100.4000 1299.0000 1101.6000 ;
	    RECT 1300.2001 1089.3000 1301.4000 1106.7001 ;
	    RECT 1302.6000 1103.4000 1303.8000 1104.6000 ;
	    RECT 1305.0000 1089.3000 1306.2001 1106.7001 ;
	    RECT 1307.4000 1086.3000 1308.6000 1106.7001 ;
	    RECT 1309.8000 1086.3000 1311.0000 1106.7001 ;
	    RECT 1312.2001 1086.3000 1313.4000 1106.7001 ;
	    RECT 1326.6000 1103.4000 1327.8000 1104.6000 ;
	    RECT 1326.7500 1092.6000 1327.6500 1103.4000 ;
	    RECT 1326.6000 1091.4000 1327.8000 1092.6000 ;
	    RECT 1269.0000 1079.4000 1270.2001 1080.6000 ;
	    RECT 1281.0000 1079.4000 1282.2001 1080.6000 ;
	    RECT 1266.6000 1064.4000 1267.8000 1065.6000 ;
	    RECT 1266.7500 1056.6000 1267.6500 1064.4000 ;
	    RECT 1266.6000 1055.4000 1267.8000 1056.6000 ;
	    RECT 1259.4000 1043.4000 1260.6000 1044.6000 ;
	    RECT 1266.7500 1041.6000 1267.6500 1055.4000 ;
	    RECT 1266.6000 1040.4000 1267.8000 1041.6000 ;
	    RECT 1261.8000 1001.4000 1263.0000 1002.6000 ;
	    RECT 1261.8000 983.4000 1263.0000 984.6000 ;
	    RECT 1261.9501 948.6000 1262.8500 983.4000 ;
	    RECT 1264.2001 980.4000 1265.4000 981.6000 ;
	    RECT 1264.3500 960.6000 1265.2500 980.4000 ;
	    RECT 1271.4000 974.4000 1272.6000 975.6000 ;
	    RECT 1271.5500 966.6000 1272.4501 974.4000 ;
	    RECT 1271.4000 965.4000 1272.6000 966.6000 ;
	    RECT 1264.2001 959.4000 1265.4000 960.6000 ;
	    RECT 1261.8000 947.4000 1263.0000 948.6000 ;
	    RECT 1261.9501 912.6000 1262.8500 947.4000 ;
	    RECT 1261.8000 911.4000 1263.0000 912.6000 ;
	    RECT 1266.6000 884.4000 1267.8000 885.6000 ;
	    RECT 1266.7500 861.6000 1267.6500 884.4000 ;
	    RECT 1266.6000 860.4000 1267.8000 861.6000 ;
	    RECT 1266.6000 833.4000 1267.8000 834.6000 ;
	    RECT 1257.1500 749.5500 1260.4501 750.4500 ;
	    RECT 1249.8000 740.4000 1251.0000 741.6000 ;
	    RECT 1252.2001 729.3000 1253.4000 746.7000 ;
	    RECT 1242.6000 725.4000 1243.8000 726.6000 ;
	    RECT 1254.6000 726.3000 1255.8000 746.7000 ;
	    RECT 1257.0000 726.3000 1258.2001 746.7000 ;
	    RECT 1259.5500 738.6000 1260.4501 749.5500 ;
	    RECT 1259.4000 737.4000 1260.6000 738.6000 ;
	    RECT 1264.2001 734.4000 1265.4000 735.6000 ;
	    RECT 1264.3500 726.6000 1265.2500 734.4000 ;
	    RECT 1264.2001 725.4000 1265.4000 726.6000 ;
	    RECT 1242.7500 708.6000 1243.6500 725.4000 ;
	    RECT 1245.0000 710.4000 1246.2001 711.6000 ;
	    RECT 1242.6000 707.4000 1243.8000 708.6000 ;
	    RECT 1225.8000 677.4000 1227.0000 678.6000 ;
	    RECT 1245.1500 660.6000 1246.0500 710.4000 ;
	    RECT 1247.4000 704.4000 1248.6000 705.6000 ;
	    RECT 1247.5500 678.6000 1248.4501 704.4000 ;
	    RECT 1266.7500 678.6000 1267.6500 833.4000 ;
	    RECT 1273.8000 737.4000 1275.0000 738.6000 ;
	    RECT 1273.9501 705.6000 1274.8500 737.4000 ;
	    RECT 1276.2001 734.4000 1277.4000 735.6000 ;
	    RECT 1273.8000 704.4000 1275.0000 705.6000 ;
	    RECT 1269.0000 698.4000 1270.2001 699.6000 ;
	    RECT 1269.1500 690.6000 1270.0500 698.4000 ;
	    RECT 1269.0000 689.4000 1270.2001 690.6000 ;
	    RECT 1247.4000 677.4000 1248.6000 678.6000 ;
	    RECT 1266.6000 677.4000 1267.8000 678.6000 ;
	    RECT 1247.5500 672.6000 1248.4501 677.4000 ;
	    RECT 1266.6000 674.4000 1267.8000 675.6000 ;
	    RECT 1247.4000 671.4000 1248.6000 672.6000 ;
	    RECT 1266.7500 660.6000 1267.6500 674.4000 ;
	    RECT 1245.0000 659.4000 1246.2001 660.6000 ;
	    RECT 1266.6000 659.4000 1267.8000 660.6000 ;
	    RECT 1221.0000 647.4000 1222.2001 648.6000 ;
	    RECT 1228.2001 647.4000 1229.4000 648.6000 ;
	    RECT 1216.2001 644.4000 1217.4000 645.6000 ;
	    RECT 1213.8000 641.4000 1215.0000 642.6000 ;
	    RECT 1213.9501 624.6000 1214.8500 641.4000 ;
	    RECT 1213.8000 623.4000 1215.0000 624.6000 ;
	    RECT 1209.0000 620.4000 1210.2001 621.6000 ;
	    RECT 1213.8000 620.4000 1215.0000 621.6000 ;
	    RECT 1206.6000 617.4000 1207.8000 618.6000 ;
	    RECT 1204.2001 614.4000 1205.4000 615.6000 ;
	    RECT 1209.1500 612.6000 1210.0500 620.4000 ;
	    RECT 1213.9501 618.6000 1214.8500 620.4000 ;
	    RECT 1213.8000 617.4000 1215.0000 618.6000 ;
	    RECT 1209.0000 611.4000 1210.2001 612.6000 ;
	    RECT 1201.8000 593.4000 1203.0000 594.6000 ;
	    RECT 1199.4000 587.4000 1200.6000 588.6000 ;
	    RECT 1189.8000 581.4000 1191.0000 582.6000 ;
	    RECT 1201.9501 555.6000 1202.8500 593.4000 ;
	    RECT 1204.2001 587.4000 1205.4000 588.6000 ;
	    RECT 1201.8000 554.4000 1203.0000 555.6000 ;
	    RECT 1204.3500 546.6000 1205.2500 587.4000 ;
	    RECT 1216.3500 585.6000 1217.2500 644.4000 ;
	    RECT 1221.1500 639.6000 1222.0500 647.4000 ;
	    RECT 1221.0000 638.4000 1222.2001 639.6000 ;
	    RECT 1223.4000 629.4000 1224.6000 630.6000 ;
	    RECT 1223.5500 618.6000 1224.4501 629.4000 ;
	    RECT 1228.3500 624.6000 1229.2500 647.4000 ;
	    RECT 1245.1500 642.6000 1246.0500 659.4000 ;
	    RECT 1269.1500 645.6000 1270.0500 689.4000 ;
	    RECT 1273.9501 684.6000 1274.8500 704.4000 ;
	    RECT 1273.8000 683.4000 1275.0000 684.6000 ;
	    RECT 1273.8000 680.4000 1275.0000 681.6000 ;
	    RECT 1273.9501 672.6000 1274.8500 680.4000 ;
	    RECT 1276.3500 678.6000 1277.2500 734.4000 ;
	    RECT 1281.1500 732.6000 1282.0500 1079.4000 ;
	    RECT 1317.0000 1067.4000 1318.2001 1068.6000 ;
	    RECT 1314.6000 1061.4000 1315.8000 1062.6000 ;
	    RECT 1283.4000 1058.4000 1284.6000 1059.6000 ;
	    RECT 1283.5500 1041.4501 1284.4501 1058.4000 ;
	    RECT 1293.0000 1043.4000 1294.2001 1044.6000 ;
	    RECT 1307.4000 1043.4000 1308.6000 1044.6000 ;
	    RECT 1285.8000 1041.4501 1287.0000 1041.6000 ;
	    RECT 1283.5500 1040.5500 1287.0000 1041.4501 ;
	    RECT 1285.8000 1040.4000 1287.0000 1040.5500 ;
	    RECT 1285.9501 978.6000 1286.8500 1040.4000 ;
	    RECT 1288.2001 1037.4000 1289.4000 1038.6000 ;
	    RECT 1293.1500 1035.6000 1294.0500 1043.4000 ;
	    RECT 1295.4000 1040.4000 1296.6000 1041.6000 ;
	    RECT 1297.8000 1040.4000 1299.0000 1041.6000 ;
	    RECT 1293.0000 1034.4000 1294.2001 1035.6000 ;
	    RECT 1295.5500 1032.6000 1296.4501 1040.4000 ;
	    RECT 1297.9501 1038.6000 1298.8500 1040.4000 ;
	    RECT 1297.8000 1037.4000 1299.0000 1038.6000 ;
	    RECT 1297.8000 1034.4000 1299.0000 1035.6000 ;
	    RECT 1295.4000 1031.4000 1296.6000 1032.6000 ;
	    RECT 1290.6000 1013.4000 1291.8000 1014.6000 ;
	    RECT 1288.2001 1010.4000 1289.4000 1011.6000 ;
	    RECT 1288.3500 1008.6000 1289.2500 1010.4000 ;
	    RECT 1290.7500 1008.6000 1291.6500 1013.4000 ;
	    RECT 1297.9501 1008.6000 1298.8500 1034.4000 ;
	    RECT 1307.5500 1026.6000 1308.4501 1043.4000 ;
	    RECT 1314.7500 1026.6000 1315.6500 1061.4000 ;
	    RECT 1307.4000 1025.4000 1308.6000 1026.6000 ;
	    RECT 1314.6000 1025.4000 1315.8000 1026.6000 ;
	    RECT 1317.1500 1008.6000 1318.0500 1067.4000 ;
	    RECT 1319.4000 1058.4000 1320.6000 1059.6000 ;
	    RECT 1319.5500 1056.6000 1320.4501 1058.4000 ;
	    RECT 1319.4000 1055.4000 1320.6000 1056.6000 ;
	    RECT 1288.2001 1007.4000 1289.4000 1008.6000 ;
	    RECT 1290.6000 1007.4000 1291.8000 1008.6000 ;
	    RECT 1297.8000 1007.4000 1299.0000 1008.6000 ;
	    RECT 1317.0000 1007.4000 1318.2001 1008.6000 ;
	    RECT 1288.3500 978.6000 1289.2500 1007.4000 ;
	    RECT 1290.7500 984.4500 1291.6500 1007.4000 ;
	    RECT 1293.0000 1004.4000 1294.2001 1005.6000 ;
	    RECT 1326.6000 1004.4000 1327.8000 1005.6000 ;
	    RECT 1293.1500 1002.6000 1294.0500 1004.4000 ;
	    RECT 1293.0000 1001.4000 1294.2001 1002.6000 ;
	    RECT 1300.2001 1001.4000 1301.4000 1002.6000 ;
	    RECT 1321.8000 1001.4000 1323.0000 1002.6000 ;
	    RECT 1293.0000 984.4500 1294.2001 984.6000 ;
	    RECT 1290.7500 983.5500 1294.2001 984.4500 ;
	    RECT 1293.0000 983.4000 1294.2001 983.5500 ;
	    RECT 1285.8000 977.4000 1287.0000 978.6000 ;
	    RECT 1288.2001 977.4000 1289.4000 978.6000 ;
	    RECT 1288.3500 741.6000 1289.2500 977.4000 ;
	    RECT 1290.6000 899.4000 1291.8000 900.6000 ;
	    RECT 1290.7500 882.6000 1291.6500 899.4000 ;
	    RECT 1290.6000 881.4000 1291.8000 882.6000 ;
	    RECT 1288.2001 740.4000 1289.4000 741.6000 ;
	    RECT 1281.0000 731.4000 1282.2001 732.6000 ;
	    RECT 1276.2001 677.4000 1277.4000 678.6000 ;
	    RECT 1278.6000 677.4000 1279.8000 678.6000 ;
	    RECT 1273.8000 671.4000 1275.0000 672.6000 ;
	    RECT 1276.2001 647.4000 1277.4000 648.6000 ;
	    RECT 1249.8000 644.4000 1251.0000 645.6000 ;
	    RECT 1269.0000 644.4000 1270.2001 645.6000 ;
	    RECT 1237.8000 641.4000 1239.0000 642.6000 ;
	    RECT 1245.0000 641.4000 1246.2001 642.6000 ;
	    RECT 1237.9501 636.6000 1238.8500 641.4000 ;
	    RECT 1249.9501 636.6000 1250.8500 644.4000 ;
	    RECT 1276.3500 642.6000 1277.2500 647.4000 ;
	    RECT 1252.2001 641.4000 1253.4000 642.6000 ;
	    RECT 1271.4000 641.4000 1272.6000 642.6000 ;
	    RECT 1276.2001 641.4000 1277.4000 642.6000 ;
	    RECT 1237.8000 635.4000 1239.0000 636.6000 ;
	    RECT 1249.8000 635.4000 1251.0000 636.6000 ;
	    RECT 1228.2001 623.4000 1229.4000 624.6000 ;
	    RECT 1230.6000 623.4000 1231.8000 624.6000 ;
	    RECT 1228.3500 618.6000 1229.2500 623.4000 ;
	    RECT 1223.4000 617.4000 1224.6000 618.6000 ;
	    RECT 1228.2001 617.4000 1229.4000 618.6000 ;
	    RECT 1216.2001 584.4000 1217.4000 585.6000 ;
	    RECT 1218.6000 581.4000 1219.8000 582.6000 ;
	    RECT 1211.4000 560.4000 1212.6000 561.6000 ;
	    RECT 1206.6000 558.4500 1207.8000 558.6000 ;
	    RECT 1209.0000 558.4500 1210.2001 558.6000 ;
	    RECT 1206.6000 557.5500 1210.2001 558.4500 ;
	    RECT 1206.6000 557.4000 1207.8000 557.5500 ;
	    RECT 1209.0000 557.4000 1210.2001 557.5500 ;
	    RECT 1211.5500 555.6000 1212.4501 560.4000 ;
	    RECT 1206.6000 554.4000 1207.8000 555.6000 ;
	    RECT 1211.4000 554.4000 1212.6000 555.6000 ;
	    RECT 1204.2001 545.4000 1205.4000 546.6000 ;
	    RECT 1199.4000 533.4000 1200.6000 534.6000 ;
	    RECT 1199.5500 525.6000 1200.4501 533.4000 ;
	    RECT 1192.2001 524.4000 1193.4000 525.6000 ;
	    RECT 1199.4000 524.4000 1200.6000 525.6000 ;
	    RECT 1204.2001 524.4000 1205.4000 525.6000 ;
	    RECT 1189.8000 503.4000 1191.0000 504.6000 ;
	    RECT 1182.6000 497.4000 1183.8000 498.6000 ;
	    RECT 1187.4000 497.4000 1188.6000 498.6000 ;
	    RECT 1185.0000 491.4000 1186.2001 492.6000 ;
	    RECT 1182.6000 485.4000 1183.8000 486.6000 ;
	    RECT 1182.7500 471.6000 1183.6500 485.4000 ;
	    RECT 1185.1500 471.6000 1186.0500 491.4000 ;
	    RECT 1187.5500 480.6000 1188.4501 497.4000 ;
	    RECT 1189.9501 495.6000 1190.8500 503.4000 ;
	    RECT 1189.8000 494.4000 1191.0000 495.6000 ;
	    RECT 1192.3500 492.6000 1193.2500 524.4000 ;
	    RECT 1204.3500 504.6000 1205.2500 524.4000 ;
	    RECT 1206.7500 522.6000 1207.6500 554.4000 ;
	    RECT 1213.8000 551.4000 1215.0000 552.6000 ;
	    RECT 1213.9501 534.6000 1214.8500 551.4000 ;
	    RECT 1218.7500 540.6000 1219.6500 581.4000 ;
	    RECT 1228.2001 569.4000 1229.4000 570.6000 ;
	    RECT 1228.3500 564.6000 1229.2500 569.4000 ;
	    RECT 1228.2001 563.4000 1229.4000 564.6000 ;
	    RECT 1218.6000 539.4000 1219.8000 540.6000 ;
	    RECT 1213.8000 533.4000 1215.0000 534.6000 ;
	    RECT 1209.0000 524.4000 1210.2001 525.6000 ;
	    RECT 1206.6000 521.4000 1207.8000 522.6000 ;
	    RECT 1199.4000 503.4000 1200.6000 504.6000 ;
	    RECT 1204.2001 503.4000 1205.4000 504.6000 ;
	    RECT 1194.6000 497.4000 1195.8000 498.6000 ;
	    RECT 1192.2001 491.4000 1193.4000 492.6000 ;
	    RECT 1194.7500 486.6000 1195.6500 497.4000 ;
	    RECT 1199.5500 495.6000 1200.4501 503.4000 ;
	    RECT 1199.4000 494.4000 1200.6000 495.6000 ;
	    RECT 1194.6000 485.4000 1195.8000 486.6000 ;
	    RECT 1187.4000 479.4000 1188.6000 480.6000 ;
	    RECT 1204.2001 479.4000 1205.4000 480.6000 ;
	    RECT 1197.0000 473.4000 1198.2001 474.6000 ;
	    RECT 1182.6000 470.4000 1183.8000 471.6000 ;
	    RECT 1185.0000 470.4000 1186.2001 471.6000 ;
	    RECT 1180.2001 467.4000 1181.4000 468.6000 ;
	    RECT 1177.8000 461.4000 1179.0000 462.6000 ;
	    RECT 1175.4000 440.4000 1176.6000 441.6000 ;
	    RECT 1163.4000 437.4000 1164.6000 438.6000 ;
	    RECT 1165.8000 437.4000 1167.0000 438.6000 ;
	    RECT 1163.5500 435.6000 1164.4501 437.4000 ;
	    RECT 1163.4000 434.4000 1164.6000 435.6000 ;
	    RECT 1156.2001 431.4000 1157.4000 432.6000 ;
	    RECT 1163.4000 425.4000 1164.6000 426.6000 ;
	    RECT 1156.2001 419.4000 1157.4000 420.6000 ;
	    RECT 1156.3500 402.6000 1157.2500 419.4000 ;
	    RECT 1163.5500 405.6000 1164.4501 425.4000 ;
	    RECT 1163.4000 404.4000 1164.6000 405.6000 ;
	    RECT 1165.9501 402.6000 1166.8500 437.4000 ;
	    RECT 1173.0000 431.4000 1174.2001 432.6000 ;
	    RECT 1170.6000 413.4000 1171.8000 414.6000 ;
	    RECT 1156.2001 401.4000 1157.4000 402.6000 ;
	    RECT 1161.0000 401.4000 1162.2001 402.6000 ;
	    RECT 1165.8000 401.4000 1167.0000 402.6000 ;
	    RECT 1153.8000 395.4000 1155.0000 396.6000 ;
	    RECT 1151.4000 383.4000 1152.6000 384.6000 ;
	    RECT 1158.6000 383.4000 1159.8000 384.6000 ;
	    RECT 1151.5500 381.6000 1152.4501 383.4000 ;
	    RECT 1151.4000 380.4000 1152.6000 381.6000 ;
	    RECT 1153.8000 380.4000 1155.0000 381.6000 ;
	    RECT 1149.0000 374.4000 1150.2001 375.6000 ;
	    RECT 1146.6000 371.4000 1147.8000 372.6000 ;
	    RECT 1146.7500 222.6000 1147.6500 371.4000 ;
	    RECT 1149.1500 345.6000 1150.0500 374.4000 ;
	    RECT 1151.4000 359.4000 1152.6000 360.6000 ;
	    RECT 1149.0000 344.4000 1150.2001 345.6000 ;
	    RECT 1151.5500 342.6000 1152.4501 359.4000 ;
	    RECT 1153.9501 351.4500 1154.8500 380.4000 ;
	    RECT 1158.7500 378.6000 1159.6500 383.4000 ;
	    RECT 1158.6000 377.4000 1159.8000 378.6000 ;
	    RECT 1153.9501 350.5500 1157.2500 351.4500 ;
	    RECT 1153.8000 347.4000 1155.0000 348.6000 ;
	    RECT 1153.9501 345.6000 1154.8500 347.4000 ;
	    RECT 1153.8000 344.4000 1155.0000 345.6000 ;
	    RECT 1151.4000 341.4000 1152.6000 342.6000 ;
	    RECT 1149.0000 317.4000 1150.2001 318.6000 ;
	    RECT 1149.1500 291.6000 1150.0500 317.4000 ;
	    RECT 1149.0000 290.4000 1150.2001 291.6000 ;
	    RECT 1149.1500 282.6000 1150.0500 290.4000 ;
	    RECT 1156.3500 288.6000 1157.2500 350.5500 ;
	    RECT 1158.6000 344.4000 1159.8000 345.6000 ;
	    RECT 1158.7500 324.6000 1159.6500 344.4000 ;
	    RECT 1158.6000 323.4000 1159.8000 324.6000 ;
	    RECT 1158.7500 321.6000 1159.6500 323.4000 ;
	    RECT 1158.6000 320.4000 1159.8000 321.6000 ;
	    RECT 1161.1500 318.6000 1162.0500 401.4000 ;
	    RECT 1165.8000 383.4000 1167.0000 384.6000 ;
	    RECT 1165.9501 360.6000 1166.8500 383.4000 ;
	    RECT 1170.7500 381.6000 1171.6500 413.4000 ;
	    RECT 1170.6000 380.4000 1171.8000 381.6000 ;
	    RECT 1165.8000 359.4000 1167.0000 360.6000 ;
	    RECT 1168.2001 329.4000 1169.4000 330.6000 ;
	    RECT 1168.3500 318.6000 1169.2500 329.4000 ;
	    RECT 1161.0000 317.4000 1162.2001 318.6000 ;
	    RECT 1168.2001 317.4000 1169.4000 318.6000 ;
	    RECT 1170.6000 317.4000 1171.8000 318.6000 ;
	    RECT 1163.4000 314.4000 1164.6000 315.6000 ;
	    RECT 1163.5500 297.6000 1164.4501 314.4000 ;
	    RECT 1168.3500 312.6000 1169.2500 317.4000 ;
	    RECT 1170.7500 315.6000 1171.6500 317.4000 ;
	    RECT 1170.6000 314.4000 1171.8000 315.6000 ;
	    RECT 1165.8000 311.4000 1167.0000 312.6000 ;
	    RECT 1168.2001 311.4000 1169.4000 312.6000 ;
	    RECT 1163.4000 296.4000 1164.6000 297.6000 ;
	    RECT 1165.9501 291.6000 1166.8500 311.4000 ;
	    RECT 1170.7500 306.6000 1171.6500 314.4000 ;
	    RECT 1170.6000 305.4000 1171.8000 306.6000 ;
	    RECT 1165.8000 290.4000 1167.0000 291.6000 ;
	    RECT 1165.9501 288.6000 1166.8500 290.4000 ;
	    RECT 1156.2001 287.4000 1157.4000 288.6000 ;
	    RECT 1165.8000 287.4000 1167.0000 288.6000 ;
	    RECT 1153.8000 285.4500 1155.0000 285.6000 ;
	    RECT 1156.3500 285.4500 1157.2500 287.4000 ;
	    RECT 1153.8000 284.5500 1157.2500 285.4500 ;
	    RECT 1153.8000 284.4000 1155.0000 284.5500 ;
	    RECT 1149.0000 281.4000 1150.2001 282.6000 ;
	    RECT 1149.1500 255.6000 1150.0500 281.4000 ;
	    RECT 1158.6000 275.4000 1159.8000 276.6000 ;
	    RECT 1158.7500 264.6000 1159.6500 275.4000 ;
	    RECT 1158.6000 263.4000 1159.8000 264.6000 ;
	    RECT 1151.4000 260.4000 1152.6000 261.6000 ;
	    RECT 1149.0000 254.4000 1150.2001 255.6000 ;
	    RECT 1146.6000 221.4000 1147.8000 222.6000 ;
	    RECT 1146.7500 186.6000 1147.6500 221.4000 ;
	    RECT 1151.5500 216.6000 1152.4501 260.4000 ;
	    RECT 1158.6000 257.4000 1159.8000 258.6000 ;
	    RECT 1156.2001 224.4000 1157.4000 225.6000 ;
	    RECT 1156.3500 222.6000 1157.2500 224.4000 ;
	    RECT 1156.2001 221.4000 1157.4000 222.6000 ;
	    RECT 1151.4000 215.4000 1152.6000 216.6000 ;
	    RECT 1153.8000 197.4000 1155.0000 198.6000 ;
	    RECT 1153.9501 192.6000 1154.8500 197.4000 ;
	    RECT 1156.3500 195.6000 1157.2500 221.4000 ;
	    RECT 1158.7500 204.6000 1159.6500 257.4000 ;
	    RECT 1170.6000 239.4000 1171.8000 240.6000 ;
	    RECT 1170.7500 234.6000 1171.6500 239.4000 ;
	    RECT 1170.6000 233.4000 1171.8000 234.6000 ;
	    RECT 1173.1500 228.6000 1174.0500 431.4000 ;
	    RECT 1175.5500 372.6000 1176.4501 440.4000 ;
	    RECT 1175.4000 371.4000 1176.6000 372.6000 ;
	    RECT 1175.4000 338.4000 1176.6000 339.6000 ;
	    RECT 1175.5500 336.6000 1176.4501 338.4000 ;
	    RECT 1175.4000 335.4000 1176.6000 336.6000 ;
	    RECT 1177.9501 330.6000 1178.8500 461.4000 ;
	    RECT 1180.3500 456.6000 1181.2500 467.4000 ;
	    RECT 1182.7500 465.6000 1183.6500 470.4000 ;
	    RECT 1197.1500 468.6000 1198.0500 473.4000 ;
	    RECT 1197.0000 467.4000 1198.2001 468.6000 ;
	    RECT 1199.4000 467.4000 1200.6000 468.6000 ;
	    RECT 1182.6000 464.4000 1183.8000 465.6000 ;
	    RECT 1180.2001 455.4000 1181.4000 456.6000 ;
	    RECT 1201.8000 455.4000 1203.0000 456.6000 ;
	    RECT 1201.9501 444.6000 1202.8500 455.4000 ;
	    RECT 1189.8000 443.4000 1191.0000 444.6000 ;
	    RECT 1201.8000 443.4000 1203.0000 444.6000 ;
	    RECT 1189.9501 438.6000 1190.8500 443.4000 ;
	    RECT 1192.2001 440.4000 1193.4000 441.6000 ;
	    RECT 1189.8000 437.4000 1191.0000 438.6000 ;
	    RECT 1192.3500 414.6000 1193.2500 440.4000 ;
	    RECT 1201.9501 438.6000 1202.8500 443.4000 ;
	    RECT 1194.6000 437.4000 1195.8000 438.6000 ;
	    RECT 1201.8000 437.4000 1203.0000 438.6000 ;
	    RECT 1192.2001 413.4000 1193.4000 414.6000 ;
	    RECT 1192.2001 404.4000 1193.4000 405.6000 ;
	    RECT 1185.0000 401.4000 1186.2001 402.6000 ;
	    RECT 1189.8000 401.4000 1191.0000 402.6000 ;
	    RECT 1180.2001 395.4000 1181.4000 396.6000 ;
	    RECT 1180.3500 384.6000 1181.2500 395.4000 ;
	    RECT 1185.1500 390.6000 1186.0500 401.4000 ;
	    RECT 1189.9501 396.6000 1190.8500 401.4000 ;
	    RECT 1189.8000 395.4000 1191.0000 396.6000 ;
	    RECT 1185.0000 389.4000 1186.2001 390.6000 ;
	    RECT 1180.2001 383.4000 1181.4000 384.6000 ;
	    RECT 1189.9501 381.6000 1190.8500 395.4000 ;
	    RECT 1192.3500 384.6000 1193.2500 404.4000 ;
	    RECT 1192.2001 383.4000 1193.4000 384.6000 ;
	    RECT 1189.8000 380.4000 1191.0000 381.6000 ;
	    RECT 1194.7500 342.6000 1195.6500 437.4000 ;
	    RECT 1197.0000 419.4000 1198.2001 420.6000 ;
	    RECT 1197.1500 408.6000 1198.0500 419.4000 ;
	    RECT 1201.8000 413.4000 1203.0000 414.6000 ;
	    RECT 1197.0000 407.4000 1198.2001 408.6000 ;
	    RECT 1201.9501 402.6000 1202.8500 413.4000 ;
	    RECT 1201.8000 401.4000 1203.0000 402.6000 ;
	    RECT 1204.3500 345.6000 1205.2500 479.4000 ;
	    RECT 1206.6000 467.4000 1207.8000 468.6000 ;
	    RECT 1206.7500 408.6000 1207.6500 467.4000 ;
	    RECT 1206.6000 407.4000 1207.8000 408.6000 ;
	    RECT 1209.1500 405.6000 1210.0500 524.4000 ;
	    RECT 1211.4000 509.4000 1212.6000 510.6000 ;
	    RECT 1211.5500 462.6000 1212.4501 509.4000 ;
	    RECT 1211.4000 461.4000 1212.6000 462.6000 ;
	    RECT 1211.5500 435.6000 1212.4501 461.4000 ;
	    RECT 1213.9501 441.6000 1214.8500 533.4000 ;
	    RECT 1213.8000 440.4000 1215.0000 441.6000 ;
	    RECT 1211.4000 434.4000 1212.6000 435.6000 ;
	    RECT 1216.2001 407.4000 1217.4000 408.6000 ;
	    RECT 1209.0000 404.4000 1210.2001 405.6000 ;
	    RECT 1216.3500 345.6000 1217.2500 407.4000 ;
	    RECT 1218.7500 399.6000 1219.6500 539.4000 ;
	    RECT 1228.2001 524.4000 1229.4000 525.6000 ;
	    RECT 1228.3500 522.6000 1229.2500 524.4000 ;
	    RECT 1228.2001 521.4000 1229.4000 522.6000 ;
	    RECT 1221.0000 509.4000 1222.2001 510.6000 ;
	    RECT 1221.1500 495.6000 1222.0500 509.4000 ;
	    RECT 1225.8000 503.4000 1227.0000 504.6000 ;
	    RECT 1223.4000 497.4000 1224.6000 498.6000 ;
	    RECT 1221.0000 494.4000 1222.2001 495.6000 ;
	    RECT 1225.9501 492.6000 1226.8500 503.4000 ;
	    RECT 1221.0000 491.4000 1222.2001 492.6000 ;
	    RECT 1225.8000 491.4000 1227.0000 492.6000 ;
	    RECT 1221.1500 456.6000 1222.0500 491.4000 ;
	    RECT 1221.0000 455.4000 1222.2001 456.6000 ;
	    RECT 1221.1500 441.6000 1222.0500 455.4000 ;
	    RECT 1221.0000 440.4000 1222.2001 441.6000 ;
	    RECT 1218.6000 398.4000 1219.8000 399.6000 ;
	    RECT 1204.2001 344.4000 1205.4000 345.6000 ;
	    RECT 1211.4000 344.4000 1212.6000 345.6000 ;
	    RECT 1216.2001 344.4000 1217.4000 345.6000 ;
	    RECT 1182.6000 341.4000 1183.8000 342.6000 ;
	    RECT 1194.6000 341.4000 1195.8000 342.6000 ;
	    RECT 1209.0000 341.4000 1210.2001 342.6000 ;
	    RECT 1177.8000 329.4000 1179.0000 330.6000 ;
	    RECT 1180.2001 299.4000 1181.4000 300.6000 ;
	    RECT 1180.3500 297.6000 1181.2500 299.4000 ;
	    RECT 1180.2001 296.4000 1181.4000 297.6000 ;
	    RECT 1175.4000 287.4000 1176.6000 288.6000 ;
	    RECT 1175.5500 261.4500 1176.4501 287.4000 ;
	    RECT 1180.2001 275.4000 1181.4000 276.6000 ;
	    RECT 1180.3500 270.6000 1181.2500 275.4000 ;
	    RECT 1180.2001 269.4000 1181.4000 270.6000 ;
	    RECT 1177.8000 261.4500 1179.0000 261.6000 ;
	    RECT 1175.5500 260.5500 1179.0000 261.4500 ;
	    RECT 1177.8000 260.4000 1179.0000 260.5500 ;
	    RECT 1177.9501 258.6000 1178.8500 260.4000 ;
	    RECT 1180.3500 258.6000 1181.2500 269.4000 ;
	    RECT 1177.8000 257.4000 1179.0000 258.6000 ;
	    RECT 1180.2001 257.4000 1181.4000 258.6000 ;
	    RECT 1173.0000 227.4000 1174.2001 228.6000 ;
	    RECT 1163.4000 221.4000 1164.6000 222.6000 ;
	    RECT 1158.6000 203.4000 1159.8000 204.6000 ;
	    RECT 1158.6000 200.4000 1159.8000 201.6000 ;
	    RECT 1161.0000 200.4000 1162.2001 201.6000 ;
	    RECT 1158.7500 198.6000 1159.6500 200.4000 ;
	    RECT 1158.6000 197.4000 1159.8000 198.6000 ;
	    RECT 1156.2001 194.4000 1157.4000 195.6000 ;
	    RECT 1153.8000 191.4000 1155.0000 192.6000 ;
	    RECT 1146.6000 185.4000 1147.8000 186.6000 ;
	    RECT 1146.6000 176.4000 1147.8000 177.6000 ;
	    RECT 1146.7500 168.6000 1147.6500 176.4000 ;
	    RECT 1146.6000 167.4000 1147.8000 168.6000 ;
	    RECT 1149.0000 167.4000 1150.2001 168.6000 ;
	    RECT 1151.4000 167.4000 1152.6000 168.6000 ;
	    RECT 1144.2001 131.4000 1145.4000 132.6000 ;
	    RECT 1149.1500 114.6000 1150.0500 167.4000 ;
	    RECT 1151.5500 144.6000 1152.4501 167.4000 ;
	    RECT 1156.3500 162.6000 1157.2500 194.4000 ;
	    RECT 1158.6000 185.4000 1159.8000 186.6000 ;
	    RECT 1158.7500 174.6000 1159.6500 185.4000 ;
	    RECT 1158.6000 173.4000 1159.8000 174.6000 ;
	    RECT 1158.7500 162.6000 1159.6500 173.4000 ;
	    RECT 1161.1500 168.6000 1162.0500 200.4000 ;
	    RECT 1163.5500 186.6000 1164.4501 221.4000 ;
	    RECT 1182.7500 216.6000 1183.6500 341.4000 ;
	    RECT 1211.5500 324.6000 1212.4501 344.4000 ;
	    RECT 1221.1500 342.6000 1222.0500 440.4000 ;
	    RECT 1213.8000 341.4000 1215.0000 342.6000 ;
	    RECT 1221.0000 341.4000 1222.2001 342.6000 ;
	    RECT 1213.9501 324.6000 1214.8500 341.4000 ;
	    RECT 1225.8000 335.4000 1227.0000 336.6000 ;
	    RECT 1216.2001 329.4000 1217.4000 330.6000 ;
	    RECT 1223.4000 329.4000 1224.6000 330.6000 ;
	    RECT 1211.4000 323.4000 1212.6000 324.6000 ;
	    RECT 1213.8000 323.4000 1215.0000 324.6000 ;
	    RECT 1194.6000 320.4000 1195.8000 321.6000 ;
	    RECT 1189.8000 317.4000 1191.0000 318.6000 ;
	    RECT 1187.4000 311.4000 1188.6000 312.6000 ;
	    RECT 1185.0000 287.4000 1186.2001 288.6000 ;
	    RECT 1187.5500 285.6000 1188.4501 311.4000 ;
	    RECT 1189.9501 291.6000 1190.8500 317.4000 ;
	    RECT 1194.7500 312.6000 1195.6500 320.4000 ;
	    RECT 1194.6000 311.4000 1195.8000 312.6000 ;
	    RECT 1189.8000 290.4000 1191.0000 291.6000 ;
	    RECT 1211.5500 288.6000 1212.4501 323.4000 ;
	    RECT 1204.2001 287.4000 1205.4000 288.6000 ;
	    RECT 1206.6000 287.4000 1207.8000 288.6000 ;
	    RECT 1211.4000 287.4000 1212.6000 288.6000 ;
	    RECT 1187.4000 284.4000 1188.6000 285.6000 ;
	    RECT 1204.3500 282.6000 1205.2500 287.4000 ;
	    RECT 1187.4000 281.4000 1188.6000 282.6000 ;
	    RECT 1204.2001 281.4000 1205.4000 282.6000 ;
	    RECT 1187.5500 270.6000 1188.4501 281.4000 ;
	    RECT 1194.6000 275.4000 1195.8000 276.6000 ;
	    RECT 1211.4000 275.4000 1212.6000 276.6000 ;
	    RECT 1213.8000 275.4000 1215.0000 276.6000 ;
	    RECT 1187.4000 269.4000 1188.6000 270.6000 ;
	    RECT 1192.2001 233.4000 1193.4000 234.6000 ;
	    RECT 1185.0000 227.4000 1186.2001 228.6000 ;
	    RECT 1170.6000 215.4000 1171.8000 216.6000 ;
	    RECT 1182.6000 215.4000 1183.8000 216.6000 ;
	    RECT 1168.2001 201.4500 1169.4000 201.6000 ;
	    RECT 1170.7500 201.4500 1171.6500 215.4000 ;
	    RECT 1185.1500 204.6000 1186.0500 227.4000 ;
	    RECT 1187.4000 224.4000 1188.6000 225.6000 ;
	    RECT 1187.5500 222.6000 1188.4501 224.4000 ;
	    RECT 1194.7500 222.6000 1195.6500 275.4000 ;
	    RECT 1206.6000 269.4000 1207.8000 270.6000 ;
	    RECT 1204.2001 263.4000 1205.4000 264.6000 ;
	    RECT 1204.3500 255.6000 1205.2500 263.4000 ;
	    RECT 1204.2001 254.4000 1205.4000 255.6000 ;
	    RECT 1206.7500 252.6000 1207.6500 269.4000 ;
	    RECT 1209.0000 257.4000 1210.2001 258.6000 ;
	    RECT 1211.5500 255.6000 1212.4501 275.4000 ;
	    RECT 1213.9501 270.6000 1214.8500 275.4000 ;
	    RECT 1213.8000 269.4000 1215.0000 270.6000 ;
	    RECT 1211.4000 254.4000 1212.6000 255.6000 ;
	    RECT 1206.6000 251.4000 1207.8000 252.6000 ;
	    RECT 1197.0000 245.4000 1198.2001 246.6000 ;
	    RECT 1206.6000 245.4000 1207.8000 246.6000 ;
	    RECT 1197.1500 228.6000 1198.0500 245.4000 ;
	    RECT 1201.8000 233.4000 1203.0000 234.6000 ;
	    RECT 1197.0000 227.4000 1198.2001 228.6000 ;
	    RECT 1201.9501 225.6000 1202.8500 233.4000 ;
	    RECT 1206.7500 228.6000 1207.6500 245.4000 ;
	    RECT 1209.0000 239.4000 1210.2001 240.6000 ;
	    RECT 1206.6000 227.4000 1207.8000 228.6000 ;
	    RECT 1209.1500 225.6000 1210.0500 239.4000 ;
	    RECT 1201.8000 224.4000 1203.0000 225.6000 ;
	    RECT 1209.0000 224.4000 1210.2001 225.6000 ;
	    RECT 1211.4000 224.4000 1212.6000 225.6000 ;
	    RECT 1187.4000 221.4000 1188.6000 222.6000 ;
	    RECT 1194.6000 221.4000 1195.8000 222.6000 ;
	    RECT 1204.2001 221.4000 1205.4000 222.6000 ;
	    RECT 1209.0000 221.4000 1210.2001 222.6000 ;
	    RECT 1199.4000 215.4000 1200.6000 216.6000 ;
	    RECT 1185.0000 203.4000 1186.2001 204.6000 ;
	    RECT 1168.2001 200.5500 1171.6500 201.4500 ;
	    RECT 1168.2001 200.4000 1169.4000 200.5500 ;
	    RECT 1163.4000 185.4000 1164.6000 186.6000 ;
	    RECT 1163.4000 179.4000 1164.6000 180.6000 ;
	    RECT 1163.5500 177.6000 1164.4501 179.4000 ;
	    RECT 1163.4000 176.4000 1164.6000 177.6000 ;
	    RECT 1180.2001 173.4000 1181.4000 174.6000 ;
	    RECT 1161.0000 167.4000 1162.2001 168.6000 ;
	    RECT 1170.6000 167.4000 1171.8000 168.6000 ;
	    RECT 1173.0000 168.4500 1174.2001 168.6000 ;
	    RECT 1173.0000 167.5500 1176.4501 168.4500 ;
	    RECT 1173.0000 167.4000 1174.2001 167.5500 ;
	    RECT 1156.2001 161.4000 1157.4000 162.6000 ;
	    RECT 1158.6000 161.4000 1159.8000 162.6000 ;
	    RECT 1165.8000 161.4000 1167.0000 162.6000 ;
	    RECT 1151.4000 143.4000 1152.6000 144.6000 ;
	    RECT 1153.8000 142.5000 1155.0000 143.7000 ;
	    RECT 1155.9000 142.5000 1162.2001 143.4000 ;
	    RECT 1163.7001 142.5000 1164.9000 143.7000 ;
	    RECT 1153.8000 141.3000 1154.7001 142.5000 ;
	    RECT 1155.9000 142.2000 1157.1000 142.5000 ;
	    RECT 1161.0000 142.2000 1162.2001 142.5000 ;
	    RECT 1153.8000 140.4000 1161.0000 141.3000 ;
	    RECT 1153.8000 135.3000 1154.7001 140.4000 ;
	    RECT 1159.8000 140.1000 1161.0000 140.4000 ;
	    RECT 1156.2001 137.4000 1157.4000 138.6000 ;
	    RECT 1153.8000 134.1000 1155.0000 135.3000 ;
	    RECT 1153.8000 131.4000 1155.0000 132.6000 ;
	    RECT 1149.0000 113.4000 1150.2001 114.6000 ;
	    RECT 1144.2001 108.4500 1145.4000 108.6000 ;
	    RECT 1144.2001 107.5500 1147.6500 108.4500 ;
	    RECT 1144.2001 107.4000 1145.4000 107.5500 ;
	    RECT 1146.7500 102.6000 1147.6500 107.5500 ;
	    RECT 1146.6000 101.4000 1147.8000 102.6000 ;
	    RECT 1153.9501 96.4500 1154.8500 131.4000 ;
	    RECT 1156.3500 105.6000 1157.2500 137.4000 ;
	    RECT 1164.0000 135.3000 1164.9000 142.5000 ;
	    RECT 1163.7001 134.1000 1164.9000 135.3000 ;
	    RECT 1156.2001 104.4000 1157.4000 105.6000 ;
	    RECT 1165.9501 102.6000 1166.8500 161.4000 ;
	    RECT 1170.7500 150.6000 1171.6500 167.4000 ;
	    RECT 1173.0000 164.4000 1174.2001 165.6000 ;
	    RECT 1173.1500 162.6000 1174.0500 164.4000 ;
	    RECT 1173.0000 161.4000 1174.2001 162.6000 ;
	    RECT 1170.6000 149.4000 1171.8000 150.6000 ;
	    RECT 1168.2001 140.4000 1169.4000 141.6000 ;
	    RECT 1168.3500 120.6000 1169.2500 140.4000 ;
	    RECT 1173.1500 138.6000 1174.0500 161.4000 ;
	    RECT 1173.0000 137.4000 1174.2001 138.6000 ;
	    RECT 1175.5500 120.6000 1176.4501 167.5500 ;
	    RECT 1180.3500 165.6000 1181.2500 173.4000 ;
	    RECT 1180.2001 164.4000 1181.4000 165.6000 ;
	    RECT 1180.3500 144.6000 1181.2500 164.4000 ;
	    RECT 1185.1500 162.6000 1186.0500 203.4000 ;
	    RECT 1187.4000 179.4000 1188.6000 180.6000 ;
	    RECT 1185.0000 161.4000 1186.2001 162.6000 ;
	    RECT 1180.2001 143.4000 1181.4000 144.6000 ;
	    RECT 1180.2001 140.4000 1181.4000 141.6000 ;
	    RECT 1168.2001 119.4000 1169.4000 120.6000 ;
	    RECT 1175.4000 119.4000 1176.6000 120.6000 ;
	    RECT 1168.3500 102.6000 1169.2500 119.4000 ;
	    RECT 1170.6000 107.4000 1171.8000 108.6000 ;
	    RECT 1158.6000 101.4000 1159.8000 102.6000 ;
	    RECT 1165.8000 101.4000 1167.0000 102.6000 ;
	    RECT 1168.2001 101.4000 1169.4000 102.6000 ;
	    RECT 1156.2001 96.4500 1157.4000 96.6000 ;
	    RECT 1153.9501 95.5500 1157.4000 96.4500 ;
	    RECT 1156.2001 95.4000 1157.4000 95.5500 ;
	    RECT 1144.2001 66.3000 1145.4000 86.7000 ;
	    RECT 1146.6000 66.3000 1147.8000 86.7000 ;
	    RECT 1149.0000 66.3000 1150.2001 86.7000 ;
	    RECT 1151.4000 69.3000 1152.6000 86.7000 ;
	    RECT 1153.8000 83.4000 1155.0000 84.6000 ;
	    RECT 1153.9501 72.6000 1154.8500 83.4000 ;
	    RECT 1153.8000 71.4000 1155.0000 72.6000 ;
	    RECT 1156.2001 69.3000 1157.4000 86.7000 ;
	    RECT 1158.7500 81.6000 1159.6500 101.4000 ;
	    RECT 1168.2001 95.4000 1169.4000 96.6000 ;
	    RECT 1158.6000 80.4000 1159.8000 81.6000 ;
	    RECT 1161.0000 69.3000 1162.2001 86.7000 ;
	    RECT 1156.2001 65.4000 1157.4000 66.6000 ;
	    RECT 1163.4000 66.3000 1164.6000 86.7000 ;
	    RECT 1165.8000 66.3000 1167.0000 86.7000 ;
	    RECT 1168.3500 78.6000 1169.2500 95.4000 ;
	    RECT 1168.2001 77.4000 1169.4000 78.6000 ;
	    RECT 1170.7500 66.6000 1171.6500 107.4000 ;
	    RECT 1180.3500 105.6000 1181.2500 140.4000 ;
	    RECT 1187.5500 138.6000 1188.4501 179.4000 ;
	    RECT 1197.0000 167.4000 1198.2001 168.6000 ;
	    RECT 1197.1500 162.6000 1198.0500 167.4000 ;
	    RECT 1199.5500 165.6000 1200.4501 215.4000 ;
	    RECT 1204.3500 210.6000 1205.2500 221.4000 ;
	    RECT 1204.2001 209.4000 1205.4000 210.6000 ;
	    RECT 1209.1500 201.6000 1210.0500 221.4000 ;
	    RECT 1209.0000 200.4000 1210.2001 201.6000 ;
	    RECT 1209.1500 198.6000 1210.0500 200.4000 ;
	    RECT 1211.5500 198.6000 1212.4501 224.4000 ;
	    RECT 1216.3500 204.4500 1217.2500 329.4000 ;
	    RECT 1221.0000 317.4000 1222.2001 318.6000 ;
	    RECT 1221.1500 294.6000 1222.0500 317.4000 ;
	    RECT 1221.0000 293.4000 1222.2001 294.6000 ;
	    RECT 1221.0000 290.4000 1222.2001 291.6000 ;
	    RECT 1218.6000 284.4000 1219.8000 285.6000 ;
	    RECT 1218.7500 258.6000 1219.6500 284.4000 ;
	    RECT 1221.1500 264.6000 1222.0500 290.4000 ;
	    RECT 1221.0000 263.4000 1222.2001 264.6000 ;
	    RECT 1218.6000 257.4000 1219.8000 258.6000 ;
	    RECT 1218.7500 252.6000 1219.6500 257.4000 ;
	    RECT 1218.6000 251.4000 1219.8000 252.6000 ;
	    RECT 1221.0000 221.4000 1222.2001 222.6000 ;
	    RECT 1213.9501 203.5500 1217.2500 204.4500 ;
	    RECT 1209.0000 197.4000 1210.2001 198.6000 ;
	    RECT 1211.4000 197.4000 1212.6000 198.6000 ;
	    RECT 1204.2001 185.4000 1205.4000 186.6000 ;
	    RECT 1201.8000 167.4000 1203.0000 168.6000 ;
	    RECT 1199.4000 164.4000 1200.6000 165.6000 ;
	    RECT 1197.0000 161.4000 1198.2001 162.6000 ;
	    RECT 1197.1500 156.6000 1198.0500 161.4000 ;
	    RECT 1197.0000 155.4000 1198.2001 156.6000 ;
	    RECT 1187.4000 137.4000 1188.6000 138.6000 ;
	    RECT 1185.0000 119.4000 1186.2001 120.6000 ;
	    RECT 1185.1500 108.6000 1186.0500 119.4000 ;
	    RECT 1185.0000 107.4000 1186.2001 108.6000 ;
	    RECT 1177.8000 104.4000 1179.0000 105.6000 ;
	    RECT 1180.2001 104.4000 1181.4000 105.6000 ;
	    RECT 1175.4000 101.4000 1176.6000 102.6000 ;
	    RECT 1175.5500 84.6000 1176.4501 101.4000 ;
	    RECT 1177.9501 90.6000 1178.8500 104.4000 ;
	    RECT 1177.8000 89.4000 1179.0000 90.6000 ;
	    RECT 1175.4000 83.4000 1176.6000 84.6000 ;
	    RECT 1180.3500 81.6000 1181.2500 104.4000 ;
	    RECT 1201.9501 96.6000 1202.8500 167.4000 ;
	    RECT 1204.3500 159.6000 1205.2500 185.4000 ;
	    RECT 1204.2001 158.4000 1205.4000 159.6000 ;
	    RECT 1211.4000 149.4000 1212.6000 150.6000 ;
	    RECT 1211.5500 144.6000 1212.4501 149.4000 ;
	    RECT 1211.4000 143.4000 1212.6000 144.6000 ;
	    RECT 1211.5500 141.6000 1212.4501 143.4000 ;
	    RECT 1211.4000 140.4000 1212.6000 141.6000 ;
	    RECT 1213.9501 141.4500 1214.8500 203.5500 ;
	    RECT 1221.1500 201.6000 1222.0500 221.4000 ;
	    RECT 1221.0000 200.4000 1222.2001 201.6000 ;
	    RECT 1216.2001 197.4000 1217.4000 198.6000 ;
	    RECT 1216.3500 195.6000 1217.2500 197.4000 ;
	    RECT 1216.2001 194.4000 1217.4000 195.6000 ;
	    RECT 1223.5500 168.6000 1224.4501 329.4000 ;
	    RECT 1225.9501 321.6000 1226.8500 335.4000 ;
	    RECT 1225.8000 320.4000 1227.0000 321.6000 ;
	    RECT 1225.9501 186.6000 1226.8500 320.4000 ;
	    RECT 1228.2001 293.4000 1229.4000 294.6000 ;
	    RECT 1228.3500 222.6000 1229.2500 293.4000 ;
	    RECT 1228.2001 221.4000 1229.4000 222.6000 ;
	    RECT 1225.8000 185.4000 1227.0000 186.6000 ;
	    RECT 1223.4000 167.4000 1224.6000 168.6000 ;
	    RECT 1218.6000 149.4000 1219.8000 150.6000 ;
	    RECT 1213.9501 140.5500 1217.2500 141.4500 ;
	    RECT 1213.8000 137.4000 1215.0000 138.6000 ;
	    RECT 1209.0000 131.4000 1210.2001 132.6000 ;
	    RECT 1209.1500 108.6000 1210.0500 131.4000 ;
	    RECT 1206.6000 107.4000 1207.8000 108.6000 ;
	    RECT 1209.0000 107.4000 1210.2001 108.6000 ;
	    RECT 1206.7500 102.6000 1207.6500 107.4000 ;
	    RECT 1213.8000 104.4000 1215.0000 105.6000 ;
	    RECT 1206.6000 101.4000 1207.8000 102.6000 ;
	    RECT 1209.0000 101.4000 1210.2001 102.6000 ;
	    RECT 1201.8000 95.4000 1203.0000 96.6000 ;
	    RECT 1185.0000 83.4000 1186.2001 84.6000 ;
	    RECT 1180.2001 80.4000 1181.4000 81.6000 ;
	    RECT 1185.1500 78.6000 1186.0500 83.4000 ;
	    RECT 1185.0000 77.4000 1186.2001 78.6000 ;
	    RECT 1173.0000 74.4000 1174.2001 75.6000 ;
	    RECT 1173.1500 66.6000 1174.0500 74.4000 ;
	    RECT 1170.6000 65.4000 1171.8000 66.6000 ;
	    RECT 1173.0000 65.4000 1174.2001 66.6000 ;
	    RECT 1177.8000 65.4000 1179.0000 66.6000 ;
	    RECT 1144.5000 47.7000 1145.7001 48.9000 ;
	    RECT 1153.8000 47.7000 1155.0000 48.9000 ;
	    RECT 1141.8000 41.4000 1143.0000 42.6000 ;
	    RECT 1144.5000 40.5000 1145.4000 47.7000 ;
	    RECT 1146.3000 44.7000 1147.5000 45.9000 ;
	    RECT 1146.6000 42.6000 1147.5000 44.7000 ;
	    RECT 1154.1000 42.6000 1155.0000 47.7000 ;
	    RECT 1156.3500 42.6000 1157.2500 65.4000 ;
	    RECT 1173.0000 62.4000 1174.2001 63.6000 ;
	    RECT 1173.1500 60.6000 1174.0500 62.4000 ;
	    RECT 1173.0000 59.4000 1174.2001 60.6000 ;
	    RECT 1173.0000 53.4000 1174.2001 54.6000 ;
	    RECT 1170.6000 47.4000 1171.8000 48.6000 ;
	    RECT 1146.6000 41.7000 1155.0000 42.6000 ;
	    RECT 1146.6000 40.5000 1147.8000 40.8000 ;
	    RECT 1151.7001 40.5000 1152.9000 40.8000 ;
	    RECT 1154.1000 40.5000 1155.0000 41.7000 ;
	    RECT 1156.2001 41.4000 1157.4000 42.6000 ;
	    RECT 1170.7500 42.4500 1171.6500 47.4000 ;
	    RECT 1173.1500 45.6000 1174.0500 53.4000 ;
	    RECT 1175.4000 47.4000 1176.6000 48.6000 ;
	    RECT 1177.9501 45.6000 1178.8500 65.4000 ;
	    RECT 1180.2001 59.4000 1181.4000 60.6000 ;
	    RECT 1173.0000 44.4000 1174.2001 45.6000 ;
	    RECT 1177.8000 44.4000 1179.0000 45.6000 ;
	    RECT 1180.3500 42.6000 1181.2500 59.4000 ;
	    RECT 1182.6000 47.4000 1183.8000 48.6000 ;
	    RECT 1173.0000 42.4500 1174.2001 42.6000 ;
	    RECT 1170.7500 41.5500 1174.2001 42.4500 ;
	    RECT 1173.0000 41.4000 1174.2001 41.5500 ;
	    RECT 1180.2001 41.4000 1181.4000 42.6000 ;
	    RECT 1144.5000 39.6000 1152.9000 40.5000 ;
	    RECT 1144.5000 39.3000 1145.7001 39.6000 ;
	    RECT 1153.8000 39.3000 1155.0000 40.5000 ;
	    RECT 1182.7500 39.6000 1183.6500 47.4000 ;
	    RECT 1206.6000 41.4000 1207.8000 42.6000 ;
	    RECT 1182.6000 38.4000 1183.8000 39.6000 ;
	    RECT 1194.6000 38.4000 1195.8000 39.6000 ;
	    RECT 1074.6000 29.4000 1075.8000 30.6000 ;
	    RECT 1194.7500 12.6000 1195.6500 38.4000 ;
	    RECT 1209.1500 24.6000 1210.0500 101.4000 ;
	    RECT 1213.9501 45.6000 1214.8500 104.4000 ;
	    RECT 1216.3500 60.6000 1217.2500 140.5500 ;
	    RECT 1218.7500 138.6000 1219.6500 149.4000 ;
	    RECT 1218.6000 137.4000 1219.8000 138.6000 ;
	    RECT 1223.4000 137.4000 1224.6000 138.6000 ;
	    RECT 1223.5500 78.6000 1224.4501 137.4000 ;
	    RECT 1230.7500 132.6000 1231.6500 623.4000 ;
	    RECT 1242.6000 617.4000 1243.8000 618.6000 ;
	    RECT 1242.7500 582.6000 1243.6500 617.4000 ;
	    RECT 1247.4000 614.4000 1248.6000 615.6000 ;
	    RECT 1247.5500 612.6000 1248.4501 614.4000 ;
	    RECT 1247.4000 611.4000 1248.6000 612.6000 ;
	    RECT 1252.3500 606.6000 1253.2500 641.4000 ;
	    RECT 1276.3500 621.6000 1277.2500 641.4000 ;
	    RECT 1278.7500 624.6000 1279.6500 677.4000 ;
	    RECT 1293.1500 675.6000 1294.0500 983.4000 ;
	    RECT 1300.3500 981.6000 1301.2500 1001.4000 ;
	    RECT 1307.4000 995.4000 1308.6000 996.6000 ;
	    RECT 1295.4000 980.4000 1296.6000 981.6000 ;
	    RECT 1300.2001 980.4000 1301.4000 981.6000 ;
	    RECT 1295.5500 930.6000 1296.4501 980.4000 ;
	    RECT 1295.4000 929.4000 1296.6000 930.6000 ;
	    RECT 1297.8000 737.4000 1299.0000 738.6000 ;
	    RECT 1300.3500 726.6000 1301.2500 980.4000 ;
	    RECT 1302.6000 977.4000 1303.8000 978.6000 ;
	    RECT 1302.6000 959.4000 1303.8000 960.6000 ;
	    RECT 1302.7500 948.6000 1303.6500 959.4000 ;
	    RECT 1307.5500 948.6000 1308.4501 995.4000 ;
	    RECT 1317.0000 980.4000 1318.2001 981.6000 ;
	    RECT 1302.6000 947.4000 1303.8000 948.6000 ;
	    RECT 1307.4000 947.4000 1308.6000 948.6000 ;
	    RECT 1307.5500 945.6000 1308.4501 947.4000 ;
	    RECT 1307.4000 944.4000 1308.6000 945.6000 ;
	    RECT 1309.8000 936.3000 1311.0000 956.7000 ;
	    RECT 1312.2001 936.3000 1313.4000 956.7000 ;
	    RECT 1314.6000 936.3000 1315.8000 953.7000 ;
	    RECT 1317.1500 942.6000 1318.0500 980.4000 ;
	    RECT 1321.9501 978.6000 1322.8500 1001.4000 ;
	    RECT 1321.8000 977.4000 1323.0000 978.6000 ;
	    RECT 1321.9501 960.6000 1322.8500 977.4000 ;
	    RECT 1326.7500 975.6000 1327.6500 1004.4000 ;
	    RECT 1329.1500 996.6000 1330.0500 1244.4000 ;
	    RECT 1343.4000 1220.4000 1344.6000 1221.6000 ;
	    RECT 1343.5500 1185.6000 1344.4501 1220.4000 ;
	    RECT 1343.4000 1184.4000 1344.6000 1185.6000 ;
	    RECT 1348.2001 1181.4000 1349.4000 1182.6000 ;
	    RECT 1343.4000 1175.4000 1344.6000 1176.6000 ;
	    RECT 1333.8000 1146.3000 1335.0000 1166.7001 ;
	    RECT 1336.2001 1146.3000 1337.4000 1166.7001 ;
	    RECT 1338.6000 1146.3000 1339.8000 1166.7001 ;
	    RECT 1341.0000 1149.3000 1342.2001 1166.7001 ;
	    RECT 1343.5500 1164.6000 1344.4501 1175.4000 ;
	    RECT 1348.3500 1170.6000 1349.2500 1181.4000 ;
	    RECT 1348.2001 1169.4000 1349.4000 1170.6000 ;
	    RECT 1343.4000 1163.4000 1344.6000 1164.6000 ;
	    RECT 1345.8000 1149.3000 1347.0000 1166.7001 ;
	    RECT 1348.2001 1160.4000 1349.4000 1161.6000 ;
	    RECT 1348.3500 1152.6000 1349.2500 1160.4000 ;
	    RECT 1348.2001 1151.4000 1349.4000 1152.6000 ;
	    RECT 1350.6000 1149.3000 1351.8000 1166.7001 ;
	    RECT 1353.0000 1146.3000 1354.2001 1166.7001 ;
	    RECT 1355.4000 1146.3000 1356.6000 1166.7001 ;
	    RECT 1357.8000 1157.4000 1359.0000 1158.6000 ;
	    RECT 1362.6000 1154.4000 1363.8000 1155.6000 ;
	    RECT 1362.7500 1143.6000 1363.6500 1154.4000 ;
	    RECT 1362.6000 1142.4000 1363.8000 1143.6000 ;
	    RECT 1362.7500 1140.6000 1363.6500 1142.4000 ;
	    RECT 1362.6000 1139.4000 1363.8000 1140.6000 ;
	    RECT 1343.4000 1127.4000 1344.6000 1128.6000 ;
	    RECT 1343.5500 1086.6000 1344.4501 1127.4000 ;
	    RECT 1362.7500 1122.6000 1363.6500 1139.4000 ;
	    RECT 1362.6000 1121.4000 1363.8000 1122.6000 ;
	    RECT 1348.2001 1100.4000 1349.4000 1101.6000 ;
	    RECT 1348.3500 1098.6000 1349.2500 1100.4000 ;
	    RECT 1367.5500 1098.6000 1368.4501 1247.4000 ;
	    RECT 1369.8000 1241.4000 1371.0000 1242.6000 ;
	    RECT 1377.0000 1241.4000 1378.2001 1242.6000 ;
	    RECT 1369.9501 1224.6000 1370.8500 1241.4000 ;
	    RECT 1379.5500 1239.4501 1380.4501 1301.4000 ;
	    RECT 1377.1500 1238.5500 1380.4501 1239.4501 ;
	    RECT 1369.8000 1223.4000 1371.0000 1224.6000 ;
	    RECT 1377.1500 1218.6000 1378.0500 1238.5500 ;
	    RECT 1391.4000 1238.4000 1392.6000 1239.6000 ;
	    RECT 1391.5500 1236.6000 1392.4501 1238.4000 ;
	    RECT 1391.4000 1235.4000 1392.6000 1236.6000 ;
	    RECT 1391.4000 1229.4000 1392.6000 1230.6000 ;
	    RECT 1377.0000 1217.4000 1378.2001 1218.6000 ;
	    RECT 1372.2001 1214.4000 1373.4000 1215.6000 ;
	    RECT 1372.3500 1206.6000 1373.2500 1214.4000 ;
	    RECT 1372.2001 1205.4000 1373.4000 1206.6000 ;
	    RECT 1374.6000 1121.4000 1375.8000 1122.6000 ;
	    RECT 1372.2001 1118.4000 1373.4000 1119.6000 ;
	    RECT 1372.3500 1104.6000 1373.2500 1118.4000 ;
	    RECT 1374.7500 1116.6000 1375.6500 1121.4000 ;
	    RECT 1374.6000 1115.4000 1375.8000 1116.6000 ;
	    RECT 1372.2001 1103.4000 1373.4000 1104.6000 ;
	    RECT 1374.6000 1100.4000 1375.8000 1101.6000 ;
	    RECT 1374.7500 1098.6000 1375.6500 1100.4000 ;
	    RECT 1348.2001 1097.4000 1349.4000 1098.6000 ;
	    RECT 1367.4000 1097.4000 1368.6000 1098.6000 ;
	    RECT 1374.6000 1097.4000 1375.8000 1098.6000 ;
	    RECT 1343.4000 1085.4000 1344.6000 1086.6000 ;
	    RECT 1345.8000 1076.4000 1347.0000 1077.6000 ;
	    RECT 1343.4000 1025.4000 1344.6000 1026.6000 ;
	    RECT 1341.0000 1007.4000 1342.2001 1008.6000 ;
	    RECT 1329.0000 995.4000 1330.2001 996.6000 ;
	    RECT 1333.8000 980.4000 1335.0000 981.6000 ;
	    RECT 1333.9501 978.6000 1334.8500 980.4000 ;
	    RECT 1333.8000 977.4000 1335.0000 978.6000 ;
	    RECT 1326.6000 974.4000 1327.8000 975.6000 ;
	    RECT 1321.8000 959.4000 1323.0000 960.6000 ;
	    RECT 1317.0000 941.4000 1318.2001 942.6000 ;
	    RECT 1317.0000 935.4000 1318.2001 936.6000 ;
	    RECT 1319.4000 936.3000 1320.6000 953.7000 ;
	    RECT 1321.8000 947.4000 1323.0000 948.6000 ;
	    RECT 1321.9501 942.6000 1322.8500 947.4000 ;
	    RECT 1321.8000 941.4000 1323.0000 942.6000 ;
	    RECT 1321.8000 938.4000 1323.0000 939.6000 ;
	    RECT 1321.9501 936.6000 1322.8500 938.4000 ;
	    RECT 1321.8000 935.4000 1323.0000 936.6000 ;
	    RECT 1324.2001 936.3000 1325.4000 953.7000 ;
	    RECT 1326.6000 936.3000 1327.8000 956.7000 ;
	    RECT 1329.0000 936.3000 1330.2001 956.7000 ;
	    RECT 1331.4000 936.3000 1332.6000 956.7000 ;
	    RECT 1333.8000 941.4000 1335.0000 942.6000 ;
	    RECT 1307.4000 906.3000 1308.6000 926.7000 ;
	    RECT 1309.8000 906.3000 1311.0000 926.7000 ;
	    RECT 1312.2001 906.3000 1313.4000 926.7000 ;
	    RECT 1314.6000 909.3000 1315.8000 926.7000 ;
	    RECT 1317.1500 924.6000 1318.0500 935.4000 ;
	    RECT 1319.4000 930.4500 1320.6000 930.6000 ;
	    RECT 1319.4000 929.5500 1322.8500 930.4500 ;
	    RECT 1319.4000 929.4000 1320.6000 929.5500 ;
	    RECT 1317.0000 923.4000 1318.2001 924.6000 ;
	    RECT 1317.1500 885.6000 1318.0500 923.4000 ;
	    RECT 1319.4000 909.3000 1320.6000 926.7000 ;
	    RECT 1321.9501 921.6000 1322.8500 929.5500 ;
	    RECT 1321.8000 920.4000 1323.0000 921.6000 ;
	    RECT 1324.2001 909.3000 1325.4000 926.7000 ;
	    RECT 1326.6000 906.3000 1327.8000 926.7000 ;
	    RECT 1329.0000 906.3000 1330.2001 926.7000 ;
	    RECT 1331.4000 918.4500 1332.6000 918.6000 ;
	    RECT 1333.9501 918.4500 1334.8500 941.4000 ;
	    RECT 1331.4000 917.5500 1334.8500 918.4500 ;
	    RECT 1331.4000 917.4000 1332.6000 917.5500 ;
	    RECT 1336.2001 914.4000 1337.4000 915.6000 ;
	    RECT 1336.3500 906.6000 1337.2500 914.4000 ;
	    RECT 1336.2001 905.4000 1337.4000 906.6000 ;
	    RECT 1321.8000 893.4000 1323.0000 894.6000 ;
	    RECT 1317.0000 884.4000 1318.2001 885.6000 ;
	    RECT 1317.1500 876.6000 1318.0500 884.4000 ;
	    RECT 1317.0000 875.4000 1318.2001 876.6000 ;
	    RECT 1319.4000 855.3000 1320.6000 863.7000 ;
	    RECT 1321.9501 861.6000 1322.8500 893.4000 ;
	    RECT 1341.1500 885.6000 1342.0500 1007.4000 ;
	    RECT 1341.0000 884.4000 1342.2001 885.6000 ;
	    RECT 1341.0000 881.4000 1342.2001 882.6000 ;
	    RECT 1341.1500 870.6000 1342.0500 881.4000 ;
	    RECT 1341.0000 869.4000 1342.2001 870.6000 ;
	    RECT 1321.8000 860.4000 1323.0000 861.6000 ;
	    RECT 1324.2001 849.3000 1325.4000 866.7000 ;
	    RECT 1329.0000 857.4000 1330.2001 858.6000 ;
	    RECT 1329.1500 837.6000 1330.0500 857.4000 ;
	    RECT 1338.6000 849.3000 1339.8000 866.7000 ;
	    RECT 1329.0000 836.4000 1330.2001 837.6000 ;
	    RECT 1341.0000 836.4000 1342.2001 837.6000 ;
	    RECT 1309.8000 797.4000 1311.0000 798.6000 ;
	    RECT 1305.0000 794.4000 1306.2001 795.6000 ;
	    RECT 1305.1500 786.6000 1306.0500 794.4000 ;
	    RECT 1305.0000 785.4000 1306.2001 786.6000 ;
	    RECT 1312.2001 786.3000 1313.4000 806.7000 ;
	    RECT 1314.6000 786.3000 1315.8000 806.7000 ;
	    RECT 1317.0000 789.3000 1318.2001 806.7000 ;
	    RECT 1319.4000 803.4000 1320.6000 804.6000 ;
	    RECT 1319.5500 801.6000 1320.4501 803.4000 ;
	    RECT 1319.4000 800.4000 1320.6000 801.6000 ;
	    RECT 1321.8000 789.3000 1323.0000 806.7000 ;
	    RECT 1324.2001 803.4000 1325.4000 804.6000 ;
	    RECT 1324.3500 786.6000 1325.2500 803.4000 ;
	    RECT 1326.6000 789.3000 1327.8000 806.7000 ;
	    RECT 1324.2001 785.4000 1325.4000 786.6000 ;
	    RECT 1329.0000 786.3000 1330.2001 806.7000 ;
	    RECT 1331.4000 786.3000 1332.6000 806.7000 ;
	    RECT 1333.8000 786.3000 1335.0000 806.7000 ;
	    RECT 1341.1500 798.6000 1342.0500 836.4000 ;
	    RECT 1341.0000 797.4000 1342.2001 798.6000 ;
	    RECT 1307.4000 759.3000 1308.6000 767.7000 ;
	    RECT 1309.8000 761.4000 1311.0000 762.6000 ;
	    RECT 1312.2001 756.3000 1313.4000 773.7000 ;
	    RECT 1314.6000 773.4000 1315.8000 774.6000 ;
	    RECT 1312.2001 741.4500 1313.4000 741.6000 ;
	    RECT 1314.7500 741.4500 1315.6500 773.4000 ;
	    RECT 1317.0000 764.4000 1318.2001 765.6000 ;
	    RECT 1317.1500 741.6000 1318.0500 764.4000 ;
	    RECT 1326.6000 756.3000 1327.8000 773.7000 ;
	    RECT 1333.8000 743.4000 1335.0000 744.6000 ;
	    RECT 1333.9501 741.6000 1334.8500 743.4000 ;
	    RECT 1343.5500 741.6000 1344.4501 1025.4000 ;
	    RECT 1345.9501 984.6000 1346.8500 1076.4000 ;
	    RECT 1350.6000 1064.4000 1351.8000 1065.6000 ;
	    RECT 1350.7500 1005.4500 1351.6500 1064.4000 ;
	    RECT 1360.5000 1043.4000 1361.7001 1043.7001 ;
	    RECT 1360.5000 1042.5000 1368.9000 1043.4000 ;
	    RECT 1369.8000 1042.5000 1371.0000 1043.7001 ;
	    RECT 1357.8000 1040.4000 1359.0000 1041.6000 ;
	    RECT 1357.9501 1005.6000 1358.8500 1040.4000 ;
	    RECT 1360.5000 1035.3000 1361.4000 1042.5000 ;
	    RECT 1362.6000 1042.2001 1363.8000 1042.5000 ;
	    RECT 1367.7001 1042.2001 1368.9000 1042.5000 ;
	    RECT 1370.1000 1041.3000 1371.0000 1042.5000 ;
	    RECT 1362.6000 1040.4000 1371.0000 1041.3000 ;
	    RECT 1372.2001 1040.4000 1373.4000 1041.6000 ;
	    RECT 1362.6000 1038.3000 1363.5000 1040.4000 ;
	    RECT 1362.3000 1037.1000 1363.5000 1038.3000 ;
	    RECT 1370.1000 1035.3000 1371.0000 1040.4000 ;
	    RECT 1360.5000 1034.1000 1361.7001 1035.3000 ;
	    RECT 1369.8000 1034.1000 1371.0000 1035.3000 ;
	    RECT 1372.3500 1032.6000 1373.2500 1040.4000 ;
	    RECT 1372.2001 1031.4000 1373.4000 1032.6000 ;
	    RECT 1350.7500 1004.5500 1354.0500 1005.4500 ;
	    RECT 1353.1500 1002.6000 1354.0500 1004.5500 ;
	    RECT 1357.8000 1004.4000 1359.0000 1005.6000 ;
	    RECT 1350.6000 1001.4000 1351.8000 1002.6000 ;
	    RECT 1353.0000 1001.4000 1354.2001 1002.6000 ;
	    RECT 1350.7500 996.6000 1351.6500 1001.4000 ;
	    RECT 1350.6000 995.4000 1351.8000 996.6000 ;
	    RECT 1345.8000 983.4000 1347.0000 984.6000 ;
	    RECT 1345.9501 951.6000 1346.8500 983.4000 ;
	    RECT 1353.0000 977.4000 1354.2001 978.6000 ;
	    RECT 1353.1500 966.6000 1354.0500 977.4000 ;
	    RECT 1353.0000 965.4000 1354.2001 966.6000 ;
	    RECT 1345.8000 950.4000 1347.0000 951.6000 ;
	    RECT 1374.7500 921.6000 1375.6500 1097.4000 ;
	    RECT 1377.1500 1047.6000 1378.0500 1217.4000 ;
	    RECT 1379.4000 1206.3000 1380.6000 1226.7001 ;
	    RECT 1381.8000 1206.3000 1383.0000 1226.7001 ;
	    RECT 1384.2001 1209.3000 1385.4000 1226.7001 ;
	    RECT 1386.6000 1223.4000 1387.8000 1224.6000 ;
	    RECT 1386.7500 1221.6000 1387.6500 1223.4000 ;
	    RECT 1386.6000 1220.4000 1387.8000 1221.6000 ;
	    RECT 1389.0000 1209.3000 1390.2001 1226.7001 ;
	    RECT 1391.5500 1224.6000 1392.4501 1229.4000 ;
	    RECT 1391.4000 1223.4000 1392.6000 1224.6000 ;
	    RECT 1391.5500 1212.6000 1392.4501 1223.4000 ;
	    RECT 1391.4000 1211.4000 1392.6000 1212.6000 ;
	    RECT 1393.8000 1209.3000 1395.0000 1226.7001 ;
	    RECT 1396.2001 1206.3000 1397.4000 1226.7001 ;
	    RECT 1398.6000 1206.3000 1399.8000 1226.7001 ;
	    RECT 1401.0000 1206.3000 1402.2001 1226.7001 ;
	    RECT 1393.8000 1187.4000 1395.0000 1188.6000 ;
	    RECT 1391.4000 1127.4000 1392.6000 1128.6000 ;
	    RECT 1391.5500 1122.6000 1392.4501 1127.4000 ;
	    RECT 1393.9501 1125.6000 1394.8500 1187.4000 ;
	    RECT 1393.8000 1124.4000 1395.0000 1125.6000 ;
	    RECT 1384.2001 1121.4000 1385.4000 1122.6000 ;
	    RECT 1391.4000 1121.4000 1392.6000 1122.6000 ;
	    RECT 1384.3500 1119.6000 1385.2500 1121.4000 ;
	    RECT 1384.2001 1118.4000 1385.4000 1119.6000 ;
	    RECT 1379.4000 1094.4000 1380.6000 1095.6000 ;
	    RECT 1377.0000 1046.4000 1378.2001 1047.6000 ;
	    RECT 1379.5500 1044.6000 1380.4501 1094.4000 ;
	    RECT 1384.3500 1077.6000 1385.2500 1118.4000 ;
	    RECT 1405.8000 1109.4000 1407.0000 1110.6000 ;
	    RECT 1386.6000 1103.4000 1387.8000 1104.6000 ;
	    RECT 1386.7500 1101.6000 1387.6500 1103.4000 ;
	    RECT 1405.9501 1101.6000 1406.8500 1109.4000 ;
	    RECT 1408.3500 1104.6000 1409.2500 1340.4000 ;
	    RECT 1413.0000 1241.4000 1414.2001 1242.6000 ;
	    RECT 1413.1500 1140.6000 1414.0500 1241.4000 ;
	    RECT 1415.4000 1235.4000 1416.6000 1236.6000 ;
	    RECT 1415.5500 1212.6000 1416.4501 1235.4000 ;
	    RECT 1417.9501 1224.6000 1418.8500 1340.4000 ;
	    RECT 1451.5500 1338.6000 1452.4501 1385.4000 ;
	    RECT 1477.8000 1379.4000 1479.0000 1380.6000 ;
	    RECT 1477.9501 1341.6000 1478.8500 1379.4000 ;
	    RECT 1480.2001 1376.4000 1481.4000 1377.6000 ;
	    RECT 1480.3500 1368.6000 1481.2500 1376.4000 ;
	    RECT 1480.2001 1367.4000 1481.4000 1368.6000 ;
	    RECT 1485.0000 1367.4000 1486.2001 1368.6000 ;
	    RECT 1485.1500 1365.6000 1486.0500 1367.4000 ;
	    RECT 1485.0000 1364.4000 1486.2001 1365.6000 ;
	    RECT 1487.4000 1356.3000 1488.6000 1376.7001 ;
	    RECT 1489.8000 1356.3000 1491.0000 1376.7001 ;
	    RECT 1492.2001 1356.3000 1493.4000 1373.7001 ;
	    RECT 1494.7500 1368.6000 1495.6500 1424.4000 ;
	    RECT 1497.1500 1404.6000 1498.0500 1439.4000 ;
	    RECT 1499.4000 1436.4000 1500.6000 1437.6000 ;
	    RECT 1499.5500 1428.6000 1500.4501 1436.4000 ;
	    RECT 1499.4000 1427.4000 1500.6000 1428.6000 ;
	    RECT 1506.6000 1421.4000 1507.8000 1422.6000 ;
	    RECT 1497.0000 1404.4501 1498.2001 1404.6000 ;
	    RECT 1497.0000 1403.5500 1500.4501 1404.4501 ;
	    RECT 1497.0000 1403.4000 1498.2001 1403.5500 ;
	    RECT 1494.6000 1367.4000 1495.8000 1368.6000 ;
	    RECT 1494.6000 1361.4000 1495.8000 1362.6000 ;
	    RECT 1494.7500 1350.6000 1495.6500 1361.4000 ;
	    RECT 1497.0000 1356.3000 1498.2001 1373.7001 ;
	    RECT 1499.5500 1359.6000 1500.4501 1403.5500 ;
	    RECT 1506.7500 1386.6000 1507.6500 1421.4000 ;
	    RECT 1523.5500 1419.6000 1524.4501 1451.4000 ;
	    RECT 1540.2001 1424.4000 1541.4000 1425.6000 ;
	    RECT 1523.4000 1418.4000 1524.6000 1419.6000 ;
	    RECT 1540.3500 1410.6000 1541.2500 1424.4000 ;
	    RECT 1513.8000 1409.4000 1515.0000 1410.6000 ;
	    RECT 1540.2001 1409.4000 1541.4000 1410.6000 ;
	    RECT 1506.6000 1385.4000 1507.8000 1386.6000 ;
	    RECT 1499.4000 1358.4000 1500.6000 1359.6000 ;
	    RECT 1499.4000 1355.4000 1500.6000 1356.6000 ;
	    RECT 1501.8000 1356.3000 1503.0000 1373.7001 ;
	    RECT 1504.2001 1356.3000 1505.4000 1376.7001 ;
	    RECT 1506.6000 1356.3000 1507.8000 1376.7001 ;
	    RECT 1509.0000 1356.3000 1510.2001 1376.7001 ;
	    RECT 1499.5500 1350.6000 1500.4501 1355.4000 ;
	    RECT 1494.6000 1349.4000 1495.8000 1350.6000 ;
	    RECT 1499.4000 1349.4000 1500.6000 1350.6000 ;
	    RECT 1513.9501 1344.6000 1514.8500 1409.4000 ;
	    RECT 1521.0000 1397.4000 1522.2001 1398.6000 ;
	    RECT 1516.2001 1394.4000 1517.4000 1395.6000 ;
	    RECT 1516.3500 1386.6000 1517.2500 1394.4000 ;
	    RECT 1516.2001 1385.4000 1517.4000 1386.6000 ;
	    RECT 1516.2001 1382.4000 1517.4000 1383.6000 ;
	    RECT 1516.3500 1374.6000 1517.2500 1382.4000 ;
	    RECT 1516.2001 1373.4000 1517.4000 1374.6000 ;
	    RECT 1521.1500 1368.6000 1522.0500 1397.4000 ;
	    RECT 1523.4000 1386.3000 1524.6000 1406.7001 ;
	    RECT 1525.8000 1386.3000 1527.0000 1406.7001 ;
	    RECT 1528.2001 1389.3000 1529.4000 1406.7001 ;
	    RECT 1530.6000 1400.4000 1531.8000 1401.6000 ;
	    RECT 1530.7500 1380.6000 1531.6500 1400.4000 ;
	    RECT 1533.0000 1389.3000 1534.2001 1406.7001 ;
	    RECT 1535.4000 1403.4000 1536.6000 1404.6000 ;
	    RECT 1537.8000 1389.3000 1539.0000 1406.7001 ;
	    RECT 1540.2001 1386.3000 1541.4000 1406.7001 ;
	    RECT 1542.6000 1386.3000 1543.8000 1406.7001 ;
	    RECT 1545.0000 1386.3000 1546.2001 1406.7001 ;
	    RECT 1530.6000 1379.4000 1531.8000 1380.6000 ;
	    RECT 1549.8000 1373.4000 1551.0000 1374.6000 ;
	    RECT 1523.4000 1370.4000 1524.6000 1371.6000 ;
	    RECT 1521.0000 1367.4000 1522.2001 1368.6000 ;
	    RECT 1516.2001 1361.4000 1517.4000 1362.6000 ;
	    RECT 1516.3500 1344.6000 1517.2500 1361.4000 ;
	    RECT 1513.8000 1343.4000 1515.0000 1344.6000 ;
	    RECT 1516.2001 1343.4000 1517.4000 1344.6000 ;
	    RECT 1453.8000 1340.4000 1455.0000 1341.6000 ;
	    RECT 1477.8000 1340.4000 1479.0000 1341.6000 ;
	    RECT 1485.0000 1340.4000 1486.2001 1341.6000 ;
	    RECT 1451.4000 1337.4000 1452.6000 1338.6000 ;
	    RECT 1444.2001 1334.4000 1445.4000 1335.6000 ;
	    RECT 1446.6000 1335.4501 1447.8000 1335.6000 ;
	    RECT 1446.6000 1334.5500 1450.0500 1335.4501 ;
	    RECT 1446.6000 1334.4000 1447.8000 1334.5500 ;
	    RECT 1444.3500 1320.6000 1445.2500 1334.4000 ;
	    RECT 1446.6000 1331.4000 1447.8000 1332.6000 ;
	    RECT 1444.2001 1319.4000 1445.4000 1320.6000 ;
	    RECT 1444.2001 1295.4000 1445.4000 1296.6000 ;
	    RECT 1427.4000 1247.4000 1428.6000 1248.6000 ;
	    RECT 1422.6000 1244.4000 1423.8000 1245.6000 ;
	    RECT 1417.8000 1223.4000 1419.0000 1224.6000 ;
	    RECT 1422.7500 1221.6000 1423.6500 1244.4000 ;
	    RECT 1444.3500 1242.6000 1445.2500 1295.4000 ;
	    RECT 1441.8000 1241.4000 1443.0000 1242.6000 ;
	    RECT 1444.2001 1241.4000 1445.4000 1242.6000 ;
	    RECT 1429.8000 1223.4000 1431.0000 1224.6000 ;
	    RECT 1422.6000 1220.4000 1423.8000 1221.6000 ;
	    RECT 1415.4000 1211.4000 1416.6000 1212.6000 ;
	    RECT 1429.9501 1191.6000 1430.8500 1223.4000 ;
	    RECT 1441.9501 1194.6000 1442.8500 1241.4000 ;
	    RECT 1441.8000 1193.4000 1443.0000 1194.6000 ;
	    RECT 1429.8000 1190.4000 1431.0000 1191.6000 ;
	    RECT 1413.0000 1139.4000 1414.2001 1140.6000 ;
	    RECT 1413.1500 1134.6000 1414.0500 1139.4000 ;
	    RECT 1413.0000 1133.4000 1414.2001 1134.6000 ;
	    RECT 1444.2001 1133.4000 1445.4000 1134.6000 ;
	    RECT 1413.1500 1122.6000 1414.0500 1133.4000 ;
	    RECT 1413.0000 1121.4000 1414.2001 1122.6000 ;
	    RECT 1427.4000 1118.4000 1428.6000 1119.6000 ;
	    RECT 1408.2001 1103.4000 1409.4000 1104.6000 ;
	    RECT 1386.6000 1100.4000 1387.8000 1101.6000 ;
	    RECT 1405.8000 1100.4000 1407.0000 1101.6000 ;
	    RECT 1386.6000 1097.4000 1387.8000 1098.6000 ;
	    RECT 1384.2001 1076.4000 1385.4000 1077.6000 ;
	    RECT 1379.4000 1043.4000 1380.6000 1044.6000 ;
	    RECT 1386.7500 1038.6000 1387.6500 1097.4000 ;
	    RECT 1393.8000 1094.4000 1395.0000 1095.6000 ;
	    RECT 1389.0000 1043.4000 1390.2001 1044.6000 ;
	    RECT 1386.6000 1037.4000 1387.8000 1038.6000 ;
	    RECT 1384.2001 1007.4000 1385.4000 1008.6000 ;
	    RECT 1379.4000 1004.4000 1380.6000 1005.6000 ;
	    RECT 1379.5500 999.4500 1380.4501 1004.4000 ;
	    RECT 1379.5500 998.5500 1382.8500 999.4500 ;
	    RECT 1379.4000 995.4000 1380.6000 996.6000 ;
	    RECT 1377.0000 980.4000 1378.2001 981.6000 ;
	    RECT 1377.1500 960.6000 1378.0500 980.4000 ;
	    RECT 1377.0000 959.4000 1378.2001 960.6000 ;
	    RECT 1379.5500 948.6000 1380.4501 995.4000 ;
	    RECT 1381.9501 984.6000 1382.8500 998.5500 ;
	    RECT 1384.3500 996.6000 1385.2500 1007.4000 ;
	    RECT 1389.1500 1002.6000 1390.0500 1043.4000 ;
	    RECT 1389.0000 1001.4000 1390.2001 1002.6000 ;
	    RECT 1386.6000 998.4000 1387.8000 999.6000 ;
	    RECT 1384.2001 996.4500 1385.4000 996.6000 ;
	    RECT 1386.7500 996.4500 1387.6500 998.4000 ;
	    RECT 1384.2001 995.5500 1387.6500 996.4500 ;
	    RECT 1384.2001 995.4000 1385.4000 995.5500 ;
	    RECT 1381.8000 983.4000 1383.0000 984.6000 ;
	    RECT 1386.6000 974.4000 1387.8000 975.6000 ;
	    RECT 1379.4000 947.4000 1380.6000 948.6000 ;
	    RECT 1384.2001 947.4000 1385.4000 948.6000 ;
	    RECT 1384.3500 945.6000 1385.2500 947.4000 ;
	    RECT 1384.2001 944.4000 1385.4000 945.6000 ;
	    RECT 1386.7500 930.6000 1387.6500 974.4000 ;
	    RECT 1389.1500 948.6000 1390.0500 1001.4000 ;
	    RECT 1391.4000 983.4000 1392.6000 984.6000 ;
	    RECT 1391.5500 972.6000 1392.4501 983.4000 ;
	    RECT 1393.9501 975.6000 1394.8500 1094.4000 ;
	    RECT 1408.3500 1071.6000 1409.2500 1103.4000 ;
	    RECT 1417.8000 1085.4000 1419.0000 1086.6000 ;
	    RECT 1417.9501 1074.6000 1418.8500 1085.4000 ;
	    RECT 1417.8000 1073.4000 1419.0000 1074.6000 ;
	    RECT 1408.2001 1070.4000 1409.4000 1071.6000 ;
	    RECT 1396.2001 1001.4000 1397.4000 1002.6000 ;
	    RECT 1396.3500 990.6000 1397.2500 1001.4000 ;
	    RECT 1396.2001 989.4000 1397.4000 990.6000 ;
	    RECT 1410.6000 977.4000 1411.8000 978.6000 ;
	    RECT 1393.8000 974.4000 1395.0000 975.6000 ;
	    RECT 1391.4000 971.4000 1392.6000 972.6000 ;
	    RECT 1408.2001 971.4000 1409.4000 972.6000 ;
	    RECT 1408.3500 951.6000 1409.2500 971.4000 ;
	    RECT 1408.2001 950.4000 1409.4000 951.6000 ;
	    RECT 1410.7500 948.6000 1411.6500 977.4000 ;
	    RECT 1413.0000 974.4000 1414.2001 975.6000 ;
	    RECT 1389.0000 947.4000 1390.2001 948.6000 ;
	    RECT 1410.6000 947.4000 1411.8000 948.6000 ;
	    RECT 1386.6000 929.4000 1387.8000 930.6000 ;
	    RECT 1389.1500 924.6000 1390.0500 947.4000 ;
	    RECT 1389.0000 923.4000 1390.2001 924.6000 ;
	    RECT 1374.6000 920.4000 1375.8000 921.6000 ;
	    RECT 1377.0000 920.4000 1378.2001 921.6000 ;
	    RECT 1367.4000 917.4000 1368.6000 918.6000 ;
	    RECT 1365.0000 863.4000 1366.2001 864.6000 ;
	    RECT 1365.1500 858.6000 1366.0500 863.4000 ;
	    RECT 1365.0000 857.4000 1366.2001 858.6000 ;
	    RECT 1348.2001 818.4000 1349.4000 819.6000 ;
	    RECT 1348.3500 792.6000 1349.2500 818.4000 ;
	    RECT 1348.2001 791.4000 1349.4000 792.6000 ;
	    RECT 1312.2001 740.5500 1315.6500 741.4500 ;
	    RECT 1312.2001 740.4000 1313.4000 740.5500 ;
	    RECT 1317.0000 740.4000 1318.2001 741.6000 ;
	    RECT 1333.8000 740.4000 1335.0000 741.6000 ;
	    RECT 1343.4000 740.4000 1344.6000 741.6000 ;
	    RECT 1300.2001 725.4000 1301.4000 726.6000 ;
	    RECT 1307.4000 725.4000 1308.6000 726.6000 ;
	    RECT 1300.2001 713.4000 1301.4000 714.6000 ;
	    RECT 1297.8000 707.4000 1299.0000 708.6000 ;
	    RECT 1300.3500 705.6000 1301.2500 713.4000 ;
	    RECT 1302.6000 711.4500 1303.8000 711.6000 ;
	    RECT 1302.6000 710.5500 1306.0500 711.4500 ;
	    RECT 1302.6000 710.4000 1303.8000 710.5500 ;
	    RECT 1300.2001 704.4000 1301.4000 705.6000 ;
	    RECT 1305.1500 702.6000 1306.0500 710.5500 ;
	    RECT 1305.0000 701.4000 1306.2001 702.6000 ;
	    RECT 1305.0000 683.4000 1306.2001 684.6000 ;
	    RECT 1297.8000 680.4000 1299.0000 681.6000 ;
	    RECT 1297.9501 678.6000 1298.8500 680.4000 ;
	    RECT 1297.8000 677.4000 1299.0000 678.6000 ;
	    RECT 1293.0000 674.4000 1294.2001 675.6000 ;
	    RECT 1305.1500 651.6000 1306.0500 683.4000 ;
	    RECT 1305.0000 650.4000 1306.2001 651.6000 ;
	    RECT 1297.8000 647.4000 1299.0000 648.6000 ;
	    RECT 1295.4000 641.4000 1296.6000 642.6000 ;
	    RECT 1285.8000 629.4000 1287.0000 630.6000 ;
	    RECT 1285.9501 624.6000 1286.8500 629.4000 ;
	    RECT 1278.6000 623.4000 1279.8000 624.6000 ;
	    RECT 1285.8000 623.4000 1287.0000 624.6000 ;
	    RECT 1276.2001 620.4000 1277.4000 621.6000 ;
	    RECT 1281.0000 620.4000 1282.2001 621.6000 ;
	    RECT 1278.6000 617.4000 1279.8000 618.6000 ;
	    RECT 1276.2001 611.4000 1277.4000 612.6000 ;
	    RECT 1245.0000 605.4000 1246.2001 606.6000 ;
	    RECT 1252.2001 605.4000 1253.4000 606.6000 ;
	    RECT 1245.1500 585.6000 1246.0500 605.4000 ;
	    RECT 1276.3500 588.6000 1277.2500 611.4000 ;
	    RECT 1278.7500 588.6000 1279.6500 617.4000 ;
	    RECT 1281.1500 594.6000 1282.0500 620.4000 ;
	    RECT 1281.0000 593.4000 1282.2001 594.6000 ;
	    RECT 1281.1500 591.6000 1282.0500 593.4000 ;
	    RECT 1281.0000 590.4000 1282.2001 591.6000 ;
	    RECT 1249.8000 587.4000 1251.0000 588.6000 ;
	    RECT 1276.2001 587.4000 1277.4000 588.6000 ;
	    RECT 1278.6000 587.4000 1279.8000 588.6000 ;
	    RECT 1283.4000 587.4000 1284.6000 588.6000 ;
	    RECT 1285.8000 587.4000 1287.0000 588.6000 ;
	    RECT 1245.0000 584.4000 1246.2001 585.6000 ;
	    RECT 1242.6000 581.4000 1243.8000 582.6000 ;
	    RECT 1249.9501 564.6000 1250.8500 587.4000 ;
	    RECT 1259.4000 584.4000 1260.6000 585.6000 ;
	    RECT 1245.0000 563.4000 1246.2001 564.6000 ;
	    RECT 1249.8000 563.4000 1251.0000 564.6000 ;
	    RECT 1240.2001 560.4000 1241.4000 561.6000 ;
	    RECT 1233.0000 557.4000 1234.2001 558.6000 ;
	    RECT 1233.1500 540.6000 1234.0500 557.4000 ;
	    RECT 1235.4000 551.4000 1236.6000 552.6000 ;
	    RECT 1233.0000 539.4000 1234.2001 540.6000 ;
	    RECT 1233.1500 402.6000 1234.0500 539.4000 ;
	    RECT 1235.5500 528.6000 1236.4501 551.4000 ;
	    RECT 1237.8000 530.4000 1239.0000 531.6000 ;
	    RECT 1235.4000 527.4000 1236.6000 528.6000 ;
	    RECT 1237.9501 504.4500 1238.8500 530.4000 ;
	    RECT 1240.3500 525.6000 1241.2500 560.4000 ;
	    RECT 1245.1500 546.6000 1246.0500 563.4000 ;
	    RECT 1249.8000 557.4000 1251.0000 558.6000 ;
	    RECT 1254.6000 557.4000 1255.8000 558.6000 ;
	    RECT 1249.9501 555.6000 1250.8500 557.4000 ;
	    RECT 1249.8000 554.4000 1251.0000 555.6000 ;
	    RECT 1252.2001 551.4000 1253.4000 552.6000 ;
	    RECT 1245.0000 545.4000 1246.2001 546.6000 ;
	    RECT 1252.3500 534.6000 1253.2500 551.4000 ;
	    RECT 1254.7500 540.6000 1255.6500 557.4000 ;
	    RECT 1259.5500 555.6000 1260.4501 584.4000 ;
	    RECT 1261.8000 581.4000 1263.0000 582.6000 ;
	    RECT 1264.2001 581.4000 1265.4000 582.6000 ;
	    RECT 1261.9501 570.6000 1262.8500 581.4000 ;
	    RECT 1261.8000 569.4000 1263.0000 570.6000 ;
	    RECT 1261.8000 560.4000 1263.0000 561.6000 ;
	    RECT 1259.4000 554.4000 1260.6000 555.6000 ;
	    RECT 1259.5500 546.6000 1260.4501 554.4000 ;
	    RECT 1261.9501 552.6000 1262.8500 560.4000 ;
	    RECT 1261.8000 551.4000 1263.0000 552.6000 ;
	    RECT 1259.4000 545.4000 1260.6000 546.6000 ;
	    RECT 1254.6000 539.4000 1255.8000 540.6000 ;
	    RECT 1252.2001 533.4000 1253.4000 534.6000 ;
	    RECT 1259.5500 528.6000 1260.4501 545.4000 ;
	    RECT 1242.6000 527.4000 1243.8000 528.6000 ;
	    RECT 1259.4000 527.4000 1260.6000 528.6000 ;
	    RECT 1240.2001 524.4000 1241.4000 525.6000 ;
	    RECT 1242.7500 522.6000 1243.6500 527.4000 ;
	    RECT 1242.6000 521.4000 1243.8000 522.6000 ;
	    RECT 1257.0000 509.4000 1258.2001 510.6000 ;
	    RECT 1235.5500 503.5500 1238.8500 504.4500 ;
	    RECT 1235.5500 468.6000 1236.4501 503.5500 ;
	    RECT 1257.1500 501.6000 1258.0500 509.4000 ;
	    RECT 1257.0000 500.4000 1258.2001 501.6000 ;
	    RECT 1254.6000 497.4000 1255.8000 498.6000 ;
	    RECT 1252.2001 494.4000 1253.4000 495.6000 ;
	    RECT 1252.3500 492.6000 1253.2500 494.4000 ;
	    RECT 1252.2001 491.4000 1253.4000 492.6000 ;
	    RECT 1245.0000 479.4000 1246.2001 480.6000 ;
	    RECT 1235.4000 467.4000 1236.6000 468.6000 ;
	    RECT 1237.8000 467.4000 1239.0000 468.6000 ;
	    RECT 1237.9501 465.4500 1238.8500 467.4000 ;
	    RECT 1235.5500 464.5500 1238.8500 465.4500 ;
	    RECT 1235.5500 462.6000 1236.4501 464.5500 ;
	    RECT 1240.2001 464.4000 1241.4000 465.6000 ;
	    RECT 1235.4000 461.4000 1236.6000 462.6000 ;
	    RECT 1240.3500 450.6000 1241.2500 464.4000 ;
	    RECT 1240.2001 449.4000 1241.4000 450.6000 ;
	    RECT 1245.1500 438.6000 1246.0500 479.4000 ;
	    RECT 1237.8000 437.4000 1239.0000 438.6000 ;
	    RECT 1245.0000 437.4000 1246.2001 438.6000 ;
	    RECT 1237.9501 435.6000 1238.8500 437.4000 ;
	    RECT 1237.8000 434.4000 1239.0000 435.6000 ;
	    RECT 1245.1500 420.6000 1246.0500 437.4000 ;
	    RECT 1254.7500 435.6000 1255.6500 497.4000 ;
	    RECT 1259.5500 462.6000 1260.4501 527.4000 ;
	    RECT 1261.8000 503.4000 1263.0000 504.6000 ;
	    RECT 1259.4000 461.4000 1260.6000 462.6000 ;
	    RECT 1261.8000 455.4000 1263.0000 456.6000 ;
	    RECT 1261.9501 435.6000 1262.8500 455.4000 ;
	    RECT 1254.6000 434.4000 1255.8000 435.6000 ;
	    RECT 1261.8000 434.4000 1263.0000 435.6000 ;
	    RECT 1247.4000 431.4000 1248.6000 432.6000 ;
	    RECT 1247.5500 426.6000 1248.4501 431.4000 ;
	    RECT 1247.4000 425.4000 1248.6000 426.6000 ;
	    RECT 1245.0000 419.4000 1246.2001 420.6000 ;
	    RECT 1237.8000 407.4000 1239.0000 408.6000 ;
	    RECT 1242.6000 404.4000 1243.8000 405.6000 ;
	    RECT 1233.0000 401.4000 1234.2001 402.6000 ;
	    RECT 1242.7500 384.6000 1243.6500 404.4000 ;
	    RECT 1245.0000 401.4000 1246.2001 402.6000 ;
	    RECT 1245.1500 396.6000 1246.0500 401.4000 ;
	    RECT 1245.0000 395.4000 1246.2001 396.6000 ;
	    RECT 1242.6000 383.4000 1243.8000 384.6000 ;
	    RECT 1240.2001 347.4000 1241.4000 348.6000 ;
	    RECT 1240.3500 324.6000 1241.2500 347.4000 ;
	    RECT 1240.2001 323.4000 1241.4000 324.6000 ;
	    RECT 1233.0000 317.4000 1234.2001 318.6000 ;
	    RECT 1233.1500 312.6000 1234.0500 317.4000 ;
	    RECT 1233.0000 311.4000 1234.2001 312.6000 ;
	    RECT 1235.4000 299.4000 1236.6000 300.6000 ;
	    RECT 1235.5500 261.6000 1236.4501 299.4000 ;
	    RECT 1242.7500 294.6000 1243.6500 383.4000 ;
	    RECT 1247.5500 348.6000 1248.4501 425.4000 ;
	    RECT 1249.8000 386.4000 1251.0000 387.6000 ;
	    RECT 1247.4000 347.4000 1248.6000 348.6000 ;
	    RECT 1245.0000 344.4000 1246.2001 345.6000 ;
	    RECT 1242.6000 293.4000 1243.8000 294.6000 ;
	    RECT 1235.4000 260.4000 1236.6000 261.6000 ;
	    RECT 1237.8000 257.4000 1239.0000 258.6000 ;
	    RECT 1233.0000 203.4000 1234.2001 204.6000 ;
	    RECT 1233.1500 186.6000 1234.0500 203.4000 ;
	    RECT 1237.9501 201.6000 1238.8500 257.4000 ;
	    RECT 1242.6000 254.4000 1243.8000 255.6000 ;
	    RECT 1242.7500 240.6000 1243.6500 254.4000 ;
	    RECT 1242.6000 239.4000 1243.8000 240.6000 ;
	    RECT 1245.1500 228.6000 1246.0500 344.4000 ;
	    RECT 1249.9501 318.6000 1250.8500 386.4000 ;
	    RECT 1257.0000 368.4000 1258.2001 369.6000 ;
	    RECT 1254.6000 320.4000 1255.8000 321.6000 ;
	    RECT 1249.8000 317.4000 1251.0000 318.6000 ;
	    RECT 1252.2001 317.4000 1253.4000 318.6000 ;
	    RECT 1247.4000 263.4000 1248.6000 264.6000 ;
	    RECT 1247.5500 258.6000 1248.4501 263.4000 ;
	    RECT 1247.4000 257.4000 1248.6000 258.6000 ;
	    RECT 1245.0000 227.4000 1246.2001 228.6000 ;
	    RECT 1249.9501 216.6000 1250.8500 317.4000 ;
	    RECT 1252.3500 285.6000 1253.2500 317.4000 ;
	    RECT 1254.7500 300.6000 1255.6500 320.4000 ;
	    RECT 1254.6000 299.4000 1255.8000 300.6000 ;
	    RECT 1252.2001 284.4000 1253.4000 285.6000 ;
	    RECT 1254.7500 282.6000 1255.6500 299.4000 ;
	    RECT 1257.1500 285.6000 1258.0500 368.4000 ;
	    RECT 1259.4000 347.4000 1260.6000 348.6000 ;
	    RECT 1259.5500 312.6000 1260.4501 347.4000 ;
	    RECT 1264.3500 342.6000 1265.2500 581.4000 ;
	    RECT 1269.0000 524.4000 1270.2001 525.6000 ;
	    RECT 1269.1500 522.6000 1270.0500 524.4000 ;
	    RECT 1269.0000 521.4000 1270.2001 522.6000 ;
	    RECT 1269.0000 473.4000 1270.2001 474.6000 ;
	    RECT 1266.6000 464.4000 1267.8000 465.6000 ;
	    RECT 1266.7500 456.6000 1267.6500 464.4000 ;
	    RECT 1269.1500 462.6000 1270.0500 473.4000 ;
	    RECT 1273.8000 467.4000 1275.0000 468.6000 ;
	    RECT 1269.0000 461.4000 1270.2001 462.6000 ;
	    RECT 1273.9501 459.6000 1274.8500 467.4000 ;
	    RECT 1273.8000 458.4000 1275.0000 459.6000 ;
	    RECT 1266.6000 455.4000 1267.8000 456.6000 ;
	    RECT 1276.3500 444.6000 1277.2500 587.4000 ;
	    RECT 1281.0000 581.4000 1282.2001 582.6000 ;
	    RECT 1281.1500 558.6000 1282.0500 581.4000 ;
	    RECT 1283.5500 561.6000 1284.4501 587.4000 ;
	    RECT 1283.4000 560.4000 1284.6000 561.6000 ;
	    RECT 1281.0000 557.4000 1282.2001 558.6000 ;
	    RECT 1278.6000 539.4000 1279.8000 540.6000 ;
	    RECT 1276.2001 443.4000 1277.4000 444.6000 ;
	    RECT 1276.2001 437.4000 1277.4000 438.6000 ;
	    RECT 1273.8000 431.4000 1275.0000 432.6000 ;
	    RECT 1273.9501 426.6000 1274.8500 431.4000 ;
	    RECT 1273.8000 425.4000 1275.0000 426.6000 ;
	    RECT 1276.3500 420.6000 1277.2500 437.4000 ;
	    RECT 1276.2001 419.4000 1277.4000 420.6000 ;
	    RECT 1273.8000 413.4000 1275.0000 414.6000 ;
	    RECT 1271.4000 407.4000 1272.6000 408.6000 ;
	    RECT 1271.5500 402.6000 1272.4501 407.4000 ;
	    RECT 1273.9501 402.6000 1274.8500 413.4000 ;
	    RECT 1276.2001 404.4000 1277.4000 405.6000 ;
	    RECT 1271.4000 401.4000 1272.6000 402.6000 ;
	    RECT 1273.8000 401.4000 1275.0000 402.6000 ;
	    RECT 1276.3500 378.6000 1277.2500 404.4000 ;
	    RECT 1278.7500 402.6000 1279.6500 539.4000 ;
	    RECT 1285.9501 528.6000 1286.8500 587.4000 ;
	    RECT 1288.2001 569.4000 1289.4000 570.6000 ;
	    RECT 1288.3500 564.6000 1289.2500 569.4000 ;
	    RECT 1288.2001 563.4000 1289.4000 564.6000 ;
	    RECT 1285.8000 527.4000 1287.0000 528.6000 ;
	    RECT 1290.6000 525.4500 1291.8000 525.6000 ;
	    RECT 1288.3500 524.5500 1291.8000 525.4500 ;
	    RECT 1283.4000 518.4000 1284.6000 519.6000 ;
	    RECT 1283.5500 498.6000 1284.4501 518.4000 ;
	    RECT 1285.8000 500.4000 1287.0000 501.6000 ;
	    RECT 1283.4000 497.4000 1284.6000 498.6000 ;
	    RECT 1285.9501 486.6000 1286.8500 500.4000 ;
	    RECT 1288.3500 498.6000 1289.2500 524.5500 ;
	    RECT 1290.6000 524.4000 1291.8000 524.5500 ;
	    RECT 1288.2001 497.4000 1289.4000 498.6000 ;
	    RECT 1293.0000 497.4000 1294.2001 498.6000 ;
	    RECT 1293.1500 495.6000 1294.0500 497.4000 ;
	    RECT 1293.0000 494.4000 1294.2001 495.6000 ;
	    RECT 1285.8000 485.4000 1287.0000 486.6000 ;
	    RECT 1285.9501 465.6000 1286.8500 485.4000 ;
	    RECT 1288.2001 467.4000 1289.4000 468.6000 ;
	    RECT 1285.8000 464.4000 1287.0000 465.6000 ;
	    RECT 1281.0000 455.4000 1282.2001 456.6000 ;
	    RECT 1281.1500 435.6000 1282.0500 455.4000 ;
	    RECT 1293.0000 443.4000 1294.2001 444.6000 ;
	    RECT 1281.0000 434.4000 1282.2001 435.6000 ;
	    RECT 1281.0000 407.4000 1282.2001 408.6000 ;
	    RECT 1281.1500 405.6000 1282.0500 407.4000 ;
	    RECT 1281.0000 404.4000 1282.2001 405.6000 ;
	    RECT 1278.6000 401.4000 1279.8000 402.6000 ;
	    RECT 1285.8000 401.4000 1287.0000 402.6000 ;
	    RECT 1276.2001 377.4000 1277.4000 378.6000 ;
	    RECT 1283.4000 377.4000 1284.6000 378.6000 ;
	    RECT 1273.8000 365.4000 1275.0000 366.6000 ;
	    RECT 1266.6000 359.4000 1267.8000 360.6000 ;
	    RECT 1264.2001 341.4000 1265.4000 342.6000 ;
	    RECT 1264.3500 336.6000 1265.2500 341.4000 ;
	    RECT 1264.2001 335.4000 1265.4000 336.6000 ;
	    RECT 1259.4000 311.4000 1260.6000 312.6000 ;
	    RECT 1257.0000 284.4000 1258.2001 285.6000 ;
	    RECT 1261.8000 284.4000 1263.0000 285.6000 ;
	    RECT 1254.6000 281.4000 1255.8000 282.6000 ;
	    RECT 1259.4000 281.4000 1260.6000 282.6000 ;
	    RECT 1257.0000 239.4000 1258.2001 240.6000 ;
	    RECT 1257.1500 222.6000 1258.0500 239.4000 ;
	    RECT 1259.5500 234.6000 1260.4501 281.4000 ;
	    RECT 1261.9501 252.6000 1262.8500 284.4000 ;
	    RECT 1266.7500 261.6000 1267.6500 359.4000 ;
	    RECT 1273.9501 345.6000 1274.8500 365.4000 ;
	    RECT 1273.8000 344.4000 1275.0000 345.6000 ;
	    RECT 1281.0000 344.4000 1282.2001 345.6000 ;
	    RECT 1278.6000 338.4000 1279.8000 339.6000 ;
	    RECT 1271.4000 335.4000 1272.6000 336.6000 ;
	    RECT 1271.5500 318.6000 1272.4501 335.4000 ;
	    RECT 1278.7500 330.6000 1279.6500 338.4000 ;
	    RECT 1278.6000 329.4000 1279.8000 330.6000 ;
	    RECT 1271.4000 317.4000 1272.6000 318.6000 ;
	    RECT 1273.8000 317.4000 1275.0000 318.6000 ;
	    RECT 1271.4000 305.4000 1272.6000 306.6000 ;
	    RECT 1271.5500 276.6000 1272.4501 305.4000 ;
	    RECT 1271.4000 275.4000 1272.6000 276.6000 ;
	    RECT 1266.6000 260.4000 1267.8000 261.6000 ;
	    RECT 1269.0000 260.4000 1270.2001 261.6000 ;
	    RECT 1269.1500 258.6000 1270.0500 260.4000 ;
	    RECT 1273.9501 258.6000 1274.8500 317.4000 ;
	    RECT 1276.2001 311.4000 1277.4000 312.6000 ;
	    RECT 1276.3500 279.6000 1277.2500 311.4000 ;
	    RECT 1276.2001 278.4000 1277.4000 279.6000 ;
	    RECT 1276.2001 275.4000 1277.4000 276.6000 ;
	    RECT 1276.3500 264.6000 1277.2500 275.4000 ;
	    RECT 1276.2001 263.4000 1277.4000 264.6000 ;
	    RECT 1269.0000 257.4000 1270.2001 258.6000 ;
	    RECT 1273.8000 257.4000 1275.0000 258.6000 ;
	    RECT 1276.3500 255.6000 1277.2500 263.4000 ;
	    RECT 1276.2001 254.4000 1277.4000 255.6000 ;
	    RECT 1261.8000 251.4000 1263.0000 252.6000 ;
	    RECT 1261.9501 246.6000 1262.8500 251.4000 ;
	    RECT 1261.8000 245.4000 1263.0000 246.6000 ;
	    RECT 1278.6000 245.4000 1279.8000 246.6000 ;
	    RECT 1278.7500 234.6000 1279.6500 245.4000 ;
	    RECT 1259.4000 233.4000 1260.6000 234.6000 ;
	    RECT 1278.6000 233.4000 1279.8000 234.6000 ;
	    RECT 1259.5500 228.6000 1260.4501 233.4000 ;
	    RECT 1261.8000 230.4000 1263.0000 231.6000 ;
	    RECT 1259.4000 227.4000 1260.6000 228.6000 ;
	    RECT 1261.9501 225.4500 1262.8500 230.4000 ;
	    RECT 1266.6000 227.4000 1267.8000 228.6000 ;
	    RECT 1259.5500 224.5500 1262.8500 225.4500 ;
	    RECT 1259.5500 222.6000 1260.4501 224.5500 ;
	    RECT 1264.2001 224.4000 1265.4000 225.6000 ;
	    RECT 1257.0000 221.4000 1258.2001 222.6000 ;
	    RECT 1259.4000 221.4000 1260.6000 222.6000 ;
	    RECT 1249.8000 215.4000 1251.0000 216.6000 ;
	    RECT 1257.0000 215.4000 1258.2001 216.6000 ;
	    RECT 1257.1500 201.6000 1258.0500 215.4000 ;
	    RECT 1264.3500 201.6000 1265.2500 224.4000 ;
	    RECT 1266.7500 216.6000 1267.6500 227.4000 ;
	    RECT 1278.6000 218.4000 1279.8000 219.6000 ;
	    RECT 1266.6000 215.4000 1267.8000 216.6000 ;
	    RECT 1276.2001 203.4000 1277.4000 204.6000 ;
	    RECT 1237.8000 200.4000 1239.0000 201.6000 ;
	    RECT 1257.0000 200.4000 1258.2001 201.6000 ;
	    RECT 1264.2001 200.4000 1265.4000 201.6000 ;
	    RECT 1257.1500 198.6000 1258.0500 200.4000 ;
	    RECT 1276.3500 198.6000 1277.2500 203.4000 ;
	    RECT 1278.7500 201.6000 1279.6500 218.4000 ;
	    RECT 1278.6000 200.4000 1279.8000 201.6000 ;
	    RECT 1257.0000 197.4000 1258.2001 198.6000 ;
	    RECT 1276.2001 197.4000 1277.4000 198.6000 ;
	    RECT 1281.1500 198.4500 1282.0500 344.4000 ;
	    RECT 1283.5500 216.6000 1284.4501 377.4000 ;
	    RECT 1285.9501 354.6000 1286.8500 401.4000 ;
	    RECT 1293.1500 399.6000 1294.0500 443.4000 ;
	    RECT 1295.5500 441.6000 1296.4501 641.4000 ;
	    RECT 1297.9501 516.6000 1298.8500 647.4000 ;
	    RECT 1302.6000 644.4000 1303.8000 645.6000 ;
	    RECT 1302.7500 642.6000 1303.6500 644.4000 ;
	    RECT 1302.6000 641.4000 1303.8000 642.6000 ;
	    RECT 1302.6000 623.4000 1303.8000 624.6000 ;
	    RECT 1305.0000 623.4000 1306.2001 624.6000 ;
	    RECT 1300.2001 614.4000 1301.4000 615.6000 ;
	    RECT 1300.3500 588.6000 1301.2500 614.4000 ;
	    RECT 1302.7500 612.6000 1303.6500 623.4000 ;
	    RECT 1305.1500 618.6000 1306.0500 623.4000 ;
	    RECT 1305.0000 617.4000 1306.2001 618.6000 ;
	    RECT 1302.6000 611.4000 1303.8000 612.6000 ;
	    RECT 1300.2001 587.4000 1301.4000 588.6000 ;
	    RECT 1300.2001 584.4000 1301.4000 585.6000 ;
	    RECT 1300.3500 576.6000 1301.2500 584.4000 ;
	    RECT 1300.2001 575.4000 1301.4000 576.6000 ;
	    RECT 1300.3500 570.6000 1301.2500 575.4000 ;
	    RECT 1300.2001 569.4000 1301.4000 570.6000 ;
	    RECT 1302.6000 521.4000 1303.8000 522.6000 ;
	    RECT 1297.8000 515.4000 1299.0000 516.6000 ;
	    RECT 1302.7500 498.6000 1303.6500 521.4000 ;
	    RECT 1302.6000 497.4000 1303.8000 498.6000 ;
	    RECT 1305.0000 473.4000 1306.2001 474.6000 ;
	    RECT 1305.1500 471.6000 1306.0500 473.4000 ;
	    RECT 1305.0000 470.4000 1306.2001 471.6000 ;
	    RECT 1302.6000 464.4000 1303.8000 465.6000 ;
	    RECT 1302.7500 456.6000 1303.6500 464.4000 ;
	    RECT 1302.6000 455.4000 1303.8000 456.6000 ;
	    RECT 1295.4000 440.4000 1296.6000 441.6000 ;
	    RECT 1293.0000 398.4000 1294.2001 399.6000 ;
	    RECT 1285.8000 353.4000 1287.0000 354.6000 ;
	    RECT 1285.9501 342.6000 1286.8500 353.4000 ;
	    RECT 1285.8000 341.4000 1287.0000 342.6000 ;
	    RECT 1295.5500 339.6000 1296.4501 440.4000 ;
	    RECT 1305.0000 434.4000 1306.2001 435.6000 ;
	    RECT 1305.1500 432.6000 1306.0500 434.4000 ;
	    RECT 1305.0000 431.4000 1306.2001 432.6000 ;
	    RECT 1297.8000 347.4000 1299.0000 348.6000 ;
	    RECT 1295.4000 338.4000 1296.6000 339.6000 ;
	    RECT 1290.6000 329.4000 1291.8000 330.6000 ;
	    RECT 1285.8000 323.4000 1287.0000 324.6000 ;
	    RECT 1285.9501 312.6000 1286.8500 323.4000 ;
	    RECT 1285.8000 311.4000 1287.0000 312.6000 ;
	    RECT 1290.7500 282.6000 1291.6500 329.4000 ;
	    RECT 1293.0000 320.4000 1294.2001 321.6000 ;
	    RECT 1293.1500 294.6000 1294.0500 320.4000 ;
	    RECT 1295.4000 317.4000 1296.6000 318.6000 ;
	    RECT 1293.0000 293.4000 1294.2001 294.6000 ;
	    RECT 1290.6000 281.4000 1291.8000 282.6000 ;
	    RECT 1285.8000 278.4000 1287.0000 279.6000 ;
	    RECT 1283.4000 215.4000 1284.6000 216.6000 ;
	    RECT 1278.7500 197.5500 1282.0500 198.4500 ;
	    RECT 1252.2001 194.4000 1253.4000 195.6000 ;
	    RECT 1233.0000 185.4000 1234.2001 186.6000 ;
	    RECT 1230.6000 131.4000 1231.8000 132.6000 ;
	    RECT 1233.1500 102.6000 1234.0500 185.4000 ;
	    RECT 1252.3500 174.6000 1253.2500 194.4000 ;
	    RECT 1252.2001 173.4000 1253.4000 174.6000 ;
	    RECT 1252.2001 143.4000 1253.4000 144.6000 ;
	    RECT 1271.4000 143.4000 1272.6000 144.6000 ;
	    RECT 1252.3500 141.6000 1253.2500 143.4000 ;
	    RECT 1242.6000 140.4000 1243.8000 141.6000 ;
	    RECT 1252.2001 140.4000 1253.4000 141.6000 ;
	    RECT 1240.2001 107.4000 1241.4000 108.6000 ;
	    RECT 1233.0000 101.4000 1234.2001 102.6000 ;
	    RECT 1235.4000 101.4000 1236.6000 102.6000 ;
	    RECT 1240.3500 96.6000 1241.2500 107.4000 ;
	    RECT 1242.7500 96.6000 1243.6500 140.4000 ;
	    RECT 1254.6000 137.4000 1255.8000 138.6000 ;
	    RECT 1259.4000 137.4000 1260.6000 138.6000 ;
	    RECT 1257.0000 131.4000 1258.2001 132.6000 ;
	    RECT 1247.4000 125.4000 1248.6000 126.6000 ;
	    RECT 1245.0000 107.4000 1246.2001 108.6000 ;
	    RECT 1240.2001 95.4000 1241.4000 96.6000 ;
	    RECT 1242.6000 95.4000 1243.8000 96.6000 ;
	    RECT 1240.2001 83.4000 1241.4000 84.6000 ;
	    RECT 1237.8000 80.4000 1239.0000 81.6000 ;
	    RECT 1223.4000 77.4000 1224.6000 78.6000 ;
	    RECT 1235.4000 71.4000 1236.6000 72.6000 ;
	    RECT 1216.2001 59.4000 1217.4000 60.6000 ;
	    RECT 1213.8000 44.4000 1215.0000 45.6000 ;
	    RECT 1209.0000 23.4000 1210.2001 24.6000 ;
	    RECT 1216.3500 18.6000 1217.2500 59.4000 ;
	    RECT 1235.5500 48.6000 1236.4501 71.4000 ;
	    RECT 1235.4000 47.4000 1236.6000 48.6000 ;
	    RECT 1237.9501 42.6000 1238.8500 80.4000 ;
	    RECT 1240.3500 78.6000 1241.2500 83.4000 ;
	    RECT 1242.7500 81.6000 1243.6500 95.4000 ;
	    RECT 1242.6000 80.4000 1243.8000 81.6000 ;
	    RECT 1245.1500 78.6000 1246.0500 107.4000 ;
	    RECT 1247.5500 102.6000 1248.4501 125.4000 ;
	    RECT 1257.1500 108.6000 1258.0500 131.4000 ;
	    RECT 1269.0000 113.4000 1270.2001 114.6000 ;
	    RECT 1257.0000 107.4000 1258.2001 108.6000 ;
	    RECT 1266.6000 107.4000 1267.8000 108.6000 ;
	    RECT 1247.4000 101.4000 1248.6000 102.6000 ;
	    RECT 1247.5500 81.6000 1248.4501 101.4000 ;
	    RECT 1249.8000 95.4000 1251.0000 96.6000 ;
	    RECT 1249.9501 81.6000 1250.8500 95.4000 ;
	    RECT 1247.4000 80.4000 1248.6000 81.6000 ;
	    RECT 1249.8000 80.4000 1251.0000 81.6000 ;
	    RECT 1240.2001 77.4000 1241.4000 78.6000 ;
	    RECT 1245.0000 77.4000 1246.2001 78.6000 ;
	    RECT 1257.1500 75.6000 1258.0500 107.4000 ;
	    RECT 1269.1500 105.6000 1270.0500 113.4000 ;
	    RECT 1266.6000 104.4000 1267.8000 105.6000 ;
	    RECT 1269.0000 104.4000 1270.2001 105.6000 ;
	    RECT 1266.7500 102.6000 1267.6500 104.4000 ;
	    RECT 1266.6000 101.4000 1267.8000 102.6000 ;
	    RECT 1269.1500 78.6000 1270.0500 104.4000 ;
	    RECT 1271.5500 102.6000 1272.4501 143.4000 ;
	    RECT 1278.7500 141.6000 1279.6500 197.5500 ;
	    RECT 1281.0000 194.4000 1282.2001 195.6000 ;
	    RECT 1281.1500 174.6000 1282.0500 194.4000 ;
	    RECT 1285.9501 186.6000 1286.8500 278.4000 ;
	    RECT 1290.7500 234.6000 1291.6500 281.4000 ;
	    RECT 1293.0000 263.4000 1294.2001 264.6000 ;
	    RECT 1293.1500 252.6000 1294.0500 263.4000 ;
	    RECT 1293.0000 251.4000 1294.2001 252.6000 ;
	    RECT 1290.6000 233.4000 1291.8000 234.6000 ;
	    RECT 1295.4000 233.4000 1296.6000 234.6000 ;
	    RECT 1290.6000 227.4000 1291.8000 228.6000 ;
	    RECT 1290.7500 222.6000 1291.6500 227.4000 ;
	    RECT 1293.0000 224.4000 1294.2001 225.6000 ;
	    RECT 1290.6000 221.4000 1291.8000 222.6000 ;
	    RECT 1288.2001 219.4500 1289.4000 219.6000 ;
	    RECT 1293.1500 219.4500 1294.0500 224.4000 ;
	    RECT 1288.2001 218.5500 1294.0500 219.4500 ;
	    RECT 1288.2001 218.4000 1289.4000 218.5500 ;
	    RECT 1288.2001 215.4000 1289.4000 216.6000 ;
	    RECT 1288.3500 201.6000 1289.2500 215.4000 ;
	    RECT 1288.2001 200.4000 1289.4000 201.6000 ;
	    RECT 1285.8000 185.4000 1287.0000 186.6000 ;
	    RECT 1281.0000 173.4000 1282.2001 174.6000 ;
	    RECT 1276.2001 140.4000 1277.4000 141.6000 ;
	    RECT 1278.6000 140.4000 1279.8000 141.6000 ;
	    RECT 1273.8000 113.4000 1275.0000 114.6000 ;
	    RECT 1273.9501 105.6000 1274.8500 113.4000 ;
	    RECT 1273.8000 104.4000 1275.0000 105.6000 ;
	    RECT 1276.3500 102.6000 1277.2500 140.4000 ;
	    RECT 1278.6000 137.4000 1279.8000 138.6000 ;
	    RECT 1278.7500 105.6000 1279.6500 137.4000 ;
	    RECT 1278.6000 104.4000 1279.8000 105.6000 ;
	    RECT 1271.4000 101.4000 1272.6000 102.6000 ;
	    RECT 1273.8000 101.4000 1275.0000 102.6000 ;
	    RECT 1276.2001 101.4000 1277.4000 102.6000 ;
	    RECT 1271.4000 95.4000 1272.6000 96.6000 ;
	    RECT 1273.9501 96.4500 1274.8500 101.4000 ;
	    RECT 1276.2001 96.4500 1277.4000 96.6000 ;
	    RECT 1273.9501 95.5500 1277.4000 96.4500 ;
	    RECT 1276.2001 95.4000 1277.4000 95.5500 ;
	    RECT 1269.0000 77.4000 1270.2001 78.6000 ;
	    RECT 1257.0000 74.4000 1258.2001 75.6000 ;
	    RECT 1245.0000 71.4000 1246.2001 72.6000 ;
	    RECT 1240.2001 47.7000 1241.4000 48.9000 ;
	    RECT 1240.2001 42.6000 1241.1000 47.7000 ;
	    RECT 1245.1500 45.6000 1246.0500 71.4000 ;
	    RECT 1249.5000 47.7000 1250.7001 48.9000 ;
	    RECT 1245.0000 44.4000 1246.2001 45.6000 ;
	    RECT 1247.7001 44.7000 1248.9000 45.9000 ;
	    RECT 1247.7001 42.6000 1248.6000 44.7000 ;
	    RECT 1237.8000 41.4000 1239.0000 42.6000 ;
	    RECT 1240.2001 41.7000 1248.6000 42.6000 ;
	    RECT 1240.2001 40.5000 1241.1000 41.7000 ;
	    RECT 1242.3000 40.5000 1243.5000 40.8000 ;
	    RECT 1247.4000 40.5000 1248.6000 40.8000 ;
	    RECT 1249.8000 40.5000 1250.7001 47.7000 ;
	    RECT 1252.2001 41.4000 1253.4000 42.6000 ;
	    RECT 1240.2001 39.3000 1241.4000 40.5000 ;
	    RECT 1242.3000 39.6000 1250.7001 40.5000 ;
	    RECT 1249.5000 39.3000 1250.7001 39.6000 ;
	    RECT 1230.6000 29.4000 1231.8000 30.6000 ;
	    RECT 1216.2001 17.4000 1217.4000 18.6000 ;
	    RECT 1211.4000 14.4000 1212.6000 15.6000 ;
	    RECT 1072.2001 11.4000 1073.4000 12.6000 ;
	    RECT 1194.6000 11.4000 1195.8000 12.6000 ;
	    RECT 1211.5500 6.6000 1212.4501 14.4000 ;
	    RECT 1026.6000 5.4000 1027.8000 5.5500 ;
	    RECT 1029.0000 5.4000 1030.2001 5.5500 ;
	    RECT 1211.4000 5.4000 1212.6000 6.6000 ;
	    RECT 1218.6000 6.3000 1219.8000 26.7000 ;
	    RECT 1221.0000 6.3000 1222.2001 26.7000 ;
	    RECT 1223.4000 9.3000 1224.6000 26.7000 ;
	    RECT 1225.8000 23.4000 1227.0000 24.6000 ;
	    RECT 1225.9501 21.6000 1226.8500 23.4000 ;
	    RECT 1225.8000 20.4000 1227.0000 21.6000 ;
	    RECT 1228.2001 9.3000 1229.4000 26.7000 ;
	    RECT 1230.7500 24.6000 1231.6500 29.4000 ;
	    RECT 1230.6000 23.4000 1231.8000 24.6000 ;
	    RECT 1233.0000 9.3000 1234.2001 26.7000 ;
	    RECT 1235.4000 6.3000 1236.6000 26.7000 ;
	    RECT 1237.8000 6.3000 1239.0000 26.7000 ;
	    RECT 1240.2001 6.3000 1241.4000 26.7000 ;
	    RECT 1271.5500 24.6000 1272.4501 95.4000 ;
	    RECT 1271.4000 23.4000 1272.6000 24.6000 ;
	    RECT 1278.7500 21.6000 1279.6500 104.4000 ;
	    RECT 1285.9501 102.6000 1286.8500 185.4000 ;
	    RECT 1288.3500 162.6000 1289.2500 200.4000 ;
	    RECT 1295.5500 198.6000 1296.4501 233.4000 ;
	    RECT 1295.4000 197.4000 1296.6000 198.6000 ;
	    RECT 1288.2001 161.4000 1289.4000 162.6000 ;
	    RECT 1285.8000 101.4000 1287.0000 102.6000 ;
	    RECT 1283.4000 83.4000 1284.6000 84.6000 ;
	    RECT 1283.5500 78.6000 1284.4501 83.4000 ;
	    RECT 1288.3500 81.6000 1289.2500 161.4000 ;
	    RECT 1297.9501 132.6000 1298.8500 347.4000 ;
	    RECT 1300.2001 323.4000 1301.4000 324.6000 ;
	    RECT 1300.3500 285.6000 1301.2500 323.4000 ;
	    RECT 1305.0000 317.4000 1306.2001 318.6000 ;
	    RECT 1300.2001 284.4000 1301.4000 285.6000 ;
	    RECT 1300.2001 257.4000 1301.4000 258.6000 ;
	    RECT 1305.0000 233.4000 1306.2001 234.6000 ;
	    RECT 1305.1500 228.6000 1306.0500 233.4000 ;
	    RECT 1305.0000 227.4000 1306.2001 228.6000 ;
	    RECT 1307.5500 222.6000 1308.4501 725.4000 ;
	    RECT 1309.8000 704.4000 1311.0000 705.6000 ;
	    RECT 1309.9501 702.6000 1310.8500 704.4000 ;
	    RECT 1309.8000 701.4000 1311.0000 702.6000 ;
	    RECT 1309.8000 690.4500 1311.0000 690.6000 ;
	    RECT 1312.3500 690.4500 1313.2500 740.4000 ;
	    RECT 1326.6000 737.4000 1327.8000 738.6000 ;
	    RECT 1331.4000 737.4000 1332.6000 738.6000 ;
	    RECT 1317.0000 734.4000 1318.2001 735.6000 ;
	    RECT 1317.1500 708.6000 1318.0500 734.4000 ;
	    RECT 1317.0000 707.4000 1318.2001 708.6000 ;
	    RECT 1309.8000 689.5500 1313.2500 690.4500 ;
	    RECT 1309.8000 689.4000 1311.0000 689.5500 ;
	    RECT 1309.9501 681.6000 1310.8500 689.4000 ;
	    RECT 1309.8000 680.4000 1311.0000 681.6000 ;
	    RECT 1326.7500 678.6000 1327.6500 737.4000 ;
	    RECT 1331.5500 732.6000 1332.4501 737.4000 ;
	    RECT 1331.4000 731.4000 1332.6000 732.6000 ;
	    RECT 1331.5500 681.6000 1332.4501 731.4000 ;
	    RECT 1333.9501 708.6000 1334.8500 740.4000 ;
	    RECT 1350.6000 734.4000 1351.8000 735.6000 ;
	    RECT 1350.7500 714.6000 1351.6500 734.4000 ;
	    RECT 1350.6000 713.4000 1351.8000 714.6000 ;
	    RECT 1333.8000 707.4000 1335.0000 708.6000 ;
	    RECT 1345.8000 701.4000 1347.0000 702.6000 ;
	    RECT 1345.9501 681.6000 1346.8500 701.4000 ;
	    RECT 1331.4000 680.4000 1332.6000 681.6000 ;
	    RECT 1345.8000 680.4000 1347.0000 681.6000 ;
	    RECT 1326.6000 677.4000 1327.8000 678.6000 ;
	    RECT 1331.4000 674.4000 1332.6000 675.6000 ;
	    RECT 1331.5500 666.6000 1332.4501 674.4000 ;
	    RECT 1326.6000 665.4000 1327.8000 666.6000 ;
	    RECT 1331.4000 665.4000 1332.6000 666.6000 ;
	    RECT 1319.4000 647.4000 1320.6000 648.6000 ;
	    RECT 1314.6000 641.4000 1315.8000 642.6000 ;
	    RECT 1312.2001 617.4000 1313.4000 618.6000 ;
	    RECT 1312.3500 594.6000 1313.2500 617.4000 ;
	    RECT 1314.7500 612.6000 1315.6500 641.4000 ;
	    RECT 1319.5500 639.6000 1320.4501 647.4000 ;
	    RECT 1319.4000 638.4000 1320.6000 639.6000 ;
	    RECT 1314.6000 611.4000 1315.8000 612.6000 ;
	    RECT 1312.2001 593.4000 1313.4000 594.6000 ;
	    RECT 1312.2001 590.4000 1313.4000 591.6000 ;
	    RECT 1312.3500 582.6000 1313.2500 590.4000 ;
	    RECT 1312.2001 581.4000 1313.4000 582.6000 ;
	    RECT 1314.6000 560.4000 1315.8000 561.6000 ;
	    RECT 1314.7500 534.6000 1315.6500 560.4000 ;
	    RECT 1326.7500 540.6000 1327.6500 665.4000 ;
	    RECT 1338.6000 650.4000 1339.8000 651.6000 ;
	    RECT 1338.7500 630.6000 1339.6500 650.4000 ;
	    RECT 1345.9501 642.6000 1346.8500 680.4000 ;
	    RECT 1350.7500 678.6000 1351.6500 713.4000 ;
	    RECT 1365.1500 684.6000 1366.0500 857.4000 ;
	    RECT 1365.0000 683.4000 1366.2001 684.6000 ;
	    RECT 1367.5500 678.6000 1368.4501 917.4000 ;
	    RECT 1374.6000 888.4500 1375.8000 888.6000 ;
	    RECT 1377.1500 888.4500 1378.0500 920.4000 ;
	    RECT 1408.2001 917.4000 1409.4000 918.6000 ;
	    RECT 1410.7500 912.6000 1411.6500 947.4000 ;
	    RECT 1413.1500 924.6000 1414.0500 974.4000 ;
	    RECT 1413.0000 923.4000 1414.2001 924.6000 ;
	    RECT 1413.1500 921.6000 1414.0500 923.4000 ;
	    RECT 1417.9501 921.6000 1418.8500 1073.4000 ;
	    RECT 1427.5500 1068.6000 1428.4501 1118.4000 ;
	    RECT 1429.8000 1115.4000 1431.0000 1116.6000 ;
	    RECT 1429.9501 1110.6000 1430.8500 1115.4000 ;
	    RECT 1429.8000 1109.4000 1431.0000 1110.6000 ;
	    RECT 1441.8000 1103.4000 1443.0000 1104.6000 ;
	    RECT 1441.9501 1101.6000 1442.8500 1103.4000 ;
	    RECT 1444.3500 1101.6000 1445.2500 1133.4000 ;
	    RECT 1429.8000 1100.4000 1431.0000 1101.6000 ;
	    RECT 1432.2001 1100.4000 1433.4000 1101.6000 ;
	    RECT 1441.8000 1100.4000 1443.0000 1101.6000 ;
	    RECT 1444.2001 1100.4000 1445.4000 1101.6000 ;
	    RECT 1429.9501 1092.6000 1430.8500 1100.4000 ;
	    RECT 1429.8000 1091.4000 1431.0000 1092.6000 ;
	    RECT 1427.4000 1067.4000 1428.6000 1068.6000 ;
	    RECT 1427.5500 1032.6000 1428.4501 1067.4000 ;
	    RECT 1432.3500 1062.6000 1433.2500 1100.4000 ;
	    RECT 1439.4000 1097.4000 1440.6000 1098.6000 ;
	    RECT 1434.6000 1094.4000 1435.8000 1095.6000 ;
	    RECT 1432.2001 1061.4000 1433.4000 1062.6000 ;
	    RECT 1429.8000 1040.4000 1431.0000 1041.6000 ;
	    RECT 1427.4000 1031.4000 1428.6000 1032.6000 ;
	    RECT 1425.0000 1013.4000 1426.2001 1014.6000 ;
	    RECT 1425.1500 1005.6000 1426.0500 1013.4000 ;
	    RECT 1425.0000 1004.4000 1426.2001 1005.6000 ;
	    RECT 1429.9501 1002.6000 1430.8500 1040.4000 ;
	    RECT 1432.2001 1007.4000 1433.4000 1008.6000 ;
	    RECT 1432.3500 1005.6000 1433.2500 1007.4000 ;
	    RECT 1432.2001 1004.4000 1433.4000 1005.6000 ;
	    RECT 1429.8000 1001.4000 1431.0000 1002.6000 ;
	    RECT 1434.7500 978.6000 1435.6500 1094.4000 ;
	    RECT 1439.5500 1092.6000 1440.4501 1097.4000 ;
	    RECT 1439.4000 1091.4000 1440.6000 1092.6000 ;
	    RECT 1444.2001 1001.4000 1445.4000 1002.6000 ;
	    RECT 1437.0000 980.4000 1438.2001 981.6000 ;
	    RECT 1434.6000 977.4000 1435.8000 978.6000 ;
	    RECT 1432.2001 950.4000 1433.4000 951.6000 ;
	    RECT 1429.8000 935.4000 1431.0000 936.6000 ;
	    RECT 1429.9501 924.6000 1430.8500 935.4000 ;
	    RECT 1429.8000 923.4000 1431.0000 924.6000 ;
	    RECT 1432.3500 921.6000 1433.2500 950.4000 ;
	    RECT 1413.0000 920.4000 1414.2001 921.6000 ;
	    RECT 1417.8000 920.4000 1419.0000 921.6000 ;
	    RECT 1432.2001 920.4000 1433.4000 921.6000 ;
	    RECT 1410.6000 911.4000 1411.8000 912.6000 ;
	    RECT 1374.6000 887.5500 1378.0500 888.4500 ;
	    RECT 1374.6000 887.4000 1375.8000 887.5500 ;
	    RECT 1415.4000 884.4000 1416.6000 885.6000 ;
	    RECT 1379.4000 869.4000 1380.6000 870.6000 ;
	    RECT 1377.0000 863.4000 1378.2001 864.6000 ;
	    RECT 1377.1500 861.6000 1378.0500 863.4000 ;
	    RECT 1377.0000 860.4000 1378.2001 861.6000 ;
	    RECT 1372.2001 857.4000 1373.4000 858.6000 ;
	    RECT 1377.0000 857.4000 1378.2001 858.6000 ;
	    RECT 1372.3500 855.6000 1373.2500 857.4000 ;
	    RECT 1372.2001 854.4000 1373.4000 855.6000 ;
	    RECT 1374.6000 836.4000 1375.8000 837.6000 ;
	    RECT 1374.7500 828.6000 1375.6500 836.4000 ;
	    RECT 1374.6000 827.4000 1375.8000 828.6000 ;
	    RECT 1377.1500 801.6000 1378.0500 857.4000 ;
	    RECT 1379.5500 825.6000 1380.4501 869.4000 ;
	    RECT 1379.4000 824.4000 1380.6000 825.6000 ;
	    RECT 1377.0000 800.4000 1378.2001 801.6000 ;
	    RECT 1374.6000 764.4000 1375.8000 765.6000 ;
	    RECT 1374.7500 738.6000 1375.6500 764.4000 ;
	    RECT 1369.8000 737.4000 1371.0000 738.6000 ;
	    RECT 1374.6000 737.4000 1375.8000 738.6000 ;
	    RECT 1369.9501 732.6000 1370.8500 737.4000 ;
	    RECT 1369.8000 731.4000 1371.0000 732.6000 ;
	    RECT 1369.9501 702.6000 1370.8500 731.4000 ;
	    RECT 1369.8000 701.4000 1371.0000 702.6000 ;
	    RECT 1369.8000 698.4000 1371.0000 699.6000 ;
	    RECT 1350.6000 677.4000 1351.8000 678.6000 ;
	    RECT 1367.4000 678.4500 1368.6000 678.6000 ;
	    RECT 1365.1500 677.5500 1368.6000 678.4500 ;
	    RECT 1348.2001 647.4000 1349.4000 648.6000 ;
	    RECT 1345.8000 641.4000 1347.0000 642.6000 ;
	    RECT 1338.6000 629.4000 1339.8000 630.6000 ;
	    RECT 1345.8000 629.4000 1347.0000 630.6000 ;
	    RECT 1336.2001 617.4000 1337.4000 618.6000 ;
	    RECT 1336.3500 594.6000 1337.2500 617.4000 ;
	    RECT 1338.7500 615.6000 1339.6500 629.4000 ;
	    RECT 1341.0000 623.4000 1342.2001 624.6000 ;
	    RECT 1345.9501 621.6000 1346.8500 629.4000 ;
	    RECT 1345.8000 620.4000 1347.0000 621.6000 ;
	    RECT 1348.3500 618.6000 1349.2500 647.4000 ;
	    RECT 1350.6000 644.4000 1351.8000 645.6000 ;
	    RECT 1350.7500 636.6000 1351.6500 644.4000 ;
	    RECT 1350.6000 635.4000 1351.8000 636.6000 ;
	    RECT 1341.0000 617.4000 1342.2001 618.6000 ;
	    RECT 1348.2001 617.4000 1349.4000 618.6000 ;
	    RECT 1338.6000 614.4000 1339.8000 615.6000 ;
	    RECT 1336.2001 593.4000 1337.4000 594.6000 ;
	    RECT 1336.2001 591.4500 1337.4000 591.6000 ;
	    RECT 1336.2001 590.5500 1339.6500 591.4500 ;
	    RECT 1336.2001 590.4000 1337.4000 590.5500 ;
	    RECT 1329.0000 587.4000 1330.2001 588.6000 ;
	    RECT 1331.4000 587.4000 1332.6000 588.6000 ;
	    RECT 1336.2001 587.4000 1337.4000 588.6000 ;
	    RECT 1329.1500 582.6000 1330.0500 587.4000 ;
	    RECT 1329.0000 581.4000 1330.2001 582.6000 ;
	    RECT 1331.5500 570.6000 1332.4501 587.4000 ;
	    RECT 1333.8000 584.4000 1335.0000 585.6000 ;
	    RECT 1333.9501 576.6000 1334.8500 584.4000 ;
	    RECT 1333.8000 575.4000 1335.0000 576.6000 ;
	    RECT 1331.4000 569.4000 1332.6000 570.6000 ;
	    RECT 1326.6000 539.4000 1327.8000 540.6000 ;
	    RECT 1333.8000 539.4000 1335.0000 540.6000 ;
	    RECT 1314.6000 533.4000 1315.8000 534.6000 ;
	    RECT 1331.4000 533.4000 1332.6000 534.6000 ;
	    RECT 1317.0000 527.4000 1318.2001 528.6000 ;
	    RECT 1319.4000 527.4000 1320.6000 528.6000 ;
	    RECT 1314.6000 524.4000 1315.8000 525.6000 ;
	    RECT 1312.2001 521.4000 1313.4000 522.6000 ;
	    RECT 1312.3500 486.6000 1313.2500 521.4000 ;
	    RECT 1314.7500 516.6000 1315.6500 524.4000 ;
	    RECT 1314.6000 515.4000 1315.8000 516.6000 ;
	    RECT 1317.1500 501.6000 1318.0500 527.4000 ;
	    RECT 1319.5500 522.6000 1320.4501 527.4000 ;
	    RECT 1319.4000 521.4000 1320.6000 522.6000 ;
	    RECT 1319.5500 504.6000 1320.4501 521.4000 ;
	    RECT 1331.5500 519.6000 1332.4501 533.4000 ;
	    RECT 1333.9501 522.6000 1334.8500 539.4000 ;
	    RECT 1336.3500 534.6000 1337.2500 587.4000 ;
	    RECT 1338.7500 576.6000 1339.6500 590.5500 ;
	    RECT 1338.6000 575.4000 1339.8000 576.6000 ;
	    RECT 1336.2001 533.4000 1337.4000 534.6000 ;
	    RECT 1341.1500 522.6000 1342.0500 617.4000 ;
	    RECT 1350.7500 612.6000 1351.6500 635.4000 ;
	    RECT 1343.4000 611.4000 1344.6000 612.6000 ;
	    RECT 1350.6000 611.4000 1351.8000 612.6000 ;
	    RECT 1343.5500 588.6000 1344.4501 611.4000 ;
	    RECT 1343.4000 587.4000 1344.6000 588.6000 ;
	    RECT 1348.2001 587.4000 1349.4000 588.6000 ;
	    RECT 1343.5500 555.6000 1344.4501 587.4000 ;
	    RECT 1348.3500 570.6000 1349.2500 587.4000 ;
	    RECT 1348.2001 569.4000 1349.4000 570.6000 ;
	    RECT 1348.2001 563.4000 1349.4000 564.6000 ;
	    RECT 1355.4000 563.4000 1356.6000 564.6000 ;
	    RECT 1362.6000 563.4000 1363.8000 564.6000 ;
	    RECT 1348.3500 561.6000 1349.2500 563.4000 ;
	    RECT 1348.2001 560.4000 1349.4000 561.6000 ;
	    RECT 1350.6000 560.4000 1351.8000 561.6000 ;
	    RECT 1345.8000 557.4000 1347.0000 558.6000 ;
	    RECT 1343.4000 554.4000 1344.6000 555.6000 ;
	    RECT 1333.8000 521.4000 1335.0000 522.6000 ;
	    RECT 1341.0000 521.4000 1342.2001 522.6000 ;
	    RECT 1331.4000 518.4000 1332.6000 519.6000 ;
	    RECT 1324.2001 515.4000 1325.4000 516.6000 ;
	    RECT 1324.3500 504.6000 1325.2500 515.4000 ;
	    RECT 1319.4000 503.4000 1320.6000 504.6000 ;
	    RECT 1324.2001 503.4000 1325.4000 504.6000 ;
	    RECT 1317.0000 500.4000 1318.2001 501.6000 ;
	    RECT 1319.4000 500.4000 1320.6000 501.6000 ;
	    RECT 1314.6000 494.4000 1315.8000 495.6000 ;
	    RECT 1312.2001 485.4000 1313.4000 486.6000 ;
	    RECT 1314.7500 468.6000 1315.6500 494.4000 ;
	    RECT 1319.5500 492.6000 1320.4501 500.4000 ;
	    RECT 1326.6000 497.4000 1327.8000 498.6000 ;
	    RECT 1319.4000 491.4000 1320.6000 492.6000 ;
	    RECT 1319.5500 471.6000 1320.4501 491.4000 ;
	    RECT 1319.4000 470.4000 1320.6000 471.6000 ;
	    RECT 1312.2001 467.4000 1313.4000 468.6000 ;
	    RECT 1314.6000 467.4000 1315.8000 468.6000 ;
	    RECT 1321.8000 434.4000 1323.0000 435.6000 ;
	    RECT 1312.2001 413.4000 1313.4000 414.6000 ;
	    RECT 1312.3500 369.6000 1313.2500 413.4000 ;
	    RECT 1314.6000 401.4000 1315.8000 402.6000 ;
	    RECT 1319.4000 401.4000 1320.6000 402.6000 ;
	    RECT 1314.7500 387.6000 1315.6500 401.4000 ;
	    RECT 1317.0000 398.4000 1318.2001 399.6000 ;
	    RECT 1317.1500 396.6000 1318.0500 398.4000 ;
	    RECT 1317.0000 395.4000 1318.2001 396.6000 ;
	    RECT 1314.6000 386.4000 1315.8000 387.6000 ;
	    RECT 1317.0000 383.4000 1318.2001 384.6000 ;
	    RECT 1317.1500 381.6000 1318.0500 383.4000 ;
	    RECT 1317.0000 380.4000 1318.2001 381.6000 ;
	    RECT 1312.2001 368.4000 1313.4000 369.6000 ;
	    RECT 1319.5500 366.6000 1320.4501 401.4000 ;
	    RECT 1321.9501 372.4500 1322.8500 434.4000 ;
	    RECT 1326.7500 426.6000 1327.6500 497.4000 ;
	    RECT 1329.0000 467.4000 1330.2001 468.6000 ;
	    RECT 1329.1500 444.6000 1330.0500 467.4000 ;
	    RECT 1329.0000 443.4000 1330.2001 444.6000 ;
	    RECT 1329.1500 441.6000 1330.0500 443.4000 ;
	    RECT 1329.0000 440.4000 1330.2001 441.6000 ;
	    RECT 1329.0000 438.4500 1330.2001 438.6000 ;
	    RECT 1331.5500 438.4500 1332.4501 518.4000 ;
	    RECT 1338.6000 485.4000 1339.8000 486.6000 ;
	    RECT 1336.2001 479.4000 1337.4000 480.6000 ;
	    RECT 1336.3500 468.6000 1337.2500 479.4000 ;
	    RECT 1336.2001 467.4000 1337.4000 468.6000 ;
	    RECT 1336.3500 465.6000 1337.2500 467.4000 ;
	    RECT 1336.2001 464.4000 1337.4000 465.6000 ;
	    RECT 1336.2001 440.4000 1337.4000 441.6000 ;
	    RECT 1336.3500 438.6000 1337.2500 440.4000 ;
	    RECT 1338.7500 438.6000 1339.6500 485.4000 ;
	    RECT 1329.0000 437.5500 1332.4501 438.4500 ;
	    RECT 1329.0000 437.4000 1330.2001 437.5500 ;
	    RECT 1333.8000 437.4000 1335.0000 438.6000 ;
	    RECT 1336.2001 437.4000 1337.4000 438.6000 ;
	    RECT 1338.6000 437.4000 1339.8000 438.6000 ;
	    RECT 1326.6000 425.4000 1327.8000 426.6000 ;
	    RECT 1324.2001 419.4000 1325.4000 420.6000 ;
	    RECT 1329.0000 419.4000 1330.2001 420.6000 ;
	    RECT 1324.3500 375.6000 1325.2500 419.4000 ;
	    RECT 1333.9501 402.6000 1334.8500 437.4000 ;
	    RECT 1341.1500 408.6000 1342.0500 521.4000 ;
	    RECT 1345.9501 516.6000 1346.8500 557.4000 ;
	    RECT 1348.2001 551.4000 1349.4000 552.6000 ;
	    RECT 1345.8000 515.4000 1347.0000 516.6000 ;
	    RECT 1345.9501 495.6000 1346.8500 515.4000 ;
	    RECT 1345.8000 494.4000 1347.0000 495.6000 ;
	    RECT 1348.3500 468.6000 1349.2500 551.4000 ;
	    RECT 1350.7500 534.6000 1351.6500 560.4000 ;
	    RECT 1362.7500 546.6000 1363.6500 563.4000 ;
	    RECT 1362.6000 545.4000 1363.8000 546.6000 ;
	    RECT 1350.6000 533.4000 1351.8000 534.6000 ;
	    RECT 1350.7500 528.6000 1351.6500 533.4000 ;
	    RECT 1350.6000 527.4000 1351.8000 528.6000 ;
	    RECT 1355.4000 503.4000 1356.6000 504.6000 ;
	    RECT 1353.0000 497.4000 1354.2001 498.6000 ;
	    RECT 1350.6000 491.4000 1351.8000 492.6000 ;
	    RECT 1353.1500 480.6000 1354.0500 497.4000 ;
	    RECT 1355.5500 495.6000 1356.4501 503.4000 ;
	    RECT 1355.4000 494.4000 1356.6000 495.6000 ;
	    RECT 1353.0000 479.4000 1354.2001 480.6000 ;
	    RECT 1348.2001 467.4000 1349.4000 468.6000 ;
	    RECT 1345.8000 443.4000 1347.0000 444.6000 ;
	    RECT 1345.9501 441.6000 1346.8500 443.4000 ;
	    RECT 1345.8000 440.4000 1347.0000 441.6000 ;
	    RECT 1343.4000 437.4000 1344.6000 438.6000 ;
	    RECT 1341.0000 407.4000 1342.2001 408.6000 ;
	    RECT 1333.8000 401.4000 1335.0000 402.6000 ;
	    RECT 1326.6000 389.4000 1327.8000 390.6000 ;
	    RECT 1324.2001 374.4000 1325.4000 375.6000 ;
	    RECT 1326.7500 372.6000 1327.6500 389.4000 ;
	    RECT 1329.0000 383.4000 1330.2001 384.6000 ;
	    RECT 1329.1500 378.6000 1330.0500 383.4000 ;
	    RECT 1329.0000 377.4000 1330.2001 378.6000 ;
	    RECT 1321.9501 371.5500 1325.2500 372.4500 ;
	    RECT 1319.4000 365.4000 1320.6000 366.6000 ;
	    RECT 1321.8000 347.4000 1323.0000 348.6000 ;
	    RECT 1309.8000 341.4000 1311.0000 342.6000 ;
	    RECT 1314.6000 341.4000 1315.8000 342.6000 ;
	    RECT 1309.9501 330.6000 1310.8500 341.4000 ;
	    RECT 1309.8000 329.4000 1311.0000 330.6000 ;
	    RECT 1309.8000 314.4000 1311.0000 315.6000 ;
	    RECT 1309.9501 312.6000 1310.8500 314.4000 ;
	    RECT 1309.8000 311.4000 1311.0000 312.6000 ;
	    RECT 1309.9501 276.6000 1310.8500 311.4000 ;
	    RECT 1309.8000 275.4000 1311.0000 276.6000 ;
	    RECT 1309.9501 258.6000 1310.8500 275.4000 ;
	    RECT 1309.8000 257.4000 1311.0000 258.6000 ;
	    RECT 1300.2001 221.4000 1301.4000 222.6000 ;
	    RECT 1307.4000 221.4000 1308.6000 222.6000 ;
	    RECT 1312.2001 218.4000 1313.4000 219.6000 ;
	    RECT 1312.3500 216.6000 1313.2500 218.4000 ;
	    RECT 1312.2001 215.4000 1313.4000 216.6000 ;
	    RECT 1302.6000 209.4000 1303.8000 210.6000 ;
	    RECT 1302.7500 195.6000 1303.6500 209.4000 ;
	    RECT 1312.2001 200.4000 1313.4000 201.6000 ;
	    RECT 1312.3500 198.6000 1313.2500 200.4000 ;
	    RECT 1312.2001 197.4000 1313.4000 198.6000 ;
	    RECT 1302.6000 194.4000 1303.8000 195.6000 ;
	    RECT 1309.8000 192.4500 1311.0000 192.6000 ;
	    RECT 1312.3500 192.4500 1313.2500 197.4000 ;
	    RECT 1309.8000 191.5500 1313.2500 192.4500 ;
	    RECT 1309.8000 191.4000 1311.0000 191.5500 ;
	    RECT 1307.4000 149.4000 1308.6000 150.6000 ;
	    RECT 1307.5500 141.6000 1308.4501 149.4000 ;
	    RECT 1305.0000 140.4000 1306.2001 141.6000 ;
	    RECT 1307.4000 140.4000 1308.6000 141.6000 ;
	    RECT 1297.8000 131.4000 1299.0000 132.6000 ;
	    RECT 1305.1500 126.6000 1306.0500 140.4000 ;
	    RECT 1309.8000 137.4000 1311.0000 138.6000 ;
	    RECT 1309.9501 132.6000 1310.8500 137.4000 ;
	    RECT 1309.8000 131.4000 1311.0000 132.6000 ;
	    RECT 1305.0000 125.4000 1306.2001 126.6000 ;
	    RECT 1309.9501 114.6000 1310.8500 131.4000 ;
	    RECT 1309.8000 113.4000 1311.0000 114.6000 ;
	    RECT 1307.4000 101.4000 1308.6000 102.6000 ;
	    RECT 1307.5500 96.6000 1308.4501 101.4000 ;
	    RECT 1307.4000 95.4000 1308.6000 96.6000 ;
	    RECT 1314.7500 81.6000 1315.6500 341.4000 ;
	    RECT 1319.4000 329.4000 1320.6000 330.6000 ;
	    RECT 1319.5500 321.6000 1320.4501 329.4000 ;
	    RECT 1319.4000 320.4000 1320.6000 321.6000 ;
	    RECT 1321.9501 270.6000 1322.8500 347.4000 ;
	    RECT 1324.3500 342.6000 1325.2500 371.5500 ;
	    RECT 1326.6000 371.4000 1327.8000 372.6000 ;
	    RECT 1331.4000 366.3000 1332.6000 386.7000 ;
	    RECT 1333.8000 366.3000 1335.0000 386.7000 ;
	    RECT 1336.2001 369.3000 1337.4000 386.7000 ;
	    RECT 1338.6000 380.4000 1339.8000 381.6000 ;
	    RECT 1338.7500 360.6000 1339.6500 380.4000 ;
	    RECT 1341.0000 369.3000 1342.2001 386.7000 ;
	    RECT 1343.5500 384.6000 1344.4501 437.4000 ;
	    RECT 1345.8000 419.4000 1347.0000 420.6000 ;
	    RECT 1360.2001 419.4000 1361.4000 420.6000 ;
	    RECT 1345.9501 405.6000 1346.8500 419.4000 ;
	    RECT 1357.8000 413.4000 1359.0000 414.6000 ;
	    RECT 1350.6000 407.4000 1351.8000 408.6000 ;
	    RECT 1345.8000 404.4000 1347.0000 405.6000 ;
	    RECT 1357.9501 402.6000 1358.8500 413.4000 ;
	    RECT 1360.3500 408.6000 1361.2500 419.4000 ;
	    RECT 1360.2001 407.4000 1361.4000 408.6000 ;
	    RECT 1350.6000 401.4000 1351.8000 402.6000 ;
	    RECT 1357.8000 401.4000 1359.0000 402.6000 ;
	    RECT 1343.4000 383.4000 1344.6000 384.6000 ;
	    RECT 1345.8000 369.3000 1347.0000 386.7000 ;
	    RECT 1348.2001 366.3000 1349.4000 386.7000 ;
	    RECT 1350.6000 366.3000 1351.8000 386.7000 ;
	    RECT 1353.0000 366.3000 1354.2001 386.7000 ;
	    RECT 1365.1500 372.4500 1366.0500 677.5500 ;
	    RECT 1367.4000 677.4000 1368.6000 677.5500 ;
	    RECT 1369.9501 675.6000 1370.8500 698.4000 ;
	    RECT 1369.8000 674.4000 1371.0000 675.6000 ;
	    RECT 1369.8000 641.4000 1371.0000 642.6000 ;
	    RECT 1367.4000 617.4000 1368.6000 618.6000 ;
	    RECT 1367.5500 540.6000 1368.4501 617.4000 ;
	    RECT 1369.9501 615.6000 1370.8500 641.4000 ;
	    RECT 1369.8000 614.4000 1371.0000 615.6000 ;
	    RECT 1369.9501 552.6000 1370.8500 614.4000 ;
	    RECT 1374.7500 612.6000 1375.6500 737.4000 ;
	    RECT 1377.0000 641.4000 1378.2001 642.6000 ;
	    RECT 1374.6000 611.4000 1375.8000 612.6000 ;
	    RECT 1377.1500 591.6000 1378.0500 641.4000 ;
	    RECT 1377.0000 590.4000 1378.2001 591.6000 ;
	    RECT 1374.6000 584.4000 1375.8000 585.6000 ;
	    RECT 1374.7500 576.6000 1375.6500 584.4000 ;
	    RECT 1374.6000 575.4000 1375.8000 576.6000 ;
	    RECT 1379.5500 555.4500 1380.4501 824.4000 ;
	    RECT 1381.8000 816.3000 1383.0000 836.7000 ;
	    RECT 1384.2001 816.3000 1385.4000 836.7000 ;
	    RECT 1386.6000 816.3000 1387.8000 833.7000 ;
	    RECT 1389.0000 821.4000 1390.2001 822.6000 ;
	    RECT 1389.1500 810.6000 1390.0500 821.4000 ;
	    RECT 1391.4000 816.3000 1392.6000 833.7000 ;
	    RECT 1393.8000 821.4000 1395.0000 822.6000 ;
	    RECT 1393.9501 819.6000 1394.8500 821.4000 ;
	    RECT 1393.8000 818.4000 1395.0000 819.6000 ;
	    RECT 1389.0000 809.4000 1390.2001 810.6000 ;
	    RECT 1393.9501 762.6000 1394.8500 818.4000 ;
	    RECT 1396.2001 816.3000 1397.4000 833.7000 ;
	    RECT 1398.6000 816.3000 1399.8000 836.7000 ;
	    RECT 1401.0000 816.3000 1402.2001 836.7000 ;
	    RECT 1403.4000 816.3000 1404.6000 836.7000 ;
	    RECT 1401.3000 803.4000 1402.5000 803.7000 ;
	    RECT 1401.3000 802.5000 1409.7001 803.4000 ;
	    RECT 1410.6000 802.5000 1411.8000 803.7000 ;
	    RECT 1401.3000 795.3000 1402.2001 802.5000 ;
	    RECT 1403.4000 802.2000 1404.6000 802.5000 ;
	    RECT 1408.5000 802.2000 1409.7001 802.5000 ;
	    RECT 1410.9000 801.3000 1411.8000 802.5000 ;
	    RECT 1415.5500 801.6000 1416.4501 884.4000 ;
	    RECT 1417.9501 858.6000 1418.8500 920.4000 ;
	    RECT 1427.4000 911.4000 1428.6000 912.6000 ;
	    RECT 1417.8000 857.4000 1419.0000 858.6000 ;
	    RECT 1425.0000 857.4000 1426.2001 858.6000 ;
	    RECT 1422.6000 830.4000 1423.8000 831.6000 ;
	    RECT 1403.4000 800.4000 1411.8000 801.3000 ;
	    RECT 1413.0000 800.4000 1414.2001 801.6000 ;
	    RECT 1415.4000 800.4000 1416.6000 801.6000 ;
	    RECT 1417.8000 800.4000 1419.0000 801.6000 ;
	    RECT 1403.4000 798.3000 1404.3000 800.4000 ;
	    RECT 1403.1000 797.1000 1404.3000 798.3000 ;
	    RECT 1405.8000 797.4000 1407.0000 798.6000 ;
	    RECT 1410.9000 795.3000 1411.8000 800.4000 ;
	    RECT 1401.3000 794.1000 1402.5000 795.3000 ;
	    RECT 1410.6000 794.1000 1411.8000 795.3000 ;
	    RECT 1405.8000 791.4000 1407.0000 792.6000 ;
	    RECT 1393.8000 761.4000 1395.0000 762.6000 ;
	    RECT 1386.6000 743.4000 1387.8000 744.6000 ;
	    RECT 1386.7500 738.6000 1387.6500 743.4000 ;
	    RECT 1401.0000 740.4000 1402.2001 741.6000 ;
	    RECT 1386.6000 737.4000 1387.8000 738.6000 ;
	    RECT 1386.6000 707.4000 1387.8000 708.6000 ;
	    RECT 1389.3000 707.7000 1390.5000 708.9000 ;
	    RECT 1384.2001 699.4500 1385.4000 699.6000 ;
	    RECT 1386.7500 699.4500 1387.6500 707.4000 ;
	    RECT 1384.2001 698.5500 1387.6500 699.4500 ;
	    RECT 1389.3000 700.5000 1390.2001 707.7000 ;
	    RECT 1393.8000 707.4000 1395.0000 708.6000 ;
	    RECT 1398.6000 707.7000 1399.8000 708.9000 ;
	    RECT 1391.1000 704.7000 1392.3000 705.9000 ;
	    RECT 1393.9501 705.6000 1394.8500 707.4000 ;
	    RECT 1391.4000 702.6000 1392.3000 704.7000 ;
	    RECT 1393.8000 704.4000 1395.0000 705.6000 ;
	    RECT 1398.9000 702.6000 1399.8000 707.7000 ;
	    RECT 1401.1500 702.6000 1402.0500 740.4000 ;
	    RECT 1405.9501 735.6000 1406.8500 791.4000 ;
	    RECT 1408.2001 785.4000 1409.4000 786.6000 ;
	    RECT 1405.8000 734.4000 1407.0000 735.6000 ;
	    RECT 1391.4000 701.7000 1399.8000 702.6000 ;
	    RECT 1391.4000 700.5000 1392.6000 700.8000 ;
	    RECT 1396.5000 700.5000 1397.7001 700.8000 ;
	    RECT 1398.9000 700.5000 1399.8000 701.7000 ;
	    RECT 1401.0000 701.4000 1402.2001 702.6000 ;
	    RECT 1389.3000 699.6000 1397.7001 700.5000 ;
	    RECT 1389.3000 699.3000 1390.5000 699.6000 ;
	    RECT 1398.6000 699.3000 1399.8000 700.5000 ;
	    RECT 1384.2001 698.4000 1385.4000 698.5500 ;
	    RECT 1386.6000 680.4000 1387.8000 681.6000 ;
	    RECT 1405.8000 680.4000 1407.0000 681.6000 ;
	    RECT 1386.7500 678.6000 1387.6500 680.4000 ;
	    RECT 1386.6000 677.4000 1387.8000 678.6000 ;
	    RECT 1405.9501 672.6000 1406.8500 680.4000 ;
	    RECT 1405.8000 671.4000 1407.0000 672.6000 ;
	    RECT 1391.4000 647.4000 1392.6000 648.6000 ;
	    RECT 1401.0000 647.4000 1402.2001 648.6000 ;
	    RECT 1381.8000 644.4000 1383.0000 645.6000 ;
	    RECT 1398.6000 644.4000 1399.8000 645.6000 ;
	    RECT 1381.9501 618.6000 1382.8500 644.4000 ;
	    RECT 1398.7500 642.6000 1399.6500 644.4000 ;
	    RECT 1401.1500 642.6000 1402.0500 647.4000 ;
	    RECT 1403.4000 644.4000 1404.6000 645.6000 ;
	    RECT 1398.6000 641.4000 1399.8000 642.6000 ;
	    RECT 1401.0000 641.4000 1402.2001 642.6000 ;
	    RECT 1386.6000 629.4000 1387.8000 630.6000 ;
	    RECT 1381.8000 617.4000 1383.0000 618.6000 ;
	    RECT 1381.8000 611.4000 1383.0000 612.6000 ;
	    RECT 1384.2001 611.4000 1385.4000 612.6000 ;
	    RECT 1377.1500 554.5500 1380.4501 555.4500 ;
	    RECT 1369.8000 551.4000 1371.0000 552.6000 ;
	    RECT 1369.8000 545.4000 1371.0000 546.6000 ;
	    RECT 1367.4000 539.4000 1368.6000 540.6000 ;
	    RECT 1369.9501 531.6000 1370.8500 545.4000 ;
	    RECT 1372.2001 533.4000 1373.4000 534.6000 ;
	    RECT 1369.8000 530.4000 1371.0000 531.6000 ;
	    RECT 1367.4000 527.4000 1368.6000 528.6000 ;
	    RECT 1372.3500 525.6000 1373.2500 533.4000 ;
	    RECT 1374.6000 527.4000 1375.8000 528.6000 ;
	    RECT 1372.2001 524.4000 1373.4000 525.6000 ;
	    RECT 1374.7500 516.6000 1375.6500 527.4000 ;
	    RECT 1374.6000 515.4000 1375.8000 516.6000 ;
	    RECT 1377.1500 462.6000 1378.0500 554.5500 ;
	    RECT 1379.4000 527.4000 1380.6000 528.6000 ;
	    RECT 1379.4000 479.4000 1380.6000 480.6000 ;
	    RECT 1377.0000 461.4000 1378.2001 462.6000 ;
	    RECT 1367.4000 458.4000 1368.6000 459.6000 ;
	    RECT 1367.5500 444.6000 1368.4501 458.4000 ;
	    RECT 1367.4000 443.4000 1368.6000 444.6000 ;
	    RECT 1367.5500 420.6000 1368.4501 443.4000 ;
	    RECT 1377.0000 440.4000 1378.2001 441.6000 ;
	    RECT 1369.8000 425.4000 1371.0000 426.6000 ;
	    RECT 1367.4000 419.4000 1368.6000 420.6000 ;
	    RECT 1367.4000 404.4000 1368.6000 405.6000 ;
	    RECT 1367.5500 390.6000 1368.4501 404.4000 ;
	    RECT 1367.4000 389.4000 1368.6000 390.6000 ;
	    RECT 1367.4000 372.4500 1368.6000 372.6000 ;
	    RECT 1365.1500 371.5500 1368.6000 372.4500 ;
	    RECT 1338.6000 359.4000 1339.8000 360.6000 ;
	    RECT 1336.2001 353.4000 1337.4000 354.6000 ;
	    RECT 1333.8000 344.4000 1335.0000 345.6000 ;
	    RECT 1333.9501 342.6000 1334.8500 344.4000 ;
	    RECT 1336.3500 342.6000 1337.2500 353.4000 ;
	    RECT 1348.2001 344.4000 1349.4000 345.6000 ;
	    RECT 1324.2001 341.4000 1325.4000 342.6000 ;
	    RECT 1333.8000 341.4000 1335.0000 342.6000 ;
	    RECT 1336.2001 341.4000 1337.4000 342.6000 ;
	    RECT 1343.4000 341.4000 1344.6000 342.6000 ;
	    RECT 1324.2001 320.4000 1325.4000 321.6000 ;
	    RECT 1324.3500 300.6000 1325.2500 320.4000 ;
	    RECT 1333.8000 314.4000 1335.0000 315.6000 ;
	    RECT 1324.2001 299.4000 1325.4000 300.6000 ;
	    RECT 1324.3500 294.6000 1325.2500 299.4000 ;
	    RECT 1324.2001 293.4000 1325.4000 294.6000 ;
	    RECT 1333.9501 291.6000 1334.8500 314.4000 ;
	    RECT 1333.8000 290.4000 1335.0000 291.6000 ;
	    RECT 1324.2001 287.4000 1325.4000 288.6000 ;
	    RECT 1331.4000 287.4000 1332.6000 288.6000 ;
	    RECT 1329.0000 284.4000 1330.2001 285.6000 ;
	    RECT 1329.1500 282.6000 1330.0500 284.4000 ;
	    RECT 1329.0000 281.4000 1330.2001 282.6000 ;
	    RECT 1321.8000 269.4000 1323.0000 270.6000 ;
	    RECT 1329.0000 260.4000 1330.2001 261.6000 ;
	    RECT 1321.8000 257.4000 1323.0000 258.6000 ;
	    RECT 1321.9501 255.6000 1322.8500 257.4000 ;
	    RECT 1321.8000 254.4000 1323.0000 255.6000 ;
	    RECT 1324.2001 254.4000 1325.4000 255.6000 ;
	    RECT 1324.3500 246.6000 1325.2500 254.4000 ;
	    RECT 1329.1500 252.6000 1330.0500 260.4000 ;
	    RECT 1331.5500 258.6000 1332.4501 287.4000 ;
	    RECT 1333.9501 264.6000 1334.8500 290.4000 ;
	    RECT 1343.5500 288.6000 1344.4501 341.4000 ;
	    RECT 1348.3500 330.6000 1349.2500 344.4000 ;
	    RECT 1350.6000 341.4000 1351.8000 342.6000 ;
	    RECT 1348.2001 329.4000 1349.4000 330.6000 ;
	    RECT 1343.4000 287.4000 1344.6000 288.6000 ;
	    RECT 1333.8000 263.4000 1335.0000 264.6000 ;
	    RECT 1333.8000 260.4000 1335.0000 261.6000 ;
	    RECT 1331.4000 257.4000 1332.6000 258.6000 ;
	    RECT 1331.5500 255.6000 1332.4501 257.4000 ;
	    RECT 1331.4000 254.4000 1332.6000 255.6000 ;
	    RECT 1329.0000 251.4000 1330.2001 252.6000 ;
	    RECT 1324.2001 245.4000 1325.4000 246.6000 ;
	    RECT 1329.1500 228.6000 1330.0500 251.4000 ;
	    RECT 1329.0000 227.4000 1330.2001 228.6000 ;
	    RECT 1333.9501 228.4500 1334.8500 260.4000 ;
	    RECT 1341.0000 239.4000 1342.2001 240.6000 ;
	    RECT 1341.1500 228.6000 1342.0500 239.4000 ;
	    RECT 1343.4000 230.4000 1344.6000 231.6000 ;
	    RECT 1331.5500 227.5500 1334.8500 228.4500 ;
	    RECT 1331.5500 144.6000 1332.4501 227.5500 ;
	    RECT 1341.0000 227.4000 1342.2001 228.6000 ;
	    RECT 1341.0000 225.4500 1342.2001 225.6000 ;
	    RECT 1333.9501 224.5500 1342.2001 225.4500 ;
	    RECT 1333.9501 222.6000 1334.8500 224.5500 ;
	    RECT 1341.0000 224.4000 1342.2001 224.5500 ;
	    RECT 1333.8000 221.4000 1335.0000 222.6000 ;
	    RECT 1343.5500 204.6000 1344.4501 230.4000 ;
	    RECT 1348.2001 209.4000 1349.4000 210.6000 ;
	    RECT 1343.4000 203.4000 1344.6000 204.6000 ;
	    RECT 1348.3500 201.6000 1349.2500 209.4000 ;
	    RECT 1348.2001 200.4000 1349.4000 201.6000 ;
	    RECT 1336.2001 191.4000 1337.4000 192.6000 ;
	    RECT 1331.4000 143.4000 1332.6000 144.6000 ;
	    RECT 1331.5500 135.6000 1332.4501 143.4000 ;
	    RECT 1336.3500 141.6000 1337.2500 191.4000 ;
	    RECT 1348.2001 179.4000 1349.4000 180.6000 ;
	    RECT 1343.4000 161.4000 1344.6000 162.6000 ;
	    RECT 1338.6000 149.4000 1339.8000 150.6000 ;
	    RECT 1338.7500 141.6000 1339.6500 149.4000 ;
	    RECT 1336.2001 140.4000 1337.4000 141.6000 ;
	    RECT 1338.6000 140.4000 1339.8000 141.6000 ;
	    RECT 1336.2001 137.4000 1337.4000 138.6000 ;
	    RECT 1331.4000 134.4000 1332.6000 135.6000 ;
	    RECT 1336.3500 132.6000 1337.2500 137.4000 ;
	    RECT 1336.2001 131.4000 1337.4000 132.6000 ;
	    RECT 1329.0000 113.4000 1330.2001 114.6000 ;
	    RECT 1324.2001 107.7000 1325.4000 108.9000 ;
	    RECT 1324.2001 102.6000 1325.1000 107.7000 ;
	    RECT 1329.1500 105.6000 1330.0500 113.4000 ;
	    RECT 1333.5000 107.7000 1334.7001 108.9000 ;
	    RECT 1329.0000 104.4000 1330.2001 105.6000 ;
	    RECT 1331.7001 104.7000 1332.9000 105.9000 ;
	    RECT 1331.7001 102.6000 1332.6000 104.7000 ;
	    RECT 1321.8000 101.4000 1323.0000 102.6000 ;
	    RECT 1324.2001 101.7000 1332.6000 102.6000 ;
	    RECT 1321.9501 81.6000 1322.8500 101.4000 ;
	    RECT 1324.2001 100.5000 1325.1000 101.7000 ;
	    RECT 1326.3000 100.5000 1327.5000 100.8000 ;
	    RECT 1331.4000 100.5000 1332.6000 100.8000 ;
	    RECT 1333.8000 100.5000 1334.7001 107.7000 ;
	    RECT 1336.2001 101.4000 1337.4000 102.6000 ;
	    RECT 1324.2001 99.3000 1325.4000 100.5000 ;
	    RECT 1326.3000 99.6000 1334.7001 100.5000 ;
	    RECT 1333.5000 99.3000 1334.7001 99.6000 ;
	    RECT 1336.3500 90.6000 1337.2500 101.4000 ;
	    RECT 1336.2001 89.4000 1337.4000 90.6000 ;
	    RECT 1288.2001 80.4000 1289.4000 81.6000 ;
	    RECT 1307.4000 80.4000 1308.6000 81.6000 ;
	    RECT 1314.6000 80.4000 1315.8000 81.6000 ;
	    RECT 1321.8000 80.4000 1323.0000 81.6000 ;
	    RECT 1281.0000 77.4000 1282.2001 78.6000 ;
	    RECT 1283.4000 77.4000 1284.6000 78.6000 ;
	    RECT 1276.2001 20.4000 1277.4000 21.6000 ;
	    RECT 1278.6000 20.4000 1279.8000 21.6000 ;
	    RECT 1276.3500 18.6000 1277.2500 20.4000 ;
	    RECT 1281.1500 18.6000 1282.0500 77.4000 ;
	    RECT 1288.3500 24.6000 1289.2500 80.4000 ;
	    RECT 1302.6000 74.4000 1303.8000 75.6000 ;
	    RECT 1302.7500 54.6000 1303.6500 74.4000 ;
	    RECT 1297.8000 53.4000 1299.0000 54.6000 ;
	    RECT 1302.6000 53.4000 1303.8000 54.6000 ;
	    RECT 1288.2001 23.4000 1289.4000 24.6000 ;
	    RECT 1276.2001 17.4000 1277.4000 18.6000 ;
	    RECT 1281.0000 17.4000 1282.2001 18.6000 ;
	    RECT 1297.9501 15.6000 1298.8500 53.4000 ;
	    RECT 1305.0000 23.4000 1306.2001 24.6000 ;
	    RECT 1305.1500 21.6000 1306.0500 23.4000 ;
	    RECT 1307.5500 21.6000 1308.4501 80.4000 ;
	    RECT 1343.5500 60.6000 1344.4501 161.4000 ;
	    RECT 1348.3500 141.6000 1349.2500 179.4000 ;
	    RECT 1348.2001 140.4000 1349.4000 141.6000 ;
	    RECT 1345.8000 134.4000 1347.0000 135.6000 ;
	    RECT 1345.9501 132.6000 1346.8500 134.4000 ;
	    RECT 1345.8000 131.4000 1347.0000 132.6000 ;
	    RECT 1350.7500 75.6000 1351.6500 341.4000 ;
	    RECT 1365.1500 324.6000 1366.0500 371.5500 ;
	    RECT 1367.4000 371.4000 1368.6000 371.5500 ;
	    RECT 1369.9501 324.6000 1370.8500 425.4000 ;
	    RECT 1377.1500 408.6000 1378.0500 440.4000 ;
	    RECT 1379.5500 435.6000 1380.4501 479.4000 ;
	    RECT 1379.4000 434.4000 1380.6000 435.6000 ;
	    RECT 1377.0000 407.4000 1378.2001 408.6000 ;
	    RECT 1377.1500 339.6000 1378.0500 407.4000 ;
	    RECT 1381.9501 342.6000 1382.8500 611.4000 ;
	    RECT 1384.3500 594.6000 1385.2500 611.4000 ;
	    RECT 1384.2001 593.4000 1385.4000 594.6000 ;
	    RECT 1386.7500 558.6000 1387.6500 629.4000 ;
	    RECT 1398.7500 621.6000 1399.6500 641.4000 ;
	    RECT 1403.5500 636.6000 1404.4501 644.4000 ;
	    RECT 1408.3500 642.6000 1409.2500 785.4000 ;
	    RECT 1413.1500 774.6000 1414.0500 800.4000 ;
	    RECT 1413.0000 773.4000 1414.2001 774.6000 ;
	    RECT 1410.6000 759.3000 1411.8000 767.7000 ;
	    RECT 1413.0000 761.4000 1414.2001 762.6000 ;
	    RECT 1415.4000 756.3000 1416.6000 773.7000 ;
	    RECT 1410.6000 749.4000 1411.8000 750.6000 ;
	    RECT 1410.7500 741.6000 1411.6500 749.4000 ;
	    RECT 1410.6000 740.4000 1411.8000 741.6000 ;
	    RECT 1415.4000 737.4000 1416.6000 738.6000 ;
	    RECT 1410.6000 725.4000 1411.8000 726.6000 ;
	    RECT 1408.2001 641.4000 1409.4000 642.6000 ;
	    RECT 1403.4000 635.4000 1404.6000 636.6000 ;
	    RECT 1389.0000 620.4000 1390.2001 621.6000 ;
	    RECT 1398.6000 620.4000 1399.8000 621.6000 ;
	    RECT 1386.6000 557.4000 1387.8000 558.6000 ;
	    RECT 1389.1500 555.6000 1390.0500 620.4000 ;
	    RECT 1408.2001 617.4000 1409.4000 618.6000 ;
	    RECT 1408.3500 615.6000 1409.2500 617.4000 ;
	    RECT 1408.2001 614.4000 1409.4000 615.6000 ;
	    RECT 1410.7500 588.6000 1411.6500 725.4000 ;
	    RECT 1415.5500 714.6000 1416.4501 737.4000 ;
	    RECT 1415.4000 713.4000 1416.6000 714.6000 ;
	    RECT 1415.5500 705.6000 1416.4501 713.4000 ;
	    RECT 1415.4000 704.4000 1416.6000 705.6000 ;
	    RECT 1413.0000 677.4000 1414.2001 678.6000 ;
	    RECT 1403.4000 587.4000 1404.6000 588.6000 ;
	    RECT 1410.6000 587.4000 1411.8000 588.6000 ;
	    RECT 1405.8000 584.4000 1407.0000 585.6000 ;
	    RECT 1405.9501 582.6000 1406.8500 584.4000 ;
	    RECT 1405.8000 581.4000 1407.0000 582.6000 ;
	    RECT 1391.4000 557.4000 1392.6000 558.6000 ;
	    RECT 1389.0000 554.4000 1390.2001 555.6000 ;
	    RECT 1386.6000 551.4000 1387.8000 552.6000 ;
	    RECT 1386.7500 531.6000 1387.6500 551.4000 ;
	    RECT 1386.6000 530.4000 1387.8000 531.6000 ;
	    RECT 1386.7500 498.6000 1387.6500 530.4000 ;
	    RECT 1389.0000 510.4500 1390.2001 510.6000 ;
	    RECT 1391.5500 510.4500 1392.4501 557.4000 ;
	    RECT 1393.8000 527.4000 1395.0000 528.6000 ;
	    RECT 1389.0000 509.5500 1392.4501 510.4500 ;
	    RECT 1389.0000 509.4000 1390.2001 509.5500 ;
	    RECT 1389.1500 501.6000 1390.0500 509.4000 ;
	    RECT 1393.9501 504.6000 1394.8500 527.4000 ;
	    RECT 1403.4000 524.4000 1404.6000 525.6000 ;
	    RECT 1403.5500 510.6000 1404.4501 524.4000 ;
	    RECT 1403.4000 509.4000 1404.6000 510.6000 ;
	    RECT 1393.8000 503.4000 1395.0000 504.6000 ;
	    RECT 1389.0000 500.4000 1390.2001 501.6000 ;
	    RECT 1386.6000 497.4000 1387.8000 498.6000 ;
	    RECT 1386.7500 468.6000 1387.6500 497.4000 ;
	    RECT 1389.0000 470.4000 1390.2001 471.6000 ;
	    RECT 1386.6000 467.4000 1387.8000 468.6000 ;
	    RECT 1384.2001 461.4000 1385.4000 462.6000 ;
	    RECT 1384.2001 440.4000 1385.4000 441.6000 ;
	    RECT 1384.3500 414.6000 1385.2500 440.4000 ;
	    RECT 1384.2001 413.4000 1385.4000 414.6000 ;
	    RECT 1386.6000 407.4000 1387.8000 408.6000 ;
	    RECT 1386.7500 381.6000 1387.6500 407.4000 ;
	    RECT 1386.6000 380.4000 1387.8000 381.6000 ;
	    RECT 1389.1500 342.6000 1390.0500 470.4000 ;
	    RECT 1393.8000 467.4000 1395.0000 468.6000 ;
	    RECT 1391.4000 464.4000 1392.6000 465.6000 ;
	    RECT 1391.5500 456.6000 1392.4501 464.4000 ;
	    RECT 1393.9501 462.6000 1394.8500 467.4000 ;
	    RECT 1393.8000 461.4000 1395.0000 462.6000 ;
	    RECT 1391.4000 455.4000 1392.6000 456.6000 ;
	    RECT 1393.8000 413.4000 1395.0000 414.6000 ;
	    RECT 1393.9501 411.6000 1394.8500 413.4000 ;
	    RECT 1393.8000 410.4000 1395.0000 411.6000 ;
	    RECT 1403.5500 408.6000 1404.4501 509.4000 ;
	    RECT 1410.6000 497.4000 1411.8000 498.6000 ;
	    RECT 1410.7500 468.6000 1411.6500 497.4000 ;
	    RECT 1410.6000 467.4000 1411.8000 468.6000 ;
	    RECT 1405.8000 437.4000 1407.0000 438.6000 ;
	    RECT 1403.4000 407.4000 1404.6000 408.6000 ;
	    RECT 1391.4000 404.4000 1392.6000 405.6000 ;
	    RECT 1391.5500 402.6000 1392.4501 404.4000 ;
	    RECT 1391.4000 401.4000 1392.6000 402.6000 ;
	    RECT 1405.9501 390.6000 1406.8500 437.4000 ;
	    RECT 1410.6000 434.4000 1411.8000 435.6000 ;
	    RECT 1410.7500 426.6000 1411.6500 434.4000 ;
	    RECT 1410.6000 425.4000 1411.8000 426.6000 ;
	    RECT 1408.2001 401.4000 1409.4000 402.6000 ;
	    RECT 1405.8000 389.4000 1407.0000 390.6000 ;
	    RECT 1393.8000 377.4000 1395.0000 378.6000 ;
	    RECT 1391.4000 347.4000 1392.6000 348.6000 ;
	    RECT 1381.8000 341.4000 1383.0000 342.6000 ;
	    RECT 1389.0000 341.4000 1390.2001 342.6000 ;
	    RECT 1391.5500 339.6000 1392.4501 347.4000 ;
	    RECT 1393.9501 345.6000 1394.8500 377.4000 ;
	    RECT 1405.9501 360.6000 1406.8500 389.4000 ;
	    RECT 1408.3500 375.6000 1409.2500 401.4000 ;
	    RECT 1408.2001 374.4000 1409.4000 375.6000 ;
	    RECT 1405.8000 359.4000 1407.0000 360.6000 ;
	    RECT 1393.8000 344.4000 1395.0000 345.6000 ;
	    RECT 1405.8000 344.4000 1407.0000 345.6000 ;
	    RECT 1377.0000 338.4000 1378.2001 339.6000 ;
	    RECT 1391.4000 338.4000 1392.6000 339.6000 ;
	    RECT 1405.9501 336.6000 1406.8500 344.4000 ;
	    RECT 1408.2001 341.4000 1409.4000 342.6000 ;
	    RECT 1396.2001 335.4000 1397.4000 336.6000 ;
	    RECT 1405.8000 335.4000 1407.0000 336.6000 ;
	    RECT 1391.4000 329.4000 1392.6000 330.6000 ;
	    RECT 1365.0000 323.4000 1366.2001 324.6000 ;
	    RECT 1369.8000 323.4000 1371.0000 324.6000 ;
	    RECT 1389.0000 323.4000 1390.2001 324.6000 ;
	    RECT 1362.6000 320.4000 1363.8000 321.6000 ;
	    RECT 1362.7500 288.6000 1363.6500 320.4000 ;
	    RECT 1389.1500 318.6000 1390.0500 323.4000 ;
	    RECT 1391.5500 318.6000 1392.4501 329.4000 ;
	    RECT 1393.8000 320.4000 1395.0000 321.6000 ;
	    RECT 1365.0000 317.4000 1366.2001 318.6000 ;
	    RECT 1389.0000 317.4000 1390.2001 318.6000 ;
	    RECT 1391.4000 317.4000 1392.6000 318.6000 ;
	    RECT 1362.6000 287.4000 1363.8000 288.6000 ;
	    RECT 1365.1500 258.6000 1366.0500 317.4000 ;
	    RECT 1393.9501 306.6000 1394.8500 320.4000 ;
	    RECT 1396.3500 318.6000 1397.2500 335.4000 ;
	    RECT 1396.2001 317.4000 1397.4000 318.6000 ;
	    RECT 1401.0000 317.4000 1402.2001 318.6000 ;
	    RECT 1401.1500 315.6000 1402.0500 317.4000 ;
	    RECT 1401.0000 314.4000 1402.2001 315.6000 ;
	    RECT 1408.3500 306.6000 1409.2500 341.4000 ;
	    RECT 1393.8000 305.4000 1395.0000 306.6000 ;
	    RECT 1408.2001 305.4000 1409.4000 306.6000 ;
	    RECT 1389.0000 299.4000 1390.2001 300.6000 ;
	    RECT 1367.4000 290.4000 1368.6000 291.6000 ;
	    RECT 1367.5500 282.6000 1368.4501 290.4000 ;
	    RECT 1372.2001 287.4000 1373.4000 288.6000 ;
	    RECT 1369.8000 284.4000 1371.0000 285.6000 ;
	    RECT 1367.4000 281.4000 1368.6000 282.6000 ;
	    RECT 1369.9501 276.6000 1370.8500 284.4000 ;
	    RECT 1369.8000 275.4000 1371.0000 276.6000 ;
	    RECT 1369.9501 261.6000 1370.8500 275.4000 ;
	    RECT 1369.8000 260.4000 1371.0000 261.6000 ;
	    RECT 1372.3500 258.6000 1373.2500 287.4000 ;
	    RECT 1389.1500 264.6000 1390.0500 299.4000 ;
	    RECT 1393.9501 285.6000 1394.8500 305.4000 ;
	    RECT 1405.8000 287.4000 1407.0000 288.6000 ;
	    RECT 1405.9501 285.6000 1406.8500 287.4000 ;
	    RECT 1393.8000 284.4000 1395.0000 285.6000 ;
	    RECT 1405.8000 284.4000 1407.0000 285.6000 ;
	    RECT 1403.4000 281.4000 1404.6000 282.6000 ;
	    RECT 1398.6000 278.4000 1399.8000 279.6000 ;
	    RECT 1398.7500 264.6000 1399.6500 278.4000 ;
	    RECT 1389.0000 263.4000 1390.2001 264.6000 ;
	    RECT 1398.6000 263.4000 1399.8000 264.6000 ;
	    RECT 1398.7500 258.6000 1399.6500 263.4000 ;
	    RECT 1403.5500 261.6000 1404.4501 281.4000 ;
	    RECT 1403.4000 260.4000 1404.6000 261.6000 ;
	    RECT 1405.9501 258.6000 1406.8500 284.4000 ;
	    RECT 1360.2001 257.4000 1361.4000 258.6000 ;
	    RECT 1365.0000 257.4000 1366.2001 258.6000 ;
	    RECT 1372.2001 257.4000 1373.4000 258.6000 ;
	    RECT 1391.4000 257.4000 1392.6000 258.6000 ;
	    RECT 1398.6000 257.4000 1399.8000 258.6000 ;
	    RECT 1405.8000 257.4000 1407.0000 258.6000 ;
	    RECT 1360.3500 255.6000 1361.2500 257.4000 ;
	    RECT 1360.2001 254.4000 1361.4000 255.6000 ;
	    RECT 1379.4000 239.4000 1380.6000 240.6000 ;
	    RECT 1377.0000 227.4000 1378.2001 228.6000 ;
	    RECT 1377.1500 216.6000 1378.0500 227.4000 ;
	    RECT 1379.5500 225.6000 1380.4501 239.4000 ;
	    RECT 1379.4000 224.4000 1380.6000 225.6000 ;
	    RECT 1386.6000 221.4000 1387.8000 222.6000 ;
	    RECT 1377.0000 215.4000 1378.2001 216.6000 ;
	    RECT 1362.3000 202.5000 1363.5000 203.7000 ;
	    RECT 1365.0000 202.5000 1371.3000 203.4000 ;
	    RECT 1372.2001 202.5000 1373.4000 203.7000 ;
	    RECT 1360.2001 197.4000 1361.4000 198.6000 ;
	    RECT 1360.3500 186.6000 1361.2500 197.4000 ;
	    RECT 1362.3000 195.3000 1363.2001 202.5000 ;
	    RECT 1365.0000 202.2000 1366.2001 202.5000 ;
	    RECT 1370.1000 202.2000 1371.3000 202.5000 ;
	    RECT 1372.5000 201.3000 1373.4000 202.5000 ;
	    RECT 1366.2001 200.4000 1373.4000 201.3000 ;
	    RECT 1374.6000 200.4000 1375.8000 201.6000 ;
	    RECT 1366.2001 200.1000 1367.4000 200.4000 ;
	    RECT 1372.5000 195.3000 1373.4000 200.4000 ;
	    RECT 1374.7500 198.6000 1375.6500 200.4000 ;
	    RECT 1374.6000 197.4000 1375.8000 198.6000 ;
	    RECT 1362.3000 194.1000 1363.5000 195.3000 ;
	    RECT 1372.2001 194.1000 1373.4000 195.3000 ;
	    RECT 1360.2001 185.4000 1361.4000 186.6000 ;
	    RECT 1355.4000 176.4000 1356.6000 177.6000 ;
	    RECT 1355.5500 168.6000 1356.4501 176.4000 ;
	    RECT 1355.4000 167.4000 1356.6000 168.6000 ;
	    RECT 1360.2001 164.4000 1361.4000 165.6000 ;
	    RECT 1360.3500 162.6000 1361.2500 164.4000 ;
	    RECT 1360.2001 161.4000 1361.4000 162.6000 ;
	    RECT 1362.6000 156.3000 1363.8000 176.7000 ;
	    RECT 1365.0000 156.3000 1366.2001 176.7000 ;
	    RECT 1367.4000 156.3000 1368.6000 173.7000 ;
	    RECT 1369.8000 167.4000 1371.0000 168.6000 ;
	    RECT 1369.9501 162.6000 1370.8500 167.4000 ;
	    RECT 1369.8000 161.4000 1371.0000 162.6000 ;
	    RECT 1372.2001 156.3000 1373.4000 173.7000 ;
	    RECT 1374.6000 173.4000 1375.8000 174.6000 ;
	    RECT 1374.7500 168.6000 1375.6500 173.4000 ;
	    RECT 1374.6000 167.4000 1375.8000 168.6000 ;
	    RECT 1374.6000 158.4000 1375.8000 159.6000 ;
	    RECT 1369.8000 101.4000 1371.0000 102.6000 ;
	    RECT 1369.9501 81.6000 1370.8500 101.4000 ;
	    RECT 1362.6000 80.4000 1363.8000 81.6000 ;
	    RECT 1369.8000 80.4000 1371.0000 81.6000 ;
	    RECT 1350.6000 74.4000 1351.8000 75.6000 ;
	    RECT 1343.4000 59.4000 1344.6000 60.6000 ;
	    RECT 1362.7500 42.6000 1363.6500 80.4000 ;
	    RECT 1372.2001 77.4000 1373.4000 78.6000 ;
	    RECT 1369.8000 47.4000 1371.0000 48.6000 ;
	    RECT 1362.6000 41.4000 1363.8000 42.6000 ;
	    RECT 1341.0000 35.4000 1342.2001 36.6000 ;
	    RECT 1341.1500 30.6000 1342.0500 35.4000 ;
	    RECT 1369.9501 30.6000 1370.8500 47.4000 ;
	    RECT 1341.0000 29.4000 1342.2001 30.6000 ;
	    RECT 1369.8000 29.4000 1371.0000 30.6000 ;
	    RECT 1372.3500 24.6000 1373.2500 77.4000 ;
	    RECT 1374.7500 36.6000 1375.6500 158.4000 ;
	    RECT 1377.0000 156.3000 1378.2001 173.7000 ;
	    RECT 1379.4000 156.3000 1380.6000 176.7000 ;
	    RECT 1381.8000 156.3000 1383.0000 176.7000 ;
	    RECT 1384.2001 156.3000 1385.4000 176.7000 ;
	    RECT 1386.7500 174.6000 1387.6500 221.4000 ;
	    RECT 1386.6000 173.4000 1387.8000 174.6000 ;
	    RECT 1379.4000 149.4000 1380.6000 150.6000 ;
	    RECT 1377.0000 143.4000 1378.2001 144.6000 ;
	    RECT 1377.1500 135.6000 1378.0500 143.4000 ;
	    RECT 1379.5500 141.6000 1380.4501 149.4000 ;
	    RECT 1379.4000 140.4000 1380.6000 141.6000 ;
	    RECT 1386.6000 140.4000 1387.8000 141.6000 ;
	    RECT 1386.7500 138.6000 1387.6500 140.4000 ;
	    RECT 1384.2001 137.4000 1385.4000 138.6000 ;
	    RECT 1386.6000 137.4000 1387.8000 138.6000 ;
	    RECT 1377.0000 134.4000 1378.2001 135.6000 ;
	    RECT 1384.3500 108.6000 1385.2500 137.4000 ;
	    RECT 1391.5500 132.6000 1392.4501 257.4000 ;
	    RECT 1405.8000 251.4000 1407.0000 252.6000 ;
	    RECT 1405.9501 228.6000 1406.8500 251.4000 ;
	    RECT 1413.1500 240.6000 1414.0500 677.4000 ;
	    RECT 1415.4000 617.4000 1416.6000 618.6000 ;
	    RECT 1415.4000 614.4000 1416.6000 615.6000 ;
	    RECT 1415.5500 504.6000 1416.4501 614.4000 ;
	    RECT 1417.9501 612.6000 1418.8500 800.4000 ;
	    RECT 1420.2001 764.4000 1421.4000 765.6000 ;
	    RECT 1420.3500 750.6000 1421.2500 764.4000 ;
	    RECT 1420.2001 749.4000 1421.4000 750.6000 ;
	    RECT 1420.2001 707.4000 1421.4000 708.6000 ;
	    RECT 1422.7500 684.6000 1423.6500 830.4000 ;
	    RECT 1425.1500 828.6000 1426.0500 857.4000 ;
	    RECT 1425.0000 827.4000 1426.2001 828.6000 ;
	    RECT 1425.1500 744.6000 1426.0500 827.4000 ;
	    RECT 1427.5500 804.6000 1428.4501 911.4000 ;
	    RECT 1437.1500 861.6000 1438.0500 980.4000 ;
	    RECT 1439.4000 977.4000 1440.6000 978.6000 ;
	    RECT 1439.5500 972.6000 1440.4501 977.4000 ;
	    RECT 1439.4000 971.4000 1440.6000 972.6000 ;
	    RECT 1444.3500 957.6000 1445.2500 1001.4000 ;
	    RECT 1444.2001 956.4000 1445.4000 957.6000 ;
	    RECT 1441.8000 923.4000 1443.0000 924.6000 ;
	    RECT 1441.9501 888.6000 1442.8500 923.4000 ;
	    RECT 1441.8000 887.4000 1443.0000 888.6000 ;
	    RECT 1441.9501 882.6000 1442.8500 887.4000 ;
	    RECT 1441.8000 881.4000 1443.0000 882.6000 ;
	    RECT 1437.0000 860.4000 1438.2001 861.6000 ;
	    RECT 1432.2001 851.4000 1433.4000 852.6000 ;
	    RECT 1432.3500 840.6000 1433.2500 851.4000 ;
	    RECT 1432.2001 839.4000 1433.4000 840.6000 ;
	    RECT 1432.3500 819.6000 1433.2500 839.4000 ;
	    RECT 1432.2001 818.4000 1433.4000 819.6000 ;
	    RECT 1427.4000 803.4000 1428.6000 804.6000 ;
	    RECT 1427.5500 795.6000 1428.4501 803.4000 ;
	    RECT 1427.4000 794.4000 1428.6000 795.6000 ;
	    RECT 1437.0000 794.4000 1438.2001 795.6000 ;
	    RECT 1427.4000 773.4000 1428.6000 774.6000 ;
	    RECT 1425.0000 743.4000 1426.2001 744.6000 ;
	    RECT 1425.1500 741.6000 1426.0500 743.4000 ;
	    RECT 1425.0000 740.4000 1426.2001 741.6000 ;
	    RECT 1422.6000 683.4000 1423.8000 684.6000 ;
	    RECT 1420.2001 641.4000 1421.4000 642.6000 ;
	    RECT 1420.3500 636.6000 1421.2500 641.4000 ;
	    RECT 1420.2001 635.4000 1421.4000 636.6000 ;
	    RECT 1417.8000 611.4000 1419.0000 612.6000 ;
	    RECT 1417.8000 599.4000 1419.0000 600.6000 ;
	    RECT 1417.9501 582.6000 1418.8500 599.4000 ;
	    RECT 1422.7500 594.6000 1423.6500 683.4000 ;
	    RECT 1425.0000 674.4000 1426.2001 675.6000 ;
	    RECT 1425.1500 666.6000 1426.0500 674.4000 ;
	    RECT 1425.0000 665.4000 1426.2001 666.6000 ;
	    RECT 1427.5500 615.6000 1428.4501 773.4000 ;
	    RECT 1429.8000 756.3000 1431.0000 773.7000 ;
	    RECT 1432.2001 761.4000 1433.4000 762.6000 ;
	    RECT 1432.3500 744.6000 1433.2500 761.4000 ;
	    RECT 1432.2001 743.4000 1433.4000 744.6000 ;
	    RECT 1432.3500 675.6000 1433.2500 743.4000 ;
	    RECT 1434.6000 707.4000 1435.8000 708.6000 ;
	    RECT 1434.7500 702.6000 1435.6500 707.4000 ;
	    RECT 1434.6000 701.4000 1435.8000 702.6000 ;
	    RECT 1432.2001 674.4000 1433.4000 675.6000 ;
	    RECT 1432.3500 666.6000 1433.2500 674.4000 ;
	    RECT 1432.2001 665.4000 1433.4000 666.6000 ;
	    RECT 1437.1500 648.6000 1438.0500 794.4000 ;
	    RECT 1439.4000 764.4000 1440.6000 765.6000 ;
	    RECT 1439.5500 762.6000 1440.4501 764.4000 ;
	    RECT 1439.4000 761.4000 1440.6000 762.6000 ;
	    RECT 1441.8000 701.4000 1443.0000 702.6000 ;
	    RECT 1439.4000 689.4000 1440.6000 690.6000 ;
	    RECT 1439.5500 681.6000 1440.4501 689.4000 ;
	    RECT 1439.4000 680.4000 1440.6000 681.6000 ;
	    RECT 1441.9501 672.6000 1442.8500 701.4000 ;
	    RECT 1441.8000 671.4000 1443.0000 672.6000 ;
	    RECT 1437.0000 647.4000 1438.2001 648.6000 ;
	    RECT 1429.8000 644.4000 1431.0000 645.6000 ;
	    RECT 1429.9501 630.6000 1430.8500 644.4000 ;
	    RECT 1429.8000 629.4000 1431.0000 630.6000 ;
	    RECT 1429.9501 618.6000 1430.8500 629.4000 ;
	    RECT 1437.1500 624.6000 1438.0500 647.4000 ;
	    RECT 1444.3500 642.6000 1445.2500 956.4000 ;
	    RECT 1446.7500 672.6000 1447.6500 1331.4000 ;
	    RECT 1449.1500 1308.6000 1450.0500 1334.5500 ;
	    RECT 1453.9501 1320.6000 1454.8500 1340.4000 ;
	    RECT 1485.1500 1338.6000 1486.0500 1340.4000 ;
	    RECT 1470.6000 1337.4000 1471.8000 1338.6000 ;
	    RECT 1485.0000 1337.4000 1486.2001 1338.6000 ;
	    RECT 1470.7500 1320.6000 1471.6500 1337.4000 ;
	    RECT 1473.0000 1334.4000 1474.2001 1335.6000 ;
	    RECT 1453.8000 1319.4000 1455.0000 1320.6000 ;
	    RECT 1470.6000 1319.4000 1471.8000 1320.6000 ;
	    RECT 1470.7500 1308.6000 1471.6500 1319.4000 ;
	    RECT 1449.0000 1307.4000 1450.2001 1308.6000 ;
	    RECT 1470.6000 1307.4000 1471.8000 1308.6000 ;
	    RECT 1463.4000 1301.4000 1464.6000 1302.6000 ;
	    RECT 1449.0000 1266.3000 1450.2001 1286.7001 ;
	    RECT 1451.4000 1266.3000 1452.6000 1286.7001 ;
	    RECT 1453.8000 1266.3000 1455.0000 1286.7001 ;
	    RECT 1456.2001 1269.3000 1457.4000 1286.7001 ;
	    RECT 1458.6000 1283.4000 1459.8000 1284.6000 ;
	    RECT 1458.7500 1266.4501 1459.6500 1283.4000 ;
	    RECT 1461.0000 1269.3000 1462.2001 1286.7001 ;
	    RECT 1463.5500 1281.6000 1464.4501 1301.4000 ;
	    RECT 1473.1500 1299.4501 1474.0500 1334.4000 ;
	    RECT 1475.4000 1304.4000 1476.6000 1305.6000 ;
	    RECT 1475.5500 1302.6000 1476.4501 1304.4000 ;
	    RECT 1475.4000 1301.4000 1476.6000 1302.6000 ;
	    RECT 1473.1500 1298.5500 1476.4501 1299.4501 ;
	    RECT 1463.4000 1280.4000 1464.6000 1281.6000 ;
	    RECT 1465.8000 1269.3000 1467.0000 1286.7001 ;
	    RECT 1458.7500 1265.5500 1462.0500 1266.4501 ;
	    RECT 1458.6000 1259.4000 1459.8000 1260.6000 ;
	    RECT 1451.4000 1248.4501 1452.6000 1248.6000 ;
	    RECT 1451.4000 1247.5500 1454.8500 1248.4501 ;
	    RECT 1451.4000 1247.4000 1452.6000 1247.5500 ;
	    RECT 1451.4000 1241.4000 1452.6000 1242.6000 ;
	    RECT 1451.5500 1221.6000 1452.4501 1241.4000 ;
	    RECT 1451.4000 1220.4000 1452.6000 1221.6000 ;
	    RECT 1449.0000 1124.4000 1450.2001 1125.6000 ;
	    RECT 1449.1500 1002.4500 1450.0500 1124.4000 ;
	    RECT 1451.5500 1104.6000 1452.4501 1220.4000 ;
	    RECT 1453.9501 1218.6000 1454.8500 1247.5500 ;
	    RECT 1458.7500 1245.6000 1459.6500 1259.4000 ;
	    RECT 1458.6000 1244.4000 1459.8000 1245.6000 ;
	    RECT 1458.6000 1241.4000 1459.8000 1242.6000 ;
	    RECT 1453.8000 1217.4000 1455.0000 1218.6000 ;
	    RECT 1461.1500 1176.6000 1462.0500 1265.5500 ;
	    RECT 1465.8000 1265.4000 1467.0000 1266.6000 ;
	    RECT 1468.2001 1266.3000 1469.4000 1286.7001 ;
	    RECT 1470.6000 1266.3000 1471.8000 1286.7001 ;
	    RECT 1473.0000 1277.4000 1474.2001 1278.6000 ;
	    RECT 1463.4000 1247.4000 1464.6000 1248.6000 ;
	    RECT 1463.5500 1242.6000 1464.4501 1247.4000 ;
	    RECT 1463.4000 1241.4000 1464.6000 1242.6000 ;
	    RECT 1463.4000 1214.4000 1464.6000 1215.6000 ;
	    RECT 1461.0000 1175.4000 1462.2001 1176.6000 ;
	    RECT 1461.1500 1164.6000 1462.0500 1175.4000 ;
	    RECT 1461.0000 1163.4000 1462.2001 1164.6000 ;
	    RECT 1451.4000 1103.4000 1452.6000 1104.6000 ;
	    RECT 1453.8000 1004.4000 1455.0000 1005.6000 ;
	    RECT 1451.4000 1002.4500 1452.6000 1002.6000 ;
	    RECT 1449.1500 1001.5500 1452.6000 1002.4500 ;
	    RECT 1451.4000 1001.4000 1452.6000 1001.5500 ;
	    RECT 1451.5500 984.6000 1452.4501 1001.4000 ;
	    RECT 1451.4000 983.4000 1452.6000 984.6000 ;
	    RECT 1453.9501 948.6000 1454.8500 1004.4000 ;
	    RECT 1453.8000 947.4000 1455.0000 948.6000 ;
	    RECT 1453.9501 774.6000 1454.8500 947.4000 ;
	    RECT 1456.2001 929.4000 1457.4000 930.6000 ;
	    RECT 1456.3500 924.6000 1457.2500 929.4000 ;
	    RECT 1456.2001 923.4000 1457.4000 924.6000 ;
	    RECT 1461.0000 821.4000 1462.2001 822.6000 ;
	    RECT 1456.2001 803.4000 1457.4000 804.6000 ;
	    RECT 1456.3500 792.6000 1457.2500 803.4000 ;
	    RECT 1458.6000 797.4000 1459.8000 798.6000 ;
	    RECT 1456.2001 791.4000 1457.4000 792.6000 ;
	    RECT 1453.8000 773.4000 1455.0000 774.6000 ;
	    RECT 1456.3500 726.6000 1457.2500 791.4000 ;
	    RECT 1458.7500 786.6000 1459.6500 797.4000 ;
	    RECT 1458.6000 785.4000 1459.8000 786.6000 ;
	    RECT 1458.6000 780.4500 1459.8000 780.6000 ;
	    RECT 1461.1500 780.4500 1462.0500 821.4000 ;
	    RECT 1463.5500 807.6000 1464.4501 1214.4000 ;
	    RECT 1465.9501 1050.6000 1466.8500 1265.4000 ;
	    RECT 1473.1500 1254.6000 1474.0500 1277.4000 ;
	    RECT 1475.5500 1266.6000 1476.4501 1298.5500 ;
	    RECT 1477.8000 1296.3000 1479.0000 1316.7001 ;
	    RECT 1480.2001 1296.3000 1481.4000 1316.7001 ;
	    RECT 1482.6000 1296.3000 1483.8000 1313.7001 ;
	    RECT 1485.0000 1301.4000 1486.2001 1302.6000 ;
	    RECT 1485.1500 1296.6000 1486.0500 1301.4000 ;
	    RECT 1485.0000 1295.4000 1486.2001 1296.6000 ;
	    RECT 1487.4000 1296.3000 1488.6000 1313.7001 ;
	    RECT 1489.8000 1298.4000 1491.0000 1299.6000 ;
	    RECT 1485.0000 1280.4000 1486.2001 1281.6000 ;
	    RECT 1477.8000 1274.4000 1479.0000 1275.6000 ;
	    RECT 1477.9501 1272.6000 1478.8500 1274.4000 ;
	    RECT 1477.8000 1271.4000 1479.0000 1272.6000 ;
	    RECT 1482.6000 1271.4000 1483.8000 1272.6000 ;
	    RECT 1477.9501 1266.6000 1478.8500 1271.4000 ;
	    RECT 1475.4000 1265.4000 1476.6000 1266.6000 ;
	    RECT 1477.8000 1265.4000 1479.0000 1266.6000 ;
	    RECT 1477.9501 1254.6000 1478.8500 1265.4000 ;
	    RECT 1482.7500 1254.6000 1483.6500 1271.4000 ;
	    RECT 1485.1500 1260.6000 1486.0500 1280.4000 ;
	    RECT 1487.4000 1265.4000 1488.6000 1266.6000 ;
	    RECT 1485.0000 1259.4000 1486.2001 1260.6000 ;
	    RECT 1473.0000 1253.4000 1474.2001 1254.6000 ;
	    RECT 1477.8000 1253.4000 1479.0000 1254.6000 ;
	    RECT 1482.6000 1253.4000 1483.8000 1254.6000 ;
	    RECT 1477.9501 1242.6000 1478.8500 1253.4000 ;
	    RECT 1482.6000 1247.4000 1483.8000 1248.6000 ;
	    RECT 1477.8000 1241.4000 1479.0000 1242.6000 ;
	    RECT 1482.7500 1236.6000 1483.6500 1247.4000 ;
	    RECT 1482.6000 1235.4000 1483.8000 1236.6000 ;
	    RECT 1477.8000 1229.4000 1479.0000 1230.6000 ;
	    RECT 1470.6000 1121.4000 1471.8000 1122.6000 ;
	    RECT 1470.7500 1098.6000 1471.6500 1121.4000 ;
	    RECT 1477.9501 1104.6000 1478.8500 1229.4000 ;
	    RECT 1487.5500 1158.4501 1488.4501 1265.4000 ;
	    RECT 1489.9501 1236.6000 1490.8500 1298.4000 ;
	    RECT 1492.2001 1296.3000 1493.4000 1313.7001 ;
	    RECT 1494.6000 1296.3000 1495.8000 1316.7001 ;
	    RECT 1497.0000 1296.3000 1498.2001 1316.7001 ;
	    RECT 1499.4000 1296.3000 1500.6000 1316.7001 ;
	    RECT 1513.8000 1310.4000 1515.0000 1311.6000 ;
	    RECT 1501.8000 1307.4000 1503.0000 1308.6000 ;
	    RECT 1501.9501 1278.6000 1502.8500 1307.4000 ;
	    RECT 1513.9501 1284.6000 1514.8500 1310.4000 ;
	    RECT 1516.3500 1305.6000 1517.2500 1343.4000 ;
	    RECT 1518.6000 1325.4000 1519.8000 1326.6000 ;
	    RECT 1516.2001 1304.4000 1517.4000 1305.6000 ;
	    RECT 1509.0000 1283.4000 1510.2001 1284.6000 ;
	    RECT 1513.8000 1283.4000 1515.0000 1284.6000 ;
	    RECT 1492.2001 1277.4000 1493.4000 1278.6000 ;
	    RECT 1501.8000 1277.4000 1503.0000 1278.6000 ;
	    RECT 1489.8000 1235.4000 1491.0000 1236.6000 ;
	    RECT 1489.9501 1230.6000 1490.8500 1235.4000 ;
	    RECT 1489.8000 1229.4000 1491.0000 1230.6000 ;
	    RECT 1489.8000 1158.4501 1491.0000 1158.6000 ;
	    RECT 1487.5500 1157.5500 1491.0000 1158.4501 ;
	    RECT 1489.8000 1157.4000 1491.0000 1157.5500 ;
	    RECT 1477.8000 1103.4000 1479.0000 1104.6000 ;
	    RECT 1470.6000 1097.4000 1471.8000 1098.6000 ;
	    RECT 1468.2001 1056.3000 1469.4000 1076.7001 ;
	    RECT 1470.6000 1056.3000 1471.8000 1076.7001 ;
	    RECT 1473.0000 1056.3000 1474.2001 1076.7001 ;
	    RECT 1475.4000 1056.3000 1476.6000 1073.7001 ;
	    RECT 1477.9501 1059.6000 1478.8500 1103.4000 ;
	    RECT 1482.6000 1100.4000 1483.8000 1101.6000 ;
	    RECT 1477.8000 1058.4000 1479.0000 1059.6000 ;
	    RECT 1465.8000 1049.4000 1467.0000 1050.6000 ;
	    RECT 1470.6000 1049.4000 1471.8000 1050.6000 ;
	    RECT 1465.8000 998.4000 1467.0000 999.6000 ;
	    RECT 1465.9501 996.6000 1466.8500 998.4000 ;
	    RECT 1465.8000 995.4000 1467.0000 996.6000 ;
	    RECT 1465.8000 980.4000 1467.0000 981.6000 ;
	    RECT 1465.9501 978.6000 1466.8500 980.4000 ;
	    RECT 1465.8000 977.4000 1467.0000 978.6000 ;
	    RECT 1468.2001 977.4000 1469.4000 978.6000 ;
	    RECT 1468.3500 951.6000 1469.2500 977.4000 ;
	    RECT 1468.2001 950.4000 1469.4000 951.6000 ;
	    RECT 1465.8000 887.4000 1467.0000 888.6000 ;
	    RECT 1463.4000 806.4000 1464.6000 807.6000 ;
	    RECT 1463.4000 803.4000 1464.6000 804.6000 ;
	    RECT 1463.5500 795.6000 1464.4501 803.4000 ;
	    RECT 1465.9501 798.6000 1466.8500 887.4000 ;
	    RECT 1468.2001 809.4000 1469.4000 810.6000 ;
	    RECT 1465.8000 797.4000 1467.0000 798.6000 ;
	    RECT 1463.4000 794.4000 1464.6000 795.6000 ;
	    RECT 1458.6000 779.5500 1462.0500 780.4500 ;
	    RECT 1458.6000 779.4000 1459.8000 779.5500 ;
	    RECT 1461.0000 758.4000 1462.2001 759.6000 ;
	    RECT 1458.6000 734.4000 1459.8000 735.6000 ;
	    RECT 1456.2001 725.4000 1457.4000 726.6000 ;
	    RECT 1458.7500 714.6000 1459.6500 734.4000 ;
	    RECT 1461.1500 732.6000 1462.0500 758.4000 ;
	    RECT 1461.0000 731.4000 1462.2001 732.6000 ;
	    RECT 1458.6000 713.4000 1459.8000 714.6000 ;
	    RECT 1449.0000 704.4000 1450.2001 705.6000 ;
	    RECT 1449.1500 702.6000 1450.0500 704.4000 ;
	    RECT 1449.0000 701.4000 1450.2001 702.6000 ;
	    RECT 1451.4000 701.4000 1452.6000 702.6000 ;
	    RECT 1458.6000 701.4000 1459.8000 702.6000 ;
	    RECT 1446.6000 671.4000 1447.8000 672.6000 ;
	    RECT 1449.1500 648.6000 1450.0500 701.4000 ;
	    RECT 1456.2001 698.4000 1457.4000 699.6000 ;
	    RECT 1456.3500 696.6000 1457.2500 698.4000 ;
	    RECT 1451.4000 695.4000 1452.6000 696.6000 ;
	    RECT 1456.2001 695.4000 1457.4000 696.6000 ;
	    RECT 1451.5500 675.6000 1452.4501 695.4000 ;
	    RECT 1453.8000 677.4000 1455.0000 678.6000 ;
	    RECT 1451.4000 674.4000 1452.6000 675.6000 ;
	    RECT 1451.4000 671.4000 1452.6000 672.6000 ;
	    RECT 1449.0000 647.4000 1450.2001 648.6000 ;
	    RECT 1444.2001 641.4000 1445.4000 642.6000 ;
	    RECT 1441.8000 635.4000 1443.0000 636.6000 ;
	    RECT 1437.0000 623.4000 1438.2001 624.6000 ;
	    RECT 1429.8000 617.4000 1431.0000 618.6000 ;
	    RECT 1427.4000 614.4000 1428.6000 615.6000 ;
	    RECT 1437.0000 614.4000 1438.2001 615.6000 ;
	    RECT 1422.6000 593.4000 1423.8000 594.6000 ;
	    RECT 1417.8000 581.4000 1419.0000 582.6000 ;
	    RECT 1420.2001 575.4000 1421.4000 576.6000 ;
	    RECT 1420.3500 555.6000 1421.2500 575.4000 ;
	    RECT 1427.5500 558.6000 1428.4501 614.4000 ;
	    RECT 1434.6000 593.4000 1435.8000 594.6000 ;
	    RECT 1434.7500 588.6000 1435.6500 593.4000 ;
	    RECT 1434.6000 587.4000 1435.8000 588.6000 ;
	    RECT 1432.2001 584.4000 1433.4000 585.6000 ;
	    RECT 1425.0000 557.4000 1426.2001 558.6000 ;
	    RECT 1427.4000 557.4000 1428.6000 558.6000 ;
	    RECT 1417.8000 554.4000 1419.0000 555.6000 ;
	    RECT 1420.2001 554.4000 1421.4000 555.6000 ;
	    RECT 1417.9501 552.6000 1418.8500 554.4000 ;
	    RECT 1417.8000 551.4000 1419.0000 552.6000 ;
	    RECT 1422.6000 551.4000 1423.8000 552.6000 ;
	    RECT 1422.7500 546.6000 1423.6500 551.4000 ;
	    RECT 1422.6000 545.4000 1423.8000 546.6000 ;
	    RECT 1425.1500 540.6000 1426.0500 557.4000 ;
	    RECT 1427.5500 555.6000 1428.4501 557.4000 ;
	    RECT 1427.4000 554.4000 1428.6000 555.6000 ;
	    RECT 1425.0000 539.4000 1426.2001 540.6000 ;
	    RECT 1415.4000 503.4000 1416.6000 504.6000 ;
	    RECT 1415.5500 495.6000 1416.4501 503.4000 ;
	    RECT 1420.2001 497.4000 1421.4000 498.6000 ;
	    RECT 1425.1500 495.6000 1426.0500 539.4000 ;
	    RECT 1415.4000 494.4000 1416.6000 495.6000 ;
	    RECT 1425.0000 494.4000 1426.2001 495.6000 ;
	    RECT 1422.6000 492.4500 1423.8000 492.6000 ;
	    RECT 1427.4000 492.4500 1428.6000 492.6000 ;
	    RECT 1422.6000 491.5500 1428.6000 492.4500 ;
	    RECT 1422.6000 491.4000 1423.8000 491.5500 ;
	    RECT 1425.1500 468.6000 1426.0500 491.5500 ;
	    RECT 1427.4000 491.4000 1428.6000 491.5500 ;
	    RECT 1415.4000 467.4000 1416.6000 468.6000 ;
	    RECT 1417.8000 467.4000 1419.0000 468.6000 ;
	    RECT 1425.0000 467.4000 1426.2001 468.6000 ;
	    RECT 1415.5500 435.6000 1416.4501 467.4000 ;
	    RECT 1417.9501 444.6000 1418.8500 467.4000 ;
	    RECT 1420.2001 464.4000 1421.4000 465.6000 ;
	    RECT 1420.3500 456.6000 1421.2500 464.4000 ;
	    RECT 1420.2001 455.4000 1421.4000 456.6000 ;
	    RECT 1417.8000 443.4000 1419.0000 444.6000 ;
	    RECT 1420.3500 441.6000 1421.2500 455.4000 ;
	    RECT 1420.2001 440.4000 1421.4000 441.6000 ;
	    RECT 1415.4000 434.4000 1416.6000 435.6000 ;
	    RECT 1427.4000 434.4000 1428.6000 435.6000 ;
	    RECT 1420.2001 431.4000 1421.4000 432.6000 ;
	    RECT 1420.3500 414.6000 1421.2500 431.4000 ;
	    RECT 1420.2001 413.4000 1421.4000 414.6000 ;
	    RECT 1417.8000 380.4000 1419.0000 381.6000 ;
	    RECT 1417.9501 336.6000 1418.8500 380.4000 ;
	    RECT 1420.3500 342.4500 1421.2500 413.4000 ;
	    RECT 1425.0000 404.4000 1426.2001 405.6000 ;
	    RECT 1422.6000 401.4000 1423.8000 402.6000 ;
	    RECT 1422.7500 396.6000 1423.6500 401.4000 ;
	    RECT 1422.6000 395.4000 1423.8000 396.6000 ;
	    RECT 1422.7500 381.6000 1423.6500 395.4000 ;
	    RECT 1422.6000 380.4000 1423.8000 381.6000 ;
	    RECT 1425.1500 378.6000 1426.0500 404.4000 ;
	    RECT 1425.0000 377.4000 1426.2001 378.6000 ;
	    RECT 1427.5500 345.6000 1428.4501 434.4000 ;
	    RECT 1432.3500 363.4500 1433.2500 584.4000 ;
	    RECT 1434.6000 528.4500 1435.8000 528.6000 ;
	    RECT 1437.1500 528.4500 1438.0500 614.4000 ;
	    RECT 1434.6000 527.5500 1438.0500 528.4500 ;
	    RECT 1434.6000 527.4000 1435.8000 527.5500 ;
	    RECT 1434.6000 524.4000 1435.8000 525.6000 ;
	    RECT 1434.7500 522.6000 1435.6500 524.4000 ;
	    RECT 1434.6000 521.4000 1435.8000 522.6000 ;
	    RECT 1441.9501 495.6000 1442.8500 635.4000 ;
	    RECT 1449.1500 588.6000 1450.0500 647.4000 ;
	    RECT 1449.0000 587.4000 1450.2001 588.6000 ;
	    RECT 1446.6000 554.4000 1447.8000 555.6000 ;
	    RECT 1446.7500 531.6000 1447.6500 554.4000 ;
	    RECT 1446.6000 530.4000 1447.8000 531.6000 ;
	    RECT 1444.2001 497.4000 1445.4000 498.6000 ;
	    RECT 1441.8000 494.4000 1443.0000 495.6000 ;
	    RECT 1437.0000 437.4000 1438.2001 438.6000 ;
	    RECT 1437.1500 402.6000 1438.0500 437.4000 ;
	    RECT 1444.3500 435.6000 1445.2500 497.4000 ;
	    RECT 1446.7500 471.6000 1447.6500 530.4000 ;
	    RECT 1449.1500 528.6000 1450.0500 587.4000 ;
	    RECT 1451.5500 576.6000 1452.4501 671.4000 ;
	    RECT 1453.9501 648.6000 1454.8500 677.4000 ;
	    RECT 1453.8000 647.4000 1455.0000 648.6000 ;
	    RECT 1451.4000 575.4000 1452.6000 576.6000 ;
	    RECT 1456.2001 557.4000 1457.4000 558.6000 ;
	    RECT 1453.8000 551.4000 1455.0000 552.6000 ;
	    RECT 1453.9501 534.4500 1454.8500 551.4000 ;
	    RECT 1451.5500 533.5500 1454.8500 534.4500 ;
	    RECT 1449.0000 527.4000 1450.2001 528.6000 ;
	    RECT 1449.0000 473.4000 1450.2001 474.6000 ;
	    RECT 1446.6000 470.4000 1447.8000 471.6000 ;
	    RECT 1449.1500 468.6000 1450.0500 473.4000 ;
	    RECT 1449.0000 467.4000 1450.2001 468.6000 ;
	    RECT 1444.2001 434.4000 1445.4000 435.6000 ;
	    RECT 1444.2001 431.4000 1445.4000 432.6000 ;
	    RECT 1439.4000 407.4000 1440.6000 408.6000 ;
	    RECT 1439.5500 402.6000 1440.4501 407.4000 ;
	    RECT 1434.6000 401.4000 1435.8000 402.6000 ;
	    RECT 1437.0000 401.4000 1438.2001 402.6000 ;
	    RECT 1439.4000 401.4000 1440.6000 402.6000 ;
	    RECT 1434.7500 381.4500 1435.6500 401.4000 ;
	    RECT 1434.7500 380.5500 1438.0500 381.4500 ;
	    RECT 1434.6000 377.4000 1435.8000 378.6000 ;
	    RECT 1429.9501 362.5500 1433.2500 363.4500 ;
	    RECT 1427.4000 344.4000 1428.6000 345.6000 ;
	    RECT 1422.6000 342.4500 1423.8000 342.6000 ;
	    RECT 1420.3500 341.5500 1423.8000 342.4500 ;
	    RECT 1422.6000 341.4000 1423.8000 341.5500 ;
	    RECT 1417.8000 335.4000 1419.0000 336.6000 ;
	    RECT 1422.7500 321.6000 1423.6500 341.4000 ;
	    RECT 1422.6000 320.4000 1423.8000 321.6000 ;
	    RECT 1427.4000 317.4000 1428.6000 318.6000 ;
	    RECT 1420.2001 314.4000 1421.4000 315.6000 ;
	    RECT 1429.9501 315.4500 1430.8500 362.5500 ;
	    RECT 1432.2001 359.4000 1433.4000 360.6000 ;
	    RECT 1427.5500 314.5500 1430.8500 315.4500 ;
	    RECT 1420.3500 282.6000 1421.2500 314.4000 ;
	    RECT 1420.2001 281.4000 1421.4000 282.6000 ;
	    RECT 1420.3500 279.6000 1421.2500 281.4000 ;
	    RECT 1420.2001 278.4000 1421.4000 279.6000 ;
	    RECT 1417.8000 245.4000 1419.0000 246.6000 ;
	    RECT 1408.2001 239.4000 1409.4000 240.6000 ;
	    RECT 1413.0000 239.4000 1414.2001 240.6000 ;
	    RECT 1408.3500 228.6000 1409.2500 239.4000 ;
	    RECT 1405.8000 227.4000 1407.0000 228.6000 ;
	    RECT 1408.2001 227.4000 1409.4000 228.6000 ;
	    RECT 1415.4000 221.4000 1416.6000 222.6000 ;
	    RECT 1408.2001 203.4000 1409.4000 204.6000 ;
	    RECT 1408.3500 198.6000 1409.2500 203.4000 ;
	    RECT 1398.6000 197.4000 1399.8000 198.6000 ;
	    RECT 1401.0000 197.4000 1402.2001 198.6000 ;
	    RECT 1408.2001 197.4000 1409.4000 198.6000 ;
	    RECT 1398.7500 195.6000 1399.6500 197.4000 ;
	    RECT 1398.6000 194.4000 1399.8000 195.6000 ;
	    RECT 1396.2001 191.4000 1397.4000 192.6000 ;
	    RECT 1396.3500 168.6000 1397.2500 191.4000 ;
	    RECT 1401.1500 180.6000 1402.0500 197.4000 ;
	    RECT 1401.0000 179.4000 1402.2001 180.6000 ;
	    RECT 1398.6000 173.4000 1399.8000 174.6000 ;
	    RECT 1398.7500 171.6000 1399.6500 173.4000 ;
	    RECT 1398.6000 170.4000 1399.8000 171.6000 ;
	    RECT 1396.2001 167.4000 1397.4000 168.6000 ;
	    RECT 1396.3500 150.6000 1397.2500 167.4000 ;
	    RECT 1405.8000 158.4000 1407.0000 159.6000 ;
	    RECT 1396.2001 149.4000 1397.4000 150.6000 ;
	    RECT 1391.4000 131.4000 1392.6000 132.6000 ;
	    RECT 1405.9501 126.6000 1406.8500 158.4000 ;
	    RECT 1413.0000 143.4000 1414.2001 144.6000 ;
	    RECT 1413.1500 141.6000 1414.0500 143.4000 ;
	    RECT 1413.0000 140.4000 1414.2001 141.6000 ;
	    RECT 1405.8000 125.4000 1407.0000 126.6000 ;
	    RECT 1384.2001 107.4000 1385.4000 108.6000 ;
	    RECT 1415.5500 102.6000 1416.4501 221.4000 ;
	    RECT 1417.9501 195.6000 1418.8500 245.4000 ;
	    RECT 1420.3500 228.6000 1421.2500 278.4000 ;
	    RECT 1420.2001 227.4000 1421.4000 228.6000 ;
	    RECT 1417.8000 194.4000 1419.0000 195.6000 ;
	    RECT 1425.0000 164.4000 1426.2001 165.6000 ;
	    RECT 1420.2001 158.4000 1421.4000 159.6000 ;
	    RECT 1420.3500 150.4500 1421.2500 158.4000 ;
	    RECT 1422.6000 150.4500 1423.8000 150.6000 ;
	    RECT 1420.3500 149.5500 1423.8000 150.4500 ;
	    RECT 1422.6000 149.4000 1423.8000 149.5500 ;
	    RECT 1425.1500 144.6000 1426.0500 164.4000 ;
	    RECT 1425.0000 143.4000 1426.2001 144.6000 ;
	    RECT 1420.2001 134.4000 1421.4000 135.6000 ;
	    RECT 1420.3500 132.6000 1421.2500 134.4000 ;
	    RECT 1420.2001 131.4000 1421.4000 132.6000 ;
	    RECT 1415.4000 101.4000 1416.6000 102.6000 ;
	    RECT 1401.0000 89.4000 1402.2001 90.6000 ;
	    RECT 1401.1500 84.6000 1402.0500 89.4000 ;
	    RECT 1427.5500 84.6000 1428.4501 314.5500 ;
	    RECT 1429.8000 311.4000 1431.0000 312.6000 ;
	    RECT 1429.8000 287.4000 1431.0000 288.6000 ;
	    RECT 1429.9501 282.6000 1430.8500 287.4000 ;
	    RECT 1429.8000 281.4000 1431.0000 282.6000 ;
	    RECT 1432.3500 258.6000 1433.2500 359.4000 ;
	    RECT 1437.1500 312.6000 1438.0500 380.5500 ;
	    RECT 1439.4000 374.4000 1440.6000 375.6000 ;
	    RECT 1439.5500 372.6000 1440.4501 374.4000 ;
	    RECT 1439.4000 371.4000 1440.6000 372.6000 ;
	    RECT 1441.8000 338.4000 1443.0000 339.6000 ;
	    RECT 1441.9501 330.6000 1442.8500 338.4000 ;
	    RECT 1441.8000 329.4000 1443.0000 330.6000 ;
	    RECT 1439.4000 314.4000 1440.6000 315.6000 ;
	    RECT 1437.0000 311.4000 1438.2001 312.6000 ;
	    RECT 1439.5500 276.6000 1440.4501 314.4000 ;
	    RECT 1441.8000 293.4000 1443.0000 294.6000 ;
	    RECT 1441.9501 282.6000 1442.8500 293.4000 ;
	    RECT 1441.8000 281.4000 1443.0000 282.6000 ;
	    RECT 1439.4000 275.4000 1440.6000 276.6000 ;
	    RECT 1441.8000 263.4000 1443.0000 264.6000 ;
	    RECT 1434.6000 260.4000 1435.8000 261.6000 ;
	    RECT 1432.2001 257.4000 1433.4000 258.6000 ;
	    RECT 1434.7500 234.6000 1435.6500 260.4000 ;
	    RECT 1441.9501 258.6000 1442.8500 263.4000 ;
	    RECT 1437.0000 257.4000 1438.2001 258.6000 ;
	    RECT 1441.8000 257.4000 1443.0000 258.6000 ;
	    RECT 1437.1500 252.6000 1438.0500 257.4000 ;
	    RECT 1437.0000 251.4000 1438.2001 252.6000 ;
	    RECT 1434.6000 233.4000 1435.8000 234.6000 ;
	    RECT 1429.8000 225.4500 1431.0000 225.6000 ;
	    RECT 1429.8000 224.5500 1435.6500 225.4500 ;
	    RECT 1429.8000 224.4000 1431.0000 224.5500 ;
	    RECT 1434.7500 222.6000 1435.6500 224.5500 ;
	    RECT 1444.3500 222.6000 1445.2500 431.4000 ;
	    RECT 1446.6000 398.4000 1447.8000 399.6000 ;
	    RECT 1446.7500 375.6000 1447.6500 398.4000 ;
	    RECT 1449.0000 380.4000 1450.2001 381.6000 ;
	    RECT 1446.6000 374.4000 1447.8000 375.6000 ;
	    RECT 1446.6000 335.4000 1447.8000 336.6000 ;
	    RECT 1446.7500 318.6000 1447.6500 335.4000 ;
	    RECT 1446.6000 317.4000 1447.8000 318.6000 ;
	    RECT 1449.1500 306.6000 1450.0500 380.4000 ;
	    RECT 1451.5500 345.6000 1452.4501 533.5500 ;
	    RECT 1453.8000 497.4000 1455.0000 498.6000 ;
	    RECT 1453.8000 491.4000 1455.0000 492.6000 ;
	    RECT 1453.9501 471.6000 1454.8500 491.4000 ;
	    RECT 1453.8000 470.4000 1455.0000 471.6000 ;
	    RECT 1453.9501 420.6000 1454.8500 470.4000 ;
	    RECT 1453.8000 419.4000 1455.0000 420.6000 ;
	    RECT 1456.3500 402.6000 1457.2500 557.4000 ;
	    RECT 1458.7500 432.6000 1459.6500 701.4000 ;
	    RECT 1461.1500 675.6000 1462.0500 731.4000 ;
	    RECT 1463.5500 702.6000 1464.4501 794.4000 ;
	    RECT 1463.4000 701.4000 1464.6000 702.6000 ;
	    RECT 1468.3500 678.6000 1469.2500 809.4000 ;
	    RECT 1468.2001 677.4000 1469.4000 678.6000 ;
	    RECT 1461.0000 674.4000 1462.2001 675.6000 ;
	    RECT 1463.4000 650.4000 1464.6000 651.6000 ;
	    RECT 1463.5500 648.6000 1464.4501 650.4000 ;
	    RECT 1463.4000 647.4000 1464.6000 648.6000 ;
	    RECT 1461.0000 644.4000 1462.2001 645.6000 ;
	    RECT 1461.1500 642.6000 1462.0500 644.4000 ;
	    RECT 1461.0000 641.4000 1462.2001 642.6000 ;
	    RECT 1463.4000 590.4000 1464.6000 591.6000 ;
	    RECT 1463.5500 588.6000 1464.4501 590.4000 ;
	    RECT 1463.4000 587.4000 1464.6000 588.6000 ;
	    RECT 1461.0000 584.4000 1462.2001 585.6000 ;
	    RECT 1461.1500 582.6000 1462.0500 584.4000 ;
	    RECT 1461.0000 581.4000 1462.2001 582.6000 ;
	    RECT 1463.5500 546.6000 1464.4501 587.4000 ;
	    RECT 1463.4000 545.4000 1464.6000 546.6000 ;
	    RECT 1465.8000 530.4000 1467.0000 531.6000 ;
	    RECT 1468.2001 530.4000 1469.4000 531.6000 ;
	    RECT 1461.0000 527.4000 1462.2001 528.6000 ;
	    RECT 1461.1500 522.6000 1462.0500 527.4000 ;
	    RECT 1465.9501 525.6000 1466.8500 530.4000 ;
	    RECT 1465.8000 524.4000 1467.0000 525.6000 ;
	    RECT 1461.0000 521.4000 1462.2001 522.6000 ;
	    RECT 1461.1500 495.6000 1462.0500 521.4000 ;
	    RECT 1461.0000 494.4000 1462.2001 495.6000 ;
	    RECT 1468.3500 492.6000 1469.2500 530.4000 ;
	    RECT 1468.2001 491.4000 1469.4000 492.6000 ;
	    RECT 1468.2001 446.4000 1469.4000 447.6000 ;
	    RECT 1461.0000 440.4000 1462.2001 441.6000 ;
	    RECT 1458.6000 431.4000 1459.8000 432.6000 ;
	    RECT 1461.1500 420.6000 1462.0500 440.4000 ;
	    RECT 1465.8000 435.4500 1467.0000 435.6000 ;
	    RECT 1463.5500 434.5500 1467.0000 435.4500 ;
	    RECT 1461.0000 419.4000 1462.2001 420.6000 ;
	    RECT 1461.0000 407.4000 1462.2001 408.6000 ;
	    RECT 1461.1500 402.6000 1462.0500 407.4000 ;
	    RECT 1456.2001 401.4000 1457.4000 402.6000 ;
	    RECT 1461.0000 401.4000 1462.2001 402.6000 ;
	    RECT 1461.0000 377.4000 1462.2001 378.6000 ;
	    RECT 1458.6000 347.4000 1459.8000 348.6000 ;
	    RECT 1458.7500 345.6000 1459.6500 347.4000 ;
	    RECT 1451.4000 344.4000 1452.6000 345.6000 ;
	    RECT 1458.6000 344.4000 1459.8000 345.6000 ;
	    RECT 1451.4000 341.4000 1452.6000 342.6000 ;
	    RECT 1449.0000 305.4000 1450.2001 306.6000 ;
	    RECT 1451.5500 303.4500 1452.4501 341.4000 ;
	    RECT 1461.1500 336.6000 1462.0500 377.4000 ;
	    RECT 1463.5500 342.6000 1464.4501 434.5500 ;
	    RECT 1465.8000 434.4000 1467.0000 434.5500 ;
	    RECT 1465.8000 404.4000 1467.0000 405.6000 ;
	    RECT 1463.4000 341.4000 1464.6000 342.6000 ;
	    RECT 1461.0000 335.4000 1462.2001 336.6000 ;
	    RECT 1461.1500 318.6000 1462.0500 335.4000 ;
	    RECT 1461.0000 317.4000 1462.2001 318.6000 ;
	    RECT 1456.2001 314.4000 1457.4000 315.6000 ;
	    RECT 1463.4000 314.4000 1464.6000 315.6000 ;
	    RECT 1453.8000 311.4000 1455.0000 312.6000 ;
	    RECT 1456.3500 306.6000 1457.2500 314.4000 ;
	    RECT 1458.6000 311.4000 1459.8000 312.6000 ;
	    RECT 1453.8000 305.4000 1455.0000 306.6000 ;
	    RECT 1456.2001 305.4000 1457.4000 306.6000 ;
	    RECT 1449.1500 302.5500 1452.4501 303.4500 ;
	    RECT 1446.6000 287.4000 1447.8000 288.6000 ;
	    RECT 1446.7500 270.6000 1447.6500 287.4000 ;
	    RECT 1446.6000 269.4000 1447.8000 270.6000 ;
	    RECT 1429.8000 221.4000 1431.0000 222.6000 ;
	    RECT 1434.6000 221.4000 1435.8000 222.6000 ;
	    RECT 1444.2001 221.4000 1445.4000 222.6000 ;
	    RECT 1446.6000 221.4000 1447.8000 222.6000 ;
	    RECT 1429.9501 219.6000 1430.8500 221.4000 ;
	    RECT 1449.1500 219.6000 1450.0500 302.5500 ;
	    RECT 1453.9501 288.6000 1454.8500 305.4000 ;
	    RECT 1456.2001 299.4000 1457.4000 300.6000 ;
	    RECT 1451.4000 287.4000 1452.6000 288.6000 ;
	    RECT 1453.8000 287.4000 1455.0000 288.6000 ;
	    RECT 1451.5500 285.6000 1452.4501 287.4000 ;
	    RECT 1451.4000 284.4000 1452.6000 285.6000 ;
	    RECT 1429.8000 218.4000 1431.0000 219.6000 ;
	    RECT 1449.0000 218.4000 1450.2001 219.6000 ;
	    RECT 1449.1500 216.6000 1450.0500 218.4000 ;
	    RECT 1434.6000 215.4000 1435.8000 216.6000 ;
	    RECT 1449.0000 215.4000 1450.2001 216.6000 ;
	    RECT 1434.7500 174.6000 1435.6500 215.4000 ;
	    RECT 1444.2001 203.4000 1445.4000 204.6000 ;
	    RECT 1451.4000 203.4000 1452.6000 204.6000 ;
	    RECT 1444.3500 201.6000 1445.2500 203.4000 ;
	    RECT 1444.2001 200.4000 1445.4000 201.6000 ;
	    RECT 1451.5500 198.6000 1452.4501 203.4000 ;
	    RECT 1451.4000 197.4000 1452.6000 198.6000 ;
	    RECT 1444.2001 194.4000 1445.4000 195.6000 ;
	    RECT 1453.8000 194.4000 1455.0000 195.6000 ;
	    RECT 1429.8000 173.4000 1431.0000 174.6000 ;
	    RECT 1434.6000 173.4000 1435.8000 174.6000 ;
	    RECT 1441.8000 173.4000 1443.0000 174.6000 ;
	    RECT 1429.9501 168.6000 1430.8500 173.4000 ;
	    RECT 1444.3500 168.6000 1445.2500 194.4000 ;
	    RECT 1453.9501 192.6000 1454.8500 194.4000 ;
	    RECT 1449.0000 191.4000 1450.2001 192.6000 ;
	    RECT 1453.8000 191.4000 1455.0000 192.6000 ;
	    RECT 1429.8000 167.4000 1431.0000 168.6000 ;
	    RECT 1444.2001 167.4000 1445.4000 168.6000 ;
	    RECT 1449.1500 162.6000 1450.0500 191.4000 ;
	    RECT 1453.9501 162.6000 1454.8500 191.4000 ;
	    RECT 1456.3500 168.6000 1457.2500 299.4000 ;
	    RECT 1463.5500 294.6000 1464.4501 314.4000 ;
	    RECT 1463.4000 293.4000 1464.6000 294.6000 ;
	    RECT 1465.9501 291.6000 1466.8500 404.4000 ;
	    RECT 1468.3500 348.6000 1469.2500 446.4000 ;
	    RECT 1470.7500 438.6000 1471.6500 1049.4000 ;
	    RECT 1475.4000 1046.4000 1476.6000 1047.6000 ;
	    RECT 1473.0000 950.4000 1474.2001 951.6000 ;
	    RECT 1473.1500 930.6000 1474.0500 950.4000 ;
	    RECT 1473.0000 929.4000 1474.2001 930.6000 ;
	    RECT 1475.5500 870.6000 1476.4501 1046.4000 ;
	    RECT 1477.9501 930.6000 1478.8500 1058.4000 ;
	    RECT 1480.2001 1056.3000 1481.4000 1073.7001 ;
	    RECT 1482.7500 1068.6000 1483.6500 1100.4000 ;
	    RECT 1489.9501 1080.6000 1490.8500 1157.4000 ;
	    RECT 1492.3500 1101.6000 1493.2500 1277.4000 ;
	    RECT 1509.1500 1275.6000 1510.0500 1283.4000 ;
	    RECT 1509.0000 1274.4000 1510.2001 1275.6000 ;
	    RECT 1513.8000 1253.4000 1515.0000 1254.6000 ;
	    RECT 1497.0000 1247.4000 1498.2001 1248.6000 ;
	    RECT 1494.6000 1241.4000 1495.8000 1242.6000 ;
	    RECT 1494.7500 1164.6000 1495.6500 1241.4000 ;
	    RECT 1494.6000 1163.4000 1495.8000 1164.6000 ;
	    RECT 1494.6000 1109.4000 1495.8000 1110.6000 ;
	    RECT 1492.2001 1100.4000 1493.4000 1101.6000 ;
	    RECT 1489.8000 1079.4000 1491.0000 1080.6000 ;
	    RECT 1482.6000 1067.4000 1483.8000 1068.6000 ;
	    RECT 1482.6000 1061.4000 1483.8000 1062.6000 ;
	    RECT 1485.0000 1056.3000 1486.2001 1073.7001 ;
	    RECT 1487.4000 1056.3000 1488.6000 1076.7001 ;
	    RECT 1489.8000 1056.3000 1491.0000 1076.7001 ;
	    RECT 1492.2001 1064.4000 1493.4000 1065.6000 ;
	    RECT 1492.3500 1047.6000 1493.2500 1064.4000 ;
	    RECT 1492.2001 1046.4000 1493.4000 1047.6000 ;
	    RECT 1489.8000 1025.4000 1491.0000 1026.6000 ;
	    RECT 1489.9501 1005.6000 1490.8500 1025.4000 ;
	    RECT 1492.2001 1007.4000 1493.4000 1008.6000 ;
	    RECT 1492.3500 1005.6000 1493.2500 1007.4000 ;
	    RECT 1489.8000 1004.4000 1491.0000 1005.6000 ;
	    RECT 1492.2001 1004.4000 1493.4000 1005.6000 ;
	    RECT 1494.7500 1005.4500 1495.6500 1109.4000 ;
	    RECT 1497.1500 1080.4501 1498.0500 1247.4000 ;
	    RECT 1513.9501 1242.6000 1514.8500 1253.4000 ;
	    RECT 1513.8000 1241.4000 1515.0000 1242.6000 ;
	    RECT 1509.0000 1211.4000 1510.2001 1212.6000 ;
	    RECT 1499.4000 1176.3000 1500.6000 1196.7001 ;
	    RECT 1501.8000 1176.3000 1503.0000 1196.7001 ;
	    RECT 1504.2001 1176.3000 1505.4000 1196.7001 ;
	    RECT 1506.6000 1176.3000 1507.8000 1193.7001 ;
	    RECT 1509.1500 1182.6000 1510.0500 1211.4000 ;
	    RECT 1518.7500 1206.6000 1519.6500 1325.4000 ;
	    RECT 1521.1500 1266.6000 1522.0500 1367.4000 ;
	    RECT 1523.5500 1362.6000 1524.4501 1370.4000 ;
	    RECT 1545.0000 1367.4000 1546.2001 1368.6000 ;
	    RECT 1523.4000 1361.4000 1524.6000 1362.6000 ;
	    RECT 1542.6000 1355.4000 1543.8000 1356.6000 ;
	    RECT 1542.7500 1341.6000 1543.6500 1355.4000 ;
	    RECT 1540.2001 1340.4000 1541.4000 1341.6000 ;
	    RECT 1542.6000 1340.4000 1543.8000 1341.6000 ;
	    RECT 1540.3500 1338.6000 1541.2500 1340.4000 ;
	    RECT 1540.2001 1337.4000 1541.4000 1338.6000 ;
	    RECT 1540.2001 1334.4000 1541.4000 1335.6000 ;
	    RECT 1523.4000 1280.4000 1524.6000 1281.6000 ;
	    RECT 1521.0000 1265.4000 1522.2001 1266.6000 ;
	    RECT 1521.0000 1260.4501 1522.2001 1260.6000 ;
	    RECT 1523.5500 1260.4501 1524.4501 1280.4000 ;
	    RECT 1540.3500 1278.6000 1541.2500 1334.4000 ;
	    RECT 1542.6000 1325.4000 1543.8000 1326.6000 ;
	    RECT 1540.2001 1277.4000 1541.4000 1278.6000 ;
	    RECT 1537.8000 1274.4000 1539.0000 1275.6000 ;
	    RECT 1521.0000 1259.5500 1524.4501 1260.4501 ;
	    RECT 1521.0000 1259.4000 1522.2001 1259.5500 ;
	    RECT 1530.6000 1253.4000 1531.8000 1254.6000 ;
	    RECT 1530.7500 1248.6000 1531.6500 1253.4000 ;
	    RECT 1530.6000 1247.4000 1531.8000 1248.6000 ;
	    RECT 1530.6000 1244.4000 1531.8000 1245.6000 ;
	    RECT 1530.7500 1242.6000 1531.6500 1244.4000 ;
	    RECT 1530.6000 1241.4000 1531.8000 1242.6000 ;
	    RECT 1528.2001 1235.4000 1529.4000 1236.6000 ;
	    RECT 1525.8000 1215.3000 1527.0000 1223.7001 ;
	    RECT 1528.3500 1221.6000 1529.2500 1235.4000 ;
	    RECT 1528.2001 1220.4000 1529.4000 1221.6000 ;
	    RECT 1523.4000 1211.4000 1524.6000 1212.6000 ;
	    RECT 1530.6000 1209.3000 1531.8000 1226.7001 ;
	    RECT 1535.4000 1217.4000 1536.6000 1218.6000 ;
	    RECT 1535.5500 1212.6000 1536.4501 1217.4000 ;
	    RECT 1535.4000 1211.4000 1536.6000 1212.6000 ;
	    RECT 1518.6000 1205.4000 1519.8000 1206.6000 ;
	    RECT 1523.4000 1205.4000 1524.6000 1206.6000 ;
	    RECT 1535.4000 1205.4000 1536.6000 1206.6000 ;
	    RECT 1523.5500 1200.6000 1524.4501 1205.4000 ;
	    RECT 1523.4000 1199.4000 1524.6000 1200.6000 ;
	    RECT 1530.6000 1199.4000 1531.8000 1200.6000 ;
	    RECT 1509.0000 1181.4000 1510.2001 1182.6000 ;
	    RECT 1509.0000 1178.4000 1510.2001 1179.6000 ;
	    RECT 1501.8000 1173.4501 1503.0000 1173.6000 ;
	    RECT 1501.8000 1172.5500 1505.2500 1173.4501 ;
	    RECT 1501.8000 1172.4000 1503.0000 1172.5500 ;
	    RECT 1504.3500 1170.6000 1505.2500 1172.5500 ;
	    RECT 1506.6000 1172.4000 1507.8000 1173.6000 ;
	    RECT 1504.2001 1169.4000 1505.4000 1170.6000 ;
	    RECT 1501.8000 1154.4000 1503.0000 1155.6000 ;
	    RECT 1506.7500 1155.4501 1507.6500 1172.4000 ;
	    RECT 1509.1500 1170.6000 1510.0500 1178.4000 ;
	    RECT 1511.4000 1176.3000 1512.6000 1193.7001 ;
	    RECT 1513.8000 1193.4000 1515.0000 1194.6000 ;
	    RECT 1513.9501 1182.6000 1514.8500 1193.4000 ;
	    RECT 1513.8000 1181.4000 1515.0000 1182.6000 ;
	    RECT 1513.8000 1175.4000 1515.0000 1176.6000 ;
	    RECT 1516.2001 1176.3000 1517.4000 1193.7001 ;
	    RECT 1518.6000 1176.3000 1519.8000 1196.7001 ;
	    RECT 1521.0000 1176.3000 1522.2001 1196.7001 ;
	    RECT 1523.5500 1185.6000 1524.4501 1199.4000 ;
	    RECT 1530.7500 1197.4501 1531.6500 1199.4000 ;
	    RECT 1530.7500 1196.5500 1534.0500 1197.4501 ;
	    RECT 1530.6000 1193.4000 1531.8000 1194.6000 ;
	    RECT 1530.7500 1188.6000 1531.6500 1193.4000 ;
	    RECT 1530.6000 1187.4000 1531.8000 1188.6000 ;
	    RECT 1523.4000 1184.4000 1524.6000 1185.6000 ;
	    RECT 1533.1500 1176.6000 1534.0500 1196.5500 ;
	    RECT 1523.4000 1175.4000 1524.6000 1176.6000 ;
	    RECT 1533.0000 1175.4000 1534.2001 1176.6000 ;
	    RECT 1513.9501 1170.6000 1514.8500 1175.4000 ;
	    RECT 1509.0000 1169.4000 1510.2001 1170.6000 ;
	    RECT 1513.8000 1169.4000 1515.0000 1170.6000 ;
	    RECT 1509.0000 1157.4000 1510.2001 1158.6000 ;
	    RECT 1506.7500 1154.5500 1510.0500 1155.4501 ;
	    RECT 1501.9501 1146.4501 1502.8500 1154.4000 ;
	    RECT 1504.2001 1146.4501 1505.4000 1146.6000 ;
	    RECT 1501.9501 1145.5500 1505.4000 1146.4501 ;
	    RECT 1504.2001 1145.4000 1505.4000 1145.5500 ;
	    RECT 1501.8000 1127.4000 1503.0000 1128.6000 ;
	    RECT 1501.9501 1104.4501 1502.8500 1127.4000 ;
	    RECT 1504.2001 1116.3000 1505.4000 1133.7001 ;
	    RECT 1499.5500 1103.5500 1502.8500 1104.4501 ;
	    RECT 1499.5500 1095.6000 1500.4501 1103.5500 ;
	    RECT 1509.1500 1101.6000 1510.0500 1154.5500 ;
	    RECT 1511.4000 1146.3000 1512.6000 1166.7001 ;
	    RECT 1513.8000 1146.3000 1515.0000 1166.7001 ;
	    RECT 1516.2001 1149.3000 1517.4000 1166.7001 ;
	    RECT 1518.6000 1163.4000 1519.8000 1164.6000 ;
	    RECT 1518.7500 1161.6000 1519.6500 1163.4000 ;
	    RECT 1518.6000 1160.4000 1519.8000 1161.6000 ;
	    RECT 1521.0000 1149.3000 1522.2001 1166.7001 ;
	    RECT 1523.5500 1164.6000 1524.4501 1175.4000 ;
	    RECT 1523.4000 1163.4000 1524.6000 1164.6000 ;
	    RECT 1523.5500 1140.6000 1524.4501 1163.4000 ;
	    RECT 1525.8000 1149.3000 1527.0000 1166.7001 ;
	    RECT 1528.2001 1146.3000 1529.4000 1166.7001 ;
	    RECT 1530.6000 1146.3000 1531.8000 1166.7001 ;
	    RECT 1533.0000 1146.3000 1534.2001 1166.7001 ;
	    RECT 1523.4000 1139.4000 1524.6000 1140.6000 ;
	    RECT 1528.2001 1139.4000 1529.4000 1140.6000 ;
	    RECT 1533.0000 1139.4000 1534.2001 1140.6000 ;
	    RECT 1513.8000 1124.4000 1515.0000 1125.6000 ;
	    RECT 1513.9501 1116.6000 1514.8500 1124.4000 ;
	    RECT 1513.8000 1115.4000 1515.0000 1116.6000 ;
	    RECT 1518.6000 1116.3000 1519.8000 1133.7001 ;
	    RECT 1521.0000 1121.4000 1522.2001 1122.6000 ;
	    RECT 1521.1500 1104.6000 1522.0500 1121.4000 ;
	    RECT 1523.4000 1119.3000 1524.6000 1127.7001 ;
	    RECT 1525.8000 1127.4000 1527.0000 1128.6000 ;
	    RECT 1525.9501 1125.6000 1526.8500 1127.4000 ;
	    RECT 1525.8000 1124.4000 1527.0000 1125.6000 ;
	    RECT 1528.3500 1122.4501 1529.2500 1139.4000 ;
	    RECT 1533.1500 1122.6000 1534.0500 1139.4000 ;
	    RECT 1525.9501 1121.5500 1529.2500 1122.4501 ;
	    RECT 1525.9501 1116.4501 1526.8500 1121.5500 ;
	    RECT 1533.0000 1121.4000 1534.2001 1122.6000 ;
	    RECT 1523.5500 1115.5500 1526.8500 1116.4501 ;
	    RECT 1521.0000 1103.4000 1522.2001 1104.6000 ;
	    RECT 1501.8000 1100.4000 1503.0000 1101.6000 ;
	    RECT 1509.0000 1100.4000 1510.2001 1101.6000 ;
	    RECT 1513.8000 1100.4000 1515.0000 1101.6000 ;
	    RECT 1499.4000 1094.4000 1500.6000 1095.6000 ;
	    RECT 1501.9501 1086.6000 1502.8500 1100.4000 ;
	    RECT 1504.2001 1097.4000 1505.4000 1098.6000 ;
	    RECT 1509.0000 1097.4000 1510.2001 1098.6000 ;
	    RECT 1504.3500 1092.6000 1505.2500 1097.4000 ;
	    RECT 1504.2001 1091.4000 1505.4000 1092.6000 ;
	    RECT 1501.8000 1085.4000 1503.0000 1086.6000 ;
	    RECT 1497.1500 1079.5500 1500.4501 1080.4501 ;
	    RECT 1497.0000 1076.4000 1498.2001 1077.6000 ;
	    RECT 1497.1500 1068.6000 1498.0500 1076.4000 ;
	    RECT 1497.0000 1067.4000 1498.2001 1068.6000 ;
	    RECT 1497.0000 1013.4000 1498.2001 1014.6000 ;
	    RECT 1497.1500 1008.6000 1498.0500 1013.4000 ;
	    RECT 1499.5500 1011.4500 1500.4501 1079.5500 ;
	    RECT 1504.2001 1079.4000 1505.4000 1080.6000 ;
	    RECT 1499.5500 1010.5500 1502.8500 1011.4500 ;
	    RECT 1497.0000 1007.4000 1498.2001 1008.6000 ;
	    RECT 1499.4000 1007.4000 1500.6000 1008.6000 ;
	    RECT 1494.7500 1004.5500 1498.0500 1005.4500 ;
	    RECT 1497.1500 1002.6000 1498.0500 1004.5500 ;
	    RECT 1499.5500 1002.6000 1500.4501 1007.4000 ;
	    RECT 1492.2001 1001.4000 1493.4000 1002.6000 ;
	    RECT 1497.0000 1001.4000 1498.2001 1002.6000 ;
	    RECT 1499.4000 1001.4000 1500.6000 1002.6000 ;
	    RECT 1492.3500 996.6000 1493.2500 1001.4000 ;
	    RECT 1492.2001 995.4000 1493.4000 996.6000 ;
	    RECT 1482.6000 980.4000 1483.8000 981.6000 ;
	    RECT 1482.7500 936.6000 1483.6500 980.4000 ;
	    RECT 1489.8000 977.4000 1491.0000 978.6000 ;
	    RECT 1482.6000 935.4000 1483.8000 936.6000 ;
	    RECT 1477.8000 930.4500 1479.0000 930.6000 ;
	    RECT 1477.8000 929.5500 1481.2500 930.4500 ;
	    RECT 1477.8000 929.4000 1479.0000 929.5500 ;
	    RECT 1477.8000 920.4000 1479.0000 921.6000 ;
	    RECT 1477.9501 912.6000 1478.8500 920.4000 ;
	    RECT 1477.8000 911.4000 1479.0000 912.6000 ;
	    RECT 1480.3500 894.6000 1481.2500 929.5500 ;
	    RECT 1482.7500 921.6000 1483.6500 935.4000 ;
	    RECT 1482.6000 920.4000 1483.8000 921.6000 ;
	    RECT 1485.0000 917.4000 1486.2001 918.6000 ;
	    RECT 1489.9501 915.6000 1490.8500 977.4000 ;
	    RECT 1492.3500 975.6000 1493.2500 995.4000 ;
	    RECT 1492.2001 974.4000 1493.4000 975.6000 ;
	    RECT 1499.4000 965.4000 1500.6000 966.6000 ;
	    RECT 1497.0000 923.4000 1498.2001 924.6000 ;
	    RECT 1492.2001 920.4000 1493.4000 921.6000 ;
	    RECT 1492.3500 918.6000 1493.2500 920.4000 ;
	    RECT 1492.2001 917.4000 1493.4000 918.6000 ;
	    RECT 1489.8000 914.4000 1491.0000 915.6000 ;
	    RECT 1480.2001 893.4000 1481.4000 894.6000 ;
	    RECT 1475.4000 869.4000 1476.6000 870.6000 ;
	    RECT 1475.4000 824.4000 1476.6000 825.6000 ;
	    RECT 1475.5500 807.6000 1476.4501 824.4000 ;
	    RECT 1475.4000 806.4000 1476.6000 807.6000 ;
	    RECT 1475.5500 708.6000 1476.4501 806.4000 ;
	    RECT 1492.2001 803.4000 1493.4000 804.6000 ;
	    RECT 1492.3500 801.6000 1493.2500 803.4000 ;
	    RECT 1492.2001 800.4000 1493.4000 801.6000 ;
	    RECT 1494.6000 797.4000 1495.8000 798.6000 ;
	    RECT 1487.4000 767.4000 1488.6000 768.6000 ;
	    RECT 1482.6000 764.4000 1483.8000 765.6000 ;
	    RECT 1482.7500 762.6000 1483.6500 764.4000 ;
	    RECT 1480.2001 761.4000 1481.4000 762.6000 ;
	    RECT 1482.6000 761.4000 1483.8000 762.6000 ;
	    RECT 1480.3500 741.6000 1481.2500 761.4000 ;
	    RECT 1485.0000 743.4000 1486.2001 744.6000 ;
	    RECT 1477.8000 740.4000 1479.0000 741.6000 ;
	    RECT 1480.2001 740.4000 1481.4000 741.6000 ;
	    RECT 1475.4000 707.4000 1476.6000 708.6000 ;
	    RECT 1475.5500 696.6000 1476.4501 707.4000 ;
	    RECT 1477.9501 705.6000 1478.8500 740.4000 ;
	    RECT 1485.1500 738.6000 1486.0500 743.4000 ;
	    RECT 1487.5500 738.6000 1488.4501 767.4000 ;
	    RECT 1492.2001 761.4000 1493.4000 762.6000 ;
	    RECT 1492.3500 759.6000 1493.2500 761.4000 ;
	    RECT 1492.2001 758.4000 1493.4000 759.6000 ;
	    RECT 1485.0000 737.4000 1486.2001 738.6000 ;
	    RECT 1487.4000 737.4000 1488.6000 738.6000 ;
	    RECT 1492.2001 734.4000 1493.4000 735.6000 ;
	    RECT 1492.3500 732.6000 1493.2500 734.4000 ;
	    RECT 1492.2001 731.4000 1493.4000 732.6000 ;
	    RECT 1480.2001 710.4000 1481.4000 711.6000 ;
	    RECT 1480.3500 708.6000 1481.2500 710.4000 ;
	    RECT 1480.2001 707.4000 1481.4000 708.6000 ;
	    RECT 1477.8000 704.4000 1479.0000 705.6000 ;
	    RECT 1475.4000 695.4000 1476.6000 696.6000 ;
	    RECT 1480.3500 648.6000 1481.2500 707.4000 ;
	    RECT 1482.6000 705.4500 1483.8000 705.6000 ;
	    RECT 1482.6000 704.5500 1490.8500 705.4500 ;
	    RECT 1482.6000 704.4000 1483.8000 704.5500 ;
	    RECT 1489.9501 702.6000 1490.8500 704.5500 ;
	    RECT 1489.8000 701.4000 1491.0000 702.6000 ;
	    RECT 1485.0000 689.4000 1486.2001 690.6000 ;
	    RECT 1482.6000 683.4000 1483.8000 684.6000 ;
	    RECT 1482.7500 681.6000 1483.6500 683.4000 ;
	    RECT 1482.6000 680.4000 1483.8000 681.6000 ;
	    RECT 1482.7500 672.6000 1483.6500 680.4000 ;
	    RECT 1485.1500 678.6000 1486.0500 689.4000 ;
	    RECT 1489.8000 680.4000 1491.0000 681.6000 ;
	    RECT 1489.9501 678.6000 1490.8500 680.4000 ;
	    RECT 1485.0000 677.4000 1486.2001 678.6000 ;
	    RECT 1489.8000 677.4000 1491.0000 678.6000 ;
	    RECT 1497.1500 675.6000 1498.0500 923.4000 ;
	    RECT 1499.5500 768.6000 1500.4501 965.4000 ;
	    RECT 1501.9501 924.6000 1502.8500 1010.5500 ;
	    RECT 1501.8000 923.4000 1503.0000 924.6000 ;
	    RECT 1501.8000 917.4000 1503.0000 918.6000 ;
	    RECT 1501.9501 894.6000 1502.8500 917.4000 ;
	    RECT 1501.8000 893.4000 1503.0000 894.6000 ;
	    RECT 1504.3500 843.4500 1505.2500 1079.4000 ;
	    RECT 1506.6000 1049.4000 1507.8000 1050.6000 ;
	    RECT 1506.7500 915.4500 1507.6500 1049.4000 ;
	    RECT 1509.1500 1008.6000 1510.0500 1097.4000 ;
	    RECT 1511.4000 1085.4000 1512.6000 1086.6000 ;
	    RECT 1509.0000 1007.4000 1510.2001 1008.6000 ;
	    RECT 1511.5500 1002.6000 1512.4501 1085.4000 ;
	    RECT 1513.9501 1050.6000 1514.8500 1100.4000 ;
	    RECT 1521.0000 1091.4000 1522.2001 1092.6000 ;
	    RECT 1521.1500 1068.6000 1522.0500 1091.4000 ;
	    RECT 1516.2001 1067.4000 1517.4000 1068.6000 ;
	    RECT 1521.0000 1067.4000 1522.2001 1068.6000 ;
	    RECT 1516.3500 1062.6000 1517.2500 1067.4000 ;
	    RECT 1521.0000 1064.4000 1522.2001 1065.6000 ;
	    RECT 1516.2001 1061.4000 1517.4000 1062.6000 ;
	    RECT 1521.1500 1050.6000 1522.0500 1064.4000 ;
	    RECT 1513.8000 1049.4000 1515.0000 1050.6000 ;
	    RECT 1521.0000 1049.4000 1522.2001 1050.6000 ;
	    RECT 1513.8000 1026.3000 1515.0000 1046.7001 ;
	    RECT 1516.2001 1026.3000 1517.4000 1046.7001 ;
	    RECT 1518.6000 1026.3000 1519.8000 1046.7001 ;
	    RECT 1521.0000 1029.3000 1522.2001 1046.7001 ;
	    RECT 1523.5500 1044.6000 1524.4501 1115.5500 ;
	    RECT 1528.2001 1115.4000 1529.4000 1116.6000 ;
	    RECT 1525.8000 1097.4000 1527.0000 1098.6000 ;
	    RECT 1525.9501 1092.6000 1526.8500 1097.4000 ;
	    RECT 1528.3500 1095.6000 1529.2500 1115.4000 ;
	    RECT 1535.5500 1095.6000 1536.4501 1205.4000 ;
	    RECT 1528.2001 1094.4000 1529.4000 1095.6000 ;
	    RECT 1533.0000 1094.4000 1534.2001 1095.6000 ;
	    RECT 1535.4000 1094.4000 1536.6000 1095.6000 ;
	    RECT 1525.8000 1091.4000 1527.0000 1092.6000 ;
	    RECT 1533.1500 1080.6000 1534.0500 1094.4000 ;
	    RECT 1535.5500 1086.6000 1536.4501 1094.4000 ;
	    RECT 1535.4000 1085.4000 1536.6000 1086.6000 ;
	    RECT 1537.9501 1080.6000 1538.8500 1274.4000 ;
	    RECT 1540.2001 1199.4000 1541.4000 1200.6000 ;
	    RECT 1540.3500 1194.6000 1541.2500 1199.4000 ;
	    RECT 1540.2001 1193.4000 1541.4000 1194.6000 ;
	    RECT 1542.7500 1179.6000 1543.6500 1325.4000 ;
	    RECT 1545.1500 1230.6000 1546.0500 1367.4000 ;
	    RECT 1549.9501 1341.6000 1550.8500 1373.4000 ;
	    RECT 1554.6000 1364.4000 1555.8000 1365.6000 ;
	    RECT 1549.8000 1340.4000 1551.0000 1341.6000 ;
	    RECT 1547.4000 1337.4000 1548.6000 1338.6000 ;
	    RECT 1554.7500 1326.6000 1555.6500 1364.4000 ;
	    RECT 1554.6000 1325.4000 1555.8000 1326.6000 ;
	    RECT 1547.4000 1319.4000 1548.6000 1320.6000 ;
	    RECT 1547.5500 1281.6000 1548.4501 1319.4000 ;
	    RECT 1554.6000 1301.4000 1555.8000 1302.6000 ;
	    RECT 1552.2001 1298.4000 1553.4000 1299.6000 ;
	    RECT 1547.4000 1280.4000 1548.6000 1281.6000 ;
	    RECT 1547.4000 1238.4000 1548.6000 1239.6000 ;
	    RECT 1545.0000 1229.4000 1546.2001 1230.6000 ;
	    RECT 1545.0000 1209.3000 1546.2001 1226.7001 ;
	    RECT 1545.0000 1193.4000 1546.2001 1194.6000 ;
	    RECT 1542.6000 1178.4000 1543.8000 1179.6000 ;
	    RECT 1540.2001 1175.4000 1541.4000 1176.6000 ;
	    RECT 1533.0000 1079.4000 1534.2001 1080.6000 ;
	    RECT 1537.8000 1079.4000 1539.0000 1080.6000 ;
	    RECT 1540.3500 1071.4501 1541.2500 1175.4000 ;
	    RECT 1545.1500 1077.4501 1546.0500 1193.4000 ;
	    RECT 1547.5500 1182.6000 1548.4501 1238.4000 ;
	    RECT 1549.8000 1229.4000 1551.0000 1230.6000 ;
	    RECT 1547.4000 1181.4000 1548.6000 1182.6000 ;
	    RECT 1547.4000 1178.4000 1548.6000 1179.6000 ;
	    RECT 1537.9501 1070.5500 1541.2500 1071.4501 ;
	    RECT 1542.7500 1076.5500 1546.0500 1077.4501 ;
	    RECT 1528.2001 1061.4000 1529.4000 1062.6000 ;
	    RECT 1523.4000 1043.4000 1524.6000 1044.6000 ;
	    RECT 1521.0000 1025.4000 1522.2001 1026.6000 ;
	    RECT 1523.5500 1026.4501 1524.4501 1043.4000 ;
	    RECT 1525.8000 1029.3000 1527.0000 1046.7001 ;
	    RECT 1528.3500 1041.6000 1529.2500 1061.4000 ;
	    RECT 1528.2001 1040.4000 1529.4000 1041.6000 ;
	    RECT 1530.6000 1029.3000 1531.8000 1046.7001 ;
	    RECT 1523.5500 1025.5500 1526.8500 1026.4501 ;
	    RECT 1533.0000 1026.3000 1534.2001 1046.7001 ;
	    RECT 1535.4000 1026.3000 1536.6000 1046.7001 ;
	    RECT 1537.9501 1038.6000 1538.8500 1070.5500 ;
	    RECT 1540.2001 1067.4000 1541.4000 1068.6000 ;
	    RECT 1537.8000 1037.4000 1539.0000 1038.6000 ;
	    RECT 1516.2001 1022.4000 1517.4000 1023.6000 ;
	    RECT 1513.8000 1019.4000 1515.0000 1020.6000 ;
	    RECT 1511.4000 1001.4000 1512.6000 1002.6000 ;
	    RECT 1509.0000 971.4000 1510.2001 972.6000 ;
	    RECT 1509.1500 957.6000 1510.0500 971.4000 ;
	    RECT 1513.9501 960.6000 1514.8500 1019.4000 ;
	    RECT 1516.3500 1014.6000 1517.2500 1022.4000 ;
	    RECT 1516.2001 1013.4000 1517.4000 1014.6000 ;
	    RECT 1521.1500 1011.6000 1522.0500 1025.4000 ;
	    RECT 1521.0000 1011.4500 1522.2001 1011.6000 ;
	    RECT 1518.7500 1010.5500 1522.2001 1011.4500 ;
	    RECT 1516.2001 1001.4000 1517.4000 1002.6000 ;
	    RECT 1516.3500 990.6000 1517.2500 1001.4000 ;
	    RECT 1516.2001 989.4000 1517.4000 990.6000 ;
	    RECT 1516.3500 978.6000 1517.2500 989.4000 ;
	    RECT 1518.7500 981.6000 1519.6500 1010.5500 ;
	    RECT 1521.0000 1010.4000 1522.2001 1010.5500 ;
	    RECT 1521.0000 1007.4000 1522.2001 1008.6000 ;
	    RECT 1521.1500 990.6000 1522.0500 1007.4000 ;
	    RECT 1523.4000 1001.4000 1524.6000 1002.6000 ;
	    RECT 1521.0000 989.4000 1522.2001 990.6000 ;
	    RECT 1518.6000 980.4000 1519.8000 981.6000 ;
	    RECT 1516.2001 977.4000 1517.4000 978.6000 ;
	    RECT 1513.8000 959.4000 1515.0000 960.6000 ;
	    RECT 1518.6000 959.4000 1519.8000 960.6000 ;
	    RECT 1509.0000 956.4000 1510.2001 957.6000 ;
	    RECT 1518.7500 921.6000 1519.6500 959.4000 ;
	    RECT 1521.1500 948.6000 1522.0500 989.4000 ;
	    RECT 1523.5500 984.6000 1524.4501 1001.4000 ;
	    RECT 1525.9501 996.6000 1526.8500 1025.5500 ;
	    RECT 1535.4000 1013.4000 1536.6000 1014.6000 ;
	    RECT 1535.5500 1008.6000 1536.4501 1013.4000 ;
	    RECT 1533.0000 1007.4000 1534.2001 1008.6000 ;
	    RECT 1535.4000 1007.4000 1536.6000 1008.6000 ;
	    RECT 1533.1500 999.6000 1534.0500 1007.4000 ;
	    RECT 1533.0000 998.4000 1534.2001 999.6000 ;
	    RECT 1537.9501 999.4500 1538.8500 1037.4000 ;
	    RECT 1540.3500 1008.6000 1541.2500 1067.4000 ;
	    RECT 1542.7500 1062.6000 1543.6500 1076.5500 ;
	    RECT 1545.0000 1073.4000 1546.2001 1074.6000 ;
	    RECT 1542.6000 1061.4000 1543.8000 1062.6000 ;
	    RECT 1545.1500 1059.4501 1546.0500 1073.4000 ;
	    RECT 1542.7500 1058.5500 1546.0500 1059.4501 ;
	    RECT 1540.2001 1007.4000 1541.4000 1008.6000 ;
	    RECT 1540.2001 1004.4000 1541.4000 1005.6000 ;
	    RECT 1540.3500 1002.6000 1541.2500 1004.4000 ;
	    RECT 1540.2001 1001.4000 1541.4000 1002.6000 ;
	    RECT 1535.5500 998.5500 1538.8500 999.4500 ;
	    RECT 1525.8000 995.4000 1527.0000 996.6000 ;
	    RECT 1523.4000 983.4000 1524.6000 984.6000 ;
	    RECT 1523.4000 977.4000 1524.6000 978.6000 ;
	    RECT 1523.5500 966.6000 1524.4501 977.4000 ;
	    RECT 1535.5500 972.6000 1536.4501 998.5500 ;
	    RECT 1537.8000 995.4000 1539.0000 996.6000 ;
	    RECT 1535.4000 971.4000 1536.6000 972.6000 ;
	    RECT 1523.4000 965.4000 1524.6000 966.6000 ;
	    RECT 1525.8000 959.4000 1527.0000 960.6000 ;
	    RECT 1521.0000 947.4000 1522.2001 948.6000 ;
	    RECT 1521.0000 929.4000 1522.2001 930.6000 ;
	    RECT 1518.6000 920.4000 1519.8000 921.6000 ;
	    RECT 1521.1500 918.6000 1522.0500 929.4000 ;
	    RECT 1521.0000 917.4000 1522.2001 918.6000 ;
	    RECT 1506.7500 914.5500 1510.0500 915.4500 ;
	    RECT 1504.3500 842.5500 1507.6500 843.4500 ;
	    RECT 1501.8000 827.4000 1503.0000 828.6000 ;
	    RECT 1504.2001 827.4000 1505.4000 828.6000 ;
	    RECT 1501.9501 768.6000 1502.8500 827.4000 ;
	    RECT 1504.3500 801.6000 1505.2500 827.4000 ;
	    RECT 1504.2001 800.4000 1505.4000 801.6000 ;
	    RECT 1504.2001 785.4000 1505.4000 786.6000 ;
	    RECT 1499.4000 767.4000 1500.6000 768.6000 ;
	    RECT 1501.8000 767.4000 1503.0000 768.6000 ;
	    RECT 1504.3500 762.6000 1505.2500 785.4000 ;
	    RECT 1504.2001 761.4000 1505.4000 762.6000 ;
	    RECT 1506.7500 741.6000 1507.6500 842.5500 ;
	    RECT 1504.2001 740.4000 1505.4000 741.6000 ;
	    RECT 1506.6000 740.4000 1507.8000 741.6000 ;
	    RECT 1504.3500 738.6000 1505.2500 740.4000 ;
	    RECT 1509.1500 738.6000 1510.0500 914.5500 ;
	    RECT 1525.9501 906.6000 1526.8500 959.4000 ;
	    RECT 1528.2001 936.3000 1529.4000 956.7000 ;
	    RECT 1530.6000 936.3000 1531.8000 956.7000 ;
	    RECT 1533.0000 936.3000 1534.2001 956.7000 ;
	    RECT 1535.4000 936.3000 1536.6000 953.7000 ;
	    RECT 1537.9501 939.6000 1538.8500 995.4000 ;
	    RECT 1542.7500 981.6000 1543.6500 1058.5500 ;
	    RECT 1545.0000 1034.4000 1546.2001 1035.6000 ;
	    RECT 1547.5500 1008.6000 1548.4501 1178.4000 ;
	    RECT 1549.9501 1116.6000 1550.8500 1229.4000 ;
	    RECT 1552.3500 1218.6000 1553.2500 1298.4000 ;
	    RECT 1552.2001 1217.4000 1553.4000 1218.6000 ;
	    RECT 1552.3500 1206.6000 1553.2500 1217.4000 ;
	    RECT 1552.2001 1205.4000 1553.4000 1206.6000 ;
	    RECT 1554.7500 1194.6000 1555.6500 1301.4000 ;
	    RECT 1554.6000 1193.4000 1555.8000 1194.6000 ;
	    RECT 1557.1500 1188.4501 1558.0500 1454.4000 ;
	    RECT 1559.4000 1409.4000 1560.6000 1410.6000 ;
	    RECT 1559.5500 1392.6000 1560.4501 1409.4000 ;
	    RECT 1559.4000 1391.4000 1560.6000 1392.6000 ;
	    RECT 1559.4000 1370.4000 1560.6000 1371.6000 ;
	    RECT 1554.7500 1187.5500 1558.0500 1188.4501 ;
	    RECT 1549.8000 1115.4000 1551.0000 1116.6000 ;
	    RECT 1549.8000 1097.4000 1551.0000 1098.6000 ;
	    RECT 1552.2001 1097.4000 1553.4000 1098.6000 ;
	    RECT 1547.4000 1007.4000 1548.6000 1008.6000 ;
	    RECT 1547.4000 989.4000 1548.6000 990.6000 ;
	    RECT 1542.6000 981.4500 1543.8000 981.6000 ;
	    RECT 1540.3500 980.5500 1543.8000 981.4500 ;
	    RECT 1540.3500 972.6000 1541.2500 980.5500 ;
	    RECT 1542.6000 980.4000 1543.8000 980.5500 ;
	    RECT 1547.5500 975.6000 1548.4501 989.4000 ;
	    RECT 1547.4000 974.4000 1548.6000 975.6000 ;
	    RECT 1540.2001 971.4000 1541.4000 972.6000 ;
	    RECT 1542.6000 971.4000 1543.8000 972.6000 ;
	    RECT 1537.8000 938.4000 1539.0000 939.6000 ;
	    RECT 1537.9501 933.4500 1538.8500 938.4000 ;
	    RECT 1540.2001 936.3000 1541.4000 953.7000 ;
	    RECT 1542.7500 948.6000 1543.6500 971.4000 ;
	    RECT 1549.9501 960.6000 1550.8500 1097.4000 ;
	    RECT 1552.3500 1068.6000 1553.2500 1097.4000 ;
	    RECT 1552.2001 1067.4000 1553.4000 1068.6000 ;
	    RECT 1552.2001 1061.4000 1553.4000 1062.6000 ;
	    RECT 1549.8000 959.4000 1551.0000 960.6000 ;
	    RECT 1542.6000 947.4000 1543.8000 948.6000 ;
	    RECT 1542.6000 941.4000 1543.8000 942.6000 ;
	    RECT 1537.9501 932.5500 1541.2500 933.4500 ;
	    RECT 1530.6000 923.4000 1531.8000 924.6000 ;
	    RECT 1530.7500 918.6000 1531.6500 923.4000 ;
	    RECT 1530.6000 917.4000 1531.8000 918.6000 ;
	    RECT 1533.0000 917.4000 1534.2001 918.6000 ;
	    RECT 1535.4000 917.4000 1536.6000 918.6000 ;
	    RECT 1525.8000 905.4000 1527.0000 906.6000 ;
	    RECT 1513.8000 896.4000 1515.0000 897.6000 ;
	    RECT 1513.9501 888.6000 1514.8500 896.4000 ;
	    RECT 1513.8000 887.4000 1515.0000 888.6000 ;
	    RECT 1518.6000 884.4000 1519.8000 885.6000 ;
	    RECT 1518.7500 870.6000 1519.6500 884.4000 ;
	    RECT 1521.0000 876.3000 1522.2001 896.7000 ;
	    RECT 1523.4000 876.3000 1524.6000 896.7000 ;
	    RECT 1525.8000 876.3000 1527.0000 893.7000 ;
	    RECT 1528.2001 893.4000 1529.4000 894.6000 ;
	    RECT 1528.3500 882.6000 1529.2500 893.4000 ;
	    RECT 1528.2001 881.4000 1529.4000 882.6000 ;
	    RECT 1530.6000 876.3000 1531.8000 893.7000 ;
	    RECT 1533.1500 879.6000 1534.0500 917.4000 ;
	    RECT 1535.5500 912.6000 1536.4501 917.4000 ;
	    RECT 1540.3500 912.6000 1541.2500 932.5500 ;
	    RECT 1542.7500 921.6000 1543.6500 941.4000 ;
	    RECT 1545.0000 936.3000 1546.2001 953.7000 ;
	    RECT 1547.4000 936.3000 1548.6000 956.7000 ;
	    RECT 1549.8000 936.3000 1551.0000 956.7000 ;
	    RECT 1552.3500 954.6000 1553.2500 1061.4000 ;
	    RECT 1552.2001 953.4000 1553.4000 954.6000 ;
	    RECT 1552.2001 947.4000 1553.4000 948.6000 ;
	    RECT 1552.3500 945.6000 1553.2500 947.4000 ;
	    RECT 1552.2001 944.4000 1553.4000 945.6000 ;
	    RECT 1542.6000 920.4000 1543.8000 921.6000 ;
	    RECT 1535.4000 911.4000 1536.6000 912.6000 ;
	    RECT 1540.2001 911.4000 1541.4000 912.6000 ;
	    RECT 1545.0000 911.4000 1546.2001 912.6000 ;
	    RECT 1533.0000 878.4000 1534.2001 879.6000 ;
	    RECT 1535.4000 876.3000 1536.6000 893.7000 ;
	    RECT 1537.8000 876.3000 1539.0000 896.7000 ;
	    RECT 1540.2001 876.3000 1541.4000 896.7000 ;
	    RECT 1542.6000 876.3000 1543.8000 896.7000 ;
	    RECT 1545.1500 870.6000 1546.0500 911.4000 ;
	    RECT 1547.4000 905.4000 1548.6000 906.6000 ;
	    RECT 1518.6000 869.4000 1519.8000 870.6000 ;
	    RECT 1530.6000 869.4000 1531.8000 870.6000 ;
	    RECT 1545.0000 869.4000 1546.2001 870.6000 ;
	    RECT 1521.0000 846.3000 1522.2001 866.7000 ;
	    RECT 1523.4000 846.3000 1524.6000 866.7000 ;
	    RECT 1525.8000 846.3000 1527.0000 866.7000 ;
	    RECT 1528.2001 849.3000 1529.4000 866.7000 ;
	    RECT 1530.7500 864.6000 1531.6500 869.4000 ;
	    RECT 1530.6000 863.4000 1531.8000 864.6000 ;
	    RECT 1518.6000 839.4000 1519.8000 840.6000 ;
	    RECT 1518.7500 765.6000 1519.6500 839.4000 ;
	    RECT 1530.7500 834.6000 1531.6500 863.4000 ;
	    RECT 1533.0000 849.3000 1534.2001 866.7000 ;
	    RECT 1535.4000 860.4000 1536.6000 861.6000 ;
	    RECT 1530.6000 833.4000 1531.8000 834.6000 ;
	    RECT 1533.0000 827.4000 1534.2001 828.6000 ;
	    RECT 1533.1500 825.6000 1534.0500 827.4000 ;
	    RECT 1533.0000 824.4000 1534.2001 825.6000 ;
	    RECT 1535.5500 822.6000 1536.4501 860.4000 ;
	    RECT 1537.8000 849.3000 1539.0000 866.7000 ;
	    RECT 1540.2001 846.3000 1541.4000 866.7000 ;
	    RECT 1542.6000 846.3000 1543.8000 866.7000 ;
	    RECT 1545.0000 857.4000 1546.2001 858.6000 ;
	    RECT 1535.4000 821.4000 1536.6000 822.6000 ;
	    RECT 1537.8000 819.3000 1539.0000 827.7000 ;
	    RECT 1540.2001 821.4000 1541.4000 822.6000 ;
	    RECT 1528.2001 809.4000 1529.4000 810.6000 ;
	    RECT 1528.3500 801.6000 1529.2500 809.4000 ;
	    RECT 1523.4000 800.4000 1524.6000 801.6000 ;
	    RECT 1528.2001 800.4000 1529.4000 801.6000 ;
	    RECT 1533.0000 800.4000 1534.2001 801.6000 ;
	    RECT 1523.5500 798.6000 1524.4501 800.4000 ;
	    RECT 1523.4000 797.4000 1524.6000 798.6000 ;
	    RECT 1525.8000 797.4000 1527.0000 798.6000 ;
	    RECT 1530.6000 797.4000 1531.8000 798.6000 ;
	    RECT 1523.5500 768.6000 1524.4501 797.4000 ;
	    RECT 1523.4000 767.4000 1524.6000 768.6000 ;
	    RECT 1511.4000 764.4000 1512.6000 765.6000 ;
	    RECT 1518.6000 764.4000 1519.8000 765.6000 ;
	    RECT 1511.5500 762.6000 1512.4501 764.4000 ;
	    RECT 1511.4000 761.4000 1512.6000 762.6000 ;
	    RECT 1516.2001 761.4000 1517.4000 762.6000 ;
	    RECT 1516.3500 744.6000 1517.2500 761.4000 ;
	    RECT 1518.7500 750.6000 1519.6500 764.4000 ;
	    RECT 1518.6000 749.4000 1519.8000 750.6000 ;
	    RECT 1516.2001 743.4000 1517.4000 744.6000 ;
	    RECT 1523.4000 743.4000 1524.6000 744.6000 ;
	    RECT 1518.6000 740.4000 1519.8000 741.6000 ;
	    RECT 1504.2001 737.4000 1505.4000 738.6000 ;
	    RECT 1506.6000 737.4000 1507.8000 738.6000 ;
	    RECT 1509.0000 737.4000 1510.2001 738.6000 ;
	    RECT 1497.0000 674.4000 1498.2001 675.6000 ;
	    RECT 1482.6000 671.4000 1483.8000 672.6000 ;
	    RECT 1504.3500 648.6000 1505.2500 737.4000 ;
	    RECT 1506.7500 720.6000 1507.6500 737.4000 ;
	    RECT 1506.6000 719.4000 1507.8000 720.6000 ;
	    RECT 1506.7500 708.6000 1507.6500 719.4000 ;
	    RECT 1506.6000 707.4000 1507.8000 708.6000 ;
	    RECT 1511.4000 707.4000 1512.6000 708.6000 ;
	    RECT 1506.6000 701.4000 1507.8000 702.6000 ;
	    RECT 1506.7500 678.6000 1507.6500 701.4000 ;
	    RECT 1511.5500 681.6000 1512.4501 707.4000 ;
	    RECT 1511.4000 680.4000 1512.6000 681.6000 ;
	    RECT 1506.6000 677.4000 1507.8000 678.6000 ;
	    RECT 1513.8000 677.4000 1515.0000 678.6000 ;
	    RECT 1480.2001 647.4000 1481.4000 648.6000 ;
	    RECT 1485.0000 647.4000 1486.2001 648.6000 ;
	    RECT 1492.2001 647.4000 1493.4000 648.6000 ;
	    RECT 1504.2001 647.4000 1505.4000 648.6000 ;
	    RECT 1482.6000 641.4000 1483.8000 642.6000 ;
	    RECT 1477.8000 635.4000 1479.0000 636.6000 ;
	    RECT 1477.9501 621.6000 1478.8500 635.4000 ;
	    RECT 1480.2001 623.4000 1481.4000 624.6000 ;
	    RECT 1477.8000 620.4000 1479.0000 621.6000 ;
	    RECT 1482.7500 618.6000 1483.6500 641.4000 ;
	    RECT 1475.4000 617.4000 1476.6000 618.6000 ;
	    RECT 1482.6000 617.4000 1483.8000 618.6000 ;
	    RECT 1485.1500 612.6000 1486.0500 647.4000 ;
	    RECT 1492.3500 645.6000 1493.2500 647.4000 ;
	    RECT 1492.2001 644.4000 1493.4000 645.6000 ;
	    RECT 1501.8000 644.4000 1503.0000 645.6000 ;
	    RECT 1504.2001 644.4000 1505.4000 645.6000 ;
	    RECT 1494.6000 641.4000 1495.8000 642.6000 ;
	    RECT 1494.7500 636.6000 1495.6500 641.4000 ;
	    RECT 1494.6000 635.4000 1495.8000 636.6000 ;
	    RECT 1487.4000 629.4000 1488.6000 630.6000 ;
	    RECT 1485.0000 611.4000 1486.2001 612.6000 ;
	    RECT 1487.5500 588.6000 1488.4501 629.4000 ;
	    RECT 1497.0000 614.4000 1498.2001 615.6000 ;
	    RECT 1492.2001 590.4000 1493.4000 591.6000 ;
	    RECT 1492.3500 588.6000 1493.2500 590.4000 ;
	    RECT 1497.1500 588.6000 1498.0500 614.4000 ;
	    RECT 1487.4000 587.4000 1488.6000 588.6000 ;
	    RECT 1489.8000 587.4000 1491.0000 588.6000 ;
	    RECT 1492.2001 587.4000 1493.4000 588.6000 ;
	    RECT 1497.0000 587.4000 1498.2001 588.6000 ;
	    RECT 1489.9501 570.6000 1490.8500 587.4000 ;
	    RECT 1494.6000 584.4000 1495.8000 585.6000 ;
	    RECT 1494.7500 582.6000 1495.6500 584.4000 ;
	    RECT 1494.6000 581.4000 1495.8000 582.6000 ;
	    RECT 1489.8000 569.4000 1491.0000 570.6000 ;
	    RECT 1482.6000 563.4000 1483.8000 564.6000 ;
	    RECT 1485.0000 563.4000 1486.2001 564.6000 ;
	    RECT 1482.7500 558.6000 1483.6500 563.4000 ;
	    RECT 1485.1500 558.6000 1486.0500 563.4000 ;
	    RECT 1494.7500 561.6000 1495.6500 581.4000 ;
	    RECT 1497.1500 564.6000 1498.0500 587.4000 ;
	    RECT 1501.9501 585.6000 1502.8500 644.4000 ;
	    RECT 1504.3500 639.6000 1505.2500 644.4000 ;
	    RECT 1504.2001 638.4000 1505.4000 639.6000 ;
	    RECT 1509.0000 617.4000 1510.2001 618.6000 ;
	    RECT 1501.8000 584.4000 1503.0000 585.6000 ;
	    RECT 1497.0000 563.4000 1498.2001 564.6000 ;
	    RECT 1489.8000 560.4000 1491.0000 561.6000 ;
	    RECT 1494.6000 560.4000 1495.8000 561.6000 ;
	    RECT 1506.6000 560.4000 1507.8000 561.6000 ;
	    RECT 1482.6000 557.4000 1483.8000 558.6000 ;
	    RECT 1485.0000 557.4000 1486.2001 558.6000 ;
	    RECT 1475.4000 554.4000 1476.6000 555.6000 ;
	    RECT 1473.0000 545.4000 1474.2001 546.6000 ;
	    RECT 1473.1500 528.6000 1474.0500 545.4000 ;
	    RECT 1473.0000 527.4000 1474.2001 528.6000 ;
	    RECT 1470.6000 437.4000 1471.8000 438.6000 ;
	    RECT 1475.5500 435.4500 1476.4501 554.4000 ;
	    RECT 1477.8000 551.4000 1479.0000 552.6000 ;
	    RECT 1477.9501 468.6000 1478.8500 551.4000 ;
	    RECT 1489.9501 546.6000 1490.8500 560.4000 ;
	    RECT 1492.2001 557.4000 1493.4000 558.6000 ;
	    RECT 1489.8000 545.4000 1491.0000 546.6000 ;
	    RECT 1492.3500 540.6000 1493.2500 557.4000 ;
	    RECT 1492.2001 539.4000 1493.4000 540.6000 ;
	    RECT 1497.0000 533.4000 1498.2001 534.6000 ;
	    RECT 1497.1500 531.6000 1498.0500 533.4000 ;
	    RECT 1497.0000 530.4000 1498.2001 531.6000 ;
	    RECT 1492.2001 527.4000 1493.4000 528.6000 ;
	    RECT 1494.6000 527.4000 1495.8000 528.6000 ;
	    RECT 1501.8000 527.4000 1503.0000 528.6000 ;
	    RECT 1482.6000 497.4000 1483.8000 498.6000 ;
	    RECT 1487.4000 497.4000 1488.6000 498.6000 ;
	    RECT 1480.2001 473.4000 1481.4000 474.6000 ;
	    RECT 1480.3500 468.6000 1481.2500 473.4000 ;
	    RECT 1477.8000 467.4000 1479.0000 468.6000 ;
	    RECT 1480.2001 467.4000 1481.4000 468.6000 ;
	    RECT 1482.7500 465.6000 1483.6500 497.4000 ;
	    RECT 1492.3500 495.6000 1493.2500 527.4000 ;
	    RECT 1494.7500 495.6000 1495.6500 527.4000 ;
	    RECT 1499.4000 524.4000 1500.6000 525.6000 ;
	    RECT 1499.5500 522.6000 1500.4501 524.4000 ;
	    RECT 1499.4000 521.4000 1500.6000 522.6000 ;
	    RECT 1492.2001 494.4000 1493.4000 495.6000 ;
	    RECT 1494.6000 494.4000 1495.8000 495.6000 ;
	    RECT 1489.8000 491.4000 1491.0000 492.6000 ;
	    RECT 1485.0000 470.4000 1486.2001 471.6000 ;
	    RECT 1485.1500 468.6000 1486.0500 470.4000 ;
	    RECT 1489.9501 468.6000 1490.8500 491.4000 ;
	    RECT 1485.0000 467.4000 1486.2001 468.6000 ;
	    RECT 1489.8000 467.4000 1491.0000 468.6000 ;
	    RECT 1482.6000 464.4000 1483.8000 465.6000 ;
	    RECT 1482.7500 447.6000 1483.6500 464.4000 ;
	    RECT 1482.6000 446.4000 1483.8000 447.6000 ;
	    RECT 1475.5500 434.5500 1478.8500 435.4500 ;
	    RECT 1470.6000 401.4000 1471.8000 402.6000 ;
	    RECT 1475.4000 401.4000 1476.6000 402.6000 ;
	    RECT 1470.7500 381.6000 1471.6500 401.4000 ;
	    RECT 1470.6000 380.4000 1471.8000 381.6000 ;
	    RECT 1473.0000 365.4000 1474.2001 366.6000 ;
	    RECT 1470.6000 350.4000 1471.8000 351.6000 ;
	    RECT 1470.7500 348.6000 1471.6500 350.4000 ;
	    RECT 1468.2001 347.4000 1469.4000 348.6000 ;
	    RECT 1470.6000 347.4000 1471.8000 348.6000 ;
	    RECT 1473.1500 345.6000 1474.0500 365.4000 ;
	    RECT 1473.0000 344.4000 1474.2001 345.6000 ;
	    RECT 1465.8000 290.4000 1467.0000 291.6000 ;
	    RECT 1470.6000 269.4000 1471.8000 270.6000 ;
	    RECT 1470.7500 255.6000 1471.6500 269.4000 ;
	    RECT 1473.1500 267.6000 1474.0500 344.4000 ;
	    RECT 1475.5500 300.6000 1476.4501 401.4000 ;
	    RECT 1477.9501 315.6000 1478.8500 434.5500 ;
	    RECT 1487.4000 413.4000 1488.6000 414.6000 ;
	    RECT 1487.5500 399.6000 1488.4501 413.4000 ;
	    RECT 1487.4000 398.4000 1488.6000 399.6000 ;
	    RECT 1482.6000 395.4000 1483.8000 396.6000 ;
	    RECT 1482.7500 384.6000 1483.6500 395.4000 ;
	    RECT 1489.9501 384.6000 1490.8500 467.4000 ;
	    RECT 1501.9501 465.6000 1502.8500 527.4000 ;
	    RECT 1504.2001 524.4000 1505.4000 525.6000 ;
	    RECT 1504.3500 522.6000 1505.2500 524.4000 ;
	    RECT 1504.2001 521.4000 1505.4000 522.6000 ;
	    RECT 1506.7500 468.6000 1507.6500 560.4000 ;
	    RECT 1509.1500 528.6000 1510.0500 617.4000 ;
	    RECT 1511.4000 611.4000 1512.6000 612.6000 ;
	    RECT 1511.5500 552.6000 1512.4501 611.4000 ;
	    RECT 1513.9501 570.4500 1514.8500 677.4000 ;
	    RECT 1518.7500 636.4500 1519.6500 740.4000 ;
	    RECT 1523.5500 738.6000 1524.4501 743.4000 ;
	    RECT 1523.4000 737.4000 1524.6000 738.6000 ;
	    RECT 1525.9501 705.6000 1526.8500 797.4000 ;
	    RECT 1528.2001 779.4000 1529.4000 780.6000 ;
	    RECT 1528.3500 738.6000 1529.2500 779.4000 ;
	    RECT 1530.7500 762.6000 1531.6500 797.4000 ;
	    RECT 1533.1500 780.6000 1534.0500 800.4000 ;
	    RECT 1535.4000 794.4000 1536.6000 795.6000 ;
	    RECT 1535.5500 792.6000 1536.4501 794.4000 ;
	    RECT 1535.4000 791.4000 1536.6000 792.6000 ;
	    RECT 1533.0000 779.4000 1534.2001 780.6000 ;
	    RECT 1533.0000 767.4000 1534.2001 768.6000 ;
	    RECT 1530.6000 761.4000 1531.8000 762.6000 ;
	    RECT 1528.2001 737.4000 1529.4000 738.6000 ;
	    RECT 1525.8000 704.4000 1527.0000 705.6000 ;
	    RECT 1523.4000 701.4000 1524.6000 702.6000 ;
	    RECT 1521.0000 695.4000 1522.2001 696.6000 ;
	    RECT 1521.1500 684.6000 1522.0500 695.4000 ;
	    RECT 1521.0000 683.4000 1522.2001 684.6000 ;
	    RECT 1523.5500 678.6000 1524.4501 701.4000 ;
	    RECT 1525.8000 683.4000 1527.0000 684.6000 ;
	    RECT 1523.4000 677.4000 1524.6000 678.6000 ;
	    RECT 1525.8000 677.4000 1527.0000 678.6000 ;
	    RECT 1523.4000 638.4000 1524.6000 639.6000 ;
	    RECT 1521.0000 636.4500 1522.2001 636.6000 ;
	    RECT 1518.7500 635.5500 1522.2001 636.4500 ;
	    RECT 1521.0000 635.4000 1522.2001 635.5500 ;
	    RECT 1521.1500 615.6000 1522.0500 635.4000 ;
	    RECT 1523.5500 624.6000 1524.4501 638.4000 ;
	    RECT 1523.4000 623.4000 1524.6000 624.6000 ;
	    RECT 1518.6000 614.4000 1519.8000 615.6000 ;
	    RECT 1521.0000 614.4000 1522.2001 615.6000 ;
	    RECT 1518.7500 612.6000 1519.6500 614.4000 ;
	    RECT 1518.6000 611.4000 1519.8000 612.6000 ;
	    RECT 1523.4000 584.4000 1524.6000 585.6000 ;
	    RECT 1521.0000 581.4000 1522.2001 582.6000 ;
	    RECT 1521.1500 576.6000 1522.0500 581.4000 ;
	    RECT 1521.0000 575.4000 1522.2001 576.6000 ;
	    RECT 1516.2001 570.4500 1517.4000 570.6000 ;
	    RECT 1513.9501 569.5500 1517.4000 570.4500 ;
	    RECT 1516.2001 569.4000 1517.4000 569.5500 ;
	    RECT 1516.3500 555.6000 1517.2500 569.4000 ;
	    RECT 1523.5500 561.6000 1524.4501 584.4000 ;
	    RECT 1523.4000 561.4500 1524.6000 561.6000 ;
	    RECT 1521.1500 560.5500 1524.6000 561.4500 ;
	    RECT 1516.2001 554.4000 1517.4000 555.6000 ;
	    RECT 1511.4000 551.4000 1512.6000 552.6000 ;
	    RECT 1521.1500 528.6000 1522.0500 560.5500 ;
	    RECT 1523.4000 560.4000 1524.6000 560.5500 ;
	    RECT 1525.9501 534.6000 1526.8500 677.4000 ;
	    RECT 1530.6000 644.4000 1531.8000 645.6000 ;
	    RECT 1528.2001 641.4000 1529.4000 642.6000 ;
	    RECT 1528.3500 612.6000 1529.2500 641.4000 ;
	    RECT 1530.7500 630.6000 1531.6500 644.4000 ;
	    RECT 1530.6000 629.4000 1531.8000 630.6000 ;
	    RECT 1530.7500 618.6000 1531.6500 629.4000 ;
	    RECT 1530.6000 617.4000 1531.8000 618.6000 ;
	    RECT 1528.2001 611.4000 1529.4000 612.6000 ;
	    RECT 1533.1500 588.6000 1534.0500 767.4000 ;
	    RECT 1537.8000 761.4000 1539.0000 762.6000 ;
	    RECT 1537.9501 705.6000 1538.8500 761.4000 ;
	    RECT 1537.8000 704.4000 1539.0000 705.6000 ;
	    RECT 1535.4000 695.4000 1536.6000 696.6000 ;
	    RECT 1535.5500 639.6000 1536.4501 695.4000 ;
	    RECT 1535.4000 638.4000 1536.6000 639.6000 ;
	    RECT 1533.0000 587.4000 1534.2001 588.6000 ;
	    RECT 1537.8000 581.4000 1539.0000 582.6000 ;
	    RECT 1535.4000 557.4000 1536.6000 558.6000 ;
	    RECT 1525.8000 533.4000 1527.0000 534.6000 ;
	    RECT 1509.0000 527.4000 1510.2001 528.6000 ;
	    RECT 1521.0000 527.4000 1522.2001 528.6000 ;
	    RECT 1516.2001 509.4000 1517.4000 510.6000 ;
	    RECT 1516.3500 501.6000 1517.2500 509.4000 ;
	    RECT 1535.5500 504.6000 1536.4501 557.4000 ;
	    RECT 1537.9501 525.6000 1538.8500 581.4000 ;
	    RECT 1537.8000 524.4000 1539.0000 525.6000 ;
	    RECT 1518.6000 503.4000 1519.8000 504.6000 ;
	    RECT 1535.4000 503.4000 1536.6000 504.6000 ;
	    RECT 1516.2001 500.4000 1517.4000 501.6000 ;
	    RECT 1506.6000 467.4000 1507.8000 468.6000 ;
	    RECT 1501.8000 464.4000 1503.0000 465.6000 ;
	    RECT 1506.6000 461.4000 1507.8000 462.6000 ;
	    RECT 1504.2001 425.4000 1505.4000 426.6000 ;
	    RECT 1504.3500 402.6000 1505.2500 425.4000 ;
	    RECT 1506.7500 408.6000 1507.6500 461.4000 ;
	    RECT 1509.0000 419.4000 1510.2001 420.6000 ;
	    RECT 1506.6000 407.4000 1507.8000 408.6000 ;
	    RECT 1504.2001 401.4000 1505.4000 402.6000 ;
	    RECT 1482.6000 383.4000 1483.8000 384.6000 ;
	    RECT 1489.8000 383.4000 1491.0000 384.6000 ;
	    RECT 1501.8000 383.4000 1503.0000 384.6000 ;
	    RECT 1487.4000 377.4000 1488.6000 378.6000 ;
	    RECT 1497.0000 377.4000 1498.2001 378.6000 ;
	    RECT 1497.1500 366.6000 1498.0500 377.4000 ;
	    RECT 1497.0000 365.4000 1498.2001 366.6000 ;
	    RECT 1492.2001 359.4000 1493.4000 360.6000 ;
	    RECT 1485.0000 347.4000 1486.2001 348.6000 ;
	    RECT 1477.8000 314.4000 1479.0000 315.6000 ;
	    RECT 1482.6000 314.4000 1483.8000 315.6000 ;
	    RECT 1477.8000 305.4000 1479.0000 306.6000 ;
	    RECT 1475.4000 299.4000 1476.6000 300.6000 ;
	    RECT 1477.9501 282.6000 1478.8500 305.4000 ;
	    RECT 1480.2001 293.4000 1481.4000 294.6000 ;
	    RECT 1480.3500 285.6000 1481.2500 293.4000 ;
	    RECT 1480.2001 284.4000 1481.4000 285.6000 ;
	    RECT 1477.8000 281.4000 1479.0000 282.6000 ;
	    RECT 1473.0000 266.4000 1474.2001 267.6000 ;
	    RECT 1480.2001 266.4000 1481.4000 267.6000 ;
	    RECT 1461.0000 254.4000 1462.2001 255.6000 ;
	    RECT 1470.6000 254.4000 1471.8000 255.6000 ;
	    RECT 1461.1500 234.6000 1462.0500 254.4000 ;
	    RECT 1470.7500 240.6000 1471.6500 254.4000 ;
	    RECT 1470.6000 239.4000 1471.8000 240.6000 ;
	    RECT 1461.0000 233.4000 1462.2001 234.6000 ;
	    RECT 1470.6000 230.4000 1471.8000 231.6000 ;
	    RECT 1463.4000 221.4000 1464.6000 222.6000 ;
	    RECT 1456.2001 167.4000 1457.4000 168.6000 ;
	    RECT 1461.0000 164.4000 1462.2001 165.6000 ;
	    RECT 1441.8000 161.4000 1443.0000 162.6000 ;
	    RECT 1444.2001 161.4000 1445.4000 162.6000 ;
	    RECT 1449.0000 161.4000 1450.2001 162.6000 ;
	    RECT 1453.8000 161.4000 1455.0000 162.6000 ;
	    RECT 1441.9501 141.6000 1442.8500 161.4000 ;
	    RECT 1444.3500 144.6000 1445.2500 161.4000 ;
	    RECT 1446.6000 149.4000 1447.8000 150.6000 ;
	    RECT 1444.2001 143.4000 1445.4000 144.6000 ;
	    RECT 1446.7500 141.6000 1447.6500 149.4000 ;
	    RECT 1441.8000 140.4000 1443.0000 141.6000 ;
	    RECT 1446.6000 140.4000 1447.8000 141.6000 ;
	    RECT 1461.1500 132.6000 1462.0500 164.4000 ;
	    RECT 1461.0000 131.4000 1462.2001 132.6000 ;
	    RECT 1444.2001 119.4000 1445.4000 120.6000 ;
	    RECT 1398.6000 83.4000 1399.8000 84.6000 ;
	    RECT 1401.0000 83.4000 1402.2001 84.6000 ;
	    RECT 1427.4000 83.4000 1428.6000 84.6000 ;
	    RECT 1434.6000 83.4000 1435.8000 84.6000 ;
	    RECT 1398.7500 66.6000 1399.6500 83.4000 ;
	    RECT 1427.4000 80.4000 1428.6000 81.6000 ;
	    RECT 1427.5500 78.6000 1428.4501 80.4000 ;
	    RECT 1427.4000 77.4000 1428.6000 78.6000 ;
	    RECT 1434.7500 75.6000 1435.6500 83.4000 ;
	    RECT 1444.3500 78.6000 1445.2500 119.4000 ;
	    RECT 1463.5500 114.6000 1464.4501 221.4000 ;
	    RECT 1468.2001 197.4000 1469.4000 198.6000 ;
	    RECT 1468.3500 195.6000 1469.2500 197.4000 ;
	    RECT 1468.2001 194.4000 1469.4000 195.6000 ;
	    RECT 1470.7500 174.6000 1471.6500 230.4000 ;
	    RECT 1480.3500 228.6000 1481.2500 266.4000 ;
	    RECT 1482.7500 246.6000 1483.6500 314.4000 ;
	    RECT 1482.6000 245.4000 1483.8000 246.6000 ;
	    RECT 1473.0000 227.4000 1474.2001 228.6000 ;
	    RECT 1480.2001 227.4000 1481.4000 228.6000 ;
	    RECT 1473.1500 180.6000 1474.0500 227.4000 ;
	    RECT 1475.4000 224.4000 1476.6000 225.6000 ;
	    RECT 1475.5500 204.6000 1476.4501 224.4000 ;
	    RECT 1475.4000 203.4000 1476.6000 204.6000 ;
	    RECT 1480.2001 197.4000 1481.4000 198.6000 ;
	    RECT 1480.3500 192.6000 1481.2500 197.4000 ;
	    RECT 1485.1500 195.6000 1486.0500 347.4000 ;
	    RECT 1492.3500 336.6000 1493.2500 359.4000 ;
	    RECT 1501.9501 342.6000 1502.8500 383.4000 ;
	    RECT 1509.1500 375.6000 1510.0500 419.4000 ;
	    RECT 1518.7500 414.6000 1519.6500 503.4000 ;
	    RECT 1530.6000 497.4000 1531.8000 498.6000 ;
	    RECT 1523.4000 461.4000 1524.6000 462.6000 ;
	    RECT 1523.5500 426.6000 1524.4501 461.4000 ;
	    RECT 1523.4000 425.4000 1524.6000 426.6000 ;
	    RECT 1518.6000 413.4000 1519.8000 414.6000 ;
	    RECT 1518.7500 408.6000 1519.6500 413.4000 ;
	    RECT 1521.0000 410.4000 1522.2001 411.6000 ;
	    RECT 1521.1500 408.6000 1522.0500 410.4000 ;
	    RECT 1518.6000 407.4000 1519.8000 408.6000 ;
	    RECT 1521.0000 407.4000 1522.2001 408.6000 ;
	    RECT 1516.2001 404.4000 1517.4000 405.6000 ;
	    RECT 1516.3500 396.6000 1517.2500 404.4000 ;
	    RECT 1523.5500 399.6000 1524.4501 425.4000 ;
	    RECT 1530.7500 420.6000 1531.6500 497.4000 ;
	    RECT 1540.3500 471.4500 1541.2500 821.4000 ;
	    RECT 1542.6000 816.3000 1543.8000 833.7000 ;
	    RECT 1547.5500 828.4500 1548.4501 905.4000 ;
	    RECT 1552.3500 858.6000 1553.2500 944.4000 ;
	    RECT 1552.2001 857.4000 1553.4000 858.6000 ;
	    RECT 1552.2001 854.4000 1553.4000 855.6000 ;
	    RECT 1552.3500 846.6000 1553.2500 854.4000 ;
	    RECT 1552.2001 845.4000 1553.4000 846.6000 ;
	    RECT 1547.5500 827.5500 1550.8500 828.4500 ;
	    RECT 1547.4000 824.4000 1548.6000 825.6000 ;
	    RECT 1547.5500 810.6000 1548.4501 824.4000 ;
	    RECT 1547.4000 809.4000 1548.6000 810.6000 ;
	    RECT 1547.4000 791.4000 1548.6000 792.6000 ;
	    RECT 1545.0000 767.4000 1546.2001 768.6000 ;
	    RECT 1542.6000 719.4000 1543.8000 720.6000 ;
	    RECT 1542.7500 708.6000 1543.6500 719.4000 ;
	    RECT 1542.6000 707.4000 1543.8000 708.6000 ;
	    RECT 1545.1500 705.6000 1546.0500 767.4000 ;
	    RECT 1547.5500 735.6000 1548.4501 791.4000 ;
	    RECT 1549.9501 765.6000 1550.8500 827.5500 ;
	    RECT 1549.8000 764.4000 1551.0000 765.6000 ;
	    RECT 1552.2001 761.4000 1553.4000 762.6000 ;
	    RECT 1549.8000 749.4000 1551.0000 750.6000 ;
	    RECT 1547.4000 734.4000 1548.6000 735.6000 ;
	    RECT 1549.9501 732.6000 1550.8500 749.4000 ;
	    RECT 1552.2001 743.4000 1553.4000 744.6000 ;
	    RECT 1552.3500 738.6000 1553.2500 743.4000 ;
	    RECT 1552.2001 737.4000 1553.4000 738.6000 ;
	    RECT 1554.7500 738.4500 1555.6500 1187.5500 ;
	    RECT 1557.0000 1184.4000 1558.2001 1185.6000 ;
	    RECT 1557.1500 1182.6000 1558.0500 1184.4000 ;
	    RECT 1557.0000 1181.4000 1558.2001 1182.6000 ;
	    RECT 1557.1500 1152.6000 1558.0500 1181.4000 ;
	    RECT 1557.0000 1151.4000 1558.2001 1152.6000 ;
	    RECT 1559.5500 1110.6000 1560.4501 1370.4000 ;
	    RECT 1561.8000 1367.4000 1563.0000 1368.6000 ;
	    RECT 1561.9501 1278.6000 1562.8500 1367.4000 ;
	    RECT 1561.8000 1277.4000 1563.0000 1278.6000 ;
	    RECT 1564.3500 1248.6000 1565.2500 1457.4000 ;
	    RECT 1566.7500 1332.6000 1567.6500 1460.4000 ;
	    RECT 1566.6000 1331.4000 1567.8000 1332.6000 ;
	    RECT 1564.2001 1247.4000 1565.4000 1248.6000 ;
	    RECT 1559.4000 1109.4000 1560.6000 1110.6000 ;
	    RECT 1561.8000 1097.4000 1563.0000 1098.6000 ;
	    RECT 1566.6000 1097.4000 1567.8000 1098.6000 ;
	    RECT 1561.9501 1074.6000 1562.8500 1097.4000 ;
	    RECT 1566.7500 1095.6000 1567.6500 1097.4000 ;
	    RECT 1566.6000 1094.4000 1567.8000 1095.6000 ;
	    RECT 1564.2001 1091.4000 1565.4000 1092.6000 ;
	    RECT 1564.2001 1079.4000 1565.4000 1080.6000 ;
	    RECT 1561.8000 1073.4000 1563.0000 1074.6000 ;
	    RECT 1561.8000 1067.4000 1563.0000 1068.6000 ;
	    RECT 1557.0000 1064.4000 1558.2001 1065.6000 ;
	    RECT 1557.1500 1014.6000 1558.0500 1064.4000 ;
	    RECT 1559.4000 1061.4000 1560.6000 1062.6000 ;
	    RECT 1557.0000 1013.4000 1558.2001 1014.6000 ;
	    RECT 1559.5500 1008.6000 1560.4501 1061.4000 ;
	    RECT 1559.4000 1007.4000 1560.6000 1008.6000 ;
	    RECT 1561.9501 978.6000 1562.8500 1067.4000 ;
	    RECT 1561.8000 977.4000 1563.0000 978.6000 ;
	    RECT 1557.0000 957.4500 1558.2001 957.6000 ;
	    RECT 1557.0000 956.5500 1560.4501 957.4500 ;
	    RECT 1557.0000 956.4000 1558.2001 956.5500 ;
	    RECT 1557.0000 953.4000 1558.2001 954.6000 ;
	    RECT 1557.1500 840.6000 1558.0500 953.4000 ;
	    RECT 1559.5500 948.6000 1560.4501 956.5500 ;
	    RECT 1559.4000 947.4000 1560.6000 948.6000 ;
	    RECT 1559.5500 921.6000 1560.4501 947.4000 ;
	    RECT 1559.4000 920.4000 1560.6000 921.6000 ;
	    RECT 1564.3500 918.6000 1565.2500 1079.4000 ;
	    RECT 1566.6000 1025.4000 1567.8000 1026.6000 ;
	    RECT 1559.4000 917.4000 1560.6000 918.6000 ;
	    RECT 1564.2001 917.4000 1565.4000 918.6000 ;
	    RECT 1559.5500 891.6000 1560.4501 917.4000 ;
	    RECT 1559.4000 890.4000 1560.6000 891.6000 ;
	    RECT 1566.6000 845.4000 1567.8000 846.6000 ;
	    RECT 1566.7500 843.6000 1567.6500 845.4000 ;
	    RECT 1566.6000 842.4000 1567.8000 843.6000 ;
	    RECT 1557.0000 839.4000 1558.2001 840.6000 ;
	    RECT 1557.0000 816.3000 1558.2001 833.7000 ;
	    RECT 1564.2001 827.4000 1565.4000 828.6000 ;
	    RECT 1564.3500 825.6000 1565.2500 827.4000 ;
	    RECT 1564.2001 824.4000 1565.4000 825.6000 ;
	    RECT 1561.8000 797.4000 1563.0000 798.6000 ;
	    RECT 1564.2001 797.4000 1565.4000 798.6000 ;
	    RECT 1561.9501 792.6000 1562.8500 797.4000 ;
	    RECT 1564.3500 795.6000 1565.2500 797.4000 ;
	    RECT 1564.2001 794.4000 1565.4000 795.6000 ;
	    RECT 1559.4000 791.4000 1560.6000 792.6000 ;
	    RECT 1561.8000 791.4000 1563.0000 792.6000 ;
	    RECT 1559.5500 786.6000 1560.4501 791.4000 ;
	    RECT 1559.4000 785.4000 1560.6000 786.6000 ;
	    RECT 1554.7500 737.5500 1558.0500 738.4500 ;
	    RECT 1554.6000 734.4000 1555.8000 735.6000 ;
	    RECT 1554.7500 732.6000 1555.6500 734.4000 ;
	    RECT 1549.8000 731.4000 1551.0000 732.6000 ;
	    RECT 1554.6000 731.4000 1555.8000 732.6000 ;
	    RECT 1545.0000 704.4000 1546.2001 705.6000 ;
	    RECT 1554.6000 701.4000 1555.8000 702.6000 ;
	    RECT 1554.7500 678.6000 1555.6500 701.4000 ;
	    RECT 1557.1500 681.6000 1558.0500 737.5500 ;
	    RECT 1566.6000 722.4000 1567.8000 723.6000 ;
	    RECT 1566.7500 720.6000 1567.6500 722.4000 ;
	    RECT 1561.8000 719.4000 1563.0000 720.6000 ;
	    RECT 1566.6000 719.4000 1567.8000 720.6000 ;
	    RECT 1561.9501 702.6000 1562.8500 719.4000 ;
	    RECT 1561.8000 701.4000 1563.0000 702.6000 ;
	    RECT 1557.0000 680.4000 1558.2001 681.6000 ;
	    RECT 1554.6000 677.4000 1555.8000 678.6000 ;
	    RECT 1547.4000 641.4000 1548.6000 642.6000 ;
	    RECT 1547.5500 624.6000 1548.4501 641.4000 ;
	    RECT 1547.4000 623.4000 1548.6000 624.6000 ;
	    RECT 1545.0000 617.4000 1546.2001 618.6000 ;
	    RECT 1547.5500 615.6000 1548.4501 623.4000 ;
	    RECT 1547.4000 614.4000 1548.6000 615.6000 ;
	    RECT 1542.6000 611.4000 1543.8000 612.6000 ;
	    RECT 1557.1500 582.6000 1558.0500 680.4000 ;
	    RECT 1542.6000 581.4000 1543.8000 582.6000 ;
	    RECT 1545.0000 581.4000 1546.2001 582.6000 ;
	    RECT 1557.0000 581.4000 1558.2001 582.6000 ;
	    RECT 1542.7500 579.6000 1543.6500 581.4000 ;
	    RECT 1542.6000 578.4000 1543.8000 579.6000 ;
	    RECT 1545.1500 576.6000 1546.0500 581.4000 ;
	    RECT 1545.0000 575.4000 1546.2001 576.6000 ;
	    RECT 1542.6000 558.4500 1543.8000 558.6000 ;
	    RECT 1545.1500 558.4500 1546.0500 575.4000 ;
	    RECT 1542.6000 557.5500 1546.0500 558.4500 ;
	    RECT 1542.6000 557.4000 1543.8000 557.5500 ;
	    RECT 1545.1500 522.6000 1546.0500 557.5500 ;
	    RECT 1542.6000 521.4000 1543.8000 522.6000 ;
	    RECT 1545.0000 521.4000 1546.2001 522.6000 ;
	    RECT 1542.7500 498.6000 1543.6500 521.4000 ;
	    RECT 1547.4000 500.4000 1548.6000 501.6000 ;
	    RECT 1542.6000 497.4000 1543.8000 498.6000 ;
	    RECT 1537.9501 470.5500 1541.2500 471.4500 ;
	    RECT 1533.0000 455.4000 1534.2001 456.6000 ;
	    RECT 1530.6000 419.4000 1531.8000 420.6000 ;
	    RECT 1523.4000 398.4000 1524.6000 399.6000 ;
	    RECT 1516.2001 395.4000 1517.4000 396.6000 ;
	    RECT 1533.1500 390.6000 1534.0500 455.4000 ;
	    RECT 1535.4000 435.3000 1536.6000 443.7000 ;
	    RECT 1537.9501 441.6000 1538.8500 470.5500 ;
	    RECT 1545.0000 470.4000 1546.2001 471.6000 ;
	    RECT 1540.2001 467.4000 1541.4000 468.6000 ;
	    RECT 1542.6000 467.4000 1543.8000 468.6000 ;
	    RECT 1540.3500 465.6000 1541.2500 467.4000 ;
	    RECT 1540.2001 464.4000 1541.4000 465.6000 ;
	    RECT 1542.7500 462.6000 1543.6500 467.4000 ;
	    RECT 1542.6000 461.4000 1543.8000 462.6000 ;
	    RECT 1545.1500 459.4500 1546.0500 470.4000 ;
	    RECT 1547.5500 468.6000 1548.4501 500.4000 ;
	    RECT 1549.8000 497.4000 1551.0000 498.6000 ;
	    RECT 1549.9501 471.6000 1550.8500 497.4000 ;
	    RECT 1549.8000 470.4000 1551.0000 471.6000 ;
	    RECT 1557.1500 468.6000 1558.0500 581.4000 ;
	    RECT 1559.4000 557.4000 1560.6000 558.6000 ;
	    RECT 1559.5500 525.6000 1560.4501 557.4000 ;
	    RECT 1559.4000 524.4000 1560.6000 525.6000 ;
	    RECT 1564.2001 524.4000 1565.4000 525.6000 ;
	    RECT 1564.3500 522.6000 1565.2500 524.4000 ;
	    RECT 1561.8000 521.4000 1563.0000 522.6000 ;
	    RECT 1564.2001 521.4000 1565.4000 522.6000 ;
	    RECT 1566.6000 521.4000 1567.8000 522.6000 ;
	    RECT 1561.9501 510.6000 1562.8500 521.4000 ;
	    RECT 1561.8000 509.4000 1563.0000 510.6000 ;
	    RECT 1547.4000 467.4000 1548.6000 468.6000 ;
	    RECT 1557.0000 467.4000 1558.2001 468.6000 ;
	    RECT 1561.8000 467.4000 1563.0000 468.6000 ;
	    RECT 1542.7500 458.5500 1546.0500 459.4500 ;
	    RECT 1537.8000 440.4000 1539.0000 441.6000 ;
	    RECT 1537.9501 438.6000 1538.8500 440.4000 ;
	    RECT 1537.8000 437.4000 1539.0000 438.6000 ;
	    RECT 1540.2001 429.3000 1541.4000 446.7000 ;
	    RECT 1540.2001 413.4000 1541.4000 414.6000 ;
	    RECT 1540.3500 405.6000 1541.2500 413.4000 ;
	    RECT 1540.2001 404.4000 1541.4000 405.6000 ;
	    RECT 1516.2001 389.4000 1517.4000 390.6000 ;
	    RECT 1533.0000 389.4000 1534.2001 390.6000 ;
	    RECT 1509.0000 374.4000 1510.2001 375.6000 ;
	    RECT 1513.8000 371.4000 1515.0000 372.6000 ;
	    RECT 1513.9501 348.6000 1514.8500 371.4000 ;
	    RECT 1513.8000 347.4000 1515.0000 348.6000 ;
	    RECT 1501.8000 341.4000 1503.0000 342.6000 ;
	    RECT 1509.0000 341.4000 1510.2001 342.6000 ;
	    RECT 1492.2001 335.4000 1493.4000 336.6000 ;
	    RECT 1489.8000 317.4000 1491.0000 318.6000 ;
	    RECT 1489.9501 300.6000 1490.8500 317.4000 ;
	    RECT 1492.3500 312.6000 1493.2500 335.4000 ;
	    RECT 1509.1500 315.6000 1510.0500 341.4000 ;
	    RECT 1509.0000 314.4000 1510.2001 315.6000 ;
	    RECT 1511.4000 314.4000 1512.6000 315.6000 ;
	    RECT 1492.2001 311.4000 1493.4000 312.6000 ;
	    RECT 1489.8000 299.4000 1491.0000 300.6000 ;
	    RECT 1506.6000 287.4000 1507.8000 288.6000 ;
	    RECT 1487.4000 281.4000 1488.6000 282.6000 ;
	    RECT 1487.5500 258.6000 1488.4501 281.4000 ;
	    RECT 1506.7500 270.6000 1507.6500 287.4000 ;
	    RECT 1506.6000 269.4000 1507.8000 270.6000 ;
	    RECT 1509.1500 258.6000 1510.0500 314.4000 ;
	    RECT 1511.5500 294.6000 1512.4501 314.4000 ;
	    RECT 1511.4000 293.4000 1512.6000 294.6000 ;
	    RECT 1511.5500 285.6000 1512.4501 293.4000 ;
	    RECT 1511.4000 284.4000 1512.6000 285.6000 ;
	    RECT 1513.8000 281.4000 1515.0000 282.6000 ;
	    RECT 1487.4000 257.4000 1488.6000 258.6000 ;
	    RECT 1509.0000 257.4000 1510.2001 258.6000 ;
	    RECT 1487.5500 234.6000 1488.4501 257.4000 ;
	    RECT 1492.2001 254.4000 1493.4000 255.6000 ;
	    RECT 1497.0000 254.4000 1498.2001 255.6000 ;
	    RECT 1489.8000 251.4000 1491.0000 252.6000 ;
	    RECT 1487.4000 233.4000 1488.6000 234.6000 ;
	    RECT 1492.3500 204.6000 1493.2500 254.4000 ;
	    RECT 1494.6000 227.4000 1495.8000 228.6000 ;
	    RECT 1492.2001 203.4000 1493.4000 204.6000 ;
	    RECT 1485.0000 194.4000 1486.2001 195.6000 ;
	    RECT 1480.2001 191.4000 1481.4000 192.6000 ;
	    RECT 1473.0000 179.4000 1474.2001 180.6000 ;
	    RECT 1470.6000 173.4000 1471.8000 174.6000 ;
	    RECT 1492.2001 173.4000 1493.4000 174.6000 ;
	    RECT 1477.8000 170.4000 1479.0000 171.6000 ;
	    RECT 1473.0000 167.4000 1474.2001 168.6000 ;
	    RECT 1465.8000 161.4000 1467.0000 162.6000 ;
	    RECT 1465.9501 138.6000 1466.8500 161.4000 ;
	    RECT 1468.2001 158.4000 1469.4000 159.6000 ;
	    RECT 1465.8000 137.4000 1467.0000 138.6000 ;
	    RECT 1463.4000 113.4000 1464.6000 114.6000 ;
	    RECT 1453.8000 110.4000 1455.0000 111.6000 ;
	    RECT 1453.9501 90.6000 1454.8500 110.4000 ;
	    RECT 1463.4000 107.4000 1464.6000 108.6000 ;
	    RECT 1453.8000 89.4000 1455.0000 90.6000 ;
	    RECT 1458.6000 89.4000 1459.8000 90.6000 ;
	    RECT 1444.2001 77.4000 1445.4000 78.6000 ;
	    RECT 1434.6000 74.4000 1435.8000 75.6000 ;
	    RECT 1398.6000 65.4000 1399.8000 66.6000 ;
	    RECT 1434.6000 65.4000 1435.8000 66.6000 ;
	    RECT 1396.2001 59.4000 1397.4000 60.6000 ;
	    RECT 1391.4000 56.4000 1392.6000 57.6000 ;
	    RECT 1391.5500 48.6000 1392.4501 56.4000 ;
	    RECT 1391.4000 47.4000 1392.6000 48.6000 ;
	    RECT 1396.3500 45.6000 1397.2500 59.4000 ;
	    RECT 1396.2001 44.4000 1397.4000 45.6000 ;
	    RECT 1374.6000 35.4000 1375.8000 36.6000 ;
	    RECT 1398.6000 36.3000 1399.8000 56.7000 ;
	    RECT 1401.0000 36.3000 1402.2001 56.7000 ;
	    RECT 1403.4000 36.3000 1404.6000 53.7000 ;
	    RECT 1405.8000 41.4000 1407.0000 42.6000 ;
	    RECT 1408.2001 36.3000 1409.4000 53.7000 ;
	    RECT 1410.6000 38.4000 1411.8000 39.6000 ;
	    RECT 1410.7500 36.6000 1411.6500 38.4000 ;
	    RECT 1410.6000 35.4000 1411.8000 36.6000 ;
	    RECT 1413.0000 36.3000 1414.2001 53.7000 ;
	    RECT 1415.4000 36.3000 1416.6000 56.7000 ;
	    RECT 1417.8000 36.3000 1419.0000 56.7000 ;
	    RECT 1420.2001 36.3000 1421.4000 56.7000 ;
	    RECT 1434.7500 51.6000 1435.6500 65.4000 ;
	    RECT 1434.6000 50.4000 1435.8000 51.6000 ;
	    RECT 1453.9501 45.6000 1454.8500 89.4000 ;
	    RECT 1456.2001 83.4000 1457.4000 84.6000 ;
	    RECT 1456.3500 72.6000 1457.2500 83.4000 ;
	    RECT 1458.7500 81.6000 1459.6500 89.4000 ;
	    RECT 1463.5500 81.6000 1464.4501 107.4000 ;
	    RECT 1465.9501 84.6000 1466.8500 137.4000 ;
	    RECT 1465.8000 83.4000 1467.0000 84.6000 ;
	    RECT 1458.6000 80.4000 1459.8000 81.6000 ;
	    RECT 1463.4000 80.4000 1464.6000 81.6000 ;
	    RECT 1458.6000 77.4000 1459.8000 78.6000 ;
	    RECT 1465.8000 77.4000 1467.0000 78.6000 ;
	    RECT 1456.2001 71.4000 1457.4000 72.6000 ;
	    RECT 1458.7500 60.6000 1459.6500 77.4000 ;
	    RECT 1458.6000 59.4000 1459.8000 60.6000 ;
	    RECT 1465.9501 51.6000 1466.8500 77.4000 ;
	    RECT 1468.3500 72.6000 1469.2500 158.4000 ;
	    RECT 1473.1500 144.6000 1474.0500 167.4000 ;
	    RECT 1473.0000 143.4000 1474.2001 144.6000 ;
	    RECT 1477.9501 138.6000 1478.8500 170.4000 ;
	    RECT 1492.3500 168.6000 1493.2500 173.4000 ;
	    RECT 1492.2001 167.4000 1493.4000 168.6000 ;
	    RECT 1494.7500 165.6000 1495.6500 227.4000 ;
	    RECT 1497.1500 171.6000 1498.0500 254.4000 ;
	    RECT 1511.4000 239.4000 1512.6000 240.6000 ;
	    RECT 1509.0000 233.4000 1510.2001 234.6000 ;
	    RECT 1509.1500 231.6000 1510.0500 233.4000 ;
	    RECT 1509.0000 230.4000 1510.2001 231.6000 ;
	    RECT 1511.5500 225.6000 1512.4501 239.4000 ;
	    RECT 1513.8000 234.4500 1515.0000 234.6000 ;
	    RECT 1516.3500 234.4500 1517.2500 389.4000 ;
	    RECT 1518.6000 380.4000 1519.8000 381.6000 ;
	    RECT 1518.7500 315.6000 1519.6500 380.4000 ;
	    RECT 1535.4000 377.4000 1536.6000 378.6000 ;
	    RECT 1537.8000 374.4000 1539.0000 375.6000 ;
	    RECT 1537.9501 372.6000 1538.8500 374.4000 ;
	    RECT 1533.0000 371.4000 1534.2001 372.6000 ;
	    RECT 1535.4000 371.4000 1536.6000 372.6000 ;
	    RECT 1537.8000 371.4000 1539.0000 372.6000 ;
	    RECT 1533.1500 360.6000 1534.0500 371.4000 ;
	    RECT 1533.0000 359.4000 1534.2001 360.6000 ;
	    RECT 1521.3000 347.7000 1522.5000 348.9000 ;
	    RECT 1530.6000 347.7000 1531.8000 348.9000 ;
	    RECT 1521.3000 340.5000 1522.2001 347.7000 ;
	    RECT 1523.1000 344.7000 1524.3000 345.9000 ;
	    RECT 1523.4000 342.6000 1524.3000 344.7000 ;
	    RECT 1530.9000 342.6000 1531.8000 347.7000 ;
	    RECT 1523.4000 341.7000 1531.8000 342.6000 ;
	    RECT 1523.4000 340.5000 1524.6000 340.8000 ;
	    RECT 1528.5000 340.5000 1529.7001 340.8000 ;
	    RECT 1530.9000 340.5000 1531.8000 341.7000 ;
	    RECT 1521.3000 339.6000 1529.7001 340.5000 ;
	    RECT 1521.3000 339.3000 1522.5000 339.6000 ;
	    RECT 1530.6000 339.3000 1531.8000 340.5000 ;
	    RECT 1521.0000 320.4000 1522.2001 321.6000 ;
	    RECT 1518.6000 314.4000 1519.8000 315.6000 ;
	    RECT 1518.6000 282.4500 1519.8000 282.6000 ;
	    RECT 1521.1500 282.4500 1522.0500 320.4000 ;
	    RECT 1535.5500 318.6000 1536.4501 371.4000 ;
	    RECT 1537.8000 353.4000 1539.0000 354.6000 ;
	    RECT 1537.9501 345.6000 1538.8500 353.4000 ;
	    RECT 1540.2001 347.4000 1541.4000 348.6000 ;
	    RECT 1537.8000 344.4000 1539.0000 345.6000 ;
	    RECT 1535.4000 317.4000 1536.6000 318.6000 ;
	    RECT 1537.9501 282.6000 1538.8500 344.4000 ;
	    RECT 1540.3500 342.6000 1541.2500 347.4000 ;
	    RECT 1540.2001 341.4000 1541.4000 342.6000 ;
	    RECT 1540.2001 329.4000 1541.4000 330.6000 ;
	    RECT 1540.3500 321.6000 1541.2500 329.4000 ;
	    RECT 1542.7500 321.6000 1543.6500 458.5500 ;
	    RECT 1545.0000 437.4000 1546.2001 438.6000 ;
	    RECT 1545.1500 420.6000 1546.0500 437.4000 ;
	    RECT 1545.0000 419.4000 1546.2001 420.6000 ;
	    RECT 1540.2001 320.4000 1541.4000 321.6000 ;
	    RECT 1542.6000 320.4000 1543.8000 321.6000 ;
	    RECT 1542.6000 317.4000 1543.8000 318.6000 ;
	    RECT 1540.2001 287.4000 1541.4000 288.6000 ;
	    RECT 1540.3500 285.6000 1541.2500 287.4000 ;
	    RECT 1540.2001 284.4000 1541.4000 285.6000 ;
	    RECT 1518.6000 281.5500 1522.0500 282.4500 ;
	    RECT 1518.6000 281.4000 1519.8000 281.5500 ;
	    RECT 1537.8000 281.4000 1539.0000 282.6000 ;
	    RECT 1540.2001 281.4000 1541.4000 282.6000 ;
	    RECT 1513.8000 233.5500 1517.2500 234.4500 ;
	    RECT 1513.8000 233.4000 1515.0000 233.5500 ;
	    RECT 1513.9501 228.6000 1514.8500 233.4000 ;
	    RECT 1513.8000 227.4000 1515.0000 228.6000 ;
	    RECT 1511.4000 224.4000 1512.6000 225.6000 ;
	    RECT 1513.9501 222.6000 1514.8500 227.4000 ;
	    RECT 1513.8000 221.4000 1515.0000 222.6000 ;
	    RECT 1518.7500 216.6000 1519.6500 281.4000 ;
	    RECT 1540.3500 279.6000 1541.2500 281.4000 ;
	    RECT 1542.7500 279.6000 1543.6500 317.4000 ;
	    RECT 1540.2001 278.4000 1541.4000 279.6000 ;
	    RECT 1542.6000 278.4000 1543.8000 279.6000 ;
	    RECT 1523.4000 275.4000 1524.6000 276.6000 ;
	    RECT 1521.0000 263.4000 1522.2001 264.6000 ;
	    RECT 1521.1500 252.6000 1522.0500 263.4000 ;
	    RECT 1523.5500 258.6000 1524.4501 275.4000 ;
	    RECT 1525.8000 269.4000 1527.0000 270.6000 ;
	    RECT 1540.2001 269.4000 1541.4000 270.6000 ;
	    RECT 1523.4000 257.4000 1524.6000 258.6000 ;
	    RECT 1521.0000 251.4000 1522.2001 252.6000 ;
	    RECT 1523.5500 240.6000 1524.4501 257.4000 ;
	    RECT 1525.9501 255.6000 1526.8500 269.4000 ;
	    RECT 1525.8000 254.4000 1527.0000 255.6000 ;
	    RECT 1523.4000 239.4000 1524.6000 240.6000 ;
	    RECT 1530.6000 227.4000 1531.8000 228.6000 ;
	    RECT 1509.0000 215.4000 1510.2001 216.6000 ;
	    RECT 1518.6000 215.4000 1519.8000 216.6000 ;
	    RECT 1506.6000 194.4000 1507.8000 195.6000 ;
	    RECT 1497.0000 170.4000 1498.2001 171.6000 ;
	    RECT 1499.4000 167.4000 1500.6000 168.6000 ;
	    RECT 1494.6000 164.4000 1495.8000 165.6000 ;
	    RECT 1480.2001 155.4000 1481.4000 156.6000 ;
	    RECT 1473.0000 137.4000 1474.2001 138.6000 ;
	    RECT 1477.8000 137.4000 1479.0000 138.6000 ;
	    RECT 1473.1500 132.6000 1474.0500 137.4000 ;
	    RECT 1477.8000 134.4000 1479.0000 135.6000 ;
	    RECT 1473.0000 131.4000 1474.2001 132.6000 ;
	    RECT 1477.9501 129.4500 1478.8500 134.4000 ;
	    RECT 1480.3500 132.6000 1481.2500 155.4000 ;
	    RECT 1494.7500 144.6000 1495.6500 164.4000 ;
	    RECT 1482.6000 143.4000 1483.8000 144.6000 ;
	    RECT 1494.6000 143.4000 1495.8000 144.6000 ;
	    RECT 1480.2001 131.4000 1481.4000 132.6000 ;
	    RECT 1482.7500 129.4500 1483.6500 143.4000 ;
	    RECT 1485.0000 134.4000 1486.2001 135.6000 ;
	    RECT 1494.6000 134.4000 1495.8000 135.6000 ;
	    RECT 1477.9501 128.5500 1483.6500 129.4500 ;
	    RECT 1485.1500 120.6000 1486.0500 134.4000 ;
	    RECT 1494.7500 132.6000 1495.6500 134.4000 ;
	    RECT 1494.6000 131.4000 1495.8000 132.6000 ;
	    RECT 1480.2001 119.4000 1481.4000 120.6000 ;
	    RECT 1485.0000 119.4000 1486.2001 120.6000 ;
	    RECT 1480.3500 72.6000 1481.2500 119.4000 ;
	    RECT 1482.6000 95.4000 1483.8000 96.6000 ;
	    RECT 1485.0000 96.3000 1486.2001 116.7000 ;
	    RECT 1487.4000 96.3000 1488.6000 116.7000 ;
	    RECT 1489.8000 96.3000 1491.0000 116.7000 ;
	    RECT 1492.2001 96.3000 1493.4000 113.7000 ;
	    RECT 1494.7500 102.6000 1495.6500 131.4000 ;
	    RECT 1494.6000 101.4000 1495.8000 102.6000 ;
	    RECT 1494.6000 98.4000 1495.8000 99.6000 ;
	    RECT 1494.7500 96.6000 1495.6500 98.4000 ;
	    RECT 1494.6000 95.4000 1495.8000 96.6000 ;
	    RECT 1497.0000 96.3000 1498.2001 113.7000 ;
	    RECT 1499.5500 108.6000 1500.4501 167.4000 ;
	    RECT 1506.7500 120.6000 1507.6500 194.4000 ;
	    RECT 1509.1500 141.6000 1510.0500 215.4000 ;
	    RECT 1511.4000 203.4000 1512.6000 204.6000 ;
	    RECT 1511.5500 192.6000 1512.4501 203.4000 ;
	    RECT 1530.7500 198.6000 1531.6500 227.4000 ;
	    RECT 1540.3500 198.6000 1541.2500 269.4000 ;
	    RECT 1545.0000 254.4000 1546.2001 255.6000 ;
	    RECT 1542.6000 239.4000 1543.8000 240.6000 ;
	    RECT 1542.7500 231.6000 1543.6500 239.4000 ;
	    RECT 1542.6000 230.4000 1543.8000 231.6000 ;
	    RECT 1545.1500 225.6000 1546.0500 254.4000 ;
	    RECT 1547.5500 252.4500 1548.4501 467.4000 ;
	    RECT 1557.0000 461.4000 1558.2001 462.6000 ;
	    RECT 1554.6000 458.4000 1555.8000 459.6000 ;
	    RECT 1554.7500 456.6000 1555.6500 458.4000 ;
	    RECT 1554.6000 455.4000 1555.8000 456.6000 ;
	    RECT 1554.6000 429.3000 1555.8000 446.7000 ;
	    RECT 1549.8000 407.4000 1551.0000 408.6000 ;
	    RECT 1549.9501 405.6000 1550.8500 407.4000 ;
	    RECT 1549.8000 404.4000 1551.0000 405.6000 ;
	    RECT 1549.9501 285.6000 1550.8500 404.4000 ;
	    RECT 1552.2001 401.4000 1553.4000 402.6000 ;
	    RECT 1552.3500 396.6000 1553.2500 401.4000 ;
	    RECT 1552.2001 395.4000 1553.4000 396.6000 ;
	    RECT 1552.3500 378.6000 1553.2500 395.4000 ;
	    RECT 1552.2001 377.4000 1553.4000 378.6000 ;
	    RECT 1554.6000 320.4000 1555.8000 321.6000 ;
	    RECT 1552.2001 317.4000 1553.4000 318.6000 ;
	    RECT 1552.3500 288.6000 1553.2500 317.4000 ;
	    RECT 1552.2001 287.4000 1553.4000 288.6000 ;
	    RECT 1549.8000 284.4000 1551.0000 285.6000 ;
	    RECT 1554.7500 270.6000 1555.6500 320.4000 ;
	    RECT 1554.6000 269.4000 1555.8000 270.6000 ;
	    RECT 1557.1500 264.6000 1558.0500 461.4000 ;
	    RECT 1561.9501 438.6000 1562.8500 467.4000 ;
	    RECT 1561.8000 437.4000 1563.0000 438.6000 ;
	    RECT 1566.7500 414.6000 1567.6500 521.4000 ;
	    RECT 1566.6000 413.4000 1567.8000 414.6000 ;
	    RECT 1561.8000 380.4000 1563.0000 381.6000 ;
	    RECT 1561.9501 354.6000 1562.8500 380.4000 ;
	    RECT 1561.8000 353.4000 1563.0000 354.6000 ;
	    RECT 1564.2001 350.4000 1565.4000 351.6000 ;
	    RECT 1559.4000 347.4000 1560.6000 348.6000 ;
	    RECT 1559.5500 282.6000 1560.4501 347.4000 ;
	    RECT 1561.8000 344.4000 1563.0000 345.6000 ;
	    RECT 1561.9501 330.6000 1562.8500 344.4000 ;
	    RECT 1561.8000 329.4000 1563.0000 330.6000 ;
	    RECT 1564.3500 294.6000 1565.2500 350.4000 ;
	    RECT 1566.6000 347.4000 1567.8000 348.6000 ;
	    RECT 1564.2001 293.4000 1565.4000 294.6000 ;
	    RECT 1559.4000 281.4000 1560.6000 282.6000 ;
	    RECT 1557.0000 263.4000 1558.2001 264.6000 ;
	    RECT 1549.8000 257.4000 1551.0000 258.6000 ;
	    RECT 1552.2001 257.4000 1553.4000 258.6000 ;
	    RECT 1554.6000 257.4000 1555.8000 258.6000 ;
	    RECT 1549.9501 255.6000 1550.8500 257.4000 ;
	    RECT 1549.8000 254.4000 1551.0000 255.6000 ;
	    RECT 1549.8000 252.4500 1551.0000 252.6000 ;
	    RECT 1547.5500 251.5500 1551.0000 252.4500 ;
	    RECT 1549.8000 251.4000 1551.0000 251.5500 ;
	    RECT 1547.4000 233.4000 1548.6000 234.6000 ;
	    RECT 1547.5500 228.6000 1548.4501 233.4000 ;
	    RECT 1547.4000 227.4000 1548.6000 228.6000 ;
	    RECT 1545.0000 224.4000 1546.2001 225.6000 ;
	    RECT 1542.6000 215.4000 1543.8000 216.6000 ;
	    RECT 1542.7500 204.6000 1543.6500 215.4000 ;
	    RECT 1552.3500 210.6000 1553.2500 257.4000 ;
	    RECT 1554.7500 252.6000 1555.6500 257.4000 ;
	    RECT 1557.0000 254.4000 1558.2001 255.6000 ;
	    RECT 1557.1500 252.6000 1558.0500 254.4000 ;
	    RECT 1554.6000 251.4000 1555.8000 252.6000 ;
	    RECT 1557.0000 251.4000 1558.2001 252.6000 ;
	    RECT 1559.5500 222.6000 1560.4501 281.4000 ;
	    RECT 1559.4000 221.4000 1560.6000 222.6000 ;
	    RECT 1561.8000 218.4000 1563.0000 219.6000 ;
	    RECT 1561.9501 216.6000 1562.8500 218.4000 ;
	    RECT 1561.8000 215.4000 1563.0000 216.6000 ;
	    RECT 1552.2001 209.4000 1553.4000 210.6000 ;
	    RECT 1561.8000 209.4000 1563.0000 210.6000 ;
	    RECT 1542.6000 203.4000 1543.8000 204.6000 ;
	    RECT 1513.8000 197.4000 1515.0000 198.6000 ;
	    RECT 1530.6000 197.4000 1531.8000 198.6000 ;
	    RECT 1540.2001 197.4000 1541.4000 198.6000 ;
	    RECT 1516.2001 194.4000 1517.4000 195.6000 ;
	    RECT 1511.4000 191.4000 1512.6000 192.6000 ;
	    RECT 1516.3500 174.6000 1517.2500 194.4000 ;
	    RECT 1528.2001 191.4000 1529.4000 192.6000 ;
	    RECT 1516.2001 173.4000 1517.4000 174.6000 ;
	    RECT 1525.8000 171.4500 1527.0000 171.6000 ;
	    RECT 1523.5500 170.5500 1527.0000 171.4500 ;
	    RECT 1518.6000 167.4000 1519.8000 168.6000 ;
	    RECT 1509.0000 140.4000 1510.2001 141.6000 ;
	    RECT 1516.2001 137.4000 1517.4000 138.6000 ;
	    RECT 1506.6000 119.4000 1507.8000 120.6000 ;
	    RECT 1511.4000 119.4000 1512.6000 120.6000 ;
	    RECT 1499.4000 107.4000 1500.6000 108.6000 ;
	    RECT 1499.4000 101.4000 1500.6000 102.6000 ;
	    RECT 1468.2001 71.4000 1469.4000 72.6000 ;
	    RECT 1480.2001 71.4000 1481.4000 72.6000 ;
	    RECT 1465.8000 50.4000 1467.0000 51.6000 ;
	    RECT 1453.8000 44.4000 1455.0000 45.6000 ;
	    RECT 1470.6000 35.4000 1471.8000 36.6000 ;
	    RECT 1470.7500 24.6000 1471.6500 35.4000 ;
	    RECT 1482.7500 30.4500 1483.6500 95.4000 ;
	    RECT 1499.5500 90.6000 1500.4501 101.4000 ;
	    RECT 1501.8000 96.3000 1503.0000 113.7000 ;
	    RECT 1504.2001 96.3000 1505.4000 116.7000 ;
	    RECT 1506.6000 96.3000 1507.8000 116.7000 ;
	    RECT 1509.0000 104.4000 1510.2001 105.6000 ;
	    RECT 1499.4000 89.4000 1500.6000 90.6000 ;
	    RECT 1489.8000 83.4000 1491.0000 84.6000 ;
	    RECT 1494.6000 83.4000 1495.8000 84.6000 ;
	    RECT 1485.0000 80.4000 1486.2001 81.6000 ;
	    RECT 1485.1500 48.6000 1486.0500 80.4000 ;
	    RECT 1489.9501 75.6000 1490.8500 83.4000 ;
	    RECT 1492.2001 77.4000 1493.4000 78.6000 ;
	    RECT 1489.8000 74.4000 1491.0000 75.6000 ;
	    RECT 1494.7500 72.6000 1495.6500 83.4000 ;
	    RECT 1487.4000 71.4000 1488.6000 72.6000 ;
	    RECT 1494.6000 71.4000 1495.8000 72.6000 ;
	    RECT 1497.0000 71.4000 1498.2001 72.6000 ;
	    RECT 1487.5500 48.6000 1488.4501 71.4000 ;
	    RECT 1497.1500 54.6000 1498.0500 71.4000 ;
	    RECT 1492.2001 53.4000 1493.4000 54.6000 ;
	    RECT 1497.0000 53.4000 1498.2001 54.6000 ;
	    RECT 1492.3500 51.6000 1493.2500 53.4000 ;
	    RECT 1492.2001 50.4000 1493.4000 51.6000 ;
	    RECT 1485.0000 47.4000 1486.2001 48.6000 ;
	    RECT 1487.4000 47.4000 1488.6000 48.6000 ;
	    RECT 1489.8000 47.4000 1491.0000 48.6000 ;
	    RECT 1489.9501 45.6000 1490.8500 47.4000 ;
	    RECT 1489.8000 44.4000 1491.0000 45.6000 ;
	    RECT 1509.1500 36.6000 1510.0500 104.4000 ;
	    RECT 1511.5500 78.6000 1512.4501 119.4000 ;
	    RECT 1513.8000 116.4000 1515.0000 117.6000 ;
	    RECT 1513.9501 108.6000 1514.8500 116.4000 ;
	    RECT 1513.8000 107.4000 1515.0000 108.6000 ;
	    RECT 1511.4000 77.4000 1512.6000 78.6000 ;
	    RECT 1513.8000 65.4000 1515.0000 66.6000 ;
	    RECT 1511.4000 53.4000 1512.6000 54.6000 ;
	    RECT 1511.5500 48.6000 1512.4501 53.4000 ;
	    RECT 1513.9501 48.6000 1514.8500 65.4000 ;
	    RECT 1516.3500 60.6000 1517.2500 137.4000 ;
	    RECT 1518.7500 72.6000 1519.6500 167.4000 ;
	    RECT 1523.5500 156.6000 1524.4501 170.5500 ;
	    RECT 1525.8000 170.4000 1527.0000 170.5500 ;
	    RECT 1528.3500 165.6000 1529.2500 191.4000 ;
	    RECT 1530.7500 168.6000 1531.6500 197.4000 ;
	    RECT 1542.7500 186.6000 1543.6500 203.4000 ;
	    RECT 1557.0000 200.4000 1558.2001 201.6000 ;
	    RECT 1554.6000 197.4000 1555.8000 198.6000 ;
	    RECT 1542.6000 185.4000 1543.8000 186.6000 ;
	    RECT 1542.7500 168.6000 1543.6500 185.4000 ;
	    RECT 1554.7500 171.6000 1555.6500 197.4000 ;
	    RECT 1554.6000 170.4000 1555.8000 171.6000 ;
	    RECT 1530.6000 167.4000 1531.8000 168.6000 ;
	    RECT 1542.6000 167.4000 1543.8000 168.6000 ;
	    RECT 1528.2001 164.4000 1529.4000 165.6000 ;
	    RECT 1545.0000 161.4000 1546.2001 162.6000 ;
	    RECT 1523.4000 155.4000 1524.6000 156.6000 ;
	    RECT 1540.2001 140.4000 1541.4000 141.6000 ;
	    RECT 1523.4000 137.4000 1524.6000 138.6000 ;
	    RECT 1521.0000 101.4000 1522.2001 102.6000 ;
	    RECT 1521.1500 75.6000 1522.0500 101.4000 ;
	    RECT 1523.5500 99.6000 1524.4501 137.4000 ;
	    RECT 1540.3500 105.6000 1541.2500 140.4000 ;
	    RECT 1540.2001 104.4000 1541.4000 105.6000 ;
	    RECT 1523.4000 98.4000 1524.6000 99.6000 ;
	    RECT 1523.4000 77.4000 1524.6000 78.6000 ;
	    RECT 1521.0000 74.4000 1522.2001 75.6000 ;
	    RECT 1518.6000 71.4000 1519.8000 72.6000 ;
	    RECT 1516.2001 59.4000 1517.4000 60.6000 ;
	    RECT 1521.1500 48.6000 1522.0500 74.4000 ;
	    RECT 1523.5500 72.6000 1524.4501 77.4000 ;
	    RECT 1545.1500 75.6000 1546.0500 161.4000 ;
	    RECT 1554.7500 141.6000 1555.6500 170.4000 ;
	    RECT 1557.1500 165.6000 1558.0500 200.4000 ;
	    RECT 1561.9501 168.6000 1562.8500 209.4000 ;
	    RECT 1561.8000 167.4000 1563.0000 168.6000 ;
	    RECT 1557.0000 164.4000 1558.2001 165.6000 ;
	    RECT 1557.1500 162.6000 1558.0500 164.4000 ;
	    RECT 1557.0000 161.4000 1558.2001 162.6000 ;
	    RECT 1554.6000 140.4000 1555.8000 141.6000 ;
	    RECT 1557.0000 134.4000 1558.2001 135.6000 ;
	    RECT 1547.4000 119.4000 1548.6000 120.6000 ;
	    RECT 1547.5500 102.6000 1548.4501 119.4000 ;
	    RECT 1549.8000 104.4000 1551.0000 105.6000 ;
	    RECT 1547.4000 101.4000 1548.6000 102.6000 ;
	    RECT 1549.9501 84.6000 1550.8500 104.4000 ;
	    RECT 1549.8000 83.4000 1551.0000 84.6000 ;
	    RECT 1554.6000 77.4000 1555.8000 78.6000 ;
	    RECT 1545.0000 74.4000 1546.2001 75.6000 ;
	    RECT 1547.4000 74.4000 1548.6000 75.6000 ;
	    RECT 1547.5500 72.6000 1548.4501 74.4000 ;
	    RECT 1523.4000 71.4000 1524.6000 72.6000 ;
	    RECT 1525.8000 71.4000 1527.0000 72.6000 ;
	    RECT 1547.4000 71.4000 1548.6000 72.6000 ;
	    RECT 1523.5500 54.6000 1524.4501 71.4000 ;
	    RECT 1525.9501 66.6000 1526.8500 71.4000 ;
	    RECT 1554.7500 66.6000 1555.6500 77.4000 ;
	    RECT 1557.1500 72.6000 1558.0500 134.4000 ;
	    RECT 1564.3500 75.6000 1565.2500 293.4000 ;
	    RECT 1566.7500 258.6000 1567.6500 347.4000 ;
	    RECT 1566.6000 257.4000 1567.8000 258.6000 ;
	    RECT 1564.2001 74.4000 1565.4000 75.6000 ;
	    RECT 1557.0000 71.4000 1558.2001 72.6000 ;
	    RECT 1525.8000 65.4000 1527.0000 66.6000 ;
	    RECT 1554.6000 65.4000 1555.8000 66.6000 ;
	    RECT 1525.8000 59.4000 1527.0000 60.6000 ;
	    RECT 1523.4000 53.4000 1524.6000 54.6000 ;
	    RECT 1511.4000 47.4000 1512.6000 48.6000 ;
	    RECT 1513.8000 47.4000 1515.0000 48.6000 ;
	    RECT 1521.0000 47.4000 1522.2001 48.6000 ;
	    RECT 1525.9501 42.6000 1526.8500 59.4000 ;
	    RECT 1554.6000 47.4000 1555.8000 48.6000 ;
	    RECT 1530.6000 44.4000 1531.8000 45.6000 ;
	    RECT 1552.2001 44.4000 1553.4000 45.6000 ;
	    RECT 1525.8000 41.4000 1527.0000 42.6000 ;
	    RECT 1509.0000 35.4000 1510.2001 36.6000 ;
	    RECT 1485.0000 30.4500 1486.2001 30.6000 ;
	    RECT 1482.7500 29.5500 1486.2001 30.4500 ;
	    RECT 1485.0000 29.4000 1486.2001 29.5500 ;
	    RECT 1329.0000 23.4000 1330.2001 24.6000 ;
	    RECT 1372.2001 23.4000 1373.4000 24.6000 ;
	    RECT 1470.6000 23.4000 1471.8000 24.6000 ;
	    RECT 1305.0000 20.4000 1306.2001 21.6000 ;
	    RECT 1307.4000 20.4000 1308.6000 21.6000 ;
	    RECT 1470.7500 18.6000 1471.6500 23.4000 ;
	    RECT 1302.6000 17.4000 1303.8000 18.6000 ;
	    RECT 1470.6000 17.4000 1471.8000 18.6000 ;
	    RECT 1297.8000 14.4000 1299.0000 15.6000 ;
	    RECT 1465.8000 14.4000 1467.0000 15.6000 ;
	    RECT 1254.6000 11.4000 1255.8000 12.6000 ;
	    RECT 1465.9501 6.6000 1466.8500 14.4000 ;
	    RECT 1465.8000 5.4000 1467.0000 6.6000 ;
	    RECT 1473.0000 6.3000 1474.2001 26.7000 ;
	    RECT 1475.4000 6.3000 1476.6000 26.7000 ;
	    RECT 1477.8000 9.3000 1479.0000 26.7000 ;
	    RECT 1480.2001 20.4000 1481.4000 21.6000 ;
	    RECT 1480.3500 18.6000 1481.2500 20.4000 ;
	    RECT 1480.2001 17.4000 1481.4000 18.6000 ;
	    RECT 1482.6000 9.3000 1483.8000 26.7000 ;
	    RECT 1485.1500 24.6000 1486.0500 29.4000 ;
	    RECT 1485.0000 23.4000 1486.2001 24.6000 ;
	    RECT 1487.4000 9.3000 1488.6000 26.7000 ;
	    RECT 1489.8000 6.3000 1491.0000 26.7000 ;
	    RECT 1492.2001 6.3000 1493.4000 26.7000 ;
	    RECT 1494.6000 6.3000 1495.8000 26.7000 ;
	    RECT 1511.4000 20.4000 1512.6000 21.6000 ;
	    RECT 1511.5500 18.6000 1512.4501 20.4000 ;
	    RECT 1511.4000 17.4000 1512.6000 18.6000 ;
	    RECT 1516.2001 17.4000 1517.4000 18.6000 ;
	    RECT 1516.3500 12.6000 1517.2500 17.4000 ;
	    RECT 1530.7500 15.6000 1531.6500 44.4000 ;
	    RECT 1552.3500 24.6000 1553.2500 44.4000 ;
	    RECT 1554.7500 39.6000 1555.6500 47.4000 ;
	    RECT 1557.1500 42.6000 1558.0500 71.4000 ;
	    RECT 1557.0000 41.4000 1558.2001 42.6000 ;
	    RECT 1554.6000 38.4000 1555.8000 39.6000 ;
	    RECT 1552.2001 23.4000 1553.4000 24.6000 ;
	    RECT 1542.6000 20.4000 1543.8000 21.6000 ;
	    RECT 1530.6000 14.4000 1531.8000 15.6000 ;
	    RECT 1516.2001 11.4000 1517.4000 12.6000 ;
	    RECT 1542.7500 6.6000 1543.6500 20.4000 ;
	    RECT 1552.3500 18.6000 1553.2500 23.4000 ;
	    RECT 1552.2001 17.4000 1553.4000 18.6000 ;
	    RECT 1542.6000 5.4000 1543.8000 6.6000 ;
	    RECT 1566.6000 5.4000 1567.8000 6.6000 ;
	    RECT 1566.7500 3.6000 1567.6500 5.4000 ;
	    RECT 1566.6000 2.4000 1567.8000 3.6000 ;
         LAYER metal3 ;
	    RECT 145.5000 1464.7500 147.3000 1464.9000 ;
	    RECT 224.7000 1464.7500 226.5000 1464.9000 ;
	    RECT 145.5000 1463.2500 226.5000 1464.7500 ;
	    RECT 145.5000 1463.1000 147.3000 1463.2500 ;
	    RECT 224.7000 1463.1000 226.5000 1463.2500 ;
	    RECT 702.3000 1464.7500 704.1000 1464.9000 ;
	    RECT 879.9000 1464.7500 881.7000 1464.9000 ;
	    RECT 702.3000 1463.2500 881.7000 1464.7500 ;
	    RECT 702.3000 1463.1000 704.1000 1463.2500 ;
	    RECT 879.9000 1463.1000 881.7000 1463.2500 ;
	    RECT 884.7000 1464.7500 886.5000 1464.9000 ;
	    RECT 906.3000 1464.7500 908.1000 1464.9000 ;
	    RECT 884.7000 1463.2500 908.1000 1464.7500 ;
	    RECT 884.7000 1463.1000 886.5000 1463.2500 ;
	    RECT 906.3000 1463.1000 908.1000 1463.2500 ;
	    RECT 1095.9000 1464.7500 1097.7001 1464.9000 ;
	    RECT 1139.1000 1464.7500 1140.9000 1464.9000 ;
	    RECT 1095.9000 1463.2500 1140.9000 1464.7500 ;
	    RECT 1095.9000 1463.1000 1097.7001 1463.2500 ;
	    RECT 1139.1000 1463.1000 1140.9000 1463.2500 ;
	    RECT 1311.9000 1464.7500 1313.7001 1464.9000 ;
	    RECT 1333.5000 1464.7500 1335.3000 1464.9000 ;
	    RECT 1311.9000 1463.2500 1335.3000 1464.7500 ;
	    RECT 1311.9000 1463.1000 1313.7001 1463.2500 ;
	    RECT 1333.5000 1463.1000 1335.3000 1463.2500 ;
	    RECT 1446.3000 1464.7500 1448.1000 1464.9000 ;
	    RECT 1487.1000 1464.7500 1488.9000 1464.9000 ;
	    RECT 1446.3000 1463.2500 1488.9000 1464.7500 ;
	    RECT 1446.3000 1463.1000 1448.1000 1463.2500 ;
	    RECT 1487.1000 1463.1000 1488.9000 1463.2500 ;
	    RECT 135.9000 1458.7500 137.7000 1458.9000 ;
	    RECT 164.7000 1458.7500 166.5000 1458.9000 ;
	    RECT 135.9000 1457.2500 166.5000 1458.7500 ;
	    RECT 135.9000 1457.1000 137.7000 1457.2500 ;
	    RECT 164.7000 1457.1000 166.5000 1457.2500 ;
	    RECT 222.3000 1458.7500 224.1000 1458.9000 ;
	    RECT 227.1000 1458.7500 228.9000 1458.9000 ;
	    RECT 222.3000 1457.2500 228.9000 1458.7500 ;
	    RECT 222.3000 1457.1000 224.1000 1457.2500 ;
	    RECT 227.1000 1457.1000 228.9000 1457.2500 ;
	    RECT 231.9000 1458.7500 233.7000 1458.9000 ;
	    RECT 255.9000 1458.7500 257.7000 1458.9000 ;
	    RECT 270.3000 1458.7500 272.1000 1458.9000 ;
	    RECT 303.9000 1458.7500 305.7000 1458.9000 ;
	    RECT 231.9000 1457.2500 305.7000 1458.7500 ;
	    RECT 231.9000 1457.1000 233.7000 1457.2500 ;
	    RECT 255.9000 1457.1000 257.7000 1457.2500 ;
	    RECT 270.3000 1457.1000 272.1000 1457.2500 ;
	    RECT 303.9000 1457.1000 305.7000 1457.2500 ;
	    RECT 651.9000 1458.7500 653.7000 1458.9000 ;
	    RECT 697.5000 1458.7500 699.3000 1458.9000 ;
	    RECT 651.9000 1457.2500 699.3000 1458.7500 ;
	    RECT 651.9000 1457.1000 653.7000 1457.2500 ;
	    RECT 697.5000 1457.1000 699.3000 1457.2500 ;
	    RECT 1043.1000 1458.7500 1044.9000 1458.9000 ;
	    RECT 1110.3000 1458.7500 1112.1000 1458.9000 ;
	    RECT 1043.1000 1457.2500 1112.1000 1458.7500 ;
	    RECT 1043.1000 1457.1000 1044.9000 1457.2500 ;
	    RECT 1110.3000 1457.1000 1112.1000 1457.2500 ;
	    RECT 191.1000 1452.7500 192.9000 1452.9000 ;
	    RECT 251.1000 1452.7500 252.9000 1452.9000 ;
	    RECT 191.1000 1451.2500 252.9000 1452.7500 ;
	    RECT 191.1000 1451.1000 192.9000 1451.2500 ;
	    RECT 251.1000 1451.1000 252.9000 1451.2500 ;
	    RECT 265.5000 1452.7500 267.3000 1452.9000 ;
	    RECT 296.7000 1452.7500 298.5000 1452.9000 ;
	    RECT 265.5000 1451.2500 298.5000 1452.7500 ;
	    RECT 265.5000 1451.1000 267.3000 1451.2500 ;
	    RECT 296.7000 1451.1000 298.5000 1451.2500 ;
	    RECT 407.1000 1452.7500 408.9000 1452.9000 ;
	    RECT 455.1000 1452.7500 456.9000 1452.9000 ;
	    RECT 407.1000 1451.2500 456.9000 1452.7500 ;
	    RECT 407.1000 1451.1000 408.9000 1451.2500 ;
	    RECT 455.1000 1451.1000 456.9000 1451.2500 ;
	    RECT 757.5000 1452.7500 759.3000 1452.9000 ;
	    RECT 894.3000 1452.7500 896.1000 1452.9000 ;
	    RECT 944.7000 1452.7500 946.5000 1452.9000 ;
	    RECT 757.5000 1451.2500 946.5000 1452.7500 ;
	    RECT 757.5000 1451.1000 759.3000 1451.2500 ;
	    RECT 894.3000 1451.1000 896.1000 1451.2500 ;
	    RECT 944.7000 1451.1000 946.5000 1451.2500 ;
	    RECT 1100.7001 1452.7500 1102.5000 1452.9000 ;
	    RECT 1110.3000 1452.7500 1112.1000 1452.9000 ;
	    RECT 1100.7001 1451.2500 1112.1000 1452.7500 ;
	    RECT 1100.7001 1451.1000 1102.5000 1451.2500 ;
	    RECT 1110.3000 1451.1000 1112.1000 1451.2500 ;
	    RECT 505.5000 1446.7500 507.3000 1446.9000 ;
	    RECT 747.9000 1446.7500 749.7000 1446.9000 ;
	    RECT 505.5000 1445.2500 749.7000 1446.7500 ;
	    RECT 505.5000 1445.1000 507.3000 1445.2500 ;
	    RECT 747.9000 1445.1000 749.7000 1445.2500 ;
	    RECT 855.9000 1446.7500 857.7000 1446.9000 ;
	    RECT 882.3000 1446.7500 884.1000 1446.9000 ;
	    RECT 855.9000 1445.2500 884.1000 1446.7500 ;
	    RECT 855.9000 1445.1000 857.7000 1445.2500 ;
	    RECT 882.3000 1445.1000 884.1000 1445.2500 ;
	    RECT 944.7000 1446.7500 946.5000 1446.9000 ;
	    RECT 1095.9000 1446.7500 1097.7001 1446.9000 ;
	    RECT 944.7000 1445.2500 1097.7001 1446.7500 ;
	    RECT 944.7000 1445.1000 946.5000 1445.2500 ;
	    RECT 1095.9000 1445.1000 1097.7001 1445.2500 ;
	    RECT 536.7000 1440.7500 538.5000 1440.9000 ;
	    RECT 654.3000 1440.7500 656.1000 1440.9000 ;
	    RECT 536.7000 1439.2500 656.1000 1440.7500 ;
	    RECT 536.7000 1439.1000 538.5000 1439.2500 ;
	    RECT 654.3000 1439.1000 656.1000 1439.2500 ;
	    RECT 899.1000 1440.7500 900.9000 1440.9000 ;
	    RECT 906.3000 1440.7500 908.1000 1440.9000 ;
	    RECT 899.1000 1439.2500 908.1000 1440.7500 ;
	    RECT 899.1000 1439.1000 900.9000 1439.2500 ;
	    RECT 906.3000 1439.1000 908.1000 1439.2500 ;
	    RECT 1067.1000 1440.7500 1068.9000 1440.9000 ;
	    RECT 1100.7001 1440.7500 1102.5000 1440.9000 ;
	    RECT 1067.1000 1439.2500 1102.5000 1440.7500 ;
	    RECT 1067.1000 1439.1000 1068.9000 1439.2500 ;
	    RECT 1100.7001 1439.1000 1102.5000 1439.2500 ;
	    RECT 1491.9000 1440.7500 1493.7001 1440.9000 ;
	    RECT 1496.7001 1440.7500 1498.5000 1440.9000 ;
	    RECT 1491.9000 1439.2500 1498.5000 1440.7500 ;
	    RECT 1491.9000 1439.1000 1493.7001 1439.2500 ;
	    RECT 1496.7001 1439.1000 1498.5000 1439.2500 ;
	    RECT 291.9000 1434.7500 293.7000 1434.9000 ;
	    RECT 337.5000 1434.7500 339.3000 1434.9000 ;
	    RECT 291.9000 1433.2500 339.3000 1434.7500 ;
	    RECT 291.9000 1433.1000 293.7000 1433.2500 ;
	    RECT 337.5000 1433.1000 339.3000 1433.2500 ;
	    RECT 1479.9000 1434.7500 1481.7001 1434.9000 ;
	    RECT 1494.3000 1434.7500 1496.1000 1434.9000 ;
	    RECT 1479.9000 1433.2500 1496.1000 1434.7500 ;
	    RECT 1479.9000 1433.1000 1481.7001 1433.2500 ;
	    RECT 1494.3000 1433.1000 1496.1000 1433.2500 ;
	    RECT 133.5000 1428.7500 135.3000 1428.9000 ;
	    RECT 347.1000 1428.7500 348.9000 1428.9000 ;
	    RECT 133.5000 1427.2500 348.9000 1428.7500 ;
	    RECT 133.5000 1427.1000 135.3000 1427.2500 ;
	    RECT 347.1000 1427.1000 348.9000 1427.2500 ;
	    RECT 380.7000 1428.7500 382.5000 1428.9000 ;
	    RECT 426.3000 1428.7500 428.1000 1428.9000 ;
	    RECT 491.1000 1428.7500 492.9000 1428.9000 ;
	    RECT 380.7000 1427.2500 492.9000 1428.7500 ;
	    RECT 380.7000 1427.1000 382.5000 1427.2500 ;
	    RECT 426.3000 1427.1000 428.1000 1427.2500 ;
	    RECT 491.1000 1427.1000 492.9000 1427.2500 ;
	    RECT 649.5000 1428.7500 651.3000 1428.9000 ;
	    RECT 659.1000 1428.7500 660.9000 1428.9000 ;
	    RECT 649.5000 1427.2500 660.9000 1428.7500 ;
	    RECT 649.5000 1427.1000 651.3000 1427.2500 ;
	    RECT 659.1000 1427.1000 660.9000 1427.2500 ;
	    RECT 675.9000 1428.7500 677.7000 1428.9000 ;
	    RECT 680.7000 1428.7500 682.5000 1428.9000 ;
	    RECT 675.9000 1427.2500 682.5000 1428.7500 ;
	    RECT 675.9000 1427.1000 677.7000 1427.2500 ;
	    RECT 680.7000 1427.1000 682.5000 1427.2500 ;
	    RECT 697.5000 1428.7500 699.3000 1428.9000 ;
	    RECT 726.3000 1428.7500 728.1000 1428.9000 ;
	    RECT 697.5000 1427.2500 728.1000 1428.7500 ;
	    RECT 697.5000 1427.1000 699.3000 1427.2500 ;
	    RECT 726.3000 1427.1000 728.1000 1427.2500 ;
	    RECT 903.9000 1428.7500 905.7000 1428.9000 ;
	    RECT 937.5000 1428.7500 939.3000 1428.9000 ;
	    RECT 903.9000 1427.2500 939.3000 1428.7500 ;
	    RECT 903.9000 1427.1000 905.7000 1427.2500 ;
	    RECT 937.5000 1427.1000 939.3000 1427.2500 ;
	    RECT 1057.5000 1428.7500 1059.3000 1428.9000 ;
	    RECT 1086.3000 1428.7500 1088.1000 1428.9000 ;
	    RECT 1057.5000 1427.2500 1088.1000 1428.7500 ;
	    RECT 1057.5000 1427.1000 1059.3000 1427.2500 ;
	    RECT 1086.3000 1427.1000 1088.1000 1427.2500 ;
	    RECT 1177.5000 1428.7500 1179.3000 1428.9000 ;
	    RECT 1302.3000 1428.7500 1304.1000 1428.9000 ;
	    RECT 1177.5000 1427.2500 1304.1000 1428.7500 ;
	    RECT 1177.5000 1427.1000 1179.3000 1427.2500 ;
	    RECT 1302.3000 1427.1000 1304.1000 1427.2500 ;
	    RECT 49.5000 1422.7500 51.3000 1422.9000 ;
	    RECT 143.1000 1422.7500 144.9000 1422.9000 ;
	    RECT 49.5000 1421.2500 144.9000 1422.7500 ;
	    RECT 49.5000 1421.1000 51.3000 1421.2500 ;
	    RECT 143.1000 1421.1000 144.9000 1421.2500 ;
	    RECT 311.1000 1422.7500 312.9000 1422.9000 ;
	    RECT 375.9000 1422.7500 377.7000 1422.9000 ;
	    RECT 311.1000 1421.2500 377.7000 1422.7500 ;
	    RECT 311.1000 1421.1000 312.9000 1421.2500 ;
	    RECT 375.9000 1421.1000 377.7000 1421.2500 ;
	    RECT 414.3000 1422.7500 416.1000 1422.9000 ;
	    RECT 459.9000 1422.7500 461.7000 1422.9000 ;
	    RECT 474.3000 1422.7500 476.1000 1422.9000 ;
	    RECT 414.3000 1421.2500 476.1000 1422.7500 ;
	    RECT 414.3000 1421.1000 416.1000 1421.2500 ;
	    RECT 459.9000 1421.1000 461.7000 1421.2500 ;
	    RECT 474.3000 1421.1000 476.1000 1421.2500 ;
	    RECT 560.7000 1422.7500 562.5000 1422.9000 ;
	    RECT 606.3000 1422.7500 608.1000 1422.9000 ;
	    RECT 560.7000 1421.2500 608.1000 1422.7500 ;
	    RECT 560.7000 1421.1000 562.5000 1421.2500 ;
	    RECT 606.3000 1421.1000 608.1000 1421.2500 ;
	    RECT 647.1000 1422.7500 648.9000 1422.9000 ;
	    RECT 675.9000 1422.7500 677.7000 1422.9000 ;
	    RECT 647.1000 1421.2500 677.7000 1422.7500 ;
	    RECT 647.1000 1421.1000 648.9000 1421.2500 ;
	    RECT 675.9000 1421.1000 677.7000 1421.2500 ;
	    RECT 1122.3000 1422.7500 1124.1000 1422.9000 ;
	    RECT 1143.9000 1422.7500 1145.7001 1422.9000 ;
	    RECT 1122.3000 1421.2500 1145.7001 1422.7500 ;
	    RECT 1122.3000 1421.1000 1124.1000 1421.2500 ;
	    RECT 1143.9000 1421.1000 1145.7001 1421.2500 ;
	    RECT 1285.5000 1422.7500 1287.3000 1422.9000 ;
	    RECT 1297.5000 1422.7500 1299.3000 1422.9000 ;
	    RECT 1285.5000 1421.2500 1299.3000 1422.7500 ;
	    RECT 1285.5000 1421.1000 1287.3000 1421.2500 ;
	    RECT 1297.5000 1421.1000 1299.3000 1421.2500 ;
	    RECT 159.9000 1416.7500 161.7000 1416.9000 ;
	    RECT 176.7000 1416.7500 178.5000 1416.9000 ;
	    RECT 159.9000 1415.2500 178.5000 1416.7500 ;
	    RECT 159.9000 1415.1000 161.7000 1415.2500 ;
	    RECT 176.7000 1415.1000 178.5000 1415.2500 ;
	    RECT 459.9000 1416.7500 461.7000 1416.9000 ;
	    RECT 505.5000 1416.7500 507.3000 1416.9000 ;
	    RECT 459.9000 1415.2500 507.3000 1416.7500 ;
	    RECT 459.9000 1415.1000 461.7000 1415.2500 ;
	    RECT 505.5000 1415.1000 507.3000 1415.2500 ;
	    RECT 577.5000 1416.7500 579.3000 1416.9000 ;
	    RECT 589.5000 1416.7500 591.3000 1416.9000 ;
	    RECT 577.5000 1415.2500 591.3000 1416.7500 ;
	    RECT 577.5000 1415.1000 579.3000 1415.2500 ;
	    RECT 589.5000 1415.1000 591.3000 1415.2500 ;
	    RECT 649.5000 1416.7500 651.3000 1416.9000 ;
	    RECT 656.7000 1416.7500 658.5000 1416.9000 ;
	    RECT 649.5000 1415.2500 658.5000 1416.7500 ;
	    RECT 649.5000 1415.1000 651.3000 1415.2500 ;
	    RECT 656.7000 1415.1000 658.5000 1415.2500 ;
	    RECT 675.9000 1416.7500 677.7000 1416.9000 ;
	    RECT 695.1000 1416.7500 696.9000 1416.9000 ;
	    RECT 675.9000 1415.2500 696.9000 1416.7500 ;
	    RECT 675.9000 1415.1000 677.7000 1415.2500 ;
	    RECT 695.1000 1415.1000 696.9000 1415.2500 ;
	    RECT 723.9000 1416.7500 725.7000 1416.9000 ;
	    RECT 848.7000 1416.7500 850.5000 1416.9000 ;
	    RECT 723.9000 1415.2500 850.5000 1416.7500 ;
	    RECT 723.9000 1415.1000 725.7000 1415.2500 ;
	    RECT 848.7000 1415.1000 850.5000 1415.2500 ;
	    RECT 853.5000 1416.7500 855.3000 1416.9000 ;
	    RECT 872.7000 1416.7500 874.5000 1416.9000 ;
	    RECT 879.9000 1416.7500 881.7000 1416.9000 ;
	    RECT 853.5000 1415.2500 881.7000 1416.7500 ;
	    RECT 853.5000 1415.1000 855.3000 1415.2500 ;
	    RECT 872.7000 1415.1000 874.5000 1415.2500 ;
	    RECT 879.9000 1415.1000 881.7000 1415.2500 ;
	    RECT 315.9000 1410.7500 317.7000 1410.9000 ;
	    RECT 380.7000 1410.7500 382.5000 1410.9000 ;
	    RECT 315.9000 1409.2500 382.5000 1410.7500 ;
	    RECT 315.9000 1409.1000 317.7000 1409.2500 ;
	    RECT 380.7000 1409.1000 382.5000 1409.2500 ;
	    RECT 471.9000 1410.7500 473.7000 1410.9000 ;
	    RECT 495.9000 1410.7500 497.7000 1410.9000 ;
	    RECT 471.9000 1409.2500 497.7000 1410.7500 ;
	    RECT 471.9000 1409.1000 473.7000 1409.2500 ;
	    RECT 495.9000 1409.1000 497.7000 1409.2500 ;
	    RECT 654.3000 1410.7500 656.1000 1410.9000 ;
	    RECT 666.3000 1410.7500 668.1000 1410.9000 ;
	    RECT 654.3000 1409.2500 668.1000 1410.7500 ;
	    RECT 654.3000 1409.1000 656.1000 1409.2500 ;
	    RECT 666.3000 1409.1000 668.1000 1409.2500 ;
	    RECT 755.1000 1410.7500 756.9000 1410.9000 ;
	    RECT 877.5000 1410.7500 879.3000 1410.9000 ;
	    RECT 755.1000 1409.2500 879.3000 1410.7500 ;
	    RECT 755.1000 1409.1000 756.9000 1409.2500 ;
	    RECT 877.5000 1409.1000 879.3000 1409.2500 ;
	    RECT 1513.5000 1410.7500 1515.3000 1410.9000 ;
	    RECT 1539.9000 1410.7500 1541.7001 1410.9000 ;
	    RECT 1559.1000 1410.7500 1560.9000 1410.9000 ;
	    RECT 1513.5000 1409.2500 1560.9000 1410.7500 ;
	    RECT 1513.5000 1409.1000 1515.3000 1409.2500 ;
	    RECT 1539.9000 1409.1000 1541.7001 1409.2500 ;
	    RECT 1559.1000 1409.1000 1560.9000 1409.2500 ;
	    RECT 462.3000 1404.7500 464.1000 1404.9000 ;
	    RECT 491.1000 1404.7500 492.9000 1404.9000 ;
	    RECT 462.3000 1403.2500 492.9000 1404.7500 ;
	    RECT 462.3000 1403.1000 464.1000 1403.2500 ;
	    RECT 491.1000 1403.1000 492.9000 1403.2500 ;
	    RECT 930.3000 1404.7500 932.1000 1404.9000 ;
	    RECT 975.9000 1404.7500 977.7000 1404.9000 ;
	    RECT 930.3000 1403.2500 977.7000 1404.7500 ;
	    RECT 930.3000 1403.1000 932.1000 1403.2500 ;
	    RECT 975.9000 1403.1000 977.7000 1403.2500 ;
	    RECT 992.7000 1404.7500 994.5000 1404.9000 ;
	    RECT 1011.9000 1404.7500 1013.7000 1404.9000 ;
	    RECT 1031.1000 1404.7500 1032.9000 1404.9000 ;
	    RECT 992.7000 1403.2500 1032.9000 1404.7500 ;
	    RECT 992.7000 1403.1000 994.5000 1403.2500 ;
	    RECT 1011.9000 1403.1000 1013.7000 1403.2500 ;
	    RECT 1031.1000 1403.1000 1032.9000 1403.2500 ;
	    RECT 1069.5000 1404.7500 1071.3000 1404.9000 ;
	    RECT 1091.1000 1404.7500 1092.9000 1404.9000 ;
	    RECT 1069.5000 1403.2500 1092.9000 1404.7500 ;
	    RECT 1069.5000 1403.1000 1071.3000 1403.2500 ;
	    RECT 1091.1000 1403.1000 1092.9000 1403.2500 ;
	    RECT 1139.1000 1404.7500 1140.9000 1404.9000 ;
	    RECT 1287.9000 1404.7500 1289.7001 1404.9000 ;
	    RECT 1316.7001 1404.7500 1318.5000 1404.9000 ;
	    RECT 1479.9000 1404.7500 1481.7001 1404.9000 ;
	    RECT 1496.7001 1404.7500 1498.5000 1404.9000 ;
	    RECT 1535.1000 1404.7500 1536.9000 1404.9000 ;
	    RECT 1139.1000 1403.2500 1536.9000 1404.7500 ;
	    RECT 1139.1000 1403.1000 1140.9000 1403.2500 ;
	    RECT 1287.9000 1403.1000 1289.7001 1403.2500 ;
	    RECT 1316.7001 1403.1000 1318.5000 1403.2500 ;
	    RECT 1479.9000 1403.1000 1481.7001 1403.2500 ;
	    RECT 1496.7001 1403.1000 1498.5000 1403.2500 ;
	    RECT 1535.1000 1403.1000 1536.9000 1403.2500 ;
	    RECT 169.5000 1398.7500 171.3000 1398.9000 ;
	    RECT 174.3000 1398.7500 176.1000 1398.9000 ;
	    RECT 169.5000 1397.2500 176.1000 1398.7500 ;
	    RECT 169.5000 1397.1000 171.3000 1397.2500 ;
	    RECT 174.3000 1397.1000 176.1000 1397.2500 ;
	    RECT 265.5000 1398.7500 267.3000 1398.9000 ;
	    RECT 284.7000 1398.7500 286.5000 1398.9000 ;
	    RECT 265.5000 1397.2500 286.5000 1398.7500 ;
	    RECT 265.5000 1397.1000 267.3000 1397.2500 ;
	    RECT 284.7000 1397.1000 286.5000 1397.2500 ;
	    RECT 428.7000 1398.7500 430.5000 1398.9000 ;
	    RECT 505.5000 1398.7500 507.3000 1398.9000 ;
	    RECT 428.7000 1397.2500 507.3000 1398.7500 ;
	    RECT 428.7000 1397.1000 430.5000 1397.2500 ;
	    RECT 505.5000 1397.1000 507.3000 1397.2500 ;
	    RECT 728.7000 1398.7500 730.5000 1398.9000 ;
	    RECT 743.1000 1398.7500 744.9000 1398.9000 ;
	    RECT 728.7000 1397.2500 744.9000 1398.7500 ;
	    RECT 728.7000 1397.1000 730.5000 1397.2500 ;
	    RECT 743.1000 1397.1000 744.9000 1397.2500 ;
	    RECT 913.5000 1398.7500 915.3000 1398.9000 ;
	    RECT 930.3000 1398.7500 932.1000 1398.9000 ;
	    RECT 913.5000 1397.2500 932.1000 1398.7500 ;
	    RECT 913.5000 1397.1000 915.3000 1397.2500 ;
	    RECT 930.3000 1397.1000 932.1000 1397.2500 ;
	    RECT 975.9000 1398.7500 977.7000 1398.9000 ;
	    RECT 992.7000 1398.7500 994.5000 1398.9000 ;
	    RECT 975.9000 1397.2500 994.5000 1398.7500 ;
	    RECT 975.9000 1397.1000 977.7000 1397.2500 ;
	    RECT 992.7000 1397.1000 994.5000 1397.2500 ;
	    RECT 1055.1000 1398.7500 1056.9000 1398.9000 ;
	    RECT 1062.3000 1398.7500 1064.1000 1398.9000 ;
	    RECT 1055.1000 1397.2500 1064.1000 1398.7500 ;
	    RECT 1055.1000 1397.1000 1056.9000 1397.2500 ;
	    RECT 1062.3000 1397.1000 1064.1000 1397.2500 ;
	    RECT 1331.1000 1398.7500 1332.9000 1398.9000 ;
	    RECT 1345.5000 1398.7500 1347.3000 1398.9000 ;
	    RECT 1331.1000 1397.2500 1347.3000 1398.7500 ;
	    RECT 1331.1000 1397.1000 1332.9000 1397.2500 ;
	    RECT 1345.5000 1397.1000 1347.3000 1397.2500 ;
	    RECT 164.7000 1392.7500 166.5000 1392.9000 ;
	    RECT 169.5000 1392.7500 171.3000 1392.9000 ;
	    RECT 164.7000 1391.2500 171.3000 1392.7500 ;
	    RECT 164.7000 1391.1000 166.5000 1391.2500 ;
	    RECT 169.5000 1391.1000 171.3000 1391.2500 ;
	    RECT 195.9000 1392.7500 197.7000 1392.9000 ;
	    RECT 203.1000 1392.7500 204.9000 1392.9000 ;
	    RECT 195.9000 1391.2500 204.9000 1392.7500 ;
	    RECT 195.9000 1391.1000 197.7000 1391.2500 ;
	    RECT 203.1000 1391.1000 204.9000 1391.2500 ;
	    RECT 315.9000 1392.7500 317.7000 1392.9000 ;
	    RECT 330.3000 1392.7500 332.1000 1392.9000 ;
	    RECT 455.1000 1392.7500 456.9000 1392.9000 ;
	    RECT 315.9000 1391.2500 456.9000 1392.7500 ;
	    RECT 315.9000 1391.1000 317.7000 1391.2500 ;
	    RECT 330.3000 1391.1000 332.1000 1391.2500 ;
	    RECT 455.1000 1391.1000 456.9000 1391.2500 ;
	    RECT 944.7000 1392.7500 946.5000 1392.9000 ;
	    RECT 968.7000 1392.7500 970.5000 1392.9000 ;
	    RECT 944.7000 1391.2500 970.5000 1392.7500 ;
	    RECT 944.7000 1391.1000 946.5000 1391.2500 ;
	    RECT 968.7000 1391.1000 970.5000 1391.2500 ;
	    RECT 1057.5000 1392.7500 1059.3000 1392.9000 ;
	    RECT 1064.7001 1392.7500 1066.5000 1392.9000 ;
	    RECT 1057.5000 1391.2500 1066.5000 1392.7500 ;
	    RECT 1057.5000 1391.1000 1059.3000 1391.2500 ;
	    RECT 1064.7001 1391.1000 1066.5000 1391.2500 ;
	    RECT 198.3000 1386.7500 200.1000 1386.9000 ;
	    RECT 234.3000 1386.7500 236.1000 1386.9000 ;
	    RECT 198.3000 1385.2500 236.1000 1386.7500 ;
	    RECT 198.3000 1385.1000 200.1000 1385.2500 ;
	    RECT 234.3000 1385.1000 236.1000 1385.2500 ;
	    RECT 644.7000 1386.7500 646.5000 1386.9000 ;
	    RECT 671.1000 1386.7500 672.9000 1386.9000 ;
	    RECT 644.7000 1385.2500 672.9000 1386.7500 ;
	    RECT 644.7000 1385.1000 646.5000 1385.2500 ;
	    RECT 671.1000 1385.1000 672.9000 1385.2500 ;
	    RECT 956.7000 1386.7500 958.5000 1386.9000 ;
	    RECT 1127.1000 1386.7500 1128.9000 1386.9000 ;
	    RECT 956.7000 1385.2500 1128.9000 1386.7500 ;
	    RECT 956.7000 1385.1000 958.5000 1385.2500 ;
	    RECT 1127.1000 1385.1000 1128.9000 1385.2500 ;
	    RECT 1307.1000 1386.7500 1308.9000 1386.9000 ;
	    RECT 1314.3000 1386.7500 1316.1000 1386.9000 ;
	    RECT 1307.1000 1385.2500 1316.1000 1386.7500 ;
	    RECT 1307.1000 1385.1000 1308.9000 1385.2500 ;
	    RECT 1314.3000 1385.1000 1316.1000 1385.2500 ;
	    RECT 23.1000 1380.7500 24.9000 1380.9000 ;
	    RECT 126.3000 1380.7500 128.1000 1380.9000 ;
	    RECT 188.7000 1380.7500 190.5000 1380.9000 ;
	    RECT 23.1000 1379.2500 190.5000 1380.7500 ;
	    RECT 23.1000 1379.1000 24.9000 1379.2500 ;
	    RECT 126.3000 1379.1000 128.1000 1379.2500 ;
	    RECT 188.7000 1379.1000 190.5000 1379.2500 ;
	    RECT 260.7000 1380.7500 262.5000 1380.9000 ;
	    RECT 368.7000 1380.7500 370.5000 1380.9000 ;
	    RECT 260.7000 1379.2500 370.5000 1380.7500 ;
	    RECT 260.7000 1379.1000 262.5000 1379.2500 ;
	    RECT 368.7000 1379.1000 370.5000 1379.2500 ;
	    RECT 375.9000 1380.7500 377.7000 1380.9000 ;
	    RECT 397.5000 1380.7500 399.3000 1380.9000 ;
	    RECT 375.9000 1379.2500 399.3000 1380.7500 ;
	    RECT 375.9000 1379.1000 377.7000 1379.2500 ;
	    RECT 397.5000 1379.1000 399.3000 1379.2500 ;
	    RECT 651.9000 1380.7500 653.7000 1380.9000 ;
	    RECT 656.7000 1380.7500 658.5000 1380.9000 ;
	    RECT 651.9000 1379.2500 658.5000 1380.7500 ;
	    RECT 651.9000 1379.1000 653.7000 1379.2500 ;
	    RECT 656.7000 1379.1000 658.5000 1379.2500 ;
	    RECT 687.9000 1380.7500 689.7000 1380.9000 ;
	    RECT 887.1000 1380.7500 888.9000 1380.9000 ;
	    RECT 687.9000 1379.2500 888.9000 1380.7500 ;
	    RECT 687.9000 1379.1000 689.7000 1379.2500 ;
	    RECT 887.1000 1379.1000 888.9000 1379.2500 ;
	    RECT 918.3000 1380.7500 920.1000 1380.9000 ;
	    RECT 923.1000 1380.7500 924.9000 1380.9000 ;
	    RECT 918.3000 1379.2500 924.9000 1380.7500 ;
	    RECT 918.3000 1379.1000 920.1000 1379.2500 ;
	    RECT 923.1000 1379.1000 924.9000 1379.2500 ;
	    RECT 968.7000 1380.7500 970.5000 1380.9000 ;
	    RECT 978.3000 1380.7500 980.1000 1380.9000 ;
	    RECT 983.1000 1380.7500 984.9000 1380.9000 ;
	    RECT 968.7000 1379.2500 984.9000 1380.7500 ;
	    RECT 968.7000 1379.1000 970.5000 1379.2500 ;
	    RECT 978.3000 1379.1000 980.1000 1379.2500 ;
	    RECT 983.1000 1379.1000 984.9000 1379.2500 ;
	    RECT 1263.9000 1380.7500 1265.7001 1380.9000 ;
	    RECT 1299.9000 1380.7500 1301.7001 1380.9000 ;
	    RECT 1263.9000 1379.2500 1301.7001 1380.7500 ;
	    RECT 1263.9000 1379.1000 1265.7001 1379.2500 ;
	    RECT 1299.9000 1379.1000 1301.7001 1379.2500 ;
	    RECT 1477.5000 1380.7500 1479.3000 1380.9000 ;
	    RECT 1530.3000 1380.7500 1532.1000 1380.9000 ;
	    RECT 1477.5000 1379.2500 1532.1000 1380.7500 ;
	    RECT 1477.5000 1379.1000 1479.3000 1379.2500 ;
	    RECT 1530.3000 1379.1000 1532.1000 1379.2500 ;
	    RECT 75.9000 1374.7500 77.7000 1374.9000 ;
	    RECT 171.9000 1374.7500 173.7000 1374.9000 ;
	    RECT 217.5000 1374.7500 219.3000 1374.9000 ;
	    RECT 75.9000 1373.2500 219.3000 1374.7500 ;
	    RECT 75.9000 1373.1000 77.7000 1373.2500 ;
	    RECT 171.9000 1373.1000 173.7000 1373.2500 ;
	    RECT 217.5000 1373.1000 219.3000 1373.2500 ;
	    RECT 431.1000 1374.7500 432.9000 1374.9000 ;
	    RECT 445.5000 1374.7500 447.3000 1374.9000 ;
	    RECT 431.1000 1373.2500 447.3000 1374.7500 ;
	    RECT 431.1000 1373.1000 432.9000 1373.2500 ;
	    RECT 445.5000 1373.1000 447.3000 1373.2500 ;
	    RECT 747.9000 1374.7500 749.7000 1374.9000 ;
	    RECT 920.7000 1374.7500 922.5000 1374.9000 ;
	    RECT 747.9000 1373.2500 922.5000 1374.7500 ;
	    RECT 747.9000 1373.1000 749.7000 1373.2500 ;
	    RECT 920.7000 1373.1000 922.5000 1373.2500 ;
	    RECT 1295.1000 1374.7500 1296.9000 1374.9000 ;
	    RECT 1311.9000 1374.7500 1313.7001 1374.9000 ;
	    RECT 1295.1000 1373.2500 1313.7001 1374.7500 ;
	    RECT 1295.1000 1373.1000 1296.9000 1373.2500 ;
	    RECT 1311.9000 1373.1000 1313.7001 1373.2500 ;
	    RECT 1515.9000 1374.7500 1517.7001 1374.9000 ;
	    RECT 1549.5000 1374.7500 1551.3000 1374.9000 ;
	    RECT 1515.9000 1373.2500 1551.3000 1374.7500 ;
	    RECT 1515.9000 1373.1000 1517.7001 1373.2500 ;
	    RECT 1549.5000 1373.1000 1551.3000 1373.2500 ;
	    RECT 457.5000 1368.7500 459.3000 1368.9000 ;
	    RECT 493.5000 1368.7500 495.3000 1368.9000 ;
	    RECT 457.5000 1367.2500 495.3000 1368.7500 ;
	    RECT 457.5000 1367.1000 459.3000 1367.2500 ;
	    RECT 493.5000 1367.1000 495.3000 1367.2500 ;
	    RECT 507.9000 1368.7500 509.7000 1368.9000 ;
	    RECT 613.5000 1368.7500 615.3000 1368.9000 ;
	    RECT 623.1000 1368.7500 624.9000 1368.9000 ;
	    RECT 507.9000 1367.2500 624.9000 1368.7500 ;
	    RECT 507.9000 1367.1000 509.7000 1367.2500 ;
	    RECT 613.5000 1367.1000 615.3000 1367.2500 ;
	    RECT 623.1000 1367.1000 624.9000 1367.2500 ;
	    RECT 637.5000 1368.7500 639.3000 1368.9000 ;
	    RECT 1016.7000 1368.7500 1018.5000 1368.9000 ;
	    RECT 637.5000 1367.2500 1018.5000 1368.7500 ;
	    RECT 637.5000 1367.1000 639.3000 1367.2500 ;
	    RECT 1016.7000 1367.1000 1018.5000 1367.2500 ;
	    RECT 1095.9000 1368.7500 1097.7001 1368.9000 ;
	    RECT 1124.7001 1368.7500 1126.5000 1368.9000 ;
	    RECT 1095.9000 1367.2500 1126.5000 1368.7500 ;
	    RECT 1095.9000 1367.1000 1097.7001 1367.2500 ;
	    RECT 1124.7001 1367.1000 1126.5000 1367.2500 ;
	    RECT 1302.3000 1368.7500 1304.1000 1368.9000 ;
	    RECT 1328.7001 1368.7500 1330.5000 1368.9000 ;
	    RECT 1302.3000 1367.2500 1330.5000 1368.7500 ;
	    RECT 1302.3000 1367.1000 1304.1000 1367.2500 ;
	    RECT 1328.7001 1367.1000 1330.5000 1367.2500 ;
	    RECT 1484.7001 1368.7500 1486.5000 1368.9000 ;
	    RECT 1494.3000 1368.7500 1496.1000 1368.9000 ;
	    RECT 1520.7001 1368.7500 1522.5000 1368.9000 ;
	    RECT 1484.7001 1367.2500 1522.5000 1368.7500 ;
	    RECT 1484.7001 1367.1000 1486.5000 1367.2500 ;
	    RECT 1494.3000 1367.1000 1496.1000 1367.2500 ;
	    RECT 1520.7001 1367.1000 1522.5000 1367.2500 ;
	    RECT 135.9000 1362.7500 137.7000 1362.9000 ;
	    RECT 167.1000 1362.7500 168.9000 1362.9000 ;
	    RECT 135.9000 1361.2500 168.9000 1362.7500 ;
	    RECT 135.9000 1361.1000 137.7000 1361.2500 ;
	    RECT 167.1000 1361.1000 168.9000 1361.2500 ;
	    RECT 241.5000 1362.7500 243.3000 1362.9000 ;
	    RECT 359.1000 1362.7500 360.9000 1362.9000 ;
	    RECT 241.5000 1361.2500 360.9000 1362.7500 ;
	    RECT 241.5000 1361.1000 243.3000 1361.2500 ;
	    RECT 359.1000 1361.1000 360.9000 1361.2500 ;
	    RECT 479.1000 1362.7500 480.9000 1362.9000 ;
	    RECT 495.9000 1362.7500 497.7000 1362.9000 ;
	    RECT 479.1000 1361.2500 497.7000 1362.7500 ;
	    RECT 479.1000 1361.1000 480.9000 1361.2500 ;
	    RECT 495.9000 1361.1000 497.7000 1361.2500 ;
	    RECT 668.7000 1362.7500 670.5000 1362.9000 ;
	    RECT 695.1000 1362.7500 696.9000 1362.9000 ;
	    RECT 668.7000 1361.2500 696.9000 1362.7500 ;
	    RECT 668.7000 1361.1000 670.5000 1361.2500 ;
	    RECT 695.1000 1361.1000 696.9000 1361.2500 ;
	    RECT 714.3000 1362.7500 716.1000 1362.9000 ;
	    RECT 750.3000 1362.7500 752.1000 1362.9000 ;
	    RECT 714.3000 1361.2500 752.1000 1362.7500 ;
	    RECT 714.3000 1361.1000 716.1000 1361.2500 ;
	    RECT 750.3000 1361.1000 752.1000 1361.2500 ;
	    RECT 911.1000 1362.7500 912.9000 1362.9000 ;
	    RECT 925.5000 1362.7500 927.3000 1362.9000 ;
	    RECT 911.1000 1361.2500 927.3000 1362.7500 ;
	    RECT 911.1000 1361.1000 912.9000 1361.2500 ;
	    RECT 925.5000 1361.1000 927.3000 1361.2500 ;
	    RECT 1016.7000 1362.7500 1018.5000 1362.9000 ;
	    RECT 1295.1000 1362.7500 1296.9000 1362.9000 ;
	    RECT 1302.3000 1362.7500 1304.1000 1362.9000 ;
	    RECT 1016.7000 1361.2500 1304.1000 1362.7500 ;
	    RECT 1016.7000 1361.1000 1018.5000 1361.2500 ;
	    RECT 1295.1000 1361.1000 1296.9000 1361.2500 ;
	    RECT 1302.3000 1361.1000 1304.1000 1361.2500 ;
	    RECT 1311.9000 1362.7500 1313.7001 1362.9000 ;
	    RECT 1347.9000 1362.7500 1349.7001 1362.9000 ;
	    RECT 1311.9000 1361.2500 1349.7001 1362.7500 ;
	    RECT 1311.9000 1361.1000 1313.7001 1361.2500 ;
	    RECT 1347.9000 1361.1000 1349.7001 1361.2500 ;
	    RECT 1515.9000 1362.7500 1517.7001 1362.9000 ;
	    RECT 1523.1000 1362.7500 1524.9000 1362.9000 ;
	    RECT 1515.9000 1361.2500 1524.9000 1362.7500 ;
	    RECT 1515.9000 1361.1000 1517.7001 1361.2500 ;
	    RECT 1523.1000 1361.1000 1524.9000 1361.2500 ;
	    RECT 104.7000 1356.7500 106.5000 1356.9000 ;
	    RECT 145.5000 1356.7500 147.3000 1356.9000 ;
	    RECT 104.7000 1355.2500 147.3000 1356.7500 ;
	    RECT 104.7000 1355.1000 106.5000 1355.2500 ;
	    RECT 145.5000 1355.1000 147.3000 1355.2500 ;
	    RECT 416.7000 1356.7500 418.5000 1356.9000 ;
	    RECT 507.9000 1356.7500 509.7000 1356.9000 ;
	    RECT 416.7000 1355.2500 509.7000 1356.7500 ;
	    RECT 416.7000 1355.1000 418.5000 1355.2500 ;
	    RECT 507.9000 1355.1000 509.7000 1355.2500 ;
	    RECT 649.5000 1356.7500 651.3000 1356.9000 ;
	    RECT 719.1000 1356.7500 720.9000 1356.9000 ;
	    RECT 649.5000 1355.2500 720.9000 1356.7500 ;
	    RECT 649.5000 1355.1000 651.3000 1355.2500 ;
	    RECT 719.1000 1355.1000 720.9000 1355.2500 ;
	    RECT 767.1000 1356.7500 768.9000 1356.9000 ;
	    RECT 877.5000 1356.7500 879.3000 1356.9000 ;
	    RECT 767.1000 1355.2500 879.3000 1356.7500 ;
	    RECT 767.1000 1355.1000 768.9000 1355.2500 ;
	    RECT 877.5000 1355.1000 879.3000 1355.2500 ;
	    RECT 973.5000 1356.7500 975.3000 1356.9000 ;
	    RECT 1124.7001 1356.7500 1126.5000 1356.9000 ;
	    RECT 973.5000 1355.2500 1126.5000 1356.7500 ;
	    RECT 973.5000 1355.1000 975.3000 1355.2500 ;
	    RECT 1124.7001 1355.1000 1126.5000 1355.2500 ;
	    RECT 1134.3000 1356.7500 1136.1000 1356.9000 ;
	    RECT 1280.7001 1356.7500 1282.5000 1356.9000 ;
	    RECT 1134.3000 1355.2500 1282.5000 1356.7500 ;
	    RECT 1134.3000 1355.1000 1136.1000 1355.2500 ;
	    RECT 1280.7001 1355.1000 1282.5000 1355.2500 ;
	    RECT 1292.7001 1356.7500 1294.5000 1356.9000 ;
	    RECT 1343.1000 1356.7500 1344.9000 1356.9000 ;
	    RECT 1292.7001 1355.2500 1344.9000 1356.7500 ;
	    RECT 1292.7001 1355.1000 1294.5000 1355.2500 ;
	    RECT 1343.1000 1355.1000 1344.9000 1355.2500 ;
	    RECT 1499.1000 1356.7500 1500.9000 1356.9000 ;
	    RECT 1542.3000 1356.7500 1544.1000 1356.9000 ;
	    RECT 1499.1000 1355.2500 1544.1000 1356.7500 ;
	    RECT 1499.1000 1355.1000 1500.9000 1355.2500 ;
	    RECT 1542.3000 1355.1000 1544.1000 1355.2500 ;
	    RECT 488.7000 1350.7500 490.5000 1350.9000 ;
	    RECT 541.5000 1350.7500 543.3000 1350.9000 ;
	    RECT 488.7000 1349.2500 543.3000 1350.7500 ;
	    RECT 488.7000 1349.1000 490.5000 1349.2500 ;
	    RECT 541.5000 1349.1000 543.3000 1349.2500 ;
	    RECT 939.9000 1350.7500 941.7000 1350.9000 ;
	    RECT 985.5000 1350.7500 987.3000 1350.9000 ;
	    RECT 939.9000 1349.2500 987.3000 1350.7500 ;
	    RECT 939.9000 1349.1000 941.7000 1349.2500 ;
	    RECT 985.5000 1349.1000 987.3000 1349.2500 ;
	    RECT 1309.5000 1350.7500 1311.3000 1350.9000 ;
	    RECT 1340.7001 1350.7500 1342.5000 1350.9000 ;
	    RECT 1309.5000 1349.2500 1342.5000 1350.7500 ;
	    RECT 1309.5000 1349.1000 1311.3000 1349.2500 ;
	    RECT 1340.7001 1349.1000 1342.5000 1349.2500 ;
	    RECT 1494.3000 1350.7500 1496.1000 1350.9000 ;
	    RECT 1499.1000 1350.7500 1500.9000 1350.9000 ;
	    RECT 1494.3000 1349.2500 1500.9000 1350.7500 ;
	    RECT 1494.3000 1349.1000 1496.1000 1349.2500 ;
	    RECT 1499.1000 1349.1000 1500.9000 1349.2500 ;
	    RECT 663.9000 1344.7500 665.7000 1344.9000 ;
	    RECT 719.1000 1344.7500 720.9000 1344.9000 ;
	    RECT 663.9000 1343.2500 720.9000 1344.7500 ;
	    RECT 663.9000 1343.1000 665.7000 1343.2500 ;
	    RECT 719.1000 1343.1000 720.9000 1343.2500 ;
	    RECT 872.7000 1344.7500 874.5000 1344.9000 ;
	    RECT 923.1000 1344.7500 924.9000 1344.9000 ;
	    RECT 872.7000 1343.2500 924.9000 1344.7500 ;
	    RECT 872.7000 1343.1000 874.5000 1343.2500 ;
	    RECT 923.1000 1343.1000 924.9000 1343.2500 ;
	    RECT 927.9000 1344.7500 929.7000 1344.9000 ;
	    RECT 949.5000 1344.7500 951.3000 1344.9000 ;
	    RECT 927.9000 1343.2500 951.3000 1344.7500 ;
	    RECT 927.9000 1343.1000 929.7000 1343.2500 ;
	    RECT 949.5000 1343.1000 951.3000 1343.2500 ;
	    RECT 1040.7001 1344.7500 1042.5000 1344.9000 ;
	    RECT 1170.3000 1344.7500 1172.1000 1344.9000 ;
	    RECT 1040.7001 1343.2500 1172.1000 1344.7500 ;
	    RECT 1040.7001 1343.1000 1042.5000 1343.2500 ;
	    RECT 1170.3000 1343.1000 1172.1000 1343.2500 ;
	    RECT 1347.9000 1344.7500 1349.7001 1344.9000 ;
	    RECT 1398.3000 1344.7500 1400.1000 1344.9000 ;
	    RECT 1347.9000 1343.2500 1400.1000 1344.7500 ;
	    RECT 1347.9000 1343.1000 1349.7001 1343.2500 ;
	    RECT 1398.3000 1343.1000 1400.1000 1343.2500 ;
	    RECT 366.3000 1338.7500 368.1000 1338.9000 ;
	    RECT 551.1000 1338.7500 552.9000 1338.9000 ;
	    RECT 366.3000 1337.2500 552.9000 1338.7500 ;
	    RECT 366.3000 1337.1000 368.1000 1337.2500 ;
	    RECT 551.1000 1337.1000 552.9000 1337.2500 ;
	    RECT 678.3000 1338.7500 680.1000 1338.9000 ;
	    RECT 704.7000 1338.7500 706.5000 1338.9000 ;
	    RECT 678.3000 1337.2500 706.5000 1338.7500 ;
	    RECT 678.3000 1337.1000 680.1000 1337.2500 ;
	    RECT 704.7000 1337.1000 706.5000 1337.2500 ;
	    RECT 911.1000 1338.7500 912.9000 1338.9000 ;
	    RECT 927.9000 1338.7500 929.7000 1338.9000 ;
	    RECT 911.1000 1337.2500 929.7000 1338.7500 ;
	    RECT 911.1000 1337.1000 912.9000 1337.2500 ;
	    RECT 927.9000 1337.1000 929.7000 1337.2500 ;
	    RECT 937.5000 1338.7500 939.3000 1338.9000 ;
	    RECT 1223.1000 1338.7500 1224.9000 1338.9000 ;
	    RECT 937.5000 1337.2500 1224.9000 1338.7500 ;
	    RECT 937.5000 1337.1000 939.3000 1337.2500 ;
	    RECT 1223.1000 1337.1000 1224.9000 1337.2500 ;
	    RECT 1295.1000 1338.7500 1296.9000 1338.9000 ;
	    RECT 1345.5000 1338.7500 1347.3000 1338.9000 ;
	    RECT 1295.1000 1337.2500 1347.3000 1338.7500 ;
	    RECT 1295.1000 1337.1000 1296.9000 1337.2500 ;
	    RECT 1345.5000 1337.1000 1347.3000 1337.2500 ;
	    RECT 1470.3000 1338.7500 1472.1000 1338.9000 ;
	    RECT 1484.7001 1338.7500 1486.5000 1338.9000 ;
	    RECT 1470.3000 1337.2500 1486.5000 1338.7500 ;
	    RECT 1470.3000 1337.1000 1472.1000 1337.2500 ;
	    RECT 1484.7001 1337.1000 1486.5000 1337.2500 ;
	    RECT 1539.9000 1338.7500 1541.7001 1338.9000 ;
	    RECT 1547.1000 1338.7500 1548.9000 1338.9000 ;
	    RECT 1539.9000 1337.2500 1548.9000 1338.7500 ;
	    RECT 1539.9000 1337.1000 1541.7001 1337.2500 ;
	    RECT 1547.1000 1337.1000 1548.9000 1337.2500 ;
	    RECT 887.1000 1332.7500 888.9000 1332.9000 ;
	    RECT 903.9000 1332.7500 905.7000 1332.9000 ;
	    RECT 975.9000 1332.7500 977.7000 1332.9000 ;
	    RECT 887.1000 1331.2500 977.7000 1332.7500 ;
	    RECT 887.1000 1331.1000 888.9000 1331.2500 ;
	    RECT 903.9000 1331.1000 905.7000 1331.2500 ;
	    RECT 975.9000 1331.1000 977.7000 1331.2500 ;
	    RECT 1170.3000 1332.7500 1172.1000 1332.9000 ;
	    RECT 1213.5000 1332.7500 1215.3000 1332.9000 ;
	    RECT 1170.3000 1331.2500 1215.3000 1332.7500 ;
	    RECT 1170.3000 1331.1000 1172.1000 1331.2500 ;
	    RECT 1213.5000 1331.1000 1215.3000 1331.2500 ;
	    RECT 1446.3000 1332.7500 1448.1000 1332.9000 ;
	    RECT 1566.3000 1332.7500 1568.1000 1332.9000 ;
	    RECT 1446.3000 1331.2500 1568.1000 1332.7500 ;
	    RECT 1446.3000 1331.1000 1448.1000 1331.2500 ;
	    RECT 1566.3000 1331.1000 1568.1000 1331.2500 ;
	    RECT 78.3000 1326.7500 80.1000 1326.9000 ;
	    RECT 152.7000 1326.7500 154.5000 1326.9000 ;
	    RECT 78.3000 1325.2500 154.5000 1326.7500 ;
	    RECT 78.3000 1325.1000 80.1000 1325.2500 ;
	    RECT 152.7000 1325.1000 154.5000 1325.2500 ;
	    RECT 169.5000 1326.7500 171.3000 1326.9000 ;
	    RECT 359.1000 1326.7500 360.9000 1326.9000 ;
	    RECT 169.5000 1325.2500 360.9000 1326.7500 ;
	    RECT 169.5000 1325.1000 171.3000 1325.2500 ;
	    RECT 359.1000 1325.1000 360.9000 1325.2500 ;
	    RECT 644.7000 1326.7500 646.5000 1326.9000 ;
	    RECT 663.9000 1326.7500 665.7000 1326.9000 ;
	    RECT 644.7000 1325.2500 665.7000 1326.7500 ;
	    RECT 644.7000 1325.1000 646.5000 1325.2500 ;
	    RECT 663.9000 1325.1000 665.7000 1325.2500 ;
	    RECT 827.1000 1326.7500 828.9000 1326.9000 ;
	    RECT 899.1000 1326.7500 900.9000 1326.9000 ;
	    RECT 942.3000 1326.7500 944.1000 1326.9000 ;
	    RECT 827.1000 1325.2500 944.1000 1326.7500 ;
	    RECT 827.1000 1325.1000 828.9000 1325.2500 ;
	    RECT 899.1000 1325.1000 900.9000 1325.2500 ;
	    RECT 942.3000 1325.1000 944.1000 1325.2500 ;
	    RECT 947.1000 1326.7500 948.9000 1326.9000 ;
	    RECT 1251.9000 1326.7500 1253.7001 1326.9000 ;
	    RECT 947.1000 1325.2500 1253.7001 1326.7500 ;
	    RECT 947.1000 1325.1000 948.9000 1325.2500 ;
	    RECT 1251.9000 1325.1000 1253.7001 1325.2500 ;
	    RECT 1302.3000 1326.7500 1304.1000 1326.9000 ;
	    RECT 1518.3000 1326.7500 1520.1000 1326.9000 ;
	    RECT 1302.3000 1325.2500 1520.1000 1326.7500 ;
	    RECT 1302.3000 1325.1000 1304.1000 1325.2500 ;
	    RECT 1518.3000 1325.1000 1520.1000 1325.2500 ;
	    RECT 1542.3000 1326.7500 1544.1000 1326.9000 ;
	    RECT 1554.3000 1326.7500 1556.1000 1326.9000 ;
	    RECT 1542.3000 1325.2500 1556.1000 1326.7500 ;
	    RECT 1542.3000 1325.1000 1544.1000 1325.2500 ;
	    RECT 1554.3000 1325.1000 1556.1000 1325.2500 ;
	    RECT 275.1000 1320.7500 276.9000 1320.9000 ;
	    RECT 351.9000 1320.7500 353.7000 1320.9000 ;
	    RECT 275.1000 1319.2500 353.7000 1320.7500 ;
	    RECT 275.1000 1319.1000 276.9000 1319.2500 ;
	    RECT 351.9000 1319.1000 353.7000 1319.2500 ;
	    RECT 359.1000 1320.7500 360.9000 1320.9000 ;
	    RECT 459.9000 1320.7500 461.7000 1320.9000 ;
	    RECT 359.1000 1319.2500 461.7000 1320.7500 ;
	    RECT 359.1000 1319.1000 360.9000 1319.2500 ;
	    RECT 459.9000 1319.1000 461.7000 1319.2500 ;
	    RECT 608.7000 1320.7500 610.5000 1320.9000 ;
	    RECT 649.5000 1320.7500 651.3000 1320.9000 ;
	    RECT 608.7000 1319.2500 651.3000 1320.7500 ;
	    RECT 608.7000 1319.1000 610.5000 1319.2500 ;
	    RECT 649.5000 1319.1000 651.3000 1319.2500 ;
	    RECT 687.9000 1320.7500 689.7000 1320.9000 ;
	    RECT 743.1000 1320.7500 744.9000 1320.9000 ;
	    RECT 687.9000 1319.2500 744.9000 1320.7500 ;
	    RECT 687.9000 1319.1000 689.7000 1319.2500 ;
	    RECT 743.1000 1319.1000 744.9000 1319.2500 ;
	    RECT 942.3000 1320.7500 944.1000 1320.9000 ;
	    RECT 951.9000 1320.7500 953.7000 1320.9000 ;
	    RECT 942.3000 1319.2500 953.7000 1320.7500 ;
	    RECT 942.3000 1319.1000 944.1000 1319.2500 ;
	    RECT 951.9000 1319.1000 953.7000 1319.2500 ;
	    RECT 1443.9000 1320.7500 1445.7001 1320.9000 ;
	    RECT 1453.5000 1320.7500 1455.3000 1320.9000 ;
	    RECT 1470.3000 1320.7500 1472.1000 1320.9000 ;
	    RECT 1443.9000 1319.2500 1472.1000 1320.7500 ;
	    RECT 1443.9000 1319.1000 1445.7001 1319.2500 ;
	    RECT 1453.5000 1319.1000 1455.3000 1319.2500 ;
	    RECT 1470.3000 1319.1000 1472.1000 1319.2500 ;
	    RECT 152.7000 1314.7500 154.5000 1314.9000 ;
	    RECT 275.1000 1314.7500 276.9000 1314.9000 ;
	    RECT 152.7000 1313.2500 276.9000 1314.7500 ;
	    RECT 152.7000 1313.1000 154.5000 1313.2500 ;
	    RECT 275.1000 1313.1000 276.9000 1313.2500 ;
	    RECT 373.5000 1314.7500 375.3000 1314.9000 ;
	    RECT 445.5000 1314.7500 447.3000 1314.9000 ;
	    RECT 491.1000 1314.7500 492.9000 1314.9000 ;
	    RECT 536.7000 1314.7500 538.5000 1314.9000 ;
	    RECT 373.5000 1313.2500 538.5000 1314.7500 ;
	    RECT 373.5000 1313.1000 375.3000 1313.2500 ;
	    RECT 445.5000 1313.1000 447.3000 1313.2500 ;
	    RECT 491.1000 1313.1000 492.9000 1313.2500 ;
	    RECT 536.7000 1313.1000 538.5000 1313.2500 ;
	    RECT 649.5000 1314.7500 651.3000 1314.9000 ;
	    RECT 663.9000 1314.7500 665.7000 1314.9000 ;
	    RECT 649.5000 1313.2500 665.7000 1314.7500 ;
	    RECT 649.5000 1313.1000 651.3000 1313.2500 ;
	    RECT 663.9000 1313.1000 665.7000 1313.2500 ;
	    RECT 731.1000 1314.7500 732.9000 1314.9000 ;
	    RECT 755.1000 1314.7500 756.9000 1314.9000 ;
	    RECT 764.7000 1314.7500 766.5000 1314.9000 ;
	    RECT 731.1000 1313.2500 766.5000 1314.7500 ;
	    RECT 731.1000 1313.1000 732.9000 1313.2500 ;
	    RECT 755.1000 1313.1000 756.9000 1313.2500 ;
	    RECT 764.7000 1313.1000 766.5000 1313.2500 ;
	    RECT 829.5000 1314.7500 831.3000 1314.9000 ;
	    RECT 997.5000 1314.7500 999.3000 1314.9000 ;
	    RECT 829.5000 1313.2500 999.3000 1314.7500 ;
	    RECT 829.5000 1313.1000 831.3000 1313.2500 ;
	    RECT 997.5000 1313.1000 999.3000 1313.2500 ;
	    RECT 1225.5000 1314.7500 1227.3000 1314.9000 ;
	    RECT 1232.7001 1314.7500 1234.5000 1314.9000 ;
	    RECT 1225.5000 1313.2500 1234.5000 1314.7500 ;
	    RECT 1225.5000 1313.1000 1227.3000 1313.2500 ;
	    RECT 1232.7001 1313.1000 1234.5000 1313.2500 ;
	    RECT 83.1000 1308.7500 84.9000 1308.9000 ;
	    RECT 181.5000 1308.7500 183.3000 1308.9000 ;
	    RECT 83.1000 1307.2500 183.3000 1308.7500 ;
	    RECT 83.1000 1307.1000 84.9000 1307.2500 ;
	    RECT 181.5000 1307.1000 183.3000 1307.2500 ;
	    RECT 195.9000 1308.7500 197.7000 1308.9000 ;
	    RECT 231.9000 1308.7500 233.7000 1308.9000 ;
	    RECT 195.9000 1307.2500 233.7000 1308.7500 ;
	    RECT 195.9000 1307.1000 197.7000 1307.2500 ;
	    RECT 231.9000 1307.1000 233.7000 1307.2500 ;
	    RECT 287.1000 1308.7500 288.9000 1308.9000 ;
	    RECT 471.9000 1308.7500 473.7000 1308.9000 ;
	    RECT 287.1000 1307.2500 473.7000 1308.7500 ;
	    RECT 287.1000 1307.1000 288.9000 1307.2500 ;
	    RECT 471.9000 1307.1000 473.7000 1307.2500 ;
	    RECT 812.7000 1308.7500 814.5000 1308.9000 ;
	    RECT 819.9000 1308.7500 821.7000 1308.9000 ;
	    RECT 812.7000 1307.2500 821.7000 1308.7500 ;
	    RECT 812.7000 1307.1000 814.5000 1307.2500 ;
	    RECT 819.9000 1307.1000 821.7000 1307.2500 ;
	    RECT 831.9000 1308.7500 833.7000 1308.9000 ;
	    RECT 860.7000 1308.7500 862.5000 1308.9000 ;
	    RECT 831.9000 1307.2500 862.5000 1308.7500 ;
	    RECT 831.9000 1307.1000 833.7000 1307.2500 ;
	    RECT 860.7000 1307.1000 862.5000 1307.2500 ;
	    RECT 951.9000 1308.7500 953.7000 1308.9000 ;
	    RECT 983.1000 1308.7500 984.9000 1308.9000 ;
	    RECT 951.9000 1307.2500 984.9000 1308.7500 ;
	    RECT 951.9000 1307.1000 953.7000 1307.2500 ;
	    RECT 983.1000 1307.1000 984.9000 1307.2500 ;
	    RECT 1191.9000 1308.7500 1193.7001 1308.9000 ;
	    RECT 1211.1000 1308.7500 1212.9000 1308.9000 ;
	    RECT 1191.9000 1307.2500 1212.9000 1308.7500 ;
	    RECT 1191.9000 1307.1000 1193.7001 1307.2500 ;
	    RECT 1211.1000 1307.1000 1212.9000 1307.2500 ;
	    RECT 1278.3000 1308.7500 1280.1000 1308.9000 ;
	    RECT 1285.5000 1308.7500 1287.3000 1308.9000 ;
	    RECT 1278.3000 1307.2500 1287.3000 1308.7500 ;
	    RECT 1278.3000 1307.1000 1280.1000 1307.2500 ;
	    RECT 1285.5000 1307.1000 1287.3000 1307.2500 ;
	    RECT 1448.7001 1308.7500 1450.5000 1308.9000 ;
	    RECT 1501.5000 1308.7500 1503.3000 1308.9000 ;
	    RECT 1448.7001 1307.2500 1503.3000 1308.7500 ;
	    RECT 1448.7001 1307.1000 1450.5000 1307.2500 ;
	    RECT 1501.5000 1307.1000 1503.3000 1307.2500 ;
	    RECT 18.3000 1302.7500 20.1000 1302.9000 ;
	    RECT 80.7000 1302.7500 82.5000 1302.9000 ;
	    RECT 107.1000 1302.7500 108.9000 1302.9000 ;
	    RECT 18.3000 1301.2500 108.9000 1302.7500 ;
	    RECT 18.3000 1301.1000 20.1000 1301.2500 ;
	    RECT 80.7000 1301.1000 82.5000 1301.2500 ;
	    RECT 107.1000 1301.1000 108.9000 1301.2500 ;
	    RECT 229.5000 1302.7500 231.3000 1302.9000 ;
	    RECT 236.7000 1302.7500 238.5000 1302.9000 ;
	    RECT 229.5000 1301.2500 238.5000 1302.7500 ;
	    RECT 229.5000 1301.1000 231.3000 1301.2500 ;
	    RECT 236.7000 1301.1000 238.5000 1301.2500 ;
	    RECT 272.7000 1302.7500 274.5000 1302.9000 ;
	    RECT 279.9000 1302.7500 281.7000 1302.9000 ;
	    RECT 272.7000 1301.2500 281.7000 1302.7500 ;
	    RECT 272.7000 1301.1000 274.5000 1301.2500 ;
	    RECT 279.9000 1301.1000 281.7000 1301.2500 ;
	    RECT 404.7000 1302.7500 406.5000 1302.9000 ;
	    RECT 450.3000 1302.7500 452.1000 1302.9000 ;
	    RECT 404.7000 1301.2500 452.1000 1302.7500 ;
	    RECT 404.7000 1301.1000 406.5000 1301.2500 ;
	    RECT 450.3000 1301.1000 452.1000 1301.2500 ;
	    RECT 1019.1000 1302.7500 1020.9000 1302.9000 ;
	    RECT 1023.9000 1302.7500 1025.7001 1302.9000 ;
	    RECT 1019.1000 1301.2500 1025.7001 1302.7500 ;
	    RECT 1019.1000 1301.1000 1020.9000 1301.2500 ;
	    RECT 1023.9000 1301.1000 1025.7001 1301.2500 ;
	    RECT 1040.7001 1302.7500 1042.5000 1302.9000 ;
	    RECT 1047.9000 1302.7500 1049.7001 1302.9000 ;
	    RECT 1040.7001 1301.2500 1049.7001 1302.7500 ;
	    RECT 1040.7001 1301.1000 1042.5000 1301.2500 ;
	    RECT 1047.9000 1301.1000 1049.7001 1301.2500 ;
	    RECT 1134.3000 1302.7500 1136.1000 1302.9000 ;
	    RECT 1220.7001 1302.7500 1222.5000 1302.9000 ;
	    RECT 1134.3000 1301.2500 1222.5000 1302.7500 ;
	    RECT 1134.3000 1301.1000 1136.1000 1301.2500 ;
	    RECT 1220.7001 1301.1000 1222.5000 1301.2500 ;
	    RECT 1379.1000 1302.7500 1380.9000 1302.9000 ;
	    RECT 1475.1000 1302.7500 1476.9000 1302.9000 ;
	    RECT 1379.1000 1301.2500 1476.9000 1302.7500 ;
	    RECT 1379.1000 1301.1000 1380.9000 1301.2500 ;
	    RECT 1475.1000 1301.1000 1476.9000 1301.2500 ;
	    RECT 133.5000 1296.7500 135.3000 1296.9000 ;
	    RECT 399.9000 1296.7500 401.7000 1296.9000 ;
	    RECT 133.5000 1295.2500 401.7000 1296.7500 ;
	    RECT 133.5000 1295.1000 135.3000 1295.2500 ;
	    RECT 399.9000 1295.1000 401.7000 1295.2500 ;
	    RECT 618.3000 1296.7500 620.1000 1296.9000 ;
	    RECT 839.1000 1296.7500 840.9000 1296.9000 ;
	    RECT 618.3000 1295.2500 840.9000 1296.7500 ;
	    RECT 618.3000 1295.1000 620.1000 1295.2500 ;
	    RECT 839.1000 1295.1000 840.9000 1295.2500 ;
	    RECT 908.7000 1296.7500 910.5000 1296.9000 ;
	    RECT 959.1000 1296.7500 960.9000 1296.9000 ;
	    RECT 908.7000 1295.2500 960.9000 1296.7500 ;
	    RECT 908.7000 1295.1000 910.5000 1295.2500 ;
	    RECT 959.1000 1295.1000 960.9000 1295.2500 ;
	    RECT 1011.9000 1296.7500 1013.7000 1296.9000 ;
	    RECT 1071.9000 1296.7500 1073.7001 1296.9000 ;
	    RECT 1011.9000 1295.2500 1073.7001 1296.7500 ;
	    RECT 1011.9000 1295.1000 1013.7000 1295.2500 ;
	    RECT 1071.9000 1295.1000 1073.7001 1295.2500 ;
	    RECT 1177.5000 1296.7500 1179.3000 1296.9000 ;
	    RECT 1191.9000 1296.7500 1193.7001 1296.9000 ;
	    RECT 1177.5000 1295.2500 1193.7001 1296.7500 ;
	    RECT 1177.5000 1295.1000 1179.3000 1295.2500 ;
	    RECT 1191.9000 1295.1000 1193.7001 1295.2500 ;
	    RECT 1443.9000 1296.7500 1445.7001 1296.9000 ;
	    RECT 1484.7001 1296.7500 1486.5000 1296.9000 ;
	    RECT 1443.9000 1295.2500 1486.5000 1296.7500 ;
	    RECT 1443.9000 1295.1000 1445.7001 1295.2500 ;
	    RECT 1484.7001 1295.1000 1486.5000 1295.2500 ;
	    RECT 107.1000 1290.7500 108.9000 1290.9000 ;
	    RECT 152.7000 1290.7500 154.5000 1290.9000 ;
	    RECT 183.9000 1290.7500 185.7000 1290.9000 ;
	    RECT 239.1000 1290.7500 240.9000 1290.9000 ;
	    RECT 272.7000 1290.7500 274.5000 1290.9000 ;
	    RECT 107.1000 1289.2500 274.5000 1290.7500 ;
	    RECT 107.1000 1289.1000 108.9000 1289.2500 ;
	    RECT 152.7000 1289.1000 154.5000 1289.2500 ;
	    RECT 183.9000 1289.1000 185.7000 1289.2500 ;
	    RECT 239.1000 1289.1000 240.9000 1289.2500 ;
	    RECT 272.7000 1289.1000 274.5000 1289.2500 ;
	    RECT 282.3000 1290.7500 284.1000 1290.9000 ;
	    RECT 291.9000 1290.7500 293.7000 1290.9000 ;
	    RECT 282.3000 1289.2500 293.7000 1290.7500 ;
	    RECT 282.3000 1289.1000 284.1000 1289.2500 ;
	    RECT 291.9000 1289.1000 293.7000 1289.2500 ;
	    RECT 311.1000 1290.7500 312.9000 1290.9000 ;
	    RECT 327.9000 1290.7500 329.7000 1290.9000 ;
	    RECT 311.1000 1289.2500 329.7000 1290.7500 ;
	    RECT 311.1000 1289.1000 312.9000 1289.2500 ;
	    RECT 327.9000 1289.1000 329.7000 1289.2500 ;
	    RECT 635.1000 1290.7500 636.9000 1290.9000 ;
	    RECT 649.5000 1290.7500 651.3000 1290.9000 ;
	    RECT 635.1000 1289.2500 651.3000 1290.7500 ;
	    RECT 635.1000 1289.1000 636.9000 1289.2500 ;
	    RECT 649.5000 1289.1000 651.3000 1289.2500 ;
	    RECT 709.5000 1290.7500 711.3000 1290.9000 ;
	    RECT 757.5000 1290.7500 759.3000 1290.9000 ;
	    RECT 709.5000 1289.2500 759.3000 1290.7500 ;
	    RECT 709.5000 1289.1000 711.3000 1289.2500 ;
	    RECT 757.5000 1289.1000 759.3000 1289.2500 ;
	    RECT 959.1000 1290.7500 960.9000 1290.9000 ;
	    RECT 995.1000 1290.7500 996.9000 1290.9000 ;
	    RECT 959.1000 1289.2500 996.9000 1290.7500 ;
	    RECT 959.1000 1289.1000 960.9000 1289.2500 ;
	    RECT 995.1000 1289.1000 996.9000 1289.2500 ;
	    RECT 1215.9000 1290.7500 1217.7001 1290.9000 ;
	    RECT 1223.1000 1290.7500 1224.9000 1290.9000 ;
	    RECT 1215.9000 1289.2500 1224.9000 1290.7500 ;
	    RECT 1215.9000 1289.1000 1217.7001 1289.2500 ;
	    RECT 1223.1000 1289.1000 1224.9000 1289.2500 ;
	    RECT 167.1000 1284.7500 168.9000 1284.9000 ;
	    RECT 241.5000 1284.7500 243.3000 1284.9000 ;
	    RECT 167.1000 1283.2500 243.3000 1284.7500 ;
	    RECT 167.1000 1283.1000 168.9000 1283.2500 ;
	    RECT 241.5000 1283.1000 243.3000 1283.2500 ;
	    RECT 620.7000 1284.7500 622.5000 1284.9000 ;
	    RECT 632.7000 1284.7500 634.5000 1284.9000 ;
	    RECT 642.3000 1284.7500 644.1000 1284.9000 ;
	    RECT 620.7000 1283.2500 644.1000 1284.7500 ;
	    RECT 620.7000 1283.1000 622.5000 1283.2500 ;
	    RECT 632.7000 1283.1000 634.5000 1283.2500 ;
	    RECT 642.3000 1283.1000 644.1000 1283.2500 ;
	    RECT 687.9000 1284.7500 689.7000 1284.9000 ;
	    RECT 699.9000 1284.7500 701.7000 1284.9000 ;
	    RECT 687.9000 1283.2500 701.7000 1284.7500 ;
	    RECT 687.9000 1283.1000 689.7000 1283.2500 ;
	    RECT 699.9000 1283.1000 701.7000 1283.2500 ;
	    RECT 884.7000 1284.7500 886.5000 1284.9000 ;
	    RECT 983.1000 1284.7500 984.9000 1284.9000 ;
	    RECT 884.7000 1283.2500 984.9000 1284.7500 ;
	    RECT 884.7000 1283.1000 886.5000 1283.2500 ;
	    RECT 983.1000 1283.1000 984.9000 1283.2500 ;
	    RECT 987.9000 1284.7500 989.7000 1284.9000 ;
	    RECT 1011.9000 1284.7500 1013.7000 1284.9000 ;
	    RECT 987.9000 1283.2500 1013.7000 1284.7500 ;
	    RECT 987.9000 1283.1000 989.7000 1283.2500 ;
	    RECT 1011.9000 1283.1000 1013.7000 1283.2500 ;
	    RECT 1033.5000 1284.7500 1035.3000 1284.9000 ;
	    RECT 1052.7001 1284.7500 1054.5000 1284.9000 ;
	    RECT 1033.5000 1283.2500 1054.5000 1284.7500 ;
	    RECT 1033.5000 1283.1000 1035.3000 1283.2500 ;
	    RECT 1052.7001 1283.1000 1054.5000 1283.2500 ;
	    RECT 1206.3000 1284.7500 1208.1000 1284.9000 ;
	    RECT 1232.7001 1284.7500 1234.5000 1284.9000 ;
	    RECT 1206.3000 1283.2500 1234.5000 1284.7500 ;
	    RECT 1206.3000 1283.1000 1208.1000 1283.2500 ;
	    RECT 1232.7001 1283.1000 1234.5000 1283.2500 ;
	    RECT 27.9000 1278.7500 29.7000 1278.9000 ;
	    RECT 35.1000 1278.7500 36.9000 1278.9000 ;
	    RECT 27.9000 1277.2500 36.9000 1278.7500 ;
	    RECT 27.9000 1277.1000 29.7000 1277.2500 ;
	    RECT 35.1000 1277.1000 36.9000 1277.2500 ;
	    RECT 323.1000 1278.7500 324.9000 1278.9000 ;
	    RECT 359.1000 1278.7500 360.9000 1278.9000 ;
	    RECT 323.1000 1277.2500 360.9000 1278.7500 ;
	    RECT 323.1000 1277.1000 324.9000 1277.2500 ;
	    RECT 359.1000 1277.1000 360.9000 1277.2500 ;
	    RECT 395.1000 1278.7500 396.9000 1278.9000 ;
	    RECT 409.5000 1278.7500 411.3000 1278.9000 ;
	    RECT 395.1000 1277.2500 411.3000 1278.7500 ;
	    RECT 395.1000 1277.1000 396.9000 1277.2500 ;
	    RECT 409.5000 1277.1000 411.3000 1277.2500 ;
	    RECT 539.1000 1278.7500 540.9000 1278.9000 ;
	    RECT 558.3000 1278.7500 560.1000 1278.9000 ;
	    RECT 539.1000 1277.2500 560.1000 1278.7500 ;
	    RECT 539.1000 1277.1000 540.9000 1277.2500 ;
	    RECT 558.3000 1277.1000 560.1000 1277.2500 ;
	    RECT 565.5000 1278.7500 567.3000 1278.9000 ;
	    RECT 644.7000 1278.7500 646.5000 1278.9000 ;
	    RECT 565.5000 1277.2500 646.5000 1278.7500 ;
	    RECT 565.5000 1277.1000 567.3000 1277.2500 ;
	    RECT 644.7000 1277.1000 646.5000 1277.2500 ;
	    RECT 695.1000 1278.7500 696.9000 1278.9000 ;
	    RECT 728.7000 1278.7500 730.5000 1278.9000 ;
	    RECT 695.1000 1277.2500 730.5000 1278.7500 ;
	    RECT 695.1000 1277.1000 696.9000 1277.2500 ;
	    RECT 728.7000 1277.1000 730.5000 1277.2500 ;
	    RECT 882.3000 1278.7500 884.1000 1278.9000 ;
	    RECT 896.7000 1278.7500 898.5000 1278.9000 ;
	    RECT 882.3000 1277.2500 898.5000 1278.7500 ;
	    RECT 882.3000 1277.1000 884.1000 1277.2500 ;
	    RECT 896.7000 1277.1000 898.5000 1277.2500 ;
	    RECT 930.3000 1278.7500 932.1000 1278.9000 ;
	    RECT 937.5000 1278.7500 939.3000 1278.9000 ;
	    RECT 930.3000 1277.2500 939.3000 1278.7500 ;
	    RECT 930.3000 1277.1000 932.1000 1277.2500 ;
	    RECT 937.5000 1277.1000 939.3000 1277.2500 ;
	    RECT 975.9000 1278.7500 977.7000 1278.9000 ;
	    RECT 1177.5000 1278.7500 1179.3000 1278.9000 ;
	    RECT 1218.3000 1278.7500 1220.1000 1278.9000 ;
	    RECT 975.9000 1277.2500 1220.1000 1278.7500 ;
	    RECT 975.9000 1277.1000 977.7000 1277.2500 ;
	    RECT 1177.5000 1277.1000 1179.3000 1277.2500 ;
	    RECT 1218.3000 1277.1000 1220.1000 1277.2500 ;
	    RECT 1491.9000 1278.7500 1493.7001 1278.9000 ;
	    RECT 1561.5000 1278.7500 1563.3000 1278.9000 ;
	    RECT 1491.9000 1277.2500 1563.3000 1278.7500 ;
	    RECT 1491.9000 1277.1000 1493.7001 1277.2500 ;
	    RECT 1561.5000 1277.1000 1563.3000 1277.2500 ;
	    RECT 35.1000 1272.7500 36.9000 1272.9000 ;
	    RECT 47.1000 1272.7500 48.9000 1272.9000 ;
	    RECT 35.1000 1271.2500 48.9000 1272.7500 ;
	    RECT 35.1000 1271.1000 36.9000 1271.2500 ;
	    RECT 47.1000 1271.1000 48.9000 1271.2500 ;
	    RECT 85.5000 1272.7500 87.3000 1272.9000 ;
	    RECT 95.1000 1272.7500 96.9000 1272.9000 ;
	    RECT 85.5000 1271.2500 96.9000 1272.7500 ;
	    RECT 85.5000 1271.1000 87.3000 1271.2500 ;
	    RECT 95.1000 1271.1000 96.9000 1271.2500 ;
	    RECT 231.9000 1272.7500 233.7000 1272.9000 ;
	    RECT 279.9000 1272.7500 281.7000 1272.9000 ;
	    RECT 231.9000 1271.2500 281.7000 1272.7500 ;
	    RECT 231.9000 1271.1000 233.7000 1271.2500 ;
	    RECT 279.9000 1271.1000 281.7000 1271.2500 ;
	    RECT 339.9000 1272.7500 341.7000 1272.9000 ;
	    RECT 363.9000 1272.7500 365.7000 1272.9000 ;
	    RECT 339.9000 1271.2500 365.7000 1272.7500 ;
	    RECT 339.9000 1271.1000 341.7000 1271.2500 ;
	    RECT 363.9000 1271.1000 365.7000 1271.2500 ;
	    RECT 419.1000 1272.7500 420.9000 1272.9000 ;
	    RECT 471.9000 1272.7500 473.7000 1272.9000 ;
	    RECT 419.1000 1271.2500 473.7000 1272.7500 ;
	    RECT 419.1000 1271.1000 420.9000 1271.2500 ;
	    RECT 471.9000 1271.1000 473.7000 1271.2500 ;
	    RECT 611.1000 1272.7500 612.9000 1272.9000 ;
	    RECT 752.7000 1272.7500 754.5000 1272.9000 ;
	    RECT 611.1000 1271.2500 754.5000 1272.7500 ;
	    RECT 611.1000 1271.1000 612.9000 1271.2500 ;
	    RECT 752.7000 1271.1000 754.5000 1271.2500 ;
	    RECT 884.7000 1272.7500 886.5000 1272.9000 ;
	    RECT 959.1000 1272.7500 960.9000 1272.9000 ;
	    RECT 884.7000 1271.2500 960.9000 1272.7500 ;
	    RECT 884.7000 1271.1000 886.5000 1271.2500 ;
	    RECT 959.1000 1271.1000 960.9000 1271.2500 ;
	    RECT 1167.9000 1272.7500 1169.7001 1272.9000 ;
	    RECT 1256.7001 1272.7500 1258.5000 1272.9000 ;
	    RECT 1167.9000 1271.2500 1258.5000 1272.7500 ;
	    RECT 1167.9000 1271.1000 1169.7001 1271.2500 ;
	    RECT 1256.7001 1271.1000 1258.5000 1271.2500 ;
	    RECT 1477.5000 1272.7500 1479.3000 1272.9000 ;
	    RECT 1482.3000 1272.7500 1484.1000 1272.9000 ;
	    RECT 1477.5000 1271.2500 1484.1000 1272.7500 ;
	    RECT 1477.5000 1271.1000 1479.3000 1271.2500 ;
	    RECT 1482.3000 1271.1000 1484.1000 1271.2500 ;
	    RECT 114.3000 1266.7500 116.1000 1266.9000 ;
	    RECT 311.1000 1266.7500 312.9000 1266.9000 ;
	    RECT 114.3000 1265.2500 312.9000 1266.7500 ;
	    RECT 114.3000 1265.1000 116.1000 1265.2500 ;
	    RECT 311.1000 1265.1000 312.9000 1265.2500 ;
	    RECT 392.7000 1266.7500 394.5000 1266.9000 ;
	    RECT 464.7000 1266.7500 466.5000 1266.9000 ;
	    RECT 392.7000 1265.2500 466.5000 1266.7500 ;
	    RECT 392.7000 1265.1000 394.5000 1265.2500 ;
	    RECT 464.7000 1265.1000 466.5000 1265.2500 ;
	    RECT 551.1000 1266.7500 552.9000 1266.9000 ;
	    RECT 563.1000 1266.7500 564.9000 1266.9000 ;
	    RECT 551.1000 1265.2500 564.9000 1266.7500 ;
	    RECT 551.1000 1265.1000 552.9000 1265.2500 ;
	    RECT 563.1000 1265.1000 564.9000 1265.2500 ;
	    RECT 851.1000 1266.7500 852.9000 1266.9000 ;
	    RECT 911.1000 1266.7500 912.9000 1266.9000 ;
	    RECT 851.1000 1265.2500 912.9000 1266.7500 ;
	    RECT 851.1000 1265.1000 852.9000 1265.2500 ;
	    RECT 911.1000 1265.1000 912.9000 1265.2500 ;
	    RECT 944.7000 1266.7500 946.5000 1266.9000 ;
	    RECT 980.7000 1266.7500 982.5000 1266.9000 ;
	    RECT 944.7000 1265.2500 982.5000 1266.7500 ;
	    RECT 944.7000 1265.1000 946.5000 1265.2500 ;
	    RECT 980.7000 1265.1000 982.5000 1265.2500 ;
	    RECT 1191.9000 1266.7500 1193.7001 1266.9000 ;
	    RECT 1227.9000 1266.7500 1229.7001 1266.9000 ;
	    RECT 1191.9000 1265.2500 1229.7001 1266.7500 ;
	    RECT 1191.9000 1265.1000 1193.7001 1265.2500 ;
	    RECT 1227.9000 1265.1000 1229.7001 1265.2500 ;
	    RECT 1465.5000 1266.7500 1467.3000 1266.9000 ;
	    RECT 1475.1000 1266.7500 1476.9000 1266.9000 ;
	    RECT 1465.5000 1265.2500 1476.9000 1266.7500 ;
	    RECT 1465.5000 1265.1000 1467.3000 1265.2500 ;
	    RECT 1475.1000 1265.1000 1476.9000 1265.2500 ;
	    RECT 1487.1000 1266.7500 1488.9000 1266.9000 ;
	    RECT 1520.7001 1266.7500 1522.5000 1266.9000 ;
	    RECT 1487.1000 1265.2500 1522.5000 1266.7500 ;
	    RECT 1487.1000 1265.1000 1488.9000 1265.2500 ;
	    RECT 1520.7001 1265.1000 1522.5000 1265.2500 ;
	    RECT 56.7000 1260.7500 58.5000 1260.9000 ;
	    RECT 121.5000 1260.7500 123.3000 1260.9000 ;
	    RECT 174.3000 1260.7500 176.1000 1260.9000 ;
	    RECT 56.7000 1259.2500 176.1000 1260.7500 ;
	    RECT 56.7000 1259.1000 58.5000 1259.2500 ;
	    RECT 121.5000 1259.1000 123.3000 1259.2500 ;
	    RECT 174.3000 1259.1000 176.1000 1259.2500 ;
	    RECT 260.7000 1260.7500 262.5000 1260.9000 ;
	    RECT 294.3000 1260.7500 296.1000 1260.9000 ;
	    RECT 260.7000 1259.2500 296.1000 1260.7500 ;
	    RECT 260.7000 1259.1000 262.5000 1259.2500 ;
	    RECT 294.3000 1259.1000 296.1000 1259.2500 ;
	    RECT 399.9000 1260.7500 401.7000 1260.9000 ;
	    RECT 467.1000 1260.7500 468.9000 1260.9000 ;
	    RECT 531.9000 1260.7500 533.7000 1260.9000 ;
	    RECT 399.9000 1259.2500 533.7000 1260.7500 ;
	    RECT 399.9000 1259.1000 401.7000 1259.2500 ;
	    RECT 467.1000 1259.1000 468.9000 1259.2500 ;
	    RECT 531.9000 1259.1000 533.7000 1259.2500 ;
	    RECT 637.5000 1260.7500 639.3000 1260.9000 ;
	    RECT 644.7000 1260.7500 646.5000 1260.9000 ;
	    RECT 637.5000 1259.2500 646.5000 1260.7500 ;
	    RECT 637.5000 1259.1000 639.3000 1259.2500 ;
	    RECT 644.7000 1259.1000 646.5000 1259.2500 ;
	    RECT 651.9000 1260.7500 653.7000 1260.9000 ;
	    RECT 656.7000 1260.7500 658.5000 1260.9000 ;
	    RECT 651.9000 1259.2500 658.5000 1260.7500 ;
	    RECT 651.9000 1259.1000 653.7000 1259.2500 ;
	    RECT 656.7000 1259.1000 658.5000 1259.2500 ;
	    RECT 978.3000 1260.7500 980.1000 1260.9000 ;
	    RECT 983.1000 1260.7500 984.9000 1260.9000 ;
	    RECT 978.3000 1259.2500 984.9000 1260.7500 ;
	    RECT 978.3000 1259.1000 980.1000 1259.2500 ;
	    RECT 983.1000 1259.1000 984.9000 1259.2500 ;
	    RECT 1326.3000 1260.7500 1328.1000 1260.9000 ;
	    RECT 1333.5000 1260.7500 1335.3000 1260.9000 ;
	    RECT 1326.3000 1259.2500 1335.3000 1260.7500 ;
	    RECT 1326.3000 1259.1000 1328.1000 1259.2500 ;
	    RECT 1333.5000 1259.1000 1335.3000 1259.2500 ;
	    RECT 1458.3000 1260.7500 1460.1000 1260.9000 ;
	    RECT 1484.7001 1260.7500 1486.5000 1260.9000 ;
	    RECT 1458.3000 1259.2500 1486.5000 1260.7500 ;
	    RECT 1458.3000 1259.1000 1460.1000 1259.2500 ;
	    RECT 1484.7001 1259.1000 1486.5000 1259.2500 ;
	    RECT 296.7000 1254.7500 298.5000 1254.9000 ;
	    RECT 325.5000 1254.7500 327.3000 1254.9000 ;
	    RECT 296.7000 1253.2500 327.3000 1254.7500 ;
	    RECT 296.7000 1253.1000 298.5000 1253.2500 ;
	    RECT 325.5000 1253.1000 327.3000 1253.2500 ;
	    RECT 692.7000 1254.7500 694.5000 1254.9000 ;
	    RECT 767.1000 1254.7500 768.9000 1254.9000 ;
	    RECT 692.7000 1253.2500 768.9000 1254.7500 ;
	    RECT 692.7000 1253.1000 694.5000 1253.2500 ;
	    RECT 767.1000 1253.1000 768.9000 1253.2500 ;
	    RECT 776.7000 1254.7500 778.5000 1254.9000 ;
	    RECT 935.1000 1254.7500 936.9000 1254.9000 ;
	    RECT 963.9000 1254.7500 965.7000 1254.9000 ;
	    RECT 776.7000 1253.2500 965.7000 1254.7500 ;
	    RECT 776.7000 1253.1000 778.5000 1253.2500 ;
	    RECT 935.1000 1253.1000 936.9000 1253.2500 ;
	    RECT 963.9000 1253.1000 965.7000 1253.2500 ;
	    RECT 968.7000 1254.7500 970.5000 1254.9000 ;
	    RECT 999.9000 1254.7500 1001.7000 1254.9000 ;
	    RECT 968.7000 1253.2500 1001.7000 1254.7500 ;
	    RECT 968.7000 1253.1000 970.5000 1253.2500 ;
	    RECT 999.9000 1253.1000 1001.7000 1253.2500 ;
	    RECT 1167.9000 1254.7500 1169.7001 1254.9000 ;
	    RECT 1302.3000 1254.7500 1304.1000 1254.9000 ;
	    RECT 1167.9000 1253.2500 1304.1000 1254.7500 ;
	    RECT 1167.9000 1253.1000 1169.7001 1253.2500 ;
	    RECT 1302.3000 1253.1000 1304.1000 1253.2500 ;
	    RECT 1328.7001 1254.7500 1330.5000 1254.9000 ;
	    RECT 1472.7001 1254.7500 1474.5000 1254.9000 ;
	    RECT 1328.7001 1253.2500 1474.5000 1254.7500 ;
	    RECT 1328.7001 1253.1000 1330.5000 1253.2500 ;
	    RECT 1472.7001 1253.1000 1474.5000 1253.2500 ;
	    RECT 1477.5000 1254.7500 1479.3000 1254.9000 ;
	    RECT 1482.3000 1254.7500 1484.1000 1254.9000 ;
	    RECT 1513.5000 1254.7500 1515.3000 1254.9000 ;
	    RECT 1530.3000 1254.7500 1532.1000 1254.9000 ;
	    RECT 1477.5000 1253.2500 1532.1000 1254.7500 ;
	    RECT 1477.5000 1253.1000 1479.3000 1253.2500 ;
	    RECT 1482.3000 1253.1000 1484.1000 1253.2500 ;
	    RECT 1513.5000 1253.1000 1515.3000 1253.2500 ;
	    RECT 1530.3000 1253.1000 1532.1000 1253.2500 ;
	    RECT 656.7000 1250.1000 658.5000 1251.9000 ;
	    RECT 123.9000 1248.7500 125.7000 1248.9000 ;
	    RECT 145.5000 1248.7500 147.3000 1248.9000 ;
	    RECT 123.9000 1247.2500 147.3000 1248.7500 ;
	    RECT 123.9000 1247.1000 125.7000 1247.2500 ;
	    RECT 145.5000 1247.1000 147.3000 1247.2500 ;
	    RECT 162.3000 1248.7500 164.1000 1248.9000 ;
	    RECT 287.1000 1248.7500 288.9000 1248.9000 ;
	    RECT 162.3000 1247.2500 288.9000 1248.7500 ;
	    RECT 162.3000 1247.1000 164.1000 1247.2500 ;
	    RECT 287.1000 1247.1000 288.9000 1247.2500 ;
	    RECT 452.7000 1248.7500 454.5000 1248.9000 ;
	    RECT 479.1000 1248.7500 480.9000 1248.9000 ;
	    RECT 452.7000 1247.2500 480.9000 1248.7500 ;
	    RECT 656.8500 1248.7500 658.3500 1250.1000 ;
	    RECT 661.5000 1248.7500 663.3000 1248.9000 ;
	    RECT 656.8500 1247.2500 663.3000 1248.7500 ;
	    RECT 452.7000 1247.1000 454.5000 1247.2500 ;
	    RECT 479.1000 1247.1000 480.9000 1247.2500 ;
	    RECT 661.5000 1247.1000 663.3000 1247.2500 ;
	    RECT 807.9000 1248.7500 809.7000 1248.9000 ;
	    RECT 831.9000 1248.7500 833.7000 1248.9000 ;
	    RECT 807.9000 1247.2500 833.7000 1248.7500 ;
	    RECT 807.9000 1247.1000 809.7000 1247.2500 ;
	    RECT 831.9000 1247.1000 833.7000 1247.2500 ;
	    RECT 870.3000 1248.7500 872.1000 1248.9000 ;
	    RECT 954.3000 1248.7500 956.1000 1248.9000 ;
	    RECT 870.3000 1247.2500 956.1000 1248.7500 ;
	    RECT 870.3000 1247.1000 872.1000 1247.2500 ;
	    RECT 954.3000 1247.1000 956.1000 1247.2500 ;
	    RECT 973.5000 1248.7500 975.3000 1248.9000 ;
	    RECT 1112.7001 1248.7500 1114.5000 1248.9000 ;
	    RECT 973.5000 1247.2500 1114.5000 1248.7500 ;
	    RECT 973.5000 1247.1000 975.3000 1247.2500 ;
	    RECT 1112.7001 1247.1000 1114.5000 1247.2500 ;
	    RECT 1122.3000 1248.7500 1124.1000 1248.9000 ;
	    RECT 1134.3000 1248.7500 1136.1000 1248.9000 ;
	    RECT 1122.3000 1247.2500 1136.1000 1248.7500 ;
	    RECT 1122.3000 1247.1000 1124.1000 1247.2500 ;
	    RECT 1134.3000 1247.1000 1136.1000 1247.2500 ;
	    RECT 1158.3000 1248.7500 1160.1000 1248.9000 ;
	    RECT 1163.1000 1248.7500 1164.9000 1248.9000 ;
	    RECT 1158.3000 1247.2500 1164.9000 1248.7500 ;
	    RECT 1158.3000 1247.1000 1160.1000 1247.2500 ;
	    RECT 1163.1000 1247.1000 1164.9000 1247.2500 ;
	    RECT 1427.1000 1248.7500 1428.9000 1248.9000 ;
	    RECT 1463.1000 1248.7500 1464.9000 1248.9000 ;
	    RECT 1427.1000 1247.2500 1464.9000 1248.7500 ;
	    RECT 1427.1000 1247.1000 1428.9000 1247.2500 ;
	    RECT 1463.1000 1247.1000 1464.9000 1247.2500 ;
	    RECT 1496.7001 1248.7500 1498.5000 1248.9000 ;
	    RECT 1563.9000 1248.7500 1565.7001 1248.9000 ;
	    RECT 1496.7001 1247.2500 1565.7001 1248.7500 ;
	    RECT 1496.7001 1247.1000 1498.5000 1247.2500 ;
	    RECT 1563.9000 1247.1000 1565.7001 1247.2500 ;
	    RECT 750.3000 1242.7500 752.1000 1242.9000 ;
	    RECT 757.5000 1242.7500 759.3000 1242.9000 ;
	    RECT 750.3000 1241.2500 759.3000 1242.7500 ;
	    RECT 750.3000 1241.1000 752.1000 1241.2500 ;
	    RECT 757.5000 1241.1000 759.3000 1241.2500 ;
	    RECT 805.5000 1242.7500 807.3000 1242.9000 ;
	    RECT 913.5000 1242.7500 915.3000 1242.9000 ;
	    RECT 949.5000 1242.7500 951.3000 1242.9000 ;
	    RECT 805.5000 1241.2500 951.3000 1242.7500 ;
	    RECT 805.5000 1241.1000 807.3000 1241.2500 ;
	    RECT 913.5000 1241.1000 915.3000 1241.2500 ;
	    RECT 949.5000 1241.1000 951.3000 1241.2500 ;
	    RECT 1297.5000 1242.7500 1299.3000 1242.9000 ;
	    RECT 1319.1000 1242.7500 1320.9000 1242.9000 ;
	    RECT 1297.5000 1241.2500 1320.9000 1242.7500 ;
	    RECT 1297.5000 1241.1000 1299.3000 1241.2500 ;
	    RECT 1319.1000 1241.1000 1320.9000 1241.2500 ;
	    RECT 1376.7001 1242.7500 1378.5000 1242.9000 ;
	    RECT 1451.1000 1242.7500 1452.9000 1242.9000 ;
	    RECT 1458.3000 1242.7500 1460.1000 1242.9000 ;
	    RECT 1376.7001 1241.2500 1460.1000 1242.7500 ;
	    RECT 1376.7001 1241.1000 1378.5000 1241.2500 ;
	    RECT 1451.1000 1241.1000 1452.9000 1241.2500 ;
	    RECT 1458.3000 1241.1000 1460.1000 1241.2500 ;
	    RECT 1463.1000 1242.7500 1464.9000 1242.9000 ;
	    RECT 1530.3000 1242.7500 1532.1000 1242.9000 ;
	    RECT 1463.1000 1241.2500 1532.1000 1242.7500 ;
	    RECT 1463.1000 1241.1000 1464.9000 1241.2500 ;
	    RECT 1530.3000 1241.1000 1532.1000 1241.2500 ;
	    RECT 258.3000 1236.7500 260.1000 1236.9000 ;
	    RECT 335.1000 1236.7500 336.9000 1236.9000 ;
	    RECT 258.3000 1235.2500 336.9000 1236.7500 ;
	    RECT 258.3000 1235.1000 260.1000 1235.2500 ;
	    RECT 335.1000 1235.1000 336.9000 1235.2500 ;
	    RECT 596.7000 1236.7500 598.5000 1236.9000 ;
	    RECT 642.3000 1236.7500 644.1000 1236.9000 ;
	    RECT 596.7000 1235.2500 644.1000 1236.7500 ;
	    RECT 596.7000 1235.1000 598.5000 1235.2500 ;
	    RECT 642.3000 1235.1000 644.1000 1235.2500 ;
	    RECT 755.1000 1236.7500 756.9000 1236.9000 ;
	    RECT 906.3000 1236.7500 908.1000 1236.9000 ;
	    RECT 755.1000 1235.2500 908.1000 1236.7500 ;
	    RECT 755.1000 1235.1000 756.9000 1235.2500 ;
	    RECT 906.3000 1235.1000 908.1000 1235.2500 ;
	    RECT 1391.1000 1236.7500 1392.9000 1236.9000 ;
	    RECT 1415.1000 1236.7500 1416.9000 1236.9000 ;
	    RECT 1482.3000 1236.7500 1484.1000 1236.9000 ;
	    RECT 1391.1000 1235.2500 1484.1000 1236.7500 ;
	    RECT 1391.1000 1235.1000 1392.9000 1235.2500 ;
	    RECT 1415.1000 1235.1000 1416.9000 1235.2500 ;
	    RECT 1482.3000 1235.1000 1484.1000 1235.2500 ;
	    RECT 1489.5000 1236.7500 1491.3000 1236.9000 ;
	    RECT 1527.9000 1236.7500 1529.7001 1236.9000 ;
	    RECT 1489.5000 1235.2500 1529.7001 1236.7500 ;
	    RECT 1489.5000 1235.1000 1491.3000 1235.2500 ;
	    RECT 1527.9000 1235.1000 1529.7001 1235.2500 ;
	    RECT 83.1000 1230.7500 84.9000 1230.9000 ;
	    RECT 143.1000 1230.7500 144.9000 1230.9000 ;
	    RECT 83.1000 1229.2500 144.9000 1230.7500 ;
	    RECT 83.1000 1229.1000 84.9000 1229.2500 ;
	    RECT 143.1000 1229.1000 144.9000 1229.2500 ;
	    RECT 335.1000 1230.7500 336.9000 1230.9000 ;
	    RECT 385.5000 1230.7500 387.3000 1230.9000 ;
	    RECT 426.3000 1230.7500 428.1000 1230.9000 ;
	    RECT 335.1000 1229.2500 428.1000 1230.7500 ;
	    RECT 335.1000 1229.1000 336.9000 1229.2500 ;
	    RECT 385.5000 1229.1000 387.3000 1229.2500 ;
	    RECT 426.3000 1229.1000 428.1000 1229.2500 ;
	    RECT 479.1000 1230.7500 480.9000 1230.9000 ;
	    RECT 553.5000 1230.7500 555.3000 1230.9000 ;
	    RECT 479.1000 1229.2500 555.3000 1230.7500 ;
	    RECT 479.1000 1229.1000 480.9000 1229.2500 ;
	    RECT 553.5000 1229.1000 555.3000 1229.2500 ;
	    RECT 623.1000 1230.7500 624.9000 1230.9000 ;
	    RECT 649.5000 1230.7500 651.3000 1230.9000 ;
	    RECT 623.1000 1229.2500 651.3000 1230.7500 ;
	    RECT 623.1000 1229.1000 624.9000 1229.2500 ;
	    RECT 649.5000 1229.1000 651.3000 1229.2500 ;
	    RECT 863.1000 1230.7500 864.9000 1230.9000 ;
	    RECT 872.7000 1230.7500 874.5000 1230.9000 ;
	    RECT 863.1000 1229.2500 874.5000 1230.7500 ;
	    RECT 863.1000 1229.1000 864.9000 1229.2500 ;
	    RECT 872.7000 1229.1000 874.5000 1229.2500 ;
	    RECT 877.5000 1230.7500 879.3000 1230.9000 ;
	    RECT 889.5000 1230.7500 891.3000 1230.9000 ;
	    RECT 877.5000 1229.2500 891.3000 1230.7500 ;
	    RECT 877.5000 1229.1000 879.3000 1229.2500 ;
	    RECT 889.5000 1229.1000 891.3000 1229.2500 ;
	    RECT 935.1000 1230.7500 936.9000 1230.9000 ;
	    RECT 1019.1000 1230.7500 1020.9000 1230.9000 ;
	    RECT 935.1000 1229.2500 1020.9000 1230.7500 ;
	    RECT 935.1000 1229.1000 936.9000 1229.2500 ;
	    RECT 1019.1000 1229.1000 1020.9000 1229.2500 ;
	    RECT 1035.9000 1230.7500 1037.7001 1230.9000 ;
	    RECT 1083.9000 1230.7500 1085.7001 1230.9000 ;
	    RECT 1035.9000 1229.2500 1085.7001 1230.7500 ;
	    RECT 1035.9000 1229.1000 1037.7001 1229.2500 ;
	    RECT 1083.9000 1229.1000 1085.7001 1229.2500 ;
	    RECT 1232.7001 1230.7500 1234.5000 1230.9000 ;
	    RECT 1295.1000 1230.7500 1296.9000 1230.9000 ;
	    RECT 1232.7001 1229.2500 1296.9000 1230.7500 ;
	    RECT 1232.7001 1229.1000 1234.5000 1229.2500 ;
	    RECT 1295.1000 1229.1000 1296.9000 1229.2500 ;
	    RECT 1391.1000 1230.7500 1392.9000 1230.9000 ;
	    RECT 1477.5000 1230.7500 1479.3000 1230.9000 ;
	    RECT 1489.5000 1230.7500 1491.3000 1230.9000 ;
	    RECT 1391.1000 1229.2500 1491.3000 1230.7500 ;
	    RECT 1391.1000 1229.1000 1392.9000 1229.2500 ;
	    RECT 1477.5000 1229.1000 1479.3000 1229.2500 ;
	    RECT 1489.5000 1229.1000 1491.3000 1229.2500 ;
	    RECT 1544.7001 1230.7500 1546.5000 1230.9000 ;
	    RECT 1549.5000 1230.7500 1551.3000 1230.9000 ;
	    RECT 1544.7001 1229.2500 1551.3000 1230.7500 ;
	    RECT 1544.7001 1229.1000 1546.5000 1229.2500 ;
	    RECT 1549.5000 1229.1000 1551.3000 1229.2500 ;
	    RECT 251.1000 1224.7500 252.9000 1224.9000 ;
	    RECT 284.7000 1224.7500 286.5000 1224.9000 ;
	    RECT 251.1000 1223.2500 286.5000 1224.7500 ;
	    RECT 251.1000 1223.1000 252.9000 1223.2500 ;
	    RECT 284.7000 1223.1000 286.5000 1223.2500 ;
	    RECT 867.9000 1224.7500 869.7000 1224.9000 ;
	    RECT 875.1000 1224.7500 876.9000 1224.9000 ;
	    RECT 867.9000 1223.2500 876.9000 1224.7500 ;
	    RECT 867.9000 1223.1000 869.7000 1223.2500 ;
	    RECT 875.1000 1223.1000 876.9000 1223.2500 ;
	    RECT 1011.9000 1224.7500 1013.7000 1224.9000 ;
	    RECT 1059.9000 1224.7500 1061.7001 1224.9000 ;
	    RECT 1011.9000 1223.2500 1061.7001 1224.7500 ;
	    RECT 1011.9000 1223.1000 1013.7000 1223.2500 ;
	    RECT 1059.9000 1223.1000 1061.7001 1223.2500 ;
	    RECT 1069.5000 1224.7500 1071.3000 1224.9000 ;
	    RECT 1165.5000 1224.7500 1167.3000 1224.9000 ;
	    RECT 1069.5000 1223.2500 1167.3000 1224.7500 ;
	    RECT 1069.5000 1223.1000 1071.3000 1223.2500 ;
	    RECT 1165.5000 1223.1000 1167.3000 1223.2500 ;
	    RECT 1369.5000 1224.7500 1371.3000 1224.9000 ;
	    RECT 1386.3000 1224.7500 1388.1000 1224.9000 ;
	    RECT 1369.5000 1223.2500 1388.1000 1224.7500 ;
	    RECT 1369.5000 1223.1000 1371.3000 1223.2500 ;
	    RECT 1386.3000 1223.1000 1388.1000 1223.2500 ;
	    RECT 308.7000 1218.7500 310.5000 1218.9000 ;
	    RECT 344.7000 1218.7500 346.5000 1218.9000 ;
	    RECT 383.1000 1218.7500 384.9000 1218.9000 ;
	    RECT 390.3000 1218.7500 392.1000 1218.9000 ;
	    RECT 308.7000 1217.2500 392.1000 1218.7500 ;
	    RECT 308.7000 1217.1000 310.5000 1217.2500 ;
	    RECT 344.7000 1217.1000 346.5000 1217.2500 ;
	    RECT 383.1000 1217.1000 384.9000 1217.2500 ;
	    RECT 390.3000 1217.1000 392.1000 1217.2500 ;
	    RECT 771.9000 1218.7500 773.7000 1218.9000 ;
	    RECT 846.3000 1218.7500 848.1000 1218.9000 ;
	    RECT 771.9000 1217.2500 848.1000 1218.7500 ;
	    RECT 771.9000 1217.1000 773.7000 1217.2500 ;
	    RECT 846.3000 1217.1000 848.1000 1217.2500 ;
	    RECT 865.5000 1218.7500 867.3000 1218.9000 ;
	    RECT 906.3000 1218.7500 908.1000 1218.9000 ;
	    RECT 865.5000 1217.2500 908.1000 1218.7500 ;
	    RECT 865.5000 1217.1000 867.3000 1217.2500 ;
	    RECT 906.3000 1217.1000 908.1000 1217.2500 ;
	    RECT 927.9000 1218.7500 929.7000 1218.9000 ;
	    RECT 949.5000 1218.7500 951.3000 1218.9000 ;
	    RECT 927.9000 1217.2500 951.3000 1218.7500 ;
	    RECT 927.9000 1217.1000 929.7000 1217.2500 ;
	    RECT 949.5000 1217.1000 951.3000 1217.2500 ;
	    RECT 971.1000 1218.7500 972.9000 1218.9000 ;
	    RECT 978.3000 1218.7500 980.1000 1218.9000 ;
	    RECT 971.1000 1217.2500 980.1000 1218.7500 ;
	    RECT 971.1000 1217.1000 972.9000 1217.2500 ;
	    RECT 978.3000 1217.1000 980.1000 1217.2500 ;
	    RECT 1196.7001 1218.7500 1198.5000 1218.9000 ;
	    RECT 1319.1000 1218.7500 1320.9000 1218.9000 ;
	    RECT 1196.7001 1217.2500 1320.9000 1218.7500 ;
	    RECT 1196.7001 1217.1000 1198.5000 1217.2500 ;
	    RECT 1319.1000 1217.1000 1320.9000 1217.2500 ;
	    RECT 246.3000 1212.7500 248.1000 1212.9000 ;
	    RECT 277.5000 1212.7500 279.3000 1212.9000 ;
	    RECT 246.3000 1211.2500 279.3000 1212.7500 ;
	    RECT 246.3000 1211.1000 248.1000 1211.2500 ;
	    RECT 277.5000 1211.1000 279.3000 1211.2500 ;
	    RECT 349.5000 1212.7500 351.3000 1212.9000 ;
	    RECT 361.5000 1212.7500 363.3000 1212.9000 ;
	    RECT 349.5000 1211.2500 363.3000 1212.7500 ;
	    RECT 349.5000 1211.1000 351.3000 1211.2500 ;
	    RECT 361.5000 1211.1000 363.3000 1211.2500 ;
	    RECT 932.7000 1212.7500 934.5000 1212.9000 ;
	    RECT 951.9000 1212.7500 953.7000 1212.9000 ;
	    RECT 932.7000 1211.2500 953.7000 1212.7500 ;
	    RECT 932.7000 1211.1000 934.5000 1211.2500 ;
	    RECT 951.9000 1211.1000 953.7000 1211.2500 ;
	    RECT 1057.5000 1212.7500 1059.3000 1212.9000 ;
	    RECT 1232.7001 1212.7500 1234.5000 1212.9000 ;
	    RECT 1057.5000 1211.2500 1234.5000 1212.7500 ;
	    RECT 1057.5000 1211.1000 1059.3000 1211.2500 ;
	    RECT 1232.7001 1211.1000 1234.5000 1211.2500 ;
	    RECT 1319.1000 1212.7500 1320.9000 1212.9000 ;
	    RECT 1391.1000 1212.7500 1392.9000 1212.9000 ;
	    RECT 1319.1000 1211.2500 1392.9000 1212.7500 ;
	    RECT 1319.1000 1211.1000 1320.9000 1211.2500 ;
	    RECT 1391.1000 1211.1000 1392.9000 1211.2500 ;
	    RECT 1523.1000 1212.7500 1524.9000 1212.9000 ;
	    RECT 1535.1000 1212.7500 1536.9000 1212.9000 ;
	    RECT 1523.1000 1211.2500 1536.9000 1212.7500 ;
	    RECT 1523.1000 1211.1000 1524.9000 1211.2500 ;
	    RECT 1535.1000 1211.1000 1536.9000 1211.2500 ;
	    RECT 251.1000 1206.7500 252.9000 1206.9000 ;
	    RECT 287.1000 1206.7500 288.9000 1206.9000 ;
	    RECT 251.1000 1205.2500 288.9000 1206.7500 ;
	    RECT 251.1000 1205.1000 252.9000 1205.2500 ;
	    RECT 287.1000 1205.1000 288.9000 1205.2500 ;
	    RECT 524.7000 1206.7500 526.5000 1206.9000 ;
	    RECT 563.1000 1206.7500 564.9000 1206.9000 ;
	    RECT 524.7000 1205.2500 564.9000 1206.7500 ;
	    RECT 524.7000 1205.1000 526.5000 1205.2500 ;
	    RECT 563.1000 1205.1000 564.9000 1205.2500 ;
	    RECT 692.7000 1206.7500 694.5000 1206.9000 ;
	    RECT 721.5000 1206.7500 723.3000 1206.9000 ;
	    RECT 692.7000 1205.2500 723.3000 1206.7500 ;
	    RECT 692.7000 1205.1000 694.5000 1205.2500 ;
	    RECT 721.5000 1205.1000 723.3000 1205.2500 ;
	    RECT 925.5000 1206.7500 927.3000 1206.9000 ;
	    RECT 973.5000 1206.7500 975.3000 1206.9000 ;
	    RECT 925.5000 1205.2500 975.3000 1206.7500 ;
	    RECT 925.5000 1205.1000 927.3000 1205.2500 ;
	    RECT 973.5000 1205.1000 975.3000 1205.2500 ;
	    RECT 1033.5000 1206.7500 1035.3000 1206.9000 ;
	    RECT 1074.3000 1206.7500 1076.1000 1206.9000 ;
	    RECT 1033.5000 1205.2500 1076.1000 1206.7500 ;
	    RECT 1033.5000 1205.1000 1035.3000 1205.2500 ;
	    RECT 1074.3000 1205.1000 1076.1000 1205.2500 ;
	    RECT 1518.3000 1206.7500 1520.1000 1206.9000 ;
	    RECT 1523.1000 1206.7500 1524.9000 1206.9000 ;
	    RECT 1518.3000 1205.2500 1524.9000 1206.7500 ;
	    RECT 1518.3000 1205.1000 1520.1000 1205.2500 ;
	    RECT 1523.1000 1205.1000 1524.9000 1205.2500 ;
	    RECT 1535.1000 1206.7500 1536.9000 1206.9000 ;
	    RECT 1551.9000 1206.7500 1553.7001 1206.9000 ;
	    RECT 1535.1000 1205.2500 1553.7001 1206.7500 ;
	    RECT 1535.1000 1205.1000 1536.9000 1205.2500 ;
	    RECT 1551.9000 1205.1000 1553.7001 1205.2500 ;
	    RECT 155.1000 1200.7500 156.9000 1200.9000 ;
	    RECT 169.5000 1200.7500 171.3000 1200.9000 ;
	    RECT 155.1000 1199.2500 171.3000 1200.7500 ;
	    RECT 155.1000 1199.1000 156.9000 1199.2500 ;
	    RECT 169.5000 1199.1000 171.3000 1199.2500 ;
	    RECT 239.1000 1200.7500 240.9000 1200.9000 ;
	    RECT 272.7000 1200.7500 274.5000 1200.9000 ;
	    RECT 239.1000 1199.2500 274.5000 1200.7500 ;
	    RECT 239.1000 1199.1000 240.9000 1199.2500 ;
	    RECT 272.7000 1199.1000 274.5000 1199.2500 ;
	    RECT 277.5000 1200.7500 279.3000 1200.9000 ;
	    RECT 308.7000 1200.7500 310.5000 1200.9000 ;
	    RECT 277.5000 1199.2500 310.5000 1200.7500 ;
	    RECT 277.5000 1199.1000 279.3000 1199.2500 ;
	    RECT 308.7000 1199.1000 310.5000 1199.2500 ;
	    RECT 459.9000 1200.7500 461.7000 1200.9000 ;
	    RECT 476.7000 1200.7500 478.5000 1200.9000 ;
	    RECT 459.9000 1199.2500 478.5000 1200.7500 ;
	    RECT 459.9000 1199.1000 461.7000 1199.2500 ;
	    RECT 476.7000 1199.1000 478.5000 1199.2500 ;
	    RECT 642.3000 1200.7500 644.1000 1200.9000 ;
	    RECT 651.9000 1200.7500 653.7000 1200.9000 ;
	    RECT 642.3000 1199.2500 653.7000 1200.7500 ;
	    RECT 642.3000 1199.1000 644.1000 1199.2500 ;
	    RECT 651.9000 1199.1000 653.7000 1199.2500 ;
	    RECT 721.5000 1200.7500 723.3000 1200.9000 ;
	    RECT 747.9000 1200.7500 749.7000 1200.9000 ;
	    RECT 721.5000 1199.2500 749.7000 1200.7500 ;
	    RECT 721.5000 1199.1000 723.3000 1199.2500 ;
	    RECT 747.9000 1199.1000 749.7000 1199.2500 ;
	    RECT 947.1000 1200.7500 948.9000 1200.9000 ;
	    RECT 956.7000 1200.7500 958.5000 1200.9000 ;
	    RECT 947.1000 1199.2500 958.5000 1200.7500 ;
	    RECT 947.1000 1199.1000 948.9000 1199.2500 ;
	    RECT 956.7000 1199.1000 958.5000 1199.2500 ;
	    RECT 1038.3000 1200.7500 1040.1000 1200.9000 ;
	    RECT 1079.1000 1200.7500 1080.9000 1200.9000 ;
	    RECT 1038.3000 1199.2500 1080.9000 1200.7500 ;
	    RECT 1038.3000 1199.1000 1040.1000 1199.2500 ;
	    RECT 1079.1000 1199.1000 1080.9000 1199.2500 ;
	    RECT 1309.5000 1200.7500 1311.3000 1200.9000 ;
	    RECT 1316.7001 1200.7500 1318.5000 1200.9000 ;
	    RECT 1309.5000 1199.2500 1318.5000 1200.7500 ;
	    RECT 1309.5000 1199.1000 1311.3000 1199.2500 ;
	    RECT 1316.7001 1199.1000 1318.5000 1199.2500 ;
	    RECT 1523.1000 1200.7500 1524.9000 1200.9000 ;
	    RECT 1530.3000 1200.7500 1532.1000 1200.9000 ;
	    RECT 1523.1000 1199.2500 1532.1000 1200.7500 ;
	    RECT 1523.1000 1199.1000 1524.9000 1199.2500 ;
	    RECT 1530.3000 1199.1000 1532.1000 1199.2500 ;
	    RECT 246.3000 1194.7500 248.1000 1194.9000 ;
	    RECT 270.3000 1194.7500 272.1000 1194.9000 ;
	    RECT 246.3000 1193.2500 272.1000 1194.7500 ;
	    RECT 246.3000 1193.1000 248.1000 1193.2500 ;
	    RECT 270.3000 1193.1000 272.1000 1193.2500 ;
	    RECT 476.7000 1194.7500 478.5000 1194.9000 ;
	    RECT 570.3000 1194.7500 572.1000 1194.9000 ;
	    RECT 476.7000 1193.2500 572.1000 1194.7500 ;
	    RECT 476.7000 1193.1000 478.5000 1193.2500 ;
	    RECT 570.3000 1193.1000 572.1000 1193.2500 ;
	    RECT 889.5000 1194.7500 891.3000 1194.9000 ;
	    RECT 1074.3000 1194.7500 1076.1000 1194.9000 ;
	    RECT 889.5000 1193.2500 1076.1000 1194.7500 ;
	    RECT 889.5000 1193.1000 891.3000 1193.2500 ;
	    RECT 1074.3000 1193.1000 1076.1000 1193.2500 ;
	    RECT 1079.1000 1194.7500 1080.9000 1194.9000 ;
	    RECT 1088.7001 1194.7500 1090.5000 1194.9000 ;
	    RECT 1155.9000 1194.7500 1157.7001 1194.9000 ;
	    RECT 1079.1000 1193.2500 1157.7001 1194.7500 ;
	    RECT 1079.1000 1193.1000 1080.9000 1193.2500 ;
	    RECT 1088.7001 1193.1000 1090.5000 1193.2500 ;
	    RECT 1155.9000 1193.1000 1157.7001 1193.2500 ;
	    RECT 1441.5000 1194.7500 1443.3000 1194.9000 ;
	    RECT 1513.5000 1194.7500 1515.3000 1194.9000 ;
	    RECT 1441.5000 1193.2500 1515.3000 1194.7500 ;
	    RECT 1441.5000 1193.1000 1443.3000 1193.2500 ;
	    RECT 1513.5000 1193.1000 1515.3000 1193.2500 ;
	    RECT 1530.3000 1194.7500 1532.1000 1194.9000 ;
	    RECT 1539.9000 1194.7500 1541.7001 1194.9000 ;
	    RECT 1530.3000 1193.2500 1541.7001 1194.7500 ;
	    RECT 1530.3000 1193.1000 1532.1000 1193.2500 ;
	    RECT 1539.9000 1193.1000 1541.7001 1193.2500 ;
	    RECT 1544.7001 1194.7500 1546.5000 1194.9000 ;
	    RECT 1554.3000 1194.7500 1556.1000 1194.9000 ;
	    RECT 1544.7001 1193.2500 1556.1000 1194.7500 ;
	    RECT 1544.7001 1193.1000 1546.5000 1193.2500 ;
	    RECT 1554.3000 1193.1000 1556.1000 1193.2500 ;
	    RECT 23.1000 1188.7500 24.9000 1188.9000 ;
	    RECT 54.3000 1188.7500 56.1000 1188.9000 ;
	    RECT 188.7000 1188.7500 190.5000 1188.9000 ;
	    RECT 23.1000 1187.2500 190.5000 1188.7500 ;
	    RECT 23.1000 1187.1000 24.9000 1187.2500 ;
	    RECT 54.3000 1187.1000 56.1000 1187.2500 ;
	    RECT 188.7000 1187.1000 190.5000 1187.2500 ;
	    RECT 255.9000 1188.7500 257.7000 1188.9000 ;
	    RECT 260.7000 1188.7500 262.5000 1188.9000 ;
	    RECT 255.9000 1187.2500 262.5000 1188.7500 ;
	    RECT 255.9000 1187.1000 257.7000 1187.2500 ;
	    RECT 260.7000 1187.1000 262.5000 1187.2500 ;
	    RECT 505.5000 1188.7500 507.3000 1188.9000 ;
	    RECT 577.5000 1188.7500 579.3000 1188.9000 ;
	    RECT 505.5000 1187.2500 579.3000 1188.7500 ;
	    RECT 505.5000 1187.1000 507.3000 1187.2500 ;
	    RECT 577.5000 1187.1000 579.3000 1187.2500 ;
	    RECT 745.5000 1188.7500 747.3000 1188.9000 ;
	    RECT 774.3000 1188.7500 776.1000 1188.9000 ;
	    RECT 745.5000 1187.2500 776.1000 1188.7500 ;
	    RECT 745.5000 1187.1000 747.3000 1187.2500 ;
	    RECT 774.3000 1187.1000 776.1000 1187.2500 ;
	    RECT 827.1000 1188.7500 828.9000 1188.9000 ;
	    RECT 839.1000 1188.7500 840.9000 1188.9000 ;
	    RECT 827.1000 1187.2500 840.9000 1188.7500 ;
	    RECT 827.1000 1187.1000 828.9000 1187.2500 ;
	    RECT 839.1000 1187.1000 840.9000 1187.2500 ;
	    RECT 843.9000 1188.7500 845.7000 1188.9000 ;
	    RECT 872.7000 1188.7500 874.5000 1188.9000 ;
	    RECT 843.9000 1187.2500 874.5000 1188.7500 ;
	    RECT 843.9000 1187.1000 845.7000 1187.2500 ;
	    RECT 872.7000 1187.1000 874.5000 1187.2500 ;
	    RECT 966.3000 1188.7500 968.1000 1188.9000 ;
	    RECT 1023.9000 1188.7500 1025.7001 1188.9000 ;
	    RECT 966.3000 1187.2500 1025.7001 1188.7500 ;
	    RECT 966.3000 1187.1000 968.1000 1187.2500 ;
	    RECT 1023.9000 1187.1000 1025.7001 1187.2500 ;
	    RECT 1079.1000 1188.7500 1080.9000 1188.9000 ;
	    RECT 1256.7001 1188.7500 1258.5000 1188.9000 ;
	    RECT 1304.7001 1188.7500 1306.5000 1188.9000 ;
	    RECT 1079.1000 1187.2500 1306.5000 1188.7500 ;
	    RECT 1079.1000 1187.1000 1080.9000 1187.2500 ;
	    RECT 1256.7001 1187.1000 1258.5000 1187.2500 ;
	    RECT 1304.7001 1187.1000 1306.5000 1187.2500 ;
	    RECT 18.3000 1182.7500 20.1000 1182.9000 ;
	    RECT 32.7000 1182.7500 34.5000 1182.9000 ;
	    RECT 18.3000 1181.2500 34.5000 1182.7500 ;
	    RECT 18.3000 1181.1000 20.1000 1181.2500 ;
	    RECT 32.7000 1181.1000 34.5000 1181.2500 ;
	    RECT 59.1000 1182.7500 60.9000 1182.9000 ;
	    RECT 80.7000 1182.7500 82.5000 1182.9000 ;
	    RECT 59.1000 1181.2500 82.5000 1182.7500 ;
	    RECT 59.1000 1181.1000 60.9000 1181.2500 ;
	    RECT 80.7000 1181.1000 82.5000 1181.2500 ;
	    RECT 90.3000 1182.7500 92.1000 1182.9000 ;
	    RECT 114.3000 1182.7500 116.1000 1182.9000 ;
	    RECT 90.3000 1181.2500 116.1000 1182.7500 ;
	    RECT 90.3000 1181.1000 92.1000 1181.2500 ;
	    RECT 114.3000 1181.1000 116.1000 1181.2500 ;
	    RECT 241.5000 1182.7500 243.3000 1182.9000 ;
	    RECT 260.7000 1182.7500 262.5000 1182.9000 ;
	    RECT 241.5000 1181.2500 262.5000 1182.7500 ;
	    RECT 241.5000 1181.1000 243.3000 1181.2500 ;
	    RECT 260.7000 1181.1000 262.5000 1181.2500 ;
	    RECT 500.7000 1182.7500 502.5000 1182.9000 ;
	    RECT 529.5000 1182.7500 531.3000 1182.9000 ;
	    RECT 500.7000 1181.2500 531.3000 1182.7500 ;
	    RECT 500.7000 1181.1000 502.5000 1181.2500 ;
	    RECT 529.5000 1181.1000 531.3000 1181.2500 ;
	    RECT 546.3000 1182.7500 548.1000 1182.9000 ;
	    RECT 579.9000 1182.7500 581.7000 1182.9000 ;
	    RECT 546.3000 1181.2500 581.7000 1182.7500 ;
	    RECT 546.3000 1181.1000 548.1000 1181.2500 ;
	    RECT 579.9000 1181.1000 581.7000 1181.2500 ;
	    RECT 695.1000 1182.7500 696.9000 1182.9000 ;
	    RECT 709.5000 1182.7500 711.3000 1182.9000 ;
	    RECT 695.1000 1181.2500 711.3000 1182.7500 ;
	    RECT 695.1000 1181.1000 696.9000 1181.2500 ;
	    RECT 709.5000 1181.1000 711.3000 1181.2500 ;
	    RECT 723.9000 1182.7500 725.7000 1182.9000 ;
	    RECT 851.1000 1182.7500 852.9000 1182.9000 ;
	    RECT 723.9000 1181.2500 852.9000 1182.7500 ;
	    RECT 723.9000 1181.1000 725.7000 1181.2500 ;
	    RECT 851.1000 1181.1000 852.9000 1181.2500 ;
	    RECT 891.9000 1182.7500 893.7000 1182.9000 ;
	    RECT 899.1000 1182.7500 900.9000 1182.9000 ;
	    RECT 891.9000 1181.2500 900.9000 1182.7500 ;
	    RECT 891.9000 1181.1000 893.7000 1181.2500 ;
	    RECT 899.1000 1181.1000 900.9000 1181.2500 ;
	    RECT 923.1000 1182.7500 924.9000 1182.9000 ;
	    RECT 963.9000 1182.7500 965.7000 1182.9000 ;
	    RECT 923.1000 1181.2500 965.7000 1182.7500 ;
	    RECT 923.1000 1181.1000 924.9000 1181.2500 ;
	    RECT 963.9000 1181.1000 965.7000 1181.2500 ;
	    RECT 975.9000 1182.7500 977.7000 1182.9000 ;
	    RECT 983.1000 1182.7500 984.9000 1182.9000 ;
	    RECT 975.9000 1181.2500 984.9000 1182.7500 ;
	    RECT 975.9000 1181.1000 977.7000 1181.2500 ;
	    RECT 983.1000 1181.1000 984.9000 1181.2500 ;
	    RECT 1071.9000 1182.7500 1073.7001 1182.9000 ;
	    RECT 1105.5000 1182.7500 1107.3000 1182.9000 ;
	    RECT 1507.2001 1182.7500 1510.5000 1182.9000 ;
	    RECT 1071.9000 1181.2500 1107.3000 1182.7500 ;
	    RECT 1071.9000 1181.1000 1073.7001 1181.2500 ;
	    RECT 1105.5000 1181.1000 1107.3000 1181.2500 ;
	    RECT 1506.4501 1181.1000 1510.5000 1182.7500 ;
	    RECT 1547.1000 1182.7500 1548.9000 1182.9000 ;
	    RECT 1556.7001 1182.7500 1558.5000 1182.9000 ;
	    RECT 1547.1000 1181.2500 1558.5000 1182.7500 ;
	    RECT 1547.1000 1181.1000 1548.9000 1181.2500 ;
	    RECT 1556.7001 1181.1000 1558.5000 1181.2500 ;
	    RECT 111.9000 1176.7500 113.7000 1176.9000 ;
	    RECT 119.1000 1176.7500 120.9000 1176.9000 ;
	    RECT 111.9000 1175.2500 120.9000 1176.7500 ;
	    RECT 111.9000 1175.1000 113.7000 1175.2500 ;
	    RECT 119.1000 1175.1000 120.9000 1175.2500 ;
	    RECT 150.3000 1176.7500 152.1000 1176.9000 ;
	    RECT 171.9000 1176.7500 173.7000 1176.9000 ;
	    RECT 150.3000 1175.2500 173.7000 1176.7500 ;
	    RECT 150.3000 1175.1000 152.1000 1175.2500 ;
	    RECT 171.9000 1175.1000 173.7000 1175.2500 ;
	    RECT 193.5000 1176.7500 195.3000 1176.9000 ;
	    RECT 275.1000 1176.7500 276.9000 1176.9000 ;
	    RECT 193.5000 1175.2500 276.9000 1176.7500 ;
	    RECT 193.5000 1175.1000 195.3000 1175.2500 ;
	    RECT 275.1000 1175.1000 276.9000 1175.2500 ;
	    RECT 344.7000 1176.7500 346.5000 1176.9000 ;
	    RECT 467.1000 1176.7500 468.9000 1176.9000 ;
	    RECT 344.7000 1175.2500 468.9000 1176.7500 ;
	    RECT 344.7000 1175.1000 346.5000 1175.2500 ;
	    RECT 467.1000 1175.1000 468.9000 1175.2500 ;
	    RECT 798.3000 1176.7500 800.1000 1176.9000 ;
	    RECT 812.7000 1176.7500 814.5000 1176.9000 ;
	    RECT 798.3000 1175.2500 814.5000 1176.7500 ;
	    RECT 798.3000 1175.1000 800.1000 1175.2500 ;
	    RECT 812.7000 1175.1000 814.5000 1175.2500 ;
	    RECT 870.3000 1176.7500 872.1000 1176.9000 ;
	    RECT 899.1000 1176.7500 900.9000 1176.9000 ;
	    RECT 870.3000 1175.2500 900.9000 1176.7500 ;
	    RECT 870.3000 1175.1000 872.1000 1175.2500 ;
	    RECT 899.1000 1175.1000 900.9000 1175.2500 ;
	    RECT 983.1000 1176.7500 984.9000 1176.9000 ;
	    RECT 1009.5000 1176.7500 1011.3000 1176.9000 ;
	    RECT 983.1000 1175.2500 1011.3000 1176.7500 ;
	    RECT 983.1000 1175.1000 984.9000 1175.2500 ;
	    RECT 1009.5000 1175.1000 1011.3000 1175.2500 ;
	    RECT 1083.9000 1176.7500 1085.7001 1176.9000 ;
	    RECT 1134.3000 1176.7500 1136.1000 1176.9000 ;
	    RECT 1196.7001 1176.7500 1198.5000 1176.9000 ;
	    RECT 1083.9000 1175.2500 1198.5000 1176.7500 ;
	    RECT 1083.9000 1175.1000 1085.7001 1175.2500 ;
	    RECT 1134.3000 1175.1000 1136.1000 1175.2500 ;
	    RECT 1196.7001 1175.1000 1198.5000 1175.2500 ;
	    RECT 1290.3000 1176.7500 1292.1000 1176.9000 ;
	    RECT 1314.3000 1176.7500 1316.1000 1176.9000 ;
	    RECT 1343.1000 1176.7500 1344.9000 1176.9000 ;
	    RECT 1290.3000 1175.2500 1344.9000 1176.7500 ;
	    RECT 1290.3000 1175.1000 1292.1000 1175.2500 ;
	    RECT 1314.3000 1175.1000 1316.1000 1175.2500 ;
	    RECT 1343.1000 1175.1000 1344.9000 1175.2500 ;
	    RECT 1460.7001 1176.7500 1462.5000 1176.9000 ;
	    RECT 1460.7001 1175.2500 1503.1500 1176.7500 ;
	    RECT 1460.7001 1175.1000 1462.5000 1175.2500 ;
	    RECT 1501.6500 1173.9000 1503.1500 1175.2500 ;
	    RECT 1506.4501 1173.9000 1507.9501 1181.1000 ;
	    RECT 1513.5000 1176.7500 1515.3000 1176.9000 ;
	    RECT 1523.1000 1176.7500 1524.9000 1176.9000 ;
	    RECT 1513.5000 1175.2500 1524.9000 1176.7500 ;
	    RECT 1513.5000 1175.1000 1515.3000 1175.2500 ;
	    RECT 1523.1000 1175.1000 1524.9000 1175.2500 ;
	    RECT 1532.7001 1176.7500 1534.5000 1176.9000 ;
	    RECT 1539.9000 1176.7500 1541.7001 1176.9000 ;
	    RECT 1532.7001 1175.2500 1541.7001 1176.7500 ;
	    RECT 1532.7001 1175.1000 1534.5000 1175.2500 ;
	    RECT 1539.9000 1175.1000 1541.7001 1175.2500 ;
	    RECT 1501.5000 1172.1000 1503.3000 1173.9000 ;
	    RECT 1506.3000 1172.1000 1508.1000 1173.9000 ;
	    RECT 71.1000 1170.7500 72.9000 1170.9000 ;
	    RECT 150.3000 1170.7500 152.1000 1170.9000 ;
	    RECT 71.1000 1169.2500 152.1000 1170.7500 ;
	    RECT 71.1000 1169.1000 72.9000 1169.2500 ;
	    RECT 150.3000 1169.1000 152.1000 1169.2500 ;
	    RECT 323.1000 1170.7500 324.9000 1170.9000 ;
	    RECT 407.1000 1170.7500 408.9000 1170.9000 ;
	    RECT 323.1000 1169.2500 408.9000 1170.7500 ;
	    RECT 323.1000 1169.1000 324.9000 1169.2500 ;
	    RECT 407.1000 1169.1000 408.9000 1169.2500 ;
	    RECT 462.3000 1170.7500 464.1000 1170.9000 ;
	    RECT 486.3000 1170.7500 488.1000 1170.9000 ;
	    RECT 462.3000 1169.2500 488.1000 1170.7500 ;
	    RECT 462.3000 1169.1000 464.1000 1169.2500 ;
	    RECT 486.3000 1169.1000 488.1000 1169.2500 ;
	    RECT 563.1000 1170.7500 564.9000 1170.9000 ;
	    RECT 615.9000 1170.7500 617.7000 1170.9000 ;
	    RECT 563.1000 1169.2500 617.7000 1170.7500 ;
	    RECT 563.1000 1169.1000 564.9000 1169.2500 ;
	    RECT 615.9000 1169.1000 617.7000 1169.2500 ;
	    RECT 848.7000 1170.7500 850.5000 1170.9000 ;
	    RECT 889.5000 1170.7500 891.3000 1170.9000 ;
	    RECT 848.7000 1169.2500 891.3000 1170.7500 ;
	    RECT 848.7000 1169.1000 850.5000 1169.2500 ;
	    RECT 889.5000 1169.1000 891.3000 1169.2500 ;
	    RECT 911.1000 1170.7500 912.9000 1170.9000 ;
	    RECT 1122.3000 1170.7500 1124.1000 1170.9000 ;
	    RECT 911.1000 1169.2500 1124.1000 1170.7500 ;
	    RECT 911.1000 1169.1000 912.9000 1169.2500 ;
	    RECT 1122.3000 1169.1000 1124.1000 1169.2500 ;
	    RECT 1155.9000 1170.7500 1157.7001 1170.9000 ;
	    RECT 1287.9000 1170.7500 1289.7001 1170.9000 ;
	    RECT 1155.9000 1169.2500 1289.7001 1170.7500 ;
	    RECT 1155.9000 1169.1000 1157.7001 1169.2500 ;
	    RECT 1287.9000 1169.1000 1289.7001 1169.2500 ;
	    RECT 1295.1000 1170.7500 1296.9000 1170.9000 ;
	    RECT 1347.9000 1170.7500 1349.7001 1170.9000 ;
	    RECT 1295.1000 1169.2500 1349.7001 1170.7500 ;
	    RECT 1295.1000 1169.1000 1296.9000 1169.2500 ;
	    RECT 1347.9000 1169.1000 1349.7001 1169.2500 ;
	    RECT 1503.9000 1170.7500 1505.7001 1170.9000 ;
	    RECT 1508.7001 1170.7500 1510.5000 1170.9000 ;
	    RECT 1513.5000 1170.7500 1515.3000 1170.9000 ;
	    RECT 1503.9000 1169.2500 1515.3000 1170.7500 ;
	    RECT 1503.9000 1169.1000 1505.7001 1169.2500 ;
	    RECT 1508.7001 1169.1000 1510.5000 1169.2500 ;
	    RECT 1513.5000 1169.1000 1515.3000 1169.2500 ;
	    RECT 150.3000 1164.7500 152.1000 1164.9000 ;
	    RECT 167.1000 1164.7500 168.9000 1164.9000 ;
	    RECT 150.3000 1163.2500 168.9000 1164.7500 ;
	    RECT 150.3000 1163.1000 152.1000 1163.2500 ;
	    RECT 167.1000 1163.1000 168.9000 1163.2500 ;
	    RECT 253.5000 1164.7500 255.3000 1164.9000 ;
	    RECT 277.5000 1164.7500 279.3000 1164.9000 ;
	    RECT 253.5000 1163.2500 279.3000 1164.7500 ;
	    RECT 253.5000 1163.1000 255.3000 1163.2500 ;
	    RECT 277.5000 1163.1000 279.3000 1163.2500 ;
	    RECT 527.1000 1164.7500 528.9000 1164.9000 ;
	    RECT 584.7000 1164.7500 586.5000 1164.9000 ;
	    RECT 527.1000 1163.2500 586.5000 1164.7500 ;
	    RECT 527.1000 1163.1000 528.9000 1163.2500 ;
	    RECT 584.7000 1163.1000 586.5000 1163.2500 ;
	    RECT 807.9000 1164.7500 809.7000 1164.9000 ;
	    RECT 819.9000 1164.7500 821.7000 1164.9000 ;
	    RECT 839.1000 1164.7500 840.9000 1164.9000 ;
	    RECT 875.1000 1164.7500 876.9000 1164.9000 ;
	    RECT 807.9000 1163.2500 876.9000 1164.7500 ;
	    RECT 807.9000 1163.1000 809.7000 1163.2500 ;
	    RECT 819.9000 1163.1000 821.7000 1163.2500 ;
	    RECT 839.1000 1163.1000 840.9000 1163.2500 ;
	    RECT 875.1000 1163.1000 876.9000 1163.2500 ;
	    RECT 891.9000 1164.7500 893.7000 1164.9000 ;
	    RECT 973.5000 1164.7500 975.3000 1164.9000 ;
	    RECT 891.9000 1163.2500 975.3000 1164.7500 ;
	    RECT 891.9000 1163.1000 893.7000 1163.2500 ;
	    RECT 973.5000 1163.1000 975.3000 1163.2500 ;
	    RECT 1086.3000 1164.7500 1088.1000 1164.9000 ;
	    RECT 1119.9000 1164.7500 1121.7001 1164.9000 ;
	    RECT 1086.3000 1163.2500 1121.7001 1164.7500 ;
	    RECT 1086.3000 1163.1000 1088.1000 1163.2500 ;
	    RECT 1119.9000 1163.1000 1121.7001 1163.2500 ;
	    RECT 1343.1000 1164.7500 1344.9000 1164.9000 ;
	    RECT 1460.7001 1164.7500 1462.5000 1164.9000 ;
	    RECT 1343.1000 1163.2500 1462.5000 1164.7500 ;
	    RECT 1343.1000 1163.1000 1344.9000 1163.2500 ;
	    RECT 1460.7001 1163.1000 1462.5000 1163.2500 ;
	    RECT 1494.3000 1164.7500 1496.1000 1164.9000 ;
	    RECT 1518.3000 1164.7500 1520.1000 1164.9000 ;
	    RECT 1494.3000 1163.2500 1520.1000 1164.7500 ;
	    RECT 1494.3000 1163.1000 1496.1000 1163.2500 ;
	    RECT 1518.3000 1163.1000 1520.1000 1163.2500 ;
	    RECT 222.3000 1158.7500 224.1000 1158.9000 ;
	    RECT 253.5000 1158.7500 255.3000 1158.9000 ;
	    RECT 222.3000 1157.2500 255.3000 1158.7500 ;
	    RECT 222.3000 1157.1000 224.1000 1157.2500 ;
	    RECT 253.5000 1157.1000 255.3000 1157.2500 ;
	    RECT 265.5000 1158.7500 267.3000 1158.9000 ;
	    RECT 378.3000 1158.7500 380.1000 1158.9000 ;
	    RECT 265.5000 1157.2500 380.1000 1158.7500 ;
	    RECT 265.5000 1157.1000 267.3000 1157.2500 ;
	    RECT 378.3000 1157.1000 380.1000 1157.2500 ;
	    RECT 565.5000 1158.7500 567.3000 1158.9000 ;
	    RECT 589.5000 1158.7500 591.3000 1158.9000 ;
	    RECT 565.5000 1157.2500 591.3000 1158.7500 ;
	    RECT 565.5000 1157.1000 567.3000 1157.2500 ;
	    RECT 589.5000 1157.1000 591.3000 1157.2500 ;
	    RECT 611.1000 1158.7500 612.9000 1158.9000 ;
	    RECT 623.1000 1158.7500 624.9000 1158.9000 ;
	    RECT 611.1000 1157.2500 624.9000 1158.7500 ;
	    RECT 611.1000 1157.1000 612.9000 1157.2500 ;
	    RECT 623.1000 1157.1000 624.9000 1157.2500 ;
	    RECT 1182.3000 1158.7500 1184.1000 1158.9000 ;
	    RECT 1189.5000 1158.7500 1191.3000 1158.9000 ;
	    RECT 1182.3000 1157.2500 1191.3000 1158.7500 ;
	    RECT 1182.3000 1157.1000 1184.1000 1157.2500 ;
	    RECT 1189.5000 1157.1000 1191.3000 1157.2500 ;
	    RECT 1304.7001 1158.7500 1306.5000 1158.9000 ;
	    RECT 1357.5000 1158.7500 1359.3000 1158.9000 ;
	    RECT 1304.7001 1157.2500 1359.3000 1158.7500 ;
	    RECT 1304.7001 1157.1000 1306.5000 1157.2500 ;
	    RECT 1357.5000 1157.1000 1359.3000 1157.2500 ;
	    RECT 1489.5000 1158.7500 1491.3000 1158.9000 ;
	    RECT 1508.7001 1158.7500 1510.5000 1158.9000 ;
	    RECT 1489.5000 1157.2500 1510.5000 1158.7500 ;
	    RECT 1489.5000 1157.1000 1491.3000 1157.2500 ;
	    RECT 1508.7001 1157.1000 1510.5000 1157.2500 ;
	    RECT 13.5000 1152.7500 15.3000 1152.9000 ;
	    RECT 85.5000 1152.7500 87.3000 1152.9000 ;
	    RECT 114.3000 1152.7500 116.1000 1152.9000 ;
	    RECT 13.5000 1151.2500 116.1000 1152.7500 ;
	    RECT 13.5000 1151.1000 15.3000 1151.2500 ;
	    RECT 85.5000 1151.1000 87.3000 1151.2500 ;
	    RECT 114.3000 1151.1000 116.1000 1151.2500 ;
	    RECT 181.5000 1152.7500 183.3000 1152.9000 ;
	    RECT 265.5000 1152.7500 267.3000 1152.9000 ;
	    RECT 181.5000 1151.2500 267.3000 1152.7500 ;
	    RECT 181.5000 1151.1000 183.3000 1151.2500 ;
	    RECT 265.5000 1151.1000 267.3000 1151.2500 ;
	    RECT 272.7000 1152.7500 274.5000 1152.9000 ;
	    RECT 287.1000 1152.7500 288.9000 1152.9000 ;
	    RECT 303.9000 1152.7500 305.7000 1152.9000 ;
	    RECT 272.7000 1151.2500 305.7000 1152.7500 ;
	    RECT 272.7000 1151.1000 274.5000 1151.2500 ;
	    RECT 287.1000 1151.1000 288.9000 1151.2500 ;
	    RECT 303.9000 1151.1000 305.7000 1151.2500 ;
	    RECT 459.9000 1152.7500 461.7000 1152.9000 ;
	    RECT 491.1000 1152.7500 492.9000 1152.9000 ;
	    RECT 459.9000 1151.2500 492.9000 1152.7500 ;
	    RECT 459.9000 1151.1000 461.7000 1151.2500 ;
	    RECT 491.1000 1151.1000 492.9000 1151.2500 ;
	    RECT 582.3000 1152.7500 584.1000 1152.9000 ;
	    RECT 709.5000 1152.7500 711.3000 1152.9000 ;
	    RECT 582.3000 1151.2500 711.3000 1152.7500 ;
	    RECT 582.3000 1151.1000 584.1000 1151.2500 ;
	    RECT 709.5000 1151.1000 711.3000 1151.2500 ;
	    RECT 743.1000 1152.7500 744.9000 1152.9000 ;
	    RECT 1098.3000 1152.7500 1100.1000 1152.9000 ;
	    RECT 743.1000 1151.2500 1100.1000 1152.7500 ;
	    RECT 743.1000 1151.1000 744.9000 1151.2500 ;
	    RECT 1098.3000 1151.1000 1100.1000 1151.2500 ;
	    RECT 1184.7001 1152.7500 1186.5000 1152.9000 ;
	    RECT 1347.9000 1152.7500 1349.7001 1152.9000 ;
	    RECT 1184.7001 1151.2500 1349.7001 1152.7500 ;
	    RECT 1184.7001 1151.1000 1186.5000 1151.2500 ;
	    RECT 1347.9000 1151.1000 1349.7001 1151.2500 ;
	    RECT 188.7000 1146.7500 190.5000 1146.9000 ;
	    RECT 258.3000 1146.7500 260.1000 1146.9000 ;
	    RECT 188.7000 1145.2500 260.1000 1146.7500 ;
	    RECT 188.7000 1145.1000 190.5000 1145.2500 ;
	    RECT 258.3000 1145.1000 260.1000 1145.2500 ;
	    RECT 289.5000 1146.7500 291.3000 1146.9000 ;
	    RECT 431.1000 1146.7500 432.9000 1146.9000 ;
	    RECT 455.1000 1146.7500 456.9000 1146.9000 ;
	    RECT 289.5000 1145.2500 456.9000 1146.7500 ;
	    RECT 289.5000 1145.1000 291.3000 1145.2500 ;
	    RECT 431.1000 1145.1000 432.9000 1145.2500 ;
	    RECT 455.1000 1145.1000 456.9000 1145.2500 ;
	    RECT 551.1000 1146.7500 552.9000 1146.9000 ;
	    RECT 589.5000 1146.7500 591.3000 1146.9000 ;
	    RECT 683.1000 1146.7500 684.9000 1146.9000 ;
	    RECT 551.1000 1145.2500 684.9000 1146.7500 ;
	    RECT 551.1000 1145.1000 552.9000 1145.2500 ;
	    RECT 589.5000 1145.1000 591.3000 1145.2500 ;
	    RECT 683.1000 1145.1000 684.9000 1145.2500 ;
	    RECT 745.5000 1146.7500 747.3000 1146.9000 ;
	    RECT 767.1000 1146.7500 768.9000 1146.9000 ;
	    RECT 745.5000 1145.2500 768.9000 1146.7500 ;
	    RECT 745.5000 1145.1000 747.3000 1145.2500 ;
	    RECT 767.1000 1145.1000 768.9000 1145.2500 ;
	    RECT 908.7000 1146.7500 910.5000 1146.9000 ;
	    RECT 968.7000 1146.7500 970.5000 1146.9000 ;
	    RECT 908.7000 1145.2500 970.5000 1146.7500 ;
	    RECT 908.7000 1145.1000 910.5000 1145.2500 ;
	    RECT 968.7000 1145.1000 970.5000 1145.2500 ;
	    RECT 997.5000 1146.7500 999.3000 1146.9000 ;
	    RECT 1057.5000 1146.7500 1059.3000 1146.9000 ;
	    RECT 997.5000 1145.2500 1059.3000 1146.7500 ;
	    RECT 997.5000 1145.1000 999.3000 1145.2500 ;
	    RECT 1057.5000 1145.1000 1059.3000 1145.2500 ;
	    RECT 1069.5000 1146.7500 1071.3000 1146.9000 ;
	    RECT 1093.5000 1146.7500 1095.3000 1146.9000 ;
	    RECT 1069.5000 1145.2500 1095.3000 1146.7500 ;
	    RECT 1069.5000 1145.1000 1071.3000 1145.2500 ;
	    RECT 1093.5000 1145.1000 1095.3000 1145.2500 ;
	    RECT 155.1000 1140.7500 156.9000 1140.9000 ;
	    RECT 164.7000 1140.7500 166.5000 1140.9000 ;
	    RECT 155.1000 1139.2500 166.5000 1140.7500 ;
	    RECT 155.1000 1139.1000 156.9000 1139.2500 ;
	    RECT 164.7000 1139.1000 166.5000 1139.2500 ;
	    RECT 229.5000 1140.7500 231.3000 1140.9000 ;
	    RECT 255.9000 1140.7500 257.7000 1140.9000 ;
	    RECT 229.5000 1139.2500 257.7000 1140.7500 ;
	    RECT 229.5000 1139.1000 231.3000 1139.2500 ;
	    RECT 255.9000 1139.1000 257.7000 1139.2500 ;
	    RECT 277.5000 1140.7500 279.3000 1140.9000 ;
	    RECT 311.1000 1140.7500 312.9000 1140.9000 ;
	    RECT 277.5000 1139.2500 312.9000 1140.7500 ;
	    RECT 277.5000 1139.1000 279.3000 1139.2500 ;
	    RECT 311.1000 1139.1000 312.9000 1139.2500 ;
	    RECT 378.3000 1140.7500 380.1000 1140.9000 ;
	    RECT 500.7000 1140.7500 502.5000 1140.9000 ;
	    RECT 378.3000 1139.2500 502.5000 1140.7500 ;
	    RECT 378.3000 1139.1000 380.1000 1139.2500 ;
	    RECT 500.7000 1139.1000 502.5000 1139.2500 ;
	    RECT 767.1000 1140.7500 768.9000 1140.9000 ;
	    RECT 781.5000 1140.7500 783.3000 1140.9000 ;
	    RECT 767.1000 1139.2500 783.3000 1140.7500 ;
	    RECT 767.1000 1139.1000 768.9000 1139.2500 ;
	    RECT 781.5000 1139.1000 783.3000 1139.2500 ;
	    RECT 851.1000 1140.7500 852.9000 1140.9000 ;
	    RECT 867.9000 1140.7500 869.7000 1140.9000 ;
	    RECT 851.1000 1139.2500 869.7000 1140.7500 ;
	    RECT 851.1000 1139.1000 852.9000 1139.2500 ;
	    RECT 867.9000 1139.1000 869.7000 1139.2500 ;
	    RECT 932.7000 1140.7500 934.5000 1140.9000 ;
	    RECT 1004.7000 1140.7500 1006.5000 1140.9000 ;
	    RECT 932.7000 1139.2500 1006.5000 1140.7500 ;
	    RECT 932.7000 1139.1000 934.5000 1139.2500 ;
	    RECT 1004.7000 1139.1000 1006.5000 1139.2500 ;
	    RECT 1091.1000 1140.7500 1092.9000 1140.9000 ;
	    RECT 1110.3000 1140.7500 1112.1000 1140.9000 ;
	    RECT 1091.1000 1139.2500 1112.1000 1140.7500 ;
	    RECT 1091.1000 1139.1000 1092.9000 1139.2500 ;
	    RECT 1110.3000 1139.1000 1112.1000 1139.2500 ;
	    RECT 1362.3000 1140.7500 1364.1000 1140.9000 ;
	    RECT 1412.7001 1140.7500 1414.5000 1140.9000 ;
	    RECT 1362.3000 1139.2500 1414.5000 1140.7500 ;
	    RECT 1362.3000 1139.1000 1364.1000 1139.2500 ;
	    RECT 1412.7001 1139.1000 1414.5000 1139.2500 ;
	    RECT 1523.1000 1140.7500 1524.9000 1140.9000 ;
	    RECT 1527.9000 1140.7500 1529.7001 1140.9000 ;
	    RECT 1523.1000 1139.2500 1529.7001 1140.7500 ;
	    RECT 1523.1000 1139.1000 1524.9000 1139.2500 ;
	    RECT 1527.9000 1139.1000 1529.7001 1139.2500 ;
	    RECT 23.1000 1134.7500 24.9000 1134.9000 ;
	    RECT 126.3000 1134.7500 128.1000 1134.9000 ;
	    RECT 23.1000 1133.2500 128.1000 1134.7500 ;
	    RECT 23.1000 1133.1000 24.9000 1133.2500 ;
	    RECT 126.3000 1133.1000 128.1000 1133.2500 ;
	    RECT 443.1000 1134.7500 444.9000 1134.9000 ;
	    RECT 452.7000 1134.7500 454.5000 1134.9000 ;
	    RECT 479.1000 1134.7500 480.9000 1134.9000 ;
	    RECT 443.1000 1133.2500 480.9000 1134.7500 ;
	    RECT 443.1000 1133.1000 444.9000 1133.2500 ;
	    RECT 452.7000 1133.1000 454.5000 1133.2500 ;
	    RECT 479.1000 1133.1000 480.9000 1133.2500 ;
	    RECT 656.7000 1134.7500 658.5000 1134.9000 ;
	    RECT 668.7000 1134.7500 670.5000 1134.9000 ;
	    RECT 863.1000 1134.7500 864.9000 1134.9000 ;
	    RECT 656.7000 1133.2500 864.9000 1134.7500 ;
	    RECT 656.7000 1133.1000 658.5000 1133.2500 ;
	    RECT 668.7000 1133.1000 670.5000 1133.2500 ;
	    RECT 863.1000 1133.1000 864.9000 1133.2500 ;
	    RECT 913.5000 1134.7500 915.3000 1134.9000 ;
	    RECT 1002.3000 1134.7500 1004.1000 1134.9000 ;
	    RECT 913.5000 1133.2500 1004.1000 1134.7500 ;
	    RECT 913.5000 1133.1000 915.3000 1133.2500 ;
	    RECT 1002.3000 1133.1000 1004.1000 1133.2500 ;
	    RECT 1014.3000 1134.7500 1016.1000 1134.9000 ;
	    RECT 1028.7001 1134.7500 1030.5000 1134.9000 ;
	    RECT 1040.7001 1134.7500 1042.5000 1134.9000 ;
	    RECT 1014.3000 1133.2500 1042.5000 1134.7500 ;
	    RECT 1014.3000 1133.1000 1016.1000 1133.2500 ;
	    RECT 1028.7001 1133.1000 1030.5000 1133.2500 ;
	    RECT 1040.7001 1133.1000 1042.5000 1133.2500 ;
	    RECT 1412.7001 1134.7500 1414.5000 1134.9000 ;
	    RECT 1443.9000 1134.7500 1445.7001 1134.9000 ;
	    RECT 1412.7001 1133.2500 1445.7001 1134.7500 ;
	    RECT 1412.7001 1133.1000 1414.5000 1133.2500 ;
	    RECT 1443.9000 1133.1000 1445.7001 1133.2500 ;
	    RECT 126.3000 1128.7500 128.1000 1128.9000 ;
	    RECT 131.1000 1128.7500 132.9000 1128.9000 ;
	    RECT 126.3000 1127.2500 132.9000 1128.7500 ;
	    RECT 126.3000 1127.1000 128.1000 1127.2500 ;
	    RECT 131.1000 1127.1000 132.9000 1127.2500 ;
	    RECT 181.5000 1128.7500 183.3000 1128.9000 ;
	    RECT 193.5000 1128.7500 195.3000 1128.9000 ;
	    RECT 181.5000 1127.2500 195.3000 1128.7500 ;
	    RECT 181.5000 1127.1000 183.3000 1127.2500 ;
	    RECT 193.5000 1127.1000 195.3000 1127.2500 ;
	    RECT 299.1000 1128.7500 300.9000 1128.9000 ;
	    RECT 303.9000 1128.7500 305.7000 1128.9000 ;
	    RECT 299.1000 1127.2500 305.7000 1128.7500 ;
	    RECT 299.1000 1127.1000 300.9000 1127.2500 ;
	    RECT 303.9000 1127.1000 305.7000 1127.2500 ;
	    RECT 500.7000 1128.7500 502.5000 1128.9000 ;
	    RECT 507.9000 1128.7500 509.7000 1128.9000 ;
	    RECT 500.7000 1127.2500 509.7000 1128.7500 ;
	    RECT 500.7000 1127.1000 502.5000 1127.2500 ;
	    RECT 507.9000 1127.1000 509.7000 1127.2500 ;
	    RECT 656.7000 1128.7500 658.5000 1128.9000 ;
	    RECT 702.3000 1128.7500 704.1000 1128.9000 ;
	    RECT 656.7000 1127.2500 704.1000 1128.7500 ;
	    RECT 656.7000 1127.1000 658.5000 1127.2500 ;
	    RECT 702.3000 1127.1000 704.1000 1127.2500 ;
	    RECT 1023.9000 1128.7500 1025.7001 1128.9000 ;
	    RECT 1045.5000 1128.7500 1047.3000 1128.9000 ;
	    RECT 1023.9000 1127.2500 1047.3000 1128.7500 ;
	    RECT 1023.9000 1127.1000 1025.7001 1127.2500 ;
	    RECT 1045.5000 1127.1000 1047.3000 1127.2500 ;
	    RECT 1052.7001 1128.7500 1054.5000 1128.9000 ;
	    RECT 1093.5000 1128.7500 1095.3000 1128.9000 ;
	    RECT 1052.7001 1127.2500 1095.3000 1128.7500 ;
	    RECT 1052.7001 1127.1000 1054.5000 1127.2500 ;
	    RECT 1093.5000 1127.1000 1095.3000 1127.2500 ;
	    RECT 1215.9000 1128.7500 1217.7001 1128.9000 ;
	    RECT 1309.5000 1128.7500 1311.3000 1128.9000 ;
	    RECT 1215.9000 1127.2500 1311.3000 1128.7500 ;
	    RECT 1215.9000 1127.1000 1217.7001 1127.2500 ;
	    RECT 1309.5000 1127.1000 1311.3000 1127.2500 ;
	    RECT 1501.5000 1128.7500 1503.3000 1128.9000 ;
	    RECT 1525.5000 1128.7500 1527.3000 1128.9000 ;
	    RECT 1501.5000 1127.2500 1527.3000 1128.7500 ;
	    RECT 1501.5000 1127.1000 1503.3000 1127.2500 ;
	    RECT 1525.5000 1127.1000 1527.3000 1127.2500 ;
	    RECT 131.1000 1122.7500 132.9000 1122.9000 ;
	    RECT 176.7000 1122.7500 178.5000 1122.9000 ;
	    RECT 131.1000 1121.2500 178.5000 1122.7500 ;
	    RECT 131.1000 1121.1000 132.9000 1121.2500 ;
	    RECT 176.7000 1121.1000 178.5000 1121.2500 ;
	    RECT 222.3000 1122.7500 224.1000 1122.9000 ;
	    RECT 231.9000 1122.7500 233.7000 1122.9000 ;
	    RECT 222.3000 1121.2500 233.7000 1122.7500 ;
	    RECT 222.3000 1121.1000 224.1000 1121.2500 ;
	    RECT 231.9000 1121.1000 233.7000 1121.2500 ;
	    RECT 270.3000 1122.7500 272.1000 1122.9000 ;
	    RECT 301.5000 1122.7500 303.3000 1122.9000 ;
	    RECT 270.3000 1121.2500 303.3000 1122.7500 ;
	    RECT 270.3000 1121.1000 272.1000 1121.2500 ;
	    RECT 301.5000 1121.1000 303.3000 1121.2500 ;
	    RECT 327.9000 1122.7500 329.7000 1122.9000 ;
	    RECT 335.1000 1122.7500 336.9000 1122.9000 ;
	    RECT 327.9000 1121.2500 336.9000 1122.7500 ;
	    RECT 327.9000 1121.1000 329.7000 1121.2500 ;
	    RECT 335.1000 1121.1000 336.9000 1121.2500 ;
	    RECT 390.3000 1122.7500 392.1000 1122.9000 ;
	    RECT 459.9000 1122.7500 461.7000 1122.9000 ;
	    RECT 390.3000 1121.2500 461.7000 1122.7500 ;
	    RECT 390.3000 1121.1000 392.1000 1121.2500 ;
	    RECT 459.9000 1121.1000 461.7000 1121.2500 ;
	    RECT 680.7000 1122.7500 682.5000 1122.9000 ;
	    RECT 711.9000 1122.7500 713.7000 1122.9000 ;
	    RECT 680.7000 1121.2500 713.7000 1122.7500 ;
	    RECT 680.7000 1121.1000 682.5000 1121.2500 ;
	    RECT 711.9000 1121.1000 713.7000 1121.2500 ;
	    RECT 716.7000 1122.7500 718.5000 1122.9000 ;
	    RECT 723.9000 1122.7500 725.7000 1122.9000 ;
	    RECT 716.7000 1121.2500 725.7000 1122.7500 ;
	    RECT 716.7000 1121.1000 718.5000 1121.2500 ;
	    RECT 723.9000 1121.1000 725.7000 1121.2500 ;
	    RECT 781.5000 1122.7500 783.3000 1122.9000 ;
	    RECT 800.7000 1122.7500 802.5000 1122.9000 ;
	    RECT 781.5000 1121.2500 802.5000 1122.7500 ;
	    RECT 781.5000 1121.1000 783.3000 1121.2500 ;
	    RECT 800.7000 1121.1000 802.5000 1121.2500 ;
	    RECT 1007.1000 1122.7500 1008.9000 1122.9000 ;
	    RECT 1083.9000 1122.7500 1085.7001 1122.9000 ;
	    RECT 1227.9000 1122.7500 1229.7001 1122.9000 ;
	    RECT 1007.1000 1121.2500 1229.7001 1122.7500 ;
	    RECT 1007.1000 1121.1000 1008.9000 1121.2500 ;
	    RECT 1083.9000 1121.1000 1085.7001 1121.2500 ;
	    RECT 1227.9000 1121.1000 1229.7001 1121.2500 ;
	    RECT 1237.5000 1122.7500 1239.3000 1122.9000 ;
	    RECT 1285.5000 1122.7500 1287.3000 1122.9000 ;
	    RECT 1237.5000 1121.2500 1287.3000 1122.7500 ;
	    RECT 1237.5000 1121.1000 1239.3000 1121.2500 ;
	    RECT 1285.5000 1121.1000 1287.3000 1121.2500 ;
	    RECT 1307.1000 1122.7500 1308.9000 1122.9000 ;
	    RECT 1314.3000 1122.7500 1316.1000 1122.9000 ;
	    RECT 1307.1000 1121.2500 1316.1000 1122.7500 ;
	    RECT 1307.1000 1121.1000 1308.9000 1121.2500 ;
	    RECT 1314.3000 1121.1000 1316.1000 1121.2500 ;
	    RECT 1383.9000 1122.7500 1385.7001 1122.9000 ;
	    RECT 1391.1000 1122.7500 1392.9000 1122.9000 ;
	    RECT 1383.9000 1121.2500 1392.9000 1122.7500 ;
	    RECT 1383.9000 1121.1000 1385.7001 1121.2500 ;
	    RECT 1391.1000 1121.1000 1392.9000 1121.2500 ;
	    RECT 155.1000 1116.7500 156.9000 1116.9000 ;
	    RECT 229.5000 1116.7500 231.3000 1116.9000 ;
	    RECT 155.1000 1115.2500 231.3000 1116.7500 ;
	    RECT 155.1000 1115.1000 156.9000 1115.2500 ;
	    RECT 229.5000 1115.1000 231.3000 1115.2500 ;
	    RECT 243.9000 1116.7500 245.7000 1116.9000 ;
	    RECT 248.7000 1116.7500 250.5000 1116.9000 ;
	    RECT 243.9000 1115.2500 250.5000 1116.7500 ;
	    RECT 243.9000 1115.1000 245.7000 1115.2500 ;
	    RECT 248.7000 1115.1000 250.5000 1115.2500 ;
	    RECT 375.9000 1116.7500 377.7000 1116.9000 ;
	    RECT 416.7000 1116.7500 418.5000 1116.9000 ;
	    RECT 445.5000 1116.7500 447.3000 1116.9000 ;
	    RECT 615.9000 1116.7500 617.7000 1116.9000 ;
	    RECT 375.9000 1115.2500 617.7000 1116.7500 ;
	    RECT 375.9000 1115.1000 377.7000 1115.2500 ;
	    RECT 416.7000 1115.1000 418.5000 1115.2500 ;
	    RECT 445.5000 1115.1000 447.3000 1115.2500 ;
	    RECT 615.9000 1115.1000 617.7000 1115.2500 ;
	    RECT 877.5000 1116.7500 879.3000 1116.9000 ;
	    RECT 923.1000 1116.7500 924.9000 1116.9000 ;
	    RECT 877.5000 1115.2500 924.9000 1116.7500 ;
	    RECT 877.5000 1115.1000 879.3000 1115.2500 ;
	    RECT 923.1000 1115.1000 924.9000 1115.2500 ;
	    RECT 944.7000 1116.7500 946.5000 1116.9000 ;
	    RECT 990.3000 1116.7500 992.1000 1116.9000 ;
	    RECT 1071.9000 1116.7500 1073.7001 1116.9000 ;
	    RECT 944.7000 1115.2500 1073.7001 1116.7500 ;
	    RECT 944.7000 1115.1000 946.5000 1115.2500 ;
	    RECT 990.3000 1115.1000 992.1000 1115.2500 ;
	    RECT 1071.9000 1115.1000 1073.7001 1115.2500 ;
	    RECT 1093.5000 1116.7500 1095.3000 1116.9000 ;
	    RECT 1374.3000 1116.7500 1376.1000 1116.9000 ;
	    RECT 1093.5000 1115.2500 1376.1000 1116.7500 ;
	    RECT 1093.5000 1115.1000 1095.3000 1115.2500 ;
	    RECT 1374.3000 1115.1000 1376.1000 1115.2500 ;
	    RECT 1429.5000 1116.7500 1431.3000 1116.9000 ;
	    RECT 1513.5000 1116.7500 1515.3000 1116.9000 ;
	    RECT 1429.5000 1115.2500 1515.3000 1116.7500 ;
	    RECT 1429.5000 1115.1000 1431.3000 1115.2500 ;
	    RECT 1513.5000 1115.1000 1515.3000 1115.2500 ;
	    RECT 1527.9000 1116.7500 1529.7001 1116.9000 ;
	    RECT 1549.5000 1116.7500 1551.3000 1116.9000 ;
	    RECT 1527.9000 1115.2500 1551.3000 1116.7500 ;
	    RECT 1527.9000 1115.1000 1529.7001 1115.2500 ;
	    RECT 1549.5000 1115.1000 1551.3000 1115.2500 ;
	    RECT 135.9000 1110.7500 137.7000 1110.9000 ;
	    RECT 159.9000 1110.7500 161.7000 1110.9000 ;
	    RECT 135.9000 1109.2500 161.7000 1110.7500 ;
	    RECT 135.9000 1109.1000 137.7000 1109.2500 ;
	    RECT 159.9000 1109.1000 161.7000 1109.2500 ;
	    RECT 246.3000 1110.7500 248.1000 1110.9000 ;
	    RECT 260.7000 1110.7500 262.5000 1110.9000 ;
	    RECT 246.3000 1109.2500 262.5000 1110.7500 ;
	    RECT 246.3000 1109.1000 248.1000 1109.2500 ;
	    RECT 260.7000 1109.1000 262.5000 1109.2500 ;
	    RECT 313.5000 1110.7500 315.3000 1110.9000 ;
	    RECT 337.5000 1110.7500 339.3000 1110.9000 ;
	    RECT 313.5000 1109.2500 339.3000 1110.7500 ;
	    RECT 313.5000 1109.1000 315.3000 1109.2500 ;
	    RECT 337.5000 1109.1000 339.3000 1109.2500 ;
	    RECT 596.7000 1110.7500 600.0000 1110.9000 ;
	    RECT 632.7000 1110.7500 634.5000 1110.9000 ;
	    RECT 707.1000 1110.7500 708.9000 1110.9000 ;
	    RECT 596.7000 1109.1000 600.7500 1110.7500 ;
	    RECT 632.7000 1109.2500 708.9000 1110.7500 ;
	    RECT 632.7000 1109.1000 634.5000 1109.2500 ;
	    RECT 707.1000 1109.1000 708.9000 1109.2500 ;
	    RECT 747.9000 1110.7500 749.7000 1110.9000 ;
	    RECT 791.1000 1110.7500 792.9000 1110.9000 ;
	    RECT 747.9000 1109.2500 792.9000 1110.7500 ;
	    RECT 747.9000 1109.1000 749.7000 1109.2500 ;
	    RECT 791.1000 1109.1000 792.9000 1109.2500 ;
	    RECT 819.9000 1110.7500 821.7000 1110.9000 ;
	    RECT 831.9000 1110.7500 833.7000 1110.9000 ;
	    RECT 819.9000 1109.2500 833.7000 1110.7500 ;
	    RECT 819.9000 1109.1000 821.7000 1109.2500 ;
	    RECT 831.9000 1109.1000 833.7000 1109.2500 ;
	    RECT 918.3000 1110.7500 920.1000 1110.9000 ;
	    RECT 930.3000 1110.7500 932.1000 1110.9000 ;
	    RECT 918.3000 1109.2500 932.1000 1110.7500 ;
	    RECT 918.3000 1109.1000 920.1000 1109.2500 ;
	    RECT 930.3000 1109.1000 932.1000 1109.2500 ;
	    RECT 999.9000 1110.7500 1001.7000 1110.9000 ;
	    RECT 1011.9000 1110.7500 1013.7000 1110.9000 ;
	    RECT 999.9000 1109.2500 1013.7000 1110.7500 ;
	    RECT 999.9000 1109.1000 1001.7000 1109.2500 ;
	    RECT 1011.9000 1109.1000 1013.7000 1109.2500 ;
	    RECT 1019.1000 1110.7500 1020.9000 1110.9000 ;
	    RECT 1112.7001 1110.7500 1114.5000 1110.9000 ;
	    RECT 1019.1000 1109.2500 1114.5000 1110.7500 ;
	    RECT 1019.1000 1109.1000 1020.9000 1109.2500 ;
	    RECT 1112.7001 1109.1000 1114.5000 1109.2500 ;
	    RECT 1218.3000 1110.7500 1220.1000 1110.9000 ;
	    RECT 1242.3000 1110.7500 1244.1000 1110.9000 ;
	    RECT 1218.3000 1109.2500 1244.1000 1110.7500 ;
	    RECT 1218.3000 1109.1000 1220.1000 1109.2500 ;
	    RECT 1242.3000 1109.1000 1244.1000 1109.2500 ;
	    RECT 1297.5000 1110.7500 1299.3000 1110.9000 ;
	    RECT 1319.1000 1110.7500 1320.9000 1110.9000 ;
	    RECT 1297.5000 1109.2500 1320.9000 1110.7500 ;
	    RECT 1297.5000 1109.1000 1299.3000 1109.2500 ;
	    RECT 1319.1000 1109.1000 1320.9000 1109.2500 ;
	    RECT 1405.5000 1110.7500 1407.3000 1110.9000 ;
	    RECT 1429.5000 1110.7500 1431.3000 1110.9000 ;
	    RECT 1405.5000 1109.2500 1431.3000 1110.7500 ;
	    RECT 1405.5000 1109.1000 1407.3000 1109.2500 ;
	    RECT 1429.5000 1109.1000 1431.3000 1109.2500 ;
	    RECT 1494.3000 1110.7500 1496.1000 1110.9000 ;
	    RECT 1559.1000 1110.7500 1560.9000 1110.9000 ;
	    RECT 1494.3000 1109.2500 1560.9000 1110.7500 ;
	    RECT 1494.3000 1109.1000 1496.1000 1109.2500 ;
	    RECT 1559.1000 1109.1000 1560.9000 1109.2500 ;
	    RECT 210.3000 1104.7500 212.1000 1104.9000 ;
	    RECT 231.9000 1104.7500 233.7000 1104.9000 ;
	    RECT 210.3000 1103.2500 233.7000 1104.7500 ;
	    RECT 210.3000 1103.1000 212.1000 1103.2500 ;
	    RECT 231.9000 1103.1000 233.7000 1103.2500 ;
	    RECT 289.5000 1104.7500 291.3000 1104.9000 ;
	    RECT 339.9000 1104.7500 341.7000 1104.9000 ;
	    RECT 289.5000 1103.2500 341.7000 1104.7500 ;
	    RECT 289.5000 1103.1000 291.3000 1103.2500 ;
	    RECT 339.9000 1103.1000 341.7000 1103.2500 ;
	    RECT 541.5000 1104.7500 543.3000 1104.9000 ;
	    RECT 548.7000 1104.7500 550.5000 1104.9000 ;
	    RECT 591.9000 1104.7500 593.7000 1104.9000 ;
	    RECT 541.5000 1103.2500 593.7000 1104.7500 ;
	    RECT 541.5000 1103.1000 543.3000 1103.2500 ;
	    RECT 548.7000 1103.1000 550.5000 1103.2500 ;
	    RECT 591.9000 1103.1000 593.7000 1103.2500 ;
	    RECT 49.5000 1098.7500 51.3000 1098.9000 ;
	    RECT 143.1000 1098.7500 144.9000 1098.9000 ;
	    RECT 49.5000 1097.2500 144.9000 1098.7500 ;
	    RECT 49.5000 1097.1000 51.3000 1097.2500 ;
	    RECT 143.1000 1097.1000 144.9000 1097.2500 ;
	    RECT 164.7000 1098.7500 166.5000 1098.9000 ;
	    RECT 169.5000 1098.7500 171.3000 1098.9000 ;
	    RECT 164.7000 1097.2500 171.3000 1098.7500 ;
	    RECT 164.7000 1097.1000 166.5000 1097.2500 ;
	    RECT 169.5000 1097.1000 171.3000 1097.2500 ;
	    RECT 260.7000 1098.7500 262.5000 1098.9000 ;
	    RECT 289.5000 1098.7500 291.3000 1098.9000 ;
	    RECT 260.7000 1097.2500 291.3000 1098.7500 ;
	    RECT 260.7000 1097.1000 262.5000 1097.2500 ;
	    RECT 289.5000 1097.1000 291.3000 1097.2500 ;
	    RECT 339.9000 1098.7500 341.7000 1098.9000 ;
	    RECT 351.9000 1098.7500 353.7000 1098.9000 ;
	    RECT 339.9000 1097.2500 353.7000 1098.7500 ;
	    RECT 339.9000 1097.1000 341.7000 1097.2500 ;
	    RECT 351.9000 1097.1000 353.7000 1097.2500 ;
	    RECT 387.9000 1098.7500 389.7000 1098.9000 ;
	    RECT 399.9000 1098.7500 401.7000 1098.9000 ;
	    RECT 387.9000 1097.2500 401.7000 1098.7500 ;
	    RECT 387.9000 1097.1000 389.7000 1097.2500 ;
	    RECT 399.9000 1097.1000 401.7000 1097.2500 ;
	    RECT 591.9000 1098.7500 593.7000 1098.9000 ;
	    RECT 599.2500 1098.7500 600.7500 1109.1000 ;
	    RECT 635.1000 1104.7500 636.9000 1104.9000 ;
	    RECT 642.3000 1104.7500 644.1000 1104.9000 ;
	    RECT 635.1000 1103.2500 644.1000 1104.7500 ;
	    RECT 635.1000 1103.1000 636.9000 1103.2500 ;
	    RECT 642.3000 1103.1000 644.1000 1103.2500 ;
	    RECT 692.7000 1104.7500 694.5000 1104.9000 ;
	    RECT 752.7000 1104.7500 754.5000 1104.9000 ;
	    RECT 692.7000 1103.2500 754.5000 1104.7500 ;
	    RECT 692.7000 1103.1000 694.5000 1103.2500 ;
	    RECT 752.7000 1103.1000 754.5000 1103.2500 ;
	    RECT 1009.5000 1104.7500 1011.3000 1104.9000 ;
	    RECT 1043.1000 1104.7500 1044.9000 1104.9000 ;
	    RECT 1009.5000 1103.2500 1044.9000 1104.7500 ;
	    RECT 1009.5000 1103.1000 1011.3000 1103.2500 ;
	    RECT 1043.1000 1103.1000 1044.9000 1103.2500 ;
	    RECT 1242.3000 1104.7500 1244.1000 1104.9000 ;
	    RECT 1302.3000 1104.7500 1304.1000 1104.9000 ;
	    RECT 1242.3000 1103.2500 1304.1000 1104.7500 ;
	    RECT 1242.3000 1103.1000 1244.1000 1103.2500 ;
	    RECT 1302.3000 1103.1000 1304.1000 1103.2500 ;
	    RECT 1326.3000 1104.7500 1328.1000 1104.9000 ;
	    RECT 1371.9000 1104.7500 1373.7001 1104.9000 ;
	    RECT 1326.3000 1103.2500 1373.7001 1104.7500 ;
	    RECT 1326.3000 1103.1000 1328.1000 1103.2500 ;
	    RECT 1371.9000 1103.1000 1373.7001 1103.2500 ;
	    RECT 1386.3000 1104.7500 1388.1000 1104.9000 ;
	    RECT 1441.5000 1104.7500 1443.3000 1104.9000 ;
	    RECT 1451.1000 1104.7500 1452.9000 1104.9000 ;
	    RECT 1386.3000 1103.2500 1452.9000 1104.7500 ;
	    RECT 1386.3000 1103.1000 1388.1000 1103.2500 ;
	    RECT 1441.5000 1103.1000 1443.3000 1103.2500 ;
	    RECT 1451.1000 1103.1000 1452.9000 1103.2500 ;
	    RECT 1477.5000 1104.7500 1479.3000 1104.9000 ;
	    RECT 1520.7001 1104.7500 1522.5000 1104.9000 ;
	    RECT 1477.5000 1103.2500 1522.5000 1104.7500 ;
	    RECT 1477.5000 1103.1000 1479.3000 1103.2500 ;
	    RECT 1520.7001 1103.1000 1522.5000 1103.2500 ;
	    RECT 591.9000 1097.2500 600.7500 1098.7500 ;
	    RECT 726.3000 1098.7500 728.1000 1098.9000 ;
	    RECT 752.7000 1098.7500 754.5000 1098.9000 ;
	    RECT 726.3000 1097.2500 754.5000 1098.7500 ;
	    RECT 591.9000 1097.1000 593.7000 1097.2500 ;
	    RECT 726.3000 1097.1000 728.1000 1097.2500 ;
	    RECT 752.7000 1097.1000 754.5000 1097.2500 ;
	    RECT 831.9000 1098.7500 833.7000 1098.9000 ;
	    RECT 913.5000 1098.7500 915.3000 1098.9000 ;
	    RECT 831.9000 1097.2500 915.3000 1098.7500 ;
	    RECT 831.9000 1097.1000 833.7000 1097.2500 ;
	    RECT 913.5000 1097.1000 915.3000 1097.2500 ;
	    RECT 1045.5000 1098.7500 1047.3000 1098.9000 ;
	    RECT 1115.1000 1098.7500 1116.9000 1098.9000 ;
	    RECT 1045.5000 1097.2500 1116.9000 1098.7500 ;
	    RECT 1045.5000 1097.1000 1047.3000 1097.2500 ;
	    RECT 1115.1000 1097.1000 1116.9000 1097.2500 ;
	    RECT 1119.9000 1098.7500 1121.7001 1098.9000 ;
	    RECT 1129.5000 1098.7500 1131.3000 1098.9000 ;
	    RECT 1119.9000 1097.2500 1131.3000 1098.7500 ;
	    RECT 1119.9000 1097.1000 1121.7001 1097.2500 ;
	    RECT 1129.5000 1097.1000 1131.3000 1097.2500 ;
	    RECT 1227.9000 1098.7500 1229.7001 1098.9000 ;
	    RECT 1287.9000 1098.7500 1289.7001 1098.9000 ;
	    RECT 1227.9000 1097.2500 1289.7001 1098.7500 ;
	    RECT 1227.9000 1097.1000 1229.7001 1097.2500 ;
	    RECT 1287.9000 1097.1000 1289.7001 1097.2500 ;
	    RECT 1347.9000 1098.7500 1349.7001 1098.9000 ;
	    RECT 1374.3000 1098.7500 1376.1000 1098.9000 ;
	    RECT 1347.9000 1097.2500 1376.1000 1098.7500 ;
	    RECT 1347.9000 1097.1000 1349.7001 1097.2500 ;
	    RECT 1374.3000 1097.1000 1376.1000 1097.2500 ;
	    RECT 1551.9000 1098.7500 1553.7001 1098.9000 ;
	    RECT 1566.3000 1098.7500 1568.1000 1098.9000 ;
	    RECT 1551.9000 1097.2500 1568.1000 1098.7500 ;
	    RECT 1551.9000 1097.1000 1553.7001 1097.2500 ;
	    RECT 1566.3000 1097.1000 1568.1000 1097.2500 ;
	    RECT 143.1000 1092.7500 144.9000 1092.9000 ;
	    RECT 159.9000 1092.7500 161.7000 1092.9000 ;
	    RECT 143.1000 1091.2500 161.7000 1092.7500 ;
	    RECT 143.1000 1091.1000 144.9000 1091.2500 ;
	    RECT 159.9000 1091.1000 161.7000 1091.2500 ;
	    RECT 248.7000 1092.7500 250.5000 1092.9000 ;
	    RECT 272.7000 1092.7500 274.5000 1092.9000 ;
	    RECT 248.7000 1091.2500 274.5000 1092.7500 ;
	    RECT 248.7000 1091.1000 250.5000 1091.2500 ;
	    RECT 272.7000 1091.1000 274.5000 1091.2500 ;
	    RECT 419.1000 1092.7500 420.9000 1092.9000 ;
	    RECT 498.3000 1092.7500 500.1000 1092.9000 ;
	    RECT 419.1000 1091.2500 500.1000 1092.7500 ;
	    RECT 419.1000 1091.1000 420.9000 1091.2500 ;
	    RECT 498.3000 1091.1000 500.1000 1091.2500 ;
	    RECT 884.7000 1092.7500 886.5000 1092.9000 ;
	    RECT 1021.5000 1092.7500 1023.3000 1092.9000 ;
	    RECT 884.7000 1091.2500 1023.3000 1092.7500 ;
	    RECT 884.7000 1091.1000 886.5000 1091.2500 ;
	    RECT 1021.5000 1091.1000 1023.3000 1091.2500 ;
	    RECT 1223.1000 1092.7500 1224.9000 1092.9000 ;
	    RECT 1326.3000 1092.7500 1328.1000 1092.9000 ;
	    RECT 1223.1000 1091.2500 1328.1000 1092.7500 ;
	    RECT 1223.1000 1091.1000 1224.9000 1091.2500 ;
	    RECT 1326.3000 1091.1000 1328.1000 1091.2500 ;
	    RECT 1429.5000 1092.7500 1431.3000 1092.9000 ;
	    RECT 1439.1000 1092.7500 1440.9000 1092.9000 ;
	    RECT 1429.5000 1091.2500 1440.9000 1092.7500 ;
	    RECT 1429.5000 1091.1000 1431.3000 1091.2500 ;
	    RECT 1439.1000 1091.1000 1440.9000 1091.2500 ;
	    RECT 1503.9000 1092.7500 1505.7001 1092.9000 ;
	    RECT 1520.7001 1092.7500 1522.5000 1092.9000 ;
	    RECT 1503.9000 1091.2500 1522.5000 1092.7500 ;
	    RECT 1503.9000 1091.1000 1505.7001 1091.2500 ;
	    RECT 1520.7001 1091.1000 1522.5000 1091.2500 ;
	    RECT 1525.5000 1092.7500 1527.3000 1092.9000 ;
	    RECT 1563.9000 1092.7500 1565.7001 1092.9000 ;
	    RECT 1525.5000 1091.2500 1565.7001 1092.7500 ;
	    RECT 1525.5000 1091.1000 1527.3000 1091.2500 ;
	    RECT 1563.9000 1091.1000 1565.7001 1091.2500 ;
	    RECT 162.3000 1086.7500 164.1000 1086.9000 ;
	    RECT 171.9000 1086.7500 173.7000 1086.9000 ;
	    RECT 162.3000 1085.2500 173.7000 1086.7500 ;
	    RECT 162.3000 1085.1000 164.1000 1085.2500 ;
	    RECT 171.9000 1085.1000 173.7000 1085.2500 ;
	    RECT 191.1000 1086.7500 192.9000 1086.9000 ;
	    RECT 222.3000 1086.7500 224.1000 1086.9000 ;
	    RECT 191.1000 1085.2500 224.1000 1086.7500 ;
	    RECT 191.1000 1085.1000 192.9000 1085.2500 ;
	    RECT 222.3000 1085.1000 224.1000 1085.2500 ;
	    RECT 258.3000 1086.7500 260.1000 1086.9000 ;
	    RECT 303.9000 1086.7500 305.7000 1086.9000 ;
	    RECT 258.3000 1085.2500 305.7000 1086.7500 ;
	    RECT 258.3000 1085.1000 260.1000 1085.2500 ;
	    RECT 303.9000 1085.1000 305.7000 1085.2500 ;
	    RECT 438.3000 1086.7500 440.1000 1086.9000 ;
	    RECT 546.3000 1086.7500 548.1000 1086.9000 ;
	    RECT 438.3000 1085.2500 548.1000 1086.7500 ;
	    RECT 438.3000 1085.1000 440.1000 1085.2500 ;
	    RECT 546.3000 1085.1000 548.1000 1085.2500 ;
	    RECT 647.1000 1086.7500 648.9000 1086.9000 ;
	    RECT 668.7000 1086.7500 670.5000 1086.9000 ;
	    RECT 647.1000 1085.2500 670.5000 1086.7500 ;
	    RECT 647.1000 1085.1000 648.9000 1085.2500 ;
	    RECT 668.7000 1085.1000 670.5000 1085.2500 ;
	    RECT 779.1000 1086.7500 780.9000 1086.9000 ;
	    RECT 822.3000 1086.7500 824.1000 1086.9000 ;
	    RECT 779.1000 1085.2500 824.1000 1086.7500 ;
	    RECT 779.1000 1085.1000 780.9000 1085.2500 ;
	    RECT 822.3000 1085.1000 824.1000 1085.2500 ;
	    RECT 990.3000 1086.7500 992.1000 1086.9000 ;
	    RECT 997.5000 1086.7500 999.3000 1086.9000 ;
	    RECT 990.3000 1085.2500 999.3000 1086.7500 ;
	    RECT 990.3000 1085.1000 992.1000 1085.2500 ;
	    RECT 997.5000 1085.1000 999.3000 1085.2500 ;
	    RECT 1035.9000 1086.7500 1037.7001 1086.9000 ;
	    RECT 1062.3000 1086.7500 1064.1000 1086.9000 ;
	    RECT 1110.3000 1086.7500 1112.1000 1086.9000 ;
	    RECT 1035.9000 1085.2500 1112.1000 1086.7500 ;
	    RECT 1035.9000 1085.1000 1037.7001 1085.2500 ;
	    RECT 1062.3000 1085.1000 1064.1000 1085.2500 ;
	    RECT 1110.3000 1085.1000 1112.1000 1085.2500 ;
	    RECT 1179.9000 1086.7500 1181.7001 1086.9000 ;
	    RECT 1343.1000 1086.7500 1344.9000 1086.9000 ;
	    RECT 1179.9000 1085.2500 1344.9000 1086.7500 ;
	    RECT 1179.9000 1085.1000 1181.7001 1085.2500 ;
	    RECT 1343.1000 1085.1000 1344.9000 1085.2500 ;
	    RECT 1417.5000 1086.7500 1419.3000 1086.9000 ;
	    RECT 1501.5000 1086.7500 1503.3000 1086.9000 ;
	    RECT 1417.5000 1085.2500 1503.3000 1086.7500 ;
	    RECT 1417.5000 1085.1000 1419.3000 1085.2500 ;
	    RECT 1501.5000 1085.1000 1503.3000 1085.2500 ;
	    RECT 1511.1000 1086.7500 1512.9000 1086.9000 ;
	    RECT 1535.1000 1086.7500 1536.9000 1086.9000 ;
	    RECT 1511.1000 1085.2500 1536.9000 1086.7500 ;
	    RECT 1511.1000 1085.1000 1512.9000 1085.2500 ;
	    RECT 1535.1000 1085.1000 1536.9000 1085.2500 ;
	    RECT 56.7000 1080.7500 58.5000 1080.9000 ;
	    RECT 191.1000 1080.7500 192.9000 1080.9000 ;
	    RECT 56.7000 1079.2500 192.9000 1080.7500 ;
	    RECT 56.7000 1079.1000 58.5000 1079.2500 ;
	    RECT 191.1000 1079.1000 192.9000 1079.2500 ;
	    RECT 299.1000 1080.7500 300.9000 1080.9000 ;
	    RECT 618.3000 1080.7500 620.1000 1080.9000 ;
	    RECT 299.1000 1079.2500 620.1000 1080.7500 ;
	    RECT 299.1000 1079.1000 300.9000 1079.2500 ;
	    RECT 618.3000 1079.1000 620.1000 1079.2500 ;
	    RECT 627.9000 1080.7500 629.7000 1080.9000 ;
	    RECT 642.3000 1080.7500 644.1000 1080.9000 ;
	    RECT 627.9000 1079.2500 644.1000 1080.7500 ;
	    RECT 627.9000 1079.1000 629.7000 1079.2500 ;
	    RECT 642.3000 1079.1000 644.1000 1079.2500 ;
	    RECT 1009.5000 1080.7500 1011.3000 1080.9000 ;
	    RECT 1021.5000 1080.7500 1023.3000 1080.9000 ;
	    RECT 1009.5000 1079.2500 1023.3000 1080.7500 ;
	    RECT 1009.5000 1079.1000 1011.3000 1079.2500 ;
	    RECT 1021.5000 1079.1000 1023.3000 1079.2500 ;
	    RECT 1095.9000 1080.7500 1097.7001 1080.9000 ;
	    RECT 1119.9000 1080.7500 1121.7001 1080.9000 ;
	    RECT 1095.9000 1079.2500 1121.7001 1080.7500 ;
	    RECT 1095.9000 1079.1000 1097.7001 1079.2500 ;
	    RECT 1119.9000 1079.1000 1121.7001 1079.2500 ;
	    RECT 1153.5000 1080.7500 1155.3000 1080.9000 ;
	    RECT 1268.7001 1080.7500 1270.5000 1080.9000 ;
	    RECT 1153.5000 1079.2500 1270.5000 1080.7500 ;
	    RECT 1153.5000 1079.1000 1155.3000 1079.2500 ;
	    RECT 1268.7001 1079.1000 1270.5000 1079.2500 ;
	    RECT 1280.7001 1080.7500 1282.5000 1080.9000 ;
	    RECT 1489.5000 1080.7500 1491.3000 1080.9000 ;
	    RECT 1280.7001 1079.2500 1491.3000 1080.7500 ;
	    RECT 1280.7001 1079.1000 1282.5000 1079.2500 ;
	    RECT 1489.5000 1079.1000 1491.3000 1079.2500 ;
	    RECT 1503.9000 1080.7500 1505.7001 1080.9000 ;
	    RECT 1532.7001 1080.7500 1534.5000 1080.9000 ;
	    RECT 1503.9000 1079.2500 1534.5000 1080.7500 ;
	    RECT 1503.9000 1079.1000 1505.7001 1079.2500 ;
	    RECT 1532.7001 1079.1000 1534.5000 1079.2500 ;
	    RECT 1537.5000 1080.7500 1539.3000 1080.9000 ;
	    RECT 1563.9000 1080.7500 1565.7001 1080.9000 ;
	    RECT 1537.5000 1079.2500 1565.7001 1080.7500 ;
	    RECT 1537.5000 1079.1000 1539.3000 1079.2500 ;
	    RECT 1563.9000 1079.1000 1565.7001 1079.2500 ;
	    RECT 133.5000 1074.7500 135.3000 1074.9000 ;
	    RECT 164.7000 1074.7500 166.5000 1074.9000 ;
	    RECT 133.5000 1073.2500 166.5000 1074.7500 ;
	    RECT 133.5000 1073.1000 135.3000 1073.2500 ;
	    RECT 164.7000 1073.1000 166.5000 1073.2500 ;
	    RECT 239.1000 1074.7500 240.9000 1074.9000 ;
	    RECT 253.5000 1074.7500 255.3000 1074.9000 ;
	    RECT 385.5000 1074.7500 387.3000 1074.9000 ;
	    RECT 239.1000 1073.2500 387.3000 1074.7500 ;
	    RECT 239.1000 1073.1000 240.9000 1073.2500 ;
	    RECT 253.5000 1073.1000 255.3000 1073.2500 ;
	    RECT 385.5000 1073.1000 387.3000 1073.2500 ;
	    RECT 846.3000 1074.7500 848.1000 1074.9000 ;
	    RECT 853.5000 1074.7500 855.3000 1074.9000 ;
	    RECT 846.3000 1073.2500 855.3000 1074.7500 ;
	    RECT 846.3000 1073.1000 848.1000 1073.2500 ;
	    RECT 853.5000 1073.1000 855.3000 1073.2500 ;
	    RECT 971.1000 1074.7500 972.9000 1074.9000 ;
	    RECT 987.9000 1074.7500 989.7000 1074.9000 ;
	    RECT 971.1000 1073.2500 989.7000 1074.7500 ;
	    RECT 971.1000 1073.1000 972.9000 1073.2500 ;
	    RECT 987.9000 1073.1000 989.7000 1073.2500 ;
	    RECT 1055.1000 1074.7500 1056.9000 1074.9000 ;
	    RECT 1067.1000 1074.7500 1068.9000 1074.9000 ;
	    RECT 1055.1000 1073.2500 1068.9000 1074.7500 ;
	    RECT 1055.1000 1073.1000 1056.9000 1073.2500 ;
	    RECT 1067.1000 1073.1000 1068.9000 1073.2500 ;
	    RECT 1182.3000 1074.7500 1184.1000 1074.9000 ;
	    RECT 1242.3000 1074.7500 1244.1000 1074.9000 ;
	    RECT 1182.3000 1073.2500 1244.1000 1074.7500 ;
	    RECT 1182.3000 1073.1000 1184.1000 1073.2500 ;
	    RECT 1242.3000 1073.1000 1244.1000 1073.2500 ;
	    RECT 1247.1000 1074.7500 1248.9000 1074.9000 ;
	    RECT 1417.5000 1074.7500 1419.3000 1074.9000 ;
	    RECT 1247.1000 1073.2500 1419.3000 1074.7500 ;
	    RECT 1247.1000 1073.1000 1248.9000 1073.2500 ;
	    RECT 1417.5000 1073.1000 1419.3000 1073.2500 ;
	    RECT 1544.7001 1074.7500 1546.5000 1074.9000 ;
	    RECT 1561.5000 1074.7500 1563.3000 1074.9000 ;
	    RECT 1544.7001 1073.2500 1563.3000 1074.7500 ;
	    RECT 1544.7001 1073.1000 1546.5000 1073.2500 ;
	    RECT 1561.5000 1073.1000 1563.3000 1073.2500 ;
	    RECT 143.1000 1068.7500 144.9000 1068.9000 ;
	    RECT 133.6500 1067.2500 144.9000 1068.7500 ;
	    RECT 133.6500 1062.9000 135.1500 1067.2500 ;
	    RECT 143.1000 1067.1000 144.9000 1067.2500 ;
	    RECT 198.3000 1068.7500 200.1000 1068.9000 ;
	    RECT 222.3000 1068.7500 224.1000 1068.9000 ;
	    RECT 198.3000 1067.2500 224.1000 1068.7500 ;
	    RECT 198.3000 1067.1000 200.1000 1067.2500 ;
	    RECT 222.3000 1067.1000 224.1000 1067.2500 ;
	    RECT 231.9000 1068.7500 233.7000 1068.9000 ;
	    RECT 258.3000 1068.7500 260.1000 1068.9000 ;
	    RECT 231.9000 1067.2500 260.1000 1068.7500 ;
	    RECT 231.9000 1067.1000 233.7000 1067.2500 ;
	    RECT 258.3000 1067.1000 260.1000 1067.2500 ;
	    RECT 327.9000 1068.7500 329.7000 1068.9000 ;
	    RECT 380.7000 1068.7500 382.5000 1068.9000 ;
	    RECT 327.9000 1067.2500 382.5000 1068.7500 ;
	    RECT 327.9000 1067.1000 329.7000 1067.2500 ;
	    RECT 380.7000 1067.1000 382.5000 1067.2500 ;
	    RECT 517.5000 1068.7500 519.3000 1068.9000 ;
	    RECT 541.5000 1068.7500 543.3000 1068.9000 ;
	    RECT 517.5000 1067.2500 543.3000 1068.7500 ;
	    RECT 517.5000 1067.1000 519.3000 1067.2500 ;
	    RECT 541.5000 1067.1000 543.3000 1067.2500 ;
	    RECT 625.5000 1068.7500 627.3000 1068.9000 ;
	    RECT 635.1000 1068.7500 636.9000 1068.9000 ;
	    RECT 625.5000 1067.2500 636.9000 1068.7500 ;
	    RECT 625.5000 1067.1000 627.3000 1067.2500 ;
	    RECT 635.1000 1067.1000 636.9000 1067.2500 ;
	    RECT 702.3000 1068.7500 704.1000 1068.9000 ;
	    RECT 747.9000 1068.7500 749.7000 1068.9000 ;
	    RECT 702.3000 1067.2500 749.7000 1068.7500 ;
	    RECT 702.3000 1067.1000 704.1000 1067.2500 ;
	    RECT 747.9000 1067.1000 749.7000 1067.2500 ;
	    RECT 915.9000 1068.7500 917.7000 1068.9000 ;
	    RECT 995.1000 1068.7500 996.9000 1068.9000 ;
	    RECT 915.9000 1067.2500 996.9000 1068.7500 ;
	    RECT 915.9000 1067.1000 917.7000 1067.2500 ;
	    RECT 995.1000 1067.1000 996.9000 1067.2500 ;
	    RECT 1191.9000 1068.7500 1193.7001 1068.9000 ;
	    RECT 1213.5000 1068.7500 1215.3000 1068.9000 ;
	    RECT 1191.9000 1067.2500 1215.3000 1068.7500 ;
	    RECT 1191.9000 1067.1000 1193.7001 1067.2500 ;
	    RECT 1213.5000 1067.1000 1215.3000 1067.2500 ;
	    RECT 1316.7001 1068.7500 1318.5000 1068.9000 ;
	    RECT 1427.1000 1068.7500 1428.9000 1068.9000 ;
	    RECT 1316.7001 1067.2500 1428.9000 1068.7500 ;
	    RECT 1316.7001 1067.1000 1318.5000 1067.2500 ;
	    RECT 1427.1000 1067.1000 1428.9000 1067.2500 ;
	    RECT 1482.3000 1068.7500 1484.1000 1068.9000 ;
	    RECT 1515.9000 1068.7500 1517.7001 1068.9000 ;
	    RECT 1482.3000 1067.2500 1517.7001 1068.7500 ;
	    RECT 1482.3000 1067.1000 1484.1000 1067.2500 ;
	    RECT 1515.9000 1067.1000 1517.7001 1067.2500 ;
	    RECT 1520.7001 1068.7500 1522.5000 1068.9000 ;
	    RECT 1561.5000 1068.7500 1563.3000 1068.9000 ;
	    RECT 1520.7001 1067.2500 1563.3000 1068.7500 ;
	    RECT 1520.7001 1067.1000 1522.5000 1067.2500 ;
	    RECT 1561.5000 1067.1000 1563.3000 1067.2500 ;
	    RECT 133.5000 1061.1000 135.3000 1062.9000 ;
	    RECT 231.9000 1062.7500 233.7000 1062.9000 ;
	    RECT 275.1000 1062.7500 276.9000 1062.9000 ;
	    RECT 231.9000 1061.2500 276.9000 1062.7500 ;
	    RECT 231.9000 1061.1000 233.7000 1061.2500 ;
	    RECT 275.1000 1061.1000 276.9000 1061.2500 ;
	    RECT 325.5000 1062.7500 327.3000 1062.9000 ;
	    RECT 373.5000 1062.7500 375.3000 1062.9000 ;
	    RECT 390.3000 1062.7500 392.1000 1062.9000 ;
	    RECT 325.5000 1061.2500 392.1000 1062.7500 ;
	    RECT 325.5000 1061.1000 327.3000 1061.2500 ;
	    RECT 373.5000 1061.1000 375.3000 1061.2500 ;
	    RECT 390.3000 1061.1000 392.1000 1061.2500 ;
	    RECT 524.7000 1062.7500 526.5000 1062.9000 ;
	    RECT 555.9000 1062.7500 557.7000 1062.9000 ;
	    RECT 524.7000 1061.2500 557.7000 1062.7500 ;
	    RECT 524.7000 1061.1000 526.5000 1061.2500 ;
	    RECT 555.9000 1061.1000 557.7000 1061.2500 ;
	    RECT 627.9000 1062.7500 629.7000 1062.9000 ;
	    RECT 651.9000 1062.7500 653.7000 1062.9000 ;
	    RECT 627.9000 1061.2500 653.7000 1062.7500 ;
	    RECT 627.9000 1061.1000 629.7000 1061.2500 ;
	    RECT 651.9000 1061.1000 653.7000 1061.2500 ;
	    RECT 1187.1000 1062.7500 1188.9000 1062.9000 ;
	    RECT 1208.7001 1062.7500 1210.5000 1062.9000 ;
	    RECT 1187.1000 1061.2500 1210.5000 1062.7500 ;
	    RECT 1187.1000 1061.1000 1188.9000 1061.2500 ;
	    RECT 1208.7001 1061.1000 1210.5000 1061.2500 ;
	    RECT 1213.5000 1062.7500 1215.3000 1062.9000 ;
	    RECT 1249.5000 1062.7500 1251.3000 1062.9000 ;
	    RECT 1213.5000 1061.2500 1251.3000 1062.7500 ;
	    RECT 1213.5000 1061.1000 1215.3000 1061.2500 ;
	    RECT 1249.5000 1061.1000 1251.3000 1061.2500 ;
	    RECT 1431.9000 1062.7500 1433.7001 1062.9000 ;
	    RECT 1482.3000 1062.7500 1484.1000 1062.9000 ;
	    RECT 1431.9000 1061.2500 1484.1000 1062.7500 ;
	    RECT 1431.9000 1061.1000 1433.7001 1061.2500 ;
	    RECT 1482.3000 1061.1000 1484.1000 1061.2500 ;
	    RECT 1515.9000 1062.7500 1517.7001 1062.9000 ;
	    RECT 1527.9000 1062.7500 1529.7001 1062.9000 ;
	    RECT 1515.9000 1061.2500 1529.7001 1062.7500 ;
	    RECT 1515.9000 1061.1000 1517.7001 1061.2500 ;
	    RECT 1527.9000 1061.1000 1529.7001 1061.2500 ;
	    RECT 176.7000 1056.7500 178.5000 1056.9000 ;
	    RECT 217.5000 1056.7500 219.3000 1056.9000 ;
	    RECT 176.7000 1055.2500 219.3000 1056.7500 ;
	    RECT 176.7000 1055.1000 178.5000 1055.2500 ;
	    RECT 217.5000 1055.1000 219.3000 1055.2500 ;
	    RECT 222.3000 1056.7500 224.1000 1056.9000 ;
	    RECT 308.7000 1056.7500 310.5000 1056.9000 ;
	    RECT 222.3000 1055.2500 310.5000 1056.7500 ;
	    RECT 222.3000 1055.1000 224.1000 1055.2500 ;
	    RECT 308.7000 1055.1000 310.5000 1055.2500 ;
	    RECT 606.3000 1056.7500 608.1000 1056.9000 ;
	    RECT 651.9000 1056.7500 653.7000 1056.9000 ;
	    RECT 606.3000 1055.2500 653.7000 1056.7500 ;
	    RECT 606.3000 1055.1000 608.1000 1055.2500 ;
	    RECT 651.9000 1055.1000 653.7000 1055.2500 ;
	    RECT 673.5000 1056.7500 675.3000 1056.9000 ;
	    RECT 733.5000 1056.7500 735.3000 1056.9000 ;
	    RECT 673.5000 1055.2500 735.3000 1056.7500 ;
	    RECT 673.5000 1055.1000 675.3000 1055.2500 ;
	    RECT 733.5000 1055.1000 735.3000 1055.2500 ;
	    RECT 745.5000 1056.7500 747.3000 1056.9000 ;
	    RECT 752.7000 1056.7500 754.5000 1056.9000 ;
	    RECT 745.5000 1055.2500 754.5000 1056.7500 ;
	    RECT 745.5000 1055.1000 747.3000 1055.2500 ;
	    RECT 752.7000 1055.1000 754.5000 1055.2500 ;
	    RECT 1266.3000 1056.7500 1268.1000 1056.9000 ;
	    RECT 1319.1000 1056.7500 1320.9000 1056.9000 ;
	    RECT 1266.3000 1055.2500 1320.9000 1056.7500 ;
	    RECT 1266.3000 1055.1000 1268.1000 1055.2500 ;
	    RECT 1319.1000 1055.1000 1320.9000 1055.2500 ;
	    RECT 83.1000 1050.7500 84.9000 1050.9000 ;
	    RECT 162.3000 1050.7500 164.1000 1050.9000 ;
	    RECT 83.1000 1049.2500 164.1000 1050.7500 ;
	    RECT 83.1000 1049.1000 84.9000 1049.2500 ;
	    RECT 162.3000 1049.1000 164.1000 1049.2500 ;
	    RECT 217.5000 1050.7500 219.3000 1050.9000 ;
	    RECT 267.9000 1050.7500 269.7000 1050.9000 ;
	    RECT 217.5000 1049.2500 269.7000 1050.7500 ;
	    RECT 217.5000 1049.1000 219.3000 1049.2500 ;
	    RECT 267.9000 1049.1000 269.7000 1049.2500 ;
	    RECT 284.7000 1050.7500 286.5000 1050.9000 ;
	    RECT 291.9000 1050.7500 293.7000 1050.9000 ;
	    RECT 284.7000 1049.2500 293.7000 1050.7500 ;
	    RECT 284.7000 1049.1000 286.5000 1049.2500 ;
	    RECT 291.9000 1049.1000 293.7000 1049.2500 ;
	    RECT 308.7000 1050.7500 310.5000 1050.9000 ;
	    RECT 363.9000 1050.7500 365.7000 1050.9000 ;
	    RECT 308.7000 1049.2500 365.7000 1050.7500 ;
	    RECT 308.7000 1049.1000 310.5000 1049.2500 ;
	    RECT 363.9000 1049.1000 365.7000 1049.2500 ;
	    RECT 471.9000 1050.7500 473.7000 1050.9000 ;
	    RECT 486.3000 1050.7500 488.1000 1050.9000 ;
	    RECT 510.3000 1050.7500 512.1000 1050.9000 ;
	    RECT 517.5000 1050.7500 519.3000 1050.9000 ;
	    RECT 471.9000 1049.2500 519.3000 1050.7500 ;
	    RECT 471.9000 1049.1000 473.7000 1049.2500 ;
	    RECT 486.3000 1049.1000 488.1000 1049.2500 ;
	    RECT 510.3000 1049.1000 512.1000 1049.2500 ;
	    RECT 517.5000 1049.1000 519.3000 1049.2500 ;
	    RECT 757.5000 1050.7500 759.3000 1050.9000 ;
	    RECT 781.5000 1050.7500 783.3000 1050.9000 ;
	    RECT 757.5000 1049.2500 783.3000 1050.7500 ;
	    RECT 757.5000 1049.1000 759.3000 1049.2500 ;
	    RECT 781.5000 1049.1000 783.3000 1049.2500 ;
	    RECT 1011.9000 1050.7500 1013.7000 1050.9000 ;
	    RECT 1081.5000 1050.7500 1083.3000 1050.9000 ;
	    RECT 1011.9000 1049.2500 1083.3000 1050.7500 ;
	    RECT 1011.9000 1049.1000 1013.7000 1049.2500 ;
	    RECT 1081.5000 1049.1000 1083.3000 1049.2500 ;
	    RECT 1465.5000 1050.7500 1467.3000 1050.9000 ;
	    RECT 1470.3000 1050.7500 1472.1000 1050.9000 ;
	    RECT 1465.5000 1049.2500 1472.1000 1050.7500 ;
	    RECT 1465.5000 1049.1000 1467.3000 1049.2500 ;
	    RECT 1470.3000 1049.1000 1472.1000 1049.2500 ;
	    RECT 1506.3000 1050.7500 1508.1000 1050.9000 ;
	    RECT 1513.5000 1050.7500 1515.3000 1050.9000 ;
	    RECT 1506.3000 1049.2500 1515.3000 1050.7500 ;
	    RECT 1506.3000 1049.1000 1508.1000 1049.2500 ;
	    RECT 1513.5000 1049.1000 1515.3000 1049.2500 ;
	    RECT 1520.7001 1049.1000 1522.5000 1050.9000 ;
	    RECT 18.3000 1044.7500 20.1000 1044.9000 ;
	    RECT 56.7000 1044.7500 58.5000 1044.9000 ;
	    RECT 18.3000 1043.2500 58.5000 1044.7500 ;
	    RECT 18.3000 1043.1000 20.1000 1043.2500 ;
	    RECT 56.7000 1043.1000 58.5000 1043.2500 ;
	    RECT 143.1000 1044.7500 144.9000 1044.9000 ;
	    RECT 183.9000 1044.7500 185.7000 1044.9000 ;
	    RECT 143.1000 1043.2500 185.7000 1044.7500 ;
	    RECT 143.1000 1043.1000 144.9000 1043.2500 ;
	    RECT 183.9000 1043.1000 185.7000 1043.2500 ;
	    RECT 270.3000 1044.7500 272.1000 1044.9000 ;
	    RECT 337.5000 1044.7500 339.3000 1044.9000 ;
	    RECT 476.7000 1044.7500 478.5000 1044.9000 ;
	    RECT 495.9000 1044.7500 497.7000 1044.9000 ;
	    RECT 270.3000 1043.2500 497.7000 1044.7500 ;
	    RECT 270.3000 1043.1000 272.1000 1043.2500 ;
	    RECT 337.5000 1043.1000 339.3000 1043.2500 ;
	    RECT 476.7000 1043.1000 478.5000 1043.2500 ;
	    RECT 495.9000 1043.1000 497.7000 1043.2500 ;
	    RECT 639.9000 1044.7500 641.7000 1044.9000 ;
	    RECT 678.3000 1044.7500 680.1000 1044.9000 ;
	    RECT 639.9000 1043.2500 680.1000 1044.7500 ;
	    RECT 639.9000 1043.1000 641.7000 1043.2500 ;
	    RECT 678.3000 1043.1000 680.1000 1043.2500 ;
	    RECT 750.3000 1044.7500 752.1000 1044.9000 ;
	    RECT 767.1000 1044.7500 768.9000 1044.9000 ;
	    RECT 750.3000 1043.2500 768.9000 1044.7500 ;
	    RECT 750.3000 1043.1000 752.1000 1043.2500 ;
	    RECT 767.1000 1043.1000 768.9000 1043.2500 ;
	    RECT 1146.3000 1044.7500 1148.1000 1044.9000 ;
	    RECT 1189.5000 1044.7500 1191.3000 1044.9000 ;
	    RECT 1146.3000 1043.2500 1191.3000 1044.7500 ;
	    RECT 1146.3000 1043.1000 1148.1000 1043.2500 ;
	    RECT 1189.5000 1043.1000 1191.3000 1043.2500 ;
	    RECT 1196.7001 1044.7500 1198.5000 1044.9000 ;
	    RECT 1215.9000 1044.7500 1217.7001 1044.9000 ;
	    RECT 1196.7001 1043.2500 1217.7001 1044.7500 ;
	    RECT 1196.7001 1043.1000 1198.5000 1043.2500 ;
	    RECT 1215.9000 1043.1000 1217.7001 1043.2500 ;
	    RECT 1237.5000 1044.7500 1239.3000 1044.9000 ;
	    RECT 1247.1000 1044.7500 1248.9000 1044.9000 ;
	    RECT 1237.5000 1043.2500 1248.9000 1044.7500 ;
	    RECT 1237.5000 1043.1000 1239.3000 1043.2500 ;
	    RECT 1247.1000 1043.1000 1248.9000 1043.2500 ;
	    RECT 1259.1000 1044.7500 1260.9000 1044.9000 ;
	    RECT 1292.7001 1044.7500 1294.5000 1044.9000 ;
	    RECT 1259.1000 1043.2500 1294.5000 1044.7500 ;
	    RECT 1259.1000 1043.1000 1260.9000 1043.2500 ;
	    RECT 1292.7001 1043.1000 1294.5000 1043.2500 ;
	    RECT 140.7000 1038.7500 142.5000 1038.9000 ;
	    RECT 167.1000 1038.7500 168.9000 1038.9000 ;
	    RECT 140.7000 1037.2500 168.9000 1038.7500 ;
	    RECT 140.7000 1037.1000 142.5000 1037.2500 ;
	    RECT 167.1000 1037.1000 168.9000 1037.2500 ;
	    RECT 181.5000 1038.7500 183.3000 1038.9000 ;
	    RECT 188.7000 1038.7500 190.5000 1038.9000 ;
	    RECT 181.5000 1037.2500 190.5000 1038.7500 ;
	    RECT 181.5000 1037.1000 183.3000 1037.2500 ;
	    RECT 188.7000 1037.1000 190.5000 1037.2500 ;
	    RECT 195.9000 1038.7500 197.7000 1038.9000 ;
	    RECT 229.5000 1038.7500 231.3000 1038.9000 ;
	    RECT 195.9000 1037.2500 231.3000 1038.7500 ;
	    RECT 195.9000 1037.1000 197.7000 1037.2500 ;
	    RECT 229.5000 1037.1000 231.3000 1037.2500 ;
	    RECT 272.7000 1038.7500 274.5000 1038.9000 ;
	    RECT 313.5000 1038.7500 315.3000 1038.9000 ;
	    RECT 272.7000 1037.2500 315.3000 1038.7500 ;
	    RECT 272.7000 1037.1000 274.5000 1037.2500 ;
	    RECT 313.5000 1037.1000 315.3000 1037.2500 ;
	    RECT 339.9000 1038.7500 341.7000 1038.9000 ;
	    RECT 344.7000 1038.7500 346.5000 1038.9000 ;
	    RECT 339.9000 1037.2500 346.5000 1038.7500 ;
	    RECT 339.9000 1037.1000 341.7000 1037.2500 ;
	    RECT 344.7000 1037.1000 346.5000 1037.2500 ;
	    RECT 671.1000 1038.7500 672.9000 1038.9000 ;
	    RECT 699.9000 1038.7500 701.7000 1038.9000 ;
	    RECT 671.1000 1037.2500 701.7000 1038.7500 ;
	    RECT 671.1000 1037.1000 672.9000 1037.2500 ;
	    RECT 699.9000 1037.1000 701.7000 1037.2500 ;
	    RECT 762.3000 1038.7500 764.1000 1038.9000 ;
	    RECT 807.9000 1038.7500 809.7000 1038.9000 ;
	    RECT 762.3000 1037.2500 809.7000 1038.7500 ;
	    RECT 762.3000 1037.1000 764.1000 1037.2500 ;
	    RECT 807.9000 1037.1000 809.7000 1037.2500 ;
	    RECT 815.1000 1038.7500 816.9000 1038.9000 ;
	    RECT 829.5000 1038.7500 831.3000 1038.9000 ;
	    RECT 841.5000 1038.7500 843.3000 1038.9000 ;
	    RECT 815.1000 1037.2500 843.3000 1038.7500 ;
	    RECT 815.1000 1037.1000 816.9000 1037.2500 ;
	    RECT 829.5000 1037.1000 831.3000 1037.2500 ;
	    RECT 841.5000 1037.1000 843.3000 1037.2500 ;
	    RECT 903.9000 1038.7500 905.7000 1038.9000 ;
	    RECT 939.9000 1038.7500 941.7000 1038.9000 ;
	    RECT 903.9000 1037.2500 941.7000 1038.7500 ;
	    RECT 903.9000 1037.1000 905.7000 1037.2500 ;
	    RECT 939.9000 1037.1000 941.7000 1037.2500 ;
	    RECT 1208.7001 1038.7500 1210.5000 1038.9000 ;
	    RECT 1287.9000 1038.7500 1289.7001 1038.9000 ;
	    RECT 1297.5000 1038.7500 1299.3000 1038.9000 ;
	    RECT 1208.7001 1037.2500 1299.3000 1038.7500 ;
	    RECT 1208.7001 1037.1000 1210.5000 1037.2500 ;
	    RECT 1287.9000 1037.1000 1289.7001 1037.2500 ;
	    RECT 1297.5000 1037.1000 1299.3000 1037.2500 ;
	    RECT 99.9000 1032.7500 101.7000 1032.9000 ;
	    RECT 145.5000 1032.7500 147.3000 1032.9000 ;
	    RECT 99.9000 1031.2500 147.3000 1032.7500 ;
	    RECT 99.9000 1031.1000 101.7000 1031.2500 ;
	    RECT 145.5000 1031.1000 147.3000 1031.2500 ;
	    RECT 150.3000 1032.7500 152.1000 1032.9000 ;
	    RECT 176.7000 1032.7500 178.5000 1032.9000 ;
	    RECT 150.3000 1031.2500 178.5000 1032.7500 ;
	    RECT 150.3000 1031.1000 152.1000 1031.2500 ;
	    RECT 176.7000 1031.1000 178.5000 1031.2500 ;
	    RECT 219.9000 1032.7500 221.7000 1032.9000 ;
	    RECT 265.5000 1032.7500 267.3000 1032.9000 ;
	    RECT 219.9000 1031.2500 267.3000 1032.7500 ;
	    RECT 219.9000 1031.1000 221.7000 1031.2500 ;
	    RECT 265.5000 1031.1000 267.3000 1031.2500 ;
	    RECT 277.5000 1032.7500 279.3000 1032.9000 ;
	    RECT 294.3000 1032.7500 296.1000 1032.9000 ;
	    RECT 277.5000 1031.2500 296.1000 1032.7500 ;
	    RECT 277.5000 1031.1000 279.3000 1031.2500 ;
	    RECT 294.3000 1031.1000 296.1000 1031.2500 ;
	    RECT 335.1000 1032.7500 336.9000 1032.9000 ;
	    RECT 409.5000 1032.7500 411.3000 1032.9000 ;
	    RECT 335.1000 1031.2500 411.3000 1032.7500 ;
	    RECT 335.1000 1031.1000 336.9000 1031.2500 ;
	    RECT 409.5000 1031.1000 411.3000 1031.2500 ;
	    RECT 714.3000 1032.7500 716.1000 1032.9000 ;
	    RECT 793.5000 1032.7500 795.3000 1032.9000 ;
	    RECT 714.3000 1031.2500 795.3000 1032.7500 ;
	    RECT 714.3000 1031.1000 716.1000 1031.2500 ;
	    RECT 793.5000 1031.1000 795.3000 1031.2500 ;
	    RECT 805.5000 1032.7500 807.3000 1032.9000 ;
	    RECT 815.1000 1032.7500 816.9000 1032.9000 ;
	    RECT 805.5000 1031.2500 816.9000 1032.7500 ;
	    RECT 805.5000 1031.1000 807.3000 1031.2500 ;
	    RECT 815.1000 1031.1000 816.9000 1031.2500 ;
	    RECT 889.5000 1032.7500 891.3000 1032.9000 ;
	    RECT 915.9000 1032.7500 917.7000 1032.9000 ;
	    RECT 889.5000 1031.2500 917.7000 1032.7500 ;
	    RECT 889.5000 1031.1000 891.3000 1031.2500 ;
	    RECT 915.9000 1031.1000 917.7000 1031.2500 ;
	    RECT 1295.1000 1032.7500 1296.9000 1032.9000 ;
	    RECT 1371.9000 1032.7500 1373.7001 1032.9000 ;
	    RECT 1295.1000 1031.2500 1373.7001 1032.7500 ;
	    RECT 1295.1000 1031.1000 1296.9000 1031.2500 ;
	    RECT 1371.9000 1031.1000 1373.7001 1031.2500 ;
	    RECT 1520.8500 1026.9000 1522.3500 1049.1000 ;
	    RECT 1544.7001 1034.1000 1546.5000 1035.9000 ;
	    RECT 1544.8500 1032.7500 1546.3500 1034.1000 ;
	    RECT 1544.8500 1031.2500 1565.5500 1032.7500 ;
	    RECT 1564.0500 1026.9000 1565.5500 1031.2500 ;
	    RECT 138.3000 1026.7500 140.1000 1026.9000 ;
	    RECT 150.3000 1026.7500 152.1000 1026.9000 ;
	    RECT 138.3000 1025.2500 152.1000 1026.7500 ;
	    RECT 138.3000 1025.1000 140.1000 1025.2500 ;
	    RECT 150.3000 1025.1000 152.1000 1025.2500 ;
	    RECT 243.9000 1026.7500 245.7000 1026.9000 ;
	    RECT 303.9000 1026.7500 305.7000 1026.9000 ;
	    RECT 243.9000 1025.2500 305.7000 1026.7500 ;
	    RECT 243.9000 1025.1000 245.7000 1025.2500 ;
	    RECT 303.9000 1025.1000 305.7000 1025.2500 ;
	    RECT 311.1000 1026.7500 312.9000 1026.9000 ;
	    RECT 349.5000 1026.7500 351.3000 1026.9000 ;
	    RECT 356.7000 1026.7500 358.5000 1026.9000 ;
	    RECT 311.1000 1025.2500 358.5000 1026.7500 ;
	    RECT 311.1000 1025.1000 312.9000 1025.2500 ;
	    RECT 349.5000 1025.1000 351.3000 1025.2500 ;
	    RECT 356.7000 1025.1000 358.5000 1025.2500 ;
	    RECT 560.7000 1026.7500 562.5000 1026.9000 ;
	    RECT 678.3000 1026.7500 680.1000 1026.9000 ;
	    RECT 560.7000 1025.2500 680.1000 1026.7500 ;
	    RECT 560.7000 1025.1000 562.5000 1025.2500 ;
	    RECT 678.3000 1025.1000 680.1000 1025.2500 ;
	    RECT 702.3000 1026.7500 704.1000 1026.9000 ;
	    RECT 755.1000 1026.7500 756.9000 1026.9000 ;
	    RECT 702.3000 1025.2500 756.9000 1026.7500 ;
	    RECT 702.3000 1025.1000 704.1000 1025.2500 ;
	    RECT 755.1000 1025.1000 756.9000 1025.2500 ;
	    RECT 803.1000 1026.7500 804.9000 1026.9000 ;
	    RECT 807.9000 1026.7500 809.7000 1026.9000 ;
	    RECT 819.9000 1026.7500 821.7000 1026.9000 ;
	    RECT 803.1000 1025.2500 821.7000 1026.7500 ;
	    RECT 803.1000 1025.1000 804.9000 1025.2500 ;
	    RECT 807.9000 1025.1000 809.7000 1025.2500 ;
	    RECT 819.9000 1025.1000 821.7000 1025.2500 ;
	    RECT 913.5000 1026.7500 915.3000 1026.9000 ;
	    RECT 1201.5000 1026.7500 1203.3000 1026.9000 ;
	    RECT 913.5000 1025.2500 1203.3000 1026.7500 ;
	    RECT 913.5000 1025.1000 915.3000 1025.2500 ;
	    RECT 1201.5000 1025.1000 1203.3000 1025.2500 ;
	    RECT 1206.3000 1026.7500 1208.1000 1026.9000 ;
	    RECT 1220.7001 1026.7500 1222.5000 1026.9000 ;
	    RECT 1206.3000 1025.2500 1222.5000 1026.7500 ;
	    RECT 1206.3000 1025.1000 1208.1000 1025.2500 ;
	    RECT 1220.7001 1025.1000 1222.5000 1025.2500 ;
	    RECT 1307.1000 1026.7500 1308.9000 1026.9000 ;
	    RECT 1314.3000 1026.7500 1316.1000 1026.9000 ;
	    RECT 1343.1000 1026.7500 1344.9000 1026.9000 ;
	    RECT 1307.1000 1025.2500 1344.9000 1026.7500 ;
	    RECT 1307.1000 1025.1000 1308.9000 1025.2500 ;
	    RECT 1314.3000 1025.1000 1316.1000 1025.2500 ;
	    RECT 1343.1000 1025.1000 1344.9000 1025.2500 ;
	    RECT 1489.5000 1026.7500 1491.3000 1026.9000 ;
	    RECT 1489.5000 1025.2500 1517.5500 1026.7500 ;
	    RECT 1489.5000 1025.1000 1491.3000 1025.2500 ;
	    RECT 1516.0500 1023.9000 1517.5500 1025.2500 ;
	    RECT 1520.7001 1025.1000 1522.5000 1026.9000 ;
	    RECT 1564.0500 1025.2500 1568.1000 1026.9000 ;
	    RECT 1564.8000 1025.1000 1568.1000 1025.2500 ;
	    RECT 1515.9000 1022.1000 1517.7001 1023.9000 ;
	    RECT 131.1000 1020.7500 132.9000 1020.9000 ;
	    RECT 135.9000 1020.7500 137.7000 1020.9000 ;
	    RECT 131.1000 1019.2500 137.7000 1020.7500 ;
	    RECT 131.1000 1019.1000 132.9000 1019.2500 ;
	    RECT 135.9000 1019.1000 137.7000 1019.2500 ;
	    RECT 143.1000 1020.7500 144.9000 1020.9000 ;
	    RECT 181.5000 1020.7500 183.3000 1020.9000 ;
	    RECT 143.1000 1019.2500 183.3000 1020.7500 ;
	    RECT 143.1000 1019.1000 144.9000 1019.2500 ;
	    RECT 181.5000 1019.1000 183.3000 1019.2500 ;
	    RECT 234.3000 1020.7500 236.1000 1020.9000 ;
	    RECT 251.1000 1020.7500 252.9000 1020.9000 ;
	    RECT 234.3000 1019.2500 252.9000 1020.7500 ;
	    RECT 234.3000 1019.1000 236.1000 1019.2500 ;
	    RECT 251.1000 1019.1000 252.9000 1019.2500 ;
	    RECT 263.1000 1020.7500 264.9000 1020.9000 ;
	    RECT 272.7000 1020.7500 274.5000 1020.9000 ;
	    RECT 263.1000 1019.2500 274.5000 1020.7500 ;
	    RECT 263.1000 1019.1000 264.9000 1019.2500 ;
	    RECT 272.7000 1019.1000 274.5000 1019.2500 ;
	    RECT 303.9000 1020.7500 305.7000 1020.9000 ;
	    RECT 335.1000 1020.7500 336.9000 1020.9000 ;
	    RECT 303.9000 1019.2500 336.9000 1020.7500 ;
	    RECT 303.9000 1019.1000 305.7000 1019.2500 ;
	    RECT 335.1000 1019.1000 336.9000 1019.2500 ;
	    RECT 459.9000 1020.7500 461.7000 1020.9000 ;
	    RECT 491.1000 1020.7500 492.9000 1020.9000 ;
	    RECT 459.9000 1019.2500 492.9000 1020.7500 ;
	    RECT 459.9000 1019.1000 461.7000 1019.2500 ;
	    RECT 491.1000 1019.1000 492.9000 1019.2500 ;
	    RECT 519.9000 1020.7500 521.7000 1020.9000 ;
	    RECT 524.7000 1020.7500 526.5000 1020.9000 ;
	    RECT 519.9000 1019.2500 526.5000 1020.7500 ;
	    RECT 519.9000 1019.1000 521.7000 1019.2500 ;
	    RECT 524.7000 1019.1000 526.5000 1019.2500 ;
	    RECT 630.3000 1020.7500 632.1000 1020.9000 ;
	    RECT 659.1000 1020.7500 660.9000 1020.9000 ;
	    RECT 630.3000 1019.2500 660.9000 1020.7500 ;
	    RECT 630.3000 1019.1000 632.1000 1019.2500 ;
	    RECT 659.1000 1019.1000 660.9000 1019.2500 ;
	    RECT 872.7000 1020.7500 874.5000 1020.9000 ;
	    RECT 887.1000 1020.7500 888.9000 1020.9000 ;
	    RECT 872.7000 1019.2500 888.9000 1020.7500 ;
	    RECT 872.7000 1019.1000 874.5000 1019.2500 ;
	    RECT 887.1000 1019.1000 888.9000 1019.2500 ;
	    RECT 920.7000 1020.7500 922.5000 1020.9000 ;
	    RECT 925.5000 1020.7500 927.3000 1020.9000 ;
	    RECT 920.7000 1019.2500 927.3000 1020.7500 ;
	    RECT 920.7000 1019.1000 922.5000 1019.2500 ;
	    RECT 925.5000 1019.1000 927.3000 1019.2500 ;
	    RECT 1035.9000 1020.7500 1037.7001 1020.9000 ;
	    RECT 1079.1000 1020.7500 1080.9000 1020.9000 ;
	    RECT 1035.9000 1019.2500 1080.9000 1020.7500 ;
	    RECT 1035.9000 1019.1000 1037.7001 1019.2500 ;
	    RECT 1079.1000 1019.1000 1080.9000 1019.2500 ;
	    RECT 167.1000 1014.7500 168.9000 1014.9000 ;
	    RECT 306.3000 1014.7500 308.1000 1014.9000 ;
	    RECT 167.1000 1013.2500 308.1000 1014.7500 ;
	    RECT 167.1000 1013.1000 168.9000 1013.2500 ;
	    RECT 306.3000 1013.1000 308.1000 1013.2500 ;
	    RECT 407.1000 1014.7500 408.9000 1014.9000 ;
	    RECT 510.3000 1014.7500 512.1000 1014.9000 ;
	    RECT 407.1000 1013.2500 512.1000 1014.7500 ;
	    RECT 407.1000 1013.1000 408.9000 1013.2500 ;
	    RECT 510.3000 1013.1000 512.1000 1013.2500 ;
	    RECT 567.9000 1014.7500 569.7000 1014.9000 ;
	    RECT 625.5000 1014.7500 627.3000 1014.9000 ;
	    RECT 567.9000 1013.2500 627.3000 1014.7500 ;
	    RECT 567.9000 1013.1000 569.7000 1013.2500 ;
	    RECT 625.5000 1013.1000 627.3000 1013.2500 ;
	    RECT 632.7000 1014.7500 634.5000 1014.9000 ;
	    RECT 639.9000 1014.7500 641.7000 1014.9000 ;
	    RECT 632.7000 1013.2500 641.7000 1014.7500 ;
	    RECT 632.7000 1013.1000 634.5000 1013.2500 ;
	    RECT 639.9000 1013.1000 641.7000 1013.2500 ;
	    RECT 747.9000 1014.7500 749.7000 1014.9000 ;
	    RECT 848.7000 1014.7500 850.5000 1014.9000 ;
	    RECT 747.9000 1013.2500 850.5000 1014.7500 ;
	    RECT 747.9000 1013.1000 749.7000 1013.2500 ;
	    RECT 848.7000 1013.1000 850.5000 1013.2500 ;
	    RECT 915.9000 1014.7500 917.7000 1014.9000 ;
	    RECT 968.7000 1014.7500 970.5000 1014.9000 ;
	    RECT 915.9000 1013.2500 970.5000 1014.7500 ;
	    RECT 915.9000 1013.1000 917.7000 1013.2500 ;
	    RECT 968.7000 1013.1000 970.5000 1013.2500 ;
	    RECT 1223.1000 1014.7500 1224.9000 1014.9000 ;
	    RECT 1290.3000 1014.7500 1292.1000 1014.9000 ;
	    RECT 1223.1000 1013.2500 1292.1000 1014.7500 ;
	    RECT 1223.1000 1013.1000 1224.9000 1013.2500 ;
	    RECT 1290.3000 1013.1000 1292.1000 1013.2500 ;
	    RECT 1424.7001 1014.7500 1426.5000 1014.9000 ;
	    RECT 1496.7001 1014.7500 1498.5000 1014.9000 ;
	    RECT 1556.7001 1014.7500 1558.5000 1014.9000 ;
	    RECT 1424.7001 1013.2500 1558.5000 1014.7500 ;
	    RECT 1424.7001 1013.1000 1426.5000 1013.2500 ;
	    RECT 1496.7001 1013.1000 1498.5000 1013.2500 ;
	    RECT 1556.7001 1013.1000 1558.5000 1013.2500 ;
	    RECT 291.9000 1008.7500 293.7000 1008.9000 ;
	    RECT 515.1000 1008.7500 516.9000 1008.9000 ;
	    RECT 291.9000 1007.2500 516.9000 1008.7500 ;
	    RECT 291.9000 1007.1000 293.7000 1007.2500 ;
	    RECT 515.1000 1007.1000 516.9000 1007.2500 ;
	    RECT 659.1000 1008.7500 660.9000 1008.9000 ;
	    RECT 671.1000 1008.7500 672.9000 1008.9000 ;
	    RECT 735.9000 1008.7500 737.7000 1008.9000 ;
	    RECT 659.1000 1007.2500 737.7000 1008.7500 ;
	    RECT 659.1000 1007.1000 660.9000 1007.2500 ;
	    RECT 671.1000 1007.1000 672.9000 1007.2500 ;
	    RECT 735.9000 1007.1000 737.7000 1007.2500 ;
	    RECT 824.7000 1008.7500 826.5000 1008.9000 ;
	    RECT 920.7000 1008.7500 922.5000 1008.9000 ;
	    RECT 824.7000 1007.2500 922.5000 1008.7500 ;
	    RECT 824.7000 1007.1000 826.5000 1007.2500 ;
	    RECT 920.7000 1007.1000 922.5000 1007.2500 ;
	    RECT 1038.3000 1008.7500 1040.1000 1008.9000 ;
	    RECT 1203.9000 1008.7500 1205.7001 1008.9000 ;
	    RECT 1038.3000 1007.2500 1205.7001 1008.7500 ;
	    RECT 1038.3000 1007.1000 1040.1000 1007.2500 ;
	    RECT 1203.9000 1007.1000 1205.7001 1007.2500 ;
	    RECT 1340.7001 1008.7500 1342.5000 1008.9000 ;
	    RECT 1431.9000 1008.7500 1433.7001 1008.9000 ;
	    RECT 1340.7001 1007.2500 1433.7001 1008.7500 ;
	    RECT 1340.7001 1007.1000 1342.5000 1007.2500 ;
	    RECT 1431.9000 1007.1000 1433.7001 1007.2500 ;
	    RECT 1491.9000 1008.7500 1493.7001 1008.9000 ;
	    RECT 1499.1000 1008.7500 1500.9000 1008.9000 ;
	    RECT 1491.9000 1007.2500 1500.9000 1008.7500 ;
	    RECT 1491.9000 1007.1000 1493.7001 1007.2500 ;
	    RECT 1499.1000 1007.1000 1500.9000 1007.2500 ;
	    RECT 1508.7001 1008.7500 1510.5000 1008.9000 ;
	    RECT 1520.7001 1008.7500 1522.5000 1008.9000 ;
	    RECT 1508.7001 1007.2500 1522.5000 1008.7500 ;
	    RECT 1508.7001 1007.1000 1510.5000 1007.2500 ;
	    RECT 1520.7001 1007.1000 1522.5000 1007.2500 ;
	    RECT 1535.1000 1008.7500 1536.9000 1008.9000 ;
	    RECT 1559.1000 1008.7500 1560.9000 1008.9000 ;
	    RECT 1535.1000 1007.2500 1560.9000 1008.7500 ;
	    RECT 1535.1000 1007.1000 1536.9000 1007.2500 ;
	    RECT 1559.1000 1007.1000 1560.9000 1007.2500 ;
	    RECT 171.9000 1002.7500 173.7000 1002.9000 ;
	    RECT 191.1000 1002.7500 192.9000 1002.9000 ;
	    RECT 171.9000 1001.2500 192.9000 1002.7500 ;
	    RECT 171.9000 1001.1000 173.7000 1001.2500 ;
	    RECT 191.1000 1001.1000 192.9000 1001.2500 ;
	    RECT 625.5000 1002.7500 627.3000 1002.9000 ;
	    RECT 642.3000 1002.7500 644.1000 1002.9000 ;
	    RECT 675.9000 1002.7500 677.7000 1002.9000 ;
	    RECT 625.5000 1001.2500 634.3500 1002.7500 ;
	    RECT 625.5000 1001.1000 627.3000 1001.2500 ;
	    RECT 632.8500 996.9000 634.3500 1001.2500 ;
	    RECT 642.3000 1001.2500 677.7000 1002.7500 ;
	    RECT 642.3000 1001.1000 644.1000 1001.2500 ;
	    RECT 675.9000 1001.1000 677.7000 1001.2500 ;
	    RECT 973.5000 1002.7500 975.3000 1002.9000 ;
	    RECT 1163.1000 1002.7500 1164.9000 1002.9000 ;
	    RECT 973.5000 1001.2500 1164.9000 1002.7500 ;
	    RECT 973.5000 1001.1000 975.3000 1001.2500 ;
	    RECT 1163.1000 1001.1000 1164.9000 1001.2500 ;
	    RECT 1201.5000 1002.7500 1203.3000 1002.9000 ;
	    RECT 1223.1000 1002.7500 1224.9000 1002.9000 ;
	    RECT 1201.5000 1001.2500 1224.9000 1002.7500 ;
	    RECT 1201.5000 1001.1000 1203.3000 1001.2500 ;
	    RECT 1223.1000 1001.1000 1224.9000 1001.2500 ;
	    RECT 1261.5000 1002.7500 1263.3000 1002.9000 ;
	    RECT 1292.7001 1002.7500 1294.5000 1002.9000 ;
	    RECT 1299.9000 1002.7500 1301.7001 1002.9000 ;
	    RECT 1261.5000 1001.2500 1301.7001 1002.7500 ;
	    RECT 1261.5000 1001.1000 1263.3000 1001.2500 ;
	    RECT 1292.7001 1001.1000 1294.5000 1001.2500 ;
	    RECT 1299.9000 1001.1000 1301.7001 1001.2500 ;
	    RECT 1388.7001 1002.7500 1390.5000 1002.9000 ;
	    RECT 1451.1000 1002.7500 1452.9000 1002.9000 ;
	    RECT 1388.7001 1001.2500 1452.9000 1002.7500 ;
	    RECT 1388.7001 1001.1000 1390.5000 1001.2500 ;
	    RECT 1451.1000 1001.1000 1452.9000 1001.2500 ;
	    RECT 1491.9000 1002.7500 1493.7001 1002.9000 ;
	    RECT 1511.1000 1002.7500 1512.9000 1002.9000 ;
	    RECT 1491.9000 1001.2500 1512.9000 1002.7500 ;
	    RECT 1491.9000 1001.1000 1493.7001 1001.2500 ;
	    RECT 1511.1000 1001.1000 1512.9000 1001.2500 ;
	    RECT 1515.9000 1002.7500 1517.7001 1002.9000 ;
	    RECT 1539.9000 1002.7500 1541.7001 1002.9000 ;
	    RECT 1515.9000 1001.2500 1541.7001 1002.7500 ;
	    RECT 1515.9000 1001.1000 1517.7001 1001.2500 ;
	    RECT 1539.9000 1001.1000 1541.7001 1001.2500 ;
	    RECT 222.3000 996.7500 224.1000 996.9000 ;
	    RECT 234.3000 996.7500 236.1000 996.9000 ;
	    RECT 222.3000 995.2500 236.1000 996.7500 ;
	    RECT 632.8500 995.2500 636.9000 996.9000 ;
	    RECT 222.3000 995.1000 224.1000 995.2500 ;
	    RECT 234.3000 995.1000 236.1000 995.2500 ;
	    RECT 633.6000 995.1000 636.9000 995.2500 ;
	    RECT 675.9000 996.7500 677.7000 996.9000 ;
	    RECT 707.1000 996.7500 708.9000 996.9000 ;
	    RECT 675.9000 995.2500 708.9000 996.7500 ;
	    RECT 675.9000 995.1000 677.7000 995.2500 ;
	    RECT 707.1000 995.1000 708.9000 995.2500 ;
	    RECT 757.5000 996.7500 759.3000 996.9000 ;
	    RECT 786.3000 996.7500 788.1000 996.9000 ;
	    RECT 757.5000 995.2500 788.1000 996.7500 ;
	    RECT 757.5000 995.1000 759.3000 995.2500 ;
	    RECT 786.3000 995.1000 788.1000 995.2500 ;
	    RECT 819.9000 996.7500 821.7000 996.9000 ;
	    RECT 839.1000 996.7500 840.9000 996.9000 ;
	    RECT 819.9000 995.2500 840.9000 996.7500 ;
	    RECT 819.9000 995.1000 821.7000 995.2500 ;
	    RECT 839.1000 995.1000 840.9000 995.2500 ;
	    RECT 1091.1000 996.7500 1092.9000 996.9000 ;
	    RECT 1232.7001 996.7500 1234.5000 996.9000 ;
	    RECT 1307.1000 996.7500 1308.9000 996.9000 ;
	    RECT 1328.7001 996.7500 1330.5000 996.9000 ;
	    RECT 1091.1000 995.2500 1330.5000 996.7500 ;
	    RECT 1091.1000 995.1000 1092.9000 995.2500 ;
	    RECT 1232.7001 995.1000 1234.5000 995.2500 ;
	    RECT 1307.1000 995.1000 1308.9000 995.2500 ;
	    RECT 1328.7001 995.1000 1330.5000 995.2500 ;
	    RECT 1350.3000 996.7500 1352.1000 996.9000 ;
	    RECT 1379.1000 996.7500 1380.9000 996.9000 ;
	    RECT 1383.9000 996.7500 1385.7001 996.9000 ;
	    RECT 1350.3000 995.2500 1385.7001 996.7500 ;
	    RECT 1350.3000 995.1000 1352.1000 995.2500 ;
	    RECT 1379.1000 995.1000 1380.9000 995.2500 ;
	    RECT 1383.9000 995.1000 1385.7001 995.2500 ;
	    RECT 1465.5000 996.7500 1467.3000 996.9000 ;
	    RECT 1491.9000 996.7500 1493.7001 996.9000 ;
	    RECT 1465.5000 995.2500 1493.7001 996.7500 ;
	    RECT 1465.5000 995.1000 1467.3000 995.2500 ;
	    RECT 1491.9000 995.1000 1493.7001 995.2500 ;
	    RECT 1525.5000 996.7500 1527.3000 996.9000 ;
	    RECT 1537.5000 996.7500 1539.3000 996.9000 ;
	    RECT 1525.5000 995.2500 1539.3000 996.7500 ;
	    RECT 1525.5000 995.1000 1527.3000 995.2500 ;
	    RECT 1537.5000 995.1000 1539.3000 995.2500 ;
	    RECT 135.9000 990.7500 137.7000 990.9000 ;
	    RECT 143.1000 990.7500 144.9000 990.9000 ;
	    RECT 135.9000 989.2500 144.9000 990.7500 ;
	    RECT 135.9000 989.1000 137.7000 989.2500 ;
	    RECT 143.1000 989.1000 144.9000 989.2500 ;
	    RECT 162.3000 990.7500 164.1000 990.9000 ;
	    RECT 188.7000 990.7500 190.5000 990.9000 ;
	    RECT 162.3000 989.2500 190.5000 990.7500 ;
	    RECT 162.3000 989.1000 164.1000 989.2500 ;
	    RECT 188.7000 989.1000 190.5000 989.2500 ;
	    RECT 217.5000 990.7500 219.3000 990.9000 ;
	    RECT 275.1000 990.7500 276.9000 990.9000 ;
	    RECT 217.5000 989.2500 276.9000 990.7500 ;
	    RECT 217.5000 989.1000 219.3000 989.2500 ;
	    RECT 275.1000 989.1000 276.9000 989.2500 ;
	    RECT 291.9000 990.7500 293.7000 990.9000 ;
	    RECT 301.5000 990.7500 303.3000 990.9000 ;
	    RECT 291.9000 989.2500 303.3000 990.7500 ;
	    RECT 291.9000 989.1000 293.7000 989.2500 ;
	    RECT 301.5000 989.1000 303.3000 989.2500 ;
	    RECT 623.1000 990.7500 624.9000 990.9000 ;
	    RECT 675.9000 990.7500 677.7000 990.9000 ;
	    RECT 623.1000 989.2500 677.7000 990.7500 ;
	    RECT 623.1000 989.1000 624.9000 989.2500 ;
	    RECT 675.9000 989.1000 677.7000 989.2500 ;
	    RECT 743.1000 990.7500 744.9000 990.9000 ;
	    RECT 781.5000 990.7500 783.3000 990.9000 ;
	    RECT 743.1000 989.2500 783.3000 990.7500 ;
	    RECT 743.1000 989.1000 744.9000 989.2500 ;
	    RECT 781.5000 989.1000 783.3000 989.2500 ;
	    RECT 908.7000 990.7500 910.5000 990.9000 ;
	    RECT 1026.3000 990.7500 1028.1000 990.9000 ;
	    RECT 908.7000 989.2500 1028.1000 990.7500 ;
	    RECT 908.7000 989.1000 910.5000 989.2500 ;
	    RECT 1026.3000 989.1000 1028.1000 989.2500 ;
	    RECT 1095.9000 990.7500 1097.7001 990.9000 ;
	    RECT 1110.3000 990.7500 1112.1000 990.9000 ;
	    RECT 1095.9000 989.2500 1112.1000 990.7500 ;
	    RECT 1095.9000 989.1000 1097.7001 989.2500 ;
	    RECT 1110.3000 989.1000 1112.1000 989.2500 ;
	    RECT 1129.5000 990.7500 1131.3000 990.9000 ;
	    RECT 1158.3000 990.7500 1160.1000 990.9000 ;
	    RECT 1129.5000 989.2500 1160.1000 990.7500 ;
	    RECT 1129.5000 989.1000 1131.3000 989.2500 ;
	    RECT 1158.3000 989.1000 1160.1000 989.2500 ;
	    RECT 1206.3000 990.7500 1208.1000 990.9000 ;
	    RECT 1220.7001 990.7500 1222.5000 990.9000 ;
	    RECT 1206.3000 989.2500 1222.5000 990.7500 ;
	    RECT 1206.3000 989.1000 1208.1000 989.2500 ;
	    RECT 1220.7001 989.1000 1222.5000 989.2500 ;
	    RECT 1395.9000 990.7500 1397.7001 990.9000 ;
	    RECT 1515.9000 990.7500 1517.7001 990.9000 ;
	    RECT 1395.9000 989.2500 1517.7001 990.7500 ;
	    RECT 1395.9000 989.1000 1397.7001 989.2500 ;
	    RECT 1515.9000 989.1000 1517.7001 989.2500 ;
	    RECT 1520.7001 990.7500 1522.5000 990.9000 ;
	    RECT 1547.1000 990.7500 1548.9000 990.9000 ;
	    RECT 1520.7001 989.2500 1548.9000 990.7500 ;
	    RECT 1520.7001 989.1000 1522.5000 989.2500 ;
	    RECT 1547.1000 989.1000 1548.9000 989.2500 ;
	    RECT 35.1000 984.7500 36.9000 984.9000 ;
	    RECT 135.9000 984.7500 137.7000 984.9000 ;
	    RECT 35.1000 983.2500 137.7000 984.7500 ;
	    RECT 35.1000 983.1000 36.9000 983.2500 ;
	    RECT 135.9000 983.1000 137.7000 983.2500 ;
	    RECT 265.5000 984.7500 267.3000 984.9000 ;
	    RECT 272.7000 984.7500 274.5000 984.9000 ;
	    RECT 265.5000 983.2500 274.5000 984.7500 ;
	    RECT 265.5000 983.1000 267.3000 983.2500 ;
	    RECT 272.7000 983.1000 274.5000 983.2500 ;
	    RECT 397.5000 984.7500 399.3000 984.9000 ;
	    RECT 524.7000 984.7500 526.5000 984.9000 ;
	    RECT 539.1000 984.7500 540.9000 984.9000 ;
	    RECT 589.5000 984.7500 591.3000 984.9000 ;
	    RECT 620.7000 984.7500 622.5000 984.9000 ;
	    RECT 397.5000 983.2500 622.5000 984.7500 ;
	    RECT 397.5000 983.1000 399.3000 983.2500 ;
	    RECT 524.7000 983.1000 526.5000 983.2500 ;
	    RECT 539.1000 983.1000 540.9000 983.2500 ;
	    RECT 589.5000 983.1000 591.3000 983.2500 ;
	    RECT 620.7000 983.1000 622.5000 983.2500 ;
	    RECT 635.1000 984.7500 636.9000 984.9000 ;
	    RECT 661.5000 984.7500 663.3000 984.9000 ;
	    RECT 635.1000 983.2500 663.3000 984.7500 ;
	    RECT 635.1000 983.1000 636.9000 983.2500 ;
	    RECT 661.5000 983.1000 663.3000 983.2500 ;
	    RECT 843.9000 984.7500 845.7000 984.9000 ;
	    RECT 951.9000 984.7500 953.7000 984.9000 ;
	    RECT 843.9000 983.2500 953.7000 984.7500 ;
	    RECT 843.9000 983.1000 845.7000 983.2500 ;
	    RECT 951.9000 983.1000 953.7000 983.2500 ;
	    RECT 1031.1000 984.7500 1032.9000 984.9000 ;
	    RECT 1062.3000 984.7500 1064.1000 984.9000 ;
	    RECT 1031.1000 983.2500 1064.1000 984.7500 ;
	    RECT 1031.1000 983.1000 1032.9000 983.2500 ;
	    RECT 1062.3000 983.1000 1064.1000 983.2500 ;
	    RECT 1088.7001 984.7500 1090.5000 984.9000 ;
	    RECT 1134.3000 984.7500 1136.1000 984.9000 ;
	    RECT 1088.7001 983.2500 1136.1000 984.7500 ;
	    RECT 1088.7001 983.1000 1090.5000 983.2500 ;
	    RECT 1134.3000 983.1000 1136.1000 983.2500 ;
	    RECT 1381.5000 984.7500 1383.3000 984.9000 ;
	    RECT 1391.1000 984.7500 1392.9000 984.9000 ;
	    RECT 1381.5000 983.2500 1392.9000 984.7500 ;
	    RECT 1381.5000 983.1000 1383.3000 983.2500 ;
	    RECT 1391.1000 983.1000 1392.9000 983.2500 ;
	    RECT 162.3000 978.7500 164.1000 978.9000 ;
	    RECT 253.5000 978.7500 255.3000 978.9000 ;
	    RECT 162.3000 977.2500 255.3000 978.7500 ;
	    RECT 162.3000 977.1000 164.1000 977.2500 ;
	    RECT 253.5000 977.1000 255.3000 977.2500 ;
	    RECT 258.3000 978.7500 260.1000 978.9000 ;
	    RECT 315.9000 978.7500 317.7000 978.9000 ;
	    RECT 258.3000 977.2500 317.7000 978.7500 ;
	    RECT 258.3000 977.1000 260.1000 977.2500 ;
	    RECT 315.9000 977.1000 317.7000 977.2500 ;
	    RECT 642.3000 978.7500 644.1000 978.9000 ;
	    RECT 668.7000 978.7500 670.5000 978.9000 ;
	    RECT 642.3000 977.2500 670.5000 978.7500 ;
	    RECT 642.3000 977.1000 644.1000 977.2500 ;
	    RECT 668.7000 977.1000 670.5000 977.2500 ;
	    RECT 817.5000 978.7500 819.3000 978.9000 ;
	    RECT 836.7000 978.7500 838.5000 978.9000 ;
	    RECT 865.5000 978.7500 867.3000 978.9000 ;
	    RECT 817.5000 977.2500 867.3000 978.7500 ;
	    RECT 817.5000 977.1000 819.3000 977.2500 ;
	    RECT 836.7000 977.1000 838.5000 977.2500 ;
	    RECT 865.5000 977.1000 867.3000 977.2500 ;
	    RECT 918.3000 978.7500 920.1000 978.9000 ;
	    RECT 930.3000 978.7500 932.1000 978.9000 ;
	    RECT 918.3000 977.2500 932.1000 978.7500 ;
	    RECT 918.3000 977.1000 920.1000 977.2500 ;
	    RECT 930.3000 977.1000 932.1000 977.2500 ;
	    RECT 949.5000 978.7500 951.3000 978.9000 ;
	    RECT 992.7000 978.7500 994.5000 978.9000 ;
	    RECT 949.5000 977.2500 994.5000 978.7500 ;
	    RECT 949.5000 977.1000 951.3000 977.2500 ;
	    RECT 992.7000 977.1000 994.5000 977.2500 ;
	    RECT 1122.3000 978.7500 1124.1000 978.9000 ;
	    RECT 1131.9000 978.7500 1133.7001 978.9000 ;
	    RECT 1122.3000 977.2500 1133.7001 978.7500 ;
	    RECT 1122.3000 977.1000 1124.1000 977.2500 ;
	    RECT 1131.9000 977.1000 1133.7001 977.2500 ;
	    RECT 1287.9000 978.7500 1289.7001 978.9000 ;
	    RECT 1302.3000 978.7500 1304.1000 978.9000 ;
	    RECT 1287.9000 977.2500 1304.1000 978.7500 ;
	    RECT 1287.9000 977.1000 1289.7001 977.2500 ;
	    RECT 1302.3000 977.1000 1304.1000 977.2500 ;
	    RECT 1321.5000 978.7500 1323.3000 978.9000 ;
	    RECT 1333.5000 978.7500 1335.3000 978.9000 ;
	    RECT 1321.5000 977.2500 1335.3000 978.7500 ;
	    RECT 1321.5000 977.1000 1323.3000 977.2500 ;
	    RECT 1333.5000 977.1000 1335.3000 977.2500 ;
	    RECT 1410.3000 978.7500 1412.1000 978.9000 ;
	    RECT 1465.5000 978.7500 1467.3000 978.9000 ;
	    RECT 1410.3000 977.2500 1467.3000 978.7500 ;
	    RECT 1410.3000 977.1000 1412.1000 977.2500 ;
	    RECT 1465.5000 977.1000 1467.3000 977.2500 ;
	    RECT 219.9000 972.7500 221.7000 972.9000 ;
	    RECT 248.7000 972.7500 250.5000 972.9000 ;
	    RECT 219.9000 971.2500 250.5000 972.7500 ;
	    RECT 219.9000 971.1000 221.7000 971.2500 ;
	    RECT 248.7000 971.1000 250.5000 971.2500 ;
	    RECT 452.7000 972.7500 454.5000 972.9000 ;
	    RECT 517.5000 972.7500 519.3000 972.9000 ;
	    RECT 452.7000 971.2500 519.3000 972.7500 ;
	    RECT 452.7000 971.1000 454.5000 971.2500 ;
	    RECT 517.5000 971.1000 519.3000 971.2500 ;
	    RECT 954.3000 972.7500 956.1000 972.9000 ;
	    RECT 1028.7001 972.7500 1030.5000 972.9000 ;
	    RECT 954.3000 971.2500 1030.5000 972.7500 ;
	    RECT 954.3000 971.1000 956.1000 971.2500 ;
	    RECT 1028.7001 971.1000 1030.5000 971.2500 ;
	    RECT 1391.1000 972.7500 1392.9000 972.9000 ;
	    RECT 1439.1000 972.7500 1440.9000 972.9000 ;
	    RECT 1391.1000 971.2500 1440.9000 972.7500 ;
	    RECT 1391.1000 971.1000 1392.9000 971.2500 ;
	    RECT 1439.1000 971.1000 1440.9000 971.2500 ;
	    RECT 1508.7001 972.7500 1510.5000 972.9000 ;
	    RECT 1539.9000 972.7500 1541.7001 972.9000 ;
	    RECT 1508.7001 971.2500 1541.7001 972.7500 ;
	    RECT 1508.7001 971.1000 1510.5000 971.2500 ;
	    RECT 1539.9000 971.1000 1541.7001 971.2500 ;
	    RECT 152.7000 966.7500 154.5000 966.9000 ;
	    RECT 258.3000 966.7500 260.1000 966.9000 ;
	    RECT 152.7000 965.2500 260.1000 966.7500 ;
	    RECT 152.7000 965.1000 154.5000 965.2500 ;
	    RECT 258.3000 965.1000 260.1000 965.2500 ;
	    RECT 282.3000 966.7500 284.1000 966.9000 ;
	    RECT 313.5000 966.7500 315.3000 966.9000 ;
	    RECT 282.3000 965.2500 315.3000 966.7500 ;
	    RECT 282.3000 965.1000 284.1000 965.2500 ;
	    RECT 313.5000 965.1000 315.3000 965.2500 ;
	    RECT 507.9000 966.7500 509.7000 966.9000 ;
	    RECT 618.3000 966.7500 620.1000 966.9000 ;
	    RECT 507.9000 965.2500 620.1000 966.7500 ;
	    RECT 507.9000 965.1000 509.7000 965.2500 ;
	    RECT 618.3000 965.1000 620.1000 965.2500 ;
	    RECT 675.9000 966.7500 677.7000 966.9000 ;
	    RECT 683.1000 966.7500 684.9000 966.9000 ;
	    RECT 675.9000 965.2500 684.9000 966.7500 ;
	    RECT 675.9000 965.1000 677.7000 965.2500 ;
	    RECT 683.1000 965.1000 684.9000 965.2500 ;
	    RECT 745.5000 966.7500 747.3000 966.9000 ;
	    RECT 759.9000 966.7500 761.7000 966.9000 ;
	    RECT 745.5000 965.2500 761.7000 966.7500 ;
	    RECT 745.5000 965.1000 747.3000 965.2500 ;
	    RECT 759.9000 965.1000 761.7000 965.2500 ;
	    RECT 786.3000 966.7500 788.1000 966.9000 ;
	    RECT 867.9000 966.7500 869.7000 966.9000 ;
	    RECT 786.3000 965.2500 869.7000 966.7500 ;
	    RECT 786.3000 965.1000 788.1000 965.2500 ;
	    RECT 867.9000 965.1000 869.7000 965.2500 ;
	    RECT 899.1000 966.7500 900.9000 966.9000 ;
	    RECT 954.3000 966.7500 956.1000 966.9000 ;
	    RECT 899.1000 965.2500 956.1000 966.7500 ;
	    RECT 899.1000 965.1000 900.9000 965.2500 ;
	    RECT 954.3000 965.1000 956.1000 965.2500 ;
	    RECT 1086.3000 966.7500 1088.1000 966.9000 ;
	    RECT 1115.1000 966.7500 1116.9000 966.9000 ;
	    RECT 1086.3000 965.2500 1116.9000 966.7500 ;
	    RECT 1086.3000 965.1000 1088.1000 965.2500 ;
	    RECT 1115.1000 965.1000 1116.9000 965.2500 ;
	    RECT 1129.5000 966.7500 1131.3000 966.9000 ;
	    RECT 1134.3000 966.7500 1136.1000 966.9000 ;
	    RECT 1129.5000 965.2500 1136.1000 966.7500 ;
	    RECT 1129.5000 965.1000 1131.3000 965.2500 ;
	    RECT 1134.3000 965.1000 1136.1000 965.2500 ;
	    RECT 1199.1000 966.7500 1200.9000 966.9000 ;
	    RECT 1227.9000 966.7500 1229.7001 966.9000 ;
	    RECT 1199.1000 965.2500 1229.7001 966.7500 ;
	    RECT 1199.1000 965.1000 1200.9000 965.2500 ;
	    RECT 1227.9000 965.1000 1229.7001 965.2500 ;
	    RECT 1271.1000 966.7500 1272.9000 966.9000 ;
	    RECT 1352.7001 966.7500 1354.5000 966.9000 ;
	    RECT 1271.1000 965.2500 1354.5000 966.7500 ;
	    RECT 1271.1000 965.1000 1272.9000 965.2500 ;
	    RECT 1352.7001 965.1000 1354.5000 965.2500 ;
	    RECT 1499.1000 966.7500 1500.9000 966.9000 ;
	    RECT 1523.1000 966.7500 1524.9000 966.9000 ;
	    RECT 1499.1000 965.2500 1524.9000 966.7500 ;
	    RECT 1499.1000 965.1000 1500.9000 965.2500 ;
	    RECT 1523.1000 965.1000 1524.9000 965.2500 ;
	    RECT 95.1000 960.7500 96.9000 960.9000 ;
	    RECT 123.9000 960.7500 125.7000 960.9000 ;
	    RECT 95.1000 959.2500 125.7000 960.7500 ;
	    RECT 95.1000 959.1000 96.9000 959.2500 ;
	    RECT 123.9000 959.1000 125.7000 959.2500 ;
	    RECT 131.1000 960.7500 132.9000 960.9000 ;
	    RECT 174.3000 960.7500 176.1000 960.9000 ;
	    RECT 131.1000 959.2500 176.1000 960.7500 ;
	    RECT 131.1000 959.1000 132.9000 959.2500 ;
	    RECT 174.3000 959.1000 176.1000 959.2500 ;
	    RECT 349.5000 960.7500 351.3000 960.9000 ;
	    RECT 371.1000 960.7500 372.9000 960.9000 ;
	    RECT 349.5000 959.2500 372.9000 960.7500 ;
	    RECT 349.5000 959.1000 351.3000 959.2500 ;
	    RECT 371.1000 959.1000 372.9000 959.2500 ;
	    RECT 385.5000 960.7500 387.3000 960.9000 ;
	    RECT 392.7000 960.7500 394.5000 960.9000 ;
	    RECT 419.1000 960.7500 420.9000 960.9000 ;
	    RECT 431.1000 960.7500 432.9000 960.9000 ;
	    RECT 455.1000 960.7500 456.9000 960.9000 ;
	    RECT 385.5000 959.2500 456.9000 960.7500 ;
	    RECT 385.5000 959.1000 387.3000 959.2500 ;
	    RECT 392.7000 959.1000 394.5000 959.2500 ;
	    RECT 419.1000 959.1000 420.9000 959.2500 ;
	    RECT 431.1000 959.1000 432.9000 959.2500 ;
	    RECT 455.1000 959.1000 456.9000 959.2500 ;
	    RECT 524.7000 960.7500 526.5000 960.9000 ;
	    RECT 536.7000 960.7500 538.5000 960.9000 ;
	    RECT 524.7000 959.2500 538.5000 960.7500 ;
	    RECT 524.7000 959.1000 526.5000 959.2500 ;
	    RECT 536.7000 959.1000 538.5000 959.2500 ;
	    RECT 591.9000 960.7500 593.7000 960.9000 ;
	    RECT 601.5000 960.7500 603.3000 960.9000 ;
	    RECT 591.9000 959.2500 603.3000 960.7500 ;
	    RECT 591.9000 959.1000 593.7000 959.2500 ;
	    RECT 601.5000 959.1000 603.3000 959.2500 ;
	    RECT 707.1000 960.7500 708.9000 960.9000 ;
	    RECT 803.1000 960.7500 804.9000 960.9000 ;
	    RECT 707.1000 959.2500 804.9000 960.7500 ;
	    RECT 707.1000 959.1000 708.9000 959.2500 ;
	    RECT 803.1000 959.1000 804.9000 959.2500 ;
	    RECT 817.5000 960.7500 819.3000 960.9000 ;
	    RECT 836.7000 960.7500 838.5000 960.9000 ;
	    RECT 817.5000 959.2500 838.5000 960.7500 ;
	    RECT 817.5000 959.1000 819.3000 959.2500 ;
	    RECT 836.7000 959.1000 838.5000 959.2500 ;
	    RECT 855.9000 960.7500 857.7000 960.9000 ;
	    RECT 863.1000 960.7500 864.9000 960.9000 ;
	    RECT 855.9000 959.2500 864.9000 960.7500 ;
	    RECT 855.9000 959.1000 857.7000 959.2500 ;
	    RECT 863.1000 959.1000 864.9000 959.2500 ;
	    RECT 906.3000 960.7500 908.1000 960.9000 ;
	    RECT 973.5000 960.7500 975.3000 960.9000 ;
	    RECT 906.3000 959.2500 975.3000 960.7500 ;
	    RECT 906.3000 959.1000 908.1000 959.2500 ;
	    RECT 973.5000 959.1000 975.3000 959.2500 ;
	    RECT 987.9000 960.7500 989.7000 960.9000 ;
	    RECT 1023.9000 960.7500 1025.7001 960.9000 ;
	    RECT 987.9000 959.2500 1025.7001 960.7500 ;
	    RECT 987.9000 959.1000 989.7000 959.2500 ;
	    RECT 1023.9000 959.1000 1025.7001 959.2500 ;
	    RECT 1263.9000 960.7500 1265.7001 960.9000 ;
	    RECT 1302.3000 960.7500 1304.1000 960.9000 ;
	    RECT 1321.5000 960.7500 1323.3000 960.9000 ;
	    RECT 1263.9000 959.2500 1323.3000 960.7500 ;
	    RECT 1263.9000 959.1000 1265.7001 959.2500 ;
	    RECT 1302.3000 959.1000 1304.1000 959.2500 ;
	    RECT 1321.5000 959.1000 1323.3000 959.2500 ;
	    RECT 1513.5000 960.7500 1515.3000 960.9000 ;
	    RECT 1518.3000 960.7500 1520.1000 960.9000 ;
	    RECT 1513.5000 959.2500 1520.1000 960.7500 ;
	    RECT 1513.5000 959.1000 1515.3000 959.2500 ;
	    RECT 1518.3000 959.1000 1520.1000 959.2500 ;
	    RECT 1525.5000 960.7500 1527.3000 960.9000 ;
	    RECT 1549.5000 960.7500 1551.3000 960.9000 ;
	    RECT 1525.5000 959.2500 1551.3000 960.7500 ;
	    RECT 1525.5000 959.1000 1527.3000 959.2500 ;
	    RECT 1549.5000 959.1000 1551.3000 959.2500 ;
	    RECT 123.9000 954.7500 125.7000 954.9000 ;
	    RECT 145.5000 954.7500 147.3000 954.9000 ;
	    RECT 123.9000 953.2500 147.3000 954.7500 ;
	    RECT 123.9000 953.1000 125.7000 953.2500 ;
	    RECT 145.5000 953.1000 147.3000 953.2500 ;
	    RECT 198.3000 954.7500 200.1000 954.9000 ;
	    RECT 222.3000 954.7500 224.1000 954.9000 ;
	    RECT 198.3000 953.2500 224.1000 954.7500 ;
	    RECT 198.3000 953.1000 200.1000 953.2500 ;
	    RECT 222.3000 953.1000 224.1000 953.2500 ;
	    RECT 255.9000 954.7500 257.7000 954.9000 ;
	    RECT 284.7000 954.7500 286.5000 954.9000 ;
	    RECT 255.9000 953.2500 286.5000 954.7500 ;
	    RECT 255.9000 953.1000 257.7000 953.2500 ;
	    RECT 284.7000 953.1000 286.5000 953.2500 ;
	    RECT 373.5000 954.7500 375.3000 954.9000 ;
	    RECT 380.7000 954.7500 382.5000 954.9000 ;
	    RECT 392.7000 954.7500 394.5000 954.9000 ;
	    RECT 433.5000 954.7500 435.3000 954.9000 ;
	    RECT 373.5000 953.2500 435.3000 954.7500 ;
	    RECT 373.5000 953.1000 375.3000 953.2500 ;
	    RECT 380.7000 953.1000 382.5000 953.2500 ;
	    RECT 392.7000 953.1000 394.5000 953.2500 ;
	    RECT 433.5000 953.1000 435.3000 953.2500 ;
	    RECT 531.9000 954.7500 533.7000 954.9000 ;
	    RECT 594.3000 954.7500 596.1000 954.9000 ;
	    RECT 606.3000 954.7500 608.1000 954.9000 ;
	    RECT 531.9000 953.2500 608.1000 954.7500 ;
	    RECT 531.9000 953.1000 533.7000 953.2500 ;
	    RECT 594.3000 953.1000 596.1000 953.2500 ;
	    RECT 606.3000 953.1000 608.1000 953.2500 ;
	    RECT 620.7000 954.7500 622.5000 954.9000 ;
	    RECT 675.9000 954.7500 677.7000 954.9000 ;
	    RECT 620.7000 953.2500 677.7000 954.7500 ;
	    RECT 620.7000 953.1000 622.5000 953.2500 ;
	    RECT 675.9000 953.1000 677.7000 953.2500 ;
	    RECT 683.1000 954.7500 684.9000 954.9000 ;
	    RECT 709.5000 954.7500 711.3000 954.9000 ;
	    RECT 767.1000 954.7500 768.9000 954.9000 ;
	    RECT 683.1000 953.2500 768.9000 954.7500 ;
	    RECT 683.1000 953.1000 684.9000 953.2500 ;
	    RECT 709.5000 953.1000 711.3000 953.2500 ;
	    RECT 767.1000 953.1000 768.9000 953.2500 ;
	    RECT 771.9000 954.7500 773.7000 954.9000 ;
	    RECT 793.5000 954.7500 795.3000 954.9000 ;
	    RECT 771.9000 953.2500 795.3000 954.7500 ;
	    RECT 771.9000 953.1000 773.7000 953.2500 ;
	    RECT 793.5000 953.1000 795.3000 953.2500 ;
	    RECT 824.7000 954.7500 826.5000 954.9000 ;
	    RECT 846.3000 954.7500 848.1000 954.9000 ;
	    RECT 824.7000 953.2500 848.1000 954.7500 ;
	    RECT 824.7000 953.1000 826.5000 953.2500 ;
	    RECT 846.3000 953.1000 848.1000 953.2500 ;
	    RECT 853.5000 954.7500 855.3000 954.9000 ;
	    RECT 899.1000 954.7500 900.9000 954.9000 ;
	    RECT 853.5000 953.2500 900.9000 954.7500 ;
	    RECT 853.5000 953.1000 855.3000 953.2500 ;
	    RECT 899.1000 953.1000 900.9000 953.2500 ;
	    RECT 1551.9000 954.7500 1553.7001 954.9000 ;
	    RECT 1556.7001 954.7500 1558.5000 954.9000 ;
	    RECT 1551.9000 953.2500 1558.5000 954.7500 ;
	    RECT 1551.9000 953.1000 1553.7001 953.2500 ;
	    RECT 1556.7001 953.1000 1558.5000 953.2500 ;
	    RECT 66.3000 948.7500 68.1000 948.9000 ;
	    RECT 133.5000 948.7500 135.3000 948.9000 ;
	    RECT 176.7000 948.7500 178.5000 948.9000 ;
	    RECT 66.3000 947.2500 178.5000 948.7500 ;
	    RECT 66.3000 947.1000 68.1000 947.2500 ;
	    RECT 133.5000 947.1000 135.3000 947.2500 ;
	    RECT 176.7000 947.1000 178.5000 947.2500 ;
	    RECT 279.9000 948.7500 281.7000 948.9000 ;
	    RECT 296.7000 948.7500 298.5000 948.9000 ;
	    RECT 301.5000 948.7500 303.3000 948.9000 ;
	    RECT 387.9000 948.7500 389.7000 948.9000 ;
	    RECT 402.3000 948.7500 404.1000 948.9000 ;
	    RECT 452.7000 948.7500 454.5000 948.9000 ;
	    RECT 279.9000 947.2500 454.5000 948.7500 ;
	    RECT 279.9000 947.1000 281.7000 947.2500 ;
	    RECT 296.7000 947.1000 298.5000 947.2500 ;
	    RECT 301.5000 947.1000 303.3000 947.2500 ;
	    RECT 387.9000 947.1000 389.7000 947.2500 ;
	    RECT 402.3000 947.1000 404.1000 947.2500 ;
	    RECT 452.7000 947.1000 454.5000 947.2500 ;
	    RECT 639.9000 948.7500 641.7000 948.9000 ;
	    RECT 680.7000 948.7500 682.5000 948.9000 ;
	    RECT 711.9000 948.7500 713.7000 948.9000 ;
	    RECT 771.9000 948.7500 773.7000 948.9000 ;
	    RECT 639.9000 947.2500 773.7000 948.7500 ;
	    RECT 639.9000 947.1000 641.7000 947.2500 ;
	    RECT 680.7000 947.1000 682.5000 947.2500 ;
	    RECT 711.9000 947.1000 713.7000 947.2500 ;
	    RECT 771.9000 947.1000 773.7000 947.2500 ;
	    RECT 795.9000 948.7500 797.7000 948.9000 ;
	    RECT 815.1000 948.7500 816.9000 948.9000 ;
	    RECT 795.9000 947.2500 816.9000 948.7500 ;
	    RECT 795.9000 947.1000 797.7000 947.2500 ;
	    RECT 815.1000 947.1000 816.9000 947.2500 ;
	    RECT 829.5000 948.7500 831.3000 948.9000 ;
	    RECT 839.1000 948.7500 840.9000 948.9000 ;
	    RECT 829.5000 947.2500 840.9000 948.7500 ;
	    RECT 829.5000 947.1000 831.3000 947.2500 ;
	    RECT 839.1000 947.1000 840.9000 947.2500 ;
	    RECT 846.3000 948.7500 848.1000 948.9000 ;
	    RECT 894.3000 948.7500 896.1000 948.9000 ;
	    RECT 846.3000 947.2500 896.1000 948.7500 ;
	    RECT 846.3000 947.1000 848.1000 947.2500 ;
	    RECT 894.3000 947.1000 896.1000 947.2500 ;
	    RECT 1119.9000 948.7500 1121.7001 948.9000 ;
	    RECT 1129.5000 948.7500 1131.3000 948.9000 ;
	    RECT 1119.9000 947.2500 1131.3000 948.7500 ;
	    RECT 1119.9000 947.1000 1121.7001 947.2500 ;
	    RECT 1129.5000 947.1000 1131.3000 947.2500 ;
	    RECT 1165.5000 948.7500 1167.3000 948.9000 ;
	    RECT 1261.5000 948.7500 1263.3000 948.9000 ;
	    RECT 1165.5000 947.2500 1263.3000 948.7500 ;
	    RECT 1165.5000 947.1000 1167.3000 947.2500 ;
	    RECT 1261.5000 947.1000 1263.3000 947.2500 ;
	    RECT 1307.1000 948.7500 1308.9000 948.9000 ;
	    RECT 1321.5000 948.7500 1323.3000 948.9000 ;
	    RECT 1307.1000 947.2500 1323.3000 948.7500 ;
	    RECT 1307.1000 947.1000 1308.9000 947.2500 ;
	    RECT 1321.5000 947.1000 1323.3000 947.2500 ;
	    RECT 1383.9000 948.7500 1385.7001 948.9000 ;
	    RECT 1410.3000 948.7500 1412.1000 948.9000 ;
	    RECT 1383.9000 947.2500 1412.1000 948.7500 ;
	    RECT 1383.9000 947.1000 1385.7001 947.2500 ;
	    RECT 1410.3000 947.1000 1412.1000 947.2500 ;
	    RECT 1453.5000 948.7500 1455.3000 948.9000 ;
	    RECT 1520.7001 948.7500 1522.5000 948.9000 ;
	    RECT 1453.5000 947.2500 1522.5000 948.7500 ;
	    RECT 1453.5000 947.1000 1455.3000 947.2500 ;
	    RECT 1520.7001 947.1000 1522.5000 947.2500 ;
	    RECT 1542.3000 948.7500 1544.1000 948.9000 ;
	    RECT 1551.9000 948.7500 1553.7001 948.9000 ;
	    RECT 1542.3000 947.2500 1553.7001 948.7500 ;
	    RECT 1542.3000 947.1000 1544.1000 947.2500 ;
	    RECT 1551.9000 947.1000 1553.7001 947.2500 ;
	    RECT 27.9000 942.7500 29.7000 942.9000 ;
	    RECT 37.5000 942.7500 39.3000 942.9000 ;
	    RECT 27.9000 941.2500 39.3000 942.7500 ;
	    RECT 27.9000 941.1000 29.7000 941.2500 ;
	    RECT 37.5000 941.1000 39.3000 941.2500 ;
	    RECT 71.1000 942.7500 72.9000 942.9000 ;
	    RECT 102.3000 942.7500 104.1000 942.9000 ;
	    RECT 71.1000 941.2500 104.1000 942.7500 ;
	    RECT 71.1000 941.1000 72.9000 941.2500 ;
	    RECT 102.3000 941.1000 104.1000 941.2500 ;
	    RECT 215.1000 942.7500 216.9000 942.9000 ;
	    RECT 248.7000 942.7500 250.5000 942.9000 ;
	    RECT 291.9000 942.7500 293.7000 942.9000 ;
	    RECT 308.7000 942.7500 310.5000 942.9000 ;
	    RECT 215.1000 941.2500 310.5000 942.7500 ;
	    RECT 215.1000 941.1000 216.9000 941.2500 ;
	    RECT 248.7000 941.1000 250.5000 941.2500 ;
	    RECT 291.9000 941.1000 293.7000 941.2500 ;
	    RECT 308.7000 941.1000 310.5000 941.2500 ;
	    RECT 313.5000 942.7500 315.3000 942.9000 ;
	    RECT 320.7000 942.7500 322.5000 942.9000 ;
	    RECT 313.5000 941.2500 322.5000 942.7500 ;
	    RECT 313.5000 941.1000 315.3000 941.2500 ;
	    RECT 320.7000 941.1000 322.5000 941.2500 ;
	    RECT 596.7000 942.7500 598.5000 942.9000 ;
	    RECT 615.9000 942.7500 617.7000 942.9000 ;
	    RECT 596.7000 941.2500 617.7000 942.7500 ;
	    RECT 596.7000 941.1000 598.5000 941.2500 ;
	    RECT 615.9000 941.1000 617.7000 941.2500 ;
	    RECT 678.3000 942.7500 680.1000 942.9000 ;
	    RECT 683.1000 942.7500 684.9000 942.9000 ;
	    RECT 678.3000 941.2500 684.9000 942.7500 ;
	    RECT 678.3000 941.1000 680.1000 941.2500 ;
	    RECT 683.1000 941.1000 684.9000 941.2500 ;
	    RECT 759.9000 942.7500 761.7000 942.9000 ;
	    RECT 798.3000 942.7500 800.1000 942.9000 ;
	    RECT 759.9000 941.2500 800.1000 942.7500 ;
	    RECT 759.9000 941.1000 761.7000 941.2500 ;
	    RECT 798.3000 941.1000 800.1000 941.2500 ;
	    RECT 834.3000 942.7500 836.1000 942.9000 ;
	    RECT 863.1000 942.7500 864.9000 942.9000 ;
	    RECT 834.3000 941.2500 864.9000 942.7500 ;
	    RECT 834.3000 941.1000 836.1000 941.2500 ;
	    RECT 863.1000 941.1000 864.9000 941.2500 ;
	    RECT 889.5000 942.7500 891.3000 942.9000 ;
	    RECT 913.5000 942.7500 915.3000 942.9000 ;
	    RECT 889.5000 941.2500 915.3000 942.7500 ;
	    RECT 889.5000 941.1000 891.3000 941.2500 ;
	    RECT 913.5000 941.1000 915.3000 941.2500 ;
	    RECT 939.9000 942.7500 941.7000 942.9000 ;
	    RECT 959.1000 942.7500 960.9000 942.9000 ;
	    RECT 939.9000 941.2500 960.9000 942.7500 ;
	    RECT 939.9000 941.1000 941.7000 941.2500 ;
	    RECT 959.1000 941.1000 960.9000 941.2500 ;
	    RECT 999.9000 942.7500 1001.7000 942.9000 ;
	    RECT 1004.7000 942.7500 1006.5000 942.9000 ;
	    RECT 999.9000 941.2500 1006.5000 942.7500 ;
	    RECT 999.9000 941.1000 1001.7000 941.2500 ;
	    RECT 1004.7000 941.1000 1006.5000 941.2500 ;
	    RECT 1103.1000 942.7500 1104.9000 942.9000 ;
	    RECT 1119.9000 942.7500 1121.7001 942.9000 ;
	    RECT 1103.1000 941.2500 1121.7001 942.7500 ;
	    RECT 1103.1000 941.1000 1104.9000 941.2500 ;
	    RECT 1119.9000 941.1000 1121.7001 941.2500 ;
	    RECT 1321.5000 942.7500 1323.3000 942.9000 ;
	    RECT 1333.5000 942.7500 1335.3000 942.9000 ;
	    RECT 1321.5000 941.2500 1335.3000 942.7500 ;
	    RECT 1321.5000 941.1000 1323.3000 941.2500 ;
	    RECT 1333.5000 941.1000 1335.3000 941.2500 ;
	    RECT 231.9000 936.7500 233.7000 936.9000 ;
	    RECT 253.5000 936.7500 255.3000 936.9000 ;
	    RECT 231.9000 935.2500 255.3000 936.7500 ;
	    RECT 231.9000 935.1000 233.7000 935.2500 ;
	    RECT 253.5000 935.1000 255.3000 935.2500 ;
	    RECT 284.7000 936.7500 286.5000 936.9000 ;
	    RECT 291.9000 936.7500 293.7000 936.9000 ;
	    RECT 284.7000 935.2500 293.7000 936.7500 ;
	    RECT 284.7000 935.1000 286.5000 935.2500 ;
	    RECT 291.9000 935.1000 293.7000 935.2500 ;
	    RECT 315.9000 936.7500 317.7000 936.9000 ;
	    RECT 347.1000 936.7500 348.9000 936.9000 ;
	    RECT 361.5000 936.7500 363.3000 936.9000 ;
	    RECT 378.3000 936.7500 380.1000 936.9000 ;
	    RECT 315.9000 935.2500 380.1000 936.7500 ;
	    RECT 315.9000 935.1000 317.7000 935.2500 ;
	    RECT 347.1000 935.1000 348.9000 935.2500 ;
	    RECT 361.5000 935.1000 363.3000 935.2500 ;
	    RECT 378.3000 935.1000 380.1000 935.2500 ;
	    RECT 560.7000 936.7500 562.5000 936.9000 ;
	    RECT 575.1000 936.7500 576.9000 936.9000 ;
	    RECT 560.7000 935.2500 576.9000 936.7500 ;
	    RECT 560.7000 935.1000 562.5000 935.2500 ;
	    RECT 575.1000 935.1000 576.9000 935.2500 ;
	    RECT 644.7000 936.7500 646.5000 936.9000 ;
	    RECT 788.7000 936.7500 790.5000 936.9000 ;
	    RECT 644.7000 935.2500 790.5000 936.7500 ;
	    RECT 644.7000 935.1000 646.5000 935.2500 ;
	    RECT 788.7000 935.1000 790.5000 935.2500 ;
	    RECT 913.5000 936.7500 915.3000 936.9000 ;
	    RECT 939.9000 936.7500 941.7000 936.9000 ;
	    RECT 913.5000 935.2500 941.7000 936.7500 ;
	    RECT 913.5000 935.1000 915.3000 935.2500 ;
	    RECT 939.9000 935.1000 941.7000 935.2500 ;
	    RECT 1115.1000 936.7500 1116.9000 936.9000 ;
	    RECT 1141.5000 936.7500 1143.3000 936.9000 ;
	    RECT 1115.1000 935.2500 1143.3000 936.7500 ;
	    RECT 1115.1000 935.1000 1116.9000 935.2500 ;
	    RECT 1141.5000 935.1000 1143.3000 935.2500 ;
	    RECT 1316.7001 936.7500 1318.5000 936.9000 ;
	    RECT 1321.5000 936.7500 1323.3000 936.9000 ;
	    RECT 1316.7001 935.2500 1323.3000 936.7500 ;
	    RECT 1316.7001 935.1000 1318.5000 935.2500 ;
	    RECT 1321.5000 935.1000 1323.3000 935.2500 ;
	    RECT 1429.5000 936.7500 1431.3000 936.9000 ;
	    RECT 1482.3000 936.7500 1484.1000 936.9000 ;
	    RECT 1429.5000 935.2500 1484.1000 936.7500 ;
	    RECT 1429.5000 935.1000 1431.3000 935.2500 ;
	    RECT 1482.3000 935.1000 1484.1000 935.2500 ;
	    RECT 80.7000 930.7500 82.5000 930.9000 ;
	    RECT 150.3000 930.7500 152.1000 930.9000 ;
	    RECT 80.7000 929.2500 152.1000 930.7500 ;
	    RECT 80.7000 929.1000 82.5000 929.2500 ;
	    RECT 150.3000 929.1000 152.1000 929.2500 ;
	    RECT 243.9000 930.7500 245.7000 930.9000 ;
	    RECT 265.5000 930.7500 267.3000 930.9000 ;
	    RECT 243.9000 929.2500 267.3000 930.7500 ;
	    RECT 243.9000 929.1000 245.7000 929.2500 ;
	    RECT 265.5000 929.1000 267.3000 929.2500 ;
	    RECT 294.3000 930.7500 296.1000 930.9000 ;
	    RECT 318.3000 930.7500 320.1000 930.9000 ;
	    RECT 294.3000 929.2500 320.1000 930.7500 ;
	    RECT 294.3000 929.1000 296.1000 929.2500 ;
	    RECT 318.3000 929.1000 320.1000 929.2500 ;
	    RECT 570.3000 930.7500 572.1000 930.9000 ;
	    RECT 587.1000 930.7500 588.9000 930.9000 ;
	    RECT 570.3000 929.2500 588.9000 930.7500 ;
	    RECT 570.3000 929.1000 572.1000 929.2500 ;
	    RECT 587.1000 929.1000 588.9000 929.2500 ;
	    RECT 615.9000 930.7500 617.7000 930.9000 ;
	    RECT 695.1000 930.7500 696.9000 930.9000 ;
	    RECT 615.9000 929.2500 696.9000 930.7500 ;
	    RECT 615.9000 929.1000 617.7000 929.2500 ;
	    RECT 695.1000 929.1000 696.9000 929.2500 ;
	    RECT 978.3000 930.7500 980.1000 930.9000 ;
	    RECT 1225.5000 930.7500 1227.3000 930.9000 ;
	    RECT 978.3000 929.2500 1227.3000 930.7500 ;
	    RECT 978.3000 929.1000 980.1000 929.2500 ;
	    RECT 1225.5000 929.1000 1227.3000 929.2500 ;
	    RECT 1295.1000 930.7500 1296.9000 930.9000 ;
	    RECT 1319.1000 930.7500 1320.9000 930.9000 ;
	    RECT 1295.1000 929.2500 1320.9000 930.7500 ;
	    RECT 1295.1000 929.1000 1296.9000 929.2500 ;
	    RECT 1319.1000 929.1000 1320.9000 929.2500 ;
	    RECT 1386.3000 930.7500 1388.1000 930.9000 ;
	    RECT 1455.9000 930.7500 1457.7001 930.9000 ;
	    RECT 1472.7001 930.7500 1474.5000 930.9000 ;
	    RECT 1386.3000 929.2500 1474.5000 930.7500 ;
	    RECT 1386.3000 929.1000 1388.1000 929.2500 ;
	    RECT 1455.9000 929.1000 1457.7001 929.2500 ;
	    RECT 1472.7001 929.1000 1474.5000 929.2500 ;
	    RECT 1477.5000 930.7500 1479.3000 930.9000 ;
	    RECT 1520.7001 930.7500 1522.5000 930.9000 ;
	    RECT 1477.5000 929.2500 1522.5000 930.7500 ;
	    RECT 1477.5000 929.1000 1479.3000 929.2500 ;
	    RECT 1520.7001 929.1000 1522.5000 929.2500 ;
	    RECT 66.3000 924.7500 68.1000 924.9000 ;
	    RECT 71.1000 924.7500 72.9000 924.9000 ;
	    RECT 66.3000 923.2500 72.9000 924.7500 ;
	    RECT 66.3000 923.1000 68.1000 923.2500 ;
	    RECT 71.1000 923.1000 72.9000 923.2500 ;
	    RECT 126.3000 924.7500 128.1000 924.9000 ;
	    RECT 243.9000 924.7500 245.7000 924.9000 ;
	    RECT 126.3000 923.2500 245.7000 924.7500 ;
	    RECT 126.3000 923.1000 128.1000 923.2500 ;
	    RECT 243.9000 923.1000 245.7000 923.2500 ;
	    RECT 253.5000 924.7500 255.3000 924.9000 ;
	    RECT 291.9000 924.7500 293.7000 924.9000 ;
	    RECT 253.5000 923.2500 293.7000 924.7500 ;
	    RECT 253.5000 923.1000 255.3000 923.2500 ;
	    RECT 291.9000 923.1000 293.7000 923.2500 ;
	    RECT 332.7000 924.7500 334.5000 924.9000 ;
	    RECT 363.9000 924.7500 365.7000 924.9000 ;
	    RECT 385.5000 924.7500 387.3000 924.9000 ;
	    RECT 332.7000 923.2500 387.3000 924.7500 ;
	    RECT 332.7000 923.1000 334.5000 923.2500 ;
	    RECT 363.9000 923.1000 365.7000 923.2500 ;
	    RECT 385.5000 923.1000 387.3000 923.2500 ;
	    RECT 491.1000 924.7500 492.9000 924.9000 ;
	    RECT 517.5000 924.7500 519.3000 924.9000 ;
	    RECT 534.3000 924.7500 536.1000 924.9000 ;
	    RECT 491.1000 923.2500 536.1000 924.7500 ;
	    RECT 491.1000 923.1000 492.9000 923.2500 ;
	    RECT 517.5000 923.1000 519.3000 923.2500 ;
	    RECT 534.3000 923.1000 536.1000 923.2500 ;
	    RECT 565.5000 924.7500 567.3000 924.9000 ;
	    RECT 714.3000 924.7500 716.1000 924.9000 ;
	    RECT 565.5000 923.2500 716.1000 924.7500 ;
	    RECT 565.5000 923.1000 567.3000 923.2500 ;
	    RECT 714.3000 923.1000 716.1000 923.2500 ;
	    RECT 774.3000 924.7500 776.1000 924.9000 ;
	    RECT 915.9000 924.7500 917.7000 924.9000 ;
	    RECT 959.1000 924.7500 960.9000 924.9000 ;
	    RECT 774.3000 923.2500 960.9000 924.7500 ;
	    RECT 774.3000 923.1000 776.1000 923.2500 ;
	    RECT 915.9000 923.1000 917.7000 923.2500 ;
	    RECT 959.1000 923.1000 960.9000 923.2500 ;
	    RECT 1083.9000 924.7500 1085.7001 924.9000 ;
	    RECT 1146.3000 924.7500 1148.1000 924.9000 ;
	    RECT 1083.9000 923.2500 1148.1000 924.7500 ;
	    RECT 1083.9000 923.1000 1085.7001 923.2500 ;
	    RECT 1146.3000 923.1000 1148.1000 923.2500 ;
	    RECT 1412.7001 924.7500 1414.5000 924.9000 ;
	    RECT 1429.5000 924.7500 1431.3000 924.9000 ;
	    RECT 1412.7001 923.2500 1431.3000 924.7500 ;
	    RECT 1412.7001 923.1000 1414.5000 923.2500 ;
	    RECT 1429.5000 923.1000 1431.3000 923.2500 ;
	    RECT 275.1000 918.7500 276.9000 918.9000 ;
	    RECT 294.3000 918.7500 296.1000 918.9000 ;
	    RECT 275.1000 917.2500 296.1000 918.7500 ;
	    RECT 275.1000 917.1000 276.9000 917.2500 ;
	    RECT 294.3000 917.1000 296.1000 917.2500 ;
	    RECT 299.1000 918.7500 300.9000 918.9000 ;
	    RECT 303.9000 918.7500 305.7000 918.9000 ;
	    RECT 332.7000 918.7500 334.5000 918.9000 ;
	    RECT 299.1000 917.2500 334.5000 918.7500 ;
	    RECT 299.1000 917.1000 300.9000 917.2500 ;
	    RECT 303.9000 917.1000 305.7000 917.2500 ;
	    RECT 332.7000 917.1000 334.5000 917.2500 ;
	    RECT 423.9000 918.7500 425.7000 918.9000 ;
	    RECT 428.7000 918.7500 430.5000 918.9000 ;
	    RECT 423.9000 917.2500 430.5000 918.7500 ;
	    RECT 423.9000 917.1000 425.7000 917.2500 ;
	    RECT 428.7000 917.1000 430.5000 917.2500 ;
	    RECT 517.5000 918.7500 519.3000 918.9000 ;
	    RECT 522.3000 918.7500 524.1000 918.9000 ;
	    RECT 517.5000 917.2500 524.1000 918.7500 ;
	    RECT 517.5000 917.1000 519.3000 917.2500 ;
	    RECT 522.3000 917.1000 524.1000 917.2500 ;
	    RECT 841.5000 918.7500 843.3000 918.9000 ;
	    RECT 870.3000 918.7500 872.1000 918.9000 ;
	    RECT 937.5000 918.7500 939.3000 918.9000 ;
	    RECT 841.5000 917.2500 939.3000 918.7500 ;
	    RECT 841.5000 917.1000 843.3000 917.2500 ;
	    RECT 870.3000 917.1000 872.1000 917.2500 ;
	    RECT 937.5000 917.1000 939.3000 917.2500 ;
	    RECT 947.1000 918.7500 948.9000 918.9000 ;
	    RECT 963.9000 918.7500 965.7000 918.9000 ;
	    RECT 947.1000 917.2500 965.7000 918.7500 ;
	    RECT 947.1000 917.1000 948.9000 917.2500 ;
	    RECT 963.9000 917.1000 965.7000 917.2500 ;
	    RECT 1367.1000 918.7500 1368.9000 918.9000 ;
	    RECT 1407.9000 918.7500 1409.7001 918.9000 ;
	    RECT 1367.1000 917.2500 1409.7001 918.7500 ;
	    RECT 1367.1000 917.1000 1368.9000 917.2500 ;
	    RECT 1407.9000 917.1000 1409.7001 917.2500 ;
	    RECT 1484.7001 918.7500 1486.5000 918.9000 ;
	    RECT 1491.9000 918.7500 1493.7001 918.9000 ;
	    RECT 1484.7001 917.2500 1493.7001 918.7500 ;
	    RECT 1484.7001 917.1000 1486.5000 917.2500 ;
	    RECT 1491.9000 917.1000 1493.7001 917.2500 ;
	    RECT 1530.3000 918.7500 1532.1000 918.9000 ;
	    RECT 1559.1000 918.7500 1560.9000 918.9000 ;
	    RECT 1563.9000 918.7500 1565.7001 918.9000 ;
	    RECT 1530.3000 917.2500 1565.7001 918.7500 ;
	    RECT 1530.3000 917.1000 1532.1000 917.2500 ;
	    RECT 1559.1000 917.1000 1560.9000 917.2500 ;
	    RECT 1563.9000 917.1000 1565.7001 917.2500 ;
	    RECT 47.1000 912.7500 48.9000 912.9000 ;
	    RECT 71.1000 912.7500 72.9000 912.9000 ;
	    RECT 47.1000 911.2500 72.9000 912.7500 ;
	    RECT 47.1000 911.1000 48.9000 911.2500 ;
	    RECT 71.1000 911.1000 72.9000 911.2500 ;
	    RECT 195.9000 912.7500 197.7000 912.9000 ;
	    RECT 212.7000 912.7500 214.5000 912.9000 ;
	    RECT 195.9000 911.2500 214.5000 912.7500 ;
	    RECT 195.9000 911.1000 197.7000 911.2500 ;
	    RECT 212.7000 911.1000 214.5000 911.2500 ;
	    RECT 654.3000 912.7500 656.1000 912.9000 ;
	    RECT 750.3000 912.7500 752.1000 912.9000 ;
	    RECT 654.3000 911.2500 752.1000 912.7500 ;
	    RECT 654.3000 911.1000 656.1000 911.2500 ;
	    RECT 750.3000 911.1000 752.1000 911.2500 ;
	    RECT 774.3000 912.7500 776.1000 912.9000 ;
	    RECT 795.9000 912.7500 797.7000 912.9000 ;
	    RECT 774.3000 911.2500 797.7000 912.7500 ;
	    RECT 774.3000 911.1000 776.1000 911.2500 ;
	    RECT 795.9000 911.1000 797.7000 911.2500 ;
	    RECT 877.5000 912.7500 879.3000 912.9000 ;
	    RECT 1167.9000 912.7500 1169.7001 912.9000 ;
	    RECT 877.5000 911.2500 1169.7001 912.7500 ;
	    RECT 877.5000 911.1000 879.3000 911.2500 ;
	    RECT 1167.9000 911.1000 1169.7001 911.2500 ;
	    RECT 1410.3000 912.7500 1412.1000 912.9000 ;
	    RECT 1427.1000 912.7500 1428.9000 912.9000 ;
	    RECT 1410.3000 911.2500 1428.9000 912.7500 ;
	    RECT 1410.3000 911.1000 1412.1000 911.2500 ;
	    RECT 1427.1000 911.1000 1428.9000 911.2500 ;
	    RECT 1477.5000 912.7500 1479.3000 912.9000 ;
	    RECT 1535.1000 912.7500 1536.9000 912.9000 ;
	    RECT 1477.5000 911.2500 1536.9000 912.7500 ;
	    RECT 1477.5000 911.1000 1479.3000 911.2500 ;
	    RECT 1535.1000 911.1000 1536.9000 911.2500 ;
	    RECT 1539.9000 912.7500 1541.7001 912.9000 ;
	    RECT 1544.7001 912.7500 1546.5000 912.9000 ;
	    RECT 1539.9000 911.2500 1546.5000 912.7500 ;
	    RECT 1539.9000 911.1000 1541.7001 911.2500 ;
	    RECT 1544.7001 911.1000 1546.5000 911.2500 ;
	    RECT 135.9000 906.7500 137.7000 906.9000 ;
	    RECT 224.7000 906.7500 226.5000 906.9000 ;
	    RECT 135.9000 905.2500 226.5000 906.7500 ;
	    RECT 135.9000 905.1000 137.7000 905.2500 ;
	    RECT 224.7000 905.1000 226.5000 905.2500 ;
	    RECT 239.1000 906.7500 240.9000 906.9000 ;
	    RECT 311.1000 906.7500 312.9000 906.9000 ;
	    RECT 239.1000 905.2500 312.9000 906.7500 ;
	    RECT 239.1000 905.1000 240.9000 905.2500 ;
	    RECT 311.1000 905.1000 312.9000 905.2500 ;
	    RECT 416.7000 906.7500 418.5000 906.9000 ;
	    RECT 572.7000 906.7500 574.5000 906.9000 ;
	    RECT 416.7000 905.2500 574.5000 906.7500 ;
	    RECT 416.7000 905.1000 418.5000 905.2500 ;
	    RECT 572.7000 905.1000 574.5000 905.2500 ;
	    RECT 956.7000 906.7500 958.5000 906.9000 ;
	    RECT 966.3000 906.7500 968.1000 906.9000 ;
	    RECT 956.7000 905.2500 968.1000 906.7500 ;
	    RECT 956.7000 905.1000 958.5000 905.2500 ;
	    RECT 966.3000 905.1000 968.1000 905.2500 ;
	    RECT 1141.5000 906.7500 1143.3000 906.9000 ;
	    RECT 1208.7001 906.7500 1210.5000 906.9000 ;
	    RECT 1218.3000 906.7500 1220.1000 906.9000 ;
	    RECT 1141.5000 905.2500 1220.1000 906.7500 ;
	    RECT 1141.5000 905.1000 1143.3000 905.2500 ;
	    RECT 1208.7001 905.1000 1210.5000 905.2500 ;
	    RECT 1218.3000 905.1000 1220.1000 905.2500 ;
	    RECT 1525.5000 906.7500 1527.3000 906.9000 ;
	    RECT 1547.1000 906.7500 1548.9000 906.9000 ;
	    RECT 1525.5000 905.2500 1548.9000 906.7500 ;
	    RECT 1525.5000 905.1000 1527.3000 905.2500 ;
	    RECT 1547.1000 905.1000 1548.9000 905.2500 ;
	    RECT 373.5000 900.7500 375.3000 900.9000 ;
	    RECT 409.5000 900.7500 411.3000 900.9000 ;
	    RECT 373.5000 899.2500 411.3000 900.7500 ;
	    RECT 373.5000 899.1000 375.3000 899.2500 ;
	    RECT 409.5000 899.1000 411.3000 899.2500 ;
	    RECT 471.9000 900.7500 473.7000 900.9000 ;
	    RECT 498.3000 900.7500 500.1000 900.9000 ;
	    RECT 572.7000 900.7500 574.5000 900.9000 ;
	    RECT 471.9000 899.2500 574.5000 900.7500 ;
	    RECT 471.9000 899.1000 473.7000 899.2500 ;
	    RECT 498.3000 899.1000 500.1000 899.2500 ;
	    RECT 572.7000 899.1000 574.5000 899.2500 ;
	    RECT 887.1000 900.7500 888.9000 900.9000 ;
	    RECT 894.3000 900.7500 896.1000 900.9000 ;
	    RECT 887.1000 899.2500 896.1000 900.7500 ;
	    RECT 887.1000 899.1000 888.9000 899.2500 ;
	    RECT 894.3000 899.1000 896.1000 899.2500 ;
	    RECT 966.3000 900.7500 968.1000 900.9000 ;
	    RECT 975.9000 900.7500 977.7000 900.9000 ;
	    RECT 966.3000 899.2500 977.7000 900.7500 ;
	    RECT 966.3000 899.1000 968.1000 899.2500 ;
	    RECT 975.9000 899.1000 977.7000 899.2500 ;
	    RECT 1155.9000 900.7500 1157.7001 900.9000 ;
	    RECT 1194.3000 900.7500 1196.1000 900.9000 ;
	    RECT 1155.9000 899.2500 1196.1000 900.7500 ;
	    RECT 1155.9000 899.1000 1157.7001 899.2500 ;
	    RECT 1194.3000 899.1000 1196.1000 899.2500 ;
	    RECT 150.3000 894.7500 152.1000 894.9000 ;
	    RECT 227.1000 894.7500 228.9000 894.9000 ;
	    RECT 299.1000 894.7500 300.9000 894.9000 ;
	    RECT 150.3000 893.2500 300.9000 894.7500 ;
	    RECT 150.3000 893.1000 152.1000 893.2500 ;
	    RECT 227.1000 893.1000 228.9000 893.2500 ;
	    RECT 299.1000 893.1000 300.9000 893.2500 ;
	    RECT 366.3000 894.7500 368.1000 894.9000 ;
	    RECT 371.1000 894.7500 372.9000 894.9000 ;
	    RECT 366.3000 893.2500 372.9000 894.7500 ;
	    RECT 366.3000 893.1000 368.1000 893.2500 ;
	    RECT 371.1000 893.1000 372.9000 893.2500 ;
	    RECT 555.9000 894.7500 557.7000 894.9000 ;
	    RECT 642.3000 894.7500 644.1000 894.9000 ;
	    RECT 555.9000 893.2500 644.1000 894.7500 ;
	    RECT 555.9000 893.1000 557.7000 893.2500 ;
	    RECT 642.3000 893.1000 644.1000 893.2500 ;
	    RECT 755.1000 894.7500 756.9000 894.9000 ;
	    RECT 764.7000 894.7500 766.5000 894.9000 ;
	    RECT 755.1000 893.2500 766.5000 894.7500 ;
	    RECT 755.1000 893.1000 756.9000 893.2500 ;
	    RECT 764.7000 893.1000 766.5000 893.2500 ;
	    RECT 937.5000 894.7500 939.3000 894.9000 ;
	    RECT 1009.5000 894.7500 1011.3000 894.9000 ;
	    RECT 937.5000 893.2500 1011.3000 894.7500 ;
	    RECT 937.5000 893.1000 939.3000 893.2500 ;
	    RECT 1009.5000 893.1000 1011.3000 893.2500 ;
	    RECT 1321.5000 894.7500 1323.3000 894.9000 ;
	    RECT 1479.9000 894.7500 1481.7001 894.9000 ;
	    RECT 1321.5000 893.2500 1481.7001 894.7500 ;
	    RECT 1321.5000 893.1000 1323.3000 893.2500 ;
	    RECT 1479.9000 893.1000 1481.7001 893.2500 ;
	    RECT 1501.5000 894.7500 1503.3000 894.9000 ;
	    RECT 1527.9000 894.7500 1529.7001 894.9000 ;
	    RECT 1501.5000 893.2500 1529.7001 894.7500 ;
	    RECT 1501.5000 893.1000 1503.3000 893.2500 ;
	    RECT 1527.9000 893.1000 1529.7001 893.2500 ;
	    RECT 303.9000 888.7500 305.7000 888.9000 ;
	    RECT 347.1000 888.7500 348.9000 888.9000 ;
	    RECT 303.9000 887.2500 348.9000 888.7500 ;
	    RECT 303.9000 887.1000 305.7000 887.2500 ;
	    RECT 347.1000 887.1000 348.9000 887.2500 ;
	    RECT 356.7000 888.7500 358.5000 888.9000 ;
	    RECT 385.5000 888.7500 387.3000 888.9000 ;
	    RECT 356.7000 887.2500 387.3000 888.7500 ;
	    RECT 356.7000 887.1000 358.5000 887.2500 ;
	    RECT 385.5000 887.1000 387.3000 887.2500 ;
	    RECT 719.1000 888.7500 720.9000 888.9000 ;
	    RECT 759.9000 888.7500 761.7000 888.9000 ;
	    RECT 719.1000 887.2500 761.7000 888.7500 ;
	    RECT 719.1000 887.1000 720.9000 887.2500 ;
	    RECT 759.9000 887.1000 761.7000 887.2500 ;
	    RECT 786.3000 888.7500 788.1000 888.9000 ;
	    RECT 829.5000 888.7500 831.3000 888.9000 ;
	    RECT 786.3000 887.2500 831.3000 888.7500 ;
	    RECT 786.3000 887.1000 788.1000 887.2500 ;
	    RECT 829.5000 887.1000 831.3000 887.2500 ;
	    RECT 889.5000 888.7500 891.3000 888.9000 ;
	    RECT 918.3000 888.7500 920.1000 888.9000 ;
	    RECT 889.5000 887.2500 920.1000 888.7500 ;
	    RECT 889.5000 887.1000 891.3000 887.2500 ;
	    RECT 918.3000 887.1000 920.1000 887.2500 ;
	    RECT 932.7000 888.7500 934.5000 888.9000 ;
	    RECT 1028.7001 888.7500 1030.5000 888.9000 ;
	    RECT 932.7000 887.2500 1030.5000 888.7500 ;
	    RECT 932.7000 887.1000 934.5000 887.2500 ;
	    RECT 1028.7001 887.1000 1030.5000 887.2500 ;
	    RECT 1223.1000 888.7500 1224.9000 888.9000 ;
	    RECT 1237.5000 888.7500 1239.3000 888.9000 ;
	    RECT 1223.1000 887.2500 1239.3000 888.7500 ;
	    RECT 1223.1000 887.1000 1224.9000 887.2500 ;
	    RECT 1237.5000 887.1000 1239.3000 887.2500 ;
	    RECT 1441.5000 888.7500 1443.3000 888.9000 ;
	    RECT 1465.5000 888.7500 1467.3000 888.9000 ;
	    RECT 1441.5000 887.2500 1467.3000 888.7500 ;
	    RECT 1441.5000 887.1000 1443.3000 887.2500 ;
	    RECT 1465.5000 887.1000 1467.3000 887.2500 ;
	    RECT 51.9000 882.7500 53.7000 882.9000 ;
	    RECT 121.5000 882.7500 123.3000 882.9000 ;
	    RECT 140.7000 882.7500 142.5000 882.9000 ;
	    RECT 51.9000 881.2500 142.5000 882.7500 ;
	    RECT 51.9000 881.1000 53.7000 881.2500 ;
	    RECT 121.5000 881.1000 123.3000 881.2500 ;
	    RECT 140.7000 881.1000 142.5000 881.2500 ;
	    RECT 167.1000 882.7500 168.9000 882.9000 ;
	    RECT 222.3000 882.7500 224.1000 882.9000 ;
	    RECT 167.1000 881.2500 224.1000 882.7500 ;
	    RECT 167.1000 881.1000 168.9000 881.2500 ;
	    RECT 222.3000 881.1000 224.1000 881.2500 ;
	    RECT 680.7000 882.7500 682.5000 882.9000 ;
	    RECT 757.5000 882.7500 759.3000 882.9000 ;
	    RECT 680.7000 881.2500 759.3000 882.7500 ;
	    RECT 680.7000 881.1000 682.5000 881.2500 ;
	    RECT 757.5000 881.1000 759.3000 881.2500 ;
	    RECT 884.7000 882.7500 886.5000 882.9000 ;
	    RECT 891.9000 882.7500 893.7000 882.9000 ;
	    RECT 884.7000 881.2500 893.7000 882.7500 ;
	    RECT 884.7000 881.1000 886.5000 881.2500 ;
	    RECT 891.9000 881.1000 893.7000 881.2500 ;
	    RECT 944.7000 882.7500 946.5000 882.9000 ;
	    RECT 959.1000 882.7500 960.9000 882.9000 ;
	    RECT 944.7000 881.2500 960.9000 882.7500 ;
	    RECT 944.7000 881.1000 946.5000 881.2500 ;
	    RECT 959.1000 881.1000 960.9000 881.2500 ;
	    RECT 1009.5000 882.7500 1011.3000 882.9000 ;
	    RECT 1033.5000 882.7500 1035.3000 882.9000 ;
	    RECT 1009.5000 881.2500 1035.3000 882.7500 ;
	    RECT 1009.5000 881.1000 1011.3000 881.2500 ;
	    RECT 1033.5000 881.1000 1035.3000 881.2500 ;
	    RECT 1203.9000 882.7500 1205.7001 882.9000 ;
	    RECT 1223.1000 882.7500 1224.9000 882.9000 ;
	    RECT 1203.9000 881.2500 1224.9000 882.7500 ;
	    RECT 1203.9000 881.1000 1205.7001 881.2500 ;
	    RECT 1223.1000 881.1000 1224.9000 881.2500 ;
	    RECT 169.5000 876.7500 171.3000 876.9000 ;
	    RECT 217.5000 876.7500 219.3000 876.9000 ;
	    RECT 169.5000 875.2500 219.3000 876.7500 ;
	    RECT 169.5000 875.1000 171.3000 875.2500 ;
	    RECT 217.5000 875.1000 219.3000 875.2500 ;
	    RECT 625.5000 876.7500 627.3000 876.9000 ;
	    RECT 654.3000 876.7500 656.1000 876.9000 ;
	    RECT 625.5000 875.2500 656.1000 876.7500 ;
	    RECT 625.5000 875.1000 627.3000 875.2500 ;
	    RECT 654.3000 875.1000 656.1000 875.2500 ;
	    RECT 726.3000 876.7500 728.1000 876.9000 ;
	    RECT 745.5000 876.7500 747.3000 876.9000 ;
	    RECT 726.3000 875.2500 747.3000 876.7500 ;
	    RECT 726.3000 875.1000 728.1000 875.2500 ;
	    RECT 745.5000 875.1000 747.3000 875.2500 ;
	    RECT 896.7000 876.7500 898.5000 876.9000 ;
	    RECT 1004.7000 876.7500 1006.5000 876.9000 ;
	    RECT 896.7000 875.2500 1006.5000 876.7500 ;
	    RECT 896.7000 875.1000 898.5000 875.2500 ;
	    RECT 1004.7000 875.1000 1006.5000 875.2500 ;
	    RECT 1026.3000 876.7500 1028.1000 876.9000 ;
	    RECT 1038.3000 876.7500 1040.1000 876.9000 ;
	    RECT 1026.3000 875.2500 1040.1000 876.7500 ;
	    RECT 1026.3000 875.1000 1028.1000 875.2500 ;
	    RECT 1038.3000 875.1000 1040.1000 875.2500 ;
	    RECT 1208.7001 876.7500 1210.5000 876.9000 ;
	    RECT 1316.7001 876.7500 1318.5000 876.9000 ;
	    RECT 1208.7001 875.2500 1318.5000 876.7500 ;
	    RECT 1208.7001 875.1000 1210.5000 875.2500 ;
	    RECT 1316.7001 875.1000 1318.5000 875.2500 ;
	    RECT 123.9000 870.7500 125.7000 870.9000 ;
	    RECT 174.3000 870.7500 176.1000 870.9000 ;
	    RECT 123.9000 869.2500 176.1000 870.7500 ;
	    RECT 123.9000 869.1000 125.7000 869.2500 ;
	    RECT 174.3000 869.1000 176.1000 869.2500 ;
	    RECT 299.1000 870.7500 300.9000 870.9000 ;
	    RECT 332.7000 870.7500 334.5000 870.9000 ;
	    RECT 299.1000 869.2500 334.5000 870.7500 ;
	    RECT 299.1000 869.1000 300.9000 869.2500 ;
	    RECT 332.7000 869.1000 334.5000 869.2500 ;
	    RECT 351.9000 870.7500 353.7000 870.9000 ;
	    RECT 373.5000 870.7500 375.3000 870.9000 ;
	    RECT 351.9000 869.2500 375.3000 870.7500 ;
	    RECT 351.9000 869.1000 353.7000 869.2500 ;
	    RECT 373.5000 869.1000 375.3000 869.2500 ;
	    RECT 591.9000 870.7500 593.7000 870.9000 ;
	    RECT 606.3000 870.7500 608.1000 870.9000 ;
	    RECT 735.9000 870.7500 737.7000 870.9000 ;
	    RECT 591.9000 869.2500 737.7000 870.7500 ;
	    RECT 591.9000 869.1000 593.7000 869.2500 ;
	    RECT 606.3000 869.1000 608.1000 869.2500 ;
	    RECT 735.9000 869.1000 737.7000 869.2500 ;
	    RECT 927.9000 870.7500 929.7000 870.9000 ;
	    RECT 932.7000 870.7500 934.5000 870.9000 ;
	    RECT 927.9000 869.2500 934.5000 870.7500 ;
	    RECT 927.9000 869.1000 929.7000 869.2500 ;
	    RECT 932.7000 869.1000 934.5000 869.2500 ;
	    RECT 1225.5000 870.7500 1227.3000 870.9000 ;
	    RECT 1340.7001 870.7500 1342.5000 870.9000 ;
	    RECT 1225.5000 869.2500 1342.5000 870.7500 ;
	    RECT 1225.5000 869.1000 1227.3000 869.2500 ;
	    RECT 1340.7001 869.1000 1342.5000 869.2500 ;
	    RECT 1379.1000 870.7500 1380.9000 870.9000 ;
	    RECT 1475.1000 870.7500 1476.9000 870.9000 ;
	    RECT 1518.3000 870.7500 1520.1000 870.9000 ;
	    RECT 1379.1000 869.2500 1520.1000 870.7500 ;
	    RECT 1379.1000 869.1000 1380.9000 869.2500 ;
	    RECT 1475.1000 869.1000 1476.9000 869.2500 ;
	    RECT 1518.3000 869.1000 1520.1000 869.2500 ;
	    RECT 1530.3000 870.7500 1532.1000 870.9000 ;
	    RECT 1544.7001 870.7500 1546.5000 870.9000 ;
	    RECT 1530.3000 869.2500 1546.5000 870.7500 ;
	    RECT 1530.3000 869.1000 1532.1000 869.2500 ;
	    RECT 1544.7001 869.1000 1546.5000 869.2500 ;
	    RECT 25.5000 864.7500 27.3000 864.9000 ;
	    RECT 54.3000 864.7500 56.1000 864.9000 ;
	    RECT 25.5000 863.2500 56.1000 864.7500 ;
	    RECT 25.5000 863.1000 27.3000 863.2500 ;
	    RECT 54.3000 863.1000 56.1000 863.2500 ;
	    RECT 102.3000 864.7500 104.1000 864.9000 ;
	    RECT 126.3000 864.7500 128.1000 864.9000 ;
	    RECT 102.3000 863.2500 128.1000 864.7500 ;
	    RECT 102.3000 863.1000 104.1000 863.2500 ;
	    RECT 126.3000 863.1000 128.1000 863.2500 ;
	    RECT 210.3000 864.7500 212.1000 864.9000 ;
	    RECT 215.1000 864.7500 216.9000 864.9000 ;
	    RECT 251.1000 864.7500 252.9000 864.9000 ;
	    RECT 301.5000 864.7500 303.3000 864.9000 ;
	    RECT 210.3000 863.2500 303.3000 864.7500 ;
	    RECT 210.3000 863.1000 212.1000 863.2500 ;
	    RECT 215.1000 863.1000 216.9000 863.2500 ;
	    RECT 251.1000 863.1000 252.9000 863.2500 ;
	    RECT 301.5000 863.1000 303.3000 863.2500 ;
	    RECT 332.7000 864.7500 334.5000 864.9000 ;
	    RECT 387.9000 864.7500 389.7000 864.9000 ;
	    RECT 332.7000 863.2500 389.7000 864.7500 ;
	    RECT 332.7000 863.1000 334.5000 863.2500 ;
	    RECT 387.9000 863.1000 389.7000 863.2500 ;
	    RECT 548.7000 864.7500 550.5000 864.9000 ;
	    RECT 572.7000 864.7500 574.5000 864.9000 ;
	    RECT 548.7000 863.2500 574.5000 864.7500 ;
	    RECT 548.7000 863.1000 550.5000 863.2500 ;
	    RECT 572.7000 863.1000 574.5000 863.2500 ;
	    RECT 577.5000 864.7500 579.3000 864.9000 ;
	    RECT 591.9000 864.7500 593.7000 864.9000 ;
	    RECT 577.5000 863.2500 593.7000 864.7500 ;
	    RECT 577.5000 863.1000 579.3000 863.2500 ;
	    RECT 591.9000 863.1000 593.7000 863.2500 ;
	    RECT 683.1000 864.7500 684.9000 864.9000 ;
	    RECT 815.1000 864.7500 816.9000 864.9000 ;
	    RECT 683.1000 863.2500 816.9000 864.7500 ;
	    RECT 683.1000 863.1000 684.9000 863.2500 ;
	    RECT 815.1000 863.1000 816.9000 863.2500 ;
	    RECT 1052.7001 864.7500 1054.5000 864.9000 ;
	    RECT 1223.1000 864.7500 1224.9000 864.9000 ;
	    RECT 1052.7001 863.2500 1224.9000 864.7500 ;
	    RECT 1052.7001 863.1000 1054.5000 863.2500 ;
	    RECT 1223.1000 863.1000 1224.9000 863.2500 ;
	    RECT 1364.7001 864.7500 1366.5000 864.9000 ;
	    RECT 1376.7001 864.7500 1378.5000 864.9000 ;
	    RECT 1364.7001 863.2500 1378.5000 864.7500 ;
	    RECT 1364.7001 863.1000 1366.5000 863.2500 ;
	    RECT 1376.7001 863.1000 1378.5000 863.2500 ;
	    RECT 18.3000 858.7500 20.1000 858.9000 ;
	    RECT 23.1000 858.7500 24.9000 858.9000 ;
	    RECT 18.3000 857.2500 24.9000 858.7500 ;
	    RECT 18.3000 857.1000 20.1000 857.2500 ;
	    RECT 23.1000 857.1000 24.9000 857.2500 ;
	    RECT 116.7000 858.7500 118.5000 858.9000 ;
	    RECT 126.3000 858.7500 128.1000 858.9000 ;
	    RECT 116.7000 857.2500 128.1000 858.7500 ;
	    RECT 116.7000 857.1000 118.5000 857.2500 ;
	    RECT 126.3000 857.1000 128.1000 857.2500 ;
	    RECT 152.7000 858.7500 154.5000 858.9000 ;
	    RECT 159.9000 858.7500 161.7000 858.9000 ;
	    RECT 152.7000 857.2500 161.7000 858.7500 ;
	    RECT 152.7000 857.1000 154.5000 857.2500 ;
	    RECT 159.9000 857.1000 161.7000 857.2500 ;
	    RECT 219.9000 858.7500 221.7000 858.9000 ;
	    RECT 306.3000 858.7500 308.1000 858.9000 ;
	    RECT 219.9000 857.2500 308.1000 858.7500 ;
	    RECT 219.9000 857.1000 221.7000 857.2500 ;
	    RECT 306.3000 857.1000 308.1000 857.2500 ;
	    RECT 601.5000 858.7500 603.3000 858.9000 ;
	    RECT 656.7000 858.7500 658.5000 858.9000 ;
	    RECT 733.5000 858.7500 735.3000 858.9000 ;
	    RECT 601.5000 857.2500 735.3000 858.7500 ;
	    RECT 601.5000 857.1000 603.3000 857.2500 ;
	    RECT 656.7000 857.1000 658.5000 857.2500 ;
	    RECT 733.5000 857.1000 735.3000 857.2500 ;
	    RECT 942.3000 858.7500 944.1000 858.9000 ;
	    RECT 983.1000 858.7500 984.9000 858.9000 ;
	    RECT 942.3000 857.2500 984.9000 858.7500 ;
	    RECT 942.3000 857.1000 944.1000 857.2500 ;
	    RECT 983.1000 857.1000 984.9000 857.2500 ;
	    RECT 1119.9000 858.7500 1121.7001 858.9000 ;
	    RECT 1177.5000 858.7500 1179.3000 858.9000 ;
	    RECT 1119.9000 857.2500 1179.3000 858.7500 ;
	    RECT 1119.9000 857.1000 1121.7001 857.2500 ;
	    RECT 1177.5000 857.1000 1179.3000 857.2500 ;
	    RECT 1223.1000 858.7500 1224.9000 858.9000 ;
	    RECT 1242.3000 858.7500 1244.1000 858.9000 ;
	    RECT 1223.1000 857.2500 1244.1000 858.7500 ;
	    RECT 1223.1000 857.1000 1224.9000 857.2500 ;
	    RECT 1242.3000 857.1000 1244.1000 857.2500 ;
	    RECT 1371.9000 858.7500 1373.7001 858.9000 ;
	    RECT 1417.5000 858.7500 1419.3000 858.9000 ;
	    RECT 1424.7001 858.7500 1426.5000 858.9000 ;
	    RECT 1371.9000 857.2500 1426.5000 858.7500 ;
	    RECT 1371.9000 857.1000 1373.7001 857.2500 ;
	    RECT 1417.5000 857.1000 1419.3000 857.2500 ;
	    RECT 1424.7001 857.1000 1426.5000 857.2500 ;
	    RECT 1544.7001 858.7500 1546.5000 858.9000 ;
	    RECT 1551.9000 858.7500 1553.7001 858.9000 ;
	    RECT 1544.7001 857.2500 1553.7001 858.7500 ;
	    RECT 1544.7001 857.1000 1546.5000 857.2500 ;
	    RECT 1551.9000 857.1000 1553.7001 857.2500 ;
	    RECT 18.3000 852.7500 20.1000 852.9000 ;
	    RECT 51.9000 852.7500 53.7000 852.9000 ;
	    RECT 18.3000 851.2500 53.7000 852.7500 ;
	    RECT 18.3000 851.1000 20.1000 851.2500 ;
	    RECT 51.9000 851.1000 53.7000 851.2500 ;
	    RECT 181.5000 852.7500 183.3000 852.9000 ;
	    RECT 215.1000 852.7500 216.9000 852.9000 ;
	    RECT 287.1000 852.7500 288.9000 852.9000 ;
	    RECT 181.5000 851.2500 288.9000 852.7500 ;
	    RECT 181.5000 851.1000 183.3000 851.2500 ;
	    RECT 215.1000 851.1000 216.9000 851.2500 ;
	    RECT 287.1000 851.1000 288.9000 851.2500 ;
	    RECT 342.3000 852.7500 344.1000 852.9000 ;
	    RECT 383.1000 852.7500 384.9000 852.9000 ;
	    RECT 342.3000 851.2500 384.9000 852.7500 ;
	    RECT 342.3000 851.1000 344.1000 851.2500 ;
	    RECT 383.1000 851.1000 384.9000 851.2500 ;
	    RECT 474.3000 852.7500 476.1000 852.9000 ;
	    RECT 483.9000 852.7500 485.7000 852.9000 ;
	    RECT 474.3000 851.2500 485.7000 852.7500 ;
	    RECT 474.3000 851.1000 476.1000 851.2500 ;
	    RECT 483.9000 851.1000 485.7000 851.2500 ;
	    RECT 613.5000 852.7500 615.3000 852.9000 ;
	    RECT 647.1000 852.7500 648.9000 852.9000 ;
	    RECT 678.3000 852.7500 680.1000 852.9000 ;
	    RECT 699.9000 852.7500 701.7000 852.9000 ;
	    RECT 613.5000 851.2500 701.7000 852.7500 ;
	    RECT 613.5000 851.1000 615.3000 851.2500 ;
	    RECT 647.1000 851.1000 648.9000 851.2500 ;
	    RECT 678.3000 851.1000 680.1000 851.2500 ;
	    RECT 699.9000 851.1000 701.7000 851.2500 ;
	    RECT 743.1000 852.7500 744.9000 852.9000 ;
	    RECT 843.9000 852.7500 845.7000 852.9000 ;
	    RECT 743.1000 851.2500 845.7000 852.7500 ;
	    RECT 743.1000 851.1000 744.9000 851.2500 ;
	    RECT 843.9000 851.1000 845.7000 851.2500 ;
	    RECT 980.7000 852.7500 982.5000 852.9000 ;
	    RECT 1167.9000 852.7500 1169.7001 852.9000 ;
	    RECT 980.7000 851.2500 1169.7001 852.7500 ;
	    RECT 980.7000 851.1000 982.5000 851.2500 ;
	    RECT 1167.9000 851.1000 1169.7001 851.2500 ;
	    RECT 164.7000 846.7500 166.5000 846.9000 ;
	    RECT 183.9000 846.7500 185.7000 846.9000 ;
	    RECT 373.5000 846.7500 375.3000 846.9000 ;
	    RECT 164.7000 845.2500 375.3000 846.7500 ;
	    RECT 164.7000 845.1000 166.5000 845.2500 ;
	    RECT 183.9000 845.1000 185.7000 845.2500 ;
	    RECT 373.5000 845.1000 375.3000 845.2500 ;
	    RECT 383.1000 846.7500 384.9000 846.9000 ;
	    RECT 411.9000 846.7500 413.7000 846.9000 ;
	    RECT 383.1000 845.2500 413.7000 846.7500 ;
	    RECT 383.1000 845.1000 384.9000 845.2500 ;
	    RECT 411.9000 845.1000 413.7000 845.2500 ;
	    RECT 517.5000 846.7500 519.3000 846.9000 ;
	    RECT 577.5000 846.7500 579.3000 846.9000 ;
	    RECT 517.5000 845.2500 579.3000 846.7500 ;
	    RECT 517.5000 845.1000 519.3000 845.2500 ;
	    RECT 577.5000 845.1000 579.3000 845.2500 ;
	    RECT 671.1000 846.7500 672.9000 846.9000 ;
	    RECT 692.7000 846.7500 694.5000 846.9000 ;
	    RECT 671.1000 845.2500 694.5000 846.7500 ;
	    RECT 671.1000 845.1000 672.9000 845.2500 ;
	    RECT 692.7000 845.1000 694.5000 845.2500 ;
	    RECT 740.7000 846.7500 742.5000 846.9000 ;
	    RECT 798.3000 846.7500 800.1000 846.9000 ;
	    RECT 740.7000 845.2500 800.1000 846.7500 ;
	    RECT 740.7000 845.1000 742.5000 845.2500 ;
	    RECT 798.3000 845.1000 800.1000 845.2500 ;
	    RECT 920.7000 846.7500 922.5000 846.9000 ;
	    RECT 1031.1000 846.7500 1032.9000 846.9000 ;
	    RECT 920.7000 845.2500 1032.9000 846.7500 ;
	    RECT 920.7000 845.1000 922.5000 845.2500 ;
	    RECT 1031.1000 845.1000 1032.9000 845.2500 ;
	    RECT 1182.3000 846.7500 1184.1000 846.9000 ;
	    RECT 1206.3000 846.7500 1208.1000 846.9000 ;
	    RECT 1213.5000 846.7500 1215.3000 846.9000 ;
	    RECT 1182.3000 845.2500 1215.3000 846.7500 ;
	    RECT 1182.3000 845.1000 1184.1000 845.2500 ;
	    RECT 1206.3000 845.1000 1208.1000 845.2500 ;
	    RECT 1213.5000 845.1000 1215.3000 845.2500 ;
	    RECT 1551.9000 846.7500 1553.7001 846.9000 ;
	    RECT 1566.3000 846.7500 1568.1000 846.9000 ;
	    RECT 1551.9000 845.2500 1568.1000 846.7500 ;
	    RECT 1551.9000 845.1000 1553.7001 845.2500 ;
	    RECT 1566.3000 845.1000 1568.1000 845.2500 ;
	    RECT 246.3000 840.7500 248.1000 840.9000 ;
	    RECT 356.7000 840.7500 358.5000 840.9000 ;
	    RECT 246.3000 839.2500 358.5000 840.7500 ;
	    RECT 246.3000 839.1000 248.1000 839.2500 ;
	    RECT 356.7000 839.1000 358.5000 839.2500 ;
	    RECT 495.9000 840.7500 497.7000 840.9000 ;
	    RECT 575.1000 840.7500 576.9000 840.9000 ;
	    RECT 495.9000 839.2500 576.9000 840.7500 ;
	    RECT 495.9000 839.1000 497.7000 839.2500 ;
	    RECT 575.1000 839.1000 576.9000 839.2500 ;
	    RECT 704.7000 840.7500 706.5000 840.9000 ;
	    RECT 755.1000 840.7500 756.9000 840.9000 ;
	    RECT 704.7000 839.2500 756.9000 840.7500 ;
	    RECT 704.7000 839.1000 706.5000 839.2500 ;
	    RECT 755.1000 839.1000 756.9000 839.2500 ;
	    RECT 887.1000 840.7500 888.9000 840.9000 ;
	    RECT 978.3000 840.7500 980.1000 840.9000 ;
	    RECT 887.1000 839.2500 980.1000 840.7500 ;
	    RECT 887.1000 839.1000 888.9000 839.2500 ;
	    RECT 978.3000 839.1000 980.1000 839.2500 ;
	    RECT 1177.5000 840.7500 1179.3000 840.9000 ;
	    RECT 1194.3000 840.7500 1196.1000 840.9000 ;
	    RECT 1177.5000 839.2500 1196.1000 840.7500 ;
	    RECT 1177.5000 839.1000 1179.3000 839.2500 ;
	    RECT 1194.3000 839.1000 1196.1000 839.2500 ;
	    RECT 1247.1000 840.7500 1248.9000 840.9000 ;
	    RECT 1431.9000 840.7500 1433.7001 840.9000 ;
	    RECT 1247.1000 839.2500 1433.7001 840.7500 ;
	    RECT 1247.1000 839.1000 1248.9000 839.2500 ;
	    RECT 1431.9000 839.1000 1433.7001 839.2500 ;
	    RECT 1518.3000 840.7500 1520.1000 840.9000 ;
	    RECT 1556.7001 840.7500 1558.5000 840.9000 ;
	    RECT 1518.3000 839.2500 1558.5000 840.7500 ;
	    RECT 1518.3000 839.1000 1520.1000 839.2500 ;
	    RECT 1556.7001 839.1000 1558.5000 839.2500 ;
	    RECT 188.7000 834.7500 190.5000 834.9000 ;
	    RECT 243.9000 834.7500 245.7000 834.9000 ;
	    RECT 188.7000 833.2500 245.7000 834.7500 ;
	    RECT 188.7000 833.1000 190.5000 833.2500 ;
	    RECT 243.9000 833.1000 245.7000 833.2500 ;
	    RECT 272.7000 834.7500 274.5000 834.9000 ;
	    RECT 366.3000 834.7500 368.1000 834.9000 ;
	    RECT 272.7000 833.2500 368.1000 834.7500 ;
	    RECT 272.7000 833.1000 274.5000 833.2500 ;
	    RECT 366.3000 833.1000 368.1000 833.2500 ;
	    RECT 553.5000 834.7500 555.3000 834.9000 ;
	    RECT 582.3000 834.7500 584.1000 834.9000 ;
	    RECT 553.5000 833.2500 584.1000 834.7500 ;
	    RECT 553.5000 833.1000 555.3000 833.2500 ;
	    RECT 582.3000 833.1000 584.1000 833.2500 ;
	    RECT 642.3000 834.7500 644.1000 834.9000 ;
	    RECT 738.3000 834.7500 740.1000 834.9000 ;
	    RECT 642.3000 833.2500 740.1000 834.7500 ;
	    RECT 642.3000 833.1000 644.1000 833.2500 ;
	    RECT 738.3000 833.1000 740.1000 833.2500 ;
	    RECT 1023.9000 834.7500 1025.7001 834.9000 ;
	    RECT 1201.5000 834.7500 1203.3000 834.9000 ;
	    RECT 1023.9000 833.2500 1203.3000 834.7500 ;
	    RECT 1023.9000 833.1000 1025.7001 833.2500 ;
	    RECT 1201.5000 833.1000 1203.3000 833.2500 ;
	    RECT 1266.3000 834.7500 1268.1000 834.9000 ;
	    RECT 1530.3000 834.7500 1532.1000 834.9000 ;
	    RECT 1266.3000 833.2500 1532.1000 834.7500 ;
	    RECT 1266.3000 833.1000 1268.1000 833.2500 ;
	    RECT 1530.3000 833.1000 1532.1000 833.2500 ;
	    RECT 155.1000 828.7500 156.9000 828.9000 ;
	    RECT 174.3000 828.7500 176.1000 828.9000 ;
	    RECT 155.1000 827.2500 176.1000 828.7500 ;
	    RECT 155.1000 827.1000 156.9000 827.2500 ;
	    RECT 174.3000 827.1000 176.1000 827.2500 ;
	    RECT 222.3000 828.7500 224.1000 828.9000 ;
	    RECT 253.5000 828.7500 255.3000 828.9000 ;
	    RECT 222.3000 827.2500 255.3000 828.7500 ;
	    RECT 222.3000 827.1000 224.1000 827.2500 ;
	    RECT 253.5000 827.1000 255.3000 827.2500 ;
	    RECT 399.9000 828.7500 401.7000 828.9000 ;
	    RECT 407.1000 828.7500 408.9000 828.9000 ;
	    RECT 399.9000 827.2500 408.9000 828.7500 ;
	    RECT 399.9000 827.1000 401.7000 827.2500 ;
	    RECT 407.1000 827.1000 408.9000 827.2500 ;
	    RECT 541.5000 828.7500 543.3000 828.9000 ;
	    RECT 577.5000 828.7500 579.3000 828.9000 ;
	    RECT 541.5000 827.2500 579.3000 828.7500 ;
	    RECT 541.5000 827.1000 543.3000 827.2500 ;
	    RECT 577.5000 827.1000 579.3000 827.2500 ;
	    RECT 731.1000 828.7500 732.9000 828.9000 ;
	    RECT 738.3000 828.7500 740.1000 828.9000 ;
	    RECT 731.1000 827.2500 740.1000 828.7500 ;
	    RECT 731.1000 827.1000 732.9000 827.2500 ;
	    RECT 738.3000 827.1000 740.1000 827.2500 ;
	    RECT 903.9000 828.7500 905.7000 828.9000 ;
	    RECT 923.1000 828.7500 924.9000 828.9000 ;
	    RECT 903.9000 827.2500 924.9000 828.7500 ;
	    RECT 903.9000 827.1000 905.7000 827.2500 ;
	    RECT 923.1000 827.1000 924.9000 827.2500 ;
	    RECT 966.3000 828.7500 968.1000 828.9000 ;
	    RECT 1050.3000 828.7500 1052.1000 828.9000 ;
	    RECT 966.3000 827.2500 1052.1000 828.7500 ;
	    RECT 966.3000 827.1000 968.1000 827.2500 ;
	    RECT 1050.3000 827.1000 1052.1000 827.2500 ;
	    RECT 1151.1000 828.7500 1152.9000 828.9000 ;
	    RECT 1167.9000 828.7500 1169.7001 828.9000 ;
	    RECT 1151.1000 827.2500 1169.7001 828.7500 ;
	    RECT 1151.1000 827.1000 1152.9000 827.2500 ;
	    RECT 1167.9000 827.1000 1169.7001 827.2500 ;
	    RECT 1424.7001 828.7500 1426.5000 828.9000 ;
	    RECT 1503.9000 828.7500 1505.7001 828.9000 ;
	    RECT 1424.7001 827.2500 1505.7001 828.7500 ;
	    RECT 1424.7001 827.1000 1426.5000 827.2500 ;
	    RECT 1503.9000 827.1000 1505.7001 827.2500 ;
	    RECT 1532.7001 828.7500 1534.5000 828.9000 ;
	    RECT 1563.9000 828.7500 1565.7001 828.9000 ;
	    RECT 1532.7001 827.2500 1565.7001 828.7500 ;
	    RECT 1532.7001 827.1000 1534.5000 827.2500 ;
	    RECT 1563.9000 827.1000 1565.7001 827.2500 ;
	    RECT 119.1000 822.7500 120.9000 822.9000 ;
	    RECT 155.1000 822.7500 156.9000 822.9000 ;
	    RECT 119.1000 821.2500 156.9000 822.7500 ;
	    RECT 119.1000 821.1000 120.9000 821.2500 ;
	    RECT 155.1000 821.1000 156.9000 821.2500 ;
	    RECT 188.7000 822.7500 190.5000 822.9000 ;
	    RECT 291.9000 822.7500 293.7000 822.9000 ;
	    RECT 188.7000 821.2500 293.7000 822.7500 ;
	    RECT 188.7000 821.1000 190.5000 821.2500 ;
	    RECT 291.9000 821.1000 293.7000 821.2500 ;
	    RECT 339.9000 822.7500 341.7000 822.9000 ;
	    RECT 407.1000 822.7500 408.9000 822.9000 ;
	    RECT 339.9000 821.2500 408.9000 822.7500 ;
	    RECT 339.9000 821.1000 341.7000 821.2500 ;
	    RECT 407.1000 821.1000 408.9000 821.2500 ;
	    RECT 551.1000 822.7500 552.9000 822.9000 ;
	    RECT 563.1000 822.7500 564.9000 822.9000 ;
	    RECT 551.1000 821.2500 564.9000 822.7500 ;
	    RECT 551.1000 821.1000 552.9000 821.2500 ;
	    RECT 563.1000 821.1000 564.9000 821.2500 ;
	    RECT 577.5000 822.7500 579.3000 822.9000 ;
	    RECT 783.9000 822.7500 785.7000 822.9000 ;
	    RECT 577.5000 821.2500 785.7000 822.7500 ;
	    RECT 577.5000 821.1000 579.3000 821.2500 ;
	    RECT 783.9000 821.1000 785.7000 821.2500 ;
	    RECT 800.7000 822.7500 802.5000 822.9000 ;
	    RECT 807.9000 822.7500 809.7000 822.9000 ;
	    RECT 819.9000 822.7500 821.7000 822.9000 ;
	    RECT 800.7000 821.2500 821.7000 822.7500 ;
	    RECT 800.7000 821.1000 802.5000 821.2500 ;
	    RECT 807.9000 821.1000 809.7000 821.2500 ;
	    RECT 819.9000 821.1000 821.7000 821.2500 ;
	    RECT 827.1000 822.7500 828.9000 822.9000 ;
	    RECT 841.5000 822.7500 843.3000 822.9000 ;
	    RECT 827.1000 821.2500 843.3000 822.7500 ;
	    RECT 827.1000 821.1000 828.9000 821.2500 ;
	    RECT 841.5000 821.1000 843.3000 821.2500 ;
	    RECT 846.3000 822.7500 848.1000 822.9000 ;
	    RECT 865.5000 822.7500 867.3000 822.9000 ;
	    RECT 846.3000 821.2500 867.3000 822.7500 ;
	    RECT 846.3000 821.1000 848.1000 821.2500 ;
	    RECT 865.5000 821.1000 867.3000 821.2500 ;
	    RECT 887.1000 822.7500 888.9000 822.9000 ;
	    RECT 918.3000 822.7500 920.1000 822.9000 ;
	    RECT 887.1000 821.2500 920.1000 822.7500 ;
	    RECT 887.1000 821.1000 888.9000 821.2500 ;
	    RECT 918.3000 821.1000 920.1000 821.2500 ;
	    RECT 973.5000 822.7500 975.3000 822.9000 ;
	    RECT 985.5000 822.7500 987.3000 822.9000 ;
	    RECT 973.5000 821.2500 987.3000 822.7500 ;
	    RECT 973.5000 821.1000 975.3000 821.2500 ;
	    RECT 985.5000 821.1000 987.3000 821.2500 ;
	    RECT 1393.5000 822.7500 1395.3000 822.9000 ;
	    RECT 1539.9000 822.7500 1541.7001 822.9000 ;
	    RECT 1393.5000 821.2500 1541.7001 822.7500 ;
	    RECT 1393.5000 821.1000 1395.3000 821.2500 ;
	    RECT 1539.9000 821.1000 1541.7001 821.2500 ;
	    RECT 138.3000 816.7500 140.1000 816.9000 ;
	    RECT 164.7000 816.7500 166.5000 816.9000 ;
	    RECT 138.3000 815.2500 166.5000 816.7500 ;
	    RECT 138.3000 815.1000 140.1000 815.2500 ;
	    RECT 164.7000 815.1000 166.5000 815.2500 ;
	    RECT 572.7000 816.7500 574.5000 816.9000 ;
	    RECT 594.3000 816.7500 596.1000 816.9000 ;
	    RECT 572.7000 815.2500 596.1000 816.7500 ;
	    RECT 572.7000 815.1000 574.5000 815.2500 ;
	    RECT 594.3000 815.1000 596.1000 815.2500 ;
	    RECT 630.3000 816.7500 632.1000 816.9000 ;
	    RECT 685.5000 816.7500 687.3000 816.9000 ;
	    RECT 630.3000 815.2500 687.3000 816.7500 ;
	    RECT 630.3000 815.1000 632.1000 815.2500 ;
	    RECT 685.5000 815.1000 687.3000 815.2500 ;
	    RECT 733.5000 816.7500 735.3000 816.9000 ;
	    RECT 740.7000 816.7500 742.5000 816.9000 ;
	    RECT 733.5000 815.2500 742.5000 816.7500 ;
	    RECT 733.5000 815.1000 735.3000 815.2500 ;
	    RECT 740.7000 815.1000 742.5000 815.2500 ;
	    RECT 750.3000 816.7500 752.1000 816.9000 ;
	    RECT 788.7000 816.7500 790.5000 816.9000 ;
	    RECT 750.3000 815.2500 790.5000 816.7500 ;
	    RECT 750.3000 815.1000 752.1000 815.2500 ;
	    RECT 788.7000 815.1000 790.5000 815.2500 ;
	    RECT 817.5000 816.7500 819.3000 816.9000 ;
	    RECT 829.5000 816.7500 831.3000 816.9000 ;
	    RECT 817.5000 815.2500 831.3000 816.7500 ;
	    RECT 817.5000 815.1000 819.3000 815.2500 ;
	    RECT 829.5000 815.1000 831.3000 815.2500 ;
	    RECT 942.3000 816.7500 944.1000 816.9000 ;
	    RECT 963.9000 816.7500 965.7000 816.9000 ;
	    RECT 942.3000 815.2500 965.7000 816.7500 ;
	    RECT 942.3000 815.1000 944.1000 815.2500 ;
	    RECT 963.9000 815.1000 965.7000 815.2500 ;
	    RECT 1117.5000 816.7500 1119.3000 816.9000 ;
	    RECT 1235.1000 816.7500 1236.9000 816.9000 ;
	    RECT 1117.5000 815.2500 1236.9000 816.7500 ;
	    RECT 1117.5000 815.1000 1119.3000 815.2500 ;
	    RECT 1235.1000 815.1000 1236.9000 815.2500 ;
	    RECT 318.3000 810.7500 320.1000 810.9000 ;
	    RECT 349.5000 810.7500 351.3000 810.9000 ;
	    RECT 368.7000 810.7500 370.5000 810.9000 ;
	    RECT 318.3000 809.2500 370.5000 810.7500 ;
	    RECT 318.3000 809.1000 320.1000 809.2500 ;
	    RECT 349.5000 809.1000 351.3000 809.2500 ;
	    RECT 368.7000 809.1000 370.5000 809.2500 ;
	    RECT 407.1000 810.7500 408.9000 810.9000 ;
	    RECT 431.1000 810.7500 432.9000 810.9000 ;
	    RECT 407.1000 809.2500 432.9000 810.7500 ;
	    RECT 407.1000 809.1000 408.9000 809.2500 ;
	    RECT 431.1000 809.1000 432.9000 809.2500 ;
	    RECT 632.7000 810.7500 634.5000 810.9000 ;
	    RECT 637.5000 810.7500 639.3000 810.9000 ;
	    RECT 632.7000 809.2500 639.3000 810.7500 ;
	    RECT 632.7000 809.1000 634.5000 809.2500 ;
	    RECT 637.5000 809.1000 639.3000 809.2500 ;
	    RECT 709.5000 810.7500 711.3000 810.9000 ;
	    RECT 716.7000 810.7500 718.5000 810.9000 ;
	    RECT 709.5000 809.2500 718.5000 810.7500 ;
	    RECT 709.5000 809.1000 711.3000 809.2500 ;
	    RECT 716.7000 809.1000 718.5000 809.2500 ;
	    RECT 731.1000 810.7500 732.9000 810.9000 ;
	    RECT 759.9000 810.7500 761.7000 810.9000 ;
	    RECT 731.1000 809.2500 761.7000 810.7500 ;
	    RECT 731.1000 809.1000 732.9000 809.2500 ;
	    RECT 759.9000 809.1000 761.7000 809.2500 ;
	    RECT 947.1000 810.7500 948.9000 810.9000 ;
	    RECT 1050.3000 810.7500 1052.1000 810.9000 ;
	    RECT 947.1000 809.2500 1052.1000 810.7500 ;
	    RECT 947.1000 809.1000 948.9000 809.2500 ;
	    RECT 1050.3000 809.1000 1052.1000 809.2500 ;
	    RECT 1059.9000 810.7500 1061.7001 810.9000 ;
	    RECT 1177.5000 810.7500 1179.3000 810.9000 ;
	    RECT 1059.9000 809.2500 1179.3000 810.7500 ;
	    RECT 1059.9000 809.1000 1061.7001 809.2500 ;
	    RECT 1177.5000 809.1000 1179.3000 809.2500 ;
	    RECT 1388.7001 810.7500 1390.5000 810.9000 ;
	    RECT 1467.9000 810.7500 1469.7001 810.9000 ;
	    RECT 1388.7001 809.2500 1469.7001 810.7500 ;
	    RECT 1388.7001 809.1000 1390.5000 809.2500 ;
	    RECT 1467.9000 809.1000 1469.7001 809.2500 ;
	    RECT 1527.9000 810.7500 1529.7001 810.9000 ;
	    RECT 1547.1000 810.7500 1548.9000 810.9000 ;
	    RECT 1527.9000 809.2500 1548.9000 810.7500 ;
	    RECT 1527.9000 809.1000 1529.7001 809.2500 ;
	    RECT 1547.1000 809.1000 1548.9000 809.2500 ;
	    RECT 128.7000 804.7500 130.5000 804.9000 ;
	    RECT 186.3000 804.7500 188.1000 804.9000 ;
	    RECT 128.7000 803.2500 188.1000 804.7500 ;
	    RECT 128.7000 803.1000 130.5000 803.2500 ;
	    RECT 186.3000 803.1000 188.1000 803.2500 ;
	    RECT 210.3000 804.7500 212.1000 804.9000 ;
	    RECT 224.7000 804.7500 226.5000 804.9000 ;
	    RECT 210.3000 803.2500 226.5000 804.7500 ;
	    RECT 210.3000 803.1000 212.1000 803.2500 ;
	    RECT 224.7000 803.1000 226.5000 803.2500 ;
	    RECT 423.9000 804.7500 425.7000 804.9000 ;
	    RECT 519.9000 804.7500 521.7000 804.9000 ;
	    RECT 423.9000 803.2500 521.7000 804.7500 ;
	    RECT 423.9000 803.1000 425.7000 803.2500 ;
	    RECT 519.9000 803.1000 521.7000 803.2500 ;
	    RECT 570.3000 804.7500 572.1000 804.9000 ;
	    RECT 582.3000 804.7500 584.1000 804.9000 ;
	    RECT 570.3000 803.2500 584.1000 804.7500 ;
	    RECT 570.3000 803.1000 572.1000 803.2500 ;
	    RECT 582.3000 803.1000 584.1000 803.2500 ;
	    RECT 606.3000 804.7500 608.1000 804.9000 ;
	    RECT 680.7000 804.7500 682.5000 804.9000 ;
	    RECT 606.3000 803.2500 682.5000 804.7500 ;
	    RECT 606.3000 803.1000 608.1000 803.2500 ;
	    RECT 680.7000 803.1000 682.5000 803.2500 ;
	    RECT 690.3000 804.7500 692.1000 804.9000 ;
	    RECT 728.7000 804.7500 730.5000 804.9000 ;
	    RECT 690.3000 803.2500 730.5000 804.7500 ;
	    RECT 690.3000 803.1000 692.1000 803.2500 ;
	    RECT 728.7000 803.1000 730.5000 803.2500 ;
	    RECT 786.3000 804.7500 788.1000 804.9000 ;
	    RECT 791.1000 804.7500 792.9000 804.9000 ;
	    RECT 786.3000 803.2500 792.9000 804.7500 ;
	    RECT 786.3000 803.1000 788.1000 803.2500 ;
	    RECT 791.1000 803.1000 792.9000 803.2500 ;
	    RECT 819.9000 804.7500 821.7000 804.9000 ;
	    RECT 851.1000 804.7500 852.9000 804.9000 ;
	    RECT 819.9000 803.2500 852.9000 804.7500 ;
	    RECT 819.9000 803.1000 821.7000 803.2500 ;
	    RECT 851.1000 803.1000 852.9000 803.2500 ;
	    RECT 858.3000 804.7500 860.1000 804.9000 ;
	    RECT 879.9000 804.7500 881.7000 804.9000 ;
	    RECT 887.1000 804.7500 888.9000 804.9000 ;
	    RECT 858.3000 803.2500 888.9000 804.7500 ;
	    RECT 858.3000 803.1000 860.1000 803.2500 ;
	    RECT 879.9000 803.1000 881.7000 803.2500 ;
	    RECT 887.1000 803.1000 888.9000 803.2500 ;
	    RECT 1098.3000 804.7500 1100.1000 804.9000 ;
	    RECT 1177.5000 804.7500 1179.3000 804.9000 ;
	    RECT 1098.3000 803.2500 1179.3000 804.7500 ;
	    RECT 1098.3000 803.1000 1100.1000 803.2500 ;
	    RECT 1177.5000 803.1000 1179.3000 803.2500 ;
	    RECT 1211.1000 804.7500 1212.9000 804.9000 ;
	    RECT 1319.1000 804.7500 1320.9000 804.9000 ;
	    RECT 1211.1000 803.2500 1320.9000 804.7500 ;
	    RECT 1211.1000 803.1000 1212.9000 803.2500 ;
	    RECT 1319.1000 803.1000 1320.9000 803.2500 ;
	    RECT 1455.9000 804.7500 1457.7001 804.9000 ;
	    RECT 1491.9000 804.7500 1493.7001 804.9000 ;
	    RECT 1455.9000 803.2500 1493.7001 804.7500 ;
	    RECT 1455.9000 803.1000 1457.7001 803.2500 ;
	    RECT 1491.9000 803.1000 1493.7001 803.2500 ;
	    RECT 47.1000 798.7500 48.9000 798.9000 ;
	    RECT 155.1000 798.7500 156.9000 798.9000 ;
	    RECT 47.1000 797.2500 156.9000 798.7500 ;
	    RECT 47.1000 797.1000 48.9000 797.2500 ;
	    RECT 155.1000 797.1000 156.9000 797.2500 ;
	    RECT 164.7000 798.7500 166.5000 798.9000 ;
	    RECT 241.5000 798.7500 243.3000 798.9000 ;
	    RECT 164.7000 797.2500 243.3000 798.7500 ;
	    RECT 164.7000 797.1000 166.5000 797.2500 ;
	    RECT 241.5000 797.1000 243.3000 797.2500 ;
	    RECT 354.3000 798.7500 356.1000 798.9000 ;
	    RECT 387.9000 798.7500 389.7000 798.9000 ;
	    RECT 354.3000 797.2500 389.7000 798.7500 ;
	    RECT 354.3000 797.1000 356.1000 797.2500 ;
	    RECT 387.9000 797.1000 389.7000 797.2500 ;
	    RECT 627.9000 798.7500 629.7000 798.9000 ;
	    RECT 671.1000 798.7500 672.9000 798.9000 ;
	    RECT 627.9000 797.2500 672.9000 798.7500 ;
	    RECT 627.9000 797.1000 629.7000 797.2500 ;
	    RECT 671.1000 797.1000 672.9000 797.2500 ;
	    RECT 735.9000 798.7500 737.7000 798.9000 ;
	    RECT 750.3000 798.7500 752.1000 798.9000 ;
	    RECT 735.9000 797.2500 752.1000 798.7500 ;
	    RECT 735.9000 797.1000 737.7000 797.2500 ;
	    RECT 750.3000 797.1000 752.1000 797.2500 ;
	    RECT 795.9000 798.7500 797.7000 798.9000 ;
	    RECT 841.5000 798.7500 843.3000 798.9000 ;
	    RECT 795.9000 797.2500 843.3000 798.7500 ;
	    RECT 795.9000 797.1000 797.7000 797.2500 ;
	    RECT 841.5000 797.1000 843.3000 797.2500 ;
	    RECT 1139.1000 798.7500 1140.9000 798.9000 ;
	    RECT 1170.3000 798.7500 1172.1000 798.9000 ;
	    RECT 1139.1000 797.2500 1172.1000 798.7500 ;
	    RECT 1139.1000 797.1000 1140.9000 797.2500 ;
	    RECT 1170.3000 797.1000 1172.1000 797.2500 ;
	    RECT 1206.3000 798.7500 1208.1000 798.9000 ;
	    RECT 1309.5000 798.7500 1311.3000 798.9000 ;
	    RECT 1206.3000 797.2500 1311.3000 798.7500 ;
	    RECT 1206.3000 797.1000 1208.1000 797.2500 ;
	    RECT 1309.5000 797.1000 1311.3000 797.2500 ;
	    RECT 1340.7001 798.7500 1342.5000 798.9000 ;
	    RECT 1405.5000 798.7500 1407.3000 798.9000 ;
	    RECT 1340.7001 797.2500 1407.3000 798.7500 ;
	    RECT 1340.7001 797.1000 1342.5000 797.2500 ;
	    RECT 1405.5000 797.1000 1407.3000 797.2500 ;
	    RECT 1458.3000 798.7500 1460.1000 798.9000 ;
	    RECT 1494.3000 798.7500 1496.1000 798.9000 ;
	    RECT 1458.3000 797.2500 1496.1000 798.7500 ;
	    RECT 1458.3000 797.1000 1460.1000 797.2500 ;
	    RECT 1494.3000 797.1000 1496.1000 797.2500 ;
	    RECT 1523.1000 798.7500 1524.9000 798.9000 ;
	    RECT 1563.9000 798.7500 1565.7001 798.9000 ;
	    RECT 1523.1000 797.2500 1565.7001 798.7500 ;
	    RECT 1523.1000 797.1000 1524.9000 797.2500 ;
	    RECT 1563.9000 797.1000 1565.7001 797.2500 ;
	    RECT 383.1000 792.7500 384.9000 792.9000 ;
	    RECT 392.7000 792.7500 394.5000 792.9000 ;
	    RECT 383.1000 791.2500 394.5000 792.7500 ;
	    RECT 383.1000 791.1000 384.9000 791.2500 ;
	    RECT 392.7000 791.1000 394.5000 791.2500 ;
	    RECT 522.3000 792.7500 524.1000 792.9000 ;
	    RECT 611.1000 792.7500 612.9000 792.9000 ;
	    RECT 522.3000 791.2500 612.9000 792.7500 ;
	    RECT 522.3000 791.1000 524.1000 791.2500 ;
	    RECT 611.1000 791.1000 612.9000 791.2500 ;
	    RECT 635.1000 792.7500 636.9000 792.9000 ;
	    RECT 678.3000 792.7500 680.1000 792.9000 ;
	    RECT 635.1000 791.2500 680.1000 792.7500 ;
	    RECT 635.1000 791.1000 636.9000 791.2500 ;
	    RECT 678.3000 791.1000 680.1000 791.2500 ;
	    RECT 757.5000 792.7500 759.3000 792.9000 ;
	    RECT 807.9000 792.7500 809.7000 792.9000 ;
	    RECT 757.5000 791.2500 809.7000 792.7500 ;
	    RECT 757.5000 791.1000 759.3000 791.2500 ;
	    RECT 807.9000 791.1000 809.7000 791.2500 ;
	    RECT 959.1000 792.7500 960.9000 792.9000 ;
	    RECT 1139.1000 792.7500 1140.9000 792.9000 ;
	    RECT 959.1000 791.2500 1140.9000 792.7500 ;
	    RECT 959.1000 791.1000 960.9000 791.2500 ;
	    RECT 1139.1000 791.1000 1140.9000 791.2500 ;
	    RECT 1405.5000 792.7500 1407.3000 792.9000 ;
	    RECT 1535.1000 792.7500 1536.9000 792.9000 ;
	    RECT 1405.5000 791.2500 1536.9000 792.7500 ;
	    RECT 1405.5000 791.1000 1407.3000 791.2500 ;
	    RECT 1535.1000 791.1000 1536.9000 791.2500 ;
	    RECT 1547.1000 792.7500 1548.9000 792.9000 ;
	    RECT 1561.5000 792.7500 1563.3000 792.9000 ;
	    RECT 1547.1000 791.2500 1563.3000 792.7500 ;
	    RECT 1547.1000 791.1000 1548.9000 791.2500 ;
	    RECT 1561.5000 791.1000 1563.3000 791.2500 ;
	    RECT 90.3000 786.7500 92.1000 786.9000 ;
	    RECT 203.1000 786.7500 204.9000 786.9000 ;
	    RECT 90.3000 785.2500 204.9000 786.7500 ;
	    RECT 90.3000 785.1000 92.1000 785.2500 ;
	    RECT 203.1000 785.1000 204.9000 785.2500 ;
	    RECT 385.5000 786.7500 387.3000 786.9000 ;
	    RECT 411.9000 786.7500 413.7000 786.9000 ;
	    RECT 385.5000 785.2500 413.7000 786.7500 ;
	    RECT 385.5000 785.1000 387.3000 785.2500 ;
	    RECT 411.9000 785.1000 413.7000 785.2500 ;
	    RECT 582.3000 786.7500 584.1000 786.9000 ;
	    RECT 599.1000 786.7500 600.9000 786.9000 ;
	    RECT 582.3000 785.2500 600.9000 786.7500 ;
	    RECT 582.3000 785.1000 584.1000 785.2500 ;
	    RECT 599.1000 785.1000 600.9000 785.2500 ;
	    RECT 740.7000 786.7500 742.5000 786.9000 ;
	    RECT 764.7000 786.7500 766.5000 786.9000 ;
	    RECT 740.7000 785.2500 766.5000 786.7500 ;
	    RECT 740.7000 785.1000 742.5000 785.2500 ;
	    RECT 764.7000 785.1000 766.5000 785.2500 ;
	    RECT 1064.7001 786.7500 1066.5000 786.9000 ;
	    RECT 1086.3000 786.7500 1088.1000 786.9000 ;
	    RECT 1093.5000 786.7500 1095.3000 786.9000 ;
	    RECT 1064.7001 785.2500 1095.3000 786.7500 ;
	    RECT 1064.7001 785.1000 1066.5000 785.2500 ;
	    RECT 1086.3000 785.1000 1088.1000 785.2500 ;
	    RECT 1093.5000 785.1000 1095.3000 785.2500 ;
	    RECT 1244.7001 786.7500 1246.5000 786.9000 ;
	    RECT 1323.9000 786.7500 1325.7001 786.9000 ;
	    RECT 1244.7001 785.2500 1325.7001 786.7500 ;
	    RECT 1244.7001 785.1000 1246.5000 785.2500 ;
	    RECT 1323.9000 785.1000 1325.7001 785.2500 ;
	    RECT 1407.9000 786.7500 1409.7001 786.9000 ;
	    RECT 1458.3000 786.7500 1460.1000 786.9000 ;
	    RECT 1407.9000 785.2500 1460.1000 786.7500 ;
	    RECT 1407.9000 785.1000 1409.7001 785.2500 ;
	    RECT 1458.3000 785.1000 1460.1000 785.2500 ;
	    RECT 1503.9000 786.7500 1505.7001 786.9000 ;
	    RECT 1559.1000 786.7500 1560.9000 786.9000 ;
	    RECT 1503.9000 785.2500 1560.9000 786.7500 ;
	    RECT 1503.9000 785.1000 1505.7001 785.2500 ;
	    RECT 1559.1000 785.1000 1560.9000 785.2500 ;
	    RECT 236.7000 780.7500 238.5000 780.9000 ;
	    RECT 251.1000 780.7500 252.9000 780.9000 ;
	    RECT 236.7000 779.2500 252.9000 780.7500 ;
	    RECT 236.7000 779.1000 238.5000 779.2500 ;
	    RECT 251.1000 779.1000 252.9000 779.2500 ;
	    RECT 366.3000 780.7500 368.1000 780.9000 ;
	    RECT 620.7000 780.7500 622.5000 780.9000 ;
	    RECT 366.3000 779.2500 622.5000 780.7500 ;
	    RECT 366.3000 779.1000 368.1000 779.2500 ;
	    RECT 620.7000 779.1000 622.5000 779.2500 ;
	    RECT 723.9000 780.7500 725.7000 780.9000 ;
	    RECT 786.3000 780.7500 788.1000 780.9000 ;
	    RECT 723.9000 779.2500 788.1000 780.7500 ;
	    RECT 723.9000 779.1000 725.7000 779.2500 ;
	    RECT 786.3000 779.1000 788.1000 779.2500 ;
	    RECT 815.1000 780.7500 816.9000 780.9000 ;
	    RECT 995.1000 780.7500 996.9000 780.9000 ;
	    RECT 815.1000 779.2500 996.9000 780.7500 ;
	    RECT 815.1000 779.1000 816.9000 779.2500 ;
	    RECT 995.1000 779.1000 996.9000 779.2500 ;
	    RECT 1038.3000 780.7500 1040.1000 780.9000 ;
	    RECT 1045.5000 780.7500 1047.3000 780.9000 ;
	    RECT 1038.3000 779.2500 1047.3000 780.7500 ;
	    RECT 1038.3000 779.1000 1040.1000 779.2500 ;
	    RECT 1045.5000 779.1000 1047.3000 779.2500 ;
	    RECT 1093.5000 780.7500 1095.3000 780.9000 ;
	    RECT 1098.3000 780.7500 1100.1000 780.9000 ;
	    RECT 1093.5000 779.2500 1100.1000 780.7500 ;
	    RECT 1093.5000 779.1000 1095.3000 779.2500 ;
	    RECT 1098.3000 779.1000 1100.1000 779.2500 ;
	    RECT 1151.1000 780.7500 1152.9000 780.9000 ;
	    RECT 1158.3000 780.7500 1160.1000 780.9000 ;
	    RECT 1151.1000 779.2500 1160.1000 780.7500 ;
	    RECT 1151.1000 779.1000 1152.9000 779.2500 ;
	    RECT 1158.3000 779.1000 1160.1000 779.2500 ;
	    RECT 1527.9000 780.7500 1529.7001 780.9000 ;
	    RECT 1532.7001 780.7500 1534.5000 780.9000 ;
	    RECT 1527.9000 779.2500 1534.5000 780.7500 ;
	    RECT 1527.9000 779.1000 1529.7001 779.2500 ;
	    RECT 1532.7001 779.1000 1534.5000 779.2500 ;
	    RECT 114.3000 774.7500 116.1000 774.9000 ;
	    RECT 191.1000 774.7500 192.9000 774.9000 ;
	    RECT 114.3000 773.2500 192.9000 774.7500 ;
	    RECT 114.3000 773.1000 116.1000 773.2500 ;
	    RECT 191.1000 773.1000 192.9000 773.2500 ;
	    RECT 361.5000 774.7500 363.3000 774.9000 ;
	    RECT 411.9000 774.7500 413.7000 774.9000 ;
	    RECT 361.5000 773.2500 413.7000 774.7500 ;
	    RECT 361.5000 773.1000 363.3000 773.2500 ;
	    RECT 411.9000 773.1000 413.7000 773.2500 ;
	    RECT 515.1000 774.7500 516.9000 774.9000 ;
	    RECT 587.1000 774.7500 588.9000 774.9000 ;
	    RECT 515.1000 773.2500 588.9000 774.7500 ;
	    RECT 515.1000 773.1000 516.9000 773.2500 ;
	    RECT 587.1000 773.1000 588.9000 773.2500 ;
	    RECT 899.1000 774.7500 900.9000 774.9000 ;
	    RECT 942.3000 774.7500 944.1000 774.9000 ;
	    RECT 899.1000 773.2500 944.1000 774.7500 ;
	    RECT 899.1000 773.1000 900.9000 773.2500 ;
	    RECT 942.3000 773.1000 944.1000 773.2500 ;
	    RECT 966.3000 774.7500 968.1000 774.9000 ;
	    RECT 999.9000 774.7500 1001.7000 774.9000 ;
	    RECT 1059.9000 774.7500 1061.7001 774.9000 ;
	    RECT 966.3000 773.2500 1061.7001 774.7500 ;
	    RECT 966.3000 773.1000 968.1000 773.2500 ;
	    RECT 999.9000 773.1000 1001.7000 773.2500 ;
	    RECT 1059.9000 773.1000 1061.7001 773.2500 ;
	    RECT 1064.7001 774.7500 1066.5000 774.9000 ;
	    RECT 1103.1000 774.7500 1104.9000 774.9000 ;
	    RECT 1064.7001 773.2500 1104.9000 774.7500 ;
	    RECT 1064.7001 773.1000 1066.5000 773.2500 ;
	    RECT 1103.1000 773.1000 1104.9000 773.2500 ;
	    RECT 1314.3000 774.7500 1316.1000 774.9000 ;
	    RECT 1412.7001 774.7500 1414.5000 774.9000 ;
	    RECT 1314.3000 773.2500 1414.5000 774.7500 ;
	    RECT 1314.3000 773.1000 1316.1000 773.2500 ;
	    RECT 1412.7001 773.1000 1414.5000 773.2500 ;
	    RECT 1427.1000 774.7500 1428.9000 774.9000 ;
	    RECT 1453.5000 774.7500 1455.3000 774.9000 ;
	    RECT 1427.1000 773.2500 1455.3000 774.7500 ;
	    RECT 1427.1000 773.1000 1428.9000 773.2500 ;
	    RECT 1453.5000 773.1000 1455.3000 773.2500 ;
	    RECT 155.1000 768.7500 156.9000 768.9000 ;
	    RECT 167.1000 768.7500 168.9000 768.9000 ;
	    RECT 155.1000 767.2500 168.9000 768.7500 ;
	    RECT 155.1000 767.1000 156.9000 767.2500 ;
	    RECT 167.1000 767.1000 168.9000 767.2500 ;
	    RECT 587.1000 768.7500 588.9000 768.9000 ;
	    RECT 644.7000 768.7500 646.5000 768.9000 ;
	    RECT 587.1000 767.2500 646.5000 768.7500 ;
	    RECT 587.1000 767.1000 588.9000 767.2500 ;
	    RECT 644.7000 767.1000 646.5000 767.2500 ;
	    RECT 661.5000 768.7500 663.3000 768.9000 ;
	    RECT 702.3000 768.7500 704.1000 768.9000 ;
	    RECT 661.5000 767.2500 704.1000 768.7500 ;
	    RECT 661.5000 767.1000 663.3000 767.2500 ;
	    RECT 702.3000 767.1000 704.1000 767.2500 ;
	    RECT 719.1000 768.7500 720.9000 768.9000 ;
	    RECT 735.9000 768.7500 737.7000 768.9000 ;
	    RECT 719.1000 767.2500 737.7000 768.7500 ;
	    RECT 719.1000 767.1000 720.9000 767.2500 ;
	    RECT 735.9000 767.1000 737.7000 767.2500 ;
	    RECT 783.9000 768.7500 785.7000 768.9000 ;
	    RECT 824.7000 768.7500 826.5000 768.9000 ;
	    RECT 855.9000 768.7500 857.7000 768.9000 ;
	    RECT 870.3000 768.7500 872.1000 768.9000 ;
	    RECT 901.5000 768.7500 903.3000 768.9000 ;
	    RECT 783.9000 767.2500 903.3000 768.7500 ;
	    RECT 783.9000 767.1000 785.7000 767.2500 ;
	    RECT 824.7000 767.1000 826.5000 767.2500 ;
	    RECT 855.9000 767.1000 857.7000 767.2500 ;
	    RECT 870.3000 767.1000 872.1000 767.2500 ;
	    RECT 901.5000 767.1000 903.3000 767.2500 ;
	    RECT 995.1000 768.7500 996.9000 768.9000 ;
	    RECT 1093.5000 768.7500 1095.3000 768.9000 ;
	    RECT 995.1000 767.2500 1095.3000 768.7500 ;
	    RECT 995.1000 767.1000 996.9000 767.2500 ;
	    RECT 1093.5000 767.1000 1095.3000 767.2500 ;
	    RECT 1100.7001 768.7500 1102.5000 768.9000 ;
	    RECT 1134.3000 768.7500 1136.1000 768.9000 ;
	    RECT 1100.7001 767.2500 1136.1000 768.7500 ;
	    RECT 1100.7001 767.1000 1102.5000 767.2500 ;
	    RECT 1134.3000 767.1000 1136.1000 767.2500 ;
	    RECT 1501.5000 768.7500 1503.3000 768.9000 ;
	    RECT 1544.7001 768.7500 1546.5000 768.9000 ;
	    RECT 1501.5000 767.2500 1546.5000 768.7500 ;
	    RECT 1501.5000 767.1000 1503.3000 767.2500 ;
	    RECT 1544.7001 767.1000 1546.5000 767.2500 ;
	    RECT 104.7000 762.7500 106.5000 762.9000 ;
	    RECT 284.7000 762.7500 286.5000 762.9000 ;
	    RECT 104.7000 761.2500 286.5000 762.7500 ;
	    RECT 104.7000 761.1000 106.5000 761.2500 ;
	    RECT 284.7000 761.1000 286.5000 761.2500 ;
	    RECT 548.7000 762.7500 550.5000 762.9000 ;
	    RECT 596.7000 762.7500 598.5000 762.9000 ;
	    RECT 548.7000 761.2500 598.5000 762.7500 ;
	    RECT 548.7000 761.1000 550.5000 761.2500 ;
	    RECT 596.7000 761.1000 598.5000 761.2500 ;
	    RECT 656.7000 762.7500 658.5000 762.9000 ;
	    RECT 663.9000 762.7500 665.7000 762.9000 ;
	    RECT 656.7000 761.2500 665.7000 762.7500 ;
	    RECT 656.7000 761.1000 658.5000 761.2500 ;
	    RECT 663.9000 761.1000 665.7000 761.2500 ;
	    RECT 687.9000 762.7500 689.7000 762.9000 ;
	    RECT 759.9000 762.7500 761.7000 762.9000 ;
	    RECT 687.9000 761.2500 761.7000 762.7500 ;
	    RECT 687.9000 761.1000 689.7000 761.2500 ;
	    RECT 759.9000 761.1000 761.7000 761.2500 ;
	    RECT 800.7000 762.7500 802.5000 762.9000 ;
	    RECT 860.7000 762.7500 862.5000 762.9000 ;
	    RECT 906.3000 762.7500 908.1000 762.9000 ;
	    RECT 800.7000 761.2500 908.1000 762.7500 ;
	    RECT 800.7000 761.1000 802.5000 761.2500 ;
	    RECT 860.7000 761.1000 862.5000 761.2500 ;
	    RECT 906.3000 761.1000 908.1000 761.2500 ;
	    RECT 911.1000 762.7500 912.9000 762.9000 ;
	    RECT 949.5000 762.7500 951.3000 762.9000 ;
	    RECT 911.1000 761.2500 951.3000 762.7500 ;
	    RECT 911.1000 761.1000 912.9000 761.2500 ;
	    RECT 949.5000 761.1000 951.3000 761.2500 ;
	    RECT 1143.9000 762.7500 1145.7001 762.9000 ;
	    RECT 1309.5000 762.7500 1311.3000 762.9000 ;
	    RECT 1393.5000 762.7500 1395.3000 762.9000 ;
	    RECT 1412.7001 762.7500 1414.5000 762.9000 ;
	    RECT 1143.9000 761.2500 1414.5000 762.7500 ;
	    RECT 1143.9000 761.1000 1145.7001 761.2500 ;
	    RECT 1309.5000 761.1000 1311.3000 761.2500 ;
	    RECT 1393.5000 761.1000 1395.3000 761.2500 ;
	    RECT 1412.7001 761.1000 1414.5000 761.2500 ;
	    RECT 1431.9000 762.7500 1433.7001 762.9000 ;
	    RECT 1439.1000 762.7500 1440.9000 762.9000 ;
	    RECT 1431.9000 761.2500 1440.9000 762.7500 ;
	    RECT 1431.9000 761.1000 1433.7001 761.2500 ;
	    RECT 1439.1000 761.1000 1440.9000 761.2500 ;
	    RECT 1482.3000 762.7500 1484.1000 762.9000 ;
	    RECT 1491.9000 762.7500 1493.7001 762.9000 ;
	    RECT 1482.3000 761.2500 1493.7001 762.7500 ;
	    RECT 1482.3000 761.1000 1484.1000 761.2500 ;
	    RECT 1491.9000 761.1000 1493.7001 761.2500 ;
	    RECT 1511.1000 762.7500 1512.9000 762.9000 ;
	    RECT 1537.5000 762.7500 1539.3000 762.9000 ;
	    RECT 1551.9000 762.7500 1553.7001 762.9000 ;
	    RECT 1511.1000 761.2500 1553.7001 762.7500 ;
	    RECT 1511.1000 761.1000 1512.9000 761.2500 ;
	    RECT 1537.5000 761.1000 1539.3000 761.2500 ;
	    RECT 1551.9000 761.1000 1553.7001 761.2500 ;
	    RECT 164.7000 756.7500 166.5000 756.9000 ;
	    RECT 171.9000 756.7500 173.7000 756.9000 ;
	    RECT 195.9000 756.7500 197.7000 756.9000 ;
	    RECT 164.7000 755.2500 197.7000 756.7500 ;
	    RECT 164.7000 755.1000 166.5000 755.2500 ;
	    RECT 171.9000 755.1000 173.7000 755.2500 ;
	    RECT 195.9000 755.1000 197.7000 755.2500 ;
	    RECT 231.9000 756.7500 233.7000 756.9000 ;
	    RECT 236.7000 756.7500 238.5000 756.9000 ;
	    RECT 231.9000 755.2500 238.5000 756.7500 ;
	    RECT 231.9000 755.1000 233.7000 755.2500 ;
	    RECT 236.7000 755.1000 238.5000 755.2500 ;
	    RECT 596.7000 756.7500 598.5000 756.9000 ;
	    RECT 639.9000 756.7500 641.7000 756.9000 ;
	    RECT 596.7000 755.2500 641.7000 756.7500 ;
	    RECT 596.7000 755.1000 598.5000 755.2500 ;
	    RECT 639.9000 755.1000 641.7000 755.2500 ;
	    RECT 747.9000 756.7500 749.7000 756.9000 ;
	    RECT 781.5000 756.7500 783.3000 756.9000 ;
	    RECT 839.1000 756.7500 840.9000 756.9000 ;
	    RECT 747.9000 755.2500 840.9000 756.7500 ;
	    RECT 747.9000 755.1000 749.7000 755.2500 ;
	    RECT 781.5000 755.1000 783.3000 755.2500 ;
	    RECT 839.1000 755.1000 840.9000 755.2500 ;
	    RECT 1004.7000 756.7500 1006.5000 756.9000 ;
	    RECT 1076.7001 756.7500 1078.5000 756.9000 ;
	    RECT 1004.7000 755.2500 1078.5000 756.7500 ;
	    RECT 1004.7000 755.1000 1006.5000 755.2500 ;
	    RECT 1076.7001 755.1000 1078.5000 755.2500 ;
	    RECT 1095.9000 756.7500 1097.7001 756.9000 ;
	    RECT 1100.7001 756.7500 1102.5000 756.9000 ;
	    RECT 1143.9000 756.7500 1145.7001 756.9000 ;
	    RECT 1095.9000 755.2500 1145.7001 756.7500 ;
	    RECT 1095.9000 755.1000 1097.7001 755.2500 ;
	    RECT 1100.7001 755.1000 1102.5000 755.2500 ;
	    RECT 1143.9000 755.1000 1145.7001 755.2500 ;
	    RECT 51.9000 750.7500 53.7000 750.9000 ;
	    RECT 176.7000 750.7500 178.5000 750.9000 ;
	    RECT 51.9000 749.2500 178.5000 750.7500 ;
	    RECT 51.9000 749.1000 53.7000 749.2500 ;
	    RECT 176.7000 749.1000 178.5000 749.2500 ;
	    RECT 193.5000 750.7500 195.3000 750.9000 ;
	    RECT 217.5000 750.7500 219.3000 750.9000 ;
	    RECT 193.5000 749.2500 219.3000 750.7500 ;
	    RECT 193.5000 749.1000 195.3000 749.2500 ;
	    RECT 217.5000 749.1000 219.3000 749.2500 ;
	    RECT 231.9000 750.7500 233.7000 750.9000 ;
	    RECT 248.7000 750.7500 250.5000 750.9000 ;
	    RECT 231.9000 749.2500 250.5000 750.7500 ;
	    RECT 231.9000 749.1000 233.7000 749.2500 ;
	    RECT 248.7000 749.1000 250.5000 749.2500 ;
	    RECT 361.5000 750.7500 363.3000 750.9000 ;
	    RECT 431.1000 750.7500 432.9000 750.9000 ;
	    RECT 361.5000 749.2500 432.9000 750.7500 ;
	    RECT 361.5000 749.1000 363.3000 749.2500 ;
	    RECT 431.1000 749.1000 432.9000 749.2500 ;
	    RECT 507.9000 750.7500 509.7000 750.9000 ;
	    RECT 539.1000 750.7500 540.9000 750.9000 ;
	    RECT 507.9000 749.2500 540.9000 750.7500 ;
	    RECT 507.9000 749.1000 509.7000 749.2500 ;
	    RECT 539.1000 749.1000 540.9000 749.2500 ;
	    RECT 603.9000 750.7500 605.7000 750.9000 ;
	    RECT 615.9000 750.7500 617.7000 750.9000 ;
	    RECT 603.9000 749.2500 617.7000 750.7500 ;
	    RECT 603.9000 749.1000 605.7000 749.2500 ;
	    RECT 615.9000 749.1000 617.7000 749.2500 ;
	    RECT 661.5000 750.7500 663.3000 750.9000 ;
	    RECT 699.9000 750.7500 701.7000 750.9000 ;
	    RECT 661.5000 749.2500 701.7000 750.7500 ;
	    RECT 661.5000 749.1000 663.3000 749.2500 ;
	    RECT 699.9000 749.1000 701.7000 749.2500 ;
	    RECT 807.9000 750.7500 809.7000 750.9000 ;
	    RECT 827.1000 750.7500 828.9000 750.9000 ;
	    RECT 807.9000 749.2500 828.9000 750.7500 ;
	    RECT 807.9000 749.1000 809.7000 749.2500 ;
	    RECT 827.1000 749.1000 828.9000 749.2500 ;
	    RECT 831.9000 750.7500 833.7000 750.9000 ;
	    RECT 839.1000 750.7500 840.9000 750.9000 ;
	    RECT 831.9000 749.2500 840.9000 750.7500 ;
	    RECT 831.9000 749.1000 833.7000 749.2500 ;
	    RECT 839.1000 749.1000 840.9000 749.2500 ;
	    RECT 1076.7001 750.7500 1078.5000 750.9000 ;
	    RECT 1117.5000 750.7500 1119.3000 750.9000 ;
	    RECT 1076.7001 749.2500 1119.3000 750.7500 ;
	    RECT 1076.7001 749.1000 1078.5000 749.2500 ;
	    RECT 1117.5000 749.1000 1119.3000 749.2500 ;
	    RECT 1199.1000 750.7500 1200.9000 750.9000 ;
	    RECT 1211.1000 750.7500 1212.9000 750.9000 ;
	    RECT 1199.1000 749.2500 1212.9000 750.7500 ;
	    RECT 1199.1000 749.1000 1200.9000 749.2500 ;
	    RECT 1211.1000 749.1000 1212.9000 749.2500 ;
	    RECT 1410.3000 750.7500 1412.1000 750.9000 ;
	    RECT 1419.9000 750.7500 1421.7001 750.9000 ;
	    RECT 1410.3000 749.2500 1421.7001 750.7500 ;
	    RECT 1410.3000 749.1000 1412.1000 749.2500 ;
	    RECT 1419.9000 749.1000 1421.7001 749.2500 ;
	    RECT 1518.3000 750.7500 1520.1000 750.9000 ;
	    RECT 1549.5000 750.7500 1551.3000 750.9000 ;
	    RECT 1518.3000 749.2500 1551.3000 750.7500 ;
	    RECT 1518.3000 749.1000 1520.1000 749.2500 ;
	    RECT 1549.5000 749.1000 1551.3000 749.2500 ;
	    RECT 167.1000 744.7500 168.9000 744.9000 ;
	    RECT 251.1000 744.7500 252.9000 744.9000 ;
	    RECT 263.1000 744.7500 264.9000 744.9000 ;
	    RECT 167.1000 743.2500 264.9000 744.7500 ;
	    RECT 167.1000 743.1000 168.9000 743.2500 ;
	    RECT 251.1000 743.1000 252.9000 743.2500 ;
	    RECT 263.1000 743.1000 264.9000 743.2500 ;
	    RECT 445.5000 744.7500 447.3000 744.9000 ;
	    RECT 510.3000 744.7500 512.1000 744.9000 ;
	    RECT 445.5000 743.2500 512.1000 744.7500 ;
	    RECT 445.5000 743.1000 447.3000 743.2500 ;
	    RECT 510.3000 743.1000 512.1000 743.2500 ;
	    RECT 673.5000 744.7500 675.3000 744.9000 ;
	    RECT 687.9000 744.7500 689.7000 744.9000 ;
	    RECT 673.5000 743.2500 689.7000 744.7500 ;
	    RECT 673.5000 743.1000 675.3000 743.2500 ;
	    RECT 687.9000 743.1000 689.7000 743.2500 ;
	    RECT 774.3000 744.7500 776.1000 744.9000 ;
	    RECT 827.1000 744.7500 828.9000 744.9000 ;
	    RECT 774.3000 743.2500 828.9000 744.7500 ;
	    RECT 774.3000 743.1000 776.1000 743.2500 ;
	    RECT 827.1000 743.1000 828.9000 743.2500 ;
	    RECT 834.3000 744.7500 836.1000 744.9000 ;
	    RECT 887.1000 744.7500 888.9000 744.9000 ;
	    RECT 834.3000 743.2500 888.9000 744.7500 ;
	    RECT 834.3000 743.1000 836.1000 743.2500 ;
	    RECT 887.1000 743.1000 888.9000 743.2500 ;
	    RECT 999.9000 744.7500 1001.7000 744.9000 ;
	    RECT 1026.3000 744.7500 1028.1000 744.9000 ;
	    RECT 999.9000 743.2500 1028.1000 744.7500 ;
	    RECT 999.9000 743.1000 1001.7000 743.2500 ;
	    RECT 1026.3000 743.1000 1028.1000 743.2500 ;
	    RECT 1333.5000 744.7500 1335.3000 744.9000 ;
	    RECT 1424.7001 744.7500 1426.5000 744.9000 ;
	    RECT 1333.5000 743.2500 1426.5000 744.7500 ;
	    RECT 1333.5000 743.1000 1335.3000 743.2500 ;
	    RECT 1424.7001 743.1000 1426.5000 743.2500 ;
	    RECT 1484.7001 744.7500 1486.5000 744.9000 ;
	    RECT 1515.9000 744.7500 1517.7001 744.9000 ;
	    RECT 1551.9000 744.7500 1553.7001 744.9000 ;
	    RECT 1484.7001 743.2500 1553.7001 744.7500 ;
	    RECT 1484.7001 743.1000 1486.5000 743.2500 ;
	    RECT 1515.9000 743.1000 1517.7001 743.2500 ;
	    RECT 1551.9000 743.1000 1553.7001 743.2500 ;
	    RECT 164.7000 738.7500 166.5000 738.9000 ;
	    RECT 291.9000 738.7500 293.7000 738.9000 ;
	    RECT 423.9000 738.7500 425.7000 738.9000 ;
	    RECT 164.7000 737.2500 425.7000 738.7500 ;
	    RECT 164.7000 737.1000 166.5000 737.2500 ;
	    RECT 291.9000 737.1000 293.7000 737.2500 ;
	    RECT 423.9000 737.1000 425.7000 737.2500 ;
	    RECT 546.3000 738.7500 548.1000 738.9000 ;
	    RECT 567.9000 738.7500 569.7000 738.9000 ;
	    RECT 546.3000 737.2500 569.7000 738.7500 ;
	    RECT 546.3000 737.1000 548.1000 737.2500 ;
	    RECT 567.9000 737.1000 569.7000 737.2500 ;
	    RECT 594.3000 738.7500 596.1000 738.9000 ;
	    RECT 627.9000 738.7500 629.7000 738.9000 ;
	    RECT 594.3000 737.2500 629.7000 738.7500 ;
	    RECT 594.3000 737.1000 596.1000 737.2500 ;
	    RECT 627.9000 737.1000 629.7000 737.2500 ;
	    RECT 649.5000 738.7500 651.3000 738.9000 ;
	    RECT 690.3000 738.7500 692.1000 738.9000 ;
	    RECT 711.9000 738.7500 713.7000 738.9000 ;
	    RECT 721.5000 738.7500 723.3000 738.9000 ;
	    RECT 649.5000 737.2500 723.3000 738.7500 ;
	    RECT 649.5000 737.1000 651.3000 737.2500 ;
	    RECT 690.3000 737.1000 692.1000 737.2500 ;
	    RECT 711.9000 737.1000 713.7000 737.2500 ;
	    RECT 721.5000 737.1000 723.3000 737.2500 ;
	    RECT 733.5000 738.7500 735.3000 738.9000 ;
	    RECT 743.1000 738.7500 744.9000 738.9000 ;
	    RECT 747.9000 738.7500 749.7000 738.9000 ;
	    RECT 733.5000 737.2500 749.7000 738.7500 ;
	    RECT 733.5000 737.1000 735.3000 737.2500 ;
	    RECT 743.1000 737.1000 744.9000 737.2500 ;
	    RECT 747.9000 737.1000 749.7000 737.2500 ;
	    RECT 786.3000 738.7500 788.1000 738.9000 ;
	    RECT 795.9000 738.7500 797.7000 738.9000 ;
	    RECT 786.3000 737.2500 797.7000 738.7500 ;
	    RECT 786.3000 737.1000 788.1000 737.2500 ;
	    RECT 795.9000 737.1000 797.7000 737.2500 ;
	    RECT 1011.9000 738.7500 1013.7000 738.9000 ;
	    RECT 1052.7001 738.7500 1054.5000 738.9000 ;
	    RECT 1059.9000 738.7500 1061.7001 738.9000 ;
	    RECT 1011.9000 737.2500 1061.7001 738.7500 ;
	    RECT 1011.9000 737.1000 1013.7000 737.2500 ;
	    RECT 1052.7001 737.1000 1054.5000 737.2500 ;
	    RECT 1059.9000 737.1000 1061.7001 737.2500 ;
	    RECT 1105.5000 738.7500 1107.3000 738.9000 ;
	    RECT 1163.1000 738.7500 1164.9000 738.9000 ;
	    RECT 1191.9000 738.7500 1193.7001 738.9000 ;
	    RECT 1244.7001 738.7500 1246.5000 738.9000 ;
	    RECT 1105.5000 737.2500 1246.5000 738.7500 ;
	    RECT 1105.5000 737.1000 1107.3000 737.2500 ;
	    RECT 1163.1000 737.1000 1164.9000 737.2500 ;
	    RECT 1191.9000 737.1000 1193.7001 737.2500 ;
	    RECT 1244.7001 737.1000 1246.5000 737.2500 ;
	    RECT 1273.5000 738.7500 1275.3000 738.9000 ;
	    RECT 1297.5000 738.7500 1299.3000 738.9000 ;
	    RECT 1273.5000 737.2500 1299.3000 738.7500 ;
	    RECT 1273.5000 737.1000 1275.3000 737.2500 ;
	    RECT 1297.5000 737.1000 1299.3000 737.2500 ;
	    RECT 1374.3000 738.7500 1376.1000 738.9000 ;
	    RECT 1386.3000 738.7500 1388.1000 738.9000 ;
	    RECT 1374.3000 737.2500 1388.1000 738.7500 ;
	    RECT 1374.3000 737.1000 1376.1000 737.2500 ;
	    RECT 1386.3000 737.1000 1388.1000 737.2500 ;
	    RECT 1503.9000 738.7500 1505.7001 738.9000 ;
	    RECT 1523.1000 738.7500 1524.9000 738.9000 ;
	    RECT 1503.9000 737.2500 1524.9000 738.7500 ;
	    RECT 1503.9000 737.1000 1505.7001 737.2500 ;
	    RECT 1523.1000 737.1000 1524.9000 737.2500 ;
	    RECT 227.1000 732.7500 228.9000 732.9000 ;
	    RECT 248.7000 732.7500 250.5000 732.9000 ;
	    RECT 227.1000 731.2500 250.5000 732.7500 ;
	    RECT 227.1000 731.1000 228.9000 731.2500 ;
	    RECT 248.7000 731.1000 250.5000 731.2500 ;
	    RECT 577.5000 732.7500 579.3000 732.9000 ;
	    RECT 620.7000 732.7500 622.5000 732.9000 ;
	    RECT 577.5000 731.2500 622.5000 732.7500 ;
	    RECT 577.5000 731.1000 579.3000 731.2500 ;
	    RECT 620.7000 731.1000 622.5000 731.2500 ;
	    RECT 651.9000 732.7500 653.7000 732.9000 ;
	    RECT 659.1000 732.7500 660.9000 732.9000 ;
	    RECT 714.3000 732.7500 716.1000 732.9000 ;
	    RECT 651.9000 731.2500 716.1000 732.7500 ;
	    RECT 651.9000 731.1000 653.7000 731.2500 ;
	    RECT 659.1000 731.1000 660.9000 731.2500 ;
	    RECT 714.3000 731.1000 716.1000 731.2500 ;
	    RECT 745.5000 732.7500 747.3000 732.9000 ;
	    RECT 750.3000 732.7500 752.1000 732.9000 ;
	    RECT 745.5000 731.2500 752.1000 732.7500 ;
	    RECT 745.5000 731.1000 747.3000 731.2500 ;
	    RECT 750.3000 731.1000 752.1000 731.2500 ;
	    RECT 774.3000 732.7500 776.1000 732.9000 ;
	    RECT 798.3000 732.7500 800.1000 732.9000 ;
	    RECT 774.3000 731.2500 800.1000 732.7500 ;
	    RECT 774.3000 731.1000 776.1000 731.2500 ;
	    RECT 798.3000 731.1000 800.1000 731.2500 ;
	    RECT 906.3000 732.7500 908.1000 732.9000 ;
	    RECT 915.9000 732.7500 917.7000 732.9000 ;
	    RECT 906.3000 731.2500 917.7000 732.7500 ;
	    RECT 906.3000 731.1000 908.1000 731.2500 ;
	    RECT 915.9000 731.1000 917.7000 731.2500 ;
	    RECT 995.1000 732.7500 996.9000 732.9000 ;
	    RECT 1038.3000 732.7500 1040.1000 732.9000 ;
	    RECT 1105.5000 732.7500 1107.3000 732.9000 ;
	    RECT 995.1000 731.2500 1107.3000 732.7500 ;
	    RECT 995.1000 731.1000 996.9000 731.2500 ;
	    RECT 1038.3000 731.1000 1040.1000 731.2500 ;
	    RECT 1105.5000 731.1000 1107.3000 731.2500 ;
	    RECT 1163.1000 732.7500 1164.9000 732.9000 ;
	    RECT 1280.7001 732.7500 1282.5000 732.9000 ;
	    RECT 1163.1000 731.2500 1282.5000 732.7500 ;
	    RECT 1163.1000 731.1000 1164.9000 731.2500 ;
	    RECT 1280.7001 731.1000 1282.5000 731.2500 ;
	    RECT 1331.1000 732.7500 1332.9000 732.9000 ;
	    RECT 1369.5000 732.7500 1371.3000 732.9000 ;
	    RECT 1331.1000 731.2500 1371.3000 732.7500 ;
	    RECT 1331.1000 731.1000 1332.9000 731.2500 ;
	    RECT 1369.5000 731.1000 1371.3000 731.2500 ;
	    RECT 1460.7001 732.7500 1462.5000 732.9000 ;
	    RECT 1491.9000 732.7500 1493.7001 732.9000 ;
	    RECT 1554.3000 732.7500 1556.1000 732.9000 ;
	    RECT 1460.7001 731.2500 1556.1000 732.7500 ;
	    RECT 1460.7001 731.1000 1462.5000 731.2500 ;
	    RECT 1491.9000 731.1000 1493.7001 731.2500 ;
	    RECT 1554.3000 731.1000 1556.1000 731.2500 ;
	    RECT 157.5000 726.7500 159.3000 726.9000 ;
	    RECT 171.9000 726.7500 173.7000 726.9000 ;
	    RECT 157.5000 725.2500 173.7000 726.7500 ;
	    RECT 157.5000 725.1000 159.3000 725.2500 ;
	    RECT 171.9000 725.1000 173.7000 725.2500 ;
	    RECT 315.9000 726.7500 317.7000 726.9000 ;
	    RECT 371.1000 726.7500 372.9000 726.9000 ;
	    RECT 404.7000 726.7500 406.5000 726.9000 ;
	    RECT 315.9000 725.2500 406.5000 726.7500 ;
	    RECT 315.9000 725.1000 317.7000 725.2500 ;
	    RECT 371.1000 725.1000 372.9000 725.2500 ;
	    RECT 404.7000 725.1000 406.5000 725.2500 ;
	    RECT 695.1000 726.7500 696.9000 726.9000 ;
	    RECT 740.7000 726.7500 742.5000 726.9000 ;
	    RECT 695.1000 725.2500 742.5000 726.7500 ;
	    RECT 695.1000 725.1000 696.9000 725.2500 ;
	    RECT 740.7000 725.1000 742.5000 725.2500 ;
	    RECT 822.3000 726.7500 824.1000 726.9000 ;
	    RECT 855.9000 726.7500 857.7000 726.9000 ;
	    RECT 822.3000 725.2500 857.7000 726.7500 ;
	    RECT 822.3000 725.1000 824.1000 725.2500 ;
	    RECT 855.9000 725.1000 857.7000 725.2500 ;
	    RECT 1242.3000 726.7500 1244.1000 726.9000 ;
	    RECT 1299.9000 726.7500 1301.7001 726.9000 ;
	    RECT 1307.1000 726.7500 1308.9000 726.9000 ;
	    RECT 1242.3000 725.2500 1308.9000 726.7500 ;
	    RECT 1242.3000 725.1000 1244.1000 725.2500 ;
	    RECT 1299.9000 725.1000 1301.7001 725.2500 ;
	    RECT 1307.1000 725.1000 1308.9000 725.2500 ;
	    RECT 1410.3000 726.7500 1412.1000 726.9000 ;
	    RECT 1455.9000 726.7500 1457.7001 726.9000 ;
	    RECT 1410.3000 725.2500 1457.7001 726.7500 ;
	    RECT 1410.3000 725.1000 1412.1000 725.2500 ;
	    RECT 1455.9000 725.1000 1457.7001 725.2500 ;
	    RECT 123.9000 720.7500 125.7000 720.9000 ;
	    RECT 162.3000 720.7500 164.1000 720.9000 ;
	    RECT 123.9000 719.2500 164.1000 720.7500 ;
	    RECT 123.9000 719.1000 125.7000 719.2500 ;
	    RECT 162.3000 719.1000 164.1000 719.2500 ;
	    RECT 253.5000 720.7500 255.3000 720.9000 ;
	    RECT 289.5000 720.7500 291.3000 720.9000 ;
	    RECT 253.5000 719.2500 291.3000 720.7500 ;
	    RECT 253.5000 719.1000 255.3000 719.2500 ;
	    RECT 289.5000 719.1000 291.3000 719.2500 ;
	    RECT 575.1000 720.7500 576.9000 720.9000 ;
	    RECT 623.1000 720.7500 624.9000 720.9000 ;
	    RECT 575.1000 719.2500 624.9000 720.7500 ;
	    RECT 575.1000 719.1000 576.9000 719.2500 ;
	    RECT 623.1000 719.1000 624.9000 719.2500 ;
	    RECT 704.7000 720.7500 706.5000 720.9000 ;
	    RECT 728.7000 720.7500 730.5000 720.9000 ;
	    RECT 704.7000 719.2500 730.5000 720.7500 ;
	    RECT 704.7000 719.1000 706.5000 719.2500 ;
	    RECT 728.7000 719.1000 730.5000 719.2500 ;
	    RECT 743.1000 720.7500 744.9000 720.9000 ;
	    RECT 779.1000 720.7500 780.9000 720.9000 ;
	    RECT 793.5000 720.7500 795.3000 720.9000 ;
	    RECT 743.1000 719.2500 795.3000 720.7500 ;
	    RECT 743.1000 719.1000 744.9000 719.2500 ;
	    RECT 779.1000 719.1000 780.9000 719.2500 ;
	    RECT 793.5000 719.1000 795.3000 719.2500 ;
	    RECT 827.1000 720.7500 828.9000 720.9000 ;
	    RECT 915.9000 720.7500 917.7000 720.9000 ;
	    RECT 827.1000 719.2500 917.7000 720.7500 ;
	    RECT 827.1000 719.1000 828.9000 719.2500 ;
	    RECT 915.9000 719.1000 917.7000 719.2500 ;
	    RECT 1026.3000 720.7500 1028.1000 720.9000 ;
	    RECT 1057.5000 720.7500 1059.3000 720.9000 ;
	    RECT 1026.3000 719.2500 1059.3000 720.7500 ;
	    RECT 1026.3000 719.1000 1028.1000 719.2500 ;
	    RECT 1057.5000 719.1000 1059.3000 719.2500 ;
	    RECT 1506.3000 720.7500 1508.1000 720.9000 ;
	    RECT 1542.3000 720.7500 1544.1000 720.9000 ;
	    RECT 1506.3000 719.2500 1544.1000 720.7500 ;
	    RECT 1506.3000 719.1000 1508.1000 719.2500 ;
	    RECT 1542.3000 719.1000 1544.1000 719.2500 ;
	    RECT 1561.5000 720.7500 1563.3000 720.9000 ;
	    RECT 1566.3000 720.7500 1568.1000 720.9000 ;
	    RECT 1561.5000 719.2500 1568.1000 720.7500 ;
	    RECT 1561.5000 719.1000 1563.3000 719.2500 ;
	    RECT 1566.3000 719.1000 1568.1000 719.2500 ;
	    RECT 18.3000 714.7500 20.1000 714.9000 ;
	    RECT 123.9000 714.7500 125.7000 714.9000 ;
	    RECT 18.3000 713.2500 125.7000 714.7500 ;
	    RECT 18.3000 713.1000 20.1000 713.2500 ;
	    RECT 123.9000 713.1000 125.7000 713.2500 ;
	    RECT 140.7000 714.7500 142.5000 714.9000 ;
	    RECT 191.1000 714.7500 192.9000 714.9000 ;
	    RECT 140.7000 713.2500 192.9000 714.7500 ;
	    RECT 140.7000 713.1000 142.5000 713.2500 ;
	    RECT 191.1000 713.1000 192.9000 713.2500 ;
	    RECT 205.5000 714.7500 207.3000 714.9000 ;
	    RECT 255.9000 714.7500 257.7000 714.9000 ;
	    RECT 205.5000 713.2500 257.7000 714.7500 ;
	    RECT 205.5000 713.1000 207.3000 713.2500 ;
	    RECT 255.9000 713.1000 257.7000 713.2500 ;
	    RECT 265.5000 714.7500 267.3000 714.9000 ;
	    RECT 347.1000 714.7500 348.9000 714.9000 ;
	    RECT 265.5000 713.2500 348.9000 714.7500 ;
	    RECT 265.5000 713.1000 267.3000 713.2500 ;
	    RECT 347.1000 713.1000 348.9000 713.2500 ;
	    RECT 459.9000 714.7500 461.7000 714.9000 ;
	    RECT 635.1000 714.7500 636.9000 714.9000 ;
	    RECT 459.9000 713.2500 636.9000 714.7500 ;
	    RECT 459.9000 713.1000 461.7000 713.2500 ;
	    RECT 635.1000 713.1000 636.9000 713.2500 ;
	    RECT 678.3000 714.7500 680.1000 714.9000 ;
	    RECT 723.9000 714.7500 725.7000 714.9000 ;
	    RECT 678.3000 713.2500 725.7000 714.7500 ;
	    RECT 678.3000 713.1000 680.1000 713.2500 ;
	    RECT 723.9000 713.1000 725.7000 713.2500 ;
	    RECT 762.3000 714.7500 764.1000 714.9000 ;
	    RECT 781.5000 714.7500 783.3000 714.9000 ;
	    RECT 762.3000 713.2500 783.3000 714.7500 ;
	    RECT 762.3000 713.1000 764.1000 713.2500 ;
	    RECT 781.5000 713.1000 783.3000 713.2500 ;
	    RECT 791.1000 714.7500 792.9000 714.9000 ;
	    RECT 810.3000 714.7500 812.1000 714.9000 ;
	    RECT 817.5000 714.7500 819.3000 714.9000 ;
	    RECT 791.1000 713.2500 819.3000 714.7500 ;
	    RECT 791.1000 713.1000 792.9000 713.2500 ;
	    RECT 810.3000 713.1000 812.1000 713.2500 ;
	    RECT 817.5000 713.1000 819.3000 713.2500 ;
	    RECT 822.3000 714.7500 824.1000 714.9000 ;
	    RECT 879.9000 714.7500 881.7000 714.9000 ;
	    RECT 822.3000 713.2500 881.7000 714.7500 ;
	    RECT 822.3000 713.1000 824.1000 713.2500 ;
	    RECT 879.9000 713.1000 881.7000 713.2500 ;
	    RECT 887.1000 714.7500 888.9000 714.9000 ;
	    RECT 913.5000 714.7500 915.3000 714.9000 ;
	    RECT 887.1000 713.2500 915.3000 714.7500 ;
	    RECT 887.1000 713.1000 888.9000 713.2500 ;
	    RECT 913.5000 713.1000 915.3000 713.2500 ;
	    RECT 985.5000 714.7500 987.3000 714.9000 ;
	    RECT 1081.5000 714.7500 1083.3000 714.9000 ;
	    RECT 985.5000 713.2500 1083.3000 714.7500 ;
	    RECT 985.5000 713.1000 987.3000 713.2500 ;
	    RECT 1081.5000 713.1000 1083.3000 713.2500 ;
	    RECT 1179.9000 714.7500 1181.7001 714.9000 ;
	    RECT 1196.7001 714.7500 1198.5000 714.9000 ;
	    RECT 1179.9000 713.2500 1198.5000 714.7500 ;
	    RECT 1179.9000 713.1000 1181.7001 713.2500 ;
	    RECT 1196.7001 713.1000 1198.5000 713.2500 ;
	    RECT 1299.9000 714.7500 1301.7001 714.9000 ;
	    RECT 1350.3000 714.7500 1352.1000 714.9000 ;
	    RECT 1299.9000 713.2500 1352.1000 714.7500 ;
	    RECT 1299.9000 713.1000 1301.7001 713.2500 ;
	    RECT 1350.3000 713.1000 1352.1000 713.2500 ;
	    RECT 1415.1000 714.7500 1416.9000 714.9000 ;
	    RECT 1458.3000 714.7500 1460.1000 714.9000 ;
	    RECT 1415.1000 713.2500 1460.1000 714.7500 ;
	    RECT 1415.1000 713.1000 1416.9000 713.2500 ;
	    RECT 1458.3000 713.1000 1460.1000 713.2500 ;
	    RECT 188.7000 708.7500 190.5000 708.9000 ;
	    RECT 172.0500 707.2500 190.5000 708.7500 ;
	    RECT 172.0500 702.9000 173.5500 707.2500 ;
	    RECT 188.7000 707.1000 190.5000 707.2500 ;
	    RECT 193.5000 708.7500 195.3000 708.9000 ;
	    RECT 205.5000 708.7500 207.3000 708.9000 ;
	    RECT 193.5000 707.2500 207.3000 708.7500 ;
	    RECT 193.5000 707.1000 195.3000 707.2500 ;
	    RECT 205.5000 707.1000 207.3000 707.2500 ;
	    RECT 347.1000 708.7500 348.9000 708.9000 ;
	    RECT 368.7000 708.7500 370.5000 708.9000 ;
	    RECT 347.1000 707.2500 370.5000 708.7500 ;
	    RECT 347.1000 707.1000 348.9000 707.2500 ;
	    RECT 368.7000 707.1000 370.5000 707.2500 ;
	    RECT 411.9000 708.7500 413.7000 708.9000 ;
	    RECT 419.1000 708.7500 420.9000 708.9000 ;
	    RECT 411.9000 707.2500 420.9000 708.7500 ;
	    RECT 411.9000 707.1000 413.7000 707.2500 ;
	    RECT 419.1000 707.1000 420.9000 707.2500 ;
	    RECT 601.5000 708.7500 603.3000 708.9000 ;
	    RECT 618.3000 708.7500 620.1000 708.9000 ;
	    RECT 647.1000 708.7500 648.9000 708.9000 ;
	    RECT 601.5000 707.2500 648.9000 708.7500 ;
	    RECT 601.5000 707.1000 603.3000 707.2500 ;
	    RECT 618.3000 707.1000 620.1000 707.2500 ;
	    RECT 647.1000 707.1000 648.9000 707.2500 ;
	    RECT 714.3000 708.7500 716.1000 708.9000 ;
	    RECT 738.3000 708.7500 740.1000 708.9000 ;
	    RECT 771.9000 708.7500 773.7000 708.9000 ;
	    RECT 714.3000 707.2500 773.7000 708.7500 ;
	    RECT 714.3000 707.1000 716.1000 707.2500 ;
	    RECT 738.3000 707.1000 740.1000 707.2500 ;
	    RECT 771.9000 707.1000 773.7000 707.2500 ;
	    RECT 798.3000 708.7500 800.1000 708.9000 ;
	    RECT 812.7000 708.7500 814.5000 708.9000 ;
	    RECT 798.3000 707.2500 814.5000 708.7500 ;
	    RECT 798.3000 707.1000 800.1000 707.2500 ;
	    RECT 812.7000 707.1000 814.5000 707.2500 ;
	    RECT 817.5000 708.7500 819.3000 708.9000 ;
	    RECT 853.5000 708.7500 855.3000 708.9000 ;
	    RECT 817.5000 707.2500 855.3000 708.7500 ;
	    RECT 817.5000 707.1000 819.3000 707.2500 ;
	    RECT 853.5000 707.1000 855.3000 707.2500 ;
	    RECT 870.3000 708.7500 872.1000 708.9000 ;
	    RECT 918.3000 708.7500 920.1000 708.9000 ;
	    RECT 870.3000 707.2500 920.1000 708.7500 ;
	    RECT 870.3000 707.1000 872.1000 707.2500 ;
	    RECT 918.3000 707.1000 920.1000 707.2500 ;
	    RECT 944.7000 708.7500 946.5000 708.9000 ;
	    RECT 975.9000 708.7500 977.7000 708.9000 ;
	    RECT 944.7000 707.2500 977.7000 708.7500 ;
	    RECT 944.7000 707.1000 946.5000 707.2500 ;
	    RECT 975.9000 707.1000 977.7000 707.2500 ;
	    RECT 980.7000 708.7500 982.5000 708.9000 ;
	    RECT 1206.3000 708.7500 1208.1000 708.9000 ;
	    RECT 980.7000 707.2500 1208.1000 708.7500 ;
	    RECT 980.7000 707.1000 982.5000 707.2500 ;
	    RECT 1206.3000 707.1000 1208.1000 707.2500 ;
	    RECT 1297.5000 708.7500 1299.3000 708.9000 ;
	    RECT 1333.5000 708.7500 1335.3000 708.9000 ;
	    RECT 1297.5000 707.2500 1335.3000 708.7500 ;
	    RECT 1297.5000 707.1000 1299.3000 707.2500 ;
	    RECT 1333.5000 707.1000 1335.3000 707.2500 ;
	    RECT 1386.3000 708.7500 1388.1000 708.9000 ;
	    RECT 1393.5000 708.7500 1395.3000 708.9000 ;
	    RECT 1386.3000 707.2500 1395.3000 708.7500 ;
	    RECT 1386.3000 707.1000 1388.1000 707.2500 ;
	    RECT 1393.5000 707.1000 1395.3000 707.2500 ;
	    RECT 1419.9000 708.7500 1421.7001 708.9000 ;
	    RECT 1434.3000 708.7500 1436.1000 708.9000 ;
	    RECT 1419.9000 707.2500 1436.1000 708.7500 ;
	    RECT 1419.9000 707.1000 1421.7001 707.2500 ;
	    RECT 1434.3000 707.1000 1436.1000 707.2500 ;
	    RECT 1479.9000 708.7500 1481.7001 708.9000 ;
	    RECT 1511.1000 708.7500 1512.9000 708.9000 ;
	    RECT 1479.9000 707.2500 1512.9000 708.7500 ;
	    RECT 1479.9000 707.1000 1481.7001 707.2500 ;
	    RECT 1511.1000 707.1000 1512.9000 707.2500 ;
	    RECT 102.3000 702.7500 104.1000 702.9000 ;
	    RECT 123.9000 702.7500 125.7000 702.9000 ;
	    RECT 102.3000 701.2500 125.7000 702.7500 ;
	    RECT 102.3000 701.1000 104.1000 701.2500 ;
	    RECT 123.9000 701.1000 125.7000 701.2500 ;
	    RECT 147.9000 702.7500 149.7000 702.9000 ;
	    RECT 164.7000 702.7500 166.5000 702.9000 ;
	    RECT 147.9000 701.2500 166.5000 702.7500 ;
	    RECT 147.9000 701.1000 149.7000 701.2500 ;
	    RECT 164.7000 701.1000 166.5000 701.2500 ;
	    RECT 169.5000 701.2500 173.5500 702.9000 ;
	    RECT 176.7000 702.7500 178.5000 702.9000 ;
	    RECT 217.5000 702.7500 219.3000 702.9000 ;
	    RECT 231.9000 702.7500 233.7000 702.9000 ;
	    RECT 176.7000 701.2500 233.7000 702.7500 ;
	    RECT 169.5000 701.1000 172.8000 701.2500 ;
	    RECT 176.7000 701.1000 178.5000 701.2500 ;
	    RECT 217.5000 701.1000 219.3000 701.2500 ;
	    RECT 231.9000 701.1000 233.7000 701.2500 ;
	    RECT 239.1000 702.7500 240.9000 702.9000 ;
	    RECT 251.1000 702.7500 252.9000 702.9000 ;
	    RECT 239.1000 701.2500 252.9000 702.7500 ;
	    RECT 239.1000 701.1000 240.9000 701.2500 ;
	    RECT 251.1000 701.1000 252.9000 701.2500 ;
	    RECT 270.3000 702.7500 272.1000 702.9000 ;
	    RECT 339.9000 702.7500 341.7000 702.9000 ;
	    RECT 270.3000 701.2500 341.7000 702.7500 ;
	    RECT 270.3000 701.1000 272.1000 701.2500 ;
	    RECT 339.9000 701.1000 341.7000 701.2500 ;
	    RECT 414.3000 702.7500 416.1000 702.9000 ;
	    RECT 421.5000 702.7500 423.3000 702.9000 ;
	    RECT 414.3000 701.2500 423.3000 702.7500 ;
	    RECT 414.3000 701.1000 416.1000 701.2500 ;
	    RECT 421.5000 701.1000 423.3000 701.2500 ;
	    RECT 587.1000 702.7500 588.9000 702.9000 ;
	    RECT 603.9000 702.7500 605.7000 702.9000 ;
	    RECT 587.1000 701.2500 605.7000 702.7500 ;
	    RECT 587.1000 701.1000 588.9000 701.2500 ;
	    RECT 603.9000 701.1000 605.7000 701.2500 ;
	    RECT 613.5000 702.7500 615.3000 702.9000 ;
	    RECT 637.5000 702.7500 639.3000 702.9000 ;
	    RECT 613.5000 701.2500 639.3000 702.7500 ;
	    RECT 613.5000 701.1000 615.3000 701.2500 ;
	    RECT 637.5000 701.1000 639.3000 701.2500 ;
	    RECT 671.1000 702.7500 672.9000 702.9000 ;
	    RECT 678.3000 702.7500 680.1000 702.9000 ;
	    RECT 671.1000 701.2500 680.1000 702.7500 ;
	    RECT 671.1000 701.1000 672.9000 701.2500 ;
	    RECT 678.3000 701.1000 680.1000 701.2500 ;
	    RECT 740.7000 702.7500 742.5000 702.9000 ;
	    RECT 774.3000 702.7500 776.1000 702.9000 ;
	    RECT 740.7000 701.2500 776.1000 702.7500 ;
	    RECT 740.7000 701.1000 742.5000 701.2500 ;
	    RECT 774.3000 701.1000 776.1000 701.2500 ;
	    RECT 798.3000 702.7500 800.1000 702.9000 ;
	    RECT 803.1000 702.7500 804.9000 702.9000 ;
	    RECT 798.3000 701.2500 804.9000 702.7500 ;
	    RECT 798.3000 701.1000 800.1000 701.2500 ;
	    RECT 803.1000 701.1000 804.9000 701.2500 ;
	    RECT 807.9000 702.7500 809.7000 702.9000 ;
	    RECT 829.5000 702.7500 831.3000 702.9000 ;
	    RECT 807.9000 701.2500 831.3000 702.7500 ;
	    RECT 807.9000 701.1000 809.7000 701.2500 ;
	    RECT 829.5000 701.1000 831.3000 701.2500 ;
	    RECT 846.3000 702.7500 848.1000 702.9000 ;
	    RECT 875.1000 702.7500 876.9000 702.9000 ;
	    RECT 846.3000 701.2500 876.9000 702.7500 ;
	    RECT 846.3000 701.1000 848.1000 701.2500 ;
	    RECT 875.1000 701.1000 876.9000 701.2500 ;
	    RECT 918.3000 702.7500 920.1000 702.9000 ;
	    RECT 968.7000 702.7500 970.5000 702.9000 ;
	    RECT 918.3000 701.2500 970.5000 702.7500 ;
	    RECT 918.3000 701.1000 920.1000 701.2500 ;
	    RECT 968.7000 701.1000 970.5000 701.2500 ;
	    RECT 1304.7001 702.7500 1306.5000 702.9000 ;
	    RECT 1309.5000 702.7500 1311.3000 702.9000 ;
	    RECT 1304.7001 701.2500 1311.3000 702.7500 ;
	    RECT 1304.7001 701.1000 1306.5000 701.2500 ;
	    RECT 1309.5000 701.1000 1311.3000 701.2500 ;
	    RECT 1434.3000 702.7500 1436.1000 702.9000 ;
	    RECT 1441.5000 702.7500 1443.3000 702.9000 ;
	    RECT 1451.1000 702.7500 1452.9000 702.9000 ;
	    RECT 1434.3000 701.2500 1452.9000 702.7500 ;
	    RECT 1434.3000 701.1000 1436.1000 701.2500 ;
	    RECT 1441.5000 701.1000 1443.3000 701.2500 ;
	    RECT 1451.1000 701.1000 1452.9000 701.2500 ;
	    RECT 1458.3000 702.7500 1460.1000 702.9000 ;
	    RECT 1463.1000 702.7500 1464.9000 702.9000 ;
	    RECT 1458.3000 701.2500 1464.9000 702.7500 ;
	    RECT 1458.3000 701.1000 1460.1000 701.2500 ;
	    RECT 1463.1000 701.1000 1464.9000 701.2500 ;
	    RECT 95.1000 696.7500 96.9000 696.9000 ;
	    RECT 147.9000 696.7500 149.7000 696.9000 ;
	    RECT 95.1000 695.2500 149.7000 696.7500 ;
	    RECT 95.1000 695.1000 96.9000 695.2500 ;
	    RECT 147.9000 695.1000 149.7000 695.2500 ;
	    RECT 155.1000 696.7500 156.9000 696.9000 ;
	    RECT 191.1000 696.7500 192.9000 696.9000 ;
	    RECT 155.1000 695.2500 192.9000 696.7500 ;
	    RECT 155.1000 695.1000 156.9000 695.2500 ;
	    RECT 191.1000 695.1000 192.9000 695.2500 ;
	    RECT 212.7000 696.7500 214.5000 696.9000 ;
	    RECT 246.3000 696.7500 248.1000 696.9000 ;
	    RECT 212.7000 695.2500 248.1000 696.7500 ;
	    RECT 212.7000 695.1000 214.5000 695.2500 ;
	    RECT 246.3000 695.1000 248.1000 695.2500 ;
	    RECT 311.1000 696.7500 312.9000 696.9000 ;
	    RECT 318.3000 696.7500 320.1000 696.9000 ;
	    RECT 311.1000 695.2500 320.1000 696.7500 ;
	    RECT 311.1000 695.1000 312.9000 695.2500 ;
	    RECT 318.3000 695.1000 320.1000 695.2500 ;
	    RECT 419.1000 696.7500 420.9000 696.9000 ;
	    RECT 447.9000 696.7500 449.7000 696.9000 ;
	    RECT 419.1000 695.2500 449.7000 696.7500 ;
	    RECT 419.1000 695.1000 420.9000 695.2500 ;
	    RECT 447.9000 695.1000 449.7000 695.2500 ;
	    RECT 589.5000 696.7500 591.3000 696.9000 ;
	    RECT 599.1000 696.7500 600.9000 696.9000 ;
	    RECT 589.5000 695.2500 600.9000 696.7500 ;
	    RECT 589.5000 695.1000 591.3000 695.2500 ;
	    RECT 599.1000 695.1000 600.9000 695.2500 ;
	    RECT 716.7000 696.7500 718.5000 696.9000 ;
	    RECT 723.9000 696.7500 725.7000 696.9000 ;
	    RECT 716.7000 695.2500 725.7000 696.7500 ;
	    RECT 716.7000 695.1000 718.5000 695.2500 ;
	    RECT 723.9000 695.1000 725.7000 695.2500 ;
	    RECT 771.9000 696.7500 773.7000 696.9000 ;
	    RECT 843.9000 696.7500 845.7000 696.9000 ;
	    RECT 771.9000 695.2500 845.7000 696.7500 ;
	    RECT 771.9000 695.1000 773.7000 695.2500 ;
	    RECT 843.9000 695.1000 845.7000 695.2500 ;
	    RECT 1451.1000 696.7500 1452.9000 696.9000 ;
	    RECT 1455.9000 696.7500 1457.7001 696.9000 ;
	    RECT 1451.1000 695.2500 1457.7001 696.7500 ;
	    RECT 1451.1000 695.1000 1452.9000 695.2500 ;
	    RECT 1455.9000 695.1000 1457.7001 695.2500 ;
	    RECT 1475.1000 696.7500 1476.9000 696.9000 ;
	    RECT 1520.7001 696.7500 1522.5000 696.9000 ;
	    RECT 1535.1000 696.7500 1536.9000 696.9000 ;
	    RECT 1475.1000 695.2500 1536.9000 696.7500 ;
	    RECT 1475.1000 695.1000 1476.9000 695.2500 ;
	    RECT 1520.7001 695.1000 1522.5000 695.2500 ;
	    RECT 1535.1000 695.1000 1536.9000 695.2500 ;
	    RECT 169.5000 690.7500 171.3000 690.9000 ;
	    RECT 195.9000 690.7500 197.7000 690.9000 ;
	    RECT 169.5000 689.2500 197.7000 690.7500 ;
	    RECT 169.5000 689.1000 171.3000 689.2500 ;
	    RECT 195.9000 689.1000 197.7000 689.2500 ;
	    RECT 224.7000 690.7500 226.5000 690.9000 ;
	    RECT 277.5000 690.7500 279.3000 690.9000 ;
	    RECT 224.7000 689.2500 279.3000 690.7500 ;
	    RECT 224.7000 689.1000 226.5000 689.2500 ;
	    RECT 277.5000 689.1000 279.3000 689.2500 ;
	    RECT 500.7000 690.7500 502.5000 690.9000 ;
	    RECT 507.9000 690.7500 509.7000 690.9000 ;
	    RECT 500.7000 689.2500 509.7000 690.7500 ;
	    RECT 500.7000 689.1000 502.5000 689.2500 ;
	    RECT 507.9000 689.1000 509.7000 689.2500 ;
	    RECT 515.1000 690.7500 516.9000 690.9000 ;
	    RECT 608.7000 690.7500 610.5000 690.9000 ;
	    RECT 515.1000 689.2500 610.5000 690.7500 ;
	    RECT 515.1000 689.1000 516.9000 689.2500 ;
	    RECT 608.7000 689.1000 610.5000 689.2500 ;
	    RECT 649.5000 690.7500 651.3000 690.9000 ;
	    RECT 716.7000 690.7500 718.5000 690.9000 ;
	    RECT 649.5000 689.2500 718.5000 690.7500 ;
	    RECT 649.5000 689.1000 651.3000 689.2500 ;
	    RECT 716.7000 689.1000 718.5000 689.2500 ;
	    RECT 723.9000 690.7500 725.7000 690.9000 ;
	    RECT 759.9000 690.7500 761.7000 690.9000 ;
	    RECT 723.9000 689.2500 761.7000 690.7500 ;
	    RECT 723.9000 689.1000 725.7000 689.2500 ;
	    RECT 759.9000 689.1000 761.7000 689.2500 ;
	    RECT 951.9000 690.7500 953.7000 690.9000 ;
	    RECT 1002.3000 690.7500 1004.1000 690.9000 ;
	    RECT 951.9000 689.2500 1004.1000 690.7500 ;
	    RECT 951.9000 689.1000 953.7000 689.2500 ;
	    RECT 1002.3000 689.1000 1004.1000 689.2500 ;
	    RECT 1199.1000 690.7500 1200.9000 690.9000 ;
	    RECT 1220.7001 690.7500 1222.5000 690.9000 ;
	    RECT 1199.1000 689.2500 1222.5000 690.7500 ;
	    RECT 1199.1000 689.1000 1200.9000 689.2500 ;
	    RECT 1220.7001 689.1000 1222.5000 689.2500 ;
	    RECT 1268.7001 690.7500 1270.5000 690.9000 ;
	    RECT 1309.5000 690.7500 1311.3000 690.9000 ;
	    RECT 1268.7001 689.2500 1311.3000 690.7500 ;
	    RECT 1268.7001 689.1000 1270.5000 689.2500 ;
	    RECT 1309.5000 689.1000 1311.3000 689.2500 ;
	    RECT 1439.1000 690.7500 1440.9000 690.9000 ;
	    RECT 1484.7001 690.7500 1486.5000 690.9000 ;
	    RECT 1439.1000 689.2500 1486.5000 690.7500 ;
	    RECT 1439.1000 689.1000 1440.9000 689.2500 ;
	    RECT 1484.7001 689.1000 1486.5000 689.2500 ;
	    RECT 212.7000 684.7500 214.5000 684.9000 ;
	    RECT 222.3000 684.7500 224.1000 684.9000 ;
	    RECT 212.7000 683.2500 224.1000 684.7500 ;
	    RECT 212.7000 683.1000 214.5000 683.2500 ;
	    RECT 222.3000 683.1000 224.1000 683.2500 ;
	    RECT 229.5000 684.7500 231.3000 684.9000 ;
	    RECT 251.1000 684.7500 252.9000 684.9000 ;
	    RECT 229.5000 683.2500 252.9000 684.7500 ;
	    RECT 229.5000 683.1000 231.3000 683.2500 ;
	    RECT 251.1000 683.1000 252.9000 683.2500 ;
	    RECT 272.7000 684.7500 274.5000 684.9000 ;
	    RECT 315.9000 684.7500 317.7000 684.9000 ;
	    RECT 272.7000 683.2500 317.7000 684.7500 ;
	    RECT 272.7000 683.1000 274.5000 683.2500 ;
	    RECT 315.9000 683.1000 317.7000 683.2500 ;
	    RECT 447.9000 684.7500 449.7000 684.9000 ;
	    RECT 606.3000 684.7500 608.1000 684.9000 ;
	    RECT 447.9000 683.2500 608.1000 684.7500 ;
	    RECT 447.9000 683.1000 449.7000 683.2500 ;
	    RECT 606.3000 683.1000 608.1000 683.2500 ;
	    RECT 642.3000 684.7500 644.1000 684.9000 ;
	    RECT 707.1000 684.7500 708.9000 684.9000 ;
	    RECT 731.1000 684.7500 732.9000 684.9000 ;
	    RECT 642.3000 683.2500 732.9000 684.7500 ;
	    RECT 642.3000 683.1000 644.1000 683.2500 ;
	    RECT 707.1000 683.1000 708.9000 683.2500 ;
	    RECT 731.1000 683.1000 732.9000 683.2500 ;
	    RECT 767.1000 684.7500 768.9000 684.9000 ;
	    RECT 795.9000 684.7500 797.7000 684.9000 ;
	    RECT 767.1000 683.2500 797.7000 684.7500 ;
	    RECT 767.1000 683.1000 768.9000 683.2500 ;
	    RECT 795.9000 683.1000 797.7000 683.2500 ;
	    RECT 944.7000 684.7500 946.5000 684.9000 ;
	    RECT 990.3000 684.7500 992.1000 684.9000 ;
	    RECT 944.7000 683.2500 992.1000 684.7500 ;
	    RECT 944.7000 683.1000 946.5000 683.2500 ;
	    RECT 990.3000 683.1000 992.1000 683.2500 ;
	    RECT 1220.7001 684.7500 1222.5000 684.9000 ;
	    RECT 1273.5000 684.7500 1275.3000 684.9000 ;
	    RECT 1220.7001 683.2500 1275.3000 684.7500 ;
	    RECT 1220.7001 683.1000 1222.5000 683.2500 ;
	    RECT 1273.5000 683.1000 1275.3000 683.2500 ;
	    RECT 1304.7001 684.7500 1306.5000 684.9000 ;
	    RECT 1364.7001 684.7500 1366.5000 684.9000 ;
	    RECT 1304.7001 683.2500 1366.5000 684.7500 ;
	    RECT 1304.7001 683.1000 1306.5000 683.2500 ;
	    RECT 1364.7001 683.1000 1366.5000 683.2500 ;
	    RECT 1482.3000 684.7500 1484.1000 684.9000 ;
	    RECT 1525.5000 684.7500 1527.3000 684.9000 ;
	    RECT 1482.3000 683.2500 1527.3000 684.7500 ;
	    RECT 1482.3000 683.1000 1484.1000 683.2500 ;
	    RECT 1525.5000 683.1000 1527.3000 683.2500 ;
	    RECT 92.7000 678.7500 94.5000 678.9000 ;
	    RECT 150.3000 678.7500 152.1000 678.9000 ;
	    RECT 92.7000 677.2500 152.1000 678.7500 ;
	    RECT 92.7000 677.1000 94.5000 677.2500 ;
	    RECT 150.3000 677.1000 152.1000 677.2500 ;
	    RECT 157.5000 678.7500 159.3000 678.9000 ;
	    RECT 215.1000 678.7500 216.9000 678.9000 ;
	    RECT 157.5000 677.2500 216.9000 678.7500 ;
	    RECT 157.5000 677.1000 159.3000 677.2500 ;
	    RECT 215.1000 677.1000 216.9000 677.2500 ;
	    RECT 219.9000 678.7500 221.7000 678.9000 ;
	    RECT 224.7000 678.7500 226.5000 678.9000 ;
	    RECT 219.9000 677.2500 226.5000 678.7500 ;
	    RECT 219.9000 677.1000 221.7000 677.2500 ;
	    RECT 224.7000 677.1000 226.5000 677.2500 ;
	    RECT 248.7000 678.7500 250.5000 678.9000 ;
	    RECT 275.1000 678.7500 276.9000 678.9000 ;
	    RECT 248.7000 677.2500 276.9000 678.7500 ;
	    RECT 248.7000 677.1000 250.5000 677.2500 ;
	    RECT 275.1000 677.1000 276.9000 677.2500 ;
	    RECT 582.3000 678.7500 584.1000 678.9000 ;
	    RECT 596.7000 678.7500 598.5000 678.9000 ;
	    RECT 582.3000 677.2500 598.5000 678.7500 ;
	    RECT 582.3000 677.1000 584.1000 677.2500 ;
	    RECT 596.7000 677.1000 598.5000 677.2500 ;
	    RECT 630.3000 678.7500 632.1000 678.9000 ;
	    RECT 692.7000 678.7500 694.5000 678.9000 ;
	    RECT 630.3000 677.2500 694.5000 678.7500 ;
	    RECT 630.3000 677.1000 632.1000 677.2500 ;
	    RECT 692.7000 677.1000 694.5000 677.2500 ;
	    RECT 716.7000 678.7500 718.5000 678.9000 ;
	    RECT 762.3000 678.7500 764.1000 678.9000 ;
	    RECT 716.7000 677.2500 764.1000 678.7500 ;
	    RECT 716.7000 677.1000 718.5000 677.2500 ;
	    RECT 762.3000 677.1000 764.1000 677.2500 ;
	    RECT 769.5000 678.7500 771.3000 678.9000 ;
	    RECT 863.1000 678.7500 864.9000 678.9000 ;
	    RECT 769.5000 677.2500 864.9000 678.7500 ;
	    RECT 769.5000 677.1000 771.3000 677.2500 ;
	    RECT 863.1000 677.1000 864.9000 677.2500 ;
	    RECT 944.7000 678.7500 946.5000 678.9000 ;
	    RECT 951.9000 678.7500 953.7000 678.9000 ;
	    RECT 944.7000 677.2500 953.7000 678.7500 ;
	    RECT 944.7000 677.1000 946.5000 677.2500 ;
	    RECT 951.9000 677.1000 953.7000 677.2500 ;
	    RECT 1203.9000 678.7500 1205.7001 678.9000 ;
	    RECT 1247.1000 678.7500 1248.9000 678.9000 ;
	    RECT 1203.9000 677.2500 1248.9000 678.7500 ;
	    RECT 1203.9000 677.1000 1205.7001 677.2500 ;
	    RECT 1247.1000 677.1000 1248.9000 677.2500 ;
	    RECT 1297.5000 678.7500 1299.3000 678.9000 ;
	    RECT 1386.3000 678.7500 1388.1000 678.9000 ;
	    RECT 1297.5000 677.2500 1388.1000 678.7500 ;
	    RECT 1297.5000 677.1000 1299.3000 677.2500 ;
	    RECT 1386.3000 677.1000 1388.1000 677.2500 ;
	    RECT 1467.9000 678.7500 1469.7001 678.9000 ;
	    RECT 1489.5000 678.7500 1491.3000 678.9000 ;
	    RECT 1467.9000 677.2500 1491.3000 678.7500 ;
	    RECT 1467.9000 677.1000 1469.7001 677.2500 ;
	    RECT 1489.5000 677.1000 1491.3000 677.2500 ;
	    RECT 152.7000 672.7500 154.5000 672.9000 ;
	    RECT 176.7000 672.7500 178.5000 672.9000 ;
	    RECT 152.7000 671.2500 178.5000 672.7500 ;
	    RECT 152.7000 671.1000 154.5000 671.2500 ;
	    RECT 176.7000 671.1000 178.5000 671.2500 ;
	    RECT 215.1000 672.7500 216.9000 672.9000 ;
	    RECT 260.7000 672.7500 262.5000 672.9000 ;
	    RECT 215.1000 671.2500 262.5000 672.7500 ;
	    RECT 215.1000 671.1000 216.9000 671.2500 ;
	    RECT 260.7000 671.1000 262.5000 671.2500 ;
	    RECT 431.1000 672.7500 432.9000 672.9000 ;
	    RECT 515.1000 672.7500 516.9000 672.9000 ;
	    RECT 431.1000 671.2500 516.9000 672.7500 ;
	    RECT 431.1000 671.1000 432.9000 671.2500 ;
	    RECT 515.1000 671.1000 516.9000 671.2500 ;
	    RECT 589.5000 672.7500 591.3000 672.9000 ;
	    RECT 611.1000 672.7500 612.9000 672.9000 ;
	    RECT 589.5000 671.2500 612.9000 672.7500 ;
	    RECT 589.5000 671.1000 591.3000 671.2500 ;
	    RECT 611.1000 671.1000 612.9000 671.2500 ;
	    RECT 651.9000 672.7500 653.7000 672.9000 ;
	    RECT 771.9000 672.7500 773.7000 672.9000 ;
	    RECT 651.9000 671.2500 773.7000 672.7500 ;
	    RECT 651.9000 671.1000 653.7000 671.2500 ;
	    RECT 771.9000 671.1000 773.7000 671.2500 ;
	    RECT 863.1000 672.7500 864.9000 672.9000 ;
	    RECT 944.7000 672.7500 946.5000 672.9000 ;
	    RECT 863.1000 671.2500 946.5000 672.7500 ;
	    RECT 863.1000 671.1000 864.9000 671.2500 ;
	    RECT 944.7000 671.1000 946.5000 671.2500 ;
	    RECT 954.3000 672.7500 956.1000 672.9000 ;
	    RECT 975.9000 672.7500 977.7000 672.9000 ;
	    RECT 954.3000 671.2500 977.7000 672.7500 ;
	    RECT 954.3000 671.1000 956.1000 671.2500 ;
	    RECT 975.9000 671.1000 977.7000 671.2500 ;
	    RECT 1110.3000 672.7500 1112.1000 672.9000 ;
	    RECT 1124.7001 672.7500 1126.5000 672.9000 ;
	    RECT 1110.3000 671.2500 1126.5000 672.7500 ;
	    RECT 1110.3000 671.1000 1112.1000 671.2500 ;
	    RECT 1124.7001 671.1000 1126.5000 671.2500 ;
	    RECT 1247.1000 672.7500 1248.9000 672.9000 ;
	    RECT 1273.5000 672.7500 1275.3000 672.9000 ;
	    RECT 1247.1000 671.2500 1275.3000 672.7500 ;
	    RECT 1247.1000 671.1000 1248.9000 671.2500 ;
	    RECT 1273.5000 671.1000 1275.3000 671.2500 ;
	    RECT 1405.5000 672.7500 1407.3000 672.9000 ;
	    RECT 1446.3000 672.7500 1448.1000 672.9000 ;
	    RECT 1482.3000 672.7500 1484.1000 672.9000 ;
	    RECT 1405.5000 671.2500 1484.1000 672.7500 ;
	    RECT 1405.5000 671.1000 1407.3000 671.2500 ;
	    RECT 1446.3000 671.1000 1448.1000 671.2500 ;
	    RECT 1482.3000 671.1000 1484.1000 671.2500 ;
	    RECT 231.9000 666.7500 233.7000 666.9000 ;
	    RECT 313.5000 666.7500 315.3000 666.9000 ;
	    RECT 231.9000 665.2500 315.3000 666.7500 ;
	    RECT 231.9000 665.1000 233.7000 665.2500 ;
	    RECT 313.5000 665.1000 315.3000 665.2500 ;
	    RECT 591.9000 666.7500 593.7000 666.9000 ;
	    RECT 613.5000 666.7500 615.3000 666.9000 ;
	    RECT 591.9000 665.2500 615.3000 666.7500 ;
	    RECT 591.9000 665.1000 593.7000 665.2500 ;
	    RECT 613.5000 665.1000 615.3000 665.2500 ;
	    RECT 702.3000 666.7500 704.1000 666.9000 ;
	    RECT 716.7000 666.7500 718.5000 666.9000 ;
	    RECT 702.3000 665.2500 718.5000 666.7500 ;
	    RECT 702.3000 665.1000 704.1000 665.2500 ;
	    RECT 716.7000 665.1000 718.5000 665.2500 ;
	    RECT 764.7000 666.7500 766.5000 666.9000 ;
	    RECT 815.1000 666.7500 816.9000 666.9000 ;
	    RECT 839.1000 666.7500 840.9000 666.9000 ;
	    RECT 853.5000 666.7500 855.3000 666.9000 ;
	    RECT 764.7000 665.2500 855.3000 666.7500 ;
	    RECT 764.7000 665.1000 766.5000 665.2500 ;
	    RECT 815.1000 665.1000 816.9000 665.2500 ;
	    RECT 839.1000 665.1000 840.9000 665.2500 ;
	    RECT 853.5000 665.1000 855.3000 665.2500 ;
	    RECT 884.7000 666.7500 886.5000 666.9000 ;
	    RECT 913.5000 666.7500 915.3000 666.9000 ;
	    RECT 1035.9000 666.7500 1037.7001 666.9000 ;
	    RECT 884.7000 665.2500 1037.7001 666.7500 ;
	    RECT 884.7000 665.1000 886.5000 665.2500 ;
	    RECT 913.5000 665.1000 915.3000 665.2500 ;
	    RECT 1035.9000 665.1000 1037.7001 665.2500 ;
	    RECT 1326.3000 666.7500 1328.1000 666.9000 ;
	    RECT 1331.1000 666.7500 1332.9000 666.9000 ;
	    RECT 1326.3000 665.2500 1332.9000 666.7500 ;
	    RECT 1326.3000 665.1000 1328.1000 665.2500 ;
	    RECT 1331.1000 665.1000 1332.9000 665.2500 ;
	    RECT 1424.7001 666.7500 1426.5000 666.9000 ;
	    RECT 1431.9000 666.7500 1433.7001 666.9000 ;
	    RECT 1424.7001 665.2500 1433.7001 666.7500 ;
	    RECT 1424.7001 665.1000 1426.5000 665.2500 ;
	    RECT 1431.9000 665.1000 1433.7001 665.2500 ;
	    RECT 212.7000 660.7500 214.5000 660.9000 ;
	    RECT 217.5000 660.7500 219.3000 660.9000 ;
	    RECT 212.7000 659.2500 219.3000 660.7500 ;
	    RECT 212.7000 659.1000 214.5000 659.2500 ;
	    RECT 217.5000 659.1000 219.3000 659.2500 ;
	    RECT 222.3000 660.7500 224.1000 660.9000 ;
	    RECT 236.7000 660.7500 238.5000 660.9000 ;
	    RECT 222.3000 659.2500 238.5000 660.7500 ;
	    RECT 222.3000 659.1000 224.1000 659.2500 ;
	    RECT 236.7000 659.1000 238.5000 659.2500 ;
	    RECT 246.3000 660.7500 248.1000 660.9000 ;
	    RECT 255.9000 660.7500 257.7000 660.9000 ;
	    RECT 246.3000 659.2500 257.7000 660.7500 ;
	    RECT 246.3000 659.1000 248.1000 659.2500 ;
	    RECT 255.9000 659.1000 257.7000 659.2500 ;
	    RECT 260.7000 660.7500 262.5000 660.9000 ;
	    RECT 308.7000 660.7500 310.5000 660.9000 ;
	    RECT 260.7000 659.2500 310.5000 660.7500 ;
	    RECT 260.7000 659.1000 262.5000 659.2500 ;
	    RECT 308.7000 659.1000 310.5000 659.2500 ;
	    RECT 515.1000 660.7500 516.9000 660.9000 ;
	    RECT 522.3000 660.7500 524.1000 660.9000 ;
	    RECT 515.1000 659.2500 524.1000 660.7500 ;
	    RECT 515.1000 659.1000 516.9000 659.2500 ;
	    RECT 522.3000 659.1000 524.1000 659.2500 ;
	    RECT 613.5000 660.7500 615.3000 660.9000 ;
	    RECT 630.3000 660.7500 632.1000 660.9000 ;
	    RECT 613.5000 659.2500 632.1000 660.7500 ;
	    RECT 613.5000 659.1000 615.3000 659.2500 ;
	    RECT 630.3000 659.1000 632.1000 659.2500 ;
	    RECT 716.7000 660.7500 718.5000 660.9000 ;
	    RECT 747.9000 660.7500 749.7000 660.9000 ;
	    RECT 716.7000 659.2500 749.7000 660.7500 ;
	    RECT 716.7000 659.1000 718.5000 659.2500 ;
	    RECT 747.9000 659.1000 749.7000 659.2500 ;
	    RECT 853.5000 660.7500 855.3000 660.9000 ;
	    RECT 947.1000 660.7500 948.9000 660.9000 ;
	    RECT 853.5000 659.2500 948.9000 660.7500 ;
	    RECT 853.5000 659.1000 855.3000 659.2500 ;
	    RECT 947.1000 659.1000 948.9000 659.2500 ;
	    RECT 973.5000 660.7500 975.3000 660.9000 ;
	    RECT 1119.9000 660.7500 1121.7001 660.9000 ;
	    RECT 973.5000 659.2500 1121.7001 660.7500 ;
	    RECT 973.5000 659.1000 975.3000 659.2500 ;
	    RECT 1119.9000 659.1000 1121.7001 659.2500 ;
	    RECT 1244.7001 660.7500 1246.5000 660.9000 ;
	    RECT 1266.3000 660.7500 1268.1000 660.9000 ;
	    RECT 1244.7001 659.2500 1268.1000 660.7500 ;
	    RECT 1244.7001 659.1000 1246.5000 659.2500 ;
	    RECT 1266.3000 659.1000 1268.1000 659.2500 ;
	    RECT 42.3000 654.7500 44.1000 654.9000 ;
	    RECT 66.3000 654.7500 68.1000 654.9000 ;
	    RECT 42.3000 653.2500 68.1000 654.7500 ;
	    RECT 42.3000 653.1000 44.1000 653.2500 ;
	    RECT 66.3000 653.1000 68.1000 653.2500 ;
	    RECT 167.1000 654.7500 168.9000 654.9000 ;
	    RECT 198.3000 654.7500 200.1000 654.9000 ;
	    RECT 167.1000 653.2500 200.1000 654.7500 ;
	    RECT 167.1000 653.1000 168.9000 653.2500 ;
	    RECT 198.3000 653.1000 200.1000 653.2500 ;
	    RECT 239.1000 654.7500 240.9000 654.9000 ;
	    RECT 255.9000 654.7500 257.7000 654.9000 ;
	    RECT 284.7000 654.7500 286.5000 654.9000 ;
	    RECT 239.1000 653.2500 286.5000 654.7500 ;
	    RECT 239.1000 653.1000 240.9000 653.2500 ;
	    RECT 255.9000 653.1000 257.7000 653.2500 ;
	    RECT 284.7000 653.1000 286.5000 653.2500 ;
	    RECT 301.5000 654.7500 303.3000 654.9000 ;
	    RECT 551.1000 654.7500 552.9000 654.9000 ;
	    RECT 582.3000 654.7500 584.1000 654.9000 ;
	    RECT 301.5000 653.2500 584.1000 654.7500 ;
	    RECT 301.5000 653.1000 303.3000 653.2500 ;
	    RECT 551.1000 653.1000 552.9000 653.2500 ;
	    RECT 582.3000 653.1000 584.1000 653.2500 ;
	    RECT 587.1000 654.7500 588.9000 654.9000 ;
	    RECT 596.7000 654.7500 598.5000 654.9000 ;
	    RECT 587.1000 653.2500 598.5000 654.7500 ;
	    RECT 587.1000 653.1000 588.9000 653.2500 ;
	    RECT 596.7000 653.1000 598.5000 653.2500 ;
	    RECT 611.1000 654.7500 612.9000 654.9000 ;
	    RECT 651.9000 654.7500 653.7000 654.9000 ;
	    RECT 611.1000 653.2500 653.7000 654.7500 ;
	    RECT 611.1000 653.1000 612.9000 653.2500 ;
	    RECT 651.9000 653.1000 653.7000 653.2500 ;
	    RECT 697.5000 654.7500 699.3000 654.9000 ;
	    RECT 707.1000 654.7500 708.9000 654.9000 ;
	    RECT 716.7000 654.7500 718.5000 654.9000 ;
	    RECT 697.5000 653.2500 718.5000 654.7500 ;
	    RECT 697.5000 653.1000 699.3000 653.2500 ;
	    RECT 707.1000 653.1000 708.9000 653.2500 ;
	    RECT 716.7000 653.1000 718.5000 653.2500 ;
	    RECT 721.5000 654.7500 723.3000 654.9000 ;
	    RECT 757.5000 654.7500 759.3000 654.9000 ;
	    RECT 721.5000 653.2500 759.3000 654.7500 ;
	    RECT 721.5000 653.1000 723.3000 653.2500 ;
	    RECT 757.5000 653.1000 759.3000 653.2500 ;
	    RECT 764.7000 654.7500 766.5000 654.9000 ;
	    RECT 819.9000 654.7500 821.7000 654.9000 ;
	    RECT 867.9000 654.7500 869.7000 654.9000 ;
	    RECT 764.7000 653.2500 869.7000 654.7500 ;
	    RECT 764.7000 653.1000 766.5000 653.2500 ;
	    RECT 819.9000 653.1000 821.7000 653.2500 ;
	    RECT 867.9000 653.1000 869.7000 653.2500 ;
	    RECT 978.3000 654.7500 980.1000 654.9000 ;
	    RECT 1019.1000 654.7500 1020.9000 654.9000 ;
	    RECT 978.3000 653.2500 1020.9000 654.7500 ;
	    RECT 978.3000 653.1000 980.1000 653.2500 ;
	    RECT 1019.1000 653.1000 1020.9000 653.2500 ;
	    RECT 275.1000 648.7500 276.9000 648.9000 ;
	    RECT 289.5000 648.7500 291.3000 648.9000 ;
	    RECT 275.1000 647.2500 291.3000 648.7500 ;
	    RECT 275.1000 647.1000 276.9000 647.2500 ;
	    RECT 289.5000 647.1000 291.3000 647.2500 ;
	    RECT 323.1000 648.7500 324.9000 648.9000 ;
	    RECT 344.7000 648.7500 346.5000 648.9000 ;
	    RECT 323.1000 647.2500 346.5000 648.7500 ;
	    RECT 323.1000 647.1000 324.9000 647.2500 ;
	    RECT 344.7000 647.1000 346.5000 647.2500 ;
	    RECT 359.1000 648.7500 360.9000 648.9000 ;
	    RECT 435.9000 648.7500 437.7000 648.9000 ;
	    RECT 359.1000 647.2500 437.7000 648.7500 ;
	    RECT 359.1000 647.1000 360.9000 647.2500 ;
	    RECT 435.9000 647.1000 437.7000 647.2500 ;
	    RECT 577.5000 648.7500 579.3000 648.9000 ;
	    RECT 642.3000 648.7500 644.1000 648.9000 ;
	    RECT 577.5000 647.2500 644.1000 648.7500 ;
	    RECT 577.5000 647.1000 579.3000 647.2500 ;
	    RECT 642.3000 647.1000 644.1000 647.2500 ;
	    RECT 656.7000 648.7500 658.5000 648.9000 ;
	    RECT 714.3000 648.7500 716.1000 648.9000 ;
	    RECT 656.7000 647.2500 716.1000 648.7500 ;
	    RECT 656.7000 647.1000 658.5000 647.2500 ;
	    RECT 714.3000 647.1000 716.1000 647.2500 ;
	    RECT 747.9000 648.7500 749.7000 648.9000 ;
	    RECT 841.5000 648.7500 843.3000 648.9000 ;
	    RECT 872.7000 648.7500 874.5000 648.9000 ;
	    RECT 747.9000 647.2500 874.5000 648.7500 ;
	    RECT 747.9000 647.1000 749.7000 647.2500 ;
	    RECT 841.5000 647.1000 843.3000 647.2500 ;
	    RECT 872.7000 647.1000 874.5000 647.2500 ;
	    RECT 1175.1000 648.7500 1176.9000 648.9000 ;
	    RECT 1220.7001 648.7500 1222.5000 648.9000 ;
	    RECT 1175.1000 647.2500 1222.5000 648.7500 ;
	    RECT 1175.1000 647.1000 1176.9000 647.2500 ;
	    RECT 1220.7001 647.1000 1222.5000 647.2500 ;
	    RECT 1391.1000 648.7500 1392.9000 648.9000 ;
	    RECT 1400.7001 648.7500 1402.5000 648.9000 ;
	    RECT 1391.1000 647.2500 1402.5000 648.7500 ;
	    RECT 1391.1000 647.1000 1392.9000 647.2500 ;
	    RECT 1400.7001 647.1000 1402.5000 647.2500 ;
	    RECT 1463.1000 648.7500 1464.9000 648.9000 ;
	    RECT 1484.7001 648.7500 1486.5000 648.9000 ;
	    RECT 1463.1000 647.2500 1486.5000 648.7500 ;
	    RECT 1463.1000 647.1000 1464.9000 647.2500 ;
	    RECT 1484.7001 647.1000 1486.5000 647.2500 ;
	    RECT 1491.9000 648.7500 1493.7001 648.9000 ;
	    RECT 1503.9000 648.7500 1505.7001 648.9000 ;
	    RECT 1491.9000 647.2500 1505.7001 648.7500 ;
	    RECT 1491.9000 647.1000 1493.7001 647.2500 ;
	    RECT 1503.9000 647.1000 1505.7001 647.2500 ;
	    RECT 39.9000 642.7500 41.7000 642.9000 ;
	    RECT 78.3000 642.7500 80.1000 642.9000 ;
	    RECT 102.3000 642.7500 104.1000 642.9000 ;
	    RECT 119.1000 642.7500 120.9000 642.9000 ;
	    RECT 248.7000 642.7500 250.5000 642.9000 ;
	    RECT 296.7000 642.7500 298.5000 642.9000 ;
	    RECT 39.9000 641.2500 298.5000 642.7500 ;
	    RECT 39.9000 641.1000 41.7000 641.2500 ;
	    RECT 78.3000 641.1000 80.1000 641.2500 ;
	    RECT 102.3000 641.1000 104.1000 641.2500 ;
	    RECT 119.1000 641.1000 120.9000 641.2500 ;
	    RECT 248.7000 641.1000 250.5000 641.2500 ;
	    RECT 296.7000 641.1000 298.5000 641.2500 ;
	    RECT 308.7000 642.7500 310.5000 642.9000 ;
	    RECT 337.5000 642.7500 339.3000 642.9000 ;
	    RECT 308.7000 641.2500 339.3000 642.7500 ;
	    RECT 308.7000 641.1000 310.5000 641.2500 ;
	    RECT 337.5000 641.1000 339.3000 641.2500 ;
	    RECT 431.1000 642.7500 432.9000 642.9000 ;
	    RECT 517.5000 642.7500 519.3000 642.9000 ;
	    RECT 431.1000 641.2500 519.3000 642.7500 ;
	    RECT 431.1000 641.1000 432.9000 641.2500 ;
	    RECT 517.5000 641.1000 519.3000 641.2500 ;
	    RECT 582.3000 642.7500 584.1000 642.9000 ;
	    RECT 654.3000 642.7500 656.1000 642.9000 ;
	    RECT 582.3000 641.2500 656.1000 642.7500 ;
	    RECT 582.3000 641.1000 584.1000 641.2500 ;
	    RECT 654.3000 641.1000 656.1000 641.2500 ;
	    RECT 659.1000 642.7500 660.9000 642.9000 ;
	    RECT 690.3000 642.7500 692.1000 642.9000 ;
	    RECT 659.1000 641.2500 692.1000 642.7500 ;
	    RECT 659.1000 641.1000 660.9000 641.2500 ;
	    RECT 690.3000 641.1000 692.1000 641.2500 ;
	    RECT 695.1000 642.7500 696.9000 642.9000 ;
	    RECT 699.9000 642.7500 701.7000 642.9000 ;
	    RECT 695.1000 641.2500 701.7000 642.7500 ;
	    RECT 695.1000 641.1000 696.9000 641.2500 ;
	    RECT 699.9000 641.1000 701.7000 641.2500 ;
	    RECT 704.7000 642.7500 706.5000 642.9000 ;
	    RECT 721.5000 642.7500 723.3000 642.9000 ;
	    RECT 704.7000 641.2500 723.3000 642.7500 ;
	    RECT 704.7000 641.1000 706.5000 641.2500 ;
	    RECT 721.5000 641.1000 723.3000 641.2500 ;
	    RECT 735.9000 642.7500 737.7000 642.9000 ;
	    RECT 779.1000 642.7500 780.9000 642.9000 ;
	    RECT 735.9000 641.2500 780.9000 642.7500 ;
	    RECT 735.9000 641.1000 737.7000 641.2500 ;
	    RECT 779.1000 641.1000 780.9000 641.2500 ;
	    RECT 783.9000 642.7500 785.7000 642.9000 ;
	    RECT 815.1000 642.7500 816.9000 642.9000 ;
	    RECT 1177.5000 642.7500 1179.3000 642.9000 ;
	    RECT 783.9000 641.2500 1179.3000 642.7500 ;
	    RECT 783.9000 641.1000 785.7000 641.2500 ;
	    RECT 815.1000 641.1000 816.9000 641.2500 ;
	    RECT 1177.5000 641.1000 1179.3000 641.2500 ;
	    RECT 1189.5000 642.7500 1191.3000 642.9000 ;
	    RECT 1271.1000 642.7500 1272.9000 642.9000 ;
	    RECT 1189.5000 641.2500 1272.9000 642.7500 ;
	    RECT 1189.5000 641.1000 1191.3000 641.2500 ;
	    RECT 1271.1000 641.1000 1272.9000 641.2500 ;
	    RECT 1275.9000 642.7500 1277.7001 642.9000 ;
	    RECT 1295.1000 642.7500 1296.9000 642.9000 ;
	    RECT 1302.3000 642.7500 1304.1000 642.9000 ;
	    RECT 1275.9000 641.2500 1304.1000 642.7500 ;
	    RECT 1275.9000 641.1000 1277.7001 641.2500 ;
	    RECT 1295.1000 641.1000 1296.9000 641.2500 ;
	    RECT 1302.3000 641.1000 1304.1000 641.2500 ;
	    RECT 1314.3000 642.7500 1316.1000 642.9000 ;
	    RECT 1376.7001 642.7500 1378.5000 642.9000 ;
	    RECT 1314.3000 641.2500 1378.5000 642.7500 ;
	    RECT 1314.3000 641.1000 1316.1000 641.2500 ;
	    RECT 1376.7001 641.1000 1378.5000 641.2500 ;
	    RECT 1398.3000 642.7500 1400.1000 642.9000 ;
	    RECT 1419.9000 642.7500 1421.7001 642.9000 ;
	    RECT 1398.3000 641.2500 1421.7001 642.7500 ;
	    RECT 1398.3000 641.1000 1400.1000 641.2500 ;
	    RECT 1419.9000 641.1000 1421.7001 641.2500 ;
	    RECT 1460.7001 642.7500 1462.5000 642.9000 ;
	    RECT 1482.3000 642.7500 1484.1000 642.9000 ;
	    RECT 1460.7001 641.2500 1484.1000 642.7500 ;
	    RECT 1460.7001 641.1000 1462.5000 641.2500 ;
	    RECT 1482.3000 641.1000 1484.1000 641.2500 ;
	    RECT 71.1000 636.7500 72.9000 636.9000 ;
	    RECT 145.5000 636.7500 147.3000 636.9000 ;
	    RECT 71.1000 635.2500 147.3000 636.7500 ;
	    RECT 71.1000 635.1000 72.9000 635.2500 ;
	    RECT 145.5000 635.1000 147.3000 635.2500 ;
	    RECT 159.9000 636.7500 161.7000 636.9000 ;
	    RECT 169.5000 636.7500 171.3000 636.9000 ;
	    RECT 159.9000 635.2500 171.3000 636.7500 ;
	    RECT 159.9000 635.1000 161.7000 635.2500 ;
	    RECT 169.5000 635.1000 171.3000 635.2500 ;
	    RECT 217.5000 636.7500 219.3000 636.9000 ;
	    RECT 239.1000 636.7500 240.9000 636.9000 ;
	    RECT 217.5000 635.2500 240.9000 636.7500 ;
	    RECT 217.5000 635.1000 219.3000 635.2500 ;
	    RECT 239.1000 635.1000 240.9000 635.2500 ;
	    RECT 627.9000 636.7500 629.7000 636.9000 ;
	    RECT 671.1000 636.7500 672.9000 636.9000 ;
	    RECT 627.9000 635.2500 672.9000 636.7500 ;
	    RECT 627.9000 635.1000 629.7000 635.2500 ;
	    RECT 671.1000 635.1000 672.9000 635.2500 ;
	    RECT 750.3000 636.7500 752.1000 636.9000 ;
	    RECT 781.5000 636.7500 783.3000 636.9000 ;
	    RECT 750.3000 635.2500 783.3000 636.7500 ;
	    RECT 750.3000 635.1000 752.1000 635.2500 ;
	    RECT 781.5000 635.1000 783.3000 635.2500 ;
	    RECT 848.7000 636.7500 850.5000 636.9000 ;
	    RECT 973.5000 636.7500 975.3000 636.9000 ;
	    RECT 848.7000 635.2500 975.3000 636.7500 ;
	    RECT 848.7000 635.1000 850.5000 635.2500 ;
	    RECT 973.5000 635.1000 975.3000 635.2500 ;
	    RECT 1237.5000 636.7500 1239.3000 636.9000 ;
	    RECT 1249.5000 636.7500 1251.3000 636.9000 ;
	    RECT 1237.5000 635.2500 1251.3000 636.7500 ;
	    RECT 1237.5000 635.1000 1239.3000 635.2500 ;
	    RECT 1249.5000 635.1000 1251.3000 635.2500 ;
	    RECT 1350.3000 636.7500 1352.1000 636.9000 ;
	    RECT 1403.1000 636.7500 1404.9000 636.9000 ;
	    RECT 1350.3000 635.2500 1404.9000 636.7500 ;
	    RECT 1350.3000 635.1000 1352.1000 635.2500 ;
	    RECT 1403.1000 635.1000 1404.9000 635.2500 ;
	    RECT 1419.9000 636.7500 1421.7001 636.9000 ;
	    RECT 1441.5000 636.7500 1443.3000 636.9000 ;
	    RECT 1477.5000 636.7500 1479.3000 636.9000 ;
	    RECT 1419.9000 635.2500 1479.3000 636.7500 ;
	    RECT 1419.9000 635.1000 1421.7001 635.2500 ;
	    RECT 1441.5000 635.1000 1443.3000 635.2500 ;
	    RECT 1477.5000 635.1000 1479.3000 635.2500 ;
	    RECT 1494.3000 636.7500 1496.1000 636.9000 ;
	    RECT 1520.7001 636.7500 1522.5000 636.9000 ;
	    RECT 1494.3000 635.2500 1522.5000 636.7500 ;
	    RECT 1494.3000 635.1000 1496.1000 635.2500 ;
	    RECT 1520.7001 635.1000 1522.5000 635.2500 ;
	    RECT 234.3000 630.7500 236.1000 630.9000 ;
	    RECT 239.1000 630.7500 240.9000 630.9000 ;
	    RECT 234.3000 629.2500 240.9000 630.7500 ;
	    RECT 234.3000 629.1000 236.1000 629.2500 ;
	    RECT 239.1000 629.1000 240.9000 629.2500 ;
	    RECT 270.3000 630.7500 272.1000 630.9000 ;
	    RECT 320.7000 630.7500 322.5000 630.9000 ;
	    RECT 270.3000 629.2500 322.5000 630.7500 ;
	    RECT 270.3000 629.1000 272.1000 629.2500 ;
	    RECT 320.7000 629.1000 322.5000 629.2500 ;
	    RECT 330.3000 630.7500 332.1000 630.9000 ;
	    RECT 399.9000 630.7500 401.7000 630.9000 ;
	    RECT 330.3000 629.2500 401.7000 630.7500 ;
	    RECT 330.3000 629.1000 332.1000 629.2500 ;
	    RECT 399.9000 629.1000 401.7000 629.2500 ;
	    RECT 721.5000 630.7500 723.3000 630.9000 ;
	    RECT 865.5000 630.7500 867.3000 630.9000 ;
	    RECT 721.5000 629.2500 867.3000 630.7500 ;
	    RECT 721.5000 629.1000 723.3000 629.2500 ;
	    RECT 865.5000 629.1000 867.3000 629.2500 ;
	    RECT 939.9000 630.7500 941.7000 630.9000 ;
	    RECT 980.7000 630.7500 982.5000 630.9000 ;
	    RECT 939.9000 629.2500 982.5000 630.7500 ;
	    RECT 939.9000 629.1000 941.7000 629.2500 ;
	    RECT 980.7000 629.1000 982.5000 629.2500 ;
	    RECT 999.9000 630.7500 1001.7000 630.9000 ;
	    RECT 1055.1000 630.7500 1056.9000 630.9000 ;
	    RECT 999.9000 629.2500 1056.9000 630.7500 ;
	    RECT 999.9000 629.1000 1001.7000 629.2500 ;
	    RECT 1055.1000 629.1000 1056.9000 629.2500 ;
	    RECT 1064.7001 630.7500 1066.5000 630.9000 ;
	    RECT 1117.5000 630.7500 1119.3000 630.9000 ;
	    RECT 1064.7001 629.2500 1119.3000 630.7500 ;
	    RECT 1064.7001 629.1000 1066.5000 629.2500 ;
	    RECT 1117.5000 629.1000 1119.3000 629.2500 ;
	    RECT 1223.1000 630.7500 1224.9000 630.9000 ;
	    RECT 1285.5000 630.7500 1287.3000 630.9000 ;
	    RECT 1223.1000 629.2500 1287.3000 630.7500 ;
	    RECT 1223.1000 629.1000 1224.9000 629.2500 ;
	    RECT 1285.5000 629.1000 1287.3000 629.2500 ;
	    RECT 1338.3000 630.7500 1340.1000 630.9000 ;
	    RECT 1345.5000 630.7500 1347.3000 630.9000 ;
	    RECT 1338.3000 629.2500 1347.3000 630.7500 ;
	    RECT 1338.3000 629.1000 1340.1000 629.2500 ;
	    RECT 1345.5000 629.1000 1347.3000 629.2500 ;
	    RECT 1386.3000 630.7500 1388.1000 630.9000 ;
	    RECT 1429.5000 630.7500 1431.3000 630.9000 ;
	    RECT 1386.3000 629.2500 1431.3000 630.7500 ;
	    RECT 1386.3000 629.1000 1388.1000 629.2500 ;
	    RECT 1429.5000 629.1000 1431.3000 629.2500 ;
	    RECT 1487.1000 630.7500 1488.9000 630.9000 ;
	    RECT 1530.3000 630.7500 1532.1000 630.9000 ;
	    RECT 1487.1000 629.2500 1532.1000 630.7500 ;
	    RECT 1487.1000 629.1000 1488.9000 629.2500 ;
	    RECT 1530.3000 629.1000 1532.1000 629.2500 ;
	    RECT 491.1000 624.7500 492.9000 624.9000 ;
	    RECT 546.3000 624.7500 548.1000 624.9000 ;
	    RECT 491.1000 623.2500 548.1000 624.7500 ;
	    RECT 491.1000 623.1000 492.9000 623.2500 ;
	    RECT 546.3000 623.1000 548.1000 623.2500 ;
	    RECT 591.9000 624.7500 593.7000 624.9000 ;
	    RECT 642.3000 624.7500 644.1000 624.9000 ;
	    RECT 591.9000 623.2500 644.1000 624.7500 ;
	    RECT 591.9000 623.1000 593.7000 623.2500 ;
	    RECT 642.3000 623.1000 644.1000 623.2500 ;
	    RECT 723.9000 624.7500 725.7000 624.9000 ;
	    RECT 752.7000 624.7500 754.5000 624.9000 ;
	    RECT 723.9000 623.2500 754.5000 624.7500 ;
	    RECT 723.9000 623.1000 725.7000 623.2500 ;
	    RECT 752.7000 623.1000 754.5000 623.2500 ;
	    RECT 776.7000 624.7500 778.5000 624.9000 ;
	    RECT 851.1000 624.7500 852.9000 624.9000 ;
	    RECT 776.7000 623.2500 852.9000 624.7500 ;
	    RECT 776.7000 623.1000 778.5000 623.2500 ;
	    RECT 851.1000 623.1000 852.9000 623.2500 ;
	    RECT 863.1000 624.7500 864.9000 624.9000 ;
	    RECT 906.3000 624.7500 908.1000 624.9000 ;
	    RECT 911.1000 624.7500 912.9000 624.9000 ;
	    RECT 863.1000 623.2500 912.9000 624.7500 ;
	    RECT 863.1000 623.1000 864.9000 623.2500 ;
	    RECT 906.3000 623.1000 908.1000 623.2500 ;
	    RECT 911.1000 623.1000 912.9000 623.2500 ;
	    RECT 1081.5000 624.7500 1083.3000 624.9000 ;
	    RECT 1107.9000 624.7500 1109.7001 624.9000 ;
	    RECT 1081.5000 623.2500 1109.7001 624.7500 ;
	    RECT 1081.5000 623.1000 1083.3000 623.2500 ;
	    RECT 1107.9000 623.1000 1109.7001 623.2500 ;
	    RECT 1230.3000 624.7500 1232.1000 624.9000 ;
	    RECT 1278.3000 624.7500 1280.1000 624.9000 ;
	    RECT 1230.3000 623.2500 1280.1000 624.7500 ;
	    RECT 1230.3000 623.1000 1232.1000 623.2500 ;
	    RECT 1278.3000 623.1000 1280.1000 623.2500 ;
	    RECT 1304.7001 624.7500 1306.5000 624.9000 ;
	    RECT 1340.7001 624.7500 1342.5000 624.9000 ;
	    RECT 1304.7001 623.2500 1342.5000 624.7500 ;
	    RECT 1304.7001 623.1000 1306.5000 623.2500 ;
	    RECT 1340.7001 623.1000 1342.5000 623.2500 ;
	    RECT 1436.7001 624.7500 1438.5000 624.9000 ;
	    RECT 1479.9000 624.7500 1481.7001 624.9000 ;
	    RECT 1436.7001 623.2500 1481.7001 624.7500 ;
	    RECT 1436.7001 623.1000 1438.5000 623.2500 ;
	    RECT 1479.9000 623.1000 1481.7001 623.2500 ;
	    RECT 1523.1000 624.7500 1524.9000 624.9000 ;
	    RECT 1547.1000 624.7500 1548.9000 624.9000 ;
	    RECT 1523.1000 623.2500 1548.9000 624.7500 ;
	    RECT 1523.1000 623.1000 1524.9000 623.2500 ;
	    RECT 1547.1000 623.1000 1548.9000 623.2500 ;
	    RECT 313.5000 618.7500 315.3000 618.9000 ;
	    RECT 342.3000 618.7500 344.1000 618.9000 ;
	    RECT 313.5000 617.2500 344.1000 618.7500 ;
	    RECT 313.5000 617.1000 315.3000 617.2500 ;
	    RECT 342.3000 617.1000 344.1000 617.2500 ;
	    RECT 387.9000 618.7500 389.7000 618.9000 ;
	    RECT 416.7000 618.7500 418.5000 618.9000 ;
	    RECT 387.9000 617.2500 418.5000 618.7500 ;
	    RECT 387.9000 617.1000 389.7000 617.2500 ;
	    RECT 416.7000 617.1000 418.5000 617.2500 ;
	    RECT 445.5000 618.7500 447.3000 618.9000 ;
	    RECT 464.7000 618.7500 466.5000 618.9000 ;
	    RECT 445.5000 617.2500 466.5000 618.7500 ;
	    RECT 445.5000 617.1000 447.3000 617.2500 ;
	    RECT 464.7000 617.1000 466.5000 617.2500 ;
	    RECT 647.1000 618.7500 648.9000 618.9000 ;
	    RECT 661.5000 618.7500 663.3000 618.9000 ;
	    RECT 687.9000 618.7500 689.7000 618.9000 ;
	    RECT 647.1000 617.2500 689.7000 618.7500 ;
	    RECT 647.1000 617.1000 648.9000 617.2500 ;
	    RECT 661.5000 617.1000 663.3000 617.2500 ;
	    RECT 687.9000 617.1000 689.7000 617.2500 ;
	    RECT 882.3000 618.7500 884.1000 618.9000 ;
	    RECT 896.7000 618.7500 898.5000 618.9000 ;
	    RECT 882.3000 617.2500 898.5000 618.7500 ;
	    RECT 882.3000 617.1000 884.1000 617.2500 ;
	    RECT 896.7000 617.1000 898.5000 617.2500 ;
	    RECT 1059.9000 618.7500 1061.7001 618.9000 ;
	    RECT 1117.5000 618.7500 1119.3000 618.9000 ;
	    RECT 1059.9000 617.2500 1119.3000 618.7500 ;
	    RECT 1059.9000 617.1000 1061.7001 617.2500 ;
	    RECT 1117.5000 617.1000 1119.3000 617.2500 ;
	    RECT 1177.5000 618.7500 1179.3000 618.9000 ;
	    RECT 1206.3000 618.7500 1208.1000 618.9000 ;
	    RECT 1213.5000 618.7500 1215.3000 618.9000 ;
	    RECT 1177.5000 617.2500 1215.3000 618.7500 ;
	    RECT 1177.5000 617.1000 1179.3000 617.2500 ;
	    RECT 1206.3000 617.1000 1208.1000 617.2500 ;
	    RECT 1213.5000 617.1000 1215.3000 617.2500 ;
	    RECT 1340.7001 618.7500 1342.5000 618.9000 ;
	    RECT 1347.9000 618.7500 1349.7001 618.9000 ;
	    RECT 1340.7001 617.2500 1349.7001 618.7500 ;
	    RECT 1340.7001 617.1000 1342.5000 617.2500 ;
	    RECT 1347.9000 617.1000 1349.7001 617.2500 ;
	    RECT 1367.1000 618.7500 1368.9000 618.9000 ;
	    RECT 1381.5000 618.7500 1383.3000 618.9000 ;
	    RECT 1367.1000 617.2500 1383.3000 618.7500 ;
	    RECT 1367.1000 617.1000 1368.9000 617.2500 ;
	    RECT 1381.5000 617.1000 1383.3000 617.2500 ;
	    RECT 1407.9000 618.7500 1409.7001 618.9000 ;
	    RECT 1415.1000 618.7500 1416.9000 618.9000 ;
	    RECT 1407.9000 617.2500 1416.9000 618.7500 ;
	    RECT 1407.9000 617.1000 1409.7001 617.2500 ;
	    RECT 1415.1000 617.1000 1416.9000 617.2500 ;
	    RECT 1429.5000 618.7500 1431.3000 618.9000 ;
	    RECT 1475.1000 618.7500 1476.9000 618.9000 ;
	    RECT 1429.5000 617.2500 1476.9000 618.7500 ;
	    RECT 1429.5000 617.1000 1431.3000 617.2500 ;
	    RECT 1475.1000 617.1000 1476.9000 617.2500 ;
	    RECT 1482.3000 618.7500 1484.1000 618.9000 ;
	    RECT 1508.7001 618.7500 1510.5000 618.9000 ;
	    RECT 1482.3000 617.2500 1510.5000 618.7500 ;
	    RECT 1482.3000 617.1000 1484.1000 617.2500 ;
	    RECT 1508.7001 617.1000 1510.5000 617.2500 ;
	    RECT 1530.3000 618.7500 1532.1000 618.9000 ;
	    RECT 1544.7001 618.7500 1546.5000 618.9000 ;
	    RECT 1530.3000 617.2500 1546.5000 618.7500 ;
	    RECT 1530.3000 617.1000 1532.1000 617.2500 ;
	    RECT 1544.7001 617.1000 1546.5000 617.2500 ;
	    RECT 111.9000 612.7500 113.7000 612.9000 ;
	    RECT 174.3000 612.7500 176.1000 612.9000 ;
	    RECT 215.1000 612.7500 216.9000 612.9000 ;
	    RECT 111.9000 611.2500 216.9000 612.7500 ;
	    RECT 111.9000 611.1000 113.7000 611.2500 ;
	    RECT 174.3000 611.1000 176.1000 611.2500 ;
	    RECT 215.1000 611.1000 216.9000 611.2500 ;
	    RECT 253.5000 612.7500 255.3000 612.9000 ;
	    RECT 260.7000 612.7500 262.5000 612.9000 ;
	    RECT 253.5000 611.2500 262.5000 612.7500 ;
	    RECT 253.5000 611.1000 255.3000 611.2500 ;
	    RECT 260.7000 611.1000 262.5000 611.2500 ;
	    RECT 356.7000 612.7500 358.5000 612.9000 ;
	    RECT 385.5000 612.7500 387.3000 612.9000 ;
	    RECT 356.7000 611.2500 387.3000 612.7500 ;
	    RECT 356.7000 611.1000 358.5000 611.2500 ;
	    RECT 385.5000 611.1000 387.3000 611.2500 ;
	    RECT 618.3000 612.7500 620.1000 612.9000 ;
	    RECT 695.1000 612.7500 696.9000 612.9000 ;
	    RECT 618.3000 611.2500 696.9000 612.7500 ;
	    RECT 618.3000 611.1000 620.1000 611.2500 ;
	    RECT 695.1000 611.1000 696.9000 611.2500 ;
	    RECT 745.5000 612.7500 747.3000 612.9000 ;
	    RECT 834.3000 612.7500 836.1000 612.9000 ;
	    RECT 745.5000 611.2500 836.1000 612.7500 ;
	    RECT 745.5000 611.1000 747.3000 611.2500 ;
	    RECT 834.3000 611.1000 836.1000 611.2500 ;
	    RECT 906.3000 612.7500 908.1000 612.9000 ;
	    RECT 935.1000 612.7500 936.9000 612.9000 ;
	    RECT 906.3000 611.2500 936.9000 612.7500 ;
	    RECT 906.3000 611.1000 908.1000 611.2500 ;
	    RECT 935.1000 611.1000 936.9000 611.2500 ;
	    RECT 1107.9000 612.7500 1109.7001 612.9000 ;
	    RECT 1143.9000 612.7500 1145.7001 612.9000 ;
	    RECT 1107.9000 611.2500 1145.7001 612.7500 ;
	    RECT 1107.9000 611.1000 1109.7001 611.2500 ;
	    RECT 1143.9000 611.1000 1145.7001 611.2500 ;
	    RECT 1175.1000 612.7500 1176.9000 612.9000 ;
	    RECT 1208.7001 612.7500 1210.5000 612.9000 ;
	    RECT 1175.1000 611.2500 1210.5000 612.7500 ;
	    RECT 1175.1000 611.1000 1176.9000 611.2500 ;
	    RECT 1208.7001 611.1000 1210.5000 611.2500 ;
	    RECT 1247.1000 612.7500 1248.9000 612.9000 ;
	    RECT 1275.9000 612.7500 1277.7001 612.9000 ;
	    RECT 1247.1000 611.2500 1277.7001 612.7500 ;
	    RECT 1247.1000 611.1000 1248.9000 611.2500 ;
	    RECT 1275.9000 611.1000 1277.7001 611.2500 ;
	    RECT 1343.1000 612.7500 1344.9000 612.9000 ;
	    RECT 1350.3000 612.7500 1352.1000 612.9000 ;
	    RECT 1343.1000 611.2500 1352.1000 612.7500 ;
	    RECT 1343.1000 611.1000 1344.9000 611.2500 ;
	    RECT 1350.3000 611.1000 1352.1000 611.2500 ;
	    RECT 1374.3000 612.7500 1376.1000 612.9000 ;
	    RECT 1381.5000 612.7500 1383.3000 612.9000 ;
	    RECT 1374.3000 611.2500 1383.3000 612.7500 ;
	    RECT 1374.3000 611.1000 1376.1000 611.2500 ;
	    RECT 1381.5000 611.1000 1383.3000 611.2500 ;
	    RECT 1518.3000 612.7500 1520.1000 612.9000 ;
	    RECT 1527.9000 612.7500 1529.7001 612.9000 ;
	    RECT 1542.3000 612.7500 1544.1000 612.9000 ;
	    RECT 1518.3000 611.2500 1544.1000 612.7500 ;
	    RECT 1518.3000 611.1000 1520.1000 611.2500 ;
	    RECT 1527.9000 611.1000 1529.7001 611.2500 ;
	    RECT 1542.3000 611.1000 1544.1000 611.2500 ;
	    RECT 198.3000 606.7500 200.1000 606.9000 ;
	    RECT 219.9000 606.7500 221.7000 606.9000 ;
	    RECT 198.3000 605.2500 221.7000 606.7500 ;
	    RECT 198.3000 605.1000 200.1000 605.2500 ;
	    RECT 219.9000 605.1000 221.7000 605.2500 ;
	    RECT 234.3000 606.7500 236.1000 606.9000 ;
	    RECT 251.1000 606.7500 252.9000 606.9000 ;
	    RECT 234.3000 605.2500 252.9000 606.7500 ;
	    RECT 234.3000 605.1000 236.1000 605.2500 ;
	    RECT 251.1000 605.1000 252.9000 605.2500 ;
	    RECT 303.9000 606.7500 305.7000 606.9000 ;
	    RECT 373.5000 606.7500 375.3000 606.9000 ;
	    RECT 303.9000 605.2500 375.3000 606.7500 ;
	    RECT 303.9000 605.1000 305.7000 605.2500 ;
	    RECT 373.5000 605.1000 375.3000 605.2500 ;
	    RECT 474.3000 606.7500 476.1000 606.9000 ;
	    RECT 575.1000 606.7500 576.9000 606.9000 ;
	    RECT 474.3000 605.2500 576.9000 606.7500 ;
	    RECT 474.3000 605.1000 476.1000 605.2500 ;
	    RECT 575.1000 605.1000 576.9000 605.2500 ;
	    RECT 707.1000 606.7500 708.9000 606.9000 ;
	    RECT 714.3000 606.7500 716.1000 606.9000 ;
	    RECT 771.9000 606.7500 773.7000 606.9000 ;
	    RECT 707.1000 605.2500 773.7000 606.7500 ;
	    RECT 707.1000 605.1000 708.9000 605.2500 ;
	    RECT 714.3000 605.1000 716.1000 605.2500 ;
	    RECT 771.9000 605.1000 773.7000 605.2500 ;
	    RECT 913.5000 606.7500 915.3000 606.9000 ;
	    RECT 1067.1000 606.7500 1068.9000 606.9000 ;
	    RECT 913.5000 605.2500 1068.9000 606.7500 ;
	    RECT 913.5000 605.1000 915.3000 605.2500 ;
	    RECT 1067.1000 605.1000 1068.9000 605.2500 ;
	    RECT 1100.7001 606.7500 1102.5000 606.9000 ;
	    RECT 1146.3000 606.7500 1148.1000 606.9000 ;
	    RECT 1244.7001 606.7500 1246.5000 606.9000 ;
	    RECT 1251.9000 606.7500 1253.7001 606.9000 ;
	    RECT 1100.7001 605.2500 1253.7001 606.7500 ;
	    RECT 1100.7001 605.1000 1102.5000 605.2500 ;
	    RECT 1146.3000 605.1000 1148.1000 605.2500 ;
	    RECT 1244.7001 605.1000 1246.5000 605.2500 ;
	    RECT 1251.9000 605.1000 1253.7001 605.2500 ;
	    RECT 95.1000 600.7500 96.9000 600.9000 ;
	    RECT 145.5000 600.7500 147.3000 600.9000 ;
	    RECT 95.1000 599.2500 147.3000 600.7500 ;
	    RECT 95.1000 599.1000 96.9000 599.2500 ;
	    RECT 145.5000 599.1000 147.3000 599.2500 ;
	    RECT 236.7000 600.7500 238.5000 600.9000 ;
	    RECT 267.9000 600.7500 269.7000 600.9000 ;
	    RECT 236.7000 599.2500 269.7000 600.7500 ;
	    RECT 236.7000 599.1000 238.5000 599.2500 ;
	    RECT 267.9000 599.1000 269.7000 599.2500 ;
	    RECT 291.9000 600.7500 293.7000 600.9000 ;
	    RECT 320.7000 600.7500 322.5000 600.9000 ;
	    RECT 291.9000 599.2500 322.5000 600.7500 ;
	    RECT 291.9000 599.1000 293.7000 599.2500 ;
	    RECT 320.7000 599.1000 322.5000 599.2500 ;
	    RECT 359.1000 600.7500 360.9000 600.9000 ;
	    RECT 383.1000 600.7500 384.9000 600.9000 ;
	    RECT 359.1000 599.2500 384.9000 600.7500 ;
	    RECT 359.1000 599.1000 360.9000 599.2500 ;
	    RECT 383.1000 599.1000 384.9000 599.2500 ;
	    RECT 627.9000 600.7500 629.7000 600.9000 ;
	    RECT 642.3000 600.7500 644.1000 600.9000 ;
	    RECT 627.9000 599.2500 644.1000 600.7500 ;
	    RECT 627.9000 599.1000 629.7000 599.2500 ;
	    RECT 642.3000 599.1000 644.1000 599.2500 ;
	    RECT 855.9000 600.7500 857.7000 600.9000 ;
	    RECT 908.7000 600.7500 910.5000 600.9000 ;
	    RECT 855.9000 599.2500 910.5000 600.7500 ;
	    RECT 855.9000 599.1000 857.7000 599.2500 ;
	    RECT 908.7000 599.1000 910.5000 599.2500 ;
	    RECT 949.5000 600.7500 951.3000 600.9000 ;
	    RECT 961.5000 600.7500 963.3000 600.9000 ;
	    RECT 1170.3000 600.7500 1172.1000 600.9000 ;
	    RECT 949.5000 599.2500 963.3000 600.7500 ;
	    RECT 949.5000 599.1000 951.3000 599.2500 ;
	    RECT 961.5000 599.1000 963.3000 599.2500 ;
	    RECT 1136.8500 599.2500 1172.1000 600.7500 ;
	    RECT 133.5000 594.7500 135.3000 594.9000 ;
	    RECT 174.3000 594.7500 176.1000 594.9000 ;
	    RECT 133.5000 593.2500 176.1000 594.7500 ;
	    RECT 133.5000 593.1000 135.3000 593.2500 ;
	    RECT 174.3000 593.1000 176.1000 593.2500 ;
	    RECT 267.9000 594.7500 269.7000 594.9000 ;
	    RECT 279.9000 594.7500 281.7000 594.9000 ;
	    RECT 267.9000 593.2500 281.7000 594.7500 ;
	    RECT 267.9000 593.1000 269.7000 593.2500 ;
	    RECT 279.9000 593.1000 281.7000 593.2500 ;
	    RECT 402.3000 594.7500 404.1000 594.9000 ;
	    RECT 488.7000 594.7500 490.5000 594.9000 ;
	    RECT 402.3000 593.2500 490.5000 594.7500 ;
	    RECT 402.3000 593.1000 404.1000 593.2500 ;
	    RECT 488.7000 593.1000 490.5000 593.2500 ;
	    RECT 728.7000 594.7500 730.5000 594.9000 ;
	    RECT 779.1000 594.7500 780.9000 594.9000 ;
	    RECT 728.7000 593.2500 780.9000 594.7500 ;
	    RECT 728.7000 593.1000 730.5000 593.2500 ;
	    RECT 779.1000 593.1000 780.9000 593.2500 ;
	    RECT 1095.9000 594.7500 1097.7001 594.9000 ;
	    RECT 1136.8500 594.7500 1138.3500 599.2500 ;
	    RECT 1170.3000 599.1000 1172.1000 599.2500 ;
	    RECT 1095.9000 593.2500 1138.3500 594.7500 ;
	    RECT 1201.5000 594.7500 1203.3000 594.9000 ;
	    RECT 1280.7001 594.7500 1282.5000 594.9000 ;
	    RECT 1311.9000 594.7500 1313.7001 594.9000 ;
	    RECT 1201.5000 593.2500 1313.7001 594.7500 ;
	    RECT 1095.9000 593.1000 1097.7001 593.2500 ;
	    RECT 1201.5000 593.1000 1203.3000 593.2500 ;
	    RECT 1280.7001 593.1000 1282.5000 593.2500 ;
	    RECT 1311.9000 593.1000 1313.7001 593.2500 ;
	    RECT 1335.9000 594.7500 1337.7001 594.9000 ;
	    RECT 1383.9000 594.7500 1385.7001 594.9000 ;
	    RECT 1335.9000 593.2500 1385.7001 594.7500 ;
	    RECT 1335.9000 593.1000 1337.7001 593.2500 ;
	    RECT 1383.9000 593.1000 1385.7001 593.2500 ;
	    RECT 1422.3000 594.7500 1424.1000 594.9000 ;
	    RECT 1434.3000 594.7500 1436.1000 594.9000 ;
	    RECT 1422.3000 593.2500 1436.1000 594.7500 ;
	    RECT 1422.3000 593.1000 1424.1000 593.2500 ;
	    RECT 1434.3000 593.1000 1436.1000 593.2500 ;
	    RECT 90.3000 588.7500 92.1000 588.9000 ;
	    RECT 181.5000 588.7500 183.3000 588.9000 ;
	    RECT 90.3000 587.2500 183.3000 588.7500 ;
	    RECT 90.3000 587.1000 92.1000 587.2500 ;
	    RECT 181.5000 587.1000 183.3000 587.2500 ;
	    RECT 347.1000 588.7500 348.9000 588.9000 ;
	    RECT 359.1000 588.7500 360.9000 588.9000 ;
	    RECT 347.1000 587.2500 360.9000 588.7500 ;
	    RECT 347.1000 587.1000 348.9000 587.2500 ;
	    RECT 359.1000 587.1000 360.9000 587.2500 ;
	    RECT 421.5000 588.7500 423.3000 588.9000 ;
	    RECT 457.5000 588.7500 459.3000 588.9000 ;
	    RECT 421.5000 587.2500 459.3000 588.7500 ;
	    RECT 421.5000 587.1000 423.3000 587.2500 ;
	    RECT 457.5000 587.1000 459.3000 587.2500 ;
	    RECT 584.7000 588.7500 586.5000 588.9000 ;
	    RECT 599.1000 588.7500 600.9000 588.9000 ;
	    RECT 584.7000 587.2500 600.9000 588.7500 ;
	    RECT 584.7000 587.1000 586.5000 587.2500 ;
	    RECT 599.1000 587.1000 600.9000 587.2500 ;
	    RECT 632.7000 588.7500 634.5000 588.9000 ;
	    RECT 733.5000 588.7500 735.3000 588.9000 ;
	    RECT 632.7000 587.2500 735.3000 588.7500 ;
	    RECT 632.7000 587.1000 634.5000 587.2500 ;
	    RECT 733.5000 587.1000 735.3000 587.2500 ;
	    RECT 788.7000 588.7500 790.5000 588.9000 ;
	    RECT 824.7000 588.7500 826.5000 588.9000 ;
	    RECT 788.7000 587.2500 826.5000 588.7500 ;
	    RECT 788.7000 587.1000 790.5000 587.2500 ;
	    RECT 824.7000 587.1000 826.5000 587.2500 ;
	    RECT 836.7000 588.7500 838.5000 588.9000 ;
	    RECT 843.9000 588.7500 845.7000 588.9000 ;
	    RECT 860.7000 588.7500 862.5000 588.9000 ;
	    RECT 836.7000 587.2500 862.5000 588.7500 ;
	    RECT 836.7000 587.1000 838.5000 587.2500 ;
	    RECT 843.9000 587.1000 845.7000 587.2500 ;
	    RECT 860.7000 587.1000 862.5000 587.2500 ;
	    RECT 1155.9000 588.7500 1157.7001 588.9000 ;
	    RECT 1167.9000 588.7500 1169.7001 588.9000 ;
	    RECT 1155.9000 587.2500 1169.7001 588.7500 ;
	    RECT 1155.9000 587.1000 1157.7001 587.2500 ;
	    RECT 1167.9000 587.1000 1169.7001 587.2500 ;
	    RECT 1283.1000 588.7500 1284.9000 588.9000 ;
	    RECT 1331.1000 588.7500 1332.9000 588.9000 ;
	    RECT 1283.1000 587.2500 1332.9000 588.7500 ;
	    RECT 1283.1000 587.1000 1284.9000 587.2500 ;
	    RECT 1331.1000 587.1000 1332.9000 587.2500 ;
	    RECT 1335.9000 588.7500 1337.7001 588.9000 ;
	    RECT 1403.1000 588.7500 1404.9000 588.9000 ;
	    RECT 1335.9000 587.2500 1404.9000 588.7500 ;
	    RECT 1335.9000 587.1000 1337.7001 587.2500 ;
	    RECT 1403.1000 587.1000 1404.9000 587.2500 ;
	    RECT 1463.1000 588.7500 1464.9000 588.9000 ;
	    RECT 1491.9000 588.7500 1493.7001 588.9000 ;
	    RECT 1463.1000 587.2500 1493.7001 588.7500 ;
	    RECT 1463.1000 587.1000 1464.9000 587.2500 ;
	    RECT 1491.9000 587.1000 1493.7001 587.2500 ;
	    RECT 584.7000 584.1000 586.5000 585.9000 ;
	    RECT 135.9000 582.7500 137.7000 582.9000 ;
	    RECT 164.7000 582.7500 166.5000 582.9000 ;
	    RECT 183.9000 582.7500 185.7000 582.9000 ;
	    RECT 135.9000 581.2500 185.7000 582.7500 ;
	    RECT 135.9000 581.1000 137.7000 581.2500 ;
	    RECT 164.7000 581.1000 166.5000 581.2500 ;
	    RECT 183.9000 581.1000 185.7000 581.2500 ;
	    RECT 210.3000 582.7500 212.1000 582.9000 ;
	    RECT 215.1000 582.7500 216.9000 582.9000 ;
	    RECT 210.3000 581.2500 216.9000 582.7500 ;
	    RECT 210.3000 581.1000 212.1000 581.2500 ;
	    RECT 215.1000 581.1000 216.9000 581.2500 ;
	    RECT 277.5000 582.7500 279.3000 582.9000 ;
	    RECT 287.1000 582.7500 288.9000 582.9000 ;
	    RECT 277.5000 581.2500 288.9000 582.7500 ;
	    RECT 277.5000 581.1000 279.3000 581.2500 ;
	    RECT 287.1000 581.1000 288.9000 581.2500 ;
	    RECT 359.1000 582.7500 360.9000 582.9000 ;
	    RECT 385.5000 582.7500 387.3000 582.9000 ;
	    RECT 359.1000 581.2500 387.3000 582.7500 ;
	    RECT 359.1000 581.1000 360.9000 581.2500 ;
	    RECT 385.5000 581.1000 387.3000 581.2500 ;
	    RECT 483.9000 582.7500 485.7000 582.9000 ;
	    RECT 536.7000 582.7500 538.5000 582.9000 ;
	    RECT 483.9000 581.2500 538.5000 582.7500 ;
	    RECT 483.9000 581.1000 485.7000 581.2500 ;
	    RECT 536.7000 581.1000 538.5000 581.2500 ;
	    RECT 107.1000 576.7500 108.9000 576.9000 ;
	    RECT 176.7000 576.7500 178.5000 576.9000 ;
	    RECT 107.1000 575.2500 178.5000 576.7500 ;
	    RECT 107.1000 575.1000 108.9000 575.2500 ;
	    RECT 176.7000 575.1000 178.5000 575.2500 ;
	    RECT 181.5000 576.7500 183.3000 576.9000 ;
	    RECT 279.9000 576.7500 281.7000 576.9000 ;
	    RECT 181.5000 575.2500 281.7000 576.7500 ;
	    RECT 181.5000 575.1000 183.3000 575.2500 ;
	    RECT 279.9000 575.1000 281.7000 575.2500 ;
	    RECT 289.5000 576.7500 291.3000 576.9000 ;
	    RECT 347.1000 576.7500 348.9000 576.9000 ;
	    RECT 289.5000 575.2500 348.9000 576.7500 ;
	    RECT 289.5000 575.1000 291.3000 575.2500 ;
	    RECT 347.1000 575.1000 348.9000 575.2500 ;
	    RECT 361.5000 576.7500 363.3000 576.9000 ;
	    RECT 426.3000 576.7500 428.1000 576.9000 ;
	    RECT 361.5000 575.2500 428.1000 576.7500 ;
	    RECT 361.5000 575.1000 363.3000 575.2500 ;
	    RECT 426.3000 575.1000 428.1000 575.2500 ;
	    RECT 486.3000 576.7500 488.1000 576.9000 ;
	    RECT 503.1000 576.7500 504.9000 576.9000 ;
	    RECT 515.1000 576.7500 516.9000 576.9000 ;
	    RECT 486.3000 575.2500 516.9000 576.7500 ;
	    RECT 486.3000 575.1000 488.1000 575.2500 ;
	    RECT 503.1000 575.1000 504.9000 575.2500 ;
	    RECT 515.1000 575.1000 516.9000 575.2500 ;
	    RECT 524.7000 576.7500 526.5000 576.9000 ;
	    RECT 536.7000 576.7500 538.5000 576.9000 ;
	    RECT 524.7000 575.2500 538.5000 576.7500 ;
	    RECT 584.8500 576.7500 586.3500 584.1000 ;
	    RECT 747.9000 582.7500 749.7000 582.9000 ;
	    RECT 759.9000 582.7500 761.7000 582.9000 ;
	    RECT 747.9000 581.2500 761.7000 582.7500 ;
	    RECT 747.9000 581.1000 749.7000 581.2500 ;
	    RECT 759.9000 581.1000 761.7000 581.2500 ;
	    RECT 817.5000 582.7500 819.3000 582.9000 ;
	    RECT 875.1000 582.7500 876.9000 582.9000 ;
	    RECT 817.5000 581.2500 876.9000 582.7500 ;
	    RECT 817.5000 581.1000 819.3000 581.2500 ;
	    RECT 875.1000 581.1000 876.9000 581.2500 ;
	    RECT 956.7000 582.7500 958.5000 582.9000 ;
	    RECT 963.9000 582.7500 965.7000 582.9000 ;
	    RECT 956.7000 581.2500 965.7000 582.7500 ;
	    RECT 956.7000 581.1000 958.5000 581.2500 ;
	    RECT 963.9000 581.1000 965.7000 581.2500 ;
	    RECT 1035.9000 582.7500 1037.7001 582.9000 ;
	    RECT 1129.5000 582.7500 1131.3000 582.9000 ;
	    RECT 1035.9000 581.2500 1131.3000 582.7500 ;
	    RECT 1035.9000 581.1000 1037.7001 581.2500 ;
	    RECT 1129.5000 581.1000 1131.3000 581.2500 ;
	    RECT 1167.9000 582.7500 1169.7001 582.9000 ;
	    RECT 1179.9000 582.7500 1181.7001 582.9000 ;
	    RECT 1263.9000 582.7500 1265.7001 582.9000 ;
	    RECT 1167.9000 581.2500 1265.7001 582.7500 ;
	    RECT 1167.9000 581.1000 1169.7001 581.2500 ;
	    RECT 1179.9000 581.1000 1181.7001 581.2500 ;
	    RECT 1263.9000 581.1000 1265.7001 581.2500 ;
	    RECT 1280.7001 582.7500 1282.5000 582.9000 ;
	    RECT 1311.9000 582.7500 1313.7001 582.9000 ;
	    RECT 1280.7001 581.2500 1313.7001 582.7500 ;
	    RECT 1280.7001 581.1000 1282.5000 581.2500 ;
	    RECT 1311.9000 581.1000 1313.7001 581.2500 ;
	    RECT 1328.7001 582.7500 1330.5000 582.9000 ;
	    RECT 1405.5000 582.7500 1407.3000 582.9000 ;
	    RECT 1328.7001 581.2500 1407.3000 582.7500 ;
	    RECT 1328.7001 581.1000 1330.5000 581.2500 ;
	    RECT 1405.5000 581.1000 1407.3000 581.2500 ;
	    RECT 1460.7001 582.7500 1462.5000 582.9000 ;
	    RECT 1494.3000 582.7500 1496.1000 582.9000 ;
	    RECT 1460.7001 581.2500 1496.1000 582.7500 ;
	    RECT 1460.7001 581.1000 1462.5000 581.2500 ;
	    RECT 1494.3000 581.1000 1496.1000 581.2500 ;
	    RECT 1542.3000 582.7500 1544.1000 582.9000 ;
	    RECT 1556.7001 582.7500 1558.5000 582.9000 ;
	    RECT 1542.3000 581.2500 1558.5000 582.7500 ;
	    RECT 1542.3000 581.1000 1544.1000 581.2500 ;
	    RECT 1556.7001 581.1000 1558.5000 581.2500 ;
	    RECT 589.5000 576.7500 591.3000 576.9000 ;
	    RECT 584.8500 575.2500 591.3000 576.7500 ;
	    RECT 524.7000 575.1000 526.5000 575.2500 ;
	    RECT 536.7000 575.1000 538.5000 575.2500 ;
	    RECT 589.5000 575.1000 591.3000 575.2500 ;
	    RECT 675.9000 576.7500 677.7000 576.9000 ;
	    RECT 743.1000 576.7500 744.9000 576.9000 ;
	    RECT 675.9000 575.2500 744.9000 576.7500 ;
	    RECT 675.9000 575.1000 677.7000 575.2500 ;
	    RECT 743.1000 575.1000 744.9000 575.2500 ;
	    RECT 759.9000 576.7500 761.7000 576.9000 ;
	    RECT 863.1000 576.7500 864.9000 576.9000 ;
	    RECT 759.9000 575.2500 864.9000 576.7500 ;
	    RECT 759.9000 575.1000 761.7000 575.2500 ;
	    RECT 863.1000 575.1000 864.9000 575.2500 ;
	    RECT 978.3000 576.7500 980.1000 576.9000 ;
	    RECT 1016.7000 576.7500 1018.5000 576.9000 ;
	    RECT 978.3000 575.2500 1018.5000 576.7500 ;
	    RECT 978.3000 575.1000 980.1000 575.2500 ;
	    RECT 1016.7000 575.1000 1018.5000 575.2500 ;
	    RECT 1043.1000 576.7500 1044.9000 576.9000 ;
	    RECT 1127.1000 576.7500 1128.9000 576.9000 ;
	    RECT 1043.1000 575.2500 1128.9000 576.7500 ;
	    RECT 1043.1000 575.1000 1044.9000 575.2500 ;
	    RECT 1127.1000 575.1000 1128.9000 575.2500 ;
	    RECT 1299.9000 576.7500 1301.7001 576.9000 ;
	    RECT 1333.5000 576.7500 1335.3000 576.9000 ;
	    RECT 1299.9000 575.2500 1335.3000 576.7500 ;
	    RECT 1299.9000 575.1000 1301.7001 575.2500 ;
	    RECT 1333.5000 575.1000 1335.3000 575.2500 ;
	    RECT 1338.3000 576.7500 1340.1000 576.9000 ;
	    RECT 1374.3000 576.7500 1376.1000 576.9000 ;
	    RECT 1338.3000 575.2500 1376.1000 576.7500 ;
	    RECT 1338.3000 575.1000 1340.1000 575.2500 ;
	    RECT 1374.3000 575.1000 1376.1000 575.2500 ;
	    RECT 1419.9000 576.7500 1421.7001 576.9000 ;
	    RECT 1451.1000 576.7500 1452.9000 576.9000 ;
	    RECT 1419.9000 575.2500 1452.9000 576.7500 ;
	    RECT 1419.9000 575.1000 1421.7001 575.2500 ;
	    RECT 1451.1000 575.1000 1452.9000 575.2500 ;
	    RECT 1520.7001 576.7500 1522.5000 576.9000 ;
	    RECT 1544.7001 576.7500 1546.5000 576.9000 ;
	    RECT 1520.7001 575.2500 1546.5000 576.7500 ;
	    RECT 1520.7001 575.1000 1522.5000 575.2500 ;
	    RECT 1544.7001 575.1000 1546.5000 575.2500 ;
	    RECT 212.7000 570.7500 214.5000 570.9000 ;
	    RECT 224.7000 570.7500 226.5000 570.9000 ;
	    RECT 212.7000 569.2500 226.5000 570.7500 ;
	    RECT 212.7000 569.1000 214.5000 569.2500 ;
	    RECT 224.7000 569.1000 226.5000 569.2500 ;
	    RECT 301.5000 570.7500 303.3000 570.9000 ;
	    RECT 409.5000 570.7500 411.3000 570.9000 ;
	    RECT 301.5000 569.2500 411.3000 570.7500 ;
	    RECT 301.5000 569.1000 303.3000 569.2500 ;
	    RECT 409.5000 569.1000 411.3000 569.2500 ;
	    RECT 510.3000 570.7500 512.1000 570.9000 ;
	    RECT 582.3000 570.7500 584.1000 570.9000 ;
	    RECT 608.7000 570.7500 610.5000 570.9000 ;
	    RECT 510.3000 569.2500 610.5000 570.7500 ;
	    RECT 510.3000 569.1000 512.1000 569.2500 ;
	    RECT 582.3000 569.1000 584.1000 569.2500 ;
	    RECT 608.7000 569.1000 610.5000 569.2500 ;
	    RECT 711.9000 570.7500 713.7000 570.9000 ;
	    RECT 726.3000 570.7500 728.1000 570.9000 ;
	    RECT 711.9000 569.2500 728.1000 570.7500 ;
	    RECT 711.9000 569.1000 713.7000 569.2500 ;
	    RECT 726.3000 569.1000 728.1000 569.2500 ;
	    RECT 971.1000 570.7500 972.9000 570.9000 ;
	    RECT 975.9000 570.7500 977.7000 570.9000 ;
	    RECT 971.1000 569.2500 977.7000 570.7500 ;
	    RECT 971.1000 569.1000 972.9000 569.2500 ;
	    RECT 975.9000 569.1000 977.7000 569.2500 ;
	    RECT 1093.5000 570.7500 1095.3000 570.9000 ;
	    RECT 1155.9000 570.7500 1157.7001 570.9000 ;
	    RECT 1093.5000 569.2500 1157.7001 570.7500 ;
	    RECT 1093.5000 569.1000 1095.3000 569.2500 ;
	    RECT 1155.9000 569.1000 1157.7001 569.2500 ;
	    RECT 1177.5000 570.7500 1179.3000 570.9000 ;
	    RECT 1227.9000 570.7500 1229.7001 570.9000 ;
	    RECT 1177.5000 569.2500 1229.7001 570.7500 ;
	    RECT 1177.5000 569.1000 1179.3000 569.2500 ;
	    RECT 1227.9000 569.1000 1229.7001 569.2500 ;
	    RECT 1261.5000 570.7500 1263.3000 570.9000 ;
	    RECT 1287.9000 570.7500 1289.7001 570.9000 ;
	    RECT 1299.9000 570.7500 1301.7001 570.9000 ;
	    RECT 1261.5000 569.2500 1301.7001 570.7500 ;
	    RECT 1261.5000 569.1000 1263.3000 569.2500 ;
	    RECT 1287.9000 569.1000 1289.7001 569.2500 ;
	    RECT 1299.9000 569.1000 1301.7001 569.2500 ;
	    RECT 1331.1000 570.7500 1332.9000 570.9000 ;
	    RECT 1347.9000 570.7500 1349.7001 570.9000 ;
	    RECT 1331.1000 569.2500 1349.7001 570.7500 ;
	    RECT 1331.1000 569.1000 1332.9000 569.2500 ;
	    RECT 1347.9000 569.1000 1349.7001 569.2500 ;
	    RECT 1489.5000 570.7500 1491.3000 570.9000 ;
	    RECT 1515.9000 570.7500 1517.7001 570.9000 ;
	    RECT 1489.5000 569.2500 1517.7001 570.7500 ;
	    RECT 1489.5000 569.1000 1491.3000 569.2500 ;
	    RECT 1515.9000 569.1000 1517.7001 569.2500 ;
	    RECT 18.3000 564.7500 20.1000 564.9000 ;
	    RECT 56.7000 564.7500 58.5000 564.9000 ;
	    RECT 78.3000 564.7500 80.1000 564.9000 ;
	    RECT 102.3000 564.7500 104.1000 564.9000 ;
	    RECT 18.3000 563.2500 104.1000 564.7500 ;
	    RECT 18.3000 563.1000 20.1000 563.2500 ;
	    RECT 56.7000 563.1000 58.5000 563.2500 ;
	    RECT 78.3000 563.1000 80.1000 563.2500 ;
	    RECT 102.3000 563.1000 104.1000 563.2500 ;
	    RECT 198.3000 564.7500 200.1000 564.9000 ;
	    RECT 275.1000 564.7500 276.9000 564.9000 ;
	    RECT 198.3000 563.2500 276.9000 564.7500 ;
	    RECT 198.3000 563.1000 200.1000 563.2500 ;
	    RECT 275.1000 563.1000 276.9000 563.2500 ;
	    RECT 315.9000 564.7500 317.7000 564.9000 ;
	    RECT 330.3000 564.7500 332.1000 564.9000 ;
	    RECT 315.9000 563.2500 332.1000 564.7500 ;
	    RECT 315.9000 563.1000 317.7000 563.2500 ;
	    RECT 330.3000 563.1000 332.1000 563.2500 ;
	    RECT 488.7000 564.7500 490.5000 564.9000 ;
	    RECT 531.9000 564.7500 533.7000 564.9000 ;
	    RECT 488.7000 563.2500 533.7000 564.7500 ;
	    RECT 488.7000 563.1000 490.5000 563.2500 ;
	    RECT 531.9000 563.1000 533.7000 563.2500 ;
	    RECT 601.5000 564.7500 603.3000 564.9000 ;
	    RECT 618.3000 564.7500 620.1000 564.9000 ;
	    RECT 601.5000 563.2500 620.1000 564.7500 ;
	    RECT 601.5000 563.1000 603.3000 563.2500 ;
	    RECT 618.3000 563.1000 620.1000 563.2500 ;
	    RECT 733.5000 564.7500 735.3000 564.9000 ;
	    RECT 889.5000 564.7500 891.3000 564.9000 ;
	    RECT 733.5000 563.2500 891.3000 564.7500 ;
	    RECT 733.5000 563.1000 735.3000 563.2500 ;
	    RECT 889.5000 563.1000 891.3000 563.2500 ;
	    RECT 959.1000 564.7500 960.9000 564.9000 ;
	    RECT 1091.1000 564.7500 1092.9000 564.9000 ;
	    RECT 959.1000 563.2500 1092.9000 564.7500 ;
	    RECT 959.1000 563.1000 960.9000 563.2500 ;
	    RECT 1091.1000 563.1000 1092.9000 563.2500 ;
	    RECT 1098.3000 564.7500 1100.1000 564.9000 ;
	    RECT 1141.5000 564.7500 1143.3000 564.9000 ;
	    RECT 1098.3000 563.2500 1143.3000 564.7500 ;
	    RECT 1098.3000 563.1000 1100.1000 563.2500 ;
	    RECT 1141.5000 563.1000 1143.3000 563.2500 ;
	    RECT 1227.9000 564.7500 1229.7001 564.9000 ;
	    RECT 1249.5000 564.7500 1251.3000 564.9000 ;
	    RECT 1227.9000 563.2500 1251.3000 564.7500 ;
	    RECT 1227.9000 563.1000 1229.7001 563.2500 ;
	    RECT 1249.5000 563.1000 1251.3000 563.2500 ;
	    RECT 1347.9000 564.7500 1349.7001 564.9000 ;
	    RECT 1355.1000 564.7500 1356.9000 564.9000 ;
	    RECT 1347.9000 563.2500 1356.9000 564.7500 ;
	    RECT 1347.9000 563.1000 1349.7001 563.2500 ;
	    RECT 1355.1000 563.1000 1356.9000 563.2500 ;
	    RECT 1484.7001 564.7500 1486.5000 564.9000 ;
	    RECT 1496.7001 564.7500 1498.5000 564.9000 ;
	    RECT 1484.7001 563.2500 1498.5000 564.7500 ;
	    RECT 1484.7001 563.1000 1486.5000 563.2500 ;
	    RECT 1496.7001 563.1000 1498.5000 563.2500 ;
	    RECT 39.9000 558.7500 41.7000 558.9000 ;
	    RECT 92.7000 558.7500 94.5000 558.9000 ;
	    RECT 131.1000 558.7500 132.9000 558.9000 ;
	    RECT 39.9000 557.2500 132.9000 558.7500 ;
	    RECT 39.9000 557.1000 41.7000 557.2500 ;
	    RECT 92.7000 557.1000 94.5000 557.2500 ;
	    RECT 131.1000 557.1000 132.9000 557.2500 ;
	    RECT 162.3000 558.7500 164.1000 558.9000 ;
	    RECT 275.1000 558.7500 276.9000 558.9000 ;
	    RECT 303.9000 558.7500 305.7000 558.9000 ;
	    RECT 162.3000 557.2500 305.7000 558.7500 ;
	    RECT 162.3000 557.1000 164.1000 557.2500 ;
	    RECT 275.1000 557.1000 276.9000 557.2500 ;
	    RECT 303.9000 557.1000 305.7000 557.2500 ;
	    RECT 330.3000 558.7500 332.1000 558.9000 ;
	    RECT 344.7000 558.7500 346.5000 558.9000 ;
	    RECT 330.3000 557.2500 346.5000 558.7500 ;
	    RECT 330.3000 557.1000 332.1000 557.2500 ;
	    RECT 344.7000 557.1000 346.5000 557.2500 ;
	    RECT 354.3000 558.7500 356.1000 558.9000 ;
	    RECT 390.3000 558.7500 392.1000 558.9000 ;
	    RECT 354.3000 557.2500 392.1000 558.7500 ;
	    RECT 354.3000 557.1000 356.1000 557.2500 ;
	    RECT 390.3000 557.1000 392.1000 557.2500 ;
	    RECT 709.5000 558.7500 711.3000 558.9000 ;
	    RECT 848.7000 558.7500 850.5000 558.9000 ;
	    RECT 709.5000 557.2500 850.5000 558.7500 ;
	    RECT 709.5000 557.1000 711.3000 557.2500 ;
	    RECT 848.7000 557.1000 850.5000 557.2500 ;
	    RECT 858.3000 558.7500 860.1000 558.9000 ;
	    RECT 863.1000 558.7500 864.9000 558.9000 ;
	    RECT 858.3000 557.2500 864.9000 558.7500 ;
	    RECT 858.3000 557.1000 860.1000 557.2500 ;
	    RECT 863.1000 557.1000 864.9000 557.2500 ;
	    RECT 1103.1000 558.7500 1104.9000 558.9000 ;
	    RECT 1143.9000 558.7500 1145.7001 558.9000 ;
	    RECT 1165.5000 558.7500 1167.3000 558.9000 ;
	    RECT 1170.3000 558.7500 1172.1000 558.9000 ;
	    RECT 1103.1000 557.2500 1172.1000 558.7500 ;
	    RECT 1103.1000 557.1000 1104.9000 557.2500 ;
	    RECT 1143.9000 557.1000 1145.7001 557.2500 ;
	    RECT 1165.5000 557.1000 1167.3000 557.2500 ;
	    RECT 1170.3000 557.1000 1172.1000 557.2500 ;
	    RECT 1208.7001 558.7500 1210.5000 558.9000 ;
	    RECT 1232.7001 558.7500 1234.5000 558.9000 ;
	    RECT 1208.7001 557.2500 1234.5000 558.7500 ;
	    RECT 1208.7001 557.1000 1210.5000 557.2500 ;
	    RECT 1232.7001 557.1000 1234.5000 557.2500 ;
	    RECT 1249.5000 558.7500 1251.3000 558.9000 ;
	    RECT 1280.7001 558.7500 1282.5000 558.9000 ;
	    RECT 1249.5000 557.2500 1282.5000 558.7500 ;
	    RECT 1249.5000 557.1000 1251.3000 557.2500 ;
	    RECT 1280.7001 557.1000 1282.5000 557.2500 ;
	    RECT 1427.1000 558.7500 1428.9000 558.9000 ;
	    RECT 1482.3000 558.7500 1484.1000 558.9000 ;
	    RECT 1427.1000 557.2500 1484.1000 558.7500 ;
	    RECT 1427.1000 557.1000 1428.9000 557.2500 ;
	    RECT 1482.3000 557.1000 1484.1000 557.2500 ;
	    RECT 327.9000 552.7500 329.7000 552.9000 ;
	    RECT 356.7000 552.7500 358.5000 552.9000 ;
	    RECT 327.9000 551.2500 358.5000 552.7500 ;
	    RECT 327.9000 551.1000 329.7000 551.2500 ;
	    RECT 356.7000 551.1000 358.5000 551.2500 ;
	    RECT 519.9000 552.7500 521.7000 552.9000 ;
	    RECT 560.7000 552.7500 562.5000 552.9000 ;
	    RECT 519.9000 551.2500 562.5000 552.7500 ;
	    RECT 519.9000 551.1000 521.7000 551.2500 ;
	    RECT 560.7000 551.1000 562.5000 551.2500 ;
	    RECT 637.5000 552.7500 639.3000 552.9000 ;
	    RECT 651.9000 552.7500 653.7000 552.9000 ;
	    RECT 711.9000 552.7500 713.7000 552.9000 ;
	    RECT 637.5000 551.2500 713.7000 552.7500 ;
	    RECT 637.5000 551.1000 639.3000 551.2500 ;
	    RECT 651.9000 551.1000 653.7000 551.2500 ;
	    RECT 711.9000 551.1000 713.7000 551.2500 ;
	    RECT 858.3000 552.7500 860.1000 552.9000 ;
	    RECT 877.5000 552.7500 879.3000 552.9000 ;
	    RECT 887.1000 552.7500 888.9000 552.9000 ;
	    RECT 858.3000 551.2500 888.9000 552.7500 ;
	    RECT 858.3000 551.1000 860.1000 551.2500 ;
	    RECT 877.5000 551.1000 879.3000 551.2500 ;
	    RECT 887.1000 551.1000 888.9000 551.2500 ;
	    RECT 968.7000 552.7500 970.5000 552.9000 ;
	    RECT 978.3000 552.7500 980.1000 552.9000 ;
	    RECT 968.7000 551.2500 980.1000 552.7500 ;
	    RECT 968.7000 551.1000 970.5000 551.2500 ;
	    RECT 978.3000 551.1000 980.1000 551.2500 ;
	    RECT 1134.3000 552.7500 1136.1000 552.9000 ;
	    RECT 1167.9000 552.7500 1169.7001 552.9000 ;
	    RECT 1134.3000 551.2500 1169.7001 552.7500 ;
	    RECT 1134.3000 551.1000 1136.1000 551.2500 ;
	    RECT 1167.9000 551.1000 1169.7001 551.2500 ;
	    RECT 1235.1000 552.7500 1236.9000 552.9000 ;
	    RECT 1261.5000 552.7500 1263.3000 552.9000 ;
	    RECT 1235.1000 551.2500 1263.3000 552.7500 ;
	    RECT 1235.1000 551.1000 1236.9000 551.2500 ;
	    RECT 1261.5000 551.1000 1263.3000 551.2500 ;
	    RECT 1347.9000 552.7500 1349.7001 552.9000 ;
	    RECT 1369.5000 552.7500 1371.3000 552.9000 ;
	    RECT 1347.9000 551.2500 1371.3000 552.7500 ;
	    RECT 1347.9000 551.1000 1349.7001 551.2500 ;
	    RECT 1369.5000 551.1000 1371.3000 551.2500 ;
	    RECT 1417.5000 552.7500 1419.3000 552.9000 ;
	    RECT 1422.3000 552.7500 1424.1000 552.9000 ;
	    RECT 1417.5000 551.2500 1424.1000 552.7500 ;
	    RECT 1417.5000 551.1000 1419.3000 551.2500 ;
	    RECT 1422.3000 551.1000 1424.1000 551.2500 ;
	    RECT 1477.5000 552.7500 1479.3000 552.9000 ;
	    RECT 1511.1000 552.7500 1512.9000 552.9000 ;
	    RECT 1477.5000 551.2500 1512.9000 552.7500 ;
	    RECT 1477.5000 551.1000 1479.3000 551.2500 ;
	    RECT 1511.1000 551.1000 1512.9000 551.2500 ;
	    RECT 241.5000 546.7500 243.3000 546.9000 ;
	    RECT 272.7000 546.7500 274.5000 546.9000 ;
	    RECT 241.5000 545.2500 274.5000 546.7500 ;
	    RECT 241.5000 545.1000 243.3000 545.2500 ;
	    RECT 272.7000 545.1000 274.5000 545.2500 ;
	    RECT 337.5000 546.7500 339.3000 546.9000 ;
	    RECT 351.9000 546.7500 353.7000 546.9000 ;
	    RECT 337.5000 545.2500 353.7000 546.7500 ;
	    RECT 337.5000 545.1000 339.3000 545.2500 ;
	    RECT 351.9000 545.1000 353.7000 545.2500 ;
	    RECT 517.5000 546.7500 519.3000 546.9000 ;
	    RECT 587.1000 546.7500 588.9000 546.9000 ;
	    RECT 517.5000 545.2500 588.9000 546.7500 ;
	    RECT 517.5000 545.1000 519.3000 545.2500 ;
	    RECT 587.1000 545.1000 588.9000 545.2500 ;
	    RECT 1141.5000 546.7500 1143.3000 546.9000 ;
	    RECT 1175.1000 546.7500 1176.9000 546.9000 ;
	    RECT 1203.9000 546.7500 1205.7001 546.9000 ;
	    RECT 1141.5000 545.2500 1205.7001 546.7500 ;
	    RECT 1141.5000 545.1000 1143.3000 545.2500 ;
	    RECT 1175.1000 545.1000 1176.9000 545.2500 ;
	    RECT 1203.9000 545.1000 1205.7001 545.2500 ;
	    RECT 1244.7001 546.7500 1246.5000 546.9000 ;
	    RECT 1259.1000 546.7500 1260.9000 546.9000 ;
	    RECT 1244.7001 545.2500 1260.9000 546.7500 ;
	    RECT 1244.7001 545.1000 1246.5000 545.2500 ;
	    RECT 1259.1000 545.1000 1260.9000 545.2500 ;
	    RECT 1422.3000 546.7500 1424.1000 546.9000 ;
	    RECT 1489.5000 546.7500 1491.3000 546.9000 ;
	    RECT 1422.3000 545.2500 1491.3000 546.7500 ;
	    RECT 1422.3000 545.1000 1424.1000 545.2500 ;
	    RECT 1489.5000 545.1000 1491.3000 545.2500 ;
	    RECT 294.3000 540.7500 296.1000 540.9000 ;
	    RECT 354.3000 540.7500 356.1000 540.9000 ;
	    RECT 294.3000 539.2500 356.1000 540.7500 ;
	    RECT 294.3000 539.1000 296.1000 539.2500 ;
	    RECT 354.3000 539.1000 356.1000 539.2500 ;
	    RECT 843.9000 540.7500 845.7000 540.9000 ;
	    RECT 870.3000 540.7500 872.1000 540.9000 ;
	    RECT 843.9000 539.2500 872.1000 540.7500 ;
	    RECT 843.9000 539.1000 845.7000 539.2500 ;
	    RECT 870.3000 539.1000 872.1000 539.2500 ;
	    RECT 1043.1000 540.7500 1044.9000 540.9000 ;
	    RECT 1050.3000 540.7500 1052.1000 540.9000 ;
	    RECT 1043.1000 539.2500 1052.1000 540.7500 ;
	    RECT 1043.1000 539.1000 1044.9000 539.2500 ;
	    RECT 1050.3000 539.1000 1052.1000 539.2500 ;
	    RECT 1059.9000 540.7500 1061.7001 540.9000 ;
	    RECT 1088.7001 540.7500 1090.5000 540.9000 ;
	    RECT 1117.5000 540.7500 1119.3000 540.9000 ;
	    RECT 1059.9000 539.2500 1119.3000 540.7500 ;
	    RECT 1059.9000 539.1000 1061.7001 539.2500 ;
	    RECT 1088.7001 539.1000 1090.5000 539.2500 ;
	    RECT 1117.5000 539.1000 1119.3000 539.2500 ;
	    RECT 1139.1000 540.7500 1140.9000 540.9000 ;
	    RECT 1218.3000 540.7500 1220.1000 540.9000 ;
	    RECT 1139.1000 539.2500 1220.1000 540.7500 ;
	    RECT 1139.1000 539.1000 1140.9000 539.2500 ;
	    RECT 1218.3000 539.1000 1220.1000 539.2500 ;
	    RECT 1232.7001 540.7500 1234.5000 540.9000 ;
	    RECT 1254.3000 540.7500 1256.1000 540.9000 ;
	    RECT 1232.7001 539.2500 1256.1000 540.7500 ;
	    RECT 1232.7001 539.1000 1234.5000 539.2500 ;
	    RECT 1254.3000 539.1000 1256.1000 539.2500 ;
	    RECT 1278.3000 540.7500 1280.1000 540.9000 ;
	    RECT 1326.3000 540.7500 1328.1000 540.9000 ;
	    RECT 1278.3000 539.2500 1328.1000 540.7500 ;
	    RECT 1278.3000 539.1000 1280.1000 539.2500 ;
	    RECT 1326.3000 539.1000 1328.1000 539.2500 ;
	    RECT 1333.5000 540.7500 1335.3000 540.9000 ;
	    RECT 1367.1000 540.7500 1368.9000 540.9000 ;
	    RECT 1333.5000 539.2500 1368.9000 540.7500 ;
	    RECT 1333.5000 539.1000 1335.3000 539.2500 ;
	    RECT 1367.1000 539.1000 1368.9000 539.2500 ;
	    RECT 1424.7001 540.7500 1426.5000 540.9000 ;
	    RECT 1491.9000 540.7500 1493.7001 540.9000 ;
	    RECT 1424.7001 539.2500 1493.7001 540.7500 ;
	    RECT 1424.7001 539.1000 1426.5000 539.2500 ;
	    RECT 1491.9000 539.1000 1493.7001 539.2500 ;
	    RECT 95.1000 534.7500 96.9000 534.9000 ;
	    RECT 143.1000 534.7500 144.9000 534.9000 ;
	    RECT 95.1000 533.2500 144.9000 534.7500 ;
	    RECT 95.1000 533.1000 96.9000 533.2500 ;
	    RECT 143.1000 533.1000 144.9000 533.2500 ;
	    RECT 323.1000 534.7500 324.9000 534.9000 ;
	    RECT 339.9000 534.7500 341.7000 534.9000 ;
	    RECT 323.1000 533.2500 341.7000 534.7500 ;
	    RECT 323.1000 533.1000 324.9000 533.2500 ;
	    RECT 339.9000 533.1000 341.7000 533.2500 ;
	    RECT 565.5000 534.7500 567.3000 534.9000 ;
	    RECT 719.1000 534.7500 720.9000 534.9000 ;
	    RECT 565.5000 533.2500 720.9000 534.7500 ;
	    RECT 565.5000 533.1000 567.3000 533.2500 ;
	    RECT 719.1000 533.1000 720.9000 533.2500 ;
	    RECT 834.3000 534.7500 836.1000 534.9000 ;
	    RECT 851.1000 534.7500 852.9000 534.9000 ;
	    RECT 834.3000 533.2500 852.9000 534.7500 ;
	    RECT 834.3000 533.1000 836.1000 533.2500 ;
	    RECT 851.1000 533.1000 852.9000 533.2500 ;
	    RECT 860.7000 534.7500 862.5000 534.9000 ;
	    RECT 930.3000 534.7500 932.1000 534.9000 ;
	    RECT 860.7000 533.2500 932.1000 534.7500 ;
	    RECT 860.7000 533.1000 862.5000 533.2500 ;
	    RECT 930.3000 533.1000 932.1000 533.2500 ;
	    RECT 973.5000 534.7500 975.3000 534.9000 ;
	    RECT 987.9000 534.7500 989.7000 534.9000 ;
	    RECT 973.5000 533.2500 989.7000 534.7500 ;
	    RECT 973.5000 533.1000 975.3000 533.2500 ;
	    RECT 987.9000 533.1000 989.7000 533.2500 ;
	    RECT 1105.5000 534.7500 1107.3000 534.9000 ;
	    RECT 1172.7001 534.7500 1174.5000 534.9000 ;
	    RECT 1199.1000 534.7500 1200.9000 534.9000 ;
	    RECT 1105.5000 533.2500 1200.9000 534.7500 ;
	    RECT 1105.5000 533.1000 1107.3000 533.2500 ;
	    RECT 1172.7001 533.1000 1174.5000 533.2500 ;
	    RECT 1199.1000 533.1000 1200.9000 533.2500 ;
	    RECT 1213.5000 534.7500 1215.3000 534.9000 ;
	    RECT 1251.9000 534.7500 1253.7001 534.9000 ;
	    RECT 1213.5000 533.2500 1253.7001 534.7500 ;
	    RECT 1213.5000 533.1000 1215.3000 533.2500 ;
	    RECT 1251.9000 533.1000 1253.7001 533.2500 ;
	    RECT 1314.3000 534.7500 1316.1000 534.9000 ;
	    RECT 1331.1000 534.7500 1332.9000 534.9000 ;
	    RECT 1335.9000 534.7500 1337.7001 534.9000 ;
	    RECT 1314.3000 533.2500 1337.7001 534.7500 ;
	    RECT 1314.3000 533.1000 1316.1000 533.2500 ;
	    RECT 1331.1000 533.1000 1332.9000 533.2500 ;
	    RECT 1335.9000 533.1000 1337.7001 533.2500 ;
	    RECT 1350.3000 534.7500 1352.1000 534.9000 ;
	    RECT 1371.9000 534.7500 1373.7001 534.9000 ;
	    RECT 1350.3000 533.2500 1373.7001 534.7500 ;
	    RECT 1350.3000 533.1000 1352.1000 533.2500 ;
	    RECT 1371.9000 533.1000 1373.7001 533.2500 ;
	    RECT 1496.7001 534.7500 1498.5000 534.9000 ;
	    RECT 1525.5000 534.7500 1527.3000 534.9000 ;
	    RECT 1496.7001 533.2500 1527.3000 534.7500 ;
	    RECT 1496.7001 533.1000 1498.5000 533.2500 ;
	    RECT 1525.5000 533.1000 1527.3000 533.2500 ;
	    RECT 133.5000 528.7500 135.3000 528.9000 ;
	    RECT 159.9000 528.7500 161.7000 528.9000 ;
	    RECT 301.5000 528.7500 303.3000 528.9000 ;
	    RECT 133.5000 527.2500 303.3000 528.7500 ;
	    RECT 133.5000 527.1000 135.3000 527.2500 ;
	    RECT 159.9000 527.1000 161.7000 527.2500 ;
	    RECT 301.5000 527.1000 303.3000 527.2500 ;
	    RECT 339.9000 528.7500 341.7000 528.9000 ;
	    RECT 349.5000 528.7500 351.3000 528.9000 ;
	    RECT 339.9000 527.2500 351.3000 528.7500 ;
	    RECT 339.9000 527.1000 341.7000 527.2500 ;
	    RECT 349.5000 527.1000 351.3000 527.2500 ;
	    RECT 781.5000 528.7500 783.3000 528.9000 ;
	    RECT 817.5000 528.7500 819.3000 528.9000 ;
	    RECT 781.5000 527.2500 819.3000 528.7500 ;
	    RECT 781.5000 527.1000 783.3000 527.2500 ;
	    RECT 817.5000 527.1000 819.3000 527.2500 ;
	    RECT 851.1000 528.7500 852.9000 528.9000 ;
	    RECT 911.1000 528.7500 912.9000 528.9000 ;
	    RECT 851.1000 527.2500 912.9000 528.7500 ;
	    RECT 851.1000 527.1000 852.9000 527.2500 ;
	    RECT 911.1000 527.1000 912.9000 527.2500 ;
	    RECT 973.5000 528.7500 975.3000 528.9000 ;
	    RECT 985.5000 528.7500 987.3000 528.9000 ;
	    RECT 973.5000 527.2500 987.3000 528.7500 ;
	    RECT 973.5000 527.1000 975.3000 527.2500 ;
	    RECT 985.5000 527.1000 987.3000 527.2500 ;
	    RECT 1021.5000 528.7500 1023.3000 528.9000 ;
	    RECT 1045.5000 528.7500 1047.3000 528.9000 ;
	    RECT 1021.5000 527.2500 1047.3000 528.7500 ;
	    RECT 1021.5000 527.1000 1023.3000 527.2500 ;
	    RECT 1045.5000 527.1000 1047.3000 527.2500 ;
	    RECT 1136.7001 528.7500 1138.5000 528.9000 ;
	    RECT 1146.3000 528.7500 1148.1000 528.9000 ;
	    RECT 1136.7001 527.2500 1148.1000 528.7500 ;
	    RECT 1136.7001 527.1000 1138.5000 527.2500 ;
	    RECT 1146.3000 527.1000 1148.1000 527.2500 ;
	    RECT 1316.7001 528.7500 1318.5000 528.9000 ;
	    RECT 1350.3000 528.7500 1352.1000 528.9000 ;
	    RECT 1316.7001 527.2500 1352.1000 528.7500 ;
	    RECT 1316.7001 527.1000 1318.5000 527.2500 ;
	    RECT 1350.3000 527.1000 1352.1000 527.2500 ;
	    RECT 1367.1000 528.7500 1368.9000 528.9000 ;
	    RECT 1379.1000 528.7500 1380.9000 528.9000 ;
	    RECT 1367.1000 527.2500 1380.9000 528.7500 ;
	    RECT 1367.1000 527.1000 1368.9000 527.2500 ;
	    RECT 1379.1000 527.1000 1380.9000 527.2500 ;
	    RECT 1491.9000 528.7500 1493.7001 528.9000 ;
	    RECT 1508.7001 528.7500 1510.5000 528.9000 ;
	    RECT 1491.9000 527.2500 1510.5000 528.7500 ;
	    RECT 1491.9000 527.1000 1493.7001 527.2500 ;
	    RECT 1508.7001 527.1000 1510.5000 527.2500 ;
	    RECT 457.5000 522.7500 459.3000 522.9000 ;
	    RECT 531.9000 522.7500 533.7000 522.9000 ;
	    RECT 457.5000 521.2500 533.7000 522.7500 ;
	    RECT 457.5000 521.1000 459.3000 521.2500 ;
	    RECT 531.9000 521.1000 533.7000 521.2500 ;
	    RECT 536.7000 522.7500 538.5000 522.9000 ;
	    RECT 649.5000 522.7500 651.3000 522.9000 ;
	    RECT 536.7000 521.2500 651.3000 522.7500 ;
	    RECT 536.7000 521.1000 538.5000 521.2500 ;
	    RECT 649.5000 521.1000 651.3000 521.2500 ;
	    RECT 786.3000 522.7500 788.1000 522.9000 ;
	    RECT 839.1000 522.7500 840.9000 522.9000 ;
	    RECT 786.3000 521.2500 840.9000 522.7500 ;
	    RECT 786.3000 521.1000 788.1000 521.2500 ;
	    RECT 839.1000 521.1000 840.9000 521.2500 ;
	    RECT 855.9000 522.7500 857.7000 522.9000 ;
	    RECT 903.9000 522.7500 905.7000 522.9000 ;
	    RECT 855.9000 521.2500 905.7000 522.7500 ;
	    RECT 855.9000 521.1000 857.7000 521.2500 ;
	    RECT 903.9000 521.1000 905.7000 521.2500 ;
	    RECT 1043.1000 522.7500 1044.9000 522.9000 ;
	    RECT 1062.3000 522.7500 1064.1000 522.9000 ;
	    RECT 1043.1000 521.2500 1064.1000 522.7500 ;
	    RECT 1043.1000 521.1000 1044.9000 521.2500 ;
	    RECT 1062.3000 521.1000 1064.1000 521.2500 ;
	    RECT 1141.5000 522.7500 1143.3000 522.9000 ;
	    RECT 1170.3000 522.7500 1172.1000 522.9000 ;
	    RECT 1141.5000 521.2500 1172.1000 522.7500 ;
	    RECT 1141.5000 521.1000 1143.3000 521.2500 ;
	    RECT 1170.3000 521.1000 1172.1000 521.2500 ;
	    RECT 1227.9000 522.7500 1229.7001 522.9000 ;
	    RECT 1242.3000 522.7500 1244.1000 522.9000 ;
	    RECT 1268.7001 522.7500 1270.5000 522.9000 ;
	    RECT 1227.9000 521.2500 1270.5000 522.7500 ;
	    RECT 1227.9000 521.1000 1229.7001 521.2500 ;
	    RECT 1242.3000 521.1000 1244.1000 521.2500 ;
	    RECT 1268.7001 521.1000 1270.5000 521.2500 ;
	    RECT 1302.3000 522.7500 1304.1000 522.9000 ;
	    RECT 1319.1000 522.7500 1320.9000 522.9000 ;
	    RECT 1302.3000 521.2500 1320.9000 522.7500 ;
	    RECT 1302.3000 521.1000 1304.1000 521.2500 ;
	    RECT 1319.1000 521.1000 1320.9000 521.2500 ;
	    RECT 1434.3000 522.7500 1436.1000 522.9000 ;
	    RECT 1460.7001 522.7500 1462.5000 522.9000 ;
	    RECT 1434.3000 521.2500 1462.5000 522.7500 ;
	    RECT 1434.3000 521.1000 1436.1000 521.2500 ;
	    RECT 1460.7001 521.1000 1462.5000 521.2500 ;
	    RECT 1499.1000 522.7500 1500.9000 522.9000 ;
	    RECT 1503.9000 522.7500 1505.7001 522.9000 ;
	    RECT 1499.1000 521.2500 1505.7001 522.7500 ;
	    RECT 1499.1000 521.1000 1500.9000 521.2500 ;
	    RECT 1503.9000 521.1000 1505.7001 521.2500 ;
	    RECT 1542.3000 522.7500 1544.1000 522.9000 ;
	    RECT 1563.9000 522.7500 1565.7001 522.9000 ;
	    RECT 1542.3000 521.2500 1565.7001 522.7500 ;
	    RECT 1542.3000 521.1000 1544.1000 521.2500 ;
	    RECT 1563.9000 521.1000 1565.7001 521.2500 ;
	    RECT 306.3000 516.7500 308.1000 516.9000 ;
	    RECT 349.5000 516.7500 351.3000 516.9000 ;
	    RECT 306.3000 515.2500 351.3000 516.7500 ;
	    RECT 306.3000 515.1000 308.1000 515.2500 ;
	    RECT 349.5000 515.1000 351.3000 515.2500 ;
	    RECT 647.1000 516.7500 648.9000 516.9000 ;
	    RECT 810.3000 516.7500 812.1000 516.9000 ;
	    RECT 647.1000 515.2500 812.1000 516.7500 ;
	    RECT 647.1000 515.1000 648.9000 515.2500 ;
	    RECT 810.3000 515.1000 812.1000 515.2500 ;
	    RECT 817.5000 516.7500 819.3000 516.9000 ;
	    RECT 843.9000 516.7500 845.7000 516.9000 ;
	    RECT 817.5000 515.2500 845.7000 516.7500 ;
	    RECT 817.5000 515.1000 819.3000 515.2500 ;
	    RECT 843.9000 515.1000 845.7000 515.2500 ;
	    RECT 1033.5000 516.7500 1035.3000 516.9000 ;
	    RECT 1127.1000 516.7500 1128.9000 516.9000 ;
	    RECT 1297.5000 516.7500 1299.3000 516.9000 ;
	    RECT 1033.5000 515.2500 1299.3000 516.7500 ;
	    RECT 1033.5000 515.1000 1035.3000 515.2500 ;
	    RECT 1127.1000 515.1000 1128.9000 515.2500 ;
	    RECT 1297.5000 515.1000 1299.3000 515.2500 ;
	    RECT 1314.3000 516.7500 1316.1000 516.9000 ;
	    RECT 1323.9000 516.7500 1325.7001 516.9000 ;
	    RECT 1314.3000 515.2500 1325.7001 516.7500 ;
	    RECT 1314.3000 515.1000 1316.1000 515.2500 ;
	    RECT 1323.9000 515.1000 1325.7001 515.2500 ;
	    RECT 1345.5000 516.7500 1347.3000 516.9000 ;
	    RECT 1374.3000 516.7500 1376.1000 516.9000 ;
	    RECT 1345.5000 515.2500 1376.1000 516.7500 ;
	    RECT 1345.5000 515.1000 1347.3000 515.2500 ;
	    RECT 1374.3000 515.1000 1376.1000 515.2500 ;
	    RECT 131.1000 510.7500 132.9000 510.9000 ;
	    RECT 174.3000 510.7500 176.1000 510.9000 ;
	    RECT 131.1000 509.2500 176.1000 510.7500 ;
	    RECT 131.1000 509.1000 132.9000 509.2500 ;
	    RECT 174.3000 509.1000 176.1000 509.2500 ;
	    RECT 445.5000 510.7500 447.3000 510.9000 ;
	    RECT 495.9000 510.7500 497.7000 510.9000 ;
	    RECT 445.5000 509.2500 497.7000 510.7500 ;
	    RECT 445.5000 509.1000 447.3000 509.2500 ;
	    RECT 495.9000 509.1000 497.7000 509.2500 ;
	    RECT 539.1000 510.7500 540.9000 510.9000 ;
	    RECT 615.9000 510.7500 617.7000 510.9000 ;
	    RECT 539.1000 509.2500 617.7000 510.7500 ;
	    RECT 539.1000 509.1000 540.9000 509.2500 ;
	    RECT 615.9000 509.1000 617.7000 509.2500 ;
	    RECT 743.1000 510.7500 744.9000 510.9000 ;
	    RECT 750.3000 510.7500 752.1000 510.9000 ;
	    RECT 743.1000 509.2500 752.1000 510.7500 ;
	    RECT 743.1000 509.1000 744.9000 509.2500 ;
	    RECT 750.3000 509.1000 752.1000 509.2500 ;
	    RECT 812.7000 510.7500 814.5000 510.9000 ;
	    RECT 824.7000 510.7500 826.5000 510.9000 ;
	    RECT 812.7000 509.2500 826.5000 510.7500 ;
	    RECT 812.7000 509.1000 814.5000 509.2500 ;
	    RECT 824.7000 509.1000 826.5000 509.2500 ;
	    RECT 1069.5000 510.7500 1071.3000 510.9000 ;
	    RECT 1107.9000 510.7500 1109.7001 510.9000 ;
	    RECT 1069.5000 509.2500 1109.7001 510.7500 ;
	    RECT 1069.5000 509.1000 1071.3000 509.2500 ;
	    RECT 1107.9000 509.1000 1109.7001 509.2500 ;
	    RECT 1134.3000 510.7500 1136.1000 510.9000 ;
	    RECT 1211.1000 510.7500 1212.9000 510.9000 ;
	    RECT 1134.3000 509.2500 1212.9000 510.7500 ;
	    RECT 1134.3000 509.1000 1136.1000 509.2500 ;
	    RECT 1211.1000 509.1000 1212.9000 509.2500 ;
	    RECT 1220.7001 510.7500 1222.5000 510.9000 ;
	    RECT 1256.7001 510.7500 1258.5000 510.9000 ;
	    RECT 1220.7001 509.2500 1258.5000 510.7500 ;
	    RECT 1220.7001 509.1000 1222.5000 509.2500 ;
	    RECT 1256.7001 509.1000 1258.5000 509.2500 ;
	    RECT 1388.7001 510.7500 1390.5000 510.9000 ;
	    RECT 1403.1000 510.7500 1404.9000 510.9000 ;
	    RECT 1388.7001 509.2500 1404.9000 510.7500 ;
	    RECT 1388.7001 509.1000 1390.5000 509.2500 ;
	    RECT 1403.1000 509.1000 1404.9000 509.2500 ;
	    RECT 1515.9000 510.7500 1517.7001 510.9000 ;
	    RECT 1561.5000 510.7500 1563.3000 510.9000 ;
	    RECT 1515.9000 509.2500 1563.3000 510.7500 ;
	    RECT 1515.9000 509.1000 1517.7001 509.2500 ;
	    RECT 1561.5000 509.1000 1563.3000 509.2500 ;
	    RECT 49.5000 504.7500 51.3000 504.9000 ;
	    RECT 145.5000 504.7500 147.3000 504.9000 ;
	    RECT 49.5000 503.2500 147.3000 504.7500 ;
	    RECT 49.5000 503.1000 51.3000 503.2500 ;
	    RECT 145.5000 503.1000 147.3000 503.2500 ;
	    RECT 193.5000 504.7500 195.3000 504.9000 ;
	    RECT 215.1000 504.7500 216.9000 504.9000 ;
	    RECT 222.3000 504.7500 224.1000 504.9000 ;
	    RECT 193.5000 503.2500 224.1000 504.7500 ;
	    RECT 193.5000 503.1000 195.3000 503.2500 ;
	    RECT 215.1000 503.1000 216.9000 503.2500 ;
	    RECT 222.3000 503.1000 224.1000 503.2500 ;
	    RECT 282.3000 504.7500 284.1000 504.9000 ;
	    RECT 315.9000 504.7500 317.7000 504.9000 ;
	    RECT 282.3000 503.2500 317.7000 504.7500 ;
	    RECT 282.3000 503.1000 284.1000 503.2500 ;
	    RECT 315.9000 503.1000 317.7000 503.2500 ;
	    RECT 495.9000 504.7500 497.7000 504.9000 ;
	    RECT 536.7000 504.7500 538.5000 504.9000 ;
	    RECT 495.9000 503.2500 538.5000 504.7500 ;
	    RECT 495.9000 503.1000 497.7000 503.2500 ;
	    RECT 536.7000 503.1000 538.5000 503.2500 ;
	    RECT 635.1000 504.7500 636.9000 504.9000 ;
	    RECT 714.3000 504.7500 716.1000 504.9000 ;
	    RECT 635.1000 503.2500 716.1000 504.7500 ;
	    RECT 635.1000 503.1000 636.9000 503.2500 ;
	    RECT 714.3000 503.1000 716.1000 503.2500 ;
	    RECT 721.5000 504.7500 723.3000 504.9000 ;
	    RECT 803.1000 504.7500 804.9000 504.9000 ;
	    RECT 721.5000 503.2500 804.9000 504.7500 ;
	    RECT 721.5000 503.1000 723.3000 503.2500 ;
	    RECT 803.1000 503.1000 804.9000 503.2500 ;
	    RECT 815.1000 504.7500 816.9000 504.9000 ;
	    RECT 819.9000 504.7500 821.7000 504.9000 ;
	    RECT 815.1000 503.2500 821.7000 504.7500 ;
	    RECT 815.1000 503.1000 816.9000 503.2500 ;
	    RECT 819.9000 503.1000 821.7000 503.2500 ;
	    RECT 1045.5000 504.7500 1047.3000 504.9000 ;
	    RECT 1064.7001 504.7500 1066.5000 504.9000 ;
	    RECT 1045.5000 503.2500 1066.5000 504.7500 ;
	    RECT 1045.5000 503.1000 1047.3000 503.2500 ;
	    RECT 1064.7001 503.1000 1066.5000 503.2500 ;
	    RECT 1076.7001 504.7500 1078.5000 504.9000 ;
	    RECT 1117.5000 504.7500 1119.3000 504.9000 ;
	    RECT 1076.7001 503.2500 1119.3000 504.7500 ;
	    RECT 1076.7001 503.1000 1078.5000 503.2500 ;
	    RECT 1117.5000 503.1000 1119.3000 503.2500 ;
	    RECT 1131.9000 504.7500 1133.7001 504.9000 ;
	    RECT 1160.7001 504.7500 1162.5000 504.9000 ;
	    RECT 1131.9000 503.2500 1162.5000 504.7500 ;
	    RECT 1131.9000 503.1000 1133.7001 503.2500 ;
	    RECT 1160.7001 503.1000 1162.5000 503.2500 ;
	    RECT 1189.5000 504.7500 1191.3000 504.9000 ;
	    RECT 1199.1000 504.7500 1200.9000 504.9000 ;
	    RECT 1189.5000 503.2500 1200.9000 504.7500 ;
	    RECT 1189.5000 503.1000 1191.3000 503.2500 ;
	    RECT 1199.1000 503.1000 1200.9000 503.2500 ;
	    RECT 1203.9000 504.7500 1205.7001 504.9000 ;
	    RECT 1225.5000 504.7500 1227.3000 504.9000 ;
	    RECT 1261.5000 504.7500 1263.3000 504.9000 ;
	    RECT 1203.9000 503.2500 1263.3000 504.7500 ;
	    RECT 1203.9000 503.1000 1205.7001 503.2500 ;
	    RECT 1225.5000 503.1000 1227.3000 503.2500 ;
	    RECT 1261.5000 503.1000 1263.3000 503.2500 ;
	    RECT 1319.1000 504.7500 1320.9000 504.9000 ;
	    RECT 1355.1000 504.7500 1356.9000 504.9000 ;
	    RECT 1319.1000 503.2500 1356.9000 504.7500 ;
	    RECT 1319.1000 503.1000 1320.9000 503.2500 ;
	    RECT 1355.1000 503.1000 1356.9000 503.2500 ;
	    RECT 135.9000 498.7500 137.7000 498.9000 ;
	    RECT 162.3000 498.7500 164.1000 498.9000 ;
	    RECT 176.7000 498.7500 178.5000 498.9000 ;
	    RECT 135.9000 497.2500 178.5000 498.7500 ;
	    RECT 135.9000 497.1000 137.7000 497.2500 ;
	    RECT 162.3000 497.1000 164.1000 497.2500 ;
	    RECT 176.7000 497.1000 178.5000 497.2500 ;
	    RECT 186.3000 498.7500 188.1000 498.9000 ;
	    RECT 251.1000 498.7500 252.9000 498.9000 ;
	    RECT 186.3000 497.2500 252.9000 498.7500 ;
	    RECT 186.3000 497.1000 188.1000 497.2500 ;
	    RECT 251.1000 497.1000 252.9000 497.2500 ;
	    RECT 263.1000 498.7500 264.9000 498.9000 ;
	    RECT 270.3000 498.7500 272.1000 498.9000 ;
	    RECT 263.1000 497.2500 272.1000 498.7500 ;
	    RECT 263.1000 497.1000 264.9000 497.2500 ;
	    RECT 270.3000 497.1000 272.1000 497.2500 ;
	    RECT 299.1000 498.7500 300.9000 498.9000 ;
	    RECT 308.7000 498.7500 310.5000 498.9000 ;
	    RECT 299.1000 497.2500 310.5000 498.7500 ;
	    RECT 299.1000 497.1000 300.9000 497.2500 ;
	    RECT 308.7000 497.1000 310.5000 497.2500 ;
	    RECT 330.3000 498.7500 332.1000 498.9000 ;
	    RECT 347.1000 498.7500 348.9000 498.9000 ;
	    RECT 330.3000 497.2500 348.9000 498.7500 ;
	    RECT 330.3000 497.1000 332.1000 497.2500 ;
	    RECT 347.1000 497.1000 348.9000 497.2500 ;
	    RECT 450.3000 498.7500 452.1000 498.9000 ;
	    RECT 500.7000 498.7500 502.5000 498.9000 ;
	    RECT 450.3000 497.2500 502.5000 498.7500 ;
	    RECT 450.3000 497.1000 452.1000 497.2500 ;
	    RECT 500.7000 497.1000 502.5000 497.2500 ;
	    RECT 611.1000 498.7500 612.9000 498.9000 ;
	    RECT 635.1000 498.7500 636.9000 498.9000 ;
	    RECT 611.1000 497.2500 636.9000 498.7500 ;
	    RECT 611.1000 497.1000 612.9000 497.2500 ;
	    RECT 635.1000 497.1000 636.9000 497.2500 ;
	    RECT 1148.7001 498.7500 1150.5000 498.9000 ;
	    RECT 1182.3000 498.7500 1184.1000 498.9000 ;
	    RECT 1148.7001 497.2500 1184.1000 498.7500 ;
	    RECT 1148.7001 497.1000 1150.5000 497.2500 ;
	    RECT 1182.3000 497.1000 1184.1000 497.2500 ;
	    RECT 1223.1000 498.7500 1224.9000 498.9000 ;
	    RECT 1254.3000 498.7500 1256.1000 498.9000 ;
	    RECT 1223.1000 497.2500 1256.1000 498.7500 ;
	    RECT 1223.1000 497.1000 1224.9000 497.2500 ;
	    RECT 1254.3000 497.1000 1256.1000 497.2500 ;
	    RECT 1283.1000 498.7500 1284.9000 498.9000 ;
	    RECT 1292.7001 498.7500 1294.5000 498.9000 ;
	    RECT 1283.1000 497.2500 1294.5000 498.7500 ;
	    RECT 1283.1000 497.1000 1284.9000 497.2500 ;
	    RECT 1292.7001 497.1000 1294.5000 497.2500 ;
	    RECT 1419.9000 498.7500 1421.7001 498.9000 ;
	    RECT 1443.9000 498.7500 1445.7001 498.9000 ;
	    RECT 1453.5000 498.7500 1455.3000 498.9000 ;
	    RECT 1419.9000 497.2500 1455.3000 498.7500 ;
	    RECT 1419.9000 497.1000 1421.7001 497.2500 ;
	    RECT 1443.9000 497.1000 1445.7001 497.2500 ;
	    RECT 1453.5000 497.1000 1455.3000 497.2500 ;
	    RECT 1482.3000 498.7500 1484.1000 498.9000 ;
	    RECT 1487.1000 498.7500 1488.9000 498.9000 ;
	    RECT 1482.3000 497.2500 1488.9000 498.7500 ;
	    RECT 1482.3000 497.1000 1484.1000 497.2500 ;
	    RECT 1487.1000 497.1000 1488.9000 497.2500 ;
	    RECT 42.3000 492.7500 44.1000 492.9000 ;
	    RECT 183.9000 492.7500 185.7000 492.9000 ;
	    RECT 42.3000 491.2500 185.7000 492.7500 ;
	    RECT 42.3000 491.1000 44.1000 491.2500 ;
	    RECT 183.9000 491.1000 185.7000 491.2500 ;
	    RECT 229.5000 492.7500 231.3000 492.9000 ;
	    RECT 272.7000 492.7500 274.5000 492.9000 ;
	    RECT 229.5000 491.2500 274.5000 492.7500 ;
	    RECT 229.5000 491.1000 231.3000 491.2500 ;
	    RECT 272.7000 491.1000 274.5000 491.2500 ;
	    RECT 289.5000 492.7500 291.3000 492.9000 ;
	    RECT 299.1000 492.7500 300.9000 492.9000 ;
	    RECT 289.5000 491.2500 300.9000 492.7500 ;
	    RECT 289.5000 491.1000 291.3000 491.2500 ;
	    RECT 299.1000 491.1000 300.9000 491.2500 ;
	    RECT 332.7000 492.7500 334.5000 492.9000 ;
	    RECT 378.3000 492.7500 380.1000 492.9000 ;
	    RECT 332.7000 491.2500 380.1000 492.7500 ;
	    RECT 332.7000 491.1000 334.5000 491.2500 ;
	    RECT 378.3000 491.1000 380.1000 491.2500 ;
	    RECT 467.1000 492.7500 468.9000 492.9000 ;
	    RECT 510.3000 492.7500 512.1000 492.9000 ;
	    RECT 467.1000 491.2500 512.1000 492.7500 ;
	    RECT 467.1000 491.1000 468.9000 491.2500 ;
	    RECT 510.3000 491.1000 512.1000 491.2500 ;
	    RECT 515.1000 492.7500 516.9000 492.9000 ;
	    RECT 577.5000 492.7500 579.3000 492.9000 ;
	    RECT 515.1000 491.2500 579.3000 492.7500 ;
	    RECT 515.1000 491.1000 516.9000 491.2500 ;
	    RECT 577.5000 491.1000 579.3000 491.2500 ;
	    RECT 582.3000 492.7500 584.1000 492.9000 ;
	    RECT 637.5000 492.7500 639.3000 492.9000 ;
	    RECT 582.3000 491.2500 639.3000 492.7500 ;
	    RECT 582.3000 491.1000 584.1000 491.2500 ;
	    RECT 637.5000 491.1000 639.3000 491.2500 ;
	    RECT 714.3000 492.7500 716.1000 492.9000 ;
	    RECT 959.1000 492.7500 960.9000 492.9000 ;
	    RECT 714.3000 491.2500 960.9000 492.7500 ;
	    RECT 714.3000 491.1000 716.1000 491.2500 ;
	    RECT 959.1000 491.1000 960.9000 491.2500 ;
	    RECT 978.3000 492.7500 980.1000 492.9000 ;
	    RECT 1050.3000 492.7500 1052.1000 492.9000 ;
	    RECT 978.3000 491.2500 1052.1000 492.7500 ;
	    RECT 978.3000 491.1000 980.1000 491.2500 ;
	    RECT 1050.3000 491.1000 1052.1000 491.2500 ;
	    RECT 1184.7001 492.7500 1186.5000 492.9000 ;
	    RECT 1191.9000 492.7500 1193.7001 492.9000 ;
	    RECT 1184.7001 491.2500 1193.7001 492.7500 ;
	    RECT 1184.7001 491.1000 1186.5000 491.2500 ;
	    RECT 1191.9000 491.1000 1193.7001 491.2500 ;
	    RECT 1251.9000 492.7500 1253.7001 492.9000 ;
	    RECT 1319.1000 492.7500 1320.9000 492.9000 ;
	    RECT 1350.3000 492.7500 1352.1000 492.9000 ;
	    RECT 1251.9000 491.2500 1352.1000 492.7500 ;
	    RECT 1251.9000 491.1000 1253.7001 491.2500 ;
	    RECT 1319.1000 491.1000 1320.9000 491.2500 ;
	    RECT 1350.3000 491.1000 1352.1000 491.2500 ;
	    RECT 1453.5000 492.7500 1455.3000 492.9000 ;
	    RECT 1467.9000 492.7500 1469.7001 492.9000 ;
	    RECT 1453.5000 491.2500 1469.7001 492.7500 ;
	    RECT 1453.5000 491.1000 1455.3000 491.2500 ;
	    RECT 1467.9000 491.1000 1469.7001 491.2500 ;
	    RECT 116.7000 486.7500 118.5000 486.9000 ;
	    RECT 171.9000 486.7500 173.7000 486.9000 ;
	    RECT 116.7000 485.2500 173.7000 486.7500 ;
	    RECT 116.7000 485.1000 118.5000 485.2500 ;
	    RECT 171.9000 485.1000 173.7000 485.2500 ;
	    RECT 219.9000 486.7500 221.7000 486.9000 ;
	    RECT 260.7000 486.7500 262.5000 486.9000 ;
	    RECT 219.9000 485.2500 262.5000 486.7500 ;
	    RECT 219.9000 485.1000 221.7000 485.2500 ;
	    RECT 260.7000 485.1000 262.5000 485.2500 ;
	    RECT 303.9000 486.7500 305.7000 486.9000 ;
	    RECT 342.3000 486.7500 344.1000 486.9000 ;
	    RECT 303.9000 485.2500 344.1000 486.7500 ;
	    RECT 303.9000 485.1000 305.7000 485.2500 ;
	    RECT 342.3000 485.1000 344.1000 485.2500 ;
	    RECT 404.7000 486.7500 406.5000 486.9000 ;
	    RECT 431.1000 486.7500 432.9000 486.9000 ;
	    RECT 404.7000 485.2500 432.9000 486.7500 ;
	    RECT 404.7000 485.1000 406.5000 485.2500 ;
	    RECT 431.1000 485.1000 432.9000 485.2500 ;
	    RECT 699.9000 486.7500 701.7000 486.9000 ;
	    RECT 872.7000 486.7500 874.5000 486.9000 ;
	    RECT 699.9000 485.2500 874.5000 486.7500 ;
	    RECT 699.9000 485.1000 701.7000 485.2500 ;
	    RECT 872.7000 485.1000 874.5000 485.2500 ;
	    RECT 1021.5000 486.7500 1023.3000 486.9000 ;
	    RECT 1047.9000 486.7500 1049.7001 486.9000 ;
	    RECT 1021.5000 485.2500 1049.7001 486.7500 ;
	    RECT 1021.5000 485.1000 1023.3000 485.2500 ;
	    RECT 1047.9000 485.1000 1049.7001 485.2500 ;
	    RECT 1074.3000 486.7500 1076.1000 486.9000 ;
	    RECT 1086.3000 486.7500 1088.1000 486.9000 ;
	    RECT 1110.3000 486.7500 1112.1000 486.9000 ;
	    RECT 1074.3000 485.2500 1112.1000 486.7500 ;
	    RECT 1074.3000 485.1000 1076.1000 485.2500 ;
	    RECT 1086.3000 485.1000 1088.1000 485.2500 ;
	    RECT 1110.3000 485.1000 1112.1000 485.2500 ;
	    RECT 1182.3000 486.7500 1184.1000 486.9000 ;
	    RECT 1194.3000 486.7500 1196.1000 486.9000 ;
	    RECT 1182.3000 485.2500 1196.1000 486.7500 ;
	    RECT 1182.3000 485.1000 1184.1000 485.2500 ;
	    RECT 1194.3000 485.1000 1196.1000 485.2500 ;
	    RECT 1285.5000 486.7500 1287.3000 486.9000 ;
	    RECT 1311.9000 486.7500 1313.7001 486.9000 ;
	    RECT 1338.3000 486.7500 1340.1000 486.9000 ;
	    RECT 1285.5000 485.2500 1340.1000 486.7500 ;
	    RECT 1285.5000 485.1000 1287.3000 485.2500 ;
	    RECT 1311.9000 485.1000 1313.7001 485.2500 ;
	    RECT 1338.3000 485.1000 1340.1000 485.2500 ;
	    RECT 318.3000 480.7500 320.1000 480.9000 ;
	    RECT 330.3000 480.7500 332.1000 480.9000 ;
	    RECT 318.3000 479.2500 332.1000 480.7500 ;
	    RECT 318.3000 479.1000 320.1000 479.2500 ;
	    RECT 330.3000 479.1000 332.1000 479.2500 ;
	    RECT 339.9000 480.7500 341.7000 480.9000 ;
	    RECT 469.5000 480.7500 471.3000 480.9000 ;
	    RECT 339.9000 479.2500 471.3000 480.7500 ;
	    RECT 339.9000 479.1000 341.7000 479.2500 ;
	    RECT 469.5000 479.1000 471.3000 479.2500 ;
	    RECT 567.9000 480.7500 569.7000 480.9000 ;
	    RECT 613.5000 480.7500 615.3000 480.9000 ;
	    RECT 567.9000 479.2500 615.3000 480.7500 ;
	    RECT 567.9000 479.1000 569.7000 479.2500 ;
	    RECT 613.5000 479.1000 615.3000 479.2500 ;
	    RECT 822.3000 480.7500 824.1000 480.9000 ;
	    RECT 831.9000 480.7500 833.7000 480.9000 ;
	    RECT 822.3000 479.2500 833.7000 480.7500 ;
	    RECT 822.3000 479.1000 824.1000 479.2500 ;
	    RECT 831.9000 479.1000 833.7000 479.2500 ;
	    RECT 839.1000 480.7500 840.9000 480.9000 ;
	    RECT 889.5000 480.7500 891.3000 480.9000 ;
	    RECT 839.1000 479.2500 891.3000 480.7500 ;
	    RECT 839.1000 479.1000 840.9000 479.2500 ;
	    RECT 889.5000 479.1000 891.3000 479.2500 ;
	    RECT 1026.3000 480.7500 1028.1000 480.9000 ;
	    RECT 1031.1000 480.7500 1032.9000 480.9000 ;
	    RECT 1026.3000 479.2500 1032.9000 480.7500 ;
	    RECT 1026.3000 479.1000 1028.1000 479.2500 ;
	    RECT 1031.1000 479.1000 1032.9000 479.2500 ;
	    RECT 1035.9000 480.7500 1037.7001 480.9000 ;
	    RECT 1040.7001 480.7500 1042.5000 480.9000 ;
	    RECT 1035.9000 479.2500 1042.5000 480.7500 ;
	    RECT 1035.9000 479.1000 1037.7001 479.2500 ;
	    RECT 1040.7001 479.1000 1042.5000 479.2500 ;
	    RECT 1045.5000 480.7500 1047.3000 480.9000 ;
	    RECT 1098.3000 480.7500 1100.1000 480.9000 ;
	    RECT 1045.5000 479.2500 1100.1000 480.7500 ;
	    RECT 1045.5000 479.1000 1047.3000 479.2500 ;
	    RECT 1098.3000 479.1000 1100.1000 479.2500 ;
	    RECT 1187.1000 480.7500 1188.9000 480.9000 ;
	    RECT 1203.9000 480.7500 1205.7001 480.9000 ;
	    RECT 1244.7001 480.7500 1246.5000 480.9000 ;
	    RECT 1187.1000 479.2500 1246.5000 480.7500 ;
	    RECT 1187.1000 479.1000 1188.9000 479.2500 ;
	    RECT 1203.9000 479.1000 1205.7001 479.2500 ;
	    RECT 1244.7001 479.1000 1246.5000 479.2500 ;
	    RECT 1335.9000 480.7500 1337.7001 480.9000 ;
	    RECT 1352.7001 480.7500 1354.5000 480.9000 ;
	    RECT 1379.1000 480.7500 1380.9000 480.9000 ;
	    RECT 1335.9000 479.2500 1380.9000 480.7500 ;
	    RECT 1335.9000 479.1000 1337.7001 479.2500 ;
	    RECT 1352.7001 479.1000 1354.5000 479.2500 ;
	    RECT 1379.1000 479.1000 1380.9000 479.2500 ;
	    RECT 131.1000 474.7500 132.9000 474.9000 ;
	    RECT 219.9000 474.7500 221.7000 474.9000 ;
	    RECT 131.1000 473.2500 221.7000 474.7500 ;
	    RECT 131.1000 473.1000 132.9000 473.2500 ;
	    RECT 219.9000 473.1000 221.7000 473.2500 ;
	    RECT 315.9000 474.7500 317.7000 474.9000 ;
	    RECT 366.3000 474.7500 368.1000 474.9000 ;
	    RECT 315.9000 473.2500 368.1000 474.7500 ;
	    RECT 315.9000 473.1000 317.7000 473.2500 ;
	    RECT 366.3000 473.1000 368.1000 473.2500 ;
	    RECT 603.9000 474.7500 605.7000 474.9000 ;
	    RECT 642.3000 474.7500 644.1000 474.9000 ;
	    RECT 603.9000 473.2500 644.1000 474.7500 ;
	    RECT 603.9000 473.1000 605.7000 473.2500 ;
	    RECT 642.3000 473.1000 644.1000 473.2500 ;
	    RECT 762.3000 474.7500 764.1000 474.9000 ;
	    RECT 810.3000 474.7500 812.1000 474.9000 ;
	    RECT 762.3000 473.2500 812.1000 474.7500 ;
	    RECT 762.3000 473.1000 764.1000 473.2500 ;
	    RECT 810.3000 473.1000 812.1000 473.2500 ;
	    RECT 843.9000 474.7500 845.7000 474.9000 ;
	    RECT 925.5000 474.7500 927.3000 474.9000 ;
	    RECT 843.9000 473.2500 927.3000 474.7500 ;
	    RECT 843.9000 473.1000 845.7000 473.2500 ;
	    RECT 925.5000 473.1000 927.3000 473.2500 ;
	    RECT 1019.1000 474.7500 1020.9000 474.9000 ;
	    RECT 1026.3000 474.7500 1028.1000 474.9000 ;
	    RECT 1019.1000 473.2500 1028.1000 474.7500 ;
	    RECT 1019.1000 473.1000 1020.9000 473.2500 ;
	    RECT 1026.3000 473.1000 1028.1000 473.2500 ;
	    RECT 1031.1000 474.7500 1032.9000 474.9000 ;
	    RECT 1035.9000 474.7500 1037.7001 474.9000 ;
	    RECT 1031.1000 473.2500 1037.7001 474.7500 ;
	    RECT 1031.1000 473.1000 1032.9000 473.2500 ;
	    RECT 1035.9000 473.1000 1037.7001 473.2500 ;
	    RECT 1196.7001 474.7500 1198.5000 474.9000 ;
	    RECT 1268.7001 474.7500 1270.5000 474.9000 ;
	    RECT 1304.7001 474.7500 1306.5000 474.9000 ;
	    RECT 1196.7001 473.2500 1306.5000 474.7500 ;
	    RECT 1196.7001 473.1000 1198.5000 473.2500 ;
	    RECT 1268.7001 473.1000 1270.5000 473.2500 ;
	    RECT 1304.7001 473.1000 1306.5000 473.2500 ;
	    RECT 1448.7001 474.7500 1450.5000 474.9000 ;
	    RECT 1479.9000 474.7500 1481.7001 474.9000 ;
	    RECT 1448.7001 473.2500 1481.7001 474.7500 ;
	    RECT 1448.7001 473.1000 1450.5000 473.2500 ;
	    RECT 1479.9000 473.1000 1481.7001 473.2500 ;
	    RECT 323.1000 468.7500 324.9000 468.9000 ;
	    RECT 339.9000 468.7500 341.7000 468.9000 ;
	    RECT 323.1000 467.2500 341.7000 468.7500 ;
	    RECT 323.1000 467.1000 324.9000 467.2500 ;
	    RECT 339.9000 467.1000 341.7000 467.2500 ;
	    RECT 392.7000 468.7500 394.5000 468.9000 ;
	    RECT 426.3000 468.7500 428.1000 468.9000 ;
	    RECT 392.7000 467.2500 428.1000 468.7500 ;
	    RECT 392.7000 467.1000 394.5000 467.2500 ;
	    RECT 426.3000 467.1000 428.1000 467.2500 ;
	    RECT 803.1000 468.7500 804.9000 468.9000 ;
	    RECT 819.9000 468.7500 821.7000 468.9000 ;
	    RECT 803.1000 467.2500 821.7000 468.7500 ;
	    RECT 803.1000 467.1000 804.9000 467.2500 ;
	    RECT 819.9000 467.1000 821.7000 467.2500 ;
	    RECT 990.3000 468.7500 992.1000 468.9000 ;
	    RECT 995.1000 468.7500 996.9000 468.9000 ;
	    RECT 1021.5000 468.7500 1023.3000 468.9000 ;
	    RECT 990.3000 467.2500 1023.3000 468.7500 ;
	    RECT 990.3000 467.1000 992.1000 467.2500 ;
	    RECT 995.1000 467.1000 996.9000 467.2500 ;
	    RECT 1021.5000 467.1000 1023.3000 467.2500 ;
	    RECT 1026.3000 468.7500 1028.1000 468.9000 ;
	    RECT 1091.1000 468.7500 1092.9000 468.9000 ;
	    RECT 1026.3000 467.2500 1092.9000 468.7500 ;
	    RECT 1026.3000 467.1000 1028.1000 467.2500 ;
	    RECT 1091.1000 467.1000 1092.9000 467.2500 ;
	    RECT 1153.5000 468.7500 1155.3000 468.9000 ;
	    RECT 1199.1000 468.7500 1200.9000 468.9000 ;
	    RECT 1153.5000 467.2500 1200.9000 468.7500 ;
	    RECT 1153.5000 467.1000 1155.3000 467.2500 ;
	    RECT 1199.1000 467.1000 1200.9000 467.2500 ;
	    RECT 1237.5000 468.7500 1239.3000 468.9000 ;
	    RECT 1273.5000 468.7500 1275.3000 468.9000 ;
	    RECT 1287.9000 468.7500 1289.7001 468.9000 ;
	    RECT 1237.5000 467.2500 1289.7001 468.7500 ;
	    RECT 1237.5000 467.1000 1239.3000 467.2500 ;
	    RECT 1273.5000 467.1000 1275.3000 467.2500 ;
	    RECT 1287.9000 467.1000 1289.7001 467.2500 ;
	    RECT 1311.9000 468.7500 1313.7001 468.9000 ;
	    RECT 1335.9000 468.7500 1337.7001 468.9000 ;
	    RECT 1311.9000 467.2500 1337.7001 468.7500 ;
	    RECT 1311.9000 467.1000 1313.7001 467.2500 ;
	    RECT 1335.9000 467.1000 1337.7001 467.2500 ;
	    RECT 1410.3000 468.7500 1412.1000 468.9000 ;
	    RECT 1448.7001 468.7500 1450.5000 468.9000 ;
	    RECT 1410.3000 467.2500 1450.5000 468.7500 ;
	    RECT 1410.3000 467.1000 1412.1000 467.2500 ;
	    RECT 1448.7001 467.1000 1450.5000 467.2500 ;
	    RECT 1484.7001 468.7500 1486.5000 468.9000 ;
	    RECT 1489.5000 468.7500 1491.3000 468.9000 ;
	    RECT 1484.7001 467.2500 1491.3000 468.7500 ;
	    RECT 1484.7001 467.1000 1486.5000 467.2500 ;
	    RECT 1489.5000 467.1000 1491.3000 467.2500 ;
	    RECT 1539.9000 468.7500 1541.7001 468.9000 ;
	    RECT 1547.1000 468.7500 1548.9000 468.9000 ;
	    RECT 1539.9000 467.2500 1548.9000 468.7500 ;
	    RECT 1539.9000 467.1000 1541.7001 467.2500 ;
	    RECT 1547.1000 467.1000 1548.9000 467.2500 ;
	    RECT 1556.7001 468.7500 1558.5000 468.9000 ;
	    RECT 1561.5000 468.7500 1563.3000 468.9000 ;
	    RECT 1556.7001 467.2500 1563.3000 468.7500 ;
	    RECT 1556.7001 467.1000 1558.5000 467.2500 ;
	    RECT 1561.5000 467.1000 1563.3000 467.2500 ;
	    RECT 133.5000 462.7500 135.3000 462.9000 ;
	    RECT 169.5000 462.7500 171.3000 462.9000 ;
	    RECT 234.3000 462.7500 236.1000 462.9000 ;
	    RECT 133.5000 461.2500 236.1000 462.7500 ;
	    RECT 133.5000 461.1000 135.3000 461.2500 ;
	    RECT 169.5000 461.1000 171.3000 461.2500 ;
	    RECT 234.3000 461.1000 236.1000 461.2500 ;
	    RECT 349.5000 462.7500 351.3000 462.9000 ;
	    RECT 452.7000 462.7500 454.5000 462.9000 ;
	    RECT 349.5000 461.2500 454.5000 462.7500 ;
	    RECT 349.5000 461.1000 351.3000 461.2500 ;
	    RECT 452.7000 461.1000 454.5000 461.2500 ;
	    RECT 618.3000 462.7500 620.1000 462.9000 ;
	    RECT 649.5000 462.7500 651.3000 462.9000 ;
	    RECT 618.3000 461.2500 651.3000 462.7500 ;
	    RECT 618.3000 461.1000 620.1000 461.2500 ;
	    RECT 649.5000 461.1000 651.3000 461.2500 ;
	    RECT 786.3000 462.7500 788.1000 462.9000 ;
	    RECT 793.5000 462.7500 795.3000 462.9000 ;
	    RECT 786.3000 461.2500 795.3000 462.7500 ;
	    RECT 786.3000 461.1000 788.1000 461.2500 ;
	    RECT 793.5000 461.1000 795.3000 461.2500 ;
	    RECT 1028.7001 462.7500 1030.5000 462.9000 ;
	    RECT 1045.5000 462.7500 1047.3000 462.9000 ;
	    RECT 1028.7001 461.2500 1047.3000 462.7500 ;
	    RECT 1028.7001 461.1000 1030.5000 461.2500 ;
	    RECT 1045.5000 461.1000 1047.3000 461.2500 ;
	    RECT 1098.3000 462.7500 1100.1000 462.9000 ;
	    RECT 1103.1000 462.7500 1104.9000 462.9000 ;
	    RECT 1115.1000 462.7500 1116.9000 462.9000 ;
	    RECT 1134.3000 462.7500 1136.1000 462.9000 ;
	    RECT 1098.3000 461.2500 1136.1000 462.7500 ;
	    RECT 1098.3000 461.1000 1100.1000 461.2500 ;
	    RECT 1103.1000 461.1000 1104.9000 461.2500 ;
	    RECT 1115.1000 461.1000 1116.9000 461.2500 ;
	    RECT 1134.3000 461.1000 1136.1000 461.2500 ;
	    RECT 1177.5000 462.7500 1179.3000 462.9000 ;
	    RECT 1376.7001 462.7500 1378.5000 462.9000 ;
	    RECT 1177.5000 461.2500 1378.5000 462.7500 ;
	    RECT 1177.5000 461.1000 1179.3000 461.2500 ;
	    RECT 1376.7001 461.1000 1378.5000 461.2500 ;
	    RECT 1383.9000 462.7500 1385.7001 462.9000 ;
	    RECT 1393.5000 462.7500 1395.3000 462.9000 ;
	    RECT 1383.9000 461.2500 1395.3000 462.7500 ;
	    RECT 1383.9000 461.1000 1385.7001 461.2500 ;
	    RECT 1393.5000 461.1000 1395.3000 461.2500 ;
	    RECT 1523.1000 462.7500 1524.9000 462.9000 ;
	    RECT 1542.3000 462.7500 1544.1000 462.9000 ;
	    RECT 1523.1000 461.2500 1544.1000 462.7500 ;
	    RECT 1523.1000 461.1000 1524.9000 461.2500 ;
	    RECT 1542.3000 461.1000 1544.1000 461.2500 ;
	    RECT 85.5000 456.7500 87.3000 456.9000 ;
	    RECT 143.1000 456.7500 144.9000 456.9000 ;
	    RECT 85.5000 455.2500 144.9000 456.7500 ;
	    RECT 85.5000 455.1000 87.3000 455.2500 ;
	    RECT 143.1000 455.1000 144.9000 455.2500 ;
	    RECT 267.9000 456.7500 269.7000 456.9000 ;
	    RECT 287.1000 456.7500 288.9000 456.9000 ;
	    RECT 267.9000 455.2500 288.9000 456.7500 ;
	    RECT 267.9000 455.1000 269.7000 455.2500 ;
	    RECT 287.1000 455.1000 288.9000 455.2500 ;
	    RECT 548.7000 456.7500 550.5000 456.9000 ;
	    RECT 572.7000 456.7500 574.5000 456.9000 ;
	    RECT 603.9000 456.7500 605.7000 456.9000 ;
	    RECT 548.7000 455.2500 605.7000 456.7500 ;
	    RECT 548.7000 455.1000 550.5000 455.2500 ;
	    RECT 572.7000 455.1000 574.5000 455.2500 ;
	    RECT 603.9000 455.1000 605.7000 455.2500 ;
	    RECT 635.1000 456.7500 636.9000 456.9000 ;
	    RECT 687.9000 456.7500 689.7000 456.9000 ;
	    RECT 635.1000 455.2500 689.7000 456.7500 ;
	    RECT 635.1000 455.1000 636.9000 455.2500 ;
	    RECT 687.9000 455.1000 689.7000 455.2500 ;
	    RECT 779.1000 456.7500 780.9000 456.9000 ;
	    RECT 954.3000 456.7500 956.1000 456.9000 ;
	    RECT 779.1000 455.2500 956.1000 456.7500 ;
	    RECT 779.1000 455.1000 780.9000 455.2500 ;
	    RECT 954.3000 455.1000 956.1000 455.2500 ;
	    RECT 1083.9000 456.7500 1085.7001 456.9000 ;
	    RECT 1100.7001 456.7500 1102.5000 456.9000 ;
	    RECT 1083.9000 455.2500 1102.5000 456.7500 ;
	    RECT 1083.9000 455.1000 1085.7001 455.2500 ;
	    RECT 1100.7001 455.1000 1102.5000 455.2500 ;
	    RECT 1110.3000 456.7500 1112.1000 456.9000 ;
	    RECT 1146.3000 456.7500 1148.1000 456.9000 ;
	    RECT 1110.3000 455.2500 1148.1000 456.7500 ;
	    RECT 1110.3000 455.1000 1112.1000 455.2500 ;
	    RECT 1146.3000 455.1000 1148.1000 455.2500 ;
	    RECT 1179.9000 456.7500 1181.7001 456.9000 ;
	    RECT 1201.5000 456.7500 1203.3000 456.9000 ;
	    RECT 1179.9000 455.2500 1203.3000 456.7500 ;
	    RECT 1179.9000 455.1000 1181.7001 455.2500 ;
	    RECT 1201.5000 455.1000 1203.3000 455.2500 ;
	    RECT 1220.7001 456.7500 1222.5000 456.9000 ;
	    RECT 1261.5000 456.7500 1263.3000 456.9000 ;
	    RECT 1220.7001 455.2500 1263.3000 456.7500 ;
	    RECT 1220.7001 455.1000 1222.5000 455.2500 ;
	    RECT 1261.5000 455.1000 1263.3000 455.2500 ;
	    RECT 1266.3000 456.7500 1268.1000 456.9000 ;
	    RECT 1280.7001 456.7500 1282.5000 456.9000 ;
	    RECT 1302.3000 456.7500 1304.1000 456.9000 ;
	    RECT 1266.3000 455.2500 1304.1000 456.7500 ;
	    RECT 1266.3000 455.1000 1268.1000 455.2500 ;
	    RECT 1280.7001 455.1000 1282.5000 455.2500 ;
	    RECT 1302.3000 455.1000 1304.1000 455.2500 ;
	    RECT 1391.1000 456.7500 1392.9000 456.9000 ;
	    RECT 1419.9000 456.7500 1421.7001 456.9000 ;
	    RECT 1391.1000 455.2500 1421.7001 456.7500 ;
	    RECT 1391.1000 455.1000 1392.9000 455.2500 ;
	    RECT 1419.9000 455.1000 1421.7001 455.2500 ;
	    RECT 1532.7001 456.7500 1534.5000 456.9000 ;
	    RECT 1554.3000 456.7500 1556.1000 456.9000 ;
	    RECT 1532.7001 455.2500 1556.1000 456.7500 ;
	    RECT 1532.7001 455.1000 1534.5000 455.2500 ;
	    RECT 1554.3000 455.1000 1556.1000 455.2500 ;
	    RECT 162.3000 450.7500 164.1000 450.9000 ;
	    RECT 198.3000 450.7500 200.1000 450.9000 ;
	    RECT 162.3000 449.2500 200.1000 450.7500 ;
	    RECT 162.3000 449.1000 164.1000 449.2500 ;
	    RECT 198.3000 449.1000 200.1000 449.2500 ;
	    RECT 627.9000 450.7500 629.7000 450.9000 ;
	    RECT 632.7000 450.7500 634.5000 450.9000 ;
	    RECT 627.9000 449.2500 634.5000 450.7500 ;
	    RECT 627.9000 449.1000 629.7000 449.2500 ;
	    RECT 632.7000 449.1000 634.5000 449.2500 ;
	    RECT 656.7000 450.7500 658.5000 450.9000 ;
	    RECT 666.3000 450.7500 668.1000 450.9000 ;
	    RECT 752.7000 450.7500 754.5000 450.9000 ;
	    RECT 656.7000 449.2500 754.5000 450.7500 ;
	    RECT 656.7000 449.1000 658.5000 449.2500 ;
	    RECT 666.3000 449.1000 668.1000 449.2500 ;
	    RECT 752.7000 449.1000 754.5000 449.2500 ;
	    RECT 870.3000 450.7500 872.1000 450.9000 ;
	    RECT 882.3000 450.7500 884.1000 450.9000 ;
	    RECT 870.3000 449.2500 884.1000 450.7500 ;
	    RECT 870.3000 449.1000 872.1000 449.2500 ;
	    RECT 882.3000 449.1000 884.1000 449.2500 ;
	    RECT 918.3000 450.7500 920.1000 450.9000 ;
	    RECT 1083.9000 450.7500 1085.7001 450.9000 ;
	    RECT 918.3000 449.2500 1085.7001 450.7500 ;
	    RECT 918.3000 449.1000 920.1000 449.2500 ;
	    RECT 1083.9000 449.1000 1085.7001 449.2500 ;
	    RECT 1167.9000 450.7500 1169.7001 450.9000 ;
	    RECT 1239.9000 450.7500 1241.7001 450.9000 ;
	    RECT 1167.9000 449.2500 1241.7001 450.7500 ;
	    RECT 1167.9000 449.1000 1169.7001 449.2500 ;
	    RECT 1239.9000 449.1000 1241.7001 449.2500 ;
	    RECT 131.1000 444.7500 132.9000 444.9000 ;
	    RECT 162.3000 444.7500 164.1000 444.9000 ;
	    RECT 131.1000 443.2500 164.1000 444.7500 ;
	    RECT 131.1000 443.1000 132.9000 443.2500 ;
	    RECT 162.3000 443.1000 164.1000 443.2500 ;
	    RECT 169.5000 444.7500 171.3000 444.9000 ;
	    RECT 193.5000 444.7500 195.3000 444.9000 ;
	    RECT 169.5000 443.2500 195.3000 444.7500 ;
	    RECT 169.5000 443.1000 171.3000 443.2500 ;
	    RECT 193.5000 443.1000 195.3000 443.2500 ;
	    RECT 258.3000 444.7500 260.1000 444.9000 ;
	    RECT 267.9000 444.7500 269.7000 444.9000 ;
	    RECT 258.3000 443.2500 269.7000 444.7500 ;
	    RECT 258.3000 443.1000 260.1000 443.2500 ;
	    RECT 267.9000 443.1000 269.7000 443.2500 ;
	    RECT 452.7000 444.7500 454.5000 444.9000 ;
	    RECT 486.3000 444.7500 488.1000 444.9000 ;
	    RECT 491.1000 444.7500 492.9000 444.9000 ;
	    RECT 452.7000 443.2500 492.9000 444.7500 ;
	    RECT 452.7000 443.1000 454.5000 443.2500 ;
	    RECT 486.3000 443.1000 488.1000 443.2500 ;
	    RECT 491.1000 443.1000 492.9000 443.2500 ;
	    RECT 637.5000 444.7500 639.3000 444.9000 ;
	    RECT 699.9000 444.7500 701.7000 444.9000 ;
	    RECT 637.5000 443.2500 701.7000 444.7500 ;
	    RECT 637.5000 443.1000 639.3000 443.2500 ;
	    RECT 699.9000 443.1000 701.7000 443.2500 ;
	    RECT 762.3000 444.7500 764.1000 444.9000 ;
	    RECT 774.3000 444.7500 776.1000 444.9000 ;
	    RECT 762.3000 443.2500 776.1000 444.7500 ;
	    RECT 762.3000 443.1000 764.1000 443.2500 ;
	    RECT 774.3000 443.1000 776.1000 443.2500 ;
	    RECT 1031.1000 444.7500 1032.9000 444.9000 ;
	    RECT 1052.7001 444.7500 1054.5000 444.9000 ;
	    RECT 1031.1000 443.2500 1054.5000 444.7500 ;
	    RECT 1031.1000 443.1000 1032.9000 443.2500 ;
	    RECT 1052.7001 443.1000 1054.5000 443.2500 ;
	    RECT 1083.9000 444.7500 1085.7001 444.9000 ;
	    RECT 1122.3000 444.7500 1124.1000 444.9000 ;
	    RECT 1083.9000 443.2500 1124.1000 444.7500 ;
	    RECT 1083.9000 443.1000 1085.7001 443.2500 ;
	    RECT 1122.3000 443.1000 1124.1000 443.2500 ;
	    RECT 1139.1000 444.7500 1140.9000 444.9000 ;
	    RECT 1167.9000 444.7500 1169.7001 444.9000 ;
	    RECT 1139.1000 443.2500 1169.7001 444.7500 ;
	    RECT 1139.1000 443.1000 1140.9000 443.2500 ;
	    RECT 1167.9000 443.1000 1169.7001 443.2500 ;
	    RECT 1189.5000 444.7500 1191.3000 444.9000 ;
	    RECT 1275.9000 444.7500 1277.7001 444.9000 ;
	    RECT 1292.7001 444.7500 1294.5000 444.9000 ;
	    RECT 1189.5000 443.2500 1294.5000 444.7500 ;
	    RECT 1189.5000 443.1000 1191.3000 443.2500 ;
	    RECT 1275.9000 443.1000 1277.7001 443.2500 ;
	    RECT 1292.7001 443.1000 1294.5000 443.2500 ;
	    RECT 1328.7001 444.7500 1330.5000 444.9000 ;
	    RECT 1345.5000 444.7500 1347.3000 444.9000 ;
	    RECT 1328.7001 443.2500 1347.3000 444.7500 ;
	    RECT 1328.7001 443.1000 1330.5000 443.2500 ;
	    RECT 1345.5000 443.1000 1347.3000 443.2500 ;
	    RECT 1367.1000 444.7500 1368.9000 444.9000 ;
	    RECT 1417.5000 444.7500 1419.3000 444.9000 ;
	    RECT 1367.1000 443.2500 1419.3000 444.7500 ;
	    RECT 1367.1000 443.1000 1368.9000 443.2500 ;
	    RECT 1417.5000 443.1000 1419.3000 443.2500 ;
	    RECT 35.1000 438.7500 36.9000 438.9000 ;
	    RECT 66.3000 438.7500 68.1000 438.9000 ;
	    RECT 35.1000 437.2500 68.1000 438.7500 ;
	    RECT 35.1000 437.1000 36.9000 437.2500 ;
	    RECT 66.3000 437.1000 68.1000 437.2500 ;
	    RECT 215.1000 438.7500 216.9000 438.9000 ;
	    RECT 255.9000 438.7500 257.7000 438.9000 ;
	    RECT 215.1000 437.2500 257.7000 438.7500 ;
	    RECT 215.1000 437.1000 216.9000 437.2500 ;
	    RECT 255.9000 437.1000 257.7000 437.2500 ;
	    RECT 769.5000 438.7500 771.3000 438.9000 ;
	    RECT 875.1000 438.7500 876.9000 438.9000 ;
	    RECT 947.1000 438.7500 948.9000 438.9000 ;
	    RECT 769.5000 437.2500 948.9000 438.7500 ;
	    RECT 769.5000 437.1000 771.3000 437.2500 ;
	    RECT 875.1000 437.1000 876.9000 437.2500 ;
	    RECT 947.1000 437.1000 948.9000 437.2500 ;
	    RECT 956.7000 438.7500 958.5000 438.9000 ;
	    RECT 1021.5000 438.7500 1023.3000 438.9000 ;
	    RECT 1040.7001 438.7500 1042.5000 438.9000 ;
	    RECT 1055.1000 438.7500 1056.9000 438.9000 ;
	    RECT 956.7000 437.2500 1056.9000 438.7500 ;
	    RECT 956.7000 437.1000 958.5000 437.2500 ;
	    RECT 1021.5000 437.1000 1023.3000 437.2500 ;
	    RECT 1040.7001 437.1000 1042.5000 437.2500 ;
	    RECT 1055.1000 437.1000 1056.9000 437.2500 ;
	    RECT 1163.1000 438.7500 1164.9000 438.9000 ;
	    RECT 1189.5000 438.7500 1191.3000 438.9000 ;
	    RECT 1163.1000 437.2500 1191.3000 438.7500 ;
	    RECT 1163.1000 437.1000 1164.9000 437.2500 ;
	    RECT 1189.5000 437.1000 1191.3000 437.2500 ;
	    RECT 1201.5000 438.7500 1203.3000 438.9000 ;
	    RECT 1237.5000 438.7500 1239.3000 438.9000 ;
	    RECT 1201.5000 437.2500 1239.3000 438.7500 ;
	    RECT 1201.5000 437.1000 1203.3000 437.2500 ;
	    RECT 1237.5000 437.1000 1239.3000 437.2500 ;
	    RECT 1328.7001 438.7500 1330.5000 438.9000 ;
	    RECT 1335.9000 438.7500 1337.7001 438.9000 ;
	    RECT 1328.7001 437.2500 1337.7001 438.7500 ;
	    RECT 1328.7001 437.1000 1330.5000 437.2500 ;
	    RECT 1335.9000 437.1000 1337.7001 437.2500 ;
	    RECT 1343.1000 438.7500 1344.9000 438.9000 ;
	    RECT 1537.5000 438.7500 1539.3000 438.9000 ;
	    RECT 1343.1000 437.2500 1539.3000 438.7500 ;
	    RECT 1343.1000 437.1000 1344.9000 437.2500 ;
	    RECT 1537.5000 437.1000 1539.3000 437.2500 ;
	    RECT 183.9000 432.7500 185.7000 432.9000 ;
	    RECT 224.7000 432.7500 226.5000 432.9000 ;
	    RECT 183.9000 431.2500 226.5000 432.7500 ;
	    RECT 183.9000 431.1000 185.7000 431.2500 ;
	    RECT 224.7000 431.1000 226.5000 431.2500 ;
	    RECT 267.9000 432.7500 269.7000 432.9000 ;
	    RECT 279.9000 432.7500 281.7000 432.9000 ;
	    RECT 267.9000 431.2500 281.7000 432.7500 ;
	    RECT 267.9000 431.1000 269.7000 431.2500 ;
	    RECT 279.9000 431.1000 281.7000 431.2500 ;
	    RECT 308.7000 432.7500 310.5000 432.9000 ;
	    RECT 325.5000 432.7500 327.3000 432.9000 ;
	    RECT 308.7000 431.2500 327.3000 432.7500 ;
	    RECT 308.7000 431.1000 310.5000 431.2500 ;
	    RECT 325.5000 431.1000 327.3000 431.2500 ;
	    RECT 627.9000 432.7500 629.7000 432.9000 ;
	    RECT 642.3000 432.7500 644.1000 432.9000 ;
	    RECT 699.9000 432.7500 701.7000 432.9000 ;
	    RECT 627.9000 431.2500 701.7000 432.7500 ;
	    RECT 627.9000 431.1000 629.7000 431.2500 ;
	    RECT 642.3000 431.1000 644.1000 431.2500 ;
	    RECT 699.9000 431.1000 701.7000 431.2500 ;
	    RECT 774.3000 432.7500 776.1000 432.9000 ;
	    RECT 824.7000 432.7500 826.5000 432.9000 ;
	    RECT 774.3000 431.2500 826.5000 432.7500 ;
	    RECT 774.3000 431.1000 776.1000 431.2500 ;
	    RECT 824.7000 431.1000 826.5000 431.2500 ;
	    RECT 1095.9000 432.7500 1097.7001 432.9000 ;
	    RECT 1139.1000 432.7500 1140.9000 432.9000 ;
	    RECT 1095.9000 431.2500 1140.9000 432.7500 ;
	    RECT 1095.9000 431.1000 1097.7001 431.2500 ;
	    RECT 1139.1000 431.1000 1140.9000 431.2500 ;
	    RECT 1155.9000 432.7500 1157.7001 432.9000 ;
	    RECT 1172.7001 432.7500 1174.5000 432.9000 ;
	    RECT 1304.7001 432.7500 1306.5000 432.9000 ;
	    RECT 1155.9000 431.2500 1306.5000 432.7500 ;
	    RECT 1155.9000 431.1000 1157.7001 431.2500 ;
	    RECT 1172.7001 431.1000 1174.5000 431.2500 ;
	    RECT 1304.7001 431.1000 1306.5000 431.2500 ;
	    RECT 1443.9000 432.7500 1445.7001 432.9000 ;
	    RECT 1458.3000 432.7500 1460.1000 432.9000 ;
	    RECT 1443.9000 431.2500 1460.1000 432.7500 ;
	    RECT 1443.9000 431.1000 1445.7001 431.2500 ;
	    RECT 1458.3000 431.1000 1460.1000 431.2500 ;
	    RECT 162.3000 426.7500 164.1000 426.9000 ;
	    RECT 193.5000 426.7500 195.3000 426.9000 ;
	    RECT 162.3000 425.2500 195.3000 426.7500 ;
	    RECT 162.3000 425.1000 164.1000 425.2500 ;
	    RECT 193.5000 425.1000 195.3000 425.2500 ;
	    RECT 311.1000 426.7500 312.9000 426.9000 ;
	    RECT 315.9000 426.7500 317.7000 426.9000 ;
	    RECT 311.1000 425.2500 317.7000 426.7500 ;
	    RECT 311.1000 425.1000 312.9000 425.2500 ;
	    RECT 315.9000 425.1000 317.7000 425.2500 ;
	    RECT 606.3000 426.7500 608.1000 426.9000 ;
	    RECT 781.5000 426.7500 783.3000 426.9000 ;
	    RECT 795.9000 426.7500 797.7000 426.9000 ;
	    RECT 606.3000 425.2500 797.7000 426.7500 ;
	    RECT 606.3000 425.1000 608.1000 425.2500 ;
	    RECT 781.5000 425.1000 783.3000 425.2500 ;
	    RECT 795.9000 425.1000 797.7000 425.2500 ;
	    RECT 877.5000 426.7500 879.3000 426.9000 ;
	    RECT 899.1000 426.7500 900.9000 426.9000 ;
	    RECT 877.5000 425.2500 900.9000 426.7500 ;
	    RECT 877.5000 425.1000 879.3000 425.2500 ;
	    RECT 899.1000 425.1000 900.9000 425.2500 ;
	    RECT 1151.1000 426.7500 1152.9000 426.9000 ;
	    RECT 1163.1000 426.7500 1164.9000 426.9000 ;
	    RECT 1151.1000 425.2500 1164.9000 426.7500 ;
	    RECT 1151.1000 425.1000 1152.9000 425.2500 ;
	    RECT 1163.1000 425.1000 1164.9000 425.2500 ;
	    RECT 1247.1000 426.7500 1248.9000 426.9000 ;
	    RECT 1273.5000 426.7500 1275.3000 426.9000 ;
	    RECT 1247.1000 425.2500 1275.3000 426.7500 ;
	    RECT 1247.1000 425.1000 1248.9000 425.2500 ;
	    RECT 1273.5000 425.1000 1275.3000 425.2500 ;
	    RECT 1326.3000 426.7500 1328.1000 426.9000 ;
	    RECT 1369.5000 426.7500 1371.3000 426.9000 ;
	    RECT 1410.3000 426.7500 1412.1000 426.9000 ;
	    RECT 1326.3000 425.2500 1412.1000 426.7500 ;
	    RECT 1326.3000 425.1000 1328.1000 425.2500 ;
	    RECT 1369.5000 425.1000 1371.3000 425.2500 ;
	    RECT 1410.3000 425.1000 1412.1000 425.2500 ;
	    RECT 35.1000 420.7500 36.9000 420.9000 ;
	    RECT 63.9000 420.7500 65.7000 420.9000 ;
	    RECT 71.1000 420.7500 72.9000 420.9000 ;
	    RECT 87.9000 420.7500 89.7000 420.9000 ;
	    RECT 35.1000 419.2500 89.7000 420.7500 ;
	    RECT 35.1000 419.1000 36.9000 419.2500 ;
	    RECT 63.9000 419.1000 65.7000 419.2500 ;
	    RECT 71.1000 419.1000 72.9000 419.2500 ;
	    RECT 87.9000 419.1000 89.7000 419.2500 ;
	    RECT 119.1000 420.7500 120.9000 420.9000 ;
	    RECT 174.3000 420.7500 176.1000 420.9000 ;
	    RECT 119.1000 419.2500 176.1000 420.7500 ;
	    RECT 119.1000 419.1000 120.9000 419.2500 ;
	    RECT 174.3000 419.1000 176.1000 419.2500 ;
	    RECT 284.7000 420.7500 286.5000 420.9000 ;
	    RECT 301.5000 420.7500 303.3000 420.9000 ;
	    RECT 284.7000 419.2500 303.3000 420.7500 ;
	    RECT 284.7000 419.1000 286.5000 419.2500 ;
	    RECT 301.5000 419.1000 303.3000 419.2500 ;
	    RECT 313.5000 420.7500 315.3000 420.9000 ;
	    RECT 330.3000 420.7500 332.1000 420.9000 ;
	    RECT 313.5000 419.2500 332.1000 420.7500 ;
	    RECT 313.5000 419.1000 315.3000 419.2500 ;
	    RECT 330.3000 419.1000 332.1000 419.2500 ;
	    RECT 399.9000 420.7500 401.7000 420.9000 ;
	    RECT 404.7000 420.7500 406.5000 420.9000 ;
	    RECT 399.9000 419.2500 406.5000 420.7500 ;
	    RECT 399.9000 419.1000 401.7000 419.2500 ;
	    RECT 404.7000 419.1000 406.5000 419.2500 ;
	    RECT 467.1000 420.7500 468.9000 420.9000 ;
	    RECT 627.9000 420.7500 629.7000 420.9000 ;
	    RECT 467.1000 419.2500 629.7000 420.7500 ;
	    RECT 467.1000 419.1000 468.9000 419.2500 ;
	    RECT 627.9000 419.1000 629.7000 419.2500 ;
	    RECT 687.9000 420.7500 689.7000 420.9000 ;
	    RECT 716.7000 420.7500 718.5000 420.9000 ;
	    RECT 738.3000 420.7500 740.1000 420.9000 ;
	    RECT 841.5000 420.7500 843.3000 420.9000 ;
	    RECT 903.9000 420.7500 905.7000 420.9000 ;
	    RECT 687.9000 419.2500 905.7000 420.7500 ;
	    RECT 687.9000 419.1000 689.7000 419.2500 ;
	    RECT 716.7000 419.1000 718.5000 419.2500 ;
	    RECT 738.3000 419.1000 740.1000 419.2500 ;
	    RECT 841.5000 419.1000 843.3000 419.2500 ;
	    RECT 903.9000 419.1000 905.7000 419.2500 ;
	    RECT 1057.5000 420.7500 1059.3000 420.9000 ;
	    RECT 1064.7001 420.7500 1066.5000 420.9000 ;
	    RECT 1057.5000 419.2500 1066.5000 420.7500 ;
	    RECT 1057.5000 419.1000 1059.3000 419.2500 ;
	    RECT 1064.7001 419.1000 1066.5000 419.2500 ;
	    RECT 1155.9000 420.7500 1157.7001 420.9000 ;
	    RECT 1196.7001 420.7500 1198.5000 420.9000 ;
	    RECT 1155.9000 419.2500 1198.5000 420.7500 ;
	    RECT 1155.9000 419.1000 1157.7001 419.2500 ;
	    RECT 1196.7001 419.1000 1198.5000 419.2500 ;
	    RECT 1244.7001 420.7500 1246.5000 420.9000 ;
	    RECT 1275.9000 420.7500 1277.7001 420.9000 ;
	    RECT 1244.7001 419.2500 1277.7001 420.7500 ;
	    RECT 1244.7001 419.1000 1246.5000 419.2500 ;
	    RECT 1275.9000 419.1000 1277.7001 419.2500 ;
	    RECT 1323.9000 420.7500 1325.7001 420.9000 ;
	    RECT 1328.7001 420.7500 1330.5000 420.9000 ;
	    RECT 1323.9000 419.2500 1330.5000 420.7500 ;
	    RECT 1323.9000 419.1000 1325.7001 419.2500 ;
	    RECT 1328.7001 419.1000 1330.5000 419.2500 ;
	    RECT 1345.5000 420.7500 1347.3000 420.9000 ;
	    RECT 1359.9000 420.7500 1361.7001 420.9000 ;
	    RECT 1367.1000 420.7500 1368.9000 420.9000 ;
	    RECT 1345.5000 419.2500 1368.9000 420.7500 ;
	    RECT 1345.5000 419.1000 1347.3000 419.2500 ;
	    RECT 1359.9000 419.1000 1361.7001 419.2500 ;
	    RECT 1367.1000 419.1000 1368.9000 419.2500 ;
	    RECT 1453.5000 420.7500 1455.3000 420.9000 ;
	    RECT 1508.7001 420.7500 1510.5000 420.9000 ;
	    RECT 1453.5000 419.2500 1510.5000 420.7500 ;
	    RECT 1453.5000 419.1000 1455.3000 419.2500 ;
	    RECT 1508.7001 419.1000 1510.5000 419.2500 ;
	    RECT 1530.3000 420.7500 1532.1000 420.9000 ;
	    RECT 1544.7001 420.7500 1546.5000 420.9000 ;
	    RECT 1530.3000 419.2500 1546.5000 420.7500 ;
	    RECT 1530.3000 419.1000 1532.1000 419.2500 ;
	    RECT 1544.7001 419.1000 1546.5000 419.2500 ;
	    RECT 32.7000 414.7500 34.5000 414.9000 ;
	    RECT 126.3000 414.7500 128.1000 414.9000 ;
	    RECT 32.7000 413.2500 128.1000 414.7500 ;
	    RECT 32.7000 413.1000 34.5000 413.2500 ;
	    RECT 126.3000 413.1000 128.1000 413.2500 ;
	    RECT 133.5000 414.7500 135.3000 414.9000 ;
	    RECT 164.7000 414.7500 166.5000 414.9000 ;
	    RECT 133.5000 413.2500 166.5000 414.7500 ;
	    RECT 133.5000 413.1000 135.3000 413.2500 ;
	    RECT 164.7000 413.1000 166.5000 413.2500 ;
	    RECT 733.5000 414.7500 735.3000 414.9000 ;
	    RECT 817.5000 414.7500 819.3000 414.9000 ;
	    RECT 733.5000 413.2500 819.3000 414.7500 ;
	    RECT 733.5000 413.1000 735.3000 413.2500 ;
	    RECT 817.5000 413.1000 819.3000 413.2500 ;
	    RECT 1052.7001 414.7500 1054.5000 414.9000 ;
	    RECT 1151.1000 414.7500 1152.9000 414.9000 ;
	    RECT 1052.7001 413.2500 1152.9000 414.7500 ;
	    RECT 1052.7001 413.1000 1054.5000 413.2500 ;
	    RECT 1151.1000 413.1000 1152.9000 413.2500 ;
	    RECT 1170.3000 414.7500 1172.1000 414.9000 ;
	    RECT 1191.9000 414.7500 1193.7001 414.9000 ;
	    RECT 1201.5000 414.7500 1203.3000 414.9000 ;
	    RECT 1273.5000 414.7500 1275.3000 414.9000 ;
	    RECT 1170.3000 413.2500 1275.3000 414.7500 ;
	    RECT 1170.3000 413.1000 1172.1000 413.2500 ;
	    RECT 1191.9000 413.1000 1193.7001 413.2500 ;
	    RECT 1201.5000 413.1000 1203.3000 413.2500 ;
	    RECT 1273.5000 413.1000 1275.3000 413.2500 ;
	    RECT 1311.9000 414.7500 1313.7001 414.9000 ;
	    RECT 1357.5000 414.7500 1359.3000 414.9000 ;
	    RECT 1383.9000 414.7500 1385.7001 414.9000 ;
	    RECT 1311.9000 413.2500 1385.7001 414.7500 ;
	    RECT 1311.9000 413.1000 1313.7001 413.2500 ;
	    RECT 1357.5000 413.1000 1359.3000 413.2500 ;
	    RECT 1383.9000 413.1000 1385.7001 413.2500 ;
	    RECT 1393.5000 414.7500 1395.3000 414.9000 ;
	    RECT 1419.9000 414.7500 1421.7001 414.9000 ;
	    RECT 1393.5000 413.2500 1421.7001 414.7500 ;
	    RECT 1393.5000 413.1000 1395.3000 413.2500 ;
	    RECT 1419.9000 413.1000 1421.7001 413.2500 ;
	    RECT 1487.1000 414.7500 1488.9000 414.9000 ;
	    RECT 1518.3000 414.7500 1520.1000 414.9000 ;
	    RECT 1487.1000 413.2500 1520.1000 414.7500 ;
	    RECT 1487.1000 413.1000 1488.9000 413.2500 ;
	    RECT 1518.3000 413.1000 1520.1000 413.2500 ;
	    RECT 1539.9000 414.7500 1541.7001 414.9000 ;
	    RECT 1566.3000 414.7500 1568.1000 414.9000 ;
	    RECT 1539.9000 413.2500 1568.1000 414.7500 ;
	    RECT 1539.9000 413.1000 1541.7001 413.2500 ;
	    RECT 1566.3000 413.1000 1568.1000 413.2500 ;
	    RECT 147.9000 408.7500 149.7000 408.9000 ;
	    RECT 299.1000 408.7500 300.9000 408.9000 ;
	    RECT 147.9000 407.2500 300.9000 408.7500 ;
	    RECT 147.9000 407.1000 149.7000 407.2500 ;
	    RECT 299.1000 407.1000 300.9000 407.2500 ;
	    RECT 462.3000 408.7500 464.1000 408.9000 ;
	    RECT 512.7000 408.7500 514.5000 408.9000 ;
	    RECT 462.3000 407.2500 514.5000 408.7500 ;
	    RECT 462.3000 407.1000 464.1000 407.2500 ;
	    RECT 512.7000 407.1000 514.5000 407.2500 ;
	    RECT 745.5000 408.7500 747.3000 408.9000 ;
	    RECT 812.7000 408.7500 814.5000 408.9000 ;
	    RECT 745.5000 407.2500 814.5000 408.7500 ;
	    RECT 745.5000 407.1000 747.3000 407.2500 ;
	    RECT 812.7000 407.1000 814.5000 407.2500 ;
	    RECT 944.7000 408.7500 946.5000 408.9000 ;
	    RECT 1040.7001 408.7500 1042.5000 408.9000 ;
	    RECT 944.7000 407.2500 1042.5000 408.7500 ;
	    RECT 944.7000 407.1000 946.5000 407.2500 ;
	    RECT 1040.7001 407.1000 1042.5000 407.2500 ;
	    RECT 1117.5000 408.7500 1119.3000 408.9000 ;
	    RECT 1148.7001 408.7500 1150.5000 408.9000 ;
	    RECT 1117.5000 407.2500 1150.5000 408.7500 ;
	    RECT 1117.5000 407.1000 1119.3000 407.2500 ;
	    RECT 1148.7001 407.1000 1150.5000 407.2500 ;
	    RECT 1206.3000 408.7500 1208.1000 408.9000 ;
	    RECT 1215.9000 408.7500 1217.7001 408.9000 ;
	    RECT 1237.5000 408.7500 1239.3000 408.9000 ;
	    RECT 1206.3000 407.2500 1239.3000 408.7500 ;
	    RECT 1206.3000 407.1000 1208.1000 407.2500 ;
	    RECT 1215.9000 407.1000 1217.7001 407.2500 ;
	    RECT 1237.5000 407.1000 1239.3000 407.2500 ;
	    RECT 1271.1000 408.7500 1272.9000 408.9000 ;
	    RECT 1280.7001 408.7500 1282.5000 408.9000 ;
	    RECT 1271.1000 407.2500 1282.5000 408.7500 ;
	    RECT 1271.1000 407.1000 1272.9000 407.2500 ;
	    RECT 1280.7001 407.1000 1282.5000 407.2500 ;
	    RECT 1350.3000 408.7500 1352.1000 408.9000 ;
	    RECT 1376.7001 408.7500 1378.5000 408.9000 ;
	    RECT 1350.3000 407.2500 1378.5000 408.7500 ;
	    RECT 1350.3000 407.1000 1352.1000 407.2500 ;
	    RECT 1376.7001 407.1000 1378.5000 407.2500 ;
	    RECT 1520.7001 408.7500 1522.5000 408.9000 ;
	    RECT 1549.5000 408.7500 1551.3000 408.9000 ;
	    RECT 1520.7001 407.2500 1551.3000 408.7500 ;
	    RECT 1520.7001 407.1000 1522.5000 407.2500 ;
	    RECT 1549.5000 407.1000 1551.3000 407.2500 ;
	    RECT 469.5000 402.7500 471.3000 402.9000 ;
	    RECT 503.1000 402.7500 504.9000 402.9000 ;
	    RECT 469.5000 401.2500 504.9000 402.7500 ;
	    RECT 469.5000 401.1000 471.3000 401.2500 ;
	    RECT 503.1000 401.1000 504.9000 401.2500 ;
	    RECT 764.7000 402.7500 766.5000 402.9000 ;
	    RECT 848.7000 402.7500 850.5000 402.9000 ;
	    RECT 939.9000 402.7500 941.7000 402.9000 ;
	    RECT 764.7000 401.2500 941.7000 402.7500 ;
	    RECT 764.7000 401.1000 766.5000 401.2500 ;
	    RECT 848.7000 401.1000 850.5000 401.2500 ;
	    RECT 939.9000 401.1000 941.7000 401.2500 ;
	    RECT 1146.3000 402.7500 1148.1000 402.9000 ;
	    RECT 1184.7001 402.7500 1186.5000 402.9000 ;
	    RECT 1146.3000 401.2500 1186.5000 402.7500 ;
	    RECT 1146.3000 401.1000 1148.1000 401.2500 ;
	    RECT 1184.7001 401.1000 1186.5000 401.2500 ;
	    RECT 1319.1000 402.7500 1320.9000 402.9000 ;
	    RECT 1333.5000 402.7500 1335.3000 402.9000 ;
	    RECT 1319.1000 401.2500 1335.3000 402.7500 ;
	    RECT 1319.1000 401.1000 1320.9000 401.2500 ;
	    RECT 1333.5000 401.1000 1335.3000 401.2500 ;
	    RECT 1350.3000 402.7500 1352.1000 402.9000 ;
	    RECT 1391.1000 402.7500 1392.9000 402.9000 ;
	    RECT 1407.9000 402.7500 1409.7001 402.9000 ;
	    RECT 1436.7001 402.7500 1438.5000 402.9000 ;
	    RECT 1350.3000 401.2500 1438.5000 402.7500 ;
	    RECT 1350.3000 401.1000 1352.1000 401.2500 ;
	    RECT 1391.1000 401.1000 1392.9000 401.2500 ;
	    RECT 1407.9000 401.1000 1409.7001 401.2500 ;
	    RECT 1436.7001 401.1000 1438.5000 401.2500 ;
	    RECT 1455.9000 402.7500 1457.7001 402.9000 ;
	    RECT 1475.1000 402.7500 1476.9000 402.9000 ;
	    RECT 1455.9000 401.2500 1476.9000 402.7500 ;
	    RECT 1455.9000 401.1000 1457.7001 401.2500 ;
	    RECT 1475.1000 401.1000 1476.9000 401.2500 ;
	    RECT 87.9000 396.7500 89.7000 396.9000 ;
	    RECT 119.1000 396.7500 120.9000 396.9000 ;
	    RECT 171.9000 396.7500 173.7000 396.9000 ;
	    RECT 87.9000 395.2500 173.7000 396.7500 ;
	    RECT 87.9000 395.1000 89.7000 395.2500 ;
	    RECT 119.1000 395.1000 120.9000 395.2500 ;
	    RECT 171.9000 395.1000 173.7000 395.2500 ;
	    RECT 275.1000 396.7500 276.9000 396.9000 ;
	    RECT 287.1000 396.7500 288.9000 396.9000 ;
	    RECT 275.1000 395.2500 288.9000 396.7500 ;
	    RECT 275.1000 395.1000 276.9000 395.2500 ;
	    RECT 287.1000 395.1000 288.9000 395.2500 ;
	    RECT 805.5000 396.7500 807.3000 396.9000 ;
	    RECT 822.3000 396.7500 824.1000 396.9000 ;
	    RECT 805.5000 395.2500 824.1000 396.7500 ;
	    RECT 805.5000 395.1000 807.3000 395.2500 ;
	    RECT 822.3000 395.1000 824.1000 395.2500 ;
	    RECT 915.9000 396.7500 917.7000 396.9000 ;
	    RECT 966.3000 396.7500 968.1000 396.9000 ;
	    RECT 915.9000 395.2500 968.1000 396.7500 ;
	    RECT 915.9000 395.1000 917.7000 395.2500 ;
	    RECT 966.3000 395.1000 968.1000 395.2500 ;
	    RECT 1033.5000 396.7500 1035.3000 396.9000 ;
	    RECT 1081.5000 396.7500 1083.3000 396.9000 ;
	    RECT 1033.5000 395.2500 1083.3000 396.7500 ;
	    RECT 1033.5000 395.1000 1035.3000 395.2500 ;
	    RECT 1081.5000 395.1000 1083.3000 395.2500 ;
	    RECT 1153.5000 396.7500 1155.3000 396.9000 ;
	    RECT 1179.9000 396.7500 1181.7001 396.9000 ;
	    RECT 1153.5000 395.2500 1181.7001 396.7500 ;
	    RECT 1153.5000 395.1000 1155.3000 395.2500 ;
	    RECT 1179.9000 395.1000 1181.7001 395.2500 ;
	    RECT 1189.5000 396.7500 1191.3000 396.9000 ;
	    RECT 1244.7001 396.7500 1246.5000 396.9000 ;
	    RECT 1189.5000 395.2500 1246.5000 396.7500 ;
	    RECT 1189.5000 395.1000 1191.3000 395.2500 ;
	    RECT 1244.7001 395.1000 1246.5000 395.2500 ;
	    RECT 1316.7001 396.7500 1318.5000 396.9000 ;
	    RECT 1422.3000 396.7500 1424.1000 396.9000 ;
	    RECT 1482.3000 396.7500 1484.1000 396.9000 ;
	    RECT 1316.7001 395.2500 1484.1000 396.7500 ;
	    RECT 1316.7001 395.1000 1318.5000 395.2500 ;
	    RECT 1422.3000 395.1000 1424.1000 395.2500 ;
	    RECT 1482.3000 395.1000 1484.1000 395.2500 ;
	    RECT 1515.9000 396.7500 1517.7001 396.9000 ;
	    RECT 1551.9000 396.7500 1553.7001 396.9000 ;
	    RECT 1515.9000 395.2500 1553.7001 396.7500 ;
	    RECT 1515.9000 395.1000 1517.7001 395.2500 ;
	    RECT 1551.9000 395.1000 1553.7001 395.2500 ;
	    RECT 107.1000 390.7500 108.9000 390.9000 ;
	    RECT 159.9000 390.7500 161.7000 390.9000 ;
	    RECT 107.1000 389.2500 161.7000 390.7500 ;
	    RECT 107.1000 389.1000 108.9000 389.2500 ;
	    RECT 159.9000 389.1000 161.7000 389.2500 ;
	    RECT 289.5000 390.7500 291.3000 390.9000 ;
	    RECT 315.9000 390.7500 317.7000 390.9000 ;
	    RECT 337.5000 390.7500 339.3000 390.9000 ;
	    RECT 289.5000 389.2500 339.3000 390.7500 ;
	    RECT 289.5000 389.1000 291.3000 389.2500 ;
	    RECT 315.9000 389.1000 317.7000 389.2500 ;
	    RECT 337.5000 389.1000 339.3000 389.2500 ;
	    RECT 498.3000 390.7500 500.1000 390.9000 ;
	    RECT 507.9000 390.7500 509.7000 390.9000 ;
	    RECT 498.3000 389.2500 509.7000 390.7500 ;
	    RECT 498.3000 389.1000 500.1000 389.2500 ;
	    RECT 507.9000 389.1000 509.7000 389.2500 ;
	    RECT 680.7000 390.7500 682.5000 390.9000 ;
	    RECT 704.7000 390.7500 706.5000 390.9000 ;
	    RECT 680.7000 389.2500 706.5000 390.7500 ;
	    RECT 680.7000 389.1000 682.5000 389.2500 ;
	    RECT 704.7000 389.1000 706.5000 389.2500 ;
	    RECT 788.7000 390.7500 790.5000 390.9000 ;
	    RECT 839.1000 390.7500 840.9000 390.9000 ;
	    RECT 788.7000 389.2500 840.9000 390.7500 ;
	    RECT 788.7000 389.1000 790.5000 389.2500 ;
	    RECT 839.1000 389.1000 840.9000 389.2500 ;
	    RECT 983.1000 390.7500 984.9000 390.9000 ;
	    RECT 1014.3000 390.7500 1016.1000 390.9000 ;
	    RECT 983.1000 389.2500 1016.1000 390.7500 ;
	    RECT 983.1000 389.1000 984.9000 389.2500 ;
	    RECT 1014.3000 389.1000 1016.1000 389.2500 ;
	    RECT 1050.3000 390.7500 1052.1000 390.9000 ;
	    RECT 1119.9000 390.7500 1121.7001 390.9000 ;
	    RECT 1050.3000 389.2500 1121.7001 390.7500 ;
	    RECT 1050.3000 389.1000 1052.1000 389.2500 ;
	    RECT 1119.9000 389.1000 1121.7001 389.2500 ;
	    RECT 1184.7001 390.7500 1186.5000 390.9000 ;
	    RECT 1326.3000 390.7500 1328.1000 390.9000 ;
	    RECT 1184.7001 389.2500 1328.1000 390.7500 ;
	    RECT 1184.7001 389.1000 1186.5000 389.2500 ;
	    RECT 1326.3000 389.1000 1328.1000 389.2500 ;
	    RECT 1367.1000 390.7500 1368.9000 390.9000 ;
	    RECT 1405.5000 390.7500 1407.3000 390.9000 ;
	    RECT 1367.1000 389.2500 1407.3000 390.7500 ;
	    RECT 1367.1000 389.1000 1368.9000 389.2500 ;
	    RECT 1405.5000 389.1000 1407.3000 389.2500 ;
	    RECT 1515.9000 390.7500 1517.7001 390.9000 ;
	    RECT 1532.7001 390.7500 1534.5000 390.9000 ;
	    RECT 1515.9000 389.2500 1534.5000 390.7500 ;
	    RECT 1515.9000 389.1000 1517.7001 389.2500 ;
	    RECT 1532.7001 389.1000 1534.5000 389.2500 ;
	    RECT 63.9000 384.7500 65.7000 384.9000 ;
	    RECT 143.1000 384.7500 144.9000 384.9000 ;
	    RECT 63.9000 383.2500 144.9000 384.7500 ;
	    RECT 63.9000 383.1000 65.7000 383.2500 ;
	    RECT 143.1000 383.1000 144.9000 383.2500 ;
	    RECT 270.3000 384.7500 272.1000 384.9000 ;
	    RECT 303.9000 384.7500 305.7000 384.9000 ;
	    RECT 270.3000 383.2500 305.7000 384.7500 ;
	    RECT 270.3000 383.1000 272.1000 383.2500 ;
	    RECT 303.9000 383.1000 305.7000 383.2500 ;
	    RECT 402.3000 384.7500 404.1000 384.9000 ;
	    RECT 512.7000 384.7500 514.5000 384.9000 ;
	    RECT 402.3000 383.2500 514.5000 384.7500 ;
	    RECT 402.3000 383.1000 404.1000 383.2500 ;
	    RECT 512.7000 383.1000 514.5000 383.2500 ;
	    RECT 563.1000 384.7500 564.9000 384.9000 ;
	    RECT 599.1000 384.7500 600.9000 384.9000 ;
	    RECT 563.1000 383.2500 600.9000 384.7500 ;
	    RECT 563.1000 383.1000 564.9000 383.2500 ;
	    RECT 599.1000 383.1000 600.9000 383.2500 ;
	    RECT 798.3000 384.7500 800.1000 384.9000 ;
	    RECT 807.9000 384.7500 809.7000 384.9000 ;
	    RECT 834.3000 384.7500 836.1000 384.9000 ;
	    RECT 798.3000 383.2500 836.1000 384.7500 ;
	    RECT 798.3000 383.1000 800.1000 383.2500 ;
	    RECT 807.9000 383.1000 809.7000 383.2500 ;
	    RECT 834.3000 383.1000 836.1000 383.2500 ;
	    RECT 1093.5000 384.7500 1095.3000 384.9000 ;
	    RECT 1112.7001 384.7500 1114.5000 384.9000 ;
	    RECT 1093.5000 383.2500 1114.5000 384.7500 ;
	    RECT 1093.5000 383.1000 1095.3000 383.2500 ;
	    RECT 1112.7001 383.1000 1114.5000 383.2500 ;
	    RECT 1151.1000 384.7500 1152.9000 384.9000 ;
	    RECT 1158.3000 384.7500 1160.1000 384.9000 ;
	    RECT 1151.1000 383.2500 1160.1000 384.7500 ;
	    RECT 1151.1000 383.1000 1152.9000 383.2500 ;
	    RECT 1158.3000 383.1000 1160.1000 383.2500 ;
	    RECT 1191.9000 384.7500 1193.7001 384.9000 ;
	    RECT 1242.3000 384.7500 1244.1000 384.9000 ;
	    RECT 1191.9000 383.2500 1244.1000 384.7500 ;
	    RECT 1191.9000 383.1000 1193.7001 383.2500 ;
	    RECT 1242.3000 383.1000 1244.1000 383.2500 ;
	    RECT 1316.7001 384.7500 1318.5000 384.9000 ;
	    RECT 1328.7001 384.7500 1330.5000 384.9000 ;
	    RECT 1316.7001 383.2500 1330.5000 384.7500 ;
	    RECT 1316.7001 383.1000 1318.5000 383.2500 ;
	    RECT 1328.7001 383.1000 1330.5000 383.2500 ;
	    RECT 191.1000 378.7500 192.9000 378.9000 ;
	    RECT 198.3000 378.7500 200.1000 378.9000 ;
	    RECT 191.1000 377.2500 200.1000 378.7500 ;
	    RECT 191.1000 377.1000 192.9000 377.2500 ;
	    RECT 198.3000 377.1000 200.1000 377.2500 ;
	    RECT 246.3000 378.7500 248.1000 378.9000 ;
	    RECT 272.7000 378.7500 274.5000 378.9000 ;
	    RECT 301.5000 378.7500 303.3000 378.9000 ;
	    RECT 342.3000 378.7500 344.1000 378.9000 ;
	    RECT 246.3000 377.2500 344.1000 378.7500 ;
	    RECT 246.3000 377.1000 248.1000 377.2500 ;
	    RECT 272.7000 377.1000 274.5000 377.2500 ;
	    RECT 301.5000 377.1000 303.3000 377.2500 ;
	    RECT 342.3000 377.1000 344.1000 377.2500 ;
	    RECT 822.3000 378.7500 824.1000 378.9000 ;
	    RECT 855.9000 378.7500 857.7000 378.9000 ;
	    RECT 822.3000 377.2500 857.7000 378.7500 ;
	    RECT 822.3000 377.1000 824.1000 377.2500 ;
	    RECT 855.9000 377.1000 857.7000 377.2500 ;
	    RECT 1158.3000 378.7500 1160.1000 378.9000 ;
	    RECT 1424.7001 378.7500 1426.5000 378.9000 ;
	    RECT 1434.3000 378.7500 1436.1000 378.9000 ;
	    RECT 1487.1000 378.7500 1488.9000 378.9000 ;
	    RECT 1158.3000 377.2500 1488.9000 378.7500 ;
	    RECT 1158.3000 377.1000 1160.1000 377.2500 ;
	    RECT 1424.7001 377.1000 1426.5000 377.2500 ;
	    RECT 1434.3000 377.1000 1436.1000 377.2500 ;
	    RECT 1487.1000 377.1000 1488.9000 377.2500 ;
	    RECT 1496.7001 378.7500 1498.5000 378.9000 ;
	    RECT 1535.1000 378.7500 1536.9000 378.9000 ;
	    RECT 1496.7001 377.2500 1536.9000 378.7500 ;
	    RECT 1496.7001 377.1000 1498.5000 377.2500 ;
	    RECT 1535.1000 377.1000 1536.9000 377.2500 ;
	    RECT 603.9000 372.7500 605.7000 372.9000 ;
	    RECT 671.1000 372.7500 672.9000 372.9000 ;
	    RECT 603.9000 371.2500 672.9000 372.7500 ;
	    RECT 603.9000 371.1000 605.7000 371.2500 ;
	    RECT 671.1000 371.1000 672.9000 371.2500 ;
	    RECT 1093.5000 372.7500 1095.3000 372.9000 ;
	    RECT 1105.5000 372.7500 1107.3000 372.9000 ;
	    RECT 1093.5000 371.2500 1107.3000 372.7500 ;
	    RECT 1093.5000 371.1000 1095.3000 371.2500 ;
	    RECT 1105.5000 371.1000 1107.3000 371.2500 ;
	    RECT 1146.3000 372.7500 1148.1000 372.9000 ;
	    RECT 1175.1000 372.7500 1176.9000 372.9000 ;
	    RECT 1146.3000 371.2500 1176.9000 372.7500 ;
	    RECT 1146.3000 371.1000 1148.1000 371.2500 ;
	    RECT 1175.1000 371.1000 1176.9000 371.2500 ;
	    RECT 1326.3000 372.7500 1328.1000 372.9000 ;
	    RECT 1439.1000 372.7500 1440.9000 372.9000 ;
	    RECT 1326.3000 371.2500 1440.9000 372.7500 ;
	    RECT 1326.3000 371.1000 1328.1000 371.2500 ;
	    RECT 1439.1000 371.1000 1440.9000 371.2500 ;
	    RECT 1513.5000 372.7500 1515.3000 372.9000 ;
	    RECT 1537.5000 372.7500 1539.3000 372.9000 ;
	    RECT 1513.5000 371.2500 1539.3000 372.7500 ;
	    RECT 1513.5000 371.1000 1515.3000 371.2500 ;
	    RECT 1537.5000 371.1000 1539.3000 371.2500 ;
	    RECT 227.1000 366.7500 228.9000 366.9000 ;
	    RECT 255.9000 366.7500 257.7000 366.9000 ;
	    RECT 227.1000 365.2500 257.7000 366.7500 ;
	    RECT 227.1000 365.1000 228.9000 365.2500 ;
	    RECT 255.9000 365.1000 257.7000 365.2500 ;
	    RECT 315.9000 366.7500 317.7000 366.9000 ;
	    RECT 349.5000 366.7500 351.3000 366.9000 ;
	    RECT 315.9000 365.2500 351.3000 366.7500 ;
	    RECT 315.9000 365.1000 317.7000 365.2500 ;
	    RECT 349.5000 365.1000 351.3000 365.2500 ;
	    RECT 601.5000 366.7500 603.3000 366.9000 ;
	    RECT 956.7000 366.7500 958.5000 366.9000 ;
	    RECT 601.5000 365.2500 958.5000 366.7500 ;
	    RECT 601.5000 365.1000 603.3000 365.2500 ;
	    RECT 956.7000 365.1000 958.5000 365.2500 ;
	    RECT 990.3000 366.7500 992.1000 366.9000 ;
	    RECT 1038.3000 366.7500 1040.1000 366.9000 ;
	    RECT 990.3000 365.2500 1040.1000 366.7500 ;
	    RECT 990.3000 365.1000 992.1000 365.2500 ;
	    RECT 1038.3000 365.1000 1040.1000 365.2500 ;
	    RECT 1273.5000 366.7500 1275.3000 366.9000 ;
	    RECT 1319.1000 366.7500 1320.9000 366.9000 ;
	    RECT 1273.5000 365.2500 1320.9000 366.7500 ;
	    RECT 1273.5000 365.1000 1275.3000 365.2500 ;
	    RECT 1319.1000 365.1000 1320.9000 365.2500 ;
	    RECT 1472.7001 366.7500 1474.5000 366.9000 ;
	    RECT 1496.7001 366.7500 1498.5000 366.9000 ;
	    RECT 1472.7001 365.2500 1498.5000 366.7500 ;
	    RECT 1472.7001 365.1000 1474.5000 365.2500 ;
	    RECT 1496.7001 365.1000 1498.5000 365.2500 ;
	    RECT 13.5000 360.7500 15.3000 360.9000 ;
	    RECT 39.9000 360.7500 41.7000 360.9000 ;
	    RECT 13.5000 359.2500 41.7000 360.7500 ;
	    RECT 13.5000 359.1000 15.3000 359.2500 ;
	    RECT 39.9000 359.1000 41.7000 359.2500 ;
	    RECT 159.9000 360.7500 161.7000 360.9000 ;
	    RECT 174.3000 360.7500 176.1000 360.9000 ;
	    RECT 159.9000 359.2500 176.1000 360.7500 ;
	    RECT 159.9000 359.1000 161.7000 359.2500 ;
	    RECT 174.3000 359.1000 176.1000 359.2500 ;
	    RECT 853.5000 360.7500 855.3000 360.9000 ;
	    RECT 858.3000 360.7500 860.1000 360.9000 ;
	    RECT 853.5000 359.2500 860.1000 360.7500 ;
	    RECT 853.5000 359.1000 855.3000 359.2500 ;
	    RECT 858.3000 359.1000 860.1000 359.2500 ;
	    RECT 1019.1000 360.7500 1020.9000 360.9000 ;
	    RECT 1033.5000 360.7500 1035.3000 360.9000 ;
	    RECT 1019.1000 359.2500 1035.3000 360.7500 ;
	    RECT 1019.1000 359.1000 1020.9000 359.2500 ;
	    RECT 1033.5000 359.1000 1035.3000 359.2500 ;
	    RECT 1059.9000 360.7500 1061.7001 360.9000 ;
	    RECT 1091.1000 360.7500 1092.9000 360.9000 ;
	    RECT 1119.9000 360.7500 1121.7001 360.9000 ;
	    RECT 1059.9000 359.2500 1121.7001 360.7500 ;
	    RECT 1059.9000 359.1000 1061.7001 359.2500 ;
	    RECT 1091.1000 359.1000 1092.9000 359.2500 ;
	    RECT 1119.9000 359.1000 1121.7001 359.2500 ;
	    RECT 1151.1000 360.7500 1152.9000 360.9000 ;
	    RECT 1165.5000 360.7500 1167.3000 360.9000 ;
	    RECT 1151.1000 359.2500 1167.3000 360.7500 ;
	    RECT 1151.1000 359.1000 1152.9000 359.2500 ;
	    RECT 1165.5000 359.1000 1167.3000 359.2500 ;
	    RECT 1266.3000 360.7500 1268.1000 360.9000 ;
	    RECT 1338.3000 360.7500 1340.1000 360.9000 ;
	    RECT 1266.3000 359.2500 1340.1000 360.7500 ;
	    RECT 1266.3000 359.1000 1268.1000 359.2500 ;
	    RECT 1338.3000 359.1000 1340.1000 359.2500 ;
	    RECT 1405.5000 360.7500 1407.3000 360.9000 ;
	    RECT 1431.9000 360.7500 1433.7001 360.9000 ;
	    RECT 1405.5000 359.2500 1433.7001 360.7500 ;
	    RECT 1405.5000 359.1000 1407.3000 359.2500 ;
	    RECT 1431.9000 359.1000 1433.7001 359.2500 ;
	    RECT 1491.9000 360.7500 1493.7001 360.9000 ;
	    RECT 1532.7001 360.7500 1534.5000 360.9000 ;
	    RECT 1491.9000 359.2500 1534.5000 360.7500 ;
	    RECT 1491.9000 359.1000 1493.7001 359.2500 ;
	    RECT 1532.7001 359.1000 1534.5000 359.2500 ;
	    RECT 431.1000 354.7500 432.9000 354.9000 ;
	    RECT 507.9000 354.7500 509.7000 354.9000 ;
	    RECT 563.1000 354.7500 564.9000 354.9000 ;
	    RECT 431.1000 353.2500 564.9000 354.7500 ;
	    RECT 431.1000 353.1000 432.9000 353.2500 ;
	    RECT 507.9000 353.1000 509.7000 353.2500 ;
	    RECT 563.1000 353.1000 564.9000 353.2500 ;
	    RECT 647.1000 354.7500 648.9000 354.9000 ;
	    RECT 654.3000 354.7500 656.1000 354.9000 ;
	    RECT 647.1000 353.2500 656.1000 354.7500 ;
	    RECT 647.1000 353.1000 648.9000 353.2500 ;
	    RECT 654.3000 353.1000 656.1000 353.2500 ;
	    RECT 805.5000 354.7500 807.3000 354.9000 ;
	    RECT 827.1000 354.7500 828.9000 354.9000 ;
	    RECT 805.5000 353.2500 828.9000 354.7500 ;
	    RECT 805.5000 353.1000 807.3000 353.2500 ;
	    RECT 827.1000 353.1000 828.9000 353.2500 ;
	    RECT 1285.5000 354.7500 1287.3000 354.9000 ;
	    RECT 1335.9000 354.7500 1337.7001 354.9000 ;
	    RECT 1285.5000 353.2500 1337.7001 354.7500 ;
	    RECT 1285.5000 353.1000 1287.3000 353.2500 ;
	    RECT 1335.9000 353.1000 1337.7001 353.2500 ;
	    RECT 1537.5000 354.7500 1539.3000 354.9000 ;
	    RECT 1561.5000 354.7500 1563.3000 354.9000 ;
	    RECT 1537.5000 353.2500 1563.3000 354.7500 ;
	    RECT 1537.5000 353.1000 1539.3000 353.2500 ;
	    RECT 1561.5000 353.1000 1563.3000 353.2500 ;
	    RECT 23.1000 348.7500 24.9000 348.9000 ;
	    RECT 66.3000 348.7500 68.1000 348.9000 ;
	    RECT 318.3000 348.7500 320.1000 348.9000 ;
	    RECT 23.1000 347.2500 320.1000 348.7500 ;
	    RECT 23.1000 347.1000 24.9000 347.2500 ;
	    RECT 66.3000 347.1000 68.1000 347.2500 ;
	    RECT 318.3000 347.1000 320.1000 347.2500 ;
	    RECT 383.1000 348.7500 384.9000 348.9000 ;
	    RECT 390.3000 348.7500 392.1000 348.9000 ;
	    RECT 383.1000 347.2500 392.1000 348.7500 ;
	    RECT 383.1000 347.1000 384.9000 347.2500 ;
	    RECT 390.3000 347.1000 392.1000 347.2500 ;
	    RECT 428.7000 348.7500 430.5000 348.9000 ;
	    RECT 474.3000 348.7500 476.1000 348.9000 ;
	    RECT 428.7000 347.2500 476.1000 348.7500 ;
	    RECT 428.7000 347.1000 430.5000 347.2500 ;
	    RECT 474.3000 347.1000 476.1000 347.2500 ;
	    RECT 642.3000 348.7500 644.1000 348.9000 ;
	    RECT 714.3000 348.7500 716.1000 348.9000 ;
	    RECT 642.3000 347.2500 716.1000 348.7500 ;
	    RECT 642.3000 347.1000 644.1000 347.2500 ;
	    RECT 714.3000 347.1000 716.1000 347.2500 ;
	    RECT 1081.5000 348.7500 1083.3000 348.9000 ;
	    RECT 1115.1000 348.7500 1116.9000 348.9000 ;
	    RECT 1136.7001 348.7500 1138.5000 348.9000 ;
	    RECT 1153.5000 348.7500 1155.3000 348.9000 ;
	    RECT 1081.5000 347.2500 1155.3000 348.7500 ;
	    RECT 1081.5000 347.1000 1083.3000 347.2500 ;
	    RECT 1115.1000 347.1000 1116.9000 347.2500 ;
	    RECT 1136.7001 347.1000 1138.5000 347.2500 ;
	    RECT 1153.5000 347.1000 1155.3000 347.2500 ;
	    RECT 1458.3000 348.7500 1460.1000 348.9000 ;
	    RECT 1470.3000 348.7500 1472.1000 348.9000 ;
	    RECT 1458.3000 347.2500 1472.1000 348.7500 ;
	    RECT 1458.3000 347.1000 1460.1000 347.2500 ;
	    RECT 1470.3000 347.1000 1472.1000 347.2500 ;
	    RECT 25.5000 342.7500 27.3000 342.9000 ;
	    RECT 47.1000 342.7500 48.9000 342.9000 ;
	    RECT 66.3000 342.7500 68.1000 342.9000 ;
	    RECT 71.1000 342.7500 72.9000 342.9000 ;
	    RECT 25.5000 341.2500 72.9000 342.7500 ;
	    RECT 25.5000 341.1000 27.3000 341.2500 ;
	    RECT 47.1000 341.1000 48.9000 341.2500 ;
	    RECT 66.3000 341.1000 68.1000 341.2500 ;
	    RECT 71.1000 341.1000 72.9000 341.2500 ;
	    RECT 111.9000 342.7500 113.7000 342.9000 ;
	    RECT 119.1000 342.7500 120.9000 342.9000 ;
	    RECT 111.9000 341.2500 120.9000 342.7500 ;
	    RECT 111.9000 341.1000 113.7000 341.2500 ;
	    RECT 119.1000 341.1000 120.9000 341.2500 ;
	    RECT 138.3000 342.7500 140.1000 342.9000 ;
	    RECT 167.1000 342.7500 168.9000 342.9000 ;
	    RECT 186.3000 342.7500 188.1000 342.9000 ;
	    RECT 138.3000 341.2500 188.1000 342.7500 ;
	    RECT 138.3000 341.1000 140.1000 341.2500 ;
	    RECT 167.1000 341.1000 168.9000 341.2500 ;
	    RECT 186.3000 341.1000 188.1000 341.2500 ;
	    RECT 380.7000 342.7500 382.5000 342.9000 ;
	    RECT 387.9000 342.7500 389.7000 342.9000 ;
	    RECT 380.7000 341.2500 389.7000 342.7500 ;
	    RECT 380.7000 341.1000 382.5000 341.2500 ;
	    RECT 387.9000 341.1000 389.7000 341.2500 ;
	    RECT 421.5000 342.7500 423.3000 342.9000 ;
	    RECT 445.5000 342.7500 447.3000 342.9000 ;
	    RECT 421.5000 341.2500 447.3000 342.7500 ;
	    RECT 421.5000 341.1000 423.3000 341.2500 ;
	    RECT 445.5000 341.1000 447.3000 341.2500 ;
	    RECT 579.9000 342.7500 581.7000 342.9000 ;
	    RECT 632.7000 342.7500 634.5000 342.9000 ;
	    RECT 579.9000 341.2500 634.5000 342.7500 ;
	    RECT 579.9000 341.1000 581.7000 341.2500 ;
	    RECT 632.7000 341.1000 634.5000 341.2500 ;
	    RECT 875.1000 342.7500 876.9000 342.9000 ;
	    RECT 882.3000 342.7500 884.1000 342.9000 ;
	    RECT 875.1000 341.2500 884.1000 342.7500 ;
	    RECT 875.1000 341.1000 876.9000 341.2500 ;
	    RECT 882.3000 341.1000 884.1000 341.2500 ;
	    RECT 1208.7001 342.7500 1210.5000 342.9000 ;
	    RECT 1220.7001 342.7500 1222.5000 342.9000 ;
	    RECT 1208.7001 341.2500 1222.5000 342.7500 ;
	    RECT 1208.7001 341.1000 1210.5000 341.2500 ;
	    RECT 1220.7001 341.1000 1222.5000 341.2500 ;
	    RECT 1309.5000 342.7500 1311.3000 342.9000 ;
	    RECT 1333.5000 342.7500 1335.3000 342.9000 ;
	    RECT 1309.5000 341.2500 1335.3000 342.7500 ;
	    RECT 1309.5000 341.1000 1311.3000 341.2500 ;
	    RECT 1333.5000 341.1000 1335.3000 341.2500 ;
	    RECT 1350.3000 342.7500 1352.1000 342.9000 ;
	    RECT 1381.5000 342.7500 1383.3000 342.9000 ;
	    RECT 1350.3000 341.2500 1383.3000 342.7500 ;
	    RECT 1350.3000 341.1000 1352.1000 341.2500 ;
	    RECT 1381.5000 341.1000 1383.3000 341.2500 ;
	    RECT 1451.1000 342.7500 1452.9000 342.9000 ;
	    RECT 1463.1000 342.7500 1464.9000 342.9000 ;
	    RECT 1451.1000 341.2500 1464.9000 342.7500 ;
	    RECT 1451.1000 341.1000 1452.9000 341.2500 ;
	    RECT 1463.1000 341.1000 1464.9000 341.2500 ;
	    RECT 71.1000 336.7500 72.9000 336.9000 ;
	    RECT 109.5000 336.7500 111.3000 336.9000 ;
	    RECT 138.3000 336.7500 140.1000 336.9000 ;
	    RECT 71.1000 335.2500 140.1000 336.7500 ;
	    RECT 71.1000 335.1000 72.9000 335.2500 ;
	    RECT 109.5000 335.1000 111.3000 335.2500 ;
	    RECT 138.3000 335.1000 140.1000 335.2500 ;
	    RECT 193.5000 336.7500 195.3000 336.9000 ;
	    RECT 198.3000 336.7500 200.1000 336.9000 ;
	    RECT 193.5000 335.2500 200.1000 336.7500 ;
	    RECT 193.5000 335.1000 195.3000 335.2500 ;
	    RECT 198.3000 335.1000 200.1000 335.2500 ;
	    RECT 407.1000 336.7500 408.9000 336.9000 ;
	    RECT 440.7000 336.7500 442.5000 336.9000 ;
	    RECT 407.1000 335.2500 442.5000 336.7500 ;
	    RECT 407.1000 335.1000 408.9000 335.2500 ;
	    RECT 440.7000 335.1000 442.5000 335.2500 ;
	    RECT 589.5000 336.7500 591.3000 336.9000 ;
	    RECT 671.1000 336.7500 672.9000 336.9000 ;
	    RECT 589.5000 335.2500 672.9000 336.7500 ;
	    RECT 589.5000 335.1000 591.3000 335.2500 ;
	    RECT 671.1000 335.1000 672.9000 335.2500 ;
	    RECT 1088.7001 336.7500 1090.5000 336.9000 ;
	    RECT 1134.3000 336.7500 1136.1000 336.9000 ;
	    RECT 1175.1000 336.7500 1176.9000 336.9000 ;
	    RECT 1088.7001 335.2500 1176.9000 336.7500 ;
	    RECT 1088.7001 335.1000 1090.5000 335.2500 ;
	    RECT 1134.3000 335.1000 1136.1000 335.2500 ;
	    RECT 1175.1000 335.1000 1176.9000 335.2500 ;
	    RECT 1225.5000 336.7500 1227.3000 336.9000 ;
	    RECT 1263.9000 336.7500 1265.7001 336.9000 ;
	    RECT 1225.5000 335.2500 1265.7001 336.7500 ;
	    RECT 1225.5000 335.1000 1227.3000 335.2500 ;
	    RECT 1263.9000 335.1000 1265.7001 335.2500 ;
	    RECT 1271.1000 336.7500 1272.9000 336.9000 ;
	    RECT 1395.9000 336.7500 1397.7001 336.9000 ;
	    RECT 1405.5000 336.7500 1407.3000 336.9000 ;
	    RECT 1271.1000 335.2500 1407.3000 336.7500 ;
	    RECT 1271.1000 335.1000 1272.9000 335.2500 ;
	    RECT 1395.9000 335.1000 1397.7001 335.2500 ;
	    RECT 1405.5000 335.1000 1407.3000 335.2500 ;
	    RECT 1417.5000 336.7500 1419.3000 336.9000 ;
	    RECT 1491.9000 336.7500 1493.7001 336.9000 ;
	    RECT 1417.5000 335.2500 1493.7001 336.7500 ;
	    RECT 1417.5000 335.1000 1419.3000 335.2500 ;
	    RECT 1491.9000 335.1000 1493.7001 335.2500 ;
	    RECT 63.9000 330.7500 65.7000 330.9000 ;
	    RECT 73.5000 330.7500 75.3000 330.9000 ;
	    RECT 63.9000 329.2500 75.3000 330.7500 ;
	    RECT 63.9000 329.1000 65.7000 329.2500 ;
	    RECT 73.5000 329.1000 75.3000 329.2500 ;
	    RECT 143.1000 330.7500 144.9000 330.9000 ;
	    RECT 229.5000 330.7500 231.3000 330.9000 ;
	    RECT 143.1000 329.2500 231.3000 330.7500 ;
	    RECT 143.1000 329.1000 144.9000 329.2500 ;
	    RECT 229.5000 329.1000 231.3000 329.2500 ;
	    RECT 383.1000 330.7500 384.9000 330.9000 ;
	    RECT 421.5000 330.7500 423.3000 330.9000 ;
	    RECT 383.1000 329.2500 423.3000 330.7500 ;
	    RECT 383.1000 329.1000 384.9000 329.2500 ;
	    RECT 421.5000 329.1000 423.3000 329.2500 ;
	    RECT 563.1000 330.7500 564.9000 330.9000 ;
	    RECT 663.9000 330.7500 665.7000 330.9000 ;
	    RECT 699.9000 330.7500 701.7000 330.9000 ;
	    RECT 563.1000 329.2500 701.7000 330.7500 ;
	    RECT 563.1000 329.1000 564.9000 329.2500 ;
	    RECT 663.9000 329.1000 665.7000 329.2500 ;
	    RECT 699.9000 329.1000 701.7000 329.2500 ;
	    RECT 942.3000 330.7500 944.1000 330.9000 ;
	    RECT 980.7000 330.7500 982.5000 330.9000 ;
	    RECT 942.3000 329.2500 982.5000 330.7500 ;
	    RECT 942.3000 329.1000 944.1000 329.2500 ;
	    RECT 980.7000 329.1000 982.5000 329.2500 ;
	    RECT 1038.3000 330.7500 1040.1000 330.9000 ;
	    RECT 1076.7001 330.7500 1078.5000 330.9000 ;
	    RECT 1038.3000 329.2500 1078.5000 330.7500 ;
	    RECT 1038.3000 329.1000 1040.1000 329.2500 ;
	    RECT 1076.7001 329.1000 1078.5000 329.2500 ;
	    RECT 1129.5000 330.7500 1131.3000 330.9000 ;
	    RECT 1167.9000 330.7500 1169.7001 330.9000 ;
	    RECT 1129.5000 329.2500 1169.7001 330.7500 ;
	    RECT 1129.5000 329.1000 1131.3000 329.2500 ;
	    RECT 1167.9000 329.1000 1169.7001 329.2500 ;
	    RECT 1177.5000 330.7500 1179.3000 330.9000 ;
	    RECT 1215.9000 330.7500 1217.7001 330.9000 ;
	    RECT 1177.5000 329.2500 1217.7001 330.7500 ;
	    RECT 1177.5000 329.1000 1179.3000 329.2500 ;
	    RECT 1215.9000 329.1000 1217.7001 329.2500 ;
	    RECT 1223.1000 330.7500 1224.9000 330.9000 ;
	    RECT 1278.3000 330.7500 1280.1000 330.9000 ;
	    RECT 1223.1000 329.2500 1280.1000 330.7500 ;
	    RECT 1223.1000 329.1000 1224.9000 329.2500 ;
	    RECT 1278.3000 329.1000 1280.1000 329.2500 ;
	    RECT 1290.3000 330.7500 1292.1000 330.9000 ;
	    RECT 1309.5000 330.7500 1311.3000 330.9000 ;
	    RECT 1290.3000 329.2500 1311.3000 330.7500 ;
	    RECT 1290.3000 329.1000 1292.1000 329.2500 ;
	    RECT 1309.5000 329.1000 1311.3000 329.2500 ;
	    RECT 1319.1000 330.7500 1320.9000 330.9000 ;
	    RECT 1347.9000 330.7500 1349.7001 330.9000 ;
	    RECT 1319.1000 329.2500 1349.7001 330.7500 ;
	    RECT 1319.1000 329.1000 1320.9000 329.2500 ;
	    RECT 1347.9000 329.1000 1349.7001 329.2500 ;
	    RECT 1391.1000 330.7500 1392.9000 330.9000 ;
	    RECT 1441.5000 330.7500 1443.3000 330.9000 ;
	    RECT 1391.1000 329.2500 1443.3000 330.7500 ;
	    RECT 1391.1000 329.1000 1392.9000 329.2500 ;
	    RECT 1441.5000 329.1000 1443.3000 329.2500 ;
	    RECT 1539.9000 330.7500 1541.7001 330.9000 ;
	    RECT 1561.5000 330.7500 1563.3000 330.9000 ;
	    RECT 1539.9000 329.2500 1563.3000 330.7500 ;
	    RECT 1539.9000 329.1000 1541.7001 329.2500 ;
	    RECT 1561.5000 329.1000 1563.3000 329.2500 ;
	    RECT 157.5000 324.7500 159.3000 324.9000 ;
	    RECT 164.7000 324.7500 166.5000 324.9000 ;
	    RECT 174.3000 324.7500 176.1000 324.9000 ;
	    RECT 157.5000 323.2500 176.1000 324.7500 ;
	    RECT 157.5000 323.1000 159.3000 323.2500 ;
	    RECT 164.7000 323.1000 166.5000 323.2500 ;
	    RECT 174.3000 323.1000 176.1000 323.2500 ;
	    RECT 239.1000 324.7500 240.9000 324.9000 ;
	    RECT 272.7000 324.7500 274.5000 324.9000 ;
	    RECT 239.1000 323.2500 274.5000 324.7500 ;
	    RECT 239.1000 323.1000 240.9000 323.2500 ;
	    RECT 272.7000 323.1000 274.5000 323.2500 ;
	    RECT 435.9000 324.7500 437.7000 324.9000 ;
	    RECT 445.5000 324.7500 447.3000 324.9000 ;
	    RECT 435.9000 323.2500 447.3000 324.7500 ;
	    RECT 435.9000 323.1000 437.7000 323.2500 ;
	    RECT 445.5000 323.1000 447.3000 323.2500 ;
	    RECT 527.1000 324.7500 528.9000 324.9000 ;
	    RECT 534.3000 324.7500 536.1000 324.9000 ;
	    RECT 527.1000 323.2500 536.1000 324.7500 ;
	    RECT 527.1000 323.1000 528.9000 323.2500 ;
	    RECT 534.3000 323.1000 536.1000 323.2500 ;
	    RECT 831.9000 324.7500 833.7000 324.9000 ;
	    RECT 942.3000 324.7500 944.1000 324.9000 ;
	    RECT 831.9000 323.2500 944.1000 324.7500 ;
	    RECT 831.9000 323.1000 833.7000 323.2500 ;
	    RECT 942.3000 323.1000 944.1000 323.2500 ;
	    RECT 997.5000 324.7500 999.3000 324.9000 ;
	    RECT 1040.7001 324.7500 1042.5000 324.9000 ;
	    RECT 997.5000 323.2500 1042.5000 324.7500 ;
	    RECT 997.5000 323.1000 999.3000 323.2500 ;
	    RECT 1040.7001 323.1000 1042.5000 323.2500 ;
	    RECT 1083.9000 324.7500 1085.7001 324.9000 ;
	    RECT 1100.7001 324.7500 1102.5000 324.9000 ;
	    RECT 1083.9000 323.2500 1102.5000 324.7500 ;
	    RECT 1083.9000 323.1000 1085.7001 323.2500 ;
	    RECT 1100.7001 323.1000 1102.5000 323.2500 ;
	    RECT 1158.3000 324.7500 1160.1000 324.9000 ;
	    RECT 1213.5000 324.7500 1215.3000 324.9000 ;
	    RECT 1239.9000 324.7500 1241.7001 324.9000 ;
	    RECT 1158.3000 323.2500 1241.7001 324.7500 ;
	    RECT 1158.3000 323.1000 1160.1000 323.2500 ;
	    RECT 1213.5000 323.1000 1215.3000 323.2500 ;
	    RECT 1239.9000 323.1000 1241.7001 323.2500 ;
	    RECT 1299.9000 324.7500 1301.7001 324.9000 ;
	    RECT 1364.7001 324.7500 1366.5000 324.9000 ;
	    RECT 1299.9000 323.2500 1366.5000 324.7500 ;
	    RECT 1299.9000 323.1000 1301.7001 323.2500 ;
	    RECT 1364.7001 323.1000 1366.5000 323.2500 ;
	    RECT 27.9000 318.7500 29.7000 318.9000 ;
	    RECT 35.1000 318.7500 36.9000 318.9000 ;
	    RECT 27.9000 317.2500 36.9000 318.7500 ;
	    RECT 27.9000 317.1000 29.7000 317.2500 ;
	    RECT 35.1000 317.1000 36.9000 317.2500 ;
	    RECT 39.9000 318.7500 41.7000 318.9000 ;
	    RECT 47.1000 318.7500 48.9000 318.9000 ;
	    RECT 39.9000 317.2500 48.9000 318.7500 ;
	    RECT 39.9000 317.1000 41.7000 317.2500 ;
	    RECT 47.1000 317.1000 48.9000 317.2500 ;
	    RECT 73.5000 318.7500 75.3000 318.9000 ;
	    RECT 90.3000 318.7500 92.1000 318.9000 ;
	    RECT 73.5000 317.2500 92.1000 318.7500 ;
	    RECT 73.5000 317.1000 75.3000 317.2500 ;
	    RECT 90.3000 317.1000 92.1000 317.2500 ;
	    RECT 445.5000 318.7500 447.3000 318.9000 ;
	    RECT 457.5000 318.7500 459.3000 318.9000 ;
	    RECT 445.5000 317.2500 459.3000 318.7500 ;
	    RECT 445.5000 317.1000 447.3000 317.2500 ;
	    RECT 457.5000 317.1000 459.3000 317.2500 ;
	    RECT 915.9000 318.7500 917.7000 318.9000 ;
	    RECT 947.1000 318.7500 948.9000 318.9000 ;
	    RECT 915.9000 317.2500 948.9000 318.7500 ;
	    RECT 915.9000 317.1000 917.7000 317.2500 ;
	    RECT 947.1000 317.1000 948.9000 317.2500 ;
	    RECT 1004.7000 318.7500 1006.5000 318.9000 ;
	    RECT 1038.3000 318.7500 1040.1000 318.9000 ;
	    RECT 1004.7000 317.2500 1040.1000 318.7500 ;
	    RECT 1004.7000 317.1000 1006.5000 317.2500 ;
	    RECT 1038.3000 317.1000 1040.1000 317.2500 ;
	    RECT 1069.5000 318.7500 1071.3000 318.9000 ;
	    RECT 1081.5000 318.7500 1083.3000 318.9000 ;
	    RECT 1069.5000 317.2500 1083.3000 318.7500 ;
	    RECT 1069.5000 317.1000 1071.3000 317.2500 ;
	    RECT 1081.5000 317.1000 1083.3000 317.2500 ;
	    RECT 1160.7001 318.7500 1162.5000 318.9000 ;
	    RECT 1170.3000 318.7500 1172.1000 318.9000 ;
	    RECT 1160.7001 317.2500 1172.1000 318.7500 ;
	    RECT 1160.7001 317.1000 1162.5000 317.2500 ;
	    RECT 1170.3000 317.1000 1172.1000 317.2500 ;
	    RECT 1295.1000 318.7500 1296.9000 318.9000 ;
	    RECT 1304.7001 318.7500 1306.5000 318.9000 ;
	    RECT 1364.7001 318.7500 1366.5000 318.9000 ;
	    RECT 1295.1000 317.2500 1366.5000 318.7500 ;
	    RECT 1295.1000 317.1000 1296.9000 317.2500 ;
	    RECT 1304.7001 317.1000 1306.5000 317.2500 ;
	    RECT 1364.7001 317.1000 1366.5000 317.2500 ;
	    RECT 1388.7001 318.7500 1390.5000 318.9000 ;
	    RECT 1400.7001 318.7500 1402.5000 318.9000 ;
	    RECT 1388.7001 317.2500 1402.5000 318.7500 ;
	    RECT 1388.7001 317.1000 1390.5000 317.2500 ;
	    RECT 1400.7001 317.1000 1402.5000 317.2500 ;
	    RECT 1427.1000 318.7500 1428.9000 318.9000 ;
	    RECT 1446.3000 318.7500 1448.1000 318.9000 ;
	    RECT 1427.1000 317.2500 1448.1000 318.7500 ;
	    RECT 1427.1000 317.1000 1428.9000 317.2500 ;
	    RECT 1446.3000 317.1000 1448.1000 317.2500 ;
	    RECT 923.1000 312.7500 924.9000 312.9000 ;
	    RECT 961.5000 312.7500 963.3000 312.9000 ;
	    RECT 923.1000 311.2500 963.3000 312.7500 ;
	    RECT 923.1000 311.1000 924.9000 311.2500 ;
	    RECT 961.5000 311.1000 963.3000 311.2500 ;
	    RECT 1112.7001 312.7500 1114.5000 312.9000 ;
	    RECT 1232.7001 312.7500 1234.5000 312.9000 ;
	    RECT 1259.1000 312.7500 1260.9000 312.9000 ;
	    RECT 1275.9000 312.7500 1277.7001 312.9000 ;
	    RECT 1112.7001 311.2500 1277.7001 312.7500 ;
	    RECT 1112.7001 311.1000 1114.5000 311.2500 ;
	    RECT 1232.7001 311.1000 1234.5000 311.2500 ;
	    RECT 1259.1000 311.1000 1260.9000 311.2500 ;
	    RECT 1275.9000 311.1000 1277.7001 311.2500 ;
	    RECT 1285.5000 312.7500 1287.3000 312.9000 ;
	    RECT 1309.5000 312.7500 1311.3000 312.9000 ;
	    RECT 1285.5000 311.2500 1311.3000 312.7500 ;
	    RECT 1285.5000 311.1000 1287.3000 311.2500 ;
	    RECT 1309.5000 311.1000 1311.3000 311.2500 ;
	    RECT 1429.5000 312.7500 1431.3000 312.9000 ;
	    RECT 1436.7001 312.7500 1438.5000 312.9000 ;
	    RECT 1429.5000 311.2500 1438.5000 312.7500 ;
	    RECT 1429.5000 311.1000 1431.3000 311.2500 ;
	    RECT 1436.7001 311.1000 1438.5000 311.2500 ;
	    RECT 1453.5000 312.7500 1455.3000 312.9000 ;
	    RECT 1458.3000 312.7500 1460.1000 312.9000 ;
	    RECT 1453.5000 311.2500 1460.1000 312.7500 ;
	    RECT 1453.5000 311.1000 1455.3000 311.2500 ;
	    RECT 1458.3000 311.1000 1460.1000 311.2500 ;
	    RECT 344.7000 306.7500 346.5000 306.9000 ;
	    RECT 419.1000 306.7500 420.9000 306.9000 ;
	    RECT 344.7000 305.2500 420.9000 306.7500 ;
	    RECT 344.7000 305.1000 346.5000 305.2500 ;
	    RECT 419.1000 305.1000 420.9000 305.2500 ;
	    RECT 687.9000 306.7500 689.7000 306.9000 ;
	    RECT 971.1000 306.7500 972.9000 306.9000 ;
	    RECT 687.9000 305.2500 972.9000 306.7500 ;
	    RECT 687.9000 305.1000 689.7000 305.2500 ;
	    RECT 971.1000 305.1000 972.9000 305.2500 ;
	    RECT 999.9000 306.7500 1001.7000 306.9000 ;
	    RECT 1019.1000 306.7500 1020.9000 306.9000 ;
	    RECT 999.9000 305.2500 1020.9000 306.7500 ;
	    RECT 999.9000 305.1000 1001.7000 305.2500 ;
	    RECT 1019.1000 305.1000 1020.9000 305.2500 ;
	    RECT 1047.9000 306.7500 1049.7001 306.9000 ;
	    RECT 1131.9000 306.7500 1133.7001 306.9000 ;
	    RECT 1047.9000 305.2500 1133.7001 306.7500 ;
	    RECT 1047.9000 305.1000 1049.7001 305.2500 ;
	    RECT 1131.9000 305.1000 1133.7001 305.2500 ;
	    RECT 1170.3000 306.7500 1172.1000 306.9000 ;
	    RECT 1271.1000 306.7500 1272.9000 306.9000 ;
	    RECT 1170.3000 305.2500 1272.9000 306.7500 ;
	    RECT 1170.3000 305.1000 1172.1000 305.2500 ;
	    RECT 1271.1000 305.1000 1272.9000 305.2500 ;
	    RECT 1393.5000 306.7500 1395.3000 306.9000 ;
	    RECT 1407.9000 306.7500 1409.7001 306.9000 ;
	    RECT 1393.5000 305.2500 1409.7001 306.7500 ;
	    RECT 1393.5000 305.1000 1395.3000 305.2500 ;
	    RECT 1407.9000 305.1000 1409.7001 305.2500 ;
	    RECT 1455.9000 306.7500 1457.7001 306.9000 ;
	    RECT 1477.5000 306.7500 1479.3000 306.9000 ;
	    RECT 1455.9000 305.2500 1479.3000 306.7500 ;
	    RECT 1455.9000 305.1000 1457.7001 305.2500 ;
	    RECT 1477.5000 305.1000 1479.3000 305.2500 ;
	    RECT 416.7000 300.7500 418.5000 300.9000 ;
	    RECT 450.3000 300.7500 452.1000 300.9000 ;
	    RECT 416.7000 299.2500 452.1000 300.7500 ;
	    RECT 416.7000 299.1000 418.5000 299.2500 ;
	    RECT 450.3000 299.1000 452.1000 299.2500 ;
	    RECT 810.3000 300.7500 812.1000 300.9000 ;
	    RECT 985.5000 300.7500 987.3000 300.9000 ;
	    RECT 810.3000 299.2500 987.3000 300.7500 ;
	    RECT 810.3000 299.1000 812.1000 299.2500 ;
	    RECT 985.5000 299.1000 987.3000 299.2500 ;
	    RECT 1071.9000 300.7500 1073.7001 300.9000 ;
	    RECT 1083.9000 300.7500 1085.7001 300.9000 ;
	    RECT 1071.9000 299.2500 1085.7001 300.7500 ;
	    RECT 1071.9000 299.1000 1073.7001 299.2500 ;
	    RECT 1083.9000 299.1000 1085.7001 299.2500 ;
	    RECT 1179.9000 300.7500 1181.7001 300.9000 ;
	    RECT 1254.3000 300.7500 1256.1000 300.9000 ;
	    RECT 1179.9000 299.2500 1256.1000 300.7500 ;
	    RECT 1179.9000 299.1000 1181.7001 299.2500 ;
	    RECT 1254.3000 299.1000 1256.1000 299.2500 ;
	    RECT 1323.9000 300.7500 1325.7001 300.9000 ;
	    RECT 1388.7001 300.7500 1390.5000 300.9000 ;
	    RECT 1323.9000 299.2500 1390.5000 300.7500 ;
	    RECT 1323.9000 299.1000 1325.7001 299.2500 ;
	    RECT 1388.7001 299.1000 1390.5000 299.2500 ;
	    RECT 1455.9000 300.7500 1457.7001 300.9000 ;
	    RECT 1475.1000 300.7500 1476.9000 300.9000 ;
	    RECT 1489.5000 300.7500 1491.3000 300.9000 ;
	    RECT 1455.9000 299.2500 1491.3000 300.7500 ;
	    RECT 1455.9000 299.1000 1457.7001 299.2500 ;
	    RECT 1475.1000 299.1000 1476.9000 299.2500 ;
	    RECT 1489.5000 299.1000 1491.3000 299.2500 ;
	    RECT 147.9000 294.7500 149.7000 294.9000 ;
	    RECT 167.1000 294.7500 168.9000 294.9000 ;
	    RECT 181.5000 294.7500 183.3000 294.9000 ;
	    RECT 147.9000 293.2500 183.3000 294.7500 ;
	    RECT 147.9000 293.1000 149.7000 293.2500 ;
	    RECT 167.1000 293.1000 168.9000 293.2500 ;
	    RECT 181.5000 293.1000 183.3000 293.2500 ;
	    RECT 198.3000 294.7500 200.1000 294.9000 ;
	    RECT 205.5000 294.7500 207.3000 294.9000 ;
	    RECT 198.3000 293.2500 207.3000 294.7500 ;
	    RECT 198.3000 293.1000 200.1000 293.2500 ;
	    RECT 205.5000 293.1000 207.3000 293.2500 ;
	    RECT 325.5000 294.7500 327.3000 294.9000 ;
	    RECT 359.1000 294.7500 360.9000 294.9000 ;
	    RECT 325.5000 293.2500 360.9000 294.7500 ;
	    RECT 325.5000 293.1000 327.3000 293.2500 ;
	    RECT 359.1000 293.1000 360.9000 293.2500 ;
	    RECT 1033.5000 294.7500 1035.3000 294.9000 ;
	    RECT 1047.9000 294.7500 1049.7001 294.9000 ;
	    RECT 1033.5000 293.2500 1049.7001 294.7500 ;
	    RECT 1033.5000 293.1000 1035.3000 293.2500 ;
	    RECT 1047.9000 293.1000 1049.7001 293.2500 ;
	    RECT 1083.9000 294.7500 1085.7001 294.9000 ;
	    RECT 1107.9000 294.7500 1109.7001 294.9000 ;
	    RECT 1083.9000 293.2500 1109.7001 294.7500 ;
	    RECT 1083.9000 293.1000 1085.7001 293.2500 ;
	    RECT 1107.9000 293.1000 1109.7001 293.2500 ;
	    RECT 1220.7001 294.7500 1222.5000 294.9000 ;
	    RECT 1292.7001 294.7500 1294.5000 294.9000 ;
	    RECT 1323.9000 294.7500 1325.7001 294.9000 ;
	    RECT 1220.7001 293.2500 1325.7001 294.7500 ;
	    RECT 1220.7001 293.1000 1222.5000 293.2500 ;
	    RECT 1292.7001 293.1000 1294.5000 293.2500 ;
	    RECT 1323.9000 293.1000 1325.7001 293.2500 ;
	    RECT 1441.5000 294.7500 1443.3000 294.9000 ;
	    RECT 1463.1000 294.7500 1464.9000 294.9000 ;
	    RECT 1479.9000 294.7500 1481.7001 294.9000 ;
	    RECT 1441.5000 293.2500 1481.7001 294.7500 ;
	    RECT 1441.5000 293.1000 1443.3000 293.2500 ;
	    RECT 1463.1000 293.1000 1464.9000 293.2500 ;
	    RECT 1479.9000 293.1000 1481.7001 293.2500 ;
	    RECT 1511.1000 294.7500 1512.9000 294.9000 ;
	    RECT 1563.9000 294.7500 1565.7001 294.9000 ;
	    RECT 1511.1000 293.2500 1565.7001 294.7500 ;
	    RECT 1511.1000 293.1000 1512.9000 293.2500 ;
	    RECT 1563.9000 293.1000 1565.7001 293.2500 ;
	    RECT 25.5000 288.7500 27.3000 288.9000 ;
	    RECT 75.9000 288.7500 77.7000 288.9000 ;
	    RECT 25.5000 287.2500 77.7000 288.7500 ;
	    RECT 25.5000 287.1000 27.3000 287.2500 ;
	    RECT 75.9000 287.1000 77.7000 287.2500 ;
	    RECT 167.1000 288.7500 168.9000 288.9000 ;
	    RECT 176.7000 288.7500 178.5000 288.9000 ;
	    RECT 167.1000 287.2500 178.5000 288.7500 ;
	    RECT 167.1000 287.1000 168.9000 287.2500 ;
	    RECT 176.7000 287.1000 178.5000 287.2500 ;
	    RECT 721.5000 288.7500 723.3000 288.9000 ;
	    RECT 747.9000 288.7500 749.7000 288.9000 ;
	    RECT 721.5000 287.2500 749.7000 288.7500 ;
	    RECT 721.5000 287.1000 723.3000 287.2500 ;
	    RECT 747.9000 287.1000 749.7000 287.2500 ;
	    RECT 968.7000 288.7500 970.5000 288.9000 ;
	    RECT 1088.7001 288.7500 1090.5000 288.9000 ;
	    RECT 968.7000 287.2500 1090.5000 288.7500 ;
	    RECT 968.7000 287.1000 970.5000 287.2500 ;
	    RECT 1088.7001 287.1000 1090.5000 287.2500 ;
	    RECT 1093.5000 288.7500 1095.3000 288.9000 ;
	    RECT 1131.9000 288.7500 1133.7001 288.9000 ;
	    RECT 1093.5000 287.2500 1133.7001 288.7500 ;
	    RECT 1093.5000 287.1000 1095.3000 287.2500 ;
	    RECT 1131.9000 287.1000 1133.7001 287.2500 ;
	    RECT 1155.9000 288.7500 1157.7001 288.9000 ;
	    RECT 1175.1000 288.7500 1176.9000 288.9000 ;
	    RECT 1155.9000 287.2500 1176.9000 288.7500 ;
	    RECT 1155.9000 287.1000 1157.7001 287.2500 ;
	    RECT 1175.1000 287.1000 1176.9000 287.2500 ;
	    RECT 1184.7001 288.7500 1186.5000 288.9000 ;
	    RECT 1206.3000 288.7500 1208.1000 288.9000 ;
	    RECT 1184.7001 287.2500 1208.1000 288.7500 ;
	    RECT 1184.7001 287.1000 1186.5000 287.2500 ;
	    RECT 1206.3000 287.1000 1208.1000 287.2500 ;
	    RECT 1323.9000 288.7500 1325.7001 288.9000 ;
	    RECT 1343.1000 288.7500 1344.9000 288.9000 ;
	    RECT 1323.9000 287.2500 1344.9000 288.7500 ;
	    RECT 1323.9000 287.1000 1325.7001 287.2500 ;
	    RECT 1343.1000 287.1000 1344.9000 287.2500 ;
	    RECT 1371.9000 288.7500 1373.7001 288.9000 ;
	    RECT 1405.5000 288.7500 1407.3000 288.9000 ;
	    RECT 1371.9000 287.2500 1407.3000 288.7500 ;
	    RECT 1371.9000 287.1000 1373.7001 287.2500 ;
	    RECT 1405.5000 287.1000 1407.3000 287.2500 ;
	    RECT 1429.5000 288.7500 1431.3000 288.9000 ;
	    RECT 1451.1000 288.7500 1452.9000 288.9000 ;
	    RECT 1429.5000 287.2500 1452.9000 288.7500 ;
	    RECT 1429.5000 287.1000 1431.3000 287.2500 ;
	    RECT 1451.1000 287.1000 1452.9000 287.2500 ;
	    RECT 1539.9000 288.7500 1541.7001 288.9000 ;
	    RECT 1551.9000 288.7500 1553.7001 288.9000 ;
	    RECT 1539.9000 287.2500 1553.7001 288.7500 ;
	    RECT 1539.9000 287.1000 1541.7001 287.2500 ;
	    RECT 1551.9000 287.1000 1553.7001 287.2500 ;
	    RECT 159.9000 282.7500 161.7000 282.9000 ;
	    RECT 176.7000 282.7500 178.5000 282.9000 ;
	    RECT 159.9000 281.2500 178.5000 282.7500 ;
	    RECT 159.9000 281.1000 161.7000 281.2500 ;
	    RECT 176.7000 281.1000 178.5000 281.2500 ;
	    RECT 567.9000 282.7500 569.7000 282.9000 ;
	    RECT 606.3000 282.7500 608.1000 282.9000 ;
	    RECT 567.9000 281.2500 608.1000 282.7500 ;
	    RECT 567.9000 281.1000 569.7000 281.2500 ;
	    RECT 606.3000 281.1000 608.1000 281.2500 ;
	    RECT 733.5000 282.7500 735.3000 282.9000 ;
	    RECT 783.9000 282.7500 785.7000 282.9000 ;
	    RECT 843.9000 282.7500 845.7000 282.9000 ;
	    RECT 733.5000 281.2500 845.7000 282.7500 ;
	    RECT 733.5000 281.1000 735.3000 281.2500 ;
	    RECT 783.9000 281.1000 785.7000 281.2500 ;
	    RECT 843.9000 281.1000 845.7000 281.2500 ;
	    RECT 872.7000 282.7500 874.5000 282.9000 ;
	    RECT 879.9000 282.7500 881.7000 282.9000 ;
	    RECT 872.7000 281.2500 881.7000 282.7500 ;
	    RECT 872.7000 281.1000 874.5000 281.2500 ;
	    RECT 879.9000 281.1000 881.7000 281.2500 ;
	    RECT 1014.3000 282.7500 1016.1000 282.9000 ;
	    RECT 1043.1000 282.7500 1044.9000 282.9000 ;
	    RECT 1014.3000 281.2500 1044.9000 282.7500 ;
	    RECT 1014.3000 281.1000 1016.1000 281.2500 ;
	    RECT 1043.1000 281.1000 1044.9000 281.2500 ;
	    RECT 1069.5000 282.7500 1071.3000 282.9000 ;
	    RECT 1110.3000 282.7500 1112.1000 282.9000 ;
	    RECT 1069.5000 281.2500 1112.1000 282.7500 ;
	    RECT 1069.5000 281.1000 1071.3000 281.2500 ;
	    RECT 1110.3000 281.1000 1112.1000 281.2500 ;
	    RECT 1148.7001 282.7500 1150.5000 282.9000 ;
	    RECT 1187.1000 282.7500 1188.9000 282.9000 ;
	    RECT 1148.7001 281.2500 1188.9000 282.7500 ;
	    RECT 1148.7001 281.1000 1150.5000 281.2500 ;
	    RECT 1187.1000 281.1000 1188.9000 281.2500 ;
	    RECT 1203.9000 282.7500 1205.7001 282.9000 ;
	    RECT 1328.7001 282.7500 1330.5000 282.9000 ;
	    RECT 1367.1000 282.7500 1368.9000 282.9000 ;
	    RECT 1403.1000 282.7500 1404.9000 282.9000 ;
	    RECT 1203.9000 281.2500 1404.9000 282.7500 ;
	    RECT 1203.9000 281.1000 1205.7001 281.2500 ;
	    RECT 1328.7001 281.1000 1330.5000 281.2500 ;
	    RECT 1367.1000 281.1000 1368.9000 281.2500 ;
	    RECT 1403.1000 281.1000 1404.9000 281.2500 ;
	    RECT 1419.9000 282.7500 1421.7001 282.9000 ;
	    RECT 1429.5000 282.7500 1431.3000 282.9000 ;
	    RECT 1419.9000 281.2500 1431.3000 282.7500 ;
	    RECT 1419.9000 281.1000 1421.7001 281.2500 ;
	    RECT 1429.5000 281.1000 1431.3000 281.2500 ;
	    RECT 1477.5000 282.7500 1479.3000 282.9000 ;
	    RECT 1487.1000 282.7500 1488.9000 282.9000 ;
	    RECT 1477.5000 281.2500 1488.9000 282.7500 ;
	    RECT 1477.5000 281.1000 1479.3000 281.2500 ;
	    RECT 1487.1000 281.1000 1488.9000 281.2500 ;
	    RECT 1513.5000 282.7500 1515.3000 282.9000 ;
	    RECT 1518.3000 282.7500 1520.1000 282.9000 ;
	    RECT 1513.5000 281.2500 1520.1000 282.7500 ;
	    RECT 1513.5000 281.1000 1515.3000 281.2500 ;
	    RECT 1518.3000 281.1000 1520.1000 281.2500 ;
	    RECT 1539.9000 282.7500 1541.7001 282.9000 ;
	    RECT 1559.1000 282.7500 1560.9000 282.9000 ;
	    RECT 1539.9000 281.2500 1560.9000 282.7500 ;
	    RECT 1539.9000 281.1000 1541.7001 281.2500 ;
	    RECT 1559.1000 281.1000 1560.9000 281.2500 ;
	    RECT 140.7000 276.7500 142.5000 276.9000 ;
	    RECT 176.7000 276.7500 178.5000 276.9000 ;
	    RECT 140.7000 275.2500 178.5000 276.7500 ;
	    RECT 140.7000 275.1000 142.5000 275.2500 ;
	    RECT 176.7000 275.1000 178.5000 275.2500 ;
	    RECT 570.3000 276.7500 572.1000 276.9000 ;
	    RECT 615.9000 276.7500 617.7000 276.9000 ;
	    RECT 570.3000 275.2500 617.7000 276.7500 ;
	    RECT 570.3000 275.1000 572.1000 275.2500 ;
	    RECT 615.9000 275.1000 617.7000 275.2500 ;
	    RECT 1134.3000 276.7500 1136.1000 276.9000 ;
	    RECT 1158.3000 276.7500 1160.1000 276.9000 ;
	    RECT 1134.3000 275.2500 1160.1000 276.7500 ;
	    RECT 1134.3000 275.1000 1136.1000 275.2500 ;
	    RECT 1158.3000 275.1000 1160.1000 275.2500 ;
	    RECT 1179.9000 276.7500 1181.7001 276.9000 ;
	    RECT 1211.1000 276.7500 1212.9000 276.9000 ;
	    RECT 1179.9000 275.2500 1212.9000 276.7500 ;
	    RECT 1179.9000 275.1000 1181.7001 275.2500 ;
	    RECT 1211.1000 275.1000 1212.9000 275.2500 ;
	    RECT 1271.1000 276.7500 1272.9000 276.9000 ;
	    RECT 1275.9000 276.7500 1277.7001 276.9000 ;
	    RECT 1271.1000 275.2500 1277.7001 276.7500 ;
	    RECT 1271.1000 275.1000 1272.9000 275.2500 ;
	    RECT 1275.9000 275.1000 1277.7001 275.2500 ;
	    RECT 1309.5000 276.7500 1311.3000 276.9000 ;
	    RECT 1369.5000 276.7500 1371.3000 276.9000 ;
	    RECT 1309.5000 275.2500 1371.3000 276.7500 ;
	    RECT 1309.5000 275.1000 1311.3000 275.2500 ;
	    RECT 1369.5000 275.1000 1371.3000 275.2500 ;
	    RECT 1439.1000 276.7500 1440.9000 276.9000 ;
	    RECT 1523.1000 276.7500 1524.9000 276.9000 ;
	    RECT 1439.1000 275.2500 1524.9000 276.7500 ;
	    RECT 1439.1000 275.1000 1440.9000 275.2500 ;
	    RECT 1523.1000 275.1000 1524.9000 275.2500 ;
	    RECT 176.7000 270.7500 178.5000 270.9000 ;
	    RECT 195.9000 270.7500 197.7000 270.9000 ;
	    RECT 176.7000 269.2500 197.7000 270.7500 ;
	    RECT 176.7000 269.1000 178.5000 269.2500 ;
	    RECT 195.9000 269.1000 197.7000 269.2500 ;
	    RECT 534.3000 270.7500 536.1000 270.9000 ;
	    RECT 558.3000 270.7500 560.1000 270.9000 ;
	    RECT 534.3000 269.2500 560.1000 270.7500 ;
	    RECT 534.3000 269.1000 536.1000 269.2500 ;
	    RECT 558.3000 269.1000 560.1000 269.2500 ;
	    RECT 1011.9000 270.7500 1013.7000 270.9000 ;
	    RECT 1021.5000 270.7500 1023.3000 270.9000 ;
	    RECT 1011.9000 269.2500 1023.3000 270.7500 ;
	    RECT 1011.9000 269.1000 1013.7000 269.2500 ;
	    RECT 1021.5000 269.1000 1023.3000 269.2500 ;
	    RECT 1095.9000 270.7500 1097.7001 270.9000 ;
	    RECT 1115.1000 270.7500 1116.9000 270.9000 ;
	    RECT 1179.9000 270.7500 1181.7001 270.9000 ;
	    RECT 1095.9000 269.2500 1181.7001 270.7500 ;
	    RECT 1095.9000 269.1000 1097.7001 269.2500 ;
	    RECT 1115.1000 269.1000 1116.9000 269.2500 ;
	    RECT 1179.9000 269.1000 1181.7001 269.2500 ;
	    RECT 1187.1000 270.7500 1188.9000 270.9000 ;
	    RECT 1206.3000 270.7500 1208.1000 270.9000 ;
	    RECT 1187.1000 269.2500 1208.1000 270.7500 ;
	    RECT 1187.1000 269.1000 1188.9000 269.2500 ;
	    RECT 1206.3000 269.1000 1208.1000 269.2500 ;
	    RECT 1213.5000 270.7500 1215.3000 270.9000 ;
	    RECT 1321.5000 270.7500 1323.3000 270.9000 ;
	    RECT 1213.5000 269.2500 1323.3000 270.7500 ;
	    RECT 1213.5000 269.1000 1215.3000 269.2500 ;
	    RECT 1321.5000 269.1000 1323.3000 269.2500 ;
	    RECT 1446.3000 270.7500 1448.1000 270.9000 ;
	    RECT 1470.3000 270.7500 1472.1000 270.9000 ;
	    RECT 1446.3000 269.2500 1472.1000 270.7500 ;
	    RECT 1446.3000 269.1000 1448.1000 269.2500 ;
	    RECT 1470.3000 269.1000 1472.1000 269.2500 ;
	    RECT 1506.3000 270.7500 1508.1000 270.9000 ;
	    RECT 1525.5000 270.7500 1527.3000 270.9000 ;
	    RECT 1506.3000 269.2500 1527.3000 270.7500 ;
	    RECT 1506.3000 269.1000 1508.1000 269.2500 ;
	    RECT 1525.5000 269.1000 1527.3000 269.2500 ;
	    RECT 1539.9000 270.7500 1541.7001 270.9000 ;
	    RECT 1554.3000 270.7500 1556.1000 270.9000 ;
	    RECT 1539.9000 269.2500 1556.1000 270.7500 ;
	    RECT 1539.9000 269.1000 1541.7001 269.2500 ;
	    RECT 1554.3000 269.1000 1556.1000 269.2500 ;
	    RECT 301.5000 264.7500 303.3000 264.9000 ;
	    RECT 339.9000 264.7500 341.7000 264.9000 ;
	    RECT 301.5000 263.2500 341.7000 264.7500 ;
	    RECT 301.5000 263.1000 303.3000 263.2500 ;
	    RECT 339.9000 263.1000 341.7000 263.2500 ;
	    RECT 395.1000 264.7500 396.9000 264.9000 ;
	    RECT 510.3000 264.7500 512.1000 264.9000 ;
	    RECT 395.1000 263.2500 512.1000 264.7500 ;
	    RECT 395.1000 263.1000 396.9000 263.2500 ;
	    RECT 510.3000 263.1000 512.1000 263.2500 ;
	    RECT 529.5000 264.7500 531.3000 264.9000 ;
	    RECT 558.3000 264.7500 560.1000 264.9000 ;
	    RECT 529.5000 263.2500 560.1000 264.7500 ;
	    RECT 529.5000 263.1000 531.3000 263.2500 ;
	    RECT 558.3000 263.1000 560.1000 263.2500 ;
	    RECT 709.5000 264.7500 711.3000 264.9000 ;
	    RECT 788.7000 264.7500 790.5000 264.9000 ;
	    RECT 815.1000 264.7500 816.9000 264.9000 ;
	    RECT 709.5000 263.2500 816.9000 264.7500 ;
	    RECT 709.5000 263.1000 711.3000 263.2500 ;
	    RECT 788.7000 263.1000 790.5000 263.2500 ;
	    RECT 815.1000 263.1000 816.9000 263.2500 ;
	    RECT 877.5000 264.7500 879.3000 264.9000 ;
	    RECT 1021.5000 264.7500 1023.3000 264.9000 ;
	    RECT 877.5000 263.2500 1023.3000 264.7500 ;
	    RECT 877.5000 263.1000 879.3000 263.2500 ;
	    RECT 1021.5000 263.1000 1023.3000 263.2500 ;
	    RECT 1040.7001 264.7500 1042.5000 264.9000 ;
	    RECT 1071.9000 264.7500 1073.7001 264.9000 ;
	    RECT 1079.1000 264.7500 1080.9000 264.9000 ;
	    RECT 1040.7001 263.2500 1080.9000 264.7500 ;
	    RECT 1040.7001 263.1000 1042.5000 263.2500 ;
	    RECT 1071.9000 263.1000 1073.7001 263.2500 ;
	    RECT 1079.1000 263.1000 1080.9000 263.2500 ;
	    RECT 1100.7001 264.7500 1102.5000 264.9000 ;
	    RECT 1105.5000 264.7500 1107.3000 264.9000 ;
	    RECT 1119.9000 264.7500 1121.7001 264.9000 ;
	    RECT 1100.7001 263.2500 1121.7001 264.7500 ;
	    RECT 1100.7001 263.1000 1102.5000 263.2500 ;
	    RECT 1105.5000 263.1000 1107.3000 263.2500 ;
	    RECT 1119.9000 263.1000 1121.7001 263.2500 ;
	    RECT 1203.9000 264.7500 1205.7001 264.9000 ;
	    RECT 1220.7001 264.7500 1222.5000 264.9000 ;
	    RECT 1247.1000 264.7500 1248.9000 264.9000 ;
	    RECT 1292.7001 264.7500 1294.5000 264.9000 ;
	    RECT 1203.9000 263.2500 1294.5000 264.7500 ;
	    RECT 1203.9000 263.1000 1205.7001 263.2500 ;
	    RECT 1220.7001 263.1000 1222.5000 263.2500 ;
	    RECT 1247.1000 263.1000 1248.9000 263.2500 ;
	    RECT 1292.7001 263.1000 1294.5000 263.2500 ;
	    RECT 1333.5000 264.7500 1335.3000 264.9000 ;
	    RECT 1398.3000 264.7500 1400.1000 264.9000 ;
	    RECT 1441.5000 264.7500 1443.3000 264.9000 ;
	    RECT 1333.5000 263.2500 1443.3000 264.7500 ;
	    RECT 1333.5000 263.1000 1335.3000 263.2500 ;
	    RECT 1398.3000 263.1000 1400.1000 263.2500 ;
	    RECT 1441.5000 263.1000 1443.3000 263.2500 ;
	    RECT 1520.7001 264.7500 1522.5000 264.9000 ;
	    RECT 1556.7001 264.7500 1558.5000 264.9000 ;
	    RECT 1520.7001 263.2500 1558.5000 264.7500 ;
	    RECT 1520.7001 263.1000 1522.5000 263.2500 ;
	    RECT 1556.7001 263.1000 1558.5000 263.2500 ;
	    RECT 368.7000 258.7500 370.5000 258.9000 ;
	    RECT 375.9000 258.7500 377.7000 258.9000 ;
	    RECT 368.7000 257.2500 377.7000 258.7500 ;
	    RECT 368.7000 257.1000 370.5000 257.2500 ;
	    RECT 375.9000 257.1000 377.7000 257.2500 ;
	    RECT 575.1000 258.7500 576.9000 258.9000 ;
	    RECT 587.1000 258.7500 588.9000 258.9000 ;
	    RECT 575.1000 257.2500 588.9000 258.7500 ;
	    RECT 575.1000 257.1000 576.9000 257.2500 ;
	    RECT 587.1000 257.1000 588.9000 257.2500 ;
	    RECT 618.3000 258.7500 620.1000 258.9000 ;
	    RECT 723.9000 258.7500 725.7000 258.9000 ;
	    RECT 618.3000 257.2500 725.7000 258.7500 ;
	    RECT 618.3000 257.1000 620.1000 257.2500 ;
	    RECT 723.9000 257.1000 725.7000 257.2500 ;
	    RECT 781.5000 258.7500 783.3000 258.9000 ;
	    RECT 819.9000 258.7500 821.7000 258.9000 ;
	    RECT 781.5000 257.2500 821.7000 258.7500 ;
	    RECT 781.5000 257.1000 783.3000 257.2500 ;
	    RECT 819.9000 257.1000 821.7000 257.2500 ;
	    RECT 1177.5000 258.7500 1179.3000 258.9000 ;
	    RECT 1208.7001 258.7500 1210.5000 258.9000 ;
	    RECT 1177.5000 257.2500 1210.5000 258.7500 ;
	    RECT 1177.5000 257.1000 1179.3000 257.2500 ;
	    RECT 1208.7001 257.1000 1210.5000 257.2500 ;
	    RECT 1218.3000 258.7500 1220.1000 258.9000 ;
	    RECT 1268.7001 258.7500 1270.5000 258.9000 ;
	    RECT 1299.9000 258.7500 1301.7001 258.9000 ;
	    RECT 1218.3000 257.2500 1301.7001 258.7500 ;
	    RECT 1218.3000 257.1000 1220.1000 257.2500 ;
	    RECT 1268.7001 257.1000 1270.5000 257.2500 ;
	    RECT 1299.9000 257.1000 1301.7001 257.2500 ;
	    RECT 1321.5000 258.7500 1323.3000 258.9000 ;
	    RECT 1331.1000 258.7500 1332.9000 258.9000 ;
	    RECT 1321.5000 257.2500 1332.9000 258.7500 ;
	    RECT 1321.5000 257.1000 1323.3000 257.2500 ;
	    RECT 1331.1000 257.1000 1332.9000 257.2500 ;
	    RECT 1359.9000 258.7500 1361.7001 258.9000 ;
	    RECT 1371.9000 258.7500 1373.7001 258.9000 ;
	    RECT 1359.9000 257.2500 1373.7001 258.7500 ;
	    RECT 1359.9000 257.1000 1361.7001 257.2500 ;
	    RECT 1371.9000 257.1000 1373.7001 257.2500 ;
	    RECT 1508.7001 258.7500 1510.5000 258.9000 ;
	    RECT 1549.5000 258.7500 1551.3000 258.9000 ;
	    RECT 1508.7001 257.2500 1551.3000 258.7500 ;
	    RECT 1508.7001 257.1000 1510.5000 257.2500 ;
	    RECT 1549.5000 257.1000 1551.3000 257.2500 ;
	    RECT 1554.3000 258.7500 1556.1000 258.9000 ;
	    RECT 1566.3000 258.7500 1568.1000 258.9000 ;
	    RECT 1554.3000 257.2500 1568.1000 258.7500 ;
	    RECT 1554.3000 257.1000 1556.1000 257.2500 ;
	    RECT 1566.3000 257.1000 1568.1000 257.2500 ;
	    RECT 162.3000 252.7500 164.1000 252.9000 ;
	    RECT 171.9000 252.7500 173.7000 252.9000 ;
	    RECT 162.3000 251.2500 173.7000 252.7500 ;
	    RECT 162.3000 251.1000 164.1000 251.2500 ;
	    RECT 171.9000 251.1000 173.7000 251.2500 ;
	    RECT 181.5000 252.7500 183.3000 252.9000 ;
	    RECT 313.5000 252.7500 315.3000 252.9000 ;
	    RECT 181.5000 251.2500 315.3000 252.7500 ;
	    RECT 181.5000 251.1000 183.3000 251.2500 ;
	    RECT 313.5000 251.1000 315.3000 251.2500 ;
	    RECT 366.3000 252.7500 368.1000 252.9000 ;
	    RECT 373.5000 252.7500 375.3000 252.9000 ;
	    RECT 366.3000 251.2500 375.3000 252.7500 ;
	    RECT 366.3000 251.1000 368.1000 251.2500 ;
	    RECT 373.5000 251.1000 375.3000 251.2500 ;
	    RECT 836.7000 252.7500 838.5000 252.9000 ;
	    RECT 1093.5000 252.7500 1095.3000 252.9000 ;
	    RECT 836.7000 251.2500 1095.3000 252.7500 ;
	    RECT 836.7000 251.1000 838.5000 251.2500 ;
	    RECT 1093.5000 251.1000 1095.3000 251.2500 ;
	    RECT 1098.3000 252.7500 1100.1000 252.9000 ;
	    RECT 1218.3000 252.7500 1220.1000 252.9000 ;
	    RECT 1098.3000 251.2500 1220.1000 252.7500 ;
	    RECT 1098.3000 251.1000 1100.1000 251.2500 ;
	    RECT 1218.3000 251.1000 1220.1000 251.2500 ;
	    RECT 1261.5000 252.7500 1263.3000 252.9000 ;
	    RECT 1328.7001 252.7500 1330.5000 252.9000 ;
	    RECT 1261.5000 251.2500 1330.5000 252.7500 ;
	    RECT 1261.5000 251.1000 1263.3000 251.2500 ;
	    RECT 1328.7001 251.1000 1330.5000 251.2500 ;
	    RECT 1405.5000 252.7500 1407.3000 252.9000 ;
	    RECT 1436.7001 252.7500 1438.5000 252.9000 ;
	    RECT 1405.5000 251.2500 1438.5000 252.7500 ;
	    RECT 1405.5000 251.1000 1407.3000 251.2500 ;
	    RECT 1436.7001 251.1000 1438.5000 251.2500 ;
	    RECT 1489.5000 252.7500 1491.3000 252.9000 ;
	    RECT 1520.7001 252.7500 1522.5000 252.9000 ;
	    RECT 1489.5000 251.2500 1522.5000 252.7500 ;
	    RECT 1489.5000 251.1000 1491.3000 251.2500 ;
	    RECT 1520.7001 251.1000 1522.5000 251.2500 ;
	    RECT 1549.5000 252.7500 1551.3000 252.9000 ;
	    RECT 1556.7001 252.7500 1558.5000 252.9000 ;
	    RECT 1549.5000 251.2500 1558.5000 252.7500 ;
	    RECT 1549.5000 251.1000 1551.3000 251.2500 ;
	    RECT 1556.7001 251.1000 1558.5000 251.2500 ;
	    RECT 133.5000 246.7500 135.3000 246.9000 ;
	    RECT 253.5000 246.7500 255.3000 246.9000 ;
	    RECT 133.5000 245.2500 255.3000 246.7500 ;
	    RECT 133.5000 245.1000 135.3000 245.2500 ;
	    RECT 253.5000 245.1000 255.3000 245.2500 ;
	    RECT 308.7000 246.7500 310.5000 246.9000 ;
	    RECT 320.7000 246.7500 322.5000 246.9000 ;
	    RECT 349.5000 246.7500 351.3000 246.9000 ;
	    RECT 443.1000 246.7500 444.9000 246.9000 ;
	    RECT 308.7000 245.2500 444.9000 246.7500 ;
	    RECT 308.7000 245.1000 310.5000 245.2500 ;
	    RECT 320.7000 245.1000 322.5000 245.2500 ;
	    RECT 349.5000 245.1000 351.3000 245.2500 ;
	    RECT 443.1000 245.1000 444.9000 245.2500 ;
	    RECT 539.1000 246.7500 540.9000 246.9000 ;
	    RECT 543.9000 246.7500 545.7000 246.9000 ;
	    RECT 539.1000 245.2500 545.7000 246.7500 ;
	    RECT 539.1000 245.1000 540.9000 245.2500 ;
	    RECT 543.9000 245.1000 545.7000 245.2500 ;
	    RECT 575.1000 246.7500 576.9000 246.9000 ;
	    RECT 747.9000 246.7500 749.7000 246.9000 ;
	    RECT 575.1000 245.2500 749.7000 246.7500 ;
	    RECT 575.1000 245.1000 576.9000 245.2500 ;
	    RECT 747.9000 245.1000 749.7000 245.2500 ;
	    RECT 1079.1000 246.7500 1080.9000 246.9000 ;
	    RECT 1196.7001 246.7500 1198.5000 246.9000 ;
	    RECT 1079.1000 245.2500 1198.5000 246.7500 ;
	    RECT 1079.1000 245.1000 1080.9000 245.2500 ;
	    RECT 1196.7001 245.1000 1198.5000 245.2500 ;
	    RECT 1206.3000 246.7500 1208.1000 246.9000 ;
	    RECT 1261.5000 246.7500 1263.3000 246.9000 ;
	    RECT 1206.3000 245.2500 1263.3000 246.7500 ;
	    RECT 1206.3000 245.1000 1208.1000 245.2500 ;
	    RECT 1261.5000 245.1000 1263.3000 245.2500 ;
	    RECT 1278.3000 246.7500 1280.1000 246.9000 ;
	    RECT 1323.9000 246.7500 1325.7001 246.9000 ;
	    RECT 1278.3000 245.2500 1325.7001 246.7500 ;
	    RECT 1278.3000 245.1000 1280.1000 245.2500 ;
	    RECT 1323.9000 245.1000 1325.7001 245.2500 ;
	    RECT 1417.5000 246.7500 1419.3000 246.9000 ;
	    RECT 1482.3000 246.7500 1484.1000 246.9000 ;
	    RECT 1417.5000 245.2500 1484.1000 246.7500 ;
	    RECT 1417.5000 245.1000 1419.3000 245.2500 ;
	    RECT 1482.3000 245.1000 1484.1000 245.2500 ;
	    RECT 164.7000 240.7500 166.5000 240.9000 ;
	    RECT 169.5000 240.7500 171.3000 240.9000 ;
	    RECT 164.7000 239.2500 171.3000 240.7500 ;
	    RECT 164.7000 239.1000 166.5000 239.2500 ;
	    RECT 169.5000 239.1000 171.3000 239.2500 ;
	    RECT 606.3000 240.7500 608.1000 240.9000 ;
	    RECT 627.9000 240.7500 629.7000 240.9000 ;
	    RECT 606.3000 239.2500 629.7000 240.7500 ;
	    RECT 606.3000 239.1000 608.1000 239.2500 ;
	    RECT 627.9000 239.1000 629.7000 239.2500 ;
	    RECT 1134.3000 240.7500 1136.1000 240.9000 ;
	    RECT 1170.3000 240.7500 1172.1000 240.9000 ;
	    RECT 1134.3000 239.2500 1172.1000 240.7500 ;
	    RECT 1134.3000 239.1000 1136.1000 239.2500 ;
	    RECT 1170.3000 239.1000 1172.1000 239.2500 ;
	    RECT 1208.7001 240.7500 1210.5000 240.9000 ;
	    RECT 1242.3000 240.7500 1244.1000 240.9000 ;
	    RECT 1208.7001 239.2500 1244.1000 240.7500 ;
	    RECT 1208.7001 239.1000 1210.5000 239.2500 ;
	    RECT 1242.3000 239.1000 1244.1000 239.2500 ;
	    RECT 1256.7001 240.7500 1258.5000 240.9000 ;
	    RECT 1340.7001 240.7500 1342.5000 240.9000 ;
	    RECT 1379.1000 240.7500 1380.9000 240.9000 ;
	    RECT 1256.7001 239.2500 1380.9000 240.7500 ;
	    RECT 1256.7001 239.1000 1258.5000 239.2500 ;
	    RECT 1340.7001 239.1000 1342.5000 239.2500 ;
	    RECT 1379.1000 239.1000 1380.9000 239.2500 ;
	    RECT 1407.9000 240.7500 1409.7001 240.9000 ;
	    RECT 1412.7001 240.7500 1414.5000 240.9000 ;
	    RECT 1407.9000 239.2500 1414.5000 240.7500 ;
	    RECT 1407.9000 239.1000 1409.7001 239.2500 ;
	    RECT 1412.7001 239.1000 1414.5000 239.2500 ;
	    RECT 1470.3000 240.7500 1472.1000 240.9000 ;
	    RECT 1511.1000 240.7500 1512.9000 240.9000 ;
	    RECT 1470.3000 239.2500 1512.9000 240.7500 ;
	    RECT 1470.3000 239.1000 1472.1000 239.2500 ;
	    RECT 1511.1000 239.1000 1512.9000 239.2500 ;
	    RECT 1523.1000 240.7500 1524.9000 240.9000 ;
	    RECT 1542.3000 240.7500 1544.1000 240.9000 ;
	    RECT 1523.1000 239.2500 1544.1000 240.7500 ;
	    RECT 1523.1000 239.1000 1524.9000 239.2500 ;
	    RECT 1542.3000 239.1000 1544.1000 239.2500 ;
	    RECT 231.9000 234.7500 233.7000 234.9000 ;
	    RECT 306.3000 234.7500 308.1000 234.9000 ;
	    RECT 231.9000 233.2500 308.1000 234.7500 ;
	    RECT 231.9000 233.1000 233.7000 233.2500 ;
	    RECT 306.3000 233.1000 308.1000 233.2500 ;
	    RECT 596.7000 234.7500 598.5000 234.9000 ;
	    RECT 925.5000 234.7500 927.3000 234.9000 ;
	    RECT 596.7000 233.2500 927.3000 234.7500 ;
	    RECT 596.7000 233.1000 598.5000 233.2500 ;
	    RECT 925.5000 233.1000 927.3000 233.2500 ;
	    RECT 1004.7000 234.7500 1006.5000 234.9000 ;
	    RECT 1052.7001 234.7500 1054.5000 234.9000 ;
	    RECT 1004.7000 233.2500 1054.5000 234.7500 ;
	    RECT 1004.7000 233.1000 1006.5000 233.2500 ;
	    RECT 1052.7001 233.1000 1054.5000 233.2500 ;
	    RECT 1093.5000 234.7500 1095.3000 234.9000 ;
	    RECT 1134.3000 234.7500 1136.1000 234.9000 ;
	    RECT 1093.5000 233.2500 1136.1000 234.7500 ;
	    RECT 1093.5000 233.1000 1095.3000 233.2500 ;
	    RECT 1134.3000 233.1000 1136.1000 233.2500 ;
	    RECT 1191.9000 234.7500 1193.7001 234.9000 ;
	    RECT 1201.5000 234.7500 1203.3000 234.9000 ;
	    RECT 1191.9000 233.2500 1203.3000 234.7500 ;
	    RECT 1191.9000 233.1000 1193.7001 233.2500 ;
	    RECT 1201.5000 233.1000 1203.3000 233.2500 ;
	    RECT 1259.1000 234.7500 1260.9000 234.9000 ;
	    RECT 1278.3000 234.7500 1280.1000 234.9000 ;
	    RECT 1259.1000 233.2500 1280.1000 234.7500 ;
	    RECT 1259.1000 233.1000 1260.9000 233.2500 ;
	    RECT 1278.3000 233.1000 1280.1000 233.2500 ;
	    RECT 1290.3000 234.7500 1292.1000 234.9000 ;
	    RECT 1295.1000 234.7500 1296.9000 234.9000 ;
	    RECT 1290.3000 233.2500 1296.9000 234.7500 ;
	    RECT 1290.3000 233.1000 1292.1000 233.2500 ;
	    RECT 1295.1000 233.1000 1296.9000 233.2500 ;
	    RECT 1304.7001 234.7500 1306.5000 234.9000 ;
	    RECT 1434.3000 234.7500 1436.1000 234.9000 ;
	    RECT 1460.7001 234.7500 1462.5000 234.9000 ;
	    RECT 1304.7001 233.2500 1462.5000 234.7500 ;
	    RECT 1304.7001 233.1000 1306.5000 233.2500 ;
	    RECT 1434.3000 233.1000 1436.1000 233.2500 ;
	    RECT 1460.7001 233.1000 1462.5000 233.2500 ;
	    RECT 1487.1000 234.7500 1488.9000 234.9000 ;
	    RECT 1508.7001 234.7500 1510.5000 234.9000 ;
	    RECT 1487.1000 233.2500 1510.5000 234.7500 ;
	    RECT 1487.1000 233.1000 1488.9000 233.2500 ;
	    RECT 1508.7001 233.1000 1510.5000 233.2500 ;
	    RECT 1513.5000 234.7500 1515.3000 234.9000 ;
	    RECT 1547.1000 234.7500 1548.9000 234.9000 ;
	    RECT 1513.5000 233.2500 1548.9000 234.7500 ;
	    RECT 1513.5000 233.1000 1515.3000 233.2500 ;
	    RECT 1547.1000 233.1000 1548.9000 233.2500 ;
	    RECT 32.7000 228.7500 34.5000 228.9000 ;
	    RECT 157.5000 228.7500 159.3000 228.9000 ;
	    RECT 32.7000 227.2500 159.3000 228.7500 ;
	    RECT 32.7000 227.1000 34.5000 227.2500 ;
	    RECT 157.5000 227.1000 159.3000 227.2500 ;
	    RECT 383.1000 228.7500 384.9000 228.9000 ;
	    RECT 421.5000 228.7500 423.3000 228.9000 ;
	    RECT 383.1000 227.2500 423.3000 228.7500 ;
	    RECT 383.1000 227.1000 384.9000 227.2500 ;
	    RECT 421.5000 227.1000 423.3000 227.2500 ;
	    RECT 495.9000 228.7500 497.7000 228.9000 ;
	    RECT 512.7000 228.7500 514.5000 228.9000 ;
	    RECT 495.9000 227.2500 514.5000 228.7500 ;
	    RECT 495.9000 227.1000 497.7000 227.2500 ;
	    RECT 512.7000 227.1000 514.5000 227.2500 ;
	    RECT 608.7000 228.7500 610.5000 228.9000 ;
	    RECT 632.7000 228.7500 634.5000 228.9000 ;
	    RECT 608.7000 227.2500 634.5000 228.7500 ;
	    RECT 608.7000 227.1000 610.5000 227.2500 ;
	    RECT 632.7000 227.1000 634.5000 227.2500 ;
	    RECT 644.7000 228.7500 646.5000 228.9000 ;
	    RECT 692.7000 228.7500 694.5000 228.9000 ;
	    RECT 644.7000 227.2500 694.5000 228.7500 ;
	    RECT 644.7000 227.1000 646.5000 227.2500 ;
	    RECT 692.7000 227.1000 694.5000 227.2500 ;
	    RECT 762.3000 228.7500 764.1000 228.9000 ;
	    RECT 908.7000 228.7500 910.5000 228.9000 ;
	    RECT 930.3000 228.7500 932.1000 228.9000 ;
	    RECT 762.3000 227.2500 932.1000 228.7500 ;
	    RECT 762.3000 227.1000 764.1000 227.2500 ;
	    RECT 908.7000 227.1000 910.5000 227.2500 ;
	    RECT 930.3000 227.1000 932.1000 227.2500 ;
	    RECT 1028.7001 228.7500 1030.5000 228.9000 ;
	    RECT 1081.5000 228.7500 1083.3000 228.9000 ;
	    RECT 1028.7001 227.2500 1083.3000 228.7500 ;
	    RECT 1028.7001 227.1000 1030.5000 227.2500 ;
	    RECT 1081.5000 227.1000 1083.3000 227.2500 ;
	    RECT 1196.7001 228.7500 1198.5000 228.9000 ;
	    RECT 1419.9000 228.7500 1421.7001 228.9000 ;
	    RECT 1196.7001 227.2500 1421.7001 228.7500 ;
	    RECT 1196.7001 227.1000 1198.5000 227.2500 ;
	    RECT 1419.9000 227.1000 1421.7001 227.2500 ;
	    RECT 318.3000 222.7500 320.1000 222.9000 ;
	    RECT 335.1000 222.7500 336.9000 222.9000 ;
	    RECT 318.3000 221.2500 336.9000 222.7500 ;
	    RECT 318.3000 221.1000 320.1000 221.2500 ;
	    RECT 335.1000 221.1000 336.9000 221.2500 ;
	    RECT 491.1000 222.7500 492.9000 222.9000 ;
	    RECT 498.3000 222.7500 500.1000 222.9000 ;
	    RECT 491.1000 221.2500 500.1000 222.7500 ;
	    RECT 491.1000 221.1000 492.9000 221.2500 ;
	    RECT 498.3000 221.1000 500.1000 221.2500 ;
	    RECT 529.5000 222.7500 531.3000 222.9000 ;
	    RECT 546.3000 222.7500 548.1000 222.9000 ;
	    RECT 529.5000 221.2500 548.1000 222.7500 ;
	    RECT 529.5000 221.1000 531.3000 221.2500 ;
	    RECT 546.3000 221.1000 548.1000 221.2500 ;
	    RECT 637.5000 222.7500 639.3000 222.9000 ;
	    RECT 675.9000 222.7500 677.7000 222.9000 ;
	    RECT 637.5000 221.2500 677.7000 222.7500 ;
	    RECT 637.5000 221.1000 639.3000 221.2500 ;
	    RECT 675.9000 221.1000 677.7000 221.2500 ;
	    RECT 683.1000 222.7500 684.9000 222.9000 ;
	    RECT 723.9000 222.7500 725.7000 222.9000 ;
	    RECT 752.7000 222.7500 754.5000 222.9000 ;
	    RECT 683.1000 221.2500 754.5000 222.7500 ;
	    RECT 683.1000 221.1000 684.9000 221.2500 ;
	    RECT 723.9000 221.1000 725.7000 221.2500 ;
	    RECT 752.7000 221.1000 754.5000 221.2500 ;
	    RECT 1033.5000 222.7500 1035.3000 222.9000 ;
	    RECT 1083.9000 222.7500 1085.7001 222.9000 ;
	    RECT 1033.5000 221.2500 1085.7001 222.7500 ;
	    RECT 1033.5000 221.1000 1035.3000 221.2500 ;
	    RECT 1083.9000 221.1000 1085.7001 221.2500 ;
	    RECT 1134.3000 222.7500 1136.1000 222.9000 ;
	    RECT 1146.3000 222.7500 1148.1000 222.9000 ;
	    RECT 1134.3000 221.2500 1148.1000 222.7500 ;
	    RECT 1134.3000 221.1000 1136.1000 221.2500 ;
	    RECT 1146.3000 221.1000 1148.1000 221.2500 ;
	    RECT 1155.9000 222.7500 1157.7001 222.9000 ;
	    RECT 1187.1000 222.7500 1188.9000 222.9000 ;
	    RECT 1155.9000 221.2500 1188.9000 222.7500 ;
	    RECT 1155.9000 221.1000 1157.7001 221.2500 ;
	    RECT 1187.1000 221.1000 1188.9000 221.2500 ;
	    RECT 1220.7001 222.7500 1222.5000 222.9000 ;
	    RECT 1259.1000 222.7500 1260.9000 222.9000 ;
	    RECT 1220.7001 221.2500 1260.9000 222.7500 ;
	    RECT 1220.7001 221.1000 1222.5000 221.2500 ;
	    RECT 1259.1000 221.1000 1260.9000 221.2500 ;
	    RECT 1290.3000 222.7500 1292.1000 222.9000 ;
	    RECT 1299.9000 222.7500 1301.7001 222.9000 ;
	    RECT 1290.3000 221.2500 1301.7001 222.7500 ;
	    RECT 1290.3000 221.1000 1292.1000 221.2500 ;
	    RECT 1299.9000 221.1000 1301.7001 221.2500 ;
	    RECT 1307.1000 222.7500 1308.9000 222.9000 ;
	    RECT 1429.5000 222.7500 1431.3000 222.9000 ;
	    RECT 1307.1000 221.2500 1431.3000 222.7500 ;
	    RECT 1307.1000 221.1000 1308.9000 221.2500 ;
	    RECT 1429.5000 221.1000 1431.3000 221.2500 ;
	    RECT 1434.3000 222.7500 1436.1000 222.9000 ;
	    RECT 1446.3000 222.7500 1448.1000 222.9000 ;
	    RECT 1434.3000 221.2500 1448.1000 222.7500 ;
	    RECT 1434.3000 221.1000 1436.1000 221.2500 ;
	    RECT 1446.3000 221.1000 1448.1000 221.2500 ;
	    RECT 1463.1000 222.7500 1464.9000 222.9000 ;
	    RECT 1513.5000 222.7500 1515.3000 222.9000 ;
	    RECT 1463.1000 221.2500 1515.3000 222.7500 ;
	    RECT 1463.1000 221.1000 1464.9000 221.2500 ;
	    RECT 1513.5000 221.1000 1515.3000 221.2500 ;
	    RECT 42.3000 216.7500 44.1000 216.9000 ;
	    RECT 71.1000 216.7500 72.9000 216.9000 ;
	    RECT 42.3000 215.2500 72.9000 216.7500 ;
	    RECT 42.3000 215.1000 44.1000 215.2500 ;
	    RECT 71.1000 215.1000 72.9000 215.2500 ;
	    RECT 193.5000 216.7500 195.3000 216.9000 ;
	    RECT 212.7000 216.7500 214.5000 216.9000 ;
	    RECT 231.9000 216.7500 233.7000 216.9000 ;
	    RECT 193.5000 215.2500 233.7000 216.7500 ;
	    RECT 193.5000 215.1000 195.3000 215.2500 ;
	    RECT 212.7000 215.1000 214.5000 215.2500 ;
	    RECT 231.9000 215.1000 233.7000 215.2500 ;
	    RECT 527.1000 216.7500 528.9000 216.9000 ;
	    RECT 563.1000 216.7500 564.9000 216.9000 ;
	    RECT 527.1000 215.2500 564.9000 216.7500 ;
	    RECT 527.1000 215.1000 528.9000 215.2500 ;
	    RECT 563.1000 215.1000 564.9000 215.2500 ;
	    RECT 572.7000 216.7500 574.5000 216.9000 ;
	    RECT 596.7000 216.7500 598.5000 216.9000 ;
	    RECT 572.7000 215.2500 598.5000 216.7500 ;
	    RECT 572.7000 215.1000 574.5000 215.2500 ;
	    RECT 596.7000 215.1000 598.5000 215.2500 ;
	    RECT 603.9000 216.7500 605.7000 216.9000 ;
	    RECT 627.9000 216.7500 629.7000 216.9000 ;
	    RECT 603.9000 215.2500 629.7000 216.7500 ;
	    RECT 603.9000 215.1000 605.7000 215.2500 ;
	    RECT 627.9000 215.1000 629.7000 215.2500 ;
	    RECT 649.5000 216.7500 651.3000 216.9000 ;
	    RECT 759.9000 216.7500 761.7000 216.9000 ;
	    RECT 649.5000 215.2500 761.7000 216.7500 ;
	    RECT 649.5000 215.1000 651.3000 215.2500 ;
	    RECT 759.9000 215.1000 761.7000 215.2500 ;
	    RECT 927.9000 216.7500 929.7000 216.9000 ;
	    RECT 959.1000 216.7500 960.9000 216.9000 ;
	    RECT 927.9000 215.2500 960.9000 216.7500 ;
	    RECT 927.9000 215.1000 929.7000 215.2500 ;
	    RECT 959.1000 215.1000 960.9000 215.2500 ;
	    RECT 1014.3000 216.7500 1016.1000 216.9000 ;
	    RECT 1059.9000 216.7500 1061.7001 216.9000 ;
	    RECT 1014.3000 215.2500 1061.7001 216.7500 ;
	    RECT 1014.3000 215.1000 1016.1000 215.2500 ;
	    RECT 1059.9000 215.1000 1061.7001 215.2500 ;
	    RECT 1100.7001 216.7500 1102.5000 216.9000 ;
	    RECT 1151.1000 216.7500 1152.9000 216.9000 ;
	    RECT 1100.7001 215.2500 1152.9000 216.7500 ;
	    RECT 1100.7001 215.1000 1102.5000 215.2500 ;
	    RECT 1151.1000 215.1000 1152.9000 215.2500 ;
	    RECT 1199.1000 216.7500 1200.9000 216.9000 ;
	    RECT 1266.3000 216.7500 1268.1000 216.9000 ;
	    RECT 1311.9000 216.7500 1313.7001 216.9000 ;
	    RECT 1376.7001 216.7500 1378.5000 216.9000 ;
	    RECT 1199.1000 215.2500 1378.5000 216.7500 ;
	    RECT 1199.1000 215.1000 1200.9000 215.2500 ;
	    RECT 1266.3000 215.1000 1268.1000 215.2500 ;
	    RECT 1311.9000 215.1000 1313.7001 215.2500 ;
	    RECT 1376.7001 215.1000 1378.5000 215.2500 ;
	    RECT 1434.3000 216.7500 1436.1000 216.9000 ;
	    RECT 1448.7001 216.7500 1450.5000 216.9000 ;
	    RECT 1434.3000 215.2500 1450.5000 216.7500 ;
	    RECT 1434.3000 215.1000 1436.1000 215.2500 ;
	    RECT 1448.7001 215.1000 1450.5000 215.2500 ;
	    RECT 1508.7001 216.7500 1510.5000 216.9000 ;
	    RECT 1518.3000 216.7500 1520.1000 216.9000 ;
	    RECT 1508.7001 215.2500 1520.1000 216.7500 ;
	    RECT 1508.7001 215.1000 1510.5000 215.2500 ;
	    RECT 1518.3000 215.1000 1520.1000 215.2500 ;
	    RECT 1542.3000 216.7500 1544.1000 216.9000 ;
	    RECT 1561.5000 216.7500 1563.3000 216.9000 ;
	    RECT 1542.3000 215.2500 1563.3000 216.7500 ;
	    RECT 1542.3000 215.1000 1544.1000 215.2500 ;
	    RECT 1561.5000 215.1000 1563.3000 215.2500 ;
	    RECT 167.1000 210.7500 168.9000 210.9000 ;
	    RECT 231.9000 210.7500 233.7000 210.9000 ;
	    RECT 167.1000 209.2500 233.7000 210.7500 ;
	    RECT 167.1000 209.1000 168.9000 209.2500 ;
	    RECT 231.9000 209.1000 233.7000 209.2500 ;
	    RECT 363.9000 210.7500 365.7000 210.9000 ;
	    RECT 380.7000 210.7500 382.5000 210.9000 ;
	    RECT 397.5000 210.7500 399.3000 210.9000 ;
	    RECT 404.7000 210.7500 406.5000 210.9000 ;
	    RECT 363.9000 209.2500 406.5000 210.7500 ;
	    RECT 363.9000 209.1000 365.7000 209.2500 ;
	    RECT 380.7000 209.1000 382.5000 209.2500 ;
	    RECT 397.5000 209.1000 399.3000 209.2500 ;
	    RECT 404.7000 209.1000 406.5000 209.2500 ;
	    RECT 685.5000 210.7500 687.3000 210.9000 ;
	    RECT 721.5000 210.7500 723.3000 210.9000 ;
	    RECT 685.5000 209.2500 723.3000 210.7500 ;
	    RECT 685.5000 209.1000 687.3000 209.2500 ;
	    RECT 721.5000 209.1000 723.3000 209.2500 ;
	    RECT 1203.9000 210.7500 1205.7001 210.9000 ;
	    RECT 1302.3000 210.7500 1304.1000 210.9000 ;
	    RECT 1347.9000 210.7500 1349.7001 210.9000 ;
	    RECT 1203.9000 209.2500 1349.7001 210.7500 ;
	    RECT 1203.9000 209.1000 1205.7001 209.2500 ;
	    RECT 1302.3000 209.1000 1304.1000 209.2500 ;
	    RECT 1347.9000 209.1000 1349.7001 209.2500 ;
	    RECT 1551.9000 210.7500 1553.7001 210.9000 ;
	    RECT 1561.5000 210.7500 1563.3000 210.9000 ;
	    RECT 1551.9000 209.2500 1563.3000 210.7500 ;
	    RECT 1551.9000 209.1000 1553.7001 209.2500 ;
	    RECT 1561.5000 209.1000 1563.3000 209.2500 ;
	    RECT 152.7000 204.7500 154.5000 204.9000 ;
	    RECT 179.1000 204.7500 180.9000 204.9000 ;
	    RECT 193.5000 204.7500 195.3000 204.9000 ;
	    RECT 152.7000 203.2500 195.3000 204.7500 ;
	    RECT 152.7000 203.1000 154.5000 203.2500 ;
	    RECT 179.1000 203.1000 180.9000 203.2500 ;
	    RECT 193.5000 203.1000 195.3000 203.2500 ;
	    RECT 558.3000 204.7500 560.1000 204.9000 ;
	    RECT 606.3000 204.7500 608.1000 204.9000 ;
	    RECT 558.3000 203.2500 608.1000 204.7500 ;
	    RECT 558.3000 203.1000 560.1000 203.2500 ;
	    RECT 606.3000 203.1000 608.1000 203.2500 ;
	    RECT 632.7000 204.7500 634.5000 204.9000 ;
	    RECT 654.3000 204.7500 656.1000 204.9000 ;
	    RECT 632.7000 203.2500 656.1000 204.7500 ;
	    RECT 632.7000 203.1000 634.5000 203.2500 ;
	    RECT 654.3000 203.1000 656.1000 203.2500 ;
	    RECT 793.5000 204.7500 795.3000 204.9000 ;
	    RECT 810.3000 204.7500 812.1000 204.9000 ;
	    RECT 829.5000 204.7500 831.3000 204.9000 ;
	    RECT 839.1000 204.7500 840.9000 204.9000 ;
	    RECT 858.3000 204.7500 860.1000 204.9000 ;
	    RECT 793.5000 203.2500 860.1000 204.7500 ;
	    RECT 793.5000 203.1000 795.3000 203.2500 ;
	    RECT 810.3000 203.1000 812.1000 203.2500 ;
	    RECT 829.5000 203.1000 831.3000 203.2500 ;
	    RECT 839.1000 203.1000 840.9000 203.2500 ;
	    RECT 858.3000 203.1000 860.1000 203.2500 ;
	    RECT 995.1000 204.7500 996.9000 204.9000 ;
	    RECT 1014.3000 204.7500 1016.1000 204.9000 ;
	    RECT 995.1000 203.2500 1016.1000 204.7500 ;
	    RECT 995.1000 203.1000 996.9000 203.2500 ;
	    RECT 1014.3000 203.1000 1016.1000 203.2500 ;
	    RECT 1023.9000 204.7500 1025.7001 204.9000 ;
	    RECT 1076.7001 204.7500 1078.5000 204.9000 ;
	    RECT 1107.9000 204.7500 1109.7001 204.9000 ;
	    RECT 1023.9000 203.2500 1109.7001 204.7500 ;
	    RECT 1023.9000 203.1000 1025.7001 203.2500 ;
	    RECT 1076.7001 203.1000 1078.5000 203.2500 ;
	    RECT 1107.9000 203.1000 1109.7001 203.2500 ;
	    RECT 1275.9000 204.7500 1277.7001 204.9000 ;
	    RECT 1343.1000 204.7500 1344.9000 204.9000 ;
	    RECT 1275.9000 203.2500 1344.9000 204.7500 ;
	    RECT 1275.9000 203.1000 1277.7001 203.2500 ;
	    RECT 1343.1000 203.1000 1344.9000 203.2500 ;
	    RECT 1443.9000 204.7500 1445.7001 204.9000 ;
	    RECT 1451.1000 204.7500 1452.9000 204.9000 ;
	    RECT 1475.1000 204.7500 1476.9000 204.9000 ;
	    RECT 1443.9000 203.2500 1476.9000 204.7500 ;
	    RECT 1443.9000 203.1000 1445.7001 203.2500 ;
	    RECT 1451.1000 203.1000 1452.9000 203.2500 ;
	    RECT 1475.1000 203.1000 1476.9000 203.2500 ;
	    RECT 1491.9000 204.7500 1493.7001 204.9000 ;
	    RECT 1511.1000 204.7500 1512.9000 204.9000 ;
	    RECT 1491.9000 203.2500 1512.9000 204.7500 ;
	    RECT 1491.9000 203.1000 1493.7001 203.2500 ;
	    RECT 1511.1000 203.1000 1512.9000 203.2500 ;
	    RECT 18.3000 198.7500 20.1000 198.9000 ;
	    RECT 54.3000 198.7500 56.1000 198.9000 ;
	    RECT 102.3000 198.7500 104.1000 198.9000 ;
	    RECT 123.9000 198.7500 125.7000 198.9000 ;
	    RECT 162.3000 198.7500 164.1000 198.9000 ;
	    RECT 215.1000 198.7500 216.9000 198.9000 ;
	    RECT 18.3000 197.2500 216.9000 198.7500 ;
	    RECT 18.3000 197.1000 20.1000 197.2500 ;
	    RECT 54.3000 197.1000 56.1000 197.2500 ;
	    RECT 102.3000 197.1000 104.1000 197.2500 ;
	    RECT 123.9000 197.1000 125.7000 197.2500 ;
	    RECT 162.3000 197.1000 164.1000 197.2500 ;
	    RECT 215.1000 197.1000 216.9000 197.2500 ;
	    RECT 577.5000 198.7500 579.3000 198.9000 ;
	    RECT 596.7000 198.7500 598.5000 198.9000 ;
	    RECT 577.5000 197.2500 598.5000 198.7500 ;
	    RECT 577.5000 197.1000 579.3000 197.2500 ;
	    RECT 596.7000 197.1000 598.5000 197.2500 ;
	    RECT 608.7000 198.7500 610.5000 198.9000 ;
	    RECT 637.5000 198.7500 639.3000 198.9000 ;
	    RECT 608.7000 197.2500 639.3000 198.7500 ;
	    RECT 608.7000 197.1000 610.5000 197.2500 ;
	    RECT 637.5000 197.1000 639.3000 197.2500 ;
	    RECT 757.5000 198.7500 759.3000 198.9000 ;
	    RECT 776.7000 198.7500 778.5000 198.9000 ;
	    RECT 757.5000 197.2500 778.5000 198.7500 ;
	    RECT 757.5000 197.1000 759.3000 197.2500 ;
	    RECT 776.7000 197.1000 778.5000 197.2500 ;
	    RECT 889.5000 198.7500 891.3000 198.9000 ;
	    RECT 911.1000 198.7500 912.9000 198.9000 ;
	    RECT 889.5000 197.2500 912.9000 198.7500 ;
	    RECT 889.5000 197.1000 891.3000 197.2500 ;
	    RECT 911.1000 197.1000 912.9000 197.2500 ;
	    RECT 961.5000 198.7500 963.3000 198.9000 ;
	    RECT 1153.5000 198.7500 1155.3000 198.9000 ;
	    RECT 961.5000 197.2500 1155.3000 198.7500 ;
	    RECT 961.5000 197.1000 963.3000 197.2500 ;
	    RECT 1153.5000 197.1000 1155.3000 197.2500 ;
	    RECT 1158.3000 198.7500 1160.1000 198.9000 ;
	    RECT 1208.7001 198.7500 1210.5000 198.9000 ;
	    RECT 1158.3000 197.2500 1210.5000 198.7500 ;
	    RECT 1158.3000 197.1000 1160.1000 197.2500 ;
	    RECT 1208.7001 197.1000 1210.5000 197.2500 ;
	    RECT 1215.9000 198.7500 1217.7001 198.9000 ;
	    RECT 1256.7001 198.7500 1258.5000 198.9000 ;
	    RECT 1215.9000 197.2500 1258.5000 198.7500 ;
	    RECT 1215.9000 197.1000 1217.7001 197.2500 ;
	    RECT 1256.7001 197.1000 1258.5000 197.2500 ;
	    RECT 1311.9000 198.7500 1313.7001 198.9000 ;
	    RECT 1374.3000 198.7500 1376.1000 198.9000 ;
	    RECT 1311.9000 197.2500 1376.1000 198.7500 ;
	    RECT 1311.9000 197.1000 1313.7001 197.2500 ;
	    RECT 1374.3000 197.1000 1376.1000 197.2500 ;
	    RECT 1398.3000 198.7500 1400.1000 198.9000 ;
	    RECT 1407.9000 198.7500 1409.7001 198.9000 ;
	    RECT 1467.9000 198.7500 1469.7001 198.9000 ;
	    RECT 1398.3000 197.2500 1469.7001 198.7500 ;
	    RECT 1398.3000 197.1000 1400.1000 197.2500 ;
	    RECT 1407.9000 197.1000 1409.7001 197.2500 ;
	    RECT 1467.9000 197.1000 1469.7001 197.2500 ;
	    RECT 1513.5000 198.7500 1515.3000 198.9000 ;
	    RECT 1530.3000 198.7500 1532.1000 198.9000 ;
	    RECT 1513.5000 197.2500 1532.1000 198.7500 ;
	    RECT 1513.5000 197.1000 1515.3000 197.2500 ;
	    RECT 1530.3000 197.1000 1532.1000 197.2500 ;
	    RECT 95.1000 192.7500 96.9000 192.9000 ;
	    RECT 119.1000 192.7500 120.9000 192.9000 ;
	    RECT 95.1000 191.2500 120.9000 192.7500 ;
	    RECT 95.1000 191.1000 96.9000 191.2500 ;
	    RECT 119.1000 191.1000 120.9000 191.2500 ;
	    RECT 572.7000 192.7500 574.5000 192.9000 ;
	    RECT 579.9000 192.7500 581.7000 192.9000 ;
	    RECT 572.7000 191.2500 581.7000 192.7500 ;
	    RECT 572.7000 191.1000 574.5000 191.2500 ;
	    RECT 579.9000 191.1000 581.7000 191.2500 ;
	    RECT 625.5000 192.7500 627.3000 192.9000 ;
	    RECT 687.9000 192.7500 689.7000 192.9000 ;
	    RECT 625.5000 191.2500 689.7000 192.7500 ;
	    RECT 625.5000 191.1000 627.3000 191.2500 ;
	    RECT 687.9000 191.1000 689.7000 191.2500 ;
	    RECT 915.9000 192.7500 917.7000 192.9000 ;
	    RECT 966.3000 192.7500 968.1000 192.9000 ;
	    RECT 1033.5000 192.7500 1035.3000 192.9000 ;
	    RECT 1050.3000 192.7500 1052.1000 192.9000 ;
	    RECT 915.9000 191.2500 1052.1000 192.7500 ;
	    RECT 915.9000 191.1000 917.7000 191.2500 ;
	    RECT 966.3000 191.1000 968.1000 191.2500 ;
	    RECT 1033.5000 191.1000 1035.3000 191.2500 ;
	    RECT 1050.3000 191.1000 1052.1000 191.2500 ;
	    RECT 1076.7001 192.7500 1078.5000 192.9000 ;
	    RECT 1105.5000 192.7500 1107.3000 192.9000 ;
	    RECT 1076.7001 191.2500 1107.3000 192.7500 ;
	    RECT 1076.7001 191.1000 1078.5000 191.2500 ;
	    RECT 1105.5000 191.1000 1107.3000 191.2500 ;
	    RECT 1110.3000 192.7500 1112.1000 192.9000 ;
	    RECT 1141.5000 192.7500 1143.3000 192.9000 ;
	    RECT 1110.3000 191.2500 1143.3000 192.7500 ;
	    RECT 1110.3000 191.1000 1112.1000 191.2500 ;
	    RECT 1141.5000 191.1000 1143.3000 191.2500 ;
	    RECT 1153.5000 192.7500 1155.3000 192.9000 ;
	    RECT 1309.5000 192.7500 1311.3000 192.9000 ;
	    RECT 1153.5000 191.2500 1311.3000 192.7500 ;
	    RECT 1153.5000 191.1000 1155.3000 191.2500 ;
	    RECT 1309.5000 191.1000 1311.3000 191.2500 ;
	    RECT 1335.9000 192.7500 1337.7001 192.9000 ;
	    RECT 1453.5000 192.7500 1455.3000 192.9000 ;
	    RECT 1479.9000 192.7500 1481.7001 192.9000 ;
	    RECT 1335.9000 191.2500 1481.7001 192.7500 ;
	    RECT 1335.9000 191.1000 1337.7001 191.2500 ;
	    RECT 1453.5000 191.1000 1455.3000 191.2500 ;
	    RECT 1479.9000 191.1000 1481.7001 191.2500 ;
	    RECT 207.9000 186.7500 209.7000 186.9000 ;
	    RECT 246.3000 186.7500 248.1000 186.9000 ;
	    RECT 207.9000 185.2500 248.1000 186.7500 ;
	    RECT 207.9000 185.1000 209.7000 185.2500 ;
	    RECT 246.3000 185.1000 248.1000 185.2500 ;
	    RECT 575.1000 186.7500 576.9000 186.9000 ;
	    RECT 625.5000 186.7500 627.3000 186.9000 ;
	    RECT 575.1000 185.2500 627.3000 186.7500 ;
	    RECT 575.1000 185.1000 576.9000 185.2500 ;
	    RECT 625.5000 185.1000 627.3000 185.2500 ;
	    RECT 853.5000 186.7500 855.3000 186.9000 ;
	    RECT 908.7000 186.7500 910.5000 186.9000 ;
	    RECT 853.5000 185.2500 910.5000 186.7500 ;
	    RECT 853.5000 185.1000 855.3000 185.2500 ;
	    RECT 908.7000 185.1000 910.5000 185.2500 ;
	    RECT 1002.3000 186.7500 1004.1000 186.9000 ;
	    RECT 1045.5000 186.7500 1047.3000 186.9000 ;
	    RECT 1002.3000 185.2500 1047.3000 186.7500 ;
	    RECT 1002.3000 185.1000 1004.1000 185.2500 ;
	    RECT 1045.5000 185.1000 1047.3000 185.2500 ;
	    RECT 1112.7001 186.7500 1114.5000 186.9000 ;
	    RECT 1163.1000 186.7500 1164.9000 186.9000 ;
	    RECT 1203.9000 186.7500 1205.7001 186.9000 ;
	    RECT 1225.5000 186.7500 1227.3000 186.9000 ;
	    RECT 1112.7001 185.2500 1227.3000 186.7500 ;
	    RECT 1112.7001 185.1000 1114.5000 185.2500 ;
	    RECT 1163.1000 185.1000 1164.9000 185.2500 ;
	    RECT 1203.9000 185.1000 1205.7001 185.2500 ;
	    RECT 1225.5000 185.1000 1227.3000 185.2500 ;
	    RECT 1232.7001 186.7500 1234.5000 186.9000 ;
	    RECT 1285.5000 186.7500 1287.3000 186.9000 ;
	    RECT 1232.7001 185.2500 1287.3000 186.7500 ;
	    RECT 1232.7001 185.1000 1234.5000 185.2500 ;
	    RECT 1285.5000 185.1000 1287.3000 185.2500 ;
	    RECT 1359.9000 186.7500 1361.7001 186.9000 ;
	    RECT 1542.3000 186.7500 1544.1000 186.9000 ;
	    RECT 1359.9000 185.2500 1544.1000 186.7500 ;
	    RECT 1359.9000 185.1000 1361.7001 185.2500 ;
	    RECT 1542.3000 185.1000 1544.1000 185.2500 ;
	    RECT 231.9000 180.7500 233.7000 180.9000 ;
	    RECT 363.9000 180.7500 365.7000 180.9000 ;
	    RECT 431.1000 180.7500 432.9000 180.9000 ;
	    RECT 231.9000 179.2500 432.9000 180.7500 ;
	    RECT 231.9000 179.1000 233.7000 179.2500 ;
	    RECT 363.9000 179.1000 365.7000 179.2500 ;
	    RECT 431.1000 179.1000 432.9000 179.2500 ;
	    RECT 908.7000 180.7500 910.5000 180.9000 ;
	    RECT 920.7000 180.7500 922.5000 180.9000 ;
	    RECT 908.7000 179.2500 922.5000 180.7500 ;
	    RECT 908.7000 179.1000 910.5000 179.2500 ;
	    RECT 920.7000 179.1000 922.5000 179.2500 ;
	    RECT 930.3000 180.7500 932.1000 180.9000 ;
	    RECT 963.9000 180.7500 965.7000 180.9000 ;
	    RECT 930.3000 179.2500 965.7000 180.7500 ;
	    RECT 930.3000 179.1000 932.1000 179.2500 ;
	    RECT 963.9000 179.1000 965.7000 179.2500 ;
	    RECT 1014.3000 180.7500 1016.1000 180.9000 ;
	    RECT 1098.3000 180.7500 1100.1000 180.9000 ;
	    RECT 1119.9000 180.7500 1121.7001 180.9000 ;
	    RECT 1014.3000 179.2500 1121.7001 180.7500 ;
	    RECT 1014.3000 179.1000 1016.1000 179.2500 ;
	    RECT 1098.3000 179.1000 1100.1000 179.2500 ;
	    RECT 1119.9000 179.1000 1121.7001 179.2500 ;
	    RECT 1163.1000 180.7500 1164.9000 180.9000 ;
	    RECT 1187.1000 180.7500 1188.9000 180.9000 ;
	    RECT 1163.1000 179.2500 1188.9000 180.7500 ;
	    RECT 1163.1000 179.1000 1164.9000 179.2500 ;
	    RECT 1187.1000 179.1000 1188.9000 179.2500 ;
	    RECT 1347.9000 180.7500 1349.7001 180.9000 ;
	    RECT 1400.7001 180.7500 1402.5000 180.9000 ;
	    RECT 1472.7001 180.7500 1474.5000 180.9000 ;
	    RECT 1347.9000 179.2500 1474.5000 180.7500 ;
	    RECT 1347.9000 179.1000 1349.7001 179.2500 ;
	    RECT 1400.7001 179.1000 1402.5000 179.2500 ;
	    RECT 1472.7001 179.1000 1474.5000 179.2500 ;
	    RECT 342.3000 174.7500 344.1000 174.9000 ;
	    RECT 457.5000 174.7500 459.3000 174.9000 ;
	    RECT 342.3000 173.2500 459.3000 174.7500 ;
	    RECT 342.3000 173.1000 344.1000 173.2500 ;
	    RECT 457.5000 173.1000 459.3000 173.2500 ;
	    RECT 721.5000 174.7500 723.3000 174.9000 ;
	    RECT 743.1000 174.7500 744.9000 174.9000 ;
	    RECT 721.5000 173.2500 744.9000 174.7500 ;
	    RECT 721.5000 173.1000 723.3000 173.2500 ;
	    RECT 743.1000 173.1000 744.9000 173.2500 ;
	    RECT 959.1000 174.7500 960.9000 174.9000 ;
	    RECT 992.7000 174.7500 994.5000 174.9000 ;
	    RECT 959.1000 173.2500 994.5000 174.7500 ;
	    RECT 959.1000 173.1000 960.9000 173.2500 ;
	    RECT 992.7000 173.1000 994.5000 173.2500 ;
	    RECT 1040.7001 174.7500 1042.5000 174.9000 ;
	    RECT 1067.1000 174.7500 1068.9000 174.9000 ;
	    RECT 1040.7001 173.2500 1068.9000 174.7500 ;
	    RECT 1040.7001 173.1000 1042.5000 173.2500 ;
	    RECT 1067.1000 173.1000 1068.9000 173.2500 ;
	    RECT 1110.3000 174.7500 1112.1000 174.9000 ;
	    RECT 1158.3000 174.7500 1160.1000 174.9000 ;
	    RECT 1110.3000 173.2500 1160.1000 174.7500 ;
	    RECT 1110.3000 173.1000 1112.1000 173.2500 ;
	    RECT 1158.3000 173.1000 1160.1000 173.2500 ;
	    RECT 1179.9000 174.7500 1181.7001 174.9000 ;
	    RECT 1251.9000 174.7500 1253.7001 174.9000 ;
	    RECT 1280.7001 174.7500 1282.5000 174.9000 ;
	    RECT 1179.9000 173.2500 1282.5000 174.7500 ;
	    RECT 1179.9000 173.1000 1181.7001 173.2500 ;
	    RECT 1251.9000 173.1000 1253.7001 173.2500 ;
	    RECT 1280.7001 173.1000 1282.5000 173.2500 ;
	    RECT 1374.3000 174.7500 1376.1000 174.9000 ;
	    RECT 1386.3000 174.7500 1388.1000 174.9000 ;
	    RECT 1374.3000 173.2500 1388.1000 174.7500 ;
	    RECT 1374.3000 173.1000 1376.1000 173.2500 ;
	    RECT 1386.3000 173.1000 1388.1000 173.2500 ;
	    RECT 1398.3000 174.7500 1400.1000 174.9000 ;
	    RECT 1434.3000 174.7500 1436.1000 174.9000 ;
	    RECT 1398.3000 173.2500 1436.1000 174.7500 ;
	    RECT 1398.3000 173.1000 1400.1000 173.2500 ;
	    RECT 1434.3000 173.1000 1436.1000 173.2500 ;
	    RECT 1441.5000 174.7500 1443.3000 174.9000 ;
	    RECT 1470.3000 174.7500 1472.1000 174.9000 ;
	    RECT 1441.5000 173.2500 1472.1000 174.7500 ;
	    RECT 1441.5000 173.1000 1443.3000 173.2500 ;
	    RECT 1470.3000 173.1000 1472.1000 173.2500 ;
	    RECT 1491.9000 174.7500 1493.7001 174.9000 ;
	    RECT 1515.9000 174.7500 1517.7001 174.9000 ;
	    RECT 1491.9000 173.2500 1517.7001 174.7500 ;
	    RECT 1491.9000 173.1000 1493.7001 173.2500 ;
	    RECT 1515.9000 173.1000 1517.7001 173.2500 ;
	    RECT 39.9000 168.7500 41.7000 168.9000 ;
	    RECT 47.1000 168.7500 48.9000 168.9000 ;
	    RECT 39.9000 167.2500 48.9000 168.7500 ;
	    RECT 39.9000 167.1000 41.7000 167.2500 ;
	    RECT 47.1000 167.1000 48.9000 167.2500 ;
	    RECT 195.9000 168.7500 197.7000 168.9000 ;
	    RECT 227.1000 168.7500 228.9000 168.9000 ;
	    RECT 251.1000 168.7500 252.9000 168.9000 ;
	    RECT 195.9000 167.2500 252.9000 168.7500 ;
	    RECT 195.9000 167.1000 197.7000 167.2500 ;
	    RECT 227.1000 167.1000 228.9000 167.2500 ;
	    RECT 251.1000 167.1000 252.9000 167.2500 ;
	    RECT 402.3000 168.7500 404.1000 168.9000 ;
	    RECT 435.9000 168.7500 437.7000 168.9000 ;
	    RECT 402.3000 167.2500 437.7000 168.7500 ;
	    RECT 402.3000 167.1000 404.1000 167.2500 ;
	    RECT 435.9000 167.1000 437.7000 167.2500 ;
	    RECT 649.5000 168.7500 651.3000 168.9000 ;
	    RECT 723.9000 168.7500 725.7000 168.9000 ;
	    RECT 649.5000 167.2500 725.7000 168.7500 ;
	    RECT 649.5000 167.1000 651.3000 167.2500 ;
	    RECT 723.9000 167.1000 725.7000 167.2500 ;
	    RECT 1095.9000 168.7500 1097.7001 168.9000 ;
	    RECT 1107.9000 168.7500 1109.7001 168.9000 ;
	    RECT 1095.9000 167.2500 1109.7001 168.7500 ;
	    RECT 1095.9000 167.1000 1097.7001 167.2500 ;
	    RECT 1107.9000 167.1000 1109.7001 167.2500 ;
	    RECT 1134.3000 168.7500 1136.1000 168.9000 ;
	    RECT 1146.3000 168.7500 1148.1000 168.9000 ;
	    RECT 1134.3000 167.2500 1148.1000 168.7500 ;
	    RECT 1134.3000 167.1000 1136.1000 167.2500 ;
	    RECT 1146.3000 167.1000 1148.1000 167.2500 ;
	    RECT 1160.7001 168.7500 1162.5000 168.9000 ;
	    RECT 1172.7001 168.7500 1174.5000 168.9000 ;
	    RECT 1160.7001 167.2500 1174.5000 168.7500 ;
	    RECT 1160.7001 167.1000 1162.5000 167.2500 ;
	    RECT 1172.7001 167.1000 1174.5000 167.2500 ;
	    RECT 1196.7001 168.7500 1198.5000 168.9000 ;
	    RECT 1223.1000 168.7500 1224.9000 168.9000 ;
	    RECT 1196.7001 167.2500 1224.9000 168.7500 ;
	    RECT 1196.7001 167.1000 1198.5000 167.2500 ;
	    RECT 1223.1000 167.1000 1224.9000 167.2500 ;
	    RECT 1369.5000 168.7500 1371.3000 168.9000 ;
	    RECT 1374.3000 168.7500 1376.1000 168.9000 ;
	    RECT 1369.5000 167.2500 1376.1000 168.7500 ;
	    RECT 1369.5000 167.1000 1371.3000 167.2500 ;
	    RECT 1374.3000 167.1000 1376.1000 167.2500 ;
	    RECT 1395.9000 168.7500 1397.7001 168.9000 ;
	    RECT 1429.5000 168.7500 1431.3000 168.9000 ;
	    RECT 1395.9000 167.2500 1431.3000 168.7500 ;
	    RECT 1395.9000 167.1000 1397.7001 167.2500 ;
	    RECT 1429.5000 167.1000 1431.3000 167.2500 ;
	    RECT 1443.9000 168.7500 1445.7001 168.9000 ;
	    RECT 1455.9000 168.7500 1457.7001 168.9000 ;
	    RECT 1443.9000 167.2500 1457.7001 168.7500 ;
	    RECT 1443.9000 167.1000 1445.7001 167.2500 ;
	    RECT 1455.9000 167.1000 1457.7001 167.2500 ;
	    RECT 15.9000 162.7500 17.7000 162.9000 ;
	    RECT 32.7000 162.7500 34.5000 162.9000 ;
	    RECT 15.9000 161.2500 34.5000 162.7500 ;
	    RECT 15.9000 161.1000 17.7000 161.2500 ;
	    RECT 32.7000 161.1000 34.5000 161.2500 ;
	    RECT 116.7000 162.7500 118.5000 162.9000 ;
	    RECT 191.1000 162.7500 192.9000 162.9000 ;
	    RECT 116.7000 161.2500 192.9000 162.7500 ;
	    RECT 116.7000 161.1000 118.5000 161.2500 ;
	    RECT 191.1000 161.1000 192.9000 161.2500 ;
	    RECT 248.7000 162.7500 250.5000 162.9000 ;
	    RECT 272.7000 162.7500 274.5000 162.9000 ;
	    RECT 248.7000 161.2500 274.5000 162.7500 ;
	    RECT 248.7000 161.1000 250.5000 161.2500 ;
	    RECT 272.7000 161.1000 274.5000 161.2500 ;
	    RECT 577.5000 162.7500 579.3000 162.9000 ;
	    RECT 608.7000 162.7500 610.5000 162.9000 ;
	    RECT 577.5000 161.2500 610.5000 162.7500 ;
	    RECT 577.5000 161.1000 579.3000 161.2500 ;
	    RECT 608.7000 161.1000 610.5000 161.2500 ;
	    RECT 1040.7001 162.7500 1042.5000 162.9000 ;
	    RECT 1112.7001 162.7500 1114.5000 162.9000 ;
	    RECT 1040.7001 161.2500 1114.5000 162.7500 ;
	    RECT 1040.7001 161.1000 1042.5000 161.2500 ;
	    RECT 1112.7001 161.1000 1114.5000 161.2500 ;
	    RECT 1141.5000 162.7500 1143.3000 162.9000 ;
	    RECT 1155.9000 162.7500 1157.7001 162.9000 ;
	    RECT 1141.5000 161.2500 1157.7001 162.7500 ;
	    RECT 1141.5000 161.1000 1143.3000 161.2500 ;
	    RECT 1155.9000 161.1000 1157.7001 161.2500 ;
	    RECT 1172.7001 162.7500 1174.5000 162.9000 ;
	    RECT 1184.7001 162.7500 1186.5000 162.9000 ;
	    RECT 1172.7001 161.2500 1186.5000 162.7500 ;
	    RECT 1172.7001 161.1000 1174.5000 161.2500 ;
	    RECT 1184.7001 161.1000 1186.5000 161.2500 ;
	    RECT 1343.1000 162.7500 1344.9000 162.9000 ;
	    RECT 1359.9000 162.7500 1361.7001 162.9000 ;
	    RECT 1343.1000 161.2500 1361.7001 162.7500 ;
	    RECT 1343.1000 161.1000 1344.9000 161.2500 ;
	    RECT 1359.9000 161.1000 1361.7001 161.2500 ;
	    RECT 1441.5000 162.7500 1443.3000 162.9000 ;
	    RECT 1448.7001 162.7500 1450.5000 162.9000 ;
	    RECT 1441.5000 161.2500 1450.5000 162.7500 ;
	    RECT 1441.5000 161.1000 1443.3000 161.2500 ;
	    RECT 1448.7001 161.1000 1450.5000 161.2500 ;
	    RECT 1544.7001 162.7500 1546.5000 162.9000 ;
	    RECT 1556.7001 162.7500 1558.5000 162.9000 ;
	    RECT 1544.7001 161.2500 1558.5000 162.7500 ;
	    RECT 1544.7001 161.1000 1546.5000 161.2500 ;
	    RECT 1556.7001 161.1000 1558.5000 161.2500 ;
	    RECT 191.1000 156.7500 192.9000 156.9000 ;
	    RECT 253.5000 156.7500 255.3000 156.9000 ;
	    RECT 191.1000 155.2500 255.3000 156.7500 ;
	    RECT 191.1000 155.1000 192.9000 155.2500 ;
	    RECT 253.5000 155.1000 255.3000 155.2500 ;
	    RECT 551.1000 156.7500 552.9000 156.9000 ;
	    RECT 603.9000 156.7500 605.7000 156.9000 ;
	    RECT 673.5000 156.7500 675.3000 156.9000 ;
	    RECT 726.3000 156.7500 728.1000 156.9000 ;
	    RECT 731.1000 156.7500 732.9000 156.9000 ;
	    RECT 755.1000 156.7500 756.9000 156.9000 ;
	    RECT 551.1000 155.2500 756.9000 156.7500 ;
	    RECT 551.1000 155.1000 552.9000 155.2500 ;
	    RECT 603.9000 155.1000 605.7000 155.2500 ;
	    RECT 673.5000 155.1000 675.3000 155.2500 ;
	    RECT 726.3000 155.1000 728.1000 155.2500 ;
	    RECT 731.1000 155.1000 732.9000 155.2500 ;
	    RECT 755.1000 155.1000 756.9000 155.2500 ;
	    RECT 882.3000 156.7500 884.1000 156.9000 ;
	    RECT 935.1000 156.7500 936.9000 156.9000 ;
	    RECT 882.3000 155.2500 936.9000 156.7500 ;
	    RECT 882.3000 155.1000 884.1000 155.2500 ;
	    RECT 935.1000 155.1000 936.9000 155.2500 ;
	    RECT 968.7000 156.7500 970.5000 156.9000 ;
	    RECT 1105.5000 156.7500 1107.3000 156.9000 ;
	    RECT 968.7000 155.2500 1107.3000 156.7500 ;
	    RECT 968.7000 155.1000 970.5000 155.2500 ;
	    RECT 1105.5000 155.1000 1107.3000 155.2500 ;
	    RECT 1131.9000 156.7500 1133.7001 156.9000 ;
	    RECT 1196.7001 156.7500 1198.5000 156.9000 ;
	    RECT 1131.9000 155.2500 1198.5000 156.7500 ;
	    RECT 1131.9000 155.1000 1133.7001 155.2500 ;
	    RECT 1196.7001 155.1000 1198.5000 155.2500 ;
	    RECT 1479.9000 156.7500 1481.7001 156.9000 ;
	    RECT 1523.1000 156.7500 1524.9000 156.9000 ;
	    RECT 1479.9000 155.2500 1524.9000 156.7500 ;
	    RECT 1479.9000 155.1000 1481.7001 155.2500 ;
	    RECT 1523.1000 155.1000 1524.9000 155.2500 ;
	    RECT 135.9000 150.7500 137.7000 150.9000 ;
	    RECT 174.3000 150.7500 176.1000 150.9000 ;
	    RECT 135.9000 149.2500 176.1000 150.7500 ;
	    RECT 135.9000 149.1000 137.7000 149.2500 ;
	    RECT 174.3000 149.1000 176.1000 149.2500 ;
	    RECT 323.1000 150.7500 324.9000 150.9000 ;
	    RECT 335.1000 150.7500 336.9000 150.9000 ;
	    RECT 351.9000 150.7500 353.7000 150.9000 ;
	    RECT 416.7000 150.7500 418.5000 150.9000 ;
	    RECT 431.1000 150.7500 432.9000 150.9000 ;
	    RECT 323.1000 149.2500 432.9000 150.7500 ;
	    RECT 323.1000 149.1000 324.9000 149.2500 ;
	    RECT 335.1000 149.1000 336.9000 149.2500 ;
	    RECT 351.9000 149.1000 353.7000 149.2500 ;
	    RECT 416.7000 149.1000 418.5000 149.2500 ;
	    RECT 431.1000 149.1000 432.9000 149.2500 ;
	    RECT 783.9000 150.7500 785.7000 150.9000 ;
	    RECT 822.3000 150.7500 824.1000 150.9000 ;
	    RECT 783.9000 149.2500 824.1000 150.7500 ;
	    RECT 783.9000 149.1000 785.7000 149.2500 ;
	    RECT 822.3000 149.1000 824.1000 149.2500 ;
	    RECT 906.3000 150.7500 908.1000 150.9000 ;
	    RECT 1002.3000 150.7500 1004.1000 150.9000 ;
	    RECT 906.3000 149.2500 1004.1000 150.7500 ;
	    RECT 906.3000 149.1000 908.1000 149.2500 ;
	    RECT 1002.3000 149.1000 1004.1000 149.2500 ;
	    RECT 1170.3000 150.7500 1172.1000 150.9000 ;
	    RECT 1211.1000 150.7500 1212.9000 150.9000 ;
	    RECT 1170.3000 149.2500 1212.9000 150.7500 ;
	    RECT 1170.3000 149.1000 1172.1000 149.2500 ;
	    RECT 1211.1000 149.1000 1212.9000 149.2500 ;
	    RECT 1218.3000 150.7500 1220.1000 150.9000 ;
	    RECT 1307.1000 150.7500 1308.9000 150.9000 ;
	    RECT 1338.3000 150.7500 1340.1000 150.9000 ;
	    RECT 1218.3000 149.2500 1340.1000 150.7500 ;
	    RECT 1218.3000 149.1000 1220.1000 149.2500 ;
	    RECT 1307.1000 149.1000 1308.9000 149.2500 ;
	    RECT 1338.3000 149.1000 1340.1000 149.2500 ;
	    RECT 1379.1000 150.7500 1380.9000 150.9000 ;
	    RECT 1395.9000 150.7500 1397.7001 150.9000 ;
	    RECT 1379.1000 149.2500 1397.7001 150.7500 ;
	    RECT 1379.1000 149.1000 1380.9000 149.2500 ;
	    RECT 1395.9000 149.1000 1397.7001 149.2500 ;
	    RECT 1422.3000 150.7500 1424.1000 150.9000 ;
	    RECT 1446.3000 150.7500 1448.1000 150.9000 ;
	    RECT 1422.3000 149.2500 1448.1000 150.7500 ;
	    RECT 1422.3000 149.1000 1424.1000 149.2500 ;
	    RECT 1446.3000 149.1000 1448.1000 149.2500 ;
	    RECT 92.7000 144.7500 94.5000 144.9000 ;
	    RECT 145.5000 144.7500 147.3000 144.9000 ;
	    RECT 92.7000 143.2500 147.3000 144.7500 ;
	    RECT 92.7000 143.1000 94.5000 143.2500 ;
	    RECT 145.5000 143.1000 147.3000 143.2500 ;
	    RECT 150.3000 144.7500 152.1000 144.9000 ;
	    RECT 195.9000 144.7500 197.7000 144.9000 ;
	    RECT 150.3000 143.2500 197.7000 144.7500 ;
	    RECT 150.3000 143.1000 152.1000 143.2500 ;
	    RECT 195.9000 143.1000 197.7000 143.2500 ;
	    RECT 291.9000 144.7500 293.7000 144.9000 ;
	    RECT 347.1000 144.7500 348.9000 144.9000 ;
	    RECT 291.9000 143.2500 348.9000 144.7500 ;
	    RECT 291.9000 143.1000 293.7000 143.2500 ;
	    RECT 347.1000 143.1000 348.9000 143.2500 ;
	    RECT 495.9000 144.7500 497.7000 144.9000 ;
	    RECT 546.3000 144.7500 548.1000 144.9000 ;
	    RECT 495.9000 143.2500 548.1000 144.7500 ;
	    RECT 495.9000 143.1000 497.7000 143.2500 ;
	    RECT 546.3000 143.1000 548.1000 143.2500 ;
	    RECT 992.7000 144.7500 994.5000 144.9000 ;
	    RECT 1023.9000 144.7500 1025.7001 144.9000 ;
	    RECT 992.7000 143.2500 1025.7001 144.7500 ;
	    RECT 992.7000 143.1000 994.5000 143.2500 ;
	    RECT 1023.9000 143.1000 1025.7001 143.2500 ;
	    RECT 1074.3000 144.7500 1076.1000 144.9000 ;
	    RECT 1088.7001 144.7500 1090.5000 144.9000 ;
	    RECT 1074.3000 143.2500 1090.5000 144.7500 ;
	    RECT 1074.3000 143.1000 1076.1000 143.2500 ;
	    RECT 1088.7001 143.1000 1090.5000 143.2500 ;
	    RECT 1103.1000 144.7500 1104.9000 144.9000 ;
	    RECT 1151.1000 144.7500 1152.9000 144.9000 ;
	    RECT 1103.1000 143.2500 1152.9000 144.7500 ;
	    RECT 1103.1000 143.1000 1104.9000 143.2500 ;
	    RECT 1151.1000 143.1000 1152.9000 143.2500 ;
	    RECT 1211.1000 144.7500 1212.9000 144.9000 ;
	    RECT 1251.9000 144.7500 1253.7001 144.9000 ;
	    RECT 1211.1000 143.2500 1253.7001 144.7500 ;
	    RECT 1211.1000 143.1000 1212.9000 143.2500 ;
	    RECT 1251.9000 143.1000 1253.7001 143.2500 ;
	    RECT 1331.1000 144.7500 1332.9000 144.9000 ;
	    RECT 1376.7001 144.7500 1378.5000 144.9000 ;
	    RECT 1331.1000 143.2500 1378.5000 144.7500 ;
	    RECT 1331.1000 143.1000 1332.9000 143.2500 ;
	    RECT 1376.7001 143.1000 1378.5000 143.2500 ;
	    RECT 1412.7001 144.7500 1414.5000 144.9000 ;
	    RECT 1424.7001 144.7500 1426.5000 144.9000 ;
	    RECT 1412.7001 143.2500 1426.5000 144.7500 ;
	    RECT 1412.7001 143.1000 1414.5000 143.2500 ;
	    RECT 1424.7001 143.1000 1426.5000 143.2500 ;
	    RECT 1443.9000 144.7500 1445.7001 144.9000 ;
	    RECT 1472.7001 144.7500 1474.5000 144.9000 ;
	    RECT 1443.9000 143.2500 1474.5000 144.7500 ;
	    RECT 1443.9000 143.1000 1445.7001 143.2500 ;
	    RECT 1472.7001 143.1000 1474.5000 143.2500 ;
	    RECT 1482.3000 144.7500 1484.1000 144.9000 ;
	    RECT 1494.3000 144.7500 1496.1000 144.9000 ;
	    RECT 1482.3000 143.2500 1496.1000 144.7500 ;
	    RECT 1482.3000 143.1000 1484.1000 143.2500 ;
	    RECT 1494.3000 143.1000 1496.1000 143.2500 ;
	    RECT 529.5000 138.7500 531.3000 138.9000 ;
	    RECT 536.7000 138.7500 538.5000 138.9000 ;
	    RECT 529.5000 137.2500 538.5000 138.7500 ;
	    RECT 529.5000 137.1000 531.3000 137.2500 ;
	    RECT 536.7000 137.1000 538.5000 137.2500 ;
	    RECT 699.9000 138.7500 701.7000 138.9000 ;
	    RECT 719.1000 138.7500 720.9000 138.9000 ;
	    RECT 699.9000 137.2500 720.9000 138.7500 ;
	    RECT 699.9000 137.1000 701.7000 137.2500 ;
	    RECT 719.1000 137.1000 720.9000 137.2500 ;
	    RECT 853.5000 138.7500 855.3000 138.9000 ;
	    RECT 860.7000 138.7500 862.5000 138.9000 ;
	    RECT 853.5000 137.2500 862.5000 138.7500 ;
	    RECT 853.5000 137.1000 855.3000 137.2500 ;
	    RECT 860.7000 137.1000 862.5000 137.2500 ;
	    RECT 959.1000 138.7500 960.9000 138.9000 ;
	    RECT 1028.7001 138.7500 1030.5000 138.9000 ;
	    RECT 1074.3000 138.7500 1076.1000 138.9000 ;
	    RECT 959.1000 137.2500 1076.1000 138.7500 ;
	    RECT 959.1000 137.1000 960.9000 137.2500 ;
	    RECT 1028.7001 137.1000 1030.5000 137.2500 ;
	    RECT 1074.3000 137.1000 1076.1000 137.2500 ;
	    RECT 1079.1000 138.7500 1080.9000 138.9000 ;
	    RECT 1103.1000 138.7500 1104.9000 138.9000 ;
	    RECT 1172.7001 138.7500 1174.5000 138.9000 ;
	    RECT 1079.1000 137.2500 1174.5000 138.7500 ;
	    RECT 1079.1000 137.1000 1080.9000 137.2500 ;
	    RECT 1103.1000 137.1000 1104.9000 137.2500 ;
	    RECT 1172.7001 137.1000 1174.5000 137.2500 ;
	    RECT 1213.5000 138.7500 1215.3000 138.9000 ;
	    RECT 1254.3000 138.7500 1256.1000 138.9000 ;
	    RECT 1213.5000 137.2500 1256.1000 138.7500 ;
	    RECT 1213.5000 137.1000 1215.3000 137.2500 ;
	    RECT 1254.3000 137.1000 1256.1000 137.2500 ;
	    RECT 1259.1000 138.7500 1260.9000 138.9000 ;
	    RECT 1386.3000 138.7500 1388.1000 138.9000 ;
	    RECT 1259.1000 137.2500 1388.1000 138.7500 ;
	    RECT 1259.1000 137.1000 1260.9000 137.2500 ;
	    RECT 1386.3000 137.1000 1388.1000 137.2500 ;
	    RECT 1465.5000 138.7500 1467.3000 138.9000 ;
	    RECT 1523.1000 138.7500 1524.9000 138.9000 ;
	    RECT 1465.5000 137.2500 1524.9000 138.7500 ;
	    RECT 1465.5000 137.1000 1467.3000 137.2500 ;
	    RECT 1523.1000 137.1000 1524.9000 137.2500 ;
	    RECT 493.5000 132.7500 495.3000 132.9000 ;
	    RECT 531.9000 132.7500 533.7000 132.9000 ;
	    RECT 493.5000 131.2500 533.7000 132.7500 ;
	    RECT 493.5000 131.1000 495.3000 131.2500 ;
	    RECT 531.9000 131.1000 533.7000 131.2500 ;
	    RECT 627.9000 132.7500 629.7000 132.9000 ;
	    RECT 771.9000 132.7500 773.7000 132.9000 ;
	    RECT 627.9000 131.2500 773.7000 132.7500 ;
	    RECT 627.9000 131.1000 629.7000 131.2500 ;
	    RECT 771.9000 131.1000 773.7000 131.2500 ;
	    RECT 990.3000 132.7500 992.1000 132.9000 ;
	    RECT 1052.7001 132.7500 1054.5000 132.9000 ;
	    RECT 990.3000 131.2500 1054.5000 132.7500 ;
	    RECT 990.3000 131.1000 992.1000 131.2500 ;
	    RECT 1052.7001 131.1000 1054.5000 131.2500 ;
	    RECT 1143.9000 132.7500 1145.7001 132.9000 ;
	    RECT 1153.5000 132.7500 1155.3000 132.9000 ;
	    RECT 1143.9000 131.2500 1155.3000 132.7500 ;
	    RECT 1143.9000 131.1000 1145.7001 131.2500 ;
	    RECT 1153.5000 131.1000 1155.3000 131.2500 ;
	    RECT 1208.7001 132.7500 1210.5000 132.9000 ;
	    RECT 1230.3000 132.7500 1232.1000 132.9000 ;
	    RECT 1208.7001 131.2500 1232.1000 132.7500 ;
	    RECT 1208.7001 131.1000 1210.5000 131.2500 ;
	    RECT 1230.3000 131.1000 1232.1000 131.2500 ;
	    RECT 1256.7001 132.7500 1258.5000 132.9000 ;
	    RECT 1297.5000 132.7500 1299.3000 132.9000 ;
	    RECT 1256.7001 131.2500 1299.3000 132.7500 ;
	    RECT 1256.7001 131.1000 1258.5000 131.2500 ;
	    RECT 1297.5000 131.1000 1299.3000 131.2500 ;
	    RECT 1309.5000 132.7500 1311.3000 132.9000 ;
	    RECT 1335.9000 132.7500 1337.7001 132.9000 ;
	    RECT 1309.5000 131.2500 1337.7001 132.7500 ;
	    RECT 1309.5000 131.1000 1311.3000 131.2500 ;
	    RECT 1335.9000 131.1000 1337.7001 131.2500 ;
	    RECT 1345.5000 132.7500 1347.3000 132.9000 ;
	    RECT 1391.1000 132.7500 1392.9000 132.9000 ;
	    RECT 1419.9000 132.7500 1421.7001 132.9000 ;
	    RECT 1345.5000 131.2500 1421.7001 132.7500 ;
	    RECT 1345.5000 131.1000 1347.3000 131.2500 ;
	    RECT 1391.1000 131.1000 1392.9000 131.2500 ;
	    RECT 1419.9000 131.1000 1421.7001 131.2500 ;
	    RECT 1460.7001 132.7500 1462.5000 132.9000 ;
	    RECT 1494.3000 132.7500 1496.1000 132.9000 ;
	    RECT 1460.7001 131.2500 1496.1000 132.7500 ;
	    RECT 1460.7001 131.1000 1462.5000 131.2500 ;
	    RECT 1494.3000 131.1000 1496.1000 131.2500 ;
	    RECT 229.5000 126.7500 231.3000 126.9000 ;
	    RECT 347.1000 126.7500 348.9000 126.9000 ;
	    RECT 229.5000 125.2500 348.9000 126.7500 ;
	    RECT 229.5000 125.1000 231.3000 125.2500 ;
	    RECT 347.1000 125.1000 348.9000 125.2500 ;
	    RECT 457.5000 126.7500 459.3000 126.9000 ;
	    RECT 469.5000 126.7500 471.3000 126.9000 ;
	    RECT 457.5000 125.2500 471.3000 126.7500 ;
	    RECT 457.5000 125.1000 459.3000 125.2500 ;
	    RECT 469.5000 125.1000 471.3000 125.2500 ;
	    RECT 486.3000 126.7500 488.1000 126.9000 ;
	    RECT 678.3000 126.7500 680.1000 126.9000 ;
	    RECT 486.3000 125.2500 680.1000 126.7500 ;
	    RECT 486.3000 125.1000 488.1000 125.2500 ;
	    RECT 678.3000 125.1000 680.1000 125.2500 ;
	    RECT 867.9000 126.7500 869.7000 126.9000 ;
	    RECT 954.3000 126.7500 956.1000 126.9000 ;
	    RECT 867.9000 125.2500 956.1000 126.7500 ;
	    RECT 867.9000 125.1000 869.7000 125.2500 ;
	    RECT 954.3000 125.1000 956.1000 125.2500 ;
	    RECT 973.5000 126.7500 975.3000 126.9000 ;
	    RECT 999.9000 126.7500 1001.7000 126.9000 ;
	    RECT 1009.5000 126.7500 1011.3000 126.9000 ;
	    RECT 973.5000 125.2500 1011.3000 126.7500 ;
	    RECT 973.5000 125.1000 975.3000 125.2500 ;
	    RECT 999.9000 125.1000 1001.7000 125.2500 ;
	    RECT 1009.5000 125.1000 1011.3000 125.2500 ;
	    RECT 1093.5000 126.7500 1095.3000 126.9000 ;
	    RECT 1247.1000 126.7500 1248.9000 126.9000 ;
	    RECT 1093.5000 125.2500 1248.9000 126.7500 ;
	    RECT 1093.5000 125.1000 1095.3000 125.2500 ;
	    RECT 1247.1000 125.1000 1248.9000 125.2500 ;
	    RECT 1304.7001 126.7500 1306.5000 126.9000 ;
	    RECT 1405.5000 126.7500 1407.3000 126.9000 ;
	    RECT 1304.7001 125.2500 1407.3000 126.7500 ;
	    RECT 1304.7001 125.1000 1306.5000 125.2500 ;
	    RECT 1405.5000 125.1000 1407.3000 125.2500 ;
	    RECT 287.1000 120.7500 288.9000 120.9000 ;
	    RECT 445.5000 120.7500 447.3000 120.9000 ;
	    RECT 287.1000 119.2500 447.3000 120.7500 ;
	    RECT 287.1000 119.1000 288.9000 119.2500 ;
	    RECT 445.5000 119.1000 447.3000 119.2500 ;
	    RECT 452.7000 120.7500 454.5000 120.9000 ;
	    RECT 488.7000 120.7500 490.5000 120.9000 ;
	    RECT 551.1000 120.7500 552.9000 120.9000 ;
	    RECT 452.7000 119.2500 552.9000 120.7500 ;
	    RECT 452.7000 119.1000 454.5000 119.2500 ;
	    RECT 488.7000 119.1000 490.5000 119.2500 ;
	    RECT 551.1000 119.1000 552.9000 119.2500 ;
	    RECT 791.1000 120.7500 792.9000 120.9000 ;
	    RECT 815.1000 120.7500 816.9000 120.9000 ;
	    RECT 791.1000 119.2500 816.9000 120.7500 ;
	    RECT 791.1000 119.1000 792.9000 119.2500 ;
	    RECT 815.1000 119.1000 816.9000 119.2500 ;
	    RECT 822.3000 120.7500 824.1000 120.9000 ;
	    RECT 959.1000 120.7500 960.9000 120.9000 ;
	    RECT 822.3000 119.2500 960.9000 120.7500 ;
	    RECT 822.3000 119.1000 824.1000 119.2500 ;
	    RECT 959.1000 119.1000 960.9000 119.2500 ;
	    RECT 980.7000 120.7500 982.5000 120.9000 ;
	    RECT 1081.5000 120.7500 1083.3000 120.9000 ;
	    RECT 980.7000 119.2500 1083.3000 120.7500 ;
	    RECT 980.7000 119.1000 982.5000 119.2500 ;
	    RECT 1081.5000 119.1000 1083.3000 119.2500 ;
	    RECT 1136.7001 120.7500 1138.5000 120.9000 ;
	    RECT 1167.9000 120.7500 1169.7001 120.9000 ;
	    RECT 1136.7001 119.2500 1169.7001 120.7500 ;
	    RECT 1136.7001 119.1000 1138.5000 119.2500 ;
	    RECT 1167.9000 119.1000 1169.7001 119.2500 ;
	    RECT 1175.1000 120.7500 1176.9000 120.9000 ;
	    RECT 1184.7001 120.7500 1186.5000 120.9000 ;
	    RECT 1175.1000 119.2500 1186.5000 120.7500 ;
	    RECT 1175.1000 119.1000 1176.9000 119.2500 ;
	    RECT 1184.7001 119.1000 1186.5000 119.2500 ;
	    RECT 1479.9000 120.7500 1481.7001 120.9000 ;
	    RECT 1484.7001 120.7500 1486.5000 120.9000 ;
	    RECT 1479.9000 119.2500 1486.5000 120.7500 ;
	    RECT 1479.9000 119.1000 1481.7001 119.2500 ;
	    RECT 1484.7001 119.1000 1486.5000 119.2500 ;
	    RECT 1506.3000 120.7500 1508.1000 120.9000 ;
	    RECT 1511.1000 120.7500 1512.9000 120.9000 ;
	    RECT 1547.1000 120.7500 1548.9000 120.9000 ;
	    RECT 1506.3000 119.2500 1548.9000 120.7500 ;
	    RECT 1506.3000 119.1000 1508.1000 119.2500 ;
	    RECT 1511.1000 119.1000 1512.9000 119.2500 ;
	    RECT 1547.1000 119.1000 1548.9000 119.2500 ;
	    RECT 13.5000 114.7500 15.3000 114.9000 ;
	    RECT 23.1000 114.7500 24.9000 114.9000 ;
	    RECT 13.5000 113.2500 24.9000 114.7500 ;
	    RECT 13.5000 113.1000 15.3000 113.2500 ;
	    RECT 23.1000 113.1000 24.9000 113.2500 ;
	    RECT 234.3000 114.7500 236.1000 114.9000 ;
	    RECT 243.9000 114.7500 245.7000 114.9000 ;
	    RECT 287.1000 114.7500 288.9000 114.9000 ;
	    RECT 234.3000 113.2500 288.9000 114.7500 ;
	    RECT 234.3000 113.1000 236.1000 113.2500 ;
	    RECT 243.9000 113.1000 245.7000 113.2500 ;
	    RECT 287.1000 113.1000 288.9000 113.2500 ;
	    RECT 347.1000 114.7500 348.9000 114.9000 ;
	    RECT 512.7000 114.7500 514.5000 114.9000 ;
	    RECT 347.1000 113.2500 514.5000 114.7500 ;
	    RECT 347.1000 113.1000 348.9000 113.2500 ;
	    RECT 512.7000 113.1000 514.5000 113.2500 ;
	    RECT 803.1000 114.7500 804.9000 114.9000 ;
	    RECT 851.1000 114.7500 852.9000 114.9000 ;
	    RECT 803.1000 113.2500 852.9000 114.7500 ;
	    RECT 803.1000 113.1000 804.9000 113.2500 ;
	    RECT 851.1000 113.1000 852.9000 113.2500 ;
	    RECT 935.1000 114.7500 936.9000 114.9000 ;
	    RECT 983.1000 114.7500 984.9000 114.9000 ;
	    RECT 935.1000 113.2500 984.9000 114.7500 ;
	    RECT 935.1000 113.1000 936.9000 113.2500 ;
	    RECT 983.1000 113.1000 984.9000 113.2500 ;
	    RECT 1148.7001 114.7500 1150.5000 114.9000 ;
	    RECT 1268.7001 114.7500 1270.5000 114.9000 ;
	    RECT 1148.7001 113.2500 1270.5000 114.7500 ;
	    RECT 1148.7001 113.1000 1150.5000 113.2500 ;
	    RECT 1268.7001 113.1000 1270.5000 113.2500 ;
	    RECT 1273.5000 114.7500 1275.3000 114.9000 ;
	    RECT 1309.5000 114.7500 1311.3000 114.9000 ;
	    RECT 1273.5000 113.2500 1311.3000 114.7500 ;
	    RECT 1273.5000 113.1000 1275.3000 113.2500 ;
	    RECT 1309.5000 113.1000 1311.3000 113.2500 ;
	    RECT 1328.7001 114.7500 1330.5000 114.9000 ;
	    RECT 1463.1000 114.7500 1464.9000 114.9000 ;
	    RECT 1328.7001 113.2500 1464.9000 114.7500 ;
	    RECT 1328.7001 113.1000 1330.5000 113.2500 ;
	    RECT 1463.1000 113.1000 1464.9000 113.2500 ;
	    RECT 380.7000 108.7500 382.5000 108.9000 ;
	    RECT 474.3000 108.7500 476.1000 108.9000 ;
	    RECT 380.7000 107.2500 476.1000 108.7500 ;
	    RECT 380.7000 107.1000 382.5000 107.2500 ;
	    RECT 474.3000 107.1000 476.1000 107.2500 ;
	    RECT 620.7000 108.7500 622.5000 108.9000 ;
	    RECT 721.5000 108.7500 723.3000 108.9000 ;
	    RECT 620.7000 107.2500 723.3000 108.7500 ;
	    RECT 620.7000 107.1000 622.5000 107.2500 ;
	    RECT 721.5000 107.1000 723.3000 107.2500 ;
	    RECT 944.7000 108.7500 946.5000 108.9000 ;
	    RECT 1011.9000 108.7500 1013.7000 108.9000 ;
	    RECT 944.7000 107.2500 1013.7000 108.7500 ;
	    RECT 944.7000 107.1000 946.5000 107.2500 ;
	    RECT 1011.9000 107.1000 1013.7000 107.2500 ;
	    RECT 1206.3000 108.7500 1208.1000 108.9000 ;
	    RECT 1256.7001 108.7500 1258.5000 108.9000 ;
	    RECT 1206.3000 107.2500 1258.5000 108.7500 ;
	    RECT 1206.3000 107.1000 1208.1000 107.2500 ;
	    RECT 1256.7001 107.1000 1258.5000 107.2500 ;
	    RECT 1266.3000 108.7500 1268.1000 108.9000 ;
	    RECT 1383.9000 108.7500 1385.7001 108.9000 ;
	    RECT 1266.3000 107.2500 1385.7001 108.7500 ;
	    RECT 1266.3000 107.1000 1268.1000 107.2500 ;
	    RECT 1383.9000 107.1000 1385.7001 107.2500 ;
	    RECT 1463.1000 108.7500 1464.9000 108.9000 ;
	    RECT 1499.1000 108.7500 1500.9000 108.9000 ;
	    RECT 1463.1000 107.2500 1500.9000 108.7500 ;
	    RECT 1463.1000 107.1000 1464.9000 107.2500 ;
	    RECT 1499.1000 107.1000 1500.9000 107.2500 ;
	    RECT 18.3000 102.7500 20.1000 102.9000 ;
	    RECT 54.3000 102.7500 56.1000 102.9000 ;
	    RECT 18.3000 101.2500 56.1000 102.7500 ;
	    RECT 18.3000 101.1000 20.1000 101.2500 ;
	    RECT 54.3000 101.1000 56.1000 101.2500 ;
	    RECT 234.3000 102.7500 236.1000 102.9000 ;
	    RECT 246.3000 102.7500 248.1000 102.9000 ;
	    RECT 234.3000 101.2500 248.1000 102.7500 ;
	    RECT 234.3000 101.1000 236.1000 101.2500 ;
	    RECT 246.3000 101.1000 248.1000 101.2500 ;
	    RECT 277.5000 102.7500 279.3000 102.9000 ;
	    RECT 318.3000 102.7500 320.1000 102.9000 ;
	    RECT 277.5000 101.2500 320.1000 102.7500 ;
	    RECT 277.5000 101.1000 279.3000 101.2500 ;
	    RECT 318.3000 101.1000 320.1000 101.2500 ;
	    RECT 421.5000 102.7500 423.3000 102.9000 ;
	    RECT 483.9000 102.7500 485.7000 102.9000 ;
	    RECT 421.5000 101.2500 485.7000 102.7500 ;
	    RECT 421.5000 101.1000 423.3000 101.2500 ;
	    RECT 483.9000 101.1000 485.7000 101.2500 ;
	    RECT 769.5000 102.7500 771.3000 102.9000 ;
	    RECT 779.1000 102.7500 780.9000 102.9000 ;
	    RECT 798.3000 102.7500 800.1000 102.9000 ;
	    RECT 769.5000 101.2500 800.1000 102.7500 ;
	    RECT 769.5000 101.1000 771.3000 101.2500 ;
	    RECT 779.1000 101.1000 780.9000 101.2500 ;
	    RECT 798.3000 101.1000 800.1000 101.2500 ;
	    RECT 1165.5000 102.7500 1167.3000 102.9000 ;
	    RECT 1235.1000 102.7500 1236.9000 102.9000 ;
	    RECT 1165.5000 101.2500 1236.9000 102.7500 ;
	    RECT 1165.5000 101.1000 1167.3000 101.2500 ;
	    RECT 1235.1000 101.1000 1236.9000 101.2500 ;
	    RECT 1266.3000 102.7500 1268.1000 102.9000 ;
	    RECT 1273.5000 102.7500 1275.3000 102.9000 ;
	    RECT 1266.3000 101.2500 1275.3000 102.7500 ;
	    RECT 1266.3000 101.1000 1268.1000 101.2500 ;
	    RECT 1273.5000 101.1000 1275.3000 101.2500 ;
	    RECT 1285.5000 102.7500 1287.3000 102.9000 ;
	    RECT 1321.5000 102.7500 1323.3000 102.9000 ;
	    RECT 1369.5000 102.7500 1371.3000 102.9000 ;
	    RECT 1415.1000 102.7500 1416.9000 102.9000 ;
	    RECT 1285.5000 101.2500 1416.9000 102.7500 ;
	    RECT 1285.5000 101.1000 1287.3000 101.2500 ;
	    RECT 1321.5000 101.1000 1323.3000 101.2500 ;
	    RECT 1369.5000 101.1000 1371.3000 101.2500 ;
	    RECT 1415.1000 101.1000 1416.9000 101.2500 ;
	    RECT 1494.3000 102.7500 1496.1000 102.9000 ;
	    RECT 1520.7001 102.7500 1522.5000 102.9000 ;
	    RECT 1494.3000 101.2500 1522.5000 102.7500 ;
	    RECT 1494.3000 101.1000 1496.1000 101.2500 ;
	    RECT 1520.7001 101.1000 1522.5000 101.2500 ;
	    RECT 337.5000 96.7500 339.3000 96.9000 ;
	    RECT 356.7000 96.7500 358.5000 96.9000 ;
	    RECT 337.5000 95.2500 358.5000 96.7500 ;
	    RECT 337.5000 95.1000 339.3000 95.2500 ;
	    RECT 356.7000 95.1000 358.5000 95.2500 ;
	    RECT 594.3000 96.7500 596.1000 96.9000 ;
	    RECT 687.9000 96.7500 689.7000 96.9000 ;
	    RECT 594.3000 95.2500 689.7000 96.7500 ;
	    RECT 594.3000 95.1000 596.1000 95.2500 ;
	    RECT 687.9000 95.1000 689.7000 95.2500 ;
	    RECT 1052.7001 96.7500 1054.5000 96.9000 ;
	    RECT 1201.5000 96.7500 1203.3000 96.9000 ;
	    RECT 1239.9000 96.7500 1241.7001 96.9000 ;
	    RECT 1271.1000 96.7500 1272.9000 96.9000 ;
	    RECT 1052.7001 95.2500 1272.9000 96.7500 ;
	    RECT 1052.7001 95.1000 1054.5000 95.2500 ;
	    RECT 1201.5000 95.1000 1203.3000 95.2500 ;
	    RECT 1239.9000 95.1000 1241.7001 95.2500 ;
	    RECT 1271.1000 95.1000 1272.9000 95.2500 ;
	    RECT 1275.9000 96.7500 1277.7001 96.9000 ;
	    RECT 1307.1000 96.7500 1308.9000 96.9000 ;
	    RECT 1275.9000 95.2500 1308.9000 96.7500 ;
	    RECT 1275.9000 95.1000 1277.7001 95.2500 ;
	    RECT 1307.1000 95.1000 1308.9000 95.2500 ;
	    RECT 1482.3000 96.7500 1484.1000 96.9000 ;
	    RECT 1494.3000 96.7500 1496.1000 96.9000 ;
	    RECT 1482.3000 95.2500 1496.1000 96.7500 ;
	    RECT 1482.3000 95.1000 1484.1000 95.2500 ;
	    RECT 1494.3000 95.1000 1496.1000 95.2500 ;
	    RECT 311.1000 90.7500 312.9000 90.9000 ;
	    RECT 339.9000 90.7500 341.7000 90.9000 ;
	    RECT 311.1000 89.2500 341.7000 90.7500 ;
	    RECT 311.1000 89.1000 312.9000 89.2500 ;
	    RECT 339.9000 89.1000 341.7000 89.2500 ;
	    RECT 349.5000 90.7500 351.3000 90.9000 ;
	    RECT 363.9000 90.7500 365.7000 90.9000 ;
	    RECT 349.5000 89.2500 365.7000 90.7500 ;
	    RECT 349.5000 89.1000 351.3000 89.2500 ;
	    RECT 363.9000 89.1000 365.7000 89.2500 ;
	    RECT 731.1000 90.7500 732.9000 90.9000 ;
	    RECT 781.5000 90.7500 783.3000 90.9000 ;
	    RECT 731.1000 89.2500 783.3000 90.7500 ;
	    RECT 731.1000 89.1000 732.9000 89.2500 ;
	    RECT 781.5000 89.1000 783.3000 89.2500 ;
	    RECT 1177.5000 90.7500 1179.3000 90.9000 ;
	    RECT 1335.9000 90.7500 1337.7001 90.9000 ;
	    RECT 1177.5000 89.2500 1337.7001 90.7500 ;
	    RECT 1177.5000 89.1000 1179.3000 89.2500 ;
	    RECT 1335.9000 89.1000 1337.7001 89.2500 ;
	    RECT 1400.7001 90.7500 1402.5000 90.9000 ;
	    RECT 1453.5000 90.7500 1455.3000 90.9000 ;
	    RECT 1400.7001 89.2500 1455.3000 90.7500 ;
	    RECT 1400.7001 89.1000 1402.5000 89.2500 ;
	    RECT 1453.5000 89.1000 1455.3000 89.2500 ;
	    RECT 1458.3000 90.7500 1460.1000 90.9000 ;
	    RECT 1499.1000 90.7500 1500.9000 90.9000 ;
	    RECT 1458.3000 89.2500 1500.9000 90.7500 ;
	    RECT 1458.3000 89.1000 1460.1000 89.2500 ;
	    RECT 1499.1000 89.1000 1500.9000 89.2500 ;
	    RECT 47.1000 84.7500 48.9000 84.9000 ;
	    RECT 143.1000 84.7500 144.9000 84.9000 ;
	    RECT 47.1000 83.2500 144.9000 84.7500 ;
	    RECT 47.1000 83.1000 48.9000 83.2500 ;
	    RECT 143.1000 83.1000 144.9000 83.2500 ;
	    RECT 596.7000 84.7500 598.5000 84.9000 ;
	    RECT 625.5000 84.7500 627.3000 84.9000 ;
	    RECT 596.7000 83.2500 627.3000 84.7500 ;
	    RECT 596.7000 83.1000 598.5000 83.2500 ;
	    RECT 625.5000 83.1000 627.3000 83.2500 ;
	    RECT 721.5000 84.7500 723.3000 84.9000 ;
	    RECT 750.3000 84.7500 752.1000 84.9000 ;
	    RECT 721.5000 83.2500 752.1000 84.7500 ;
	    RECT 721.5000 83.1000 723.3000 83.2500 ;
	    RECT 750.3000 83.1000 752.1000 83.2500 ;
	    RECT 1175.1000 84.7500 1176.9000 84.9000 ;
	    RECT 1184.7001 84.7500 1186.5000 84.9000 ;
	    RECT 1175.1000 83.2500 1186.5000 84.7500 ;
	    RECT 1175.1000 83.1000 1176.9000 83.2500 ;
	    RECT 1184.7001 83.1000 1186.5000 83.2500 ;
	    RECT 1239.9000 84.7500 1241.7001 84.9000 ;
	    RECT 1283.1000 84.7500 1284.9000 84.9000 ;
	    RECT 1239.9000 83.2500 1284.9000 84.7500 ;
	    RECT 1239.9000 83.1000 1241.7001 83.2500 ;
	    RECT 1283.1000 83.1000 1284.9000 83.2500 ;
	    RECT 1427.1000 84.7500 1428.9000 84.9000 ;
	    RECT 1434.3000 84.7500 1436.1000 84.9000 ;
	    RECT 1427.1000 83.2500 1436.1000 84.7500 ;
	    RECT 1427.1000 83.1000 1428.9000 83.2500 ;
	    RECT 1434.3000 83.1000 1436.1000 83.2500 ;
	    RECT 1465.5000 84.7500 1467.3000 84.9000 ;
	    RECT 1489.5000 84.7500 1491.3000 84.9000 ;
	    RECT 1465.5000 83.2500 1491.3000 84.7500 ;
	    RECT 1465.5000 83.1000 1467.3000 83.2500 ;
	    RECT 1489.5000 83.1000 1491.3000 83.2500 ;
	    RECT 1494.3000 84.7500 1496.1000 84.9000 ;
	    RECT 1549.5000 84.7500 1551.3000 84.9000 ;
	    RECT 1494.3000 83.2500 1551.3000 84.7500 ;
	    RECT 1494.3000 83.1000 1496.1000 83.2500 ;
	    RECT 1549.5000 83.1000 1551.3000 83.2500 ;
	    RECT 133.5000 78.7500 135.3000 78.9000 ;
	    RECT 243.9000 78.7500 245.7000 78.9000 ;
	    RECT 133.5000 77.2500 245.7000 78.7500 ;
	    RECT 133.5000 77.1000 135.3000 77.2500 ;
	    RECT 243.9000 77.1000 245.7000 77.2500 ;
	    RECT 491.1000 78.7500 492.9000 78.9000 ;
	    RECT 522.3000 78.7500 524.1000 78.9000 ;
	    RECT 491.1000 77.2500 524.1000 78.7500 ;
	    RECT 491.1000 77.1000 492.9000 77.2500 ;
	    RECT 522.3000 77.1000 524.1000 77.2500 ;
	    RECT 728.7000 78.7500 730.5000 78.9000 ;
	    RECT 740.7000 78.7500 742.5000 78.9000 ;
	    RECT 728.7000 77.2500 742.5000 78.7500 ;
	    RECT 728.7000 77.1000 730.5000 77.2500 ;
	    RECT 740.7000 77.1000 742.5000 77.2500 ;
	    RECT 1167.9000 78.7500 1169.7001 78.9000 ;
	    RECT 1371.9000 78.7500 1373.7001 78.9000 ;
	    RECT 1167.9000 77.2500 1373.7001 78.7500 ;
	    RECT 1167.9000 77.1000 1169.7001 77.2500 ;
	    RECT 1371.9000 77.1000 1373.7001 77.2500 ;
	    RECT 1427.1000 78.7500 1428.9000 78.9000 ;
	    RECT 1443.9000 78.7500 1445.7001 78.9000 ;
	    RECT 1427.1000 77.2500 1445.7001 78.7500 ;
	    RECT 1427.1000 77.1000 1428.9000 77.2500 ;
	    RECT 1443.9000 77.1000 1445.7001 77.2500 ;
	    RECT 1491.9000 78.7500 1493.7001 78.9000 ;
	    RECT 1511.1000 78.7500 1512.9000 78.9000 ;
	    RECT 1491.9000 77.2500 1512.9000 78.7500 ;
	    RECT 1491.9000 77.1000 1493.7001 77.2500 ;
	    RECT 1511.1000 77.1000 1512.9000 77.2500 ;
	    RECT 311.1000 72.7500 312.9000 72.9000 ;
	    RECT 320.7000 72.7500 322.5000 72.9000 ;
	    RECT 311.1000 71.2500 322.5000 72.7500 ;
	    RECT 311.1000 71.1000 312.9000 71.2500 ;
	    RECT 320.7000 71.1000 322.5000 71.2500 ;
	    RECT 534.3000 72.7500 536.1000 72.9000 ;
	    RECT 723.9000 72.7500 725.7000 72.9000 ;
	    RECT 534.3000 71.2500 725.7000 72.7500 ;
	    RECT 534.3000 71.1000 536.1000 71.2500 ;
	    RECT 723.9000 71.1000 725.7000 71.2500 ;
	    RECT 1047.9000 72.7500 1049.7001 72.9000 ;
	    RECT 1153.5000 72.7500 1155.3000 72.9000 ;
	    RECT 1235.1000 72.7500 1236.9000 72.9000 ;
	    RECT 1047.9000 71.2500 1236.9000 72.7500 ;
	    RECT 1047.9000 71.1000 1049.7001 71.2500 ;
	    RECT 1153.5000 71.1000 1155.3000 71.2500 ;
	    RECT 1235.1000 71.1000 1236.9000 71.2500 ;
	    RECT 1244.7001 72.7500 1246.5000 72.9000 ;
	    RECT 1455.9000 72.7500 1457.7001 72.9000 ;
	    RECT 1467.9000 72.7500 1469.7001 72.9000 ;
	    RECT 1487.1000 72.7500 1488.9000 72.9000 ;
	    RECT 1244.7001 71.2500 1488.9000 72.7500 ;
	    RECT 1244.7001 71.1000 1246.5000 71.2500 ;
	    RECT 1455.9000 71.1000 1457.7001 71.2500 ;
	    RECT 1467.9000 71.1000 1469.7001 71.2500 ;
	    RECT 1487.1000 71.1000 1488.9000 71.2500 ;
	    RECT 1496.7001 72.7500 1498.5000 72.9000 ;
	    RECT 1518.3000 72.7500 1520.1000 72.9000 ;
	    RECT 1496.7001 71.2500 1520.1000 72.7500 ;
	    RECT 1496.7001 71.1000 1498.5000 71.2500 ;
	    RECT 1518.3000 71.1000 1520.1000 71.2500 ;
	    RECT 1523.1000 72.7500 1524.9000 72.9000 ;
	    RECT 1547.1000 72.7500 1548.9000 72.9000 ;
	    RECT 1523.1000 71.2500 1548.9000 72.7500 ;
	    RECT 1523.1000 71.1000 1524.9000 71.2500 ;
	    RECT 1547.1000 71.1000 1548.9000 71.2500 ;
	    RECT 536.7000 66.7500 538.5000 66.9000 ;
	    RECT 558.3000 66.7500 560.1000 66.9000 ;
	    RECT 565.5000 66.7500 567.3000 66.9000 ;
	    RECT 536.7000 65.2500 567.3000 66.7500 ;
	    RECT 536.7000 65.1000 538.5000 65.2500 ;
	    RECT 558.3000 65.1000 560.1000 65.2500 ;
	    RECT 565.5000 65.1000 567.3000 65.2500 ;
	    RECT 723.9000 66.7500 725.7000 66.9000 ;
	    RECT 973.5000 66.7500 975.3000 66.9000 ;
	    RECT 723.9000 65.2500 975.3000 66.7500 ;
	    RECT 723.9000 65.1000 725.7000 65.2500 ;
	    RECT 973.5000 65.1000 975.3000 65.2500 ;
	    RECT 1098.3000 66.7500 1100.1000 66.9000 ;
	    RECT 1155.9000 66.7500 1157.7001 66.9000 ;
	    RECT 1098.3000 65.2500 1157.7001 66.7500 ;
	    RECT 1098.3000 65.1000 1100.1000 65.2500 ;
	    RECT 1155.9000 65.1000 1157.7001 65.2500 ;
	    RECT 1170.3000 66.7500 1172.1000 66.9000 ;
	    RECT 1177.5000 66.7500 1179.3000 66.9000 ;
	    RECT 1170.3000 65.2500 1179.3000 66.7500 ;
	    RECT 1170.3000 65.1000 1172.1000 65.2500 ;
	    RECT 1177.5000 65.1000 1179.3000 65.2500 ;
	    RECT 1398.3000 66.7500 1400.1000 66.9000 ;
	    RECT 1434.3000 66.7500 1436.1000 66.9000 ;
	    RECT 1513.5000 66.7500 1515.3000 66.9000 ;
	    RECT 1398.3000 65.2500 1515.3000 66.7500 ;
	    RECT 1398.3000 65.1000 1400.1000 65.2500 ;
	    RECT 1434.3000 65.1000 1436.1000 65.2500 ;
	    RECT 1513.5000 65.1000 1515.3000 65.2500 ;
	    RECT 1525.5000 66.7500 1527.3000 66.9000 ;
	    RECT 1554.3000 66.7500 1556.1000 66.9000 ;
	    RECT 1525.5000 65.2500 1556.1000 66.7500 ;
	    RECT 1525.5000 65.1000 1527.3000 65.2500 ;
	    RECT 1554.3000 65.1000 1556.1000 65.2500 ;
	    RECT 335.1000 60.7500 336.9000 60.9000 ;
	    RECT 349.5000 60.7500 351.3000 60.9000 ;
	    RECT 368.7000 60.7500 370.5000 60.9000 ;
	    RECT 335.1000 59.2500 370.5000 60.7500 ;
	    RECT 335.1000 59.1000 336.9000 59.2500 ;
	    RECT 349.5000 59.1000 351.3000 59.2500 ;
	    RECT 368.7000 59.1000 370.5000 59.2500 ;
	    RECT 493.5000 60.7500 495.3000 60.9000 ;
	    RECT 543.9000 60.7500 545.7000 60.9000 ;
	    RECT 493.5000 59.2500 545.7000 60.7500 ;
	    RECT 493.5000 59.1000 495.3000 59.2500 ;
	    RECT 543.9000 59.1000 545.7000 59.2500 ;
	    RECT 690.3000 60.7500 692.1000 60.9000 ;
	    RECT 855.9000 60.7500 857.7000 60.9000 ;
	    RECT 690.3000 59.2500 857.7000 60.7500 ;
	    RECT 690.3000 59.1000 692.1000 59.2500 ;
	    RECT 855.9000 59.1000 857.7000 59.2500 ;
	    RECT 1172.7001 60.7500 1174.5000 60.9000 ;
	    RECT 1179.9000 60.7500 1181.7001 60.9000 ;
	    RECT 1172.7001 59.2500 1181.7001 60.7500 ;
	    RECT 1172.7001 59.1000 1174.5000 59.2500 ;
	    RECT 1179.9000 59.1000 1181.7001 59.2500 ;
	    RECT 1215.9000 60.7500 1217.7001 60.9000 ;
	    RECT 1343.1000 60.7500 1344.9000 60.9000 ;
	    RECT 1395.9000 60.7500 1397.7001 60.9000 ;
	    RECT 1215.9000 59.2500 1397.7001 60.7500 ;
	    RECT 1215.9000 59.1000 1217.7001 59.2500 ;
	    RECT 1343.1000 59.1000 1344.9000 59.2500 ;
	    RECT 1395.9000 59.1000 1397.7001 59.2500 ;
	    RECT 1458.3000 60.7500 1460.1000 60.9000 ;
	    RECT 1515.9000 60.7500 1517.7001 60.9000 ;
	    RECT 1458.3000 59.2500 1517.7001 60.7500 ;
	    RECT 1458.3000 59.1000 1460.1000 59.2500 ;
	    RECT 1515.9000 59.1000 1517.7001 59.2500 ;
	    RECT 308.7000 54.7500 310.5000 54.9000 ;
	    RECT 337.5000 54.7500 339.3000 54.9000 ;
	    RECT 308.7000 53.2500 339.3000 54.7500 ;
	    RECT 308.7000 53.1000 310.5000 53.2500 ;
	    RECT 337.5000 53.1000 339.3000 53.2500 ;
	    RECT 519.9000 54.7500 521.7000 54.9000 ;
	    RECT 539.1000 54.7500 540.9000 54.9000 ;
	    RECT 519.9000 53.2500 540.9000 54.7500 ;
	    RECT 519.9000 53.1000 521.7000 53.2500 ;
	    RECT 539.1000 53.1000 540.9000 53.2500 ;
	    RECT 625.5000 54.7500 627.3000 54.9000 ;
	    RECT 731.1000 54.7500 732.9000 54.9000 ;
	    RECT 625.5000 53.2500 732.9000 54.7500 ;
	    RECT 625.5000 53.1000 627.3000 53.2500 ;
	    RECT 731.1000 53.1000 732.9000 53.2500 ;
	    RECT 963.9000 54.7500 965.7000 54.9000 ;
	    RECT 1055.1000 54.7500 1056.9000 54.9000 ;
	    RECT 963.9000 53.2500 1056.9000 54.7500 ;
	    RECT 963.9000 53.1000 965.7000 53.2500 ;
	    RECT 1055.1000 53.1000 1056.9000 53.2500 ;
	    RECT 1172.7001 54.7500 1174.5000 54.9000 ;
	    RECT 1297.5000 54.7500 1299.3000 54.9000 ;
	    RECT 1302.3000 54.7500 1304.1000 54.9000 ;
	    RECT 1172.7001 53.2500 1304.1000 54.7500 ;
	    RECT 1172.7001 53.1000 1174.5000 53.2500 ;
	    RECT 1297.5000 53.1000 1299.3000 53.2500 ;
	    RECT 1302.3000 53.1000 1304.1000 53.2500 ;
	    RECT 1491.9000 54.7500 1493.7001 54.9000 ;
	    RECT 1496.7001 54.7500 1498.5000 54.9000 ;
	    RECT 1491.9000 53.2500 1498.5000 54.7500 ;
	    RECT 1491.9000 53.1000 1493.7001 53.2500 ;
	    RECT 1496.7001 53.1000 1498.5000 53.2500 ;
	    RECT 1511.1000 54.7500 1512.9000 54.9000 ;
	    RECT 1523.1000 54.7500 1524.9000 54.9000 ;
	    RECT 1511.1000 53.2500 1524.9000 54.7500 ;
	    RECT 1511.1000 53.1000 1512.9000 53.2500 ;
	    RECT 1523.1000 53.1000 1524.9000 53.2500 ;
	    RECT 164.7000 48.7500 166.5000 48.9000 ;
	    RECT 181.5000 48.7500 183.3000 48.9000 ;
	    RECT 164.7000 47.2500 183.3000 48.7500 ;
	    RECT 164.7000 47.1000 166.5000 47.2500 ;
	    RECT 181.5000 47.1000 183.3000 47.2500 ;
	    RECT 282.3000 48.7500 284.1000 48.9000 ;
	    RECT 347.1000 48.7500 348.9000 48.9000 ;
	    RECT 282.3000 47.2500 348.9000 48.7500 ;
	    RECT 282.3000 47.1000 284.1000 47.2500 ;
	    RECT 347.1000 47.1000 348.9000 47.2500 ;
	    RECT 493.5000 48.7500 495.3000 48.9000 ;
	    RECT 500.7000 48.7500 502.5000 48.9000 ;
	    RECT 493.5000 47.2500 502.5000 48.7500 ;
	    RECT 493.5000 47.1000 495.3000 47.2500 ;
	    RECT 500.7000 47.1000 502.5000 47.2500 ;
	    RECT 702.3000 48.7500 704.1000 48.9000 ;
	    RECT 769.5000 48.7500 771.3000 48.9000 ;
	    RECT 702.3000 47.2500 771.3000 48.7500 ;
	    RECT 702.3000 47.1000 704.1000 47.2500 ;
	    RECT 769.5000 47.1000 771.3000 47.2500 ;
	    RECT 1086.3000 48.7500 1088.1000 48.9000 ;
	    RECT 1170.3000 48.7500 1172.1000 48.9000 ;
	    RECT 1086.3000 47.2500 1172.1000 48.7500 ;
	    RECT 1086.3000 47.1000 1088.1000 47.2500 ;
	    RECT 1170.3000 47.1000 1172.1000 47.2500 ;
	    RECT 1175.1000 48.7500 1176.9000 48.9000 ;
	    RECT 1182.3000 48.7500 1184.1000 48.9000 ;
	    RECT 1175.1000 47.2500 1184.1000 48.7500 ;
	    RECT 1175.1000 47.1000 1176.9000 47.2500 ;
	    RECT 1182.3000 47.1000 1184.1000 47.2500 ;
	    RECT 1235.1000 48.7500 1236.9000 48.9000 ;
	    RECT 1369.5000 48.7500 1371.3000 48.9000 ;
	    RECT 1235.1000 47.2500 1371.3000 48.7500 ;
	    RECT 1235.1000 47.1000 1236.9000 47.2500 ;
	    RECT 1369.5000 47.1000 1371.3000 47.2500 ;
	    RECT 1484.7001 48.7500 1486.5000 48.9000 ;
	    RECT 1489.5000 48.7500 1491.3000 48.9000 ;
	    RECT 1484.7001 47.2500 1491.3000 48.7500 ;
	    RECT 1484.7001 47.1000 1486.5000 47.2500 ;
	    RECT 1489.5000 47.1000 1491.3000 47.2500 ;
	    RECT 1520.7001 48.7500 1522.5000 48.9000 ;
	    RECT 1554.3000 48.7500 1556.1000 48.9000 ;
	    RECT 1520.7001 47.2500 1556.1000 48.7500 ;
	    RECT 1520.7001 47.1000 1522.5000 47.2500 ;
	    RECT 1554.3000 47.1000 1556.1000 47.2500 ;
	    RECT 126.3000 42.7500 128.1000 42.9000 ;
	    RECT 155.1000 42.7500 156.9000 42.9000 ;
	    RECT 126.3000 41.2500 156.9000 42.7500 ;
	    RECT 126.3000 41.1000 128.1000 41.2500 ;
	    RECT 155.1000 41.1000 156.9000 41.2500 ;
	    RECT 229.5000 42.7500 231.3000 42.9000 ;
	    RECT 332.7000 42.7500 334.5000 42.9000 ;
	    RECT 229.5000 41.2500 334.5000 42.7500 ;
	    RECT 229.5000 41.1000 231.3000 41.2500 ;
	    RECT 332.7000 41.1000 334.5000 41.2500 ;
	    RECT 498.3000 42.7500 500.1000 42.9000 ;
	    RECT 524.7000 42.7500 526.5000 42.9000 ;
	    RECT 498.3000 41.2500 526.5000 42.7500 ;
	    RECT 498.3000 41.1000 500.1000 41.2500 ;
	    RECT 524.7000 41.1000 526.5000 41.2500 ;
	    RECT 711.9000 42.7500 713.7000 42.9000 ;
	    RECT 723.9000 42.7500 725.7000 42.9000 ;
	    RECT 711.9000 41.2500 725.7000 42.7500 ;
	    RECT 711.9000 41.1000 713.7000 41.2500 ;
	    RECT 723.9000 41.1000 725.7000 41.2500 ;
	    RECT 947.1000 42.7500 948.9000 42.9000 ;
	    RECT 959.1000 42.7500 960.9000 42.9000 ;
	    RECT 947.1000 41.2500 960.9000 42.7500 ;
	    RECT 947.1000 41.1000 948.9000 41.2500 ;
	    RECT 959.1000 41.1000 960.9000 41.2500 ;
	    RECT 1050.3000 42.7500 1052.1000 42.9000 ;
	    RECT 1069.5000 42.7500 1071.3000 42.9000 ;
	    RECT 1050.3000 41.2500 1071.3000 42.7500 ;
	    RECT 1050.3000 41.1000 1052.1000 41.2500 ;
	    RECT 1069.5000 41.1000 1071.3000 41.2500 ;
	    RECT 1172.7001 42.7500 1174.5000 42.9000 ;
	    RECT 1206.3000 42.7500 1208.1000 42.9000 ;
	    RECT 1172.7001 41.2500 1208.1000 42.7500 ;
	    RECT 1172.7001 41.1000 1174.5000 41.2500 ;
	    RECT 1206.3000 41.1000 1208.1000 41.2500 ;
	    RECT 1237.5000 42.7500 1239.3000 42.9000 ;
	    RECT 1251.9000 42.7500 1253.7001 42.9000 ;
	    RECT 1237.5000 41.2500 1253.7001 42.7500 ;
	    RECT 1237.5000 41.1000 1239.3000 41.2500 ;
	    RECT 1251.9000 41.1000 1253.7001 41.2500 ;
	    RECT 1362.3000 42.7500 1364.1000 42.9000 ;
	    RECT 1405.5000 42.7500 1407.3000 42.9000 ;
	    RECT 1362.3000 41.2500 1407.3000 42.7500 ;
	    RECT 1362.3000 41.1000 1364.1000 41.2500 ;
	    RECT 1405.5000 41.1000 1407.3000 41.2500 ;
	    RECT 306.3000 36.7500 308.1000 36.9000 ;
	    RECT 337.5000 36.7500 339.3000 36.9000 ;
	    RECT 306.3000 35.2500 339.3000 36.7500 ;
	    RECT 306.3000 35.1000 308.1000 35.2500 ;
	    RECT 337.5000 35.1000 339.3000 35.2500 ;
	    RECT 469.5000 36.7500 471.3000 36.9000 ;
	    RECT 541.5000 36.7500 543.3000 36.9000 ;
	    RECT 469.5000 35.2500 543.3000 36.7500 ;
	    RECT 469.5000 35.1000 471.3000 35.2500 ;
	    RECT 541.5000 35.1000 543.3000 35.2500 ;
	    RECT 697.5000 36.7500 699.3000 36.9000 ;
	    RECT 755.1000 36.7500 756.9000 36.9000 ;
	    RECT 697.5000 35.2500 756.9000 36.7500 ;
	    RECT 697.5000 35.1000 699.3000 35.2500 ;
	    RECT 755.1000 35.1000 756.9000 35.2500 ;
	    RECT 1340.7001 36.7500 1342.5000 36.9000 ;
	    RECT 1374.3000 36.7500 1376.1000 36.9000 ;
	    RECT 1410.3000 36.7500 1412.1000 36.9000 ;
	    RECT 1340.7001 35.2500 1412.1000 36.7500 ;
	    RECT 1340.7001 35.1000 1342.5000 35.2500 ;
	    RECT 1374.3000 35.1000 1376.1000 35.2500 ;
	    RECT 1410.3000 35.1000 1412.1000 35.2500 ;
	    RECT 1470.3000 36.7500 1472.1000 36.9000 ;
	    RECT 1508.7001 36.7500 1510.5000 36.9000 ;
	    RECT 1470.3000 35.2500 1510.5000 36.7500 ;
	    RECT 1470.3000 35.1000 1472.1000 35.2500 ;
	    RECT 1508.7001 35.1000 1510.5000 35.2500 ;
	    RECT 347.1000 30.7500 348.9000 30.9000 ;
	    RECT 356.7000 30.7500 358.5000 30.9000 ;
	    RECT 347.1000 29.2500 358.5000 30.7500 ;
	    RECT 347.1000 29.1000 348.9000 29.2500 ;
	    RECT 356.7000 29.1000 358.5000 29.2500 ;
	    RECT 488.7000 30.7500 490.5000 30.9000 ;
	    RECT 515.1000 30.7500 516.9000 30.9000 ;
	    RECT 488.7000 29.2500 516.9000 30.7500 ;
	    RECT 488.7000 29.1000 490.5000 29.2500 ;
	    RECT 515.1000 29.1000 516.9000 29.2500 ;
	    RECT 563.1000 30.7500 564.9000 30.9000 ;
	    RECT 584.7000 30.7500 586.5000 30.9000 ;
	    RECT 563.1000 29.2500 586.5000 30.7500 ;
	    RECT 563.1000 29.1000 564.9000 29.2500 ;
	    RECT 584.7000 29.1000 586.5000 29.2500 ;
	    RECT 726.3000 30.7500 728.1000 30.9000 ;
	    RECT 764.7000 30.7500 766.5000 30.9000 ;
	    RECT 726.3000 29.2500 766.5000 30.7500 ;
	    RECT 726.3000 29.1000 728.1000 29.2500 ;
	    RECT 764.7000 29.1000 766.5000 29.2500 ;
	    RECT 774.3000 30.7500 776.1000 30.9000 ;
	    RECT 800.7000 30.7500 802.5000 30.9000 ;
	    RECT 774.3000 29.2500 802.5000 30.7500 ;
	    RECT 774.3000 29.1000 776.1000 29.2500 ;
	    RECT 800.7000 29.1000 802.5000 29.2500 ;
	    RECT 959.1000 30.7500 960.9000 30.9000 ;
	    RECT 1047.9000 30.7500 1049.7001 30.9000 ;
	    RECT 959.1000 29.2500 1049.7001 30.7500 ;
	    RECT 959.1000 29.1000 960.9000 29.2500 ;
	    RECT 1047.9000 29.1000 1049.7001 29.2500 ;
	    RECT 1074.3000 30.7500 1076.1000 30.9000 ;
	    RECT 1230.3000 30.7500 1232.1000 30.9000 ;
	    RECT 1340.7001 30.7500 1342.5000 30.9000 ;
	    RECT 1074.3000 29.2500 1342.5000 30.7500 ;
	    RECT 1074.3000 29.1000 1076.1000 29.2500 ;
	    RECT 1230.3000 29.1000 1232.1000 29.2500 ;
	    RECT 1340.7001 29.1000 1342.5000 29.2500 ;
	    RECT 1369.5000 30.7500 1371.3000 30.9000 ;
	    RECT 1484.7001 30.7500 1486.5000 30.9000 ;
	    RECT 1369.5000 29.2500 1486.5000 30.7500 ;
	    RECT 1369.5000 29.1000 1371.3000 29.2500 ;
	    RECT 1484.7001 29.1000 1486.5000 29.2500 ;
	    RECT 49.5000 24.7500 51.3000 24.9000 ;
	    RECT 155.1000 24.7500 156.9000 24.9000 ;
	    RECT 49.5000 23.2500 156.9000 24.7500 ;
	    RECT 49.5000 23.1000 51.3000 23.2500 ;
	    RECT 155.1000 23.1000 156.9000 23.2500 ;
	    RECT 332.7000 24.7500 334.5000 24.9000 ;
	    RECT 349.5000 24.7500 351.3000 24.9000 ;
	    RECT 332.7000 23.2500 351.3000 24.7500 ;
	    RECT 332.7000 23.1000 334.5000 23.2500 ;
	    RECT 349.5000 23.1000 351.3000 23.2500 ;
	    RECT 486.3000 24.7500 488.1000 24.9000 ;
	    RECT 519.9000 24.7500 521.7000 24.9000 ;
	    RECT 486.3000 23.2500 521.7000 24.7500 ;
	    RECT 486.3000 23.1000 488.1000 23.2500 ;
	    RECT 519.9000 23.1000 521.7000 23.2500 ;
	    RECT 577.5000 24.7500 579.3000 24.9000 ;
	    RECT 582.3000 24.7500 584.1000 24.9000 ;
	    RECT 577.5000 23.2500 584.1000 24.7500 ;
	    RECT 577.5000 23.1000 579.3000 23.2500 ;
	    RECT 582.3000 23.1000 584.1000 23.2500 ;
	    RECT 747.9000 24.7500 749.7000 24.9000 ;
	    RECT 771.9000 24.7500 773.7000 24.9000 ;
	    RECT 747.9000 23.2500 773.7000 24.7500 ;
	    RECT 747.9000 23.1000 749.7000 23.2500 ;
	    RECT 771.9000 23.1000 773.7000 23.2500 ;
	    RECT 1007.1000 24.7500 1008.9000 24.9000 ;
	    RECT 1043.1000 24.7500 1044.9000 24.9000 ;
	    RECT 1007.1000 23.2500 1044.9000 24.7500 ;
	    RECT 1007.1000 23.1000 1008.9000 23.2500 ;
	    RECT 1043.1000 23.1000 1044.9000 23.2500 ;
	    RECT 1208.7001 24.7500 1210.5000 24.9000 ;
	    RECT 1225.5000 24.7500 1227.3000 24.9000 ;
	    RECT 1208.7001 23.2500 1227.3000 24.7500 ;
	    RECT 1208.7001 23.1000 1210.5000 23.2500 ;
	    RECT 1225.5000 23.1000 1227.3000 23.2500 ;
	    RECT 1287.9000 24.7500 1289.7001 24.9000 ;
	    RECT 1304.7001 24.7500 1306.5000 24.9000 ;
	    RECT 1328.7001 24.7500 1330.5000 24.9000 ;
	    RECT 1287.9000 23.2500 1330.5000 24.7500 ;
	    RECT 1287.9000 23.1000 1289.7001 23.2500 ;
	    RECT 1304.7001 23.1000 1306.5000 23.2500 ;
	    RECT 1328.7001 23.1000 1330.5000 23.2500 ;
	    RECT 1371.9000 24.7500 1373.7001 24.9000 ;
	    RECT 1470.3000 24.7500 1472.1000 24.9000 ;
	    RECT 1371.9000 23.2500 1472.1000 24.7500 ;
	    RECT 1371.9000 23.1000 1373.7001 23.2500 ;
	    RECT 1470.3000 23.1000 1472.1000 23.2500 ;
	    RECT 164.7000 18.7500 166.5000 18.9000 ;
	    RECT 347.1000 18.7500 348.9000 18.9000 ;
	    RECT 164.7000 17.2500 348.9000 18.7500 ;
	    RECT 164.7000 17.1000 166.5000 17.2500 ;
	    RECT 347.1000 17.1000 348.9000 17.2500 ;
	    RECT 594.3000 18.7500 596.1000 18.9000 ;
	    RECT 738.3000 18.7500 740.1000 18.9000 ;
	    RECT 594.3000 17.2500 740.1000 18.7500 ;
	    RECT 594.3000 17.1000 596.1000 17.2500 ;
	    RECT 738.3000 17.1000 740.1000 17.2500 ;
	    RECT 855.9000 18.7500 857.7000 18.9000 ;
	    RECT 891.9000 18.7500 893.7000 18.9000 ;
	    RECT 855.9000 17.2500 893.7000 18.7500 ;
	    RECT 855.9000 17.1000 857.7000 17.2500 ;
	    RECT 891.9000 17.1000 893.7000 17.2500 ;
	    RECT 987.9000 18.7500 989.7000 18.9000 ;
	    RECT 1033.5000 18.7500 1035.3000 18.9000 ;
	    RECT 987.9000 17.2500 1035.3000 18.7500 ;
	    RECT 987.9000 17.1000 989.7000 17.2500 ;
	    RECT 1033.5000 17.1000 1035.3000 17.2500 ;
	    RECT 1275.9000 18.7500 1277.7001 18.9000 ;
	    RECT 1280.7001 18.7500 1282.5000 18.9000 ;
	    RECT 1302.3000 18.7500 1304.1000 18.9000 ;
	    RECT 1275.9000 17.2500 1304.1000 18.7500 ;
	    RECT 1275.9000 17.1000 1277.7001 17.2500 ;
	    RECT 1280.7001 17.1000 1282.5000 17.2500 ;
	    RECT 1302.3000 17.1000 1304.1000 17.2500 ;
	    RECT 1479.9000 18.7500 1481.7001 18.9000 ;
	    RECT 1511.1000 18.7500 1512.9000 18.9000 ;
	    RECT 1479.9000 17.2500 1512.9000 18.7500 ;
	    RECT 1479.9000 17.1000 1481.7001 17.2500 ;
	    RECT 1511.1000 17.1000 1512.9000 17.2500 ;
	    RECT 1515.9000 18.7500 1517.7001 18.9000 ;
	    RECT 1551.9000 18.7500 1553.7001 18.9000 ;
	    RECT 1515.9000 17.2500 1553.7001 18.7500 ;
	    RECT 1515.9000 17.1000 1517.7001 17.2500 ;
	    RECT 1551.9000 17.1000 1553.7001 17.2500 ;
	    RECT 395.1000 12.7500 396.9000 12.9000 ;
	    RECT 529.5000 12.7500 531.3000 12.9000 ;
	    RECT 395.1000 11.2500 531.3000 12.7500 ;
	    RECT 395.1000 11.1000 396.9000 11.2500 ;
	    RECT 529.5000 11.1000 531.3000 11.2500 ;
	    RECT 776.7000 12.7500 778.5000 12.9000 ;
	    RECT 795.9000 12.7500 797.7000 12.9000 ;
	    RECT 776.7000 11.2500 797.7000 12.7500 ;
	    RECT 776.7000 11.1000 778.5000 11.2500 ;
	    RECT 795.9000 11.1000 797.7000 11.2500 ;
	    RECT 1194.3000 12.7500 1196.1000 12.9000 ;
	    RECT 1254.3000 12.7500 1256.1000 12.9000 ;
	    RECT 1194.3000 11.2500 1256.1000 12.7500 ;
	    RECT 1194.3000 11.1000 1196.1000 11.2500 ;
	    RECT 1254.3000 11.1000 1256.1000 11.2500 ;
	    RECT 829.5000 6.7500 831.3000 6.9000 ;
	    RECT 1026.3000 6.7500 1028.1000 6.9000 ;
	    RECT 829.5000 5.2500 1028.1000 6.7500 ;
	    RECT 829.5000 5.1000 831.3000 5.2500 ;
	    RECT 1026.3000 5.1000 1028.1000 5.2500 ;
	    RECT 1542.3000 6.7500 1544.1000 6.9000 ;
	    RECT 1566.3000 6.7500 1568.1000 6.9000 ;
	    RECT 1542.3000 5.2500 1568.1000 6.7500 ;
	    RECT 1542.3000 5.1000 1544.1000 5.2500 ;
	    RECT 1566.3000 5.1000 1568.1000 5.2500 ;
   END
END FIR
