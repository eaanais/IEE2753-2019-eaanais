module FIR ( gnd, vdd, clk, rst, din, dout);

input gnd, vdd;
input clk;
input rst;
input [7:0] din;
output [7:0] dout;

CLKBUF1 CLKBUF1_1 ( .gnd(gnd), .vdd(vdd), .A(asr2_clk), .Y(asr2_clk_bF_buf7) );
CLKBUF1 CLKBUF1_2 ( .gnd(gnd), .vdd(vdd), .A(asr2_clk), .Y(asr2_clk_bF_buf6) );
CLKBUF1 CLKBUF1_3 ( .gnd(gnd), .vdd(vdd), .A(asr2_clk), .Y(asr2_clk_bF_buf5) );
CLKBUF1 CLKBUF1_4 ( .gnd(gnd), .vdd(vdd), .A(asr2_clk), .Y(asr2_clk_bF_buf4) );
CLKBUF1 CLKBUF1_5 ( .gnd(gnd), .vdd(vdd), .A(asr2_clk), .Y(asr2_clk_bF_buf3) );
CLKBUF1 CLKBUF1_6 ( .gnd(gnd), .vdd(vdd), .A(asr2_clk), .Y(asr2_clk_bF_buf2) );
CLKBUF1 CLKBUF1_7 ( .gnd(gnd), .vdd(vdd), .A(asr2_clk), .Y(asr2_clk_bF_buf1) );
CLKBUF1 CLKBUF1_8 ( .gnd(gnd), .vdd(vdd), .A(asr2_clk), .Y(asr2_clk_bF_buf0) );
CLKBUF1 CLKBUF1_9 ( .gnd(gnd), .vdd(vdd), .A(clk), .Y(clk_bF_buf7) );
CLKBUF1 CLKBUF1_10 ( .gnd(gnd), .vdd(vdd), .A(clk), .Y(clk_bF_buf6) );
CLKBUF1 CLKBUF1_11 ( .gnd(gnd), .vdd(vdd), .A(clk), .Y(clk_bF_buf5) );
CLKBUF1 CLKBUF1_12 ( .gnd(gnd), .vdd(vdd), .A(clk), .Y(clk_bF_buf4) );
CLKBUF1 CLKBUF1_13 ( .gnd(gnd), .vdd(vdd), .A(clk), .Y(clk_bF_buf3) );
CLKBUF1 CLKBUF1_14 ( .gnd(gnd), .vdd(vdd), .A(clk), .Y(clk_bF_buf2) );
CLKBUF1 CLKBUF1_15 ( .gnd(gnd), .vdd(vdd), .A(clk), .Y(clk_bF_buf1) );
CLKBUF1 CLKBUF1_16 ( .gnd(gnd), .vdd(vdd), .A(clk), .Y(clk_bF_buf0) );
BUFX2 BUFX2_1 ( .gnd(gnd), .vdd(vdd), .A(MAC_clr), .Y(MAC_clr_bF_buf3) );
BUFX2 BUFX2_2 ( .gnd(gnd), .vdd(vdd), .A(MAC_clr), .Y(MAC_clr_bF_buf2) );
BUFX2 BUFX2_3 ( .gnd(gnd), .vdd(vdd), .A(MAC_clr), .Y(MAC_clr_bF_buf1) );
BUFX2 BUFX2_4 ( .gnd(gnd), .vdd(vdd), .A(MAC_clr), .Y(MAC_clr_bF_buf0) );
CLKBUF1 CLKBUF1_17 ( .gnd(gnd), .vdd(vdd), .A(asr1_clk), .Y(asr1_clk_bF_buf8) );
CLKBUF1 CLKBUF1_18 ( .gnd(gnd), .vdd(vdd), .A(asr1_clk), .Y(asr1_clk_bF_buf7) );
CLKBUF1 CLKBUF1_19 ( .gnd(gnd), .vdd(vdd), .A(asr1_clk), .Y(asr1_clk_bF_buf6) );
CLKBUF1 CLKBUF1_20 ( .gnd(gnd), .vdd(vdd), .A(asr1_clk), .Y(asr1_clk_bF_buf5) );
CLKBUF1 CLKBUF1_21 ( .gnd(gnd), .vdd(vdd), .A(asr1_clk), .Y(asr1_clk_bF_buf4) );
CLKBUF1 CLKBUF1_22 ( .gnd(gnd), .vdd(vdd), .A(asr1_clk), .Y(asr1_clk_bF_buf3) );
CLKBUF1 CLKBUF1_23 ( .gnd(gnd), .vdd(vdd), .A(asr1_clk), .Y(asr1_clk_bF_buf2) );
CLKBUF1 CLKBUF1_24 ( .gnd(gnd), .vdd(vdd), .A(asr1_clk), .Y(asr1_clk_bF_buf1) );
CLKBUF1 CLKBUF1_25 ( .gnd(gnd), .vdd(vdd), .A(asr1_clk), .Y(asr1_clk_bF_buf0) );
BUFX2 BUFX2_5 ( .gnd(gnd), .vdd(vdd), .A(rst), .Y(rst_bF_buf5) );
BUFX2 BUFX2_6 ( .gnd(gnd), .vdd(vdd), .A(rst), .Y(rst_bF_buf4) );
BUFX2 BUFX2_7 ( .gnd(gnd), .vdd(vdd), .A(rst), .Y(rst_bF_buf3) );
BUFX2 BUFX2_8 ( .gnd(gnd), .vdd(vdd), .A(rst), .Y(rst_bF_buf2) );
BUFX2 BUFX2_9 ( .gnd(gnd), .vdd(vdd), .A(rst), .Y(rst_bF_buf1) );
BUFX2 BUFX2_10 ( .gnd(gnd), .vdd(vdd), .A(rst), .Y(rst_bF_buf0) );
BUFX2 BUFX2_11 ( .gnd(gnd), .vdd(vdd), .A(MAC_ROM_0_), .Y(MAC_ROM_0_bF_buf3_) );
BUFX2 BUFX2_12 ( .gnd(gnd), .vdd(vdd), .A(MAC_ROM_0_), .Y(MAC_ROM_0_bF_buf2_) );
BUFX2 BUFX2_13 ( .gnd(gnd), .vdd(vdd), .A(MAC_ROM_0_), .Y(MAC_ROM_0_bF_buf1_) );
BUFX2 BUFX2_14 ( .gnd(gnd), .vdd(vdd), .A(MAC_ROM_0_), .Y(MAC_ROM_0_bF_buf0_) );
BUFX2 BUFX2_15 ( .gnd(gnd), .vdd(vdd), .A(asr2_en), .Y(asr2_en_bF_buf10) );
BUFX2 BUFX2_16 ( .gnd(gnd), .vdd(vdd), .A(asr2_en), .Y(asr2_en_bF_buf9) );
BUFX2 BUFX2_17 ( .gnd(gnd), .vdd(vdd), .A(asr2_en), .Y(asr2_en_bF_buf8) );
BUFX2 BUFX2_18 ( .gnd(gnd), .vdd(vdd), .A(asr2_en), .Y(asr2_en_bF_buf7) );
BUFX2 BUFX2_19 ( .gnd(gnd), .vdd(vdd), .A(asr2_en), .Y(asr2_en_bF_buf6) );
BUFX2 BUFX2_20 ( .gnd(gnd), .vdd(vdd), .A(asr2_en), .Y(asr2_en_bF_buf5) );
BUFX2 BUFX2_21 ( .gnd(gnd), .vdd(vdd), .A(asr2_en), .Y(asr2_en_bF_buf4) );
BUFX2 BUFX2_22 ( .gnd(gnd), .vdd(vdd), .A(asr2_en), .Y(asr2_en_bF_buf3) );
BUFX2 BUFX2_23 ( .gnd(gnd), .vdd(vdd), .A(asr2_en), .Y(asr2_en_bF_buf2) );
BUFX2 BUFX2_24 ( .gnd(gnd), .vdd(vdd), .A(asr2_en), .Y(asr2_en_bF_buf1) );
BUFX2 BUFX2_25 ( .gnd(gnd), .vdd(vdd), .A(asr2_en), .Y(asr2_en_bF_buf0) );
NOR2X1 NOR2X1_1 ( .gnd(gnd), .vdd(vdd), .A(up_counter_contador_1_), .B(up_counter_contador_0_), .Y(_1_) );
NOR2X1 NOR2X1_2 ( .gnd(gnd), .vdd(vdd), .A(up_counter_contador_2_), .B(rst_bF_buf1), .Y(_2_) );
AND2X2 AND2X2_1 ( .gnd(gnd), .vdd(vdd), .A(_1_), .B(_2_), .Y(_0_) );
INVX1 INVX1_1 ( .gnd(gnd), .vdd(vdd), .A(asr1_clk_bF_buf6), .Y(asr2_en) );
BUFX2 BUFX2_26 ( .gnd(gnd), .vdd(vdd), .A(_3__0_), .Y(dout[0]) );
BUFX2 BUFX2_27 ( .gnd(gnd), .vdd(vdd), .A(_3__1_), .Y(dout[1]) );
BUFX2 BUFX2_28 ( .gnd(gnd), .vdd(vdd), .A(_3__2_), .Y(dout[2]) );
BUFX2 BUFX2_29 ( .gnd(gnd), .vdd(vdd), .A(_3__3_), .Y(dout[3]) );
BUFX2 BUFX2_30 ( .gnd(gnd), .vdd(vdd), .A(_3__4_), .Y(dout[4]) );
BUFX2 BUFX2_31 ( .gnd(gnd), .vdd(vdd), .A(_3__5_), .Y(dout[5]) );
BUFX2 BUFX2_32 ( .gnd(gnd), .vdd(vdd), .A(_3__6_), .Y(dout[6]) );
BUFX2 BUFX2_33 ( .gnd(gnd), .vdd(vdd), .A(_3__7_), .Y(dout[7]) );
DFFPOSX1 DFFPOSX1_1 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf4), .D(_0_), .Q(enable_asr) );
INVX1 INVX1_2 ( .gnd(gnd), .vdd(vdd), .A(asr1_cables_1__0_), .Y(_6_) );
NAND2X1 NAND2X1_1 ( .gnd(gnd), .vdd(vdd), .A(asr1_cables_0__0_), .B(vdd), .Y(_7_) );
OAI21X1 OAI21X1_1 ( .gnd(gnd), .vdd(vdd), .A(vdd), .B(_6_), .C(_7_), .Y(_4__0_) );
INVX1 INVX1_3 ( .gnd(gnd), .vdd(vdd), .A(asr1_cables_1__1_), .Y(_8_) );
NAND2X1 NAND2X1_2 ( .gnd(gnd), .vdd(vdd), .A(vdd), .B(asr1_cables_0__1_), .Y(_9_) );
OAI21X1 OAI21X1_2 ( .gnd(gnd), .vdd(vdd), .A(vdd), .B(_8_), .C(_9_), .Y(_4__1_) );
INVX1 INVX1_4 ( .gnd(gnd), .vdd(vdd), .A(asr1_cables_1__2_), .Y(_10_) );
NAND2X1 NAND2X1_3 ( .gnd(gnd), .vdd(vdd), .A(vdd), .B(asr1_cables_0__2_), .Y(_11_) );
OAI21X1 OAI21X1_3 ( .gnd(gnd), .vdd(vdd), .A(vdd), .B(_10_), .C(_11_), .Y(_4__2_) );
INVX1 INVX1_5 ( .gnd(gnd), .vdd(vdd), .A(asr1_cables_1__3_), .Y(_12_) );
NAND2X1 NAND2X1_4 ( .gnd(gnd), .vdd(vdd), .A(vdd), .B(asr1_cables_0__3_), .Y(_13_) );
OAI21X1 OAI21X1_4 ( .gnd(gnd), .vdd(vdd), .A(vdd), .B(_12_), .C(_13_), .Y(_4__3_) );
INVX1 INVX1_6 ( .gnd(gnd), .vdd(vdd), .A(asr1_cables_1__4_), .Y(_14_) );
NAND2X1 NAND2X1_5 ( .gnd(gnd), .vdd(vdd), .A(vdd), .B(asr1_cables_0__4_), .Y(_15_) );
OAI21X1 OAI21X1_5 ( .gnd(gnd), .vdd(vdd), .A(vdd), .B(_14_), .C(_15_), .Y(_4__4_) );
INVX1 INVX1_7 ( .gnd(gnd), .vdd(vdd), .A(asr1_cables_1__5_), .Y(_16_) );
NAND2X1 NAND2X1_6 ( .gnd(gnd), .vdd(vdd), .A(vdd), .B(asr1_cables_0__5_), .Y(_17_) );
OAI21X1 OAI21X1_6 ( .gnd(gnd), .vdd(vdd), .A(vdd), .B(_16_), .C(_17_), .Y(_4__5_) );
INVX1 INVX1_8 ( .gnd(gnd), .vdd(vdd), .A(asr1_cables_1__6_), .Y(_18_) );
NAND2X1 NAND2X1_7 ( .gnd(gnd), .vdd(vdd), .A(vdd), .B(asr1_cables_0__6_), .Y(_19_) );
OAI21X1 OAI21X1_7 ( .gnd(gnd), .vdd(vdd), .A(vdd), .B(_18_), .C(_19_), .Y(_4__6_) );
INVX1 INVX1_9 ( .gnd(gnd), .vdd(vdd), .A(asr1_cables_1__7_), .Y(_20_) );
NAND2X1 NAND2X1_8 ( .gnd(gnd), .vdd(vdd), .A(vdd), .B(asr1_cables_0__7_), .Y(_21_) );
OAI21X1 OAI21X1_8 ( .gnd(gnd), .vdd(vdd), .A(vdd), .B(_20_), .C(_21_), .Y(_4__7_) );
INVX1 INVX1_10 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf2), .Y(_5_) );
DFFSR DFFSR_1 ( .gnd(gnd), .vdd(vdd), .CLK(asr1_clk_bF_buf4), .D(_4__0_), .Q(asr1_cables_1__0_), .R(_5_), .S(vdd) );
DFFSR DFFSR_2 ( .gnd(gnd), .vdd(vdd), .CLK(asr1_clk_bF_buf8), .D(_4__1_), .Q(asr1_cables_1__1_), .R(_5_), .S(vdd) );
DFFSR DFFSR_3 ( .gnd(gnd), .vdd(vdd), .CLK(asr1_clk_bF_buf5), .D(_4__2_), .Q(asr1_cables_1__2_), .R(_5_), .S(vdd) );
DFFSR DFFSR_4 ( .gnd(gnd), .vdd(vdd), .CLK(asr1_clk_bF_buf8), .D(_4__3_), .Q(asr1_cables_1__3_), .R(_5_), .S(vdd) );
DFFSR DFFSR_5 ( .gnd(gnd), .vdd(vdd), .CLK(asr1_clk_bF_buf7), .D(_4__4_), .Q(asr1_cables_1__4_), .R(_5_), .S(vdd) );
DFFSR DFFSR_6 ( .gnd(gnd), .vdd(vdd), .CLK(asr1_clk_bF_buf8), .D(_4__5_), .Q(asr1_cables_1__5_), .R(_5_), .S(vdd) );
DFFSR DFFSR_7 ( .gnd(gnd), .vdd(vdd), .CLK(asr1_clk_bF_buf6), .D(_4__6_), .Q(asr1_cables_1__6_), .R(_5_), .S(vdd) );
DFFSR DFFSR_8 ( .gnd(gnd), .vdd(vdd), .CLK(asr1_clk_bF_buf4), .D(_4__7_), .Q(asr1_cables_1__7_), .R(_5_), .S(vdd) );
INVX1 INVX1_11 ( .gnd(gnd), .vdd(vdd), .A(asr1_cables_2__0_), .Y(_24_) );
NAND2X1 NAND2X1_9 ( .gnd(gnd), .vdd(vdd), .A(asr1_cables_1__0_), .B(vdd), .Y(_25_) );
OAI21X1 OAI21X1_9 ( .gnd(gnd), .vdd(vdd), .A(vdd), .B(_24_), .C(_25_), .Y(_22__0_) );
INVX1 INVX1_12 ( .gnd(gnd), .vdd(vdd), .A(asr1_cables_2__1_), .Y(_26_) );
NAND2X1 NAND2X1_10 ( .gnd(gnd), .vdd(vdd), .A(vdd), .B(asr1_cables_1__1_), .Y(_27_) );
OAI21X1 OAI21X1_10 ( .gnd(gnd), .vdd(vdd), .A(vdd), .B(_26_), .C(_27_), .Y(_22__1_) );
INVX1 INVX1_13 ( .gnd(gnd), .vdd(vdd), .A(asr1_cables_2__2_), .Y(_28_) );
NAND2X1 NAND2X1_11 ( .gnd(gnd), .vdd(vdd), .A(vdd), .B(asr1_cables_1__2_), .Y(_29_) );
OAI21X1 OAI21X1_11 ( .gnd(gnd), .vdd(vdd), .A(vdd), .B(_28_), .C(_29_), .Y(_22__2_) );
INVX1 INVX1_14 ( .gnd(gnd), .vdd(vdd), .A(asr1_cables_2__3_), .Y(_30_) );
NAND2X1 NAND2X1_12 ( .gnd(gnd), .vdd(vdd), .A(vdd), .B(asr1_cables_1__3_), .Y(_31_) );
OAI21X1 OAI21X1_12 ( .gnd(gnd), .vdd(vdd), .A(vdd), .B(_30_), .C(_31_), .Y(_22__3_) );
INVX1 INVX1_15 ( .gnd(gnd), .vdd(vdd), .A(asr1_cables_2__4_), .Y(_32_) );
NAND2X1 NAND2X1_13 ( .gnd(gnd), .vdd(vdd), .A(vdd), .B(asr1_cables_1__4_), .Y(_33_) );
OAI21X1 OAI21X1_13 ( .gnd(gnd), .vdd(vdd), .A(vdd), .B(_32_), .C(_33_), .Y(_22__4_) );
INVX1 INVX1_16 ( .gnd(gnd), .vdd(vdd), .A(asr1_cables_2__5_), .Y(_34_) );
NAND2X1 NAND2X1_14 ( .gnd(gnd), .vdd(vdd), .A(vdd), .B(asr1_cables_1__5_), .Y(_35_) );
OAI21X1 OAI21X1_14 ( .gnd(gnd), .vdd(vdd), .A(vdd), .B(_34_), .C(_35_), .Y(_22__5_) );
INVX1 INVX1_17 ( .gnd(gnd), .vdd(vdd), .A(asr1_cables_2__6_), .Y(_36_) );
NAND2X1 NAND2X1_15 ( .gnd(gnd), .vdd(vdd), .A(vdd), .B(asr1_cables_1__6_), .Y(_37_) );
OAI21X1 OAI21X1_15 ( .gnd(gnd), .vdd(vdd), .A(vdd), .B(_36_), .C(_37_), .Y(_22__6_) );
INVX1 INVX1_18 ( .gnd(gnd), .vdd(vdd), .A(asr1_cables_2__7_), .Y(_38_) );
NAND2X1 NAND2X1_16 ( .gnd(gnd), .vdd(vdd), .A(vdd), .B(asr1_cables_1__7_), .Y(_39_) );
OAI21X1 OAI21X1_16 ( .gnd(gnd), .vdd(vdd), .A(vdd), .B(_38_), .C(_39_), .Y(_22__7_) );
INVX1 INVX1_19 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf2), .Y(_23_) );
DFFSR DFFSR_9 ( .gnd(gnd), .vdd(vdd), .CLK(asr1_clk_bF_buf1), .D(_22__0_), .Q(asr1_cables_2__0_), .R(_23_), .S(vdd) );
DFFSR DFFSR_10 ( .gnd(gnd), .vdd(vdd), .CLK(asr1_clk_bF_buf7), .D(_22__1_), .Q(asr1_cables_2__1_), .R(_23_), .S(vdd) );
DFFSR DFFSR_11 ( .gnd(gnd), .vdd(vdd), .CLK(asr1_clk_bF_buf3), .D(_22__2_), .Q(asr1_cables_2__2_), .R(_23_), .S(vdd) );
DFFSR DFFSR_12 ( .gnd(gnd), .vdd(vdd), .CLK(asr1_clk_bF_buf2), .D(_22__3_), .Q(asr1_cables_2__3_), .R(_23_), .S(vdd) );
DFFSR DFFSR_13 ( .gnd(gnd), .vdd(vdd), .CLK(asr1_clk_bF_buf7), .D(_22__4_), .Q(asr1_cables_2__4_), .R(_23_), .S(vdd) );
DFFSR DFFSR_14 ( .gnd(gnd), .vdd(vdd), .CLK(asr1_clk_bF_buf8), .D(_22__5_), .Q(asr1_cables_2__5_), .R(_23_), .S(vdd) );
DFFSR DFFSR_15 ( .gnd(gnd), .vdd(vdd), .CLK(asr1_clk_bF_buf6), .D(_22__6_), .Q(asr1_cables_2__6_), .R(_23_), .S(vdd) );
DFFSR DFFSR_16 ( .gnd(gnd), .vdd(vdd), .CLK(asr1_clk_bF_buf2), .D(_22__7_), .Q(asr1_cables_2__7_), .R(_23_), .S(vdd) );
INVX1 INVX1_20 ( .gnd(gnd), .vdd(vdd), .A(asr1_cables_3__0_), .Y(_42_) );
NAND2X1 NAND2X1_17 ( .gnd(gnd), .vdd(vdd), .A(asr1_cables_2__0_), .B(vdd), .Y(_43_) );
OAI21X1 OAI21X1_17 ( .gnd(gnd), .vdd(vdd), .A(vdd), .B(_42_), .C(_43_), .Y(_40__0_) );
INVX1 INVX1_21 ( .gnd(gnd), .vdd(vdd), .A(asr1_cables_3__1_), .Y(_44_) );
NAND2X1 NAND2X1_18 ( .gnd(gnd), .vdd(vdd), .A(vdd), .B(asr1_cables_2__1_), .Y(_45_) );
OAI21X1 OAI21X1_18 ( .gnd(gnd), .vdd(vdd), .A(vdd), .B(_44_), .C(_45_), .Y(_40__1_) );
INVX1 INVX1_22 ( .gnd(gnd), .vdd(vdd), .A(asr1_cables_3__2_), .Y(_46_) );
NAND2X1 NAND2X1_19 ( .gnd(gnd), .vdd(vdd), .A(vdd), .B(asr1_cables_2__2_), .Y(_47_) );
OAI21X1 OAI21X1_19 ( .gnd(gnd), .vdd(vdd), .A(vdd), .B(_46_), .C(_47_), .Y(_40__2_) );
INVX1 INVX1_23 ( .gnd(gnd), .vdd(vdd), .A(asr1_cables_3__3_), .Y(_48_) );
NAND2X1 NAND2X1_20 ( .gnd(gnd), .vdd(vdd), .A(vdd), .B(asr1_cables_2__3_), .Y(_49_) );
OAI21X1 OAI21X1_20 ( .gnd(gnd), .vdd(vdd), .A(vdd), .B(_48_), .C(_49_), .Y(_40__3_) );
INVX1 INVX1_24 ( .gnd(gnd), .vdd(vdd), .A(asr1_cables_3__4_), .Y(_50_) );
NAND2X1 NAND2X1_21 ( .gnd(gnd), .vdd(vdd), .A(vdd), .B(asr1_cables_2__4_), .Y(_51_) );
OAI21X1 OAI21X1_21 ( .gnd(gnd), .vdd(vdd), .A(vdd), .B(_50_), .C(_51_), .Y(_40__4_) );
INVX1 INVX1_25 ( .gnd(gnd), .vdd(vdd), .A(asr1_cables_3__5_), .Y(_52_) );
NAND2X1 NAND2X1_22 ( .gnd(gnd), .vdd(vdd), .A(vdd), .B(asr1_cables_2__5_), .Y(_53_) );
OAI21X1 OAI21X1_22 ( .gnd(gnd), .vdd(vdd), .A(vdd), .B(_52_), .C(_53_), .Y(_40__5_) );
INVX1 INVX1_26 ( .gnd(gnd), .vdd(vdd), .A(asr1_cables_3__6_), .Y(_54_) );
NAND2X1 NAND2X1_23 ( .gnd(gnd), .vdd(vdd), .A(vdd), .B(asr1_cables_2__6_), .Y(_55_) );
OAI21X1 OAI21X1_23 ( .gnd(gnd), .vdd(vdd), .A(vdd), .B(_54_), .C(_55_), .Y(_40__6_) );
INVX1 INVX1_27 ( .gnd(gnd), .vdd(vdd), .A(asr1_cables_3__7_), .Y(_56_) );
NAND2X1 NAND2X1_24 ( .gnd(gnd), .vdd(vdd), .A(vdd), .B(asr1_cables_2__7_), .Y(_57_) );
OAI21X1 OAI21X1_24 ( .gnd(gnd), .vdd(vdd), .A(vdd), .B(_56_), .C(_57_), .Y(_40__7_) );
INVX1 INVX1_28 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf2), .Y(_41_) );
DFFSR DFFSR_17 ( .gnd(gnd), .vdd(vdd), .CLK(asr1_clk_bF_buf1), .D(_40__0_), .Q(asr1_cables_3__0_), .R(_41_), .S(vdd) );
DFFSR DFFSR_18 ( .gnd(gnd), .vdd(vdd), .CLK(asr1_clk_bF_buf3), .D(_40__1_), .Q(asr1_cables_3__1_), .R(_41_), .S(vdd) );
DFFSR DFFSR_19 ( .gnd(gnd), .vdd(vdd), .CLK(asr1_clk_bF_buf3), .D(_40__2_), .Q(asr1_cables_3__2_), .R(_41_), .S(vdd) );
DFFSR DFFSR_20 ( .gnd(gnd), .vdd(vdd), .CLK(asr1_clk_bF_buf5), .D(_40__3_), .Q(asr1_cables_3__3_), .R(_41_), .S(vdd) );
DFFSR DFFSR_21 ( .gnd(gnd), .vdd(vdd), .CLK(asr1_clk_bF_buf8), .D(_40__4_), .Q(asr1_cables_3__4_), .R(_41_), .S(vdd) );
DFFSR DFFSR_22 ( .gnd(gnd), .vdd(vdd), .CLK(asr1_clk_bF_buf8), .D(_40__5_), .Q(asr1_cables_3__5_), .R(_41_), .S(vdd) );
DFFSR DFFSR_23 ( .gnd(gnd), .vdd(vdd), .CLK(asr1_clk_bF_buf4), .D(_40__6_), .Q(asr1_cables_3__6_), .R(_41_), .S(vdd) );
DFFSR DFFSR_24 ( .gnd(gnd), .vdd(vdd), .CLK(asr1_clk_bF_buf5), .D(_40__7_), .Q(asr1_cables_3__7_), .R(_41_), .S(vdd) );
INVX1 INVX1_29 ( .gnd(gnd), .vdd(vdd), .A(asr1_cables_4_), .Y(_60_) );
NAND2X1 NAND2X1_25 ( .gnd(gnd), .vdd(vdd), .A(asr1_cables_3__0_), .B(vdd), .Y(_61_) );
OAI21X1 OAI21X1_25 ( .gnd(gnd), .vdd(vdd), .A(vdd), .B(_60_), .C(_61_), .Y(_58__0_) );
INVX1 INVX1_30 ( .gnd(gnd), .vdd(vdd), .A(_76_), .Y(_62_) );
NAND2X1 NAND2X1_26 ( .gnd(gnd), .vdd(vdd), .A(vdd), .B(asr1_cables_3__1_), .Y(_63_) );
OAI21X1 OAI21X1_26 ( .gnd(gnd), .vdd(vdd), .A(vdd), .B(_62_), .C(_63_), .Y(_58__1_) );
INVX1 INVX1_31 ( .gnd(gnd), .vdd(vdd), .A(_82_), .Y(_64_) );
NAND2X1 NAND2X1_27 ( .gnd(gnd), .vdd(vdd), .A(vdd), .B(asr1_cables_3__2_), .Y(_65_) );
OAI21X1 OAI21X1_27 ( .gnd(gnd), .vdd(vdd), .A(vdd), .B(_64_), .C(_65_), .Y(_58__2_) );
INVX1 INVX1_32 ( .gnd(gnd), .vdd(vdd), .A(_77_), .Y(_66_) );
NAND2X1 NAND2X1_28 ( .gnd(gnd), .vdd(vdd), .A(vdd), .B(asr1_cables_3__3_), .Y(_67_) );
OAI21X1 OAI21X1_28 ( .gnd(gnd), .vdd(vdd), .A(vdd), .B(_66_), .C(_67_), .Y(_58__3_) );
INVX1 INVX1_33 ( .gnd(gnd), .vdd(vdd), .A(_78_), .Y(_68_) );
NAND2X1 NAND2X1_29 ( .gnd(gnd), .vdd(vdd), .A(vdd), .B(asr1_cables_3__4_), .Y(_69_) );
OAI21X1 OAI21X1_29 ( .gnd(gnd), .vdd(vdd), .A(vdd), .B(_68_), .C(_69_), .Y(_58__4_) );
INVX1 INVX1_34 ( .gnd(gnd), .vdd(vdd), .A(_79_), .Y(_70_) );
NAND2X1 NAND2X1_30 ( .gnd(gnd), .vdd(vdd), .A(vdd), .B(asr1_cables_3__5_), .Y(_71_) );
OAI21X1 OAI21X1_30 ( .gnd(gnd), .vdd(vdd), .A(vdd), .B(_70_), .C(_71_), .Y(_58__5_) );
INVX1 INVX1_35 ( .gnd(gnd), .vdd(vdd), .A(_80_), .Y(_72_) );
NAND2X1 NAND2X1_31 ( .gnd(gnd), .vdd(vdd), .A(vdd), .B(asr1_cables_3__6_), .Y(_73_) );
OAI21X1 OAI21X1_31 ( .gnd(gnd), .vdd(vdd), .A(vdd), .B(_72_), .C(_73_), .Y(_58__6_) );
INVX1 INVX1_36 ( .gnd(gnd), .vdd(vdd), .A(_81_), .Y(_74_) );
NAND2X1 NAND2X1_32 ( .gnd(gnd), .vdd(vdd), .A(vdd), .B(asr1_cables_3__7_), .Y(_75_) );
OAI21X1 OAI21X1_32 ( .gnd(gnd), .vdd(vdd), .A(vdd), .B(_74_), .C(_75_), .Y(_58__7_) );
INVX1 INVX1_37 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf2), .Y(_59_) );
DFFSR DFFSR_25 ( .gnd(gnd), .vdd(vdd), .CLK(asr1_clk_bF_buf1), .D(_58__0_), .Q(asr1_cables_4_), .R(_59_), .S(vdd) );
DFFSR DFFSR_26 ( .gnd(gnd), .vdd(vdd), .CLK(asr1_clk_bF_buf5), .D(_58__1_), .Q(_76_), .R(_59_), .S(vdd) );
DFFSR DFFSR_27 ( .gnd(gnd), .vdd(vdd), .CLK(asr1_clk_bF_buf2), .D(_58__2_), .Q(_82_), .R(_59_), .S(vdd) );
DFFSR DFFSR_28 ( .gnd(gnd), .vdd(vdd), .CLK(asr1_clk_bF_buf3), .D(_58__3_), .Q(_77_), .R(_59_), .S(vdd) );
DFFSR DFFSR_29 ( .gnd(gnd), .vdd(vdd), .CLK(asr1_clk_bF_buf5), .D(_58__4_), .Q(_78_), .R(_59_), .S(vdd) );
DFFSR DFFSR_30 ( .gnd(gnd), .vdd(vdd), .CLK(asr1_clk_bF_buf7), .D(_58__5_), .Q(_79_), .R(_59_), .S(vdd) );
DFFSR DFFSR_31 ( .gnd(gnd), .vdd(vdd), .CLK(asr1_clk_bF_buf1), .D(_58__6_), .Q(_80_), .R(_59_), .S(vdd) );
DFFSR DFFSR_32 ( .gnd(gnd), .vdd(vdd), .CLK(asr1_clk_bF_buf5), .D(_58__7_), .Q(_81_), .R(_59_), .S(vdd) );
INVX1 INVX1_38 ( .gnd(gnd), .vdd(vdd), .A(asr1_cables_5__0_), .Y(_85_) );
NAND2X1 NAND2X1_33 ( .gnd(gnd), .vdd(vdd), .A(asr1_cables_4_), .B(vdd), .Y(_86_) );
OAI21X1 OAI21X1_33 ( .gnd(gnd), .vdd(vdd), .A(vdd), .B(_85_), .C(_86_), .Y(_83__0_) );
INVX1 INVX1_39 ( .gnd(gnd), .vdd(vdd), .A(asr1_cables_5__1_), .Y(_87_) );
NAND2X1 NAND2X1_34 ( .gnd(gnd), .vdd(vdd), .A(vdd), .B(_76_), .Y(_88_) );
OAI21X1 OAI21X1_34 ( .gnd(gnd), .vdd(vdd), .A(vdd), .B(_87_), .C(_88_), .Y(_83__1_) );
INVX1 INVX1_40 ( .gnd(gnd), .vdd(vdd), .A(asr1_cables_5__2_), .Y(_89_) );
NAND2X1 NAND2X1_35 ( .gnd(gnd), .vdd(vdd), .A(vdd), .B(_82_), .Y(_90_) );
OAI21X1 OAI21X1_35 ( .gnd(gnd), .vdd(vdd), .A(vdd), .B(_89_), .C(_90_), .Y(_83__2_) );
INVX1 INVX1_41 ( .gnd(gnd), .vdd(vdd), .A(asr1_cables_5__3_), .Y(_91_) );
NAND2X1 NAND2X1_36 ( .gnd(gnd), .vdd(vdd), .A(vdd), .B(_77_), .Y(_92_) );
OAI21X1 OAI21X1_36 ( .gnd(gnd), .vdd(vdd), .A(vdd), .B(_91_), .C(_92_), .Y(_83__3_) );
INVX1 INVX1_42 ( .gnd(gnd), .vdd(vdd), .A(asr1_cables_5__4_), .Y(_93_) );
NAND2X1 NAND2X1_37 ( .gnd(gnd), .vdd(vdd), .A(vdd), .B(_78_), .Y(_94_) );
OAI21X1 OAI21X1_37 ( .gnd(gnd), .vdd(vdd), .A(vdd), .B(_93_), .C(_94_), .Y(_83__4_) );
INVX1 INVX1_43 ( .gnd(gnd), .vdd(vdd), .A(asr1_cables_5__5_), .Y(_95_) );
NAND2X1 NAND2X1_38 ( .gnd(gnd), .vdd(vdd), .A(vdd), .B(_79_), .Y(_96_) );
OAI21X1 OAI21X1_38 ( .gnd(gnd), .vdd(vdd), .A(vdd), .B(_95_), .C(_96_), .Y(_83__5_) );
INVX1 INVX1_44 ( .gnd(gnd), .vdd(vdd), .A(asr1_cables_5__6_), .Y(_97_) );
NAND2X1 NAND2X1_39 ( .gnd(gnd), .vdd(vdd), .A(vdd), .B(_80_), .Y(_98_) );
OAI21X1 OAI21X1_39 ( .gnd(gnd), .vdd(vdd), .A(vdd), .B(_97_), .C(_98_), .Y(_83__6_) );
INVX1 INVX1_45 ( .gnd(gnd), .vdd(vdd), .A(asr1_cables_5__7_), .Y(_99_) );
NAND2X1 NAND2X1_40 ( .gnd(gnd), .vdd(vdd), .A(vdd), .B(_81_), .Y(_100_) );
OAI21X1 OAI21X1_40 ( .gnd(gnd), .vdd(vdd), .A(vdd), .B(_99_), .C(_100_), .Y(_83__7_) );
INVX1 INVX1_46 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf2), .Y(_84_) );
DFFSR DFFSR_33 ( .gnd(gnd), .vdd(vdd), .CLK(asr1_clk_bF_buf1), .D(_83__0_), .Q(asr1_cables_5__0_), .R(_84_), .S(vdd) );
DFFSR DFFSR_34 ( .gnd(gnd), .vdd(vdd), .CLK(asr1_clk_bF_buf2), .D(_83__1_), .Q(asr1_cables_5__1_), .R(_84_), .S(vdd) );
DFFSR DFFSR_35 ( .gnd(gnd), .vdd(vdd), .CLK(asr1_clk_bF_buf2), .D(_83__2_), .Q(asr1_cables_5__2_), .R(_84_), .S(vdd) );
DFFSR DFFSR_36 ( .gnd(gnd), .vdd(vdd), .CLK(asr1_clk_bF_buf6), .D(_83__3_), .Q(asr1_cables_5__3_), .R(_84_), .S(vdd) );
DFFSR DFFSR_37 ( .gnd(gnd), .vdd(vdd), .CLK(asr1_clk_bF_buf7), .D(_83__4_), .Q(asr1_cables_5__4_), .R(_84_), .S(vdd) );
DFFSR DFFSR_38 ( .gnd(gnd), .vdd(vdd), .CLK(asr1_clk_bF_buf7), .D(_83__5_), .Q(asr1_cables_5__5_), .R(_84_), .S(vdd) );
DFFSR DFFSR_39 ( .gnd(gnd), .vdd(vdd), .CLK(asr1_clk_bF_buf1), .D(_83__6_), .Q(asr1_cables_5__6_), .R(_84_), .S(vdd) );
DFFSR DFFSR_40 ( .gnd(gnd), .vdd(vdd), .CLK(asr1_clk_bF_buf2), .D(_83__7_), .Q(asr1_cables_5__7_), .R(_84_), .S(vdd) );
INVX1 INVX1_47 ( .gnd(gnd), .vdd(vdd), .A(asr1_cables_6__0_), .Y(_103_) );
NAND2X1 NAND2X1_41 ( .gnd(gnd), .vdd(vdd), .A(asr1_cables_5__0_), .B(vdd), .Y(_104_) );
OAI21X1 OAI21X1_41 ( .gnd(gnd), .vdd(vdd), .A(vdd), .B(_103_), .C(_104_), .Y(_101__0_) );
INVX1 INVX1_48 ( .gnd(gnd), .vdd(vdd), .A(asr1_cables_6__1_), .Y(_105_) );
NAND2X1 NAND2X1_42 ( .gnd(gnd), .vdd(vdd), .A(vdd), .B(asr1_cables_5__1_), .Y(_106_) );
OAI21X1 OAI21X1_42 ( .gnd(gnd), .vdd(vdd), .A(vdd), .B(_105_), .C(_106_), .Y(_101__1_) );
INVX1 INVX1_49 ( .gnd(gnd), .vdd(vdd), .A(asr1_cables_6__2_), .Y(_107_) );
NAND2X1 NAND2X1_43 ( .gnd(gnd), .vdd(vdd), .A(vdd), .B(asr1_cables_5__2_), .Y(_108_) );
OAI21X1 OAI21X1_43 ( .gnd(gnd), .vdd(vdd), .A(vdd), .B(_107_), .C(_108_), .Y(_101__2_) );
INVX1 INVX1_50 ( .gnd(gnd), .vdd(vdd), .A(asr1_cables_6__3_), .Y(_109_) );
NAND2X1 NAND2X1_44 ( .gnd(gnd), .vdd(vdd), .A(vdd), .B(asr1_cables_5__3_), .Y(_110_) );
OAI21X1 OAI21X1_44 ( .gnd(gnd), .vdd(vdd), .A(vdd), .B(_109_), .C(_110_), .Y(_101__3_) );
INVX1 INVX1_51 ( .gnd(gnd), .vdd(vdd), .A(asr1_cables_6__4_), .Y(_111_) );
NAND2X1 NAND2X1_45 ( .gnd(gnd), .vdd(vdd), .A(vdd), .B(asr1_cables_5__4_), .Y(_112_) );
OAI21X1 OAI21X1_45 ( .gnd(gnd), .vdd(vdd), .A(vdd), .B(_111_), .C(_112_), .Y(_101__4_) );
INVX1 INVX1_52 ( .gnd(gnd), .vdd(vdd), .A(asr1_cables_6__5_), .Y(_113_) );
NAND2X1 NAND2X1_46 ( .gnd(gnd), .vdd(vdd), .A(vdd), .B(asr1_cables_5__5_), .Y(_114_) );
OAI21X1 OAI21X1_46 ( .gnd(gnd), .vdd(vdd), .A(vdd), .B(_113_), .C(_114_), .Y(_101__5_) );
INVX1 INVX1_53 ( .gnd(gnd), .vdd(vdd), .A(asr1_cables_6__6_), .Y(_115_) );
NAND2X1 NAND2X1_47 ( .gnd(gnd), .vdd(vdd), .A(vdd), .B(asr1_cables_5__6_), .Y(_116_) );
OAI21X1 OAI21X1_47 ( .gnd(gnd), .vdd(vdd), .A(vdd), .B(_115_), .C(_116_), .Y(_101__6_) );
INVX1 INVX1_54 ( .gnd(gnd), .vdd(vdd), .A(asr1_cables_6__7_), .Y(_117_) );
NAND2X1 NAND2X1_48 ( .gnd(gnd), .vdd(vdd), .A(vdd), .B(asr1_cables_5__7_), .Y(_118_) );
OAI21X1 OAI21X1_48 ( .gnd(gnd), .vdd(vdd), .A(vdd), .B(_117_), .C(_118_), .Y(_101__7_) );
INVX1 INVX1_55 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf2), .Y(_102_) );
DFFSR DFFSR_41 ( .gnd(gnd), .vdd(vdd), .CLK(asr1_clk_bF_buf3), .D(_101__0_), .Q(asr1_cables_6__0_), .R(_102_), .S(vdd) );
DFFSR DFFSR_42 ( .gnd(gnd), .vdd(vdd), .CLK(asr1_clk_bF_buf2), .D(_101__1_), .Q(asr1_cables_6__1_), .R(_102_), .S(vdd) );
DFFSR DFFSR_43 ( .gnd(gnd), .vdd(vdd), .CLK(asr1_clk_bF_buf2), .D(_101__2_), .Q(asr1_cables_6__2_), .R(_102_), .S(vdd) );
DFFSR DFFSR_44 ( .gnd(gnd), .vdd(vdd), .CLK(asr1_clk_bF_buf3), .D(_101__3_), .Q(asr1_cables_6__3_), .R(_102_), .S(vdd) );
DFFSR DFFSR_45 ( .gnd(gnd), .vdd(vdd), .CLK(asr1_clk_bF_buf8), .D(_101__4_), .Q(asr1_cables_6__4_), .R(_102_), .S(vdd) );
DFFSR DFFSR_46 ( .gnd(gnd), .vdd(vdd), .CLK(asr1_clk_bF_buf3), .D(_101__5_), .Q(asr1_cables_6__5_), .R(_102_), .S(vdd) );
DFFSR DFFSR_47 ( .gnd(gnd), .vdd(vdd), .CLK(asr1_clk_bF_buf1), .D(_101__6_), .Q(asr1_cables_6__6_), .R(_102_), .S(vdd) );
DFFSR DFFSR_48 ( .gnd(gnd), .vdd(vdd), .CLK(asr1_clk_bF_buf5), .D(_101__7_), .Q(asr1_cables_6__7_), .R(_102_), .S(vdd) );
INVX1 INVX1_56 ( .gnd(gnd), .vdd(vdd), .A(asr1_cables_7__0_), .Y(_121_) );
NAND2X1 NAND2X1_49 ( .gnd(gnd), .vdd(vdd), .A(asr1_cables_6__0_), .B(vdd), .Y(_122_) );
OAI21X1 OAI21X1_49 ( .gnd(gnd), .vdd(vdd), .A(vdd), .B(_121_), .C(_122_), .Y(_119__0_) );
INVX1 INVX1_57 ( .gnd(gnd), .vdd(vdd), .A(asr1_cables_7__1_), .Y(_123_) );
NAND2X1 NAND2X1_50 ( .gnd(gnd), .vdd(vdd), .A(vdd), .B(asr1_cables_6__1_), .Y(_124_) );
OAI21X1 OAI21X1_50 ( .gnd(gnd), .vdd(vdd), .A(vdd), .B(_123_), .C(_124_), .Y(_119__1_) );
INVX1 INVX1_58 ( .gnd(gnd), .vdd(vdd), .A(asr1_cables_7__2_), .Y(_125_) );
NAND2X1 NAND2X1_51 ( .gnd(gnd), .vdd(vdd), .A(vdd), .B(asr1_cables_6__2_), .Y(_126_) );
OAI21X1 OAI21X1_51 ( .gnd(gnd), .vdd(vdd), .A(vdd), .B(_125_), .C(_126_), .Y(_119__2_) );
INVX1 INVX1_59 ( .gnd(gnd), .vdd(vdd), .A(asr1_cables_7__3_), .Y(_127_) );
NAND2X1 NAND2X1_52 ( .gnd(gnd), .vdd(vdd), .A(vdd), .B(asr1_cables_6__3_), .Y(_128_) );
OAI21X1 OAI21X1_52 ( .gnd(gnd), .vdd(vdd), .A(vdd), .B(_127_), .C(_128_), .Y(_119__3_) );
INVX1 INVX1_60 ( .gnd(gnd), .vdd(vdd), .A(asr1_cables_7__4_), .Y(_129_) );
NAND2X1 NAND2X1_53 ( .gnd(gnd), .vdd(vdd), .A(vdd), .B(asr1_cables_6__4_), .Y(_130_) );
OAI21X1 OAI21X1_53 ( .gnd(gnd), .vdd(vdd), .A(vdd), .B(_129_), .C(_130_), .Y(_119__4_) );
INVX1 INVX1_61 ( .gnd(gnd), .vdd(vdd), .A(asr1_cables_7__5_), .Y(_131_) );
NAND2X1 NAND2X1_54 ( .gnd(gnd), .vdd(vdd), .A(vdd), .B(asr1_cables_6__5_), .Y(_132_) );
OAI21X1 OAI21X1_54 ( .gnd(gnd), .vdd(vdd), .A(vdd), .B(_131_), .C(_132_), .Y(_119__5_) );
INVX1 INVX1_62 ( .gnd(gnd), .vdd(vdd), .A(asr1_cables_7__6_), .Y(_133_) );
NAND2X1 NAND2X1_55 ( .gnd(gnd), .vdd(vdd), .A(vdd), .B(asr1_cables_6__6_), .Y(_134_) );
OAI21X1 OAI21X1_55 ( .gnd(gnd), .vdd(vdd), .A(vdd), .B(_133_), .C(_134_), .Y(_119__6_) );
INVX1 INVX1_63 ( .gnd(gnd), .vdd(vdd), .A(asr1_cables_7__7_), .Y(_135_) );
NAND2X1 NAND2X1_56 ( .gnd(gnd), .vdd(vdd), .A(vdd), .B(asr1_cables_6__7_), .Y(_136_) );
OAI21X1 OAI21X1_56 ( .gnd(gnd), .vdd(vdd), .A(vdd), .B(_135_), .C(_136_), .Y(_119__7_) );
INVX1 INVX1_64 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf2), .Y(_120_) );
DFFSR DFFSR_49 ( .gnd(gnd), .vdd(vdd), .CLK(asr1_clk_bF_buf3), .D(_119__0_), .Q(asr1_cables_7__0_), .R(_120_), .S(vdd) );
DFFSR DFFSR_50 ( .gnd(gnd), .vdd(vdd), .CLK(asr1_clk_bF_buf4), .D(_119__1_), .Q(asr1_cables_7__1_), .R(_120_), .S(vdd) );
DFFSR DFFSR_51 ( .gnd(gnd), .vdd(vdd), .CLK(asr1_clk_bF_buf4), .D(_119__2_), .Q(asr1_cables_7__2_), .R(_120_), .S(vdd) );
DFFSR DFFSR_52 ( .gnd(gnd), .vdd(vdd), .CLK(asr1_clk_bF_buf6), .D(_119__3_), .Q(asr1_cables_7__3_), .R(_120_), .S(vdd) );
DFFSR DFFSR_53 ( .gnd(gnd), .vdd(vdd), .CLK(asr1_clk_bF_buf7), .D(_119__4_), .Q(asr1_cables_7__4_), .R(_120_), .S(vdd) );
DFFSR DFFSR_54 ( .gnd(gnd), .vdd(vdd), .CLK(asr1_clk_bF_buf3), .D(_119__5_), .Q(asr1_cables_7__5_), .R(_120_), .S(vdd) );
DFFSR DFFSR_55 ( .gnd(gnd), .vdd(vdd), .CLK(asr1_clk_bF_buf4), .D(_119__6_), .Q(asr1_cables_7__6_), .R(_120_), .S(vdd) );
DFFSR DFFSR_56 ( .gnd(gnd), .vdd(vdd), .CLK(asr1_clk_bF_buf7), .D(_119__7_), .Q(asr1_cables_7__7_), .R(_120_), .S(vdd) );
INVX1 INVX1_65 ( .gnd(gnd), .vdd(vdd), .A(asr1_cables_8__0_), .Y(_139_) );
NAND2X1 NAND2X1_57 ( .gnd(gnd), .vdd(vdd), .A(asr1_cables_7__0_), .B(vdd), .Y(_140_) );
OAI21X1 OAI21X1_57 ( .gnd(gnd), .vdd(vdd), .A(vdd), .B(_139_), .C(_140_), .Y(_137__0_) );
INVX1 INVX1_66 ( .gnd(gnd), .vdd(vdd), .A(asr1_cables_8__1_), .Y(_141_) );
NAND2X1 NAND2X1_58 ( .gnd(gnd), .vdd(vdd), .A(vdd), .B(asr1_cables_7__1_), .Y(_142_) );
OAI21X1 OAI21X1_58 ( .gnd(gnd), .vdd(vdd), .A(vdd), .B(_141_), .C(_142_), .Y(_137__1_) );
INVX1 INVX1_67 ( .gnd(gnd), .vdd(vdd), .A(asr1_cables_8__2_), .Y(_143_) );
NAND2X1 NAND2X1_59 ( .gnd(gnd), .vdd(vdd), .A(vdd), .B(asr1_cables_7__2_), .Y(_144_) );
OAI21X1 OAI21X1_59 ( .gnd(gnd), .vdd(vdd), .A(vdd), .B(_143_), .C(_144_), .Y(_137__2_) );
INVX1 INVX1_68 ( .gnd(gnd), .vdd(vdd), .A(asr1_cables_8__3_), .Y(_145_) );
NAND2X1 NAND2X1_60 ( .gnd(gnd), .vdd(vdd), .A(vdd), .B(asr1_cables_7__3_), .Y(_146_) );
OAI21X1 OAI21X1_60 ( .gnd(gnd), .vdd(vdd), .A(vdd), .B(_145_), .C(_146_), .Y(_137__3_) );
INVX1 INVX1_69 ( .gnd(gnd), .vdd(vdd), .A(asr1_cables_8__4_), .Y(_147_) );
NAND2X1 NAND2X1_61 ( .gnd(gnd), .vdd(vdd), .A(vdd), .B(asr1_cables_7__4_), .Y(_148_) );
OAI21X1 OAI21X1_61 ( .gnd(gnd), .vdd(vdd), .A(vdd), .B(_147_), .C(_148_), .Y(_137__4_) );
INVX1 INVX1_70 ( .gnd(gnd), .vdd(vdd), .A(asr1_cables_8__5_), .Y(_149_) );
NAND2X1 NAND2X1_62 ( .gnd(gnd), .vdd(vdd), .A(vdd), .B(asr1_cables_7__5_), .Y(_150_) );
OAI21X1 OAI21X1_62 ( .gnd(gnd), .vdd(vdd), .A(vdd), .B(_149_), .C(_150_), .Y(_137__5_) );
INVX1 INVX1_71 ( .gnd(gnd), .vdd(vdd), .A(asr1_cables_8__6_), .Y(_151_) );
NAND2X1 NAND2X1_63 ( .gnd(gnd), .vdd(vdd), .A(vdd), .B(asr1_cables_7__6_), .Y(_152_) );
OAI21X1 OAI21X1_63 ( .gnd(gnd), .vdd(vdd), .A(vdd), .B(_151_), .C(_152_), .Y(_137__6_) );
INVX1 INVX1_72 ( .gnd(gnd), .vdd(vdd), .A(asr1_cables_8__7_), .Y(_153_) );
NAND2X1 NAND2X1_64 ( .gnd(gnd), .vdd(vdd), .A(vdd), .B(asr1_cables_7__7_), .Y(_154_) );
OAI21X1 OAI21X1_64 ( .gnd(gnd), .vdd(vdd), .A(vdd), .B(_153_), .C(_154_), .Y(_137__7_) );
INVX1 INVX1_73 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf5), .Y(_138_) );
DFFSR DFFSR_57 ( .gnd(gnd), .vdd(vdd), .CLK(asr1_clk_bF_buf6), .D(_137__0_), .Q(asr1_cables_8__0_), .R(_138_), .S(vdd) );
DFFSR DFFSR_58 ( .gnd(gnd), .vdd(vdd), .CLK(asr1_clk_bF_buf1), .D(_137__1_), .Q(asr1_cables_8__1_), .R(_138_), .S(vdd) );
DFFSR DFFSR_59 ( .gnd(gnd), .vdd(vdd), .CLK(asr1_clk_bF_buf4), .D(_137__2_), .Q(asr1_cables_8__2_), .R(_138_), .S(vdd) );
DFFSR DFFSR_60 ( .gnd(gnd), .vdd(vdd), .CLK(asr1_clk_bF_buf6), .D(_137__3_), .Q(asr1_cables_8__3_), .R(_138_), .S(vdd) );
DFFSR DFFSR_61 ( .gnd(gnd), .vdd(vdd), .CLK(asr1_clk_bF_buf5), .D(_137__4_), .Q(asr1_cables_8__4_), .R(_138_), .S(vdd) );
DFFSR DFFSR_62 ( .gnd(gnd), .vdd(vdd), .CLK(asr1_clk_bF_buf1), .D(_137__5_), .Q(asr1_cables_8__5_), .R(_138_), .S(vdd) );
DFFSR DFFSR_63 ( .gnd(gnd), .vdd(vdd), .CLK(asr1_clk_bF_buf6), .D(_137__6_), .Q(asr1_cables_8__6_), .R(_138_), .S(vdd) );
DFFSR DFFSR_64 ( .gnd(gnd), .vdd(vdd), .CLK(asr1_clk_bF_buf5), .D(_137__7_), .Q(asr1_cables_8__7_), .R(_138_), .S(vdd) );
INVX1 INVX1_74 ( .gnd(gnd), .vdd(vdd), .A(asr2_cables_1__0_), .Y(_157_) );
NAND2X1 NAND2X1_65 ( .gnd(gnd), .vdd(vdd), .A(asr1_q_0_), .B(asr2_en_bF_buf5), .Y(_158_) );
OAI21X1 OAI21X1_65 ( .gnd(gnd), .vdd(vdd), .A(asr2_en_bF_buf5), .B(_157_), .C(_158_), .Y(_155__0_) );
INVX1 INVX1_75 ( .gnd(gnd), .vdd(vdd), .A(asr2_cables_1__1_), .Y(_159_) );
NAND2X1 NAND2X1_66 ( .gnd(gnd), .vdd(vdd), .A(asr2_en_bF_buf2), .B(asr1_q_1_), .Y(_160_) );
OAI21X1 OAI21X1_66 ( .gnd(gnd), .vdd(vdd), .A(asr2_en_bF_buf2), .B(_159_), .C(_160_), .Y(_155__1_) );
INVX1 INVX1_76 ( .gnd(gnd), .vdd(vdd), .A(asr2_cables_1__2_), .Y(_161_) );
NAND2X1 NAND2X1_67 ( .gnd(gnd), .vdd(vdd), .A(asr2_en_bF_buf2), .B(asr1_q_2_), .Y(_162_) );
OAI21X1 OAI21X1_67 ( .gnd(gnd), .vdd(vdd), .A(asr2_en_bF_buf2), .B(_161_), .C(_162_), .Y(_155__2_) );
INVX1 INVX1_77 ( .gnd(gnd), .vdd(vdd), .A(asr2_cables_1__3_), .Y(_163_) );
NAND2X1 NAND2X1_68 ( .gnd(gnd), .vdd(vdd), .A(asr2_en_bF_buf5), .B(asr1_q_3_), .Y(_164_) );
OAI21X1 OAI21X1_68 ( .gnd(gnd), .vdd(vdd), .A(asr2_en_bF_buf5), .B(_163_), .C(_164_), .Y(_155__3_) );
INVX1 INVX1_78 ( .gnd(gnd), .vdd(vdd), .A(asr2_cables_1__4_), .Y(_165_) );
NAND2X1 NAND2X1_69 ( .gnd(gnd), .vdd(vdd), .A(asr2_en_bF_buf5), .B(asr1_q_4_), .Y(_166_) );
OAI21X1 OAI21X1_69 ( .gnd(gnd), .vdd(vdd), .A(asr2_en_bF_buf5), .B(_165_), .C(_166_), .Y(_155__4_) );
INVX1 INVX1_79 ( .gnd(gnd), .vdd(vdd), .A(asr2_cables_1__5_), .Y(_167_) );
NAND2X1 NAND2X1_70 ( .gnd(gnd), .vdd(vdd), .A(asr2_en_bF_buf2), .B(asr1_q_5_), .Y(_168_) );
OAI21X1 OAI21X1_70 ( .gnd(gnd), .vdd(vdd), .A(asr2_en_bF_buf2), .B(_167_), .C(_168_), .Y(_155__5_) );
INVX1 INVX1_80 ( .gnd(gnd), .vdd(vdd), .A(asr2_cables_1__6_), .Y(_169_) );
NAND2X1 NAND2X1_71 ( .gnd(gnd), .vdd(vdd), .A(asr2_en_bF_buf5), .B(asr1_q_6_), .Y(_170_) );
OAI21X1 OAI21X1_71 ( .gnd(gnd), .vdd(vdd), .A(asr2_en_bF_buf5), .B(_169_), .C(_170_), .Y(_155__6_) );
INVX1 INVX1_81 ( .gnd(gnd), .vdd(vdd), .A(asr2_cables_1__7_), .Y(_171_) );
NAND2X1 NAND2X1_72 ( .gnd(gnd), .vdd(vdd), .A(asr2_en_bF_buf2), .B(asr1_q_7_), .Y(_172_) );
OAI21X1 OAI21X1_72 ( .gnd(gnd), .vdd(vdd), .A(asr2_en_bF_buf2), .B(_171_), .C(_172_), .Y(_155__7_) );
INVX1 INVX1_82 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf5), .Y(_156_) );
DFFSR DFFSR_65 ( .gnd(gnd), .vdd(vdd), .CLK(asr2_clk_bF_buf7), .D(_155__0_), .Q(asr2_cables_1__0_), .R(_156_), .S(vdd) );
DFFSR DFFSR_66 ( .gnd(gnd), .vdd(vdd), .CLK(asr2_clk_bF_buf4), .D(_155__1_), .Q(asr2_cables_1__1_), .R(_156_), .S(vdd) );
DFFSR DFFSR_67 ( .gnd(gnd), .vdd(vdd), .CLK(asr2_clk_bF_buf4), .D(_155__2_), .Q(asr2_cables_1__2_), .R(_156_), .S(vdd) );
DFFSR DFFSR_68 ( .gnd(gnd), .vdd(vdd), .CLK(asr2_clk_bF_buf7), .D(_155__3_), .Q(asr2_cables_1__3_), .R(_156_), .S(vdd) );
DFFSR DFFSR_69 ( .gnd(gnd), .vdd(vdd), .CLK(asr2_clk_bF_buf7), .D(_155__4_), .Q(asr2_cables_1__4_), .R(_156_), .S(vdd) );
DFFSR DFFSR_70 ( .gnd(gnd), .vdd(vdd), .CLK(asr2_clk_bF_buf4), .D(_155__5_), .Q(asr2_cables_1__5_), .R(_156_), .S(vdd) );
DFFSR DFFSR_71 ( .gnd(gnd), .vdd(vdd), .CLK(asr2_clk_bF_buf7), .D(_155__6_), .Q(asr2_cables_1__6_), .R(_156_), .S(vdd) );
DFFSR DFFSR_72 ( .gnd(gnd), .vdd(vdd), .CLK(asr2_clk_bF_buf4), .D(_155__7_), .Q(asr2_cables_1__7_), .R(_156_), .S(vdd) );
INVX1 INVX1_83 ( .gnd(gnd), .vdd(vdd), .A(asr2_cables_2__0_), .Y(_175_) );
NAND2X1 NAND2X1_73 ( .gnd(gnd), .vdd(vdd), .A(asr2_cables_1__0_), .B(asr2_en_bF_buf4), .Y(_176_) );
OAI21X1 OAI21X1_73 ( .gnd(gnd), .vdd(vdd), .A(asr2_en_bF_buf4), .B(_175_), .C(_176_), .Y(_173__0_) );
INVX1 INVX1_84 ( .gnd(gnd), .vdd(vdd), .A(asr2_cables_2__1_), .Y(_177_) );
NAND2X1 NAND2X1_74 ( .gnd(gnd), .vdd(vdd), .A(asr2_en_bF_buf2), .B(asr2_cables_1__1_), .Y(_178_) );
OAI21X1 OAI21X1_74 ( .gnd(gnd), .vdd(vdd), .A(asr2_en_bF_buf5), .B(_177_), .C(_178_), .Y(_173__1_) );
INVX1 INVX1_85 ( .gnd(gnd), .vdd(vdd), .A(asr2_cables_2__2_), .Y(_179_) );
NAND2X1 NAND2X1_75 ( .gnd(gnd), .vdd(vdd), .A(asr2_en_bF_buf8), .B(asr2_cables_1__2_), .Y(_180_) );
OAI21X1 OAI21X1_75 ( .gnd(gnd), .vdd(vdd), .A(asr2_en_bF_buf8), .B(_179_), .C(_180_), .Y(_173__2_) );
INVX1 INVX1_86 ( .gnd(gnd), .vdd(vdd), .A(asr2_cables_2__3_), .Y(_181_) );
NAND2X1 NAND2X1_76 ( .gnd(gnd), .vdd(vdd), .A(asr2_en_bF_buf4), .B(asr2_cables_1__3_), .Y(_182_) );
OAI21X1 OAI21X1_76 ( .gnd(gnd), .vdd(vdd), .A(asr2_en_bF_buf4), .B(_181_), .C(_182_), .Y(_173__3_) );
INVX1 INVX1_87 ( .gnd(gnd), .vdd(vdd), .A(asr2_cables_2__4_), .Y(_183_) );
NAND2X1 NAND2X1_77 ( .gnd(gnd), .vdd(vdd), .A(asr2_en_bF_buf10), .B(asr2_cables_1__4_), .Y(_184_) );
OAI21X1 OAI21X1_77 ( .gnd(gnd), .vdd(vdd), .A(asr2_en_bF_buf10), .B(_183_), .C(_184_), .Y(_173__4_) );
INVX1 INVX1_88 ( .gnd(gnd), .vdd(vdd), .A(asr2_cables_2__5_), .Y(_185_) );
NAND2X1 NAND2X1_78 ( .gnd(gnd), .vdd(vdd), .A(asr2_en_bF_buf2), .B(asr2_cables_1__5_), .Y(_186_) );
OAI21X1 OAI21X1_78 ( .gnd(gnd), .vdd(vdd), .A(asr2_en_bF_buf2), .B(_185_), .C(_186_), .Y(_173__5_) );
INVX1 INVX1_89 ( .gnd(gnd), .vdd(vdd), .A(asr2_cables_2__6_), .Y(_187_) );
NAND2X1 NAND2X1_79 ( .gnd(gnd), .vdd(vdd), .A(asr2_en_bF_buf4), .B(asr2_cables_1__6_), .Y(_188_) );
OAI21X1 OAI21X1_79 ( .gnd(gnd), .vdd(vdd), .A(asr2_en_bF_buf4), .B(_187_), .C(_188_), .Y(_173__6_) );
INVX1 INVX1_90 ( .gnd(gnd), .vdd(vdd), .A(asr2_cables_2__7_), .Y(_189_) );
NAND2X1 NAND2X1_80 ( .gnd(gnd), .vdd(vdd), .A(asr2_en_bF_buf5), .B(asr2_cables_1__7_), .Y(_190_) );
OAI21X1 OAI21X1_80 ( .gnd(gnd), .vdd(vdd), .A(asr2_en_bF_buf5), .B(_189_), .C(_190_), .Y(_173__7_) );
INVX1 INVX1_91 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf3), .Y(_174_) );
DFFSR DFFSR_73 ( .gnd(gnd), .vdd(vdd), .CLK(asr2_clk_bF_buf7), .D(_173__0_), .Q(asr2_cables_2__0_), .R(_174_), .S(vdd) );
DFFSR DFFSR_74 ( .gnd(gnd), .vdd(vdd), .CLK(asr2_clk_bF_buf4), .D(_173__1_), .Q(asr2_cables_2__1_), .R(_174_), .S(vdd) );
DFFSR DFFSR_75 ( .gnd(gnd), .vdd(vdd), .CLK(asr2_clk_bF_buf5), .D(_173__2_), .Q(asr2_cables_2__2_), .R(_174_), .S(vdd) );
DFFSR DFFSR_76 ( .gnd(gnd), .vdd(vdd), .CLK(asr2_clk_bF_buf0), .D(_173__3_), .Q(asr2_cables_2__3_), .R(_174_), .S(vdd) );
DFFSR DFFSR_77 ( .gnd(gnd), .vdd(vdd), .CLK(asr2_clk_bF_buf0), .D(_173__4_), .Q(asr2_cables_2__4_), .R(_174_), .S(vdd) );
DFFSR DFFSR_78 ( .gnd(gnd), .vdd(vdd), .CLK(asr2_clk_bF_buf4), .D(_173__5_), .Q(asr2_cables_2__5_), .R(_174_), .S(vdd) );
DFFSR DFFSR_79 ( .gnd(gnd), .vdd(vdd), .CLK(asr2_clk_bF_buf7), .D(_173__6_), .Q(asr2_cables_2__6_), .R(_174_), .S(vdd) );
DFFSR DFFSR_80 ( .gnd(gnd), .vdd(vdd), .CLK(asr2_clk_bF_buf4), .D(_173__7_), .Q(asr2_cables_2__7_), .R(_174_), .S(vdd) );
INVX1 INVX1_92 ( .gnd(gnd), .vdd(vdd), .A(asr2_cables_3__0_), .Y(_193_) );
NAND2X1 NAND2X1_81 ( .gnd(gnd), .vdd(vdd), .A(asr2_cables_2__0_), .B(asr2_en_bF_buf4), .Y(_194_) );
OAI21X1 OAI21X1_81 ( .gnd(gnd), .vdd(vdd), .A(asr2_en_bF_buf4), .B(_193_), .C(_194_), .Y(_191__0_) );
INVX1 INVX1_93 ( .gnd(gnd), .vdd(vdd), .A(asr2_cables_3__1_), .Y(_195_) );
NAND2X1 NAND2X1_82 ( .gnd(gnd), .vdd(vdd), .A(asr2_en_bF_buf10), .B(asr2_cables_2__1_), .Y(_196_) );
OAI21X1 OAI21X1_82 ( .gnd(gnd), .vdd(vdd), .A(asr2_en_bF_buf10), .B(_195_), .C(_196_), .Y(_191__1_) );
INVX1 INVX1_94 ( .gnd(gnd), .vdd(vdd), .A(asr2_cables_3__2_), .Y(_197_) );
NAND2X1 NAND2X1_83 ( .gnd(gnd), .vdd(vdd), .A(asr2_en_bF_buf9), .B(asr2_cables_2__2_), .Y(_198_) );
OAI21X1 OAI21X1_83 ( .gnd(gnd), .vdd(vdd), .A(asr2_en_bF_buf0), .B(_197_), .C(_198_), .Y(_191__2_) );
INVX1 INVX1_95 ( .gnd(gnd), .vdd(vdd), .A(asr2_cables_3__3_), .Y(_199_) );
NAND2X1 NAND2X1_84 ( .gnd(gnd), .vdd(vdd), .A(asr2_en_bF_buf4), .B(asr2_cables_2__3_), .Y(_200_) );
OAI21X1 OAI21X1_84 ( .gnd(gnd), .vdd(vdd), .A(asr2_en_bF_buf4), .B(_199_), .C(_200_), .Y(_191__3_) );
INVX1 INVX1_96 ( .gnd(gnd), .vdd(vdd), .A(asr2_cables_3__4_), .Y(_201_) );
NAND2X1 NAND2X1_85 ( .gnd(gnd), .vdd(vdd), .A(asr2_en_bF_buf10), .B(asr2_cables_2__4_), .Y(_202_) );
OAI21X1 OAI21X1_85 ( .gnd(gnd), .vdd(vdd), .A(asr2_en_bF_buf6), .B(_201_), .C(_202_), .Y(_191__4_) );
INVX1 INVX1_97 ( .gnd(gnd), .vdd(vdd), .A(asr2_cables_3__5_), .Y(_203_) );
NAND2X1 NAND2X1_86 ( .gnd(gnd), .vdd(vdd), .A(asr2_en_bF_buf3), .B(asr2_cables_2__5_), .Y(_204_) );
OAI21X1 OAI21X1_86 ( .gnd(gnd), .vdd(vdd), .A(asr2_en_bF_buf3), .B(_203_), .C(_204_), .Y(_191__5_) );
INVX1 INVX1_98 ( .gnd(gnd), .vdd(vdd), .A(asr2_cables_3__6_), .Y(_205_) );
NAND2X1 NAND2X1_87 ( .gnd(gnd), .vdd(vdd), .A(asr2_en_bF_buf10), .B(asr2_cables_2__6_), .Y(_206_) );
OAI21X1 OAI21X1_87 ( .gnd(gnd), .vdd(vdd), .A(asr2_en_bF_buf10), .B(_205_), .C(_206_), .Y(_191__6_) );
INVX1 INVX1_99 ( .gnd(gnd), .vdd(vdd), .A(asr2_cables_3__7_), .Y(_207_) );
NAND2X1 NAND2X1_88 ( .gnd(gnd), .vdd(vdd), .A(asr2_en_bF_buf5), .B(asr2_cables_2__7_), .Y(_208_) );
OAI21X1 OAI21X1_88 ( .gnd(gnd), .vdd(vdd), .A(asr2_en_bF_buf4), .B(_207_), .C(_208_), .Y(_191__7_) );
INVX1 INVX1_100 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf5), .Y(_192_) );
DFFSR DFFSR_81 ( .gnd(gnd), .vdd(vdd), .CLK(asr2_clk_bF_buf7), .D(_191__0_), .Q(asr2_cables_3__0_), .R(_192_), .S(vdd) );
DFFSR DFFSR_82 ( .gnd(gnd), .vdd(vdd), .CLK(asr2_clk_bF_buf0), .D(_191__1_), .Q(asr2_cables_3__1_), .R(_192_), .S(vdd) );
DFFSR DFFSR_83 ( .gnd(gnd), .vdd(vdd), .CLK(asr2_clk_bF_buf6), .D(_191__2_), .Q(asr2_cables_3__2_), .R(_192_), .S(vdd) );
DFFSR DFFSR_84 ( .gnd(gnd), .vdd(vdd), .CLK(asr2_clk_bF_buf7), .D(_191__3_), .Q(asr2_cables_3__3_), .R(_192_), .S(vdd) );
DFFSR DFFSR_85 ( .gnd(gnd), .vdd(vdd), .CLK(asr2_clk_bF_buf6), .D(_191__4_), .Q(asr2_cables_3__4_), .R(_192_), .S(vdd) );
DFFSR DFFSR_86 ( .gnd(gnd), .vdd(vdd), .CLK(asr2_clk_bF_buf3), .D(_191__5_), .Q(asr2_cables_3__5_), .R(_192_), .S(vdd) );
DFFSR DFFSR_87 ( .gnd(gnd), .vdd(vdd), .CLK(asr2_clk_bF_buf0), .D(_191__6_), .Q(asr2_cables_3__6_), .R(_192_), .S(vdd) );
DFFSR DFFSR_88 ( .gnd(gnd), .vdd(vdd), .CLK(asr2_clk_bF_buf7), .D(_191__7_), .Q(asr2_cables_3__7_), .R(_192_), .S(vdd) );
INVX1 INVX1_101 ( .gnd(gnd), .vdd(vdd), .A(asr2_cables_4_), .Y(_211_) );
NAND2X1 NAND2X1_89 ( .gnd(gnd), .vdd(vdd), .A(asr2_cables_3__0_), .B(asr2_en_bF_buf4), .Y(_212_) );
OAI21X1 OAI21X1_89 ( .gnd(gnd), .vdd(vdd), .A(asr2_en_bF_buf10), .B(_211_), .C(_212_), .Y(_209__0_) );
INVX1 INVX1_102 ( .gnd(gnd), .vdd(vdd), .A(_227_), .Y(_213_) );
NAND2X1 NAND2X1_90 ( .gnd(gnd), .vdd(vdd), .A(asr2_en_bF_buf10), .B(asr2_cables_3__1_), .Y(_214_) );
OAI21X1 OAI21X1_90 ( .gnd(gnd), .vdd(vdd), .A(asr2_en_bF_buf8), .B(_213_), .C(_214_), .Y(_209__1_) );
INVX1 INVX1_103 ( .gnd(gnd), .vdd(vdd), .A(_233_), .Y(_215_) );
NAND2X1 NAND2X1_91 ( .gnd(gnd), .vdd(vdd), .A(asr2_en_bF_buf7), .B(asr2_cables_3__2_), .Y(_216_) );
OAI21X1 OAI21X1_91 ( .gnd(gnd), .vdd(vdd), .A(asr2_en_bF_buf7), .B(_215_), .C(_216_), .Y(_209__2_) );
INVX1 INVX1_104 ( .gnd(gnd), .vdd(vdd), .A(_228_), .Y(_217_) );
NAND2X1 NAND2X1_92 ( .gnd(gnd), .vdd(vdd), .A(asr2_en_bF_buf9), .B(asr2_cables_3__3_), .Y(_218_) );
OAI21X1 OAI21X1_92 ( .gnd(gnd), .vdd(vdd), .A(asr2_en_bF_buf3), .B(_217_), .C(_218_), .Y(_209__3_) );
INVX1 INVX1_105 ( .gnd(gnd), .vdd(vdd), .A(_229_), .Y(_219_) );
NAND2X1 NAND2X1_93 ( .gnd(gnd), .vdd(vdd), .A(asr2_en_bF_buf7), .B(asr2_cables_3__4_), .Y(_220_) );
OAI21X1 OAI21X1_93 ( .gnd(gnd), .vdd(vdd), .A(asr2_en_bF_buf7), .B(_219_), .C(_220_), .Y(_209__4_) );
INVX1 INVX1_106 ( .gnd(gnd), .vdd(vdd), .A(_230_), .Y(_221_) );
NAND2X1 NAND2X1_94 ( .gnd(gnd), .vdd(vdd), .A(asr2_en_bF_buf1), .B(asr2_cables_3__5_), .Y(_222_) );
OAI21X1 OAI21X1_94 ( .gnd(gnd), .vdd(vdd), .A(asr2_en_bF_buf1), .B(_221_), .C(_222_), .Y(_209__5_) );
INVX1 INVX1_107 ( .gnd(gnd), .vdd(vdd), .A(_231_), .Y(_223_) );
NAND2X1 NAND2X1_95 ( .gnd(gnd), .vdd(vdd), .A(asr2_en_bF_buf6), .B(asr2_cables_3__6_), .Y(_224_) );
OAI21X1 OAI21X1_95 ( .gnd(gnd), .vdd(vdd), .A(asr2_en_bF_buf7), .B(_223_), .C(_224_), .Y(_209__6_) );
INVX1 INVX1_108 ( .gnd(gnd), .vdd(vdd), .A(_232_), .Y(_225_) );
NAND2X1 NAND2X1_96 ( .gnd(gnd), .vdd(vdd), .A(asr2_en_bF_buf10), .B(asr2_cables_3__7_), .Y(_226_) );
OAI21X1 OAI21X1_96 ( .gnd(gnd), .vdd(vdd), .A(asr2_en_bF_buf9), .B(_225_), .C(_226_), .Y(_209__7_) );
INVX1 INVX1_109 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf3), .Y(_210_) );
DFFSR DFFSR_89 ( .gnd(gnd), .vdd(vdd), .CLK(asr2_clk_bF_buf0), .D(_209__0_), .Q(asr2_cables_4_), .R(_210_), .S(vdd) );
DFFSR DFFSR_90 ( .gnd(gnd), .vdd(vdd), .CLK(asr2_clk_bF_buf5), .D(_209__1_), .Q(_227_), .R(_210_), .S(vdd) );
DFFSR DFFSR_91 ( .gnd(gnd), .vdd(vdd), .CLK(asr2_clk_bF_buf1), .D(_209__2_), .Q(_233_), .R(_210_), .S(vdd) );
DFFSR DFFSR_92 ( .gnd(gnd), .vdd(vdd), .CLK(asr2_clk_bF_buf3), .D(_209__3_), .Q(_228_), .R(_210_), .S(vdd) );
DFFSR DFFSR_93 ( .gnd(gnd), .vdd(vdd), .CLK(asr2_clk_bF_buf1), .D(_209__4_), .Q(_229_), .R(_210_), .S(vdd) );
DFFSR DFFSR_94 ( .gnd(gnd), .vdd(vdd), .CLK(asr2_clk_bF_buf2), .D(_209__5_), .Q(_230_), .R(_210_), .S(vdd) );
DFFSR DFFSR_95 ( .gnd(gnd), .vdd(vdd), .CLK(asr2_clk_bF_buf1), .D(_209__6_), .Q(_231_), .R(_210_), .S(vdd) );
DFFSR DFFSR_96 ( .gnd(gnd), .vdd(vdd), .CLK(asr2_clk_bF_buf6), .D(_209__7_), .Q(_232_), .R(_210_), .S(vdd) );
INVX1 INVX1_110 ( .gnd(gnd), .vdd(vdd), .A(asr2_cables_5__0_), .Y(_236_) );
NAND2X1 NAND2X1_97 ( .gnd(gnd), .vdd(vdd), .A(asr2_cables_4_), .B(asr2_en_bF_buf6), .Y(_237_) );
OAI21X1 OAI21X1_97 ( .gnd(gnd), .vdd(vdd), .A(asr2_en_bF_buf6), .B(_236_), .C(_237_), .Y(_234__0_) );
INVX1 INVX1_111 ( .gnd(gnd), .vdd(vdd), .A(asr2_cables_5__1_), .Y(_238_) );
NAND2X1 NAND2X1_98 ( .gnd(gnd), .vdd(vdd), .A(asr2_en_bF_buf0), .B(_227_), .Y(_239_) );
OAI21X1 OAI21X1_98 ( .gnd(gnd), .vdd(vdd), .A(asr2_en_bF_buf0), .B(_238_), .C(_239_), .Y(_234__1_) );
INVX1 INVX1_112 ( .gnd(gnd), .vdd(vdd), .A(asr2_cables_5__2_), .Y(_240_) );
NAND2X1 NAND2X1_99 ( .gnd(gnd), .vdd(vdd), .A(asr2_en_bF_buf1), .B(_233_), .Y(_241_) );
OAI21X1 OAI21X1_99 ( .gnd(gnd), .vdd(vdd), .A(asr2_en_bF_buf1), .B(_240_), .C(_241_), .Y(_234__2_) );
INVX1 INVX1_113 ( .gnd(gnd), .vdd(vdd), .A(asr2_cables_5__3_), .Y(_242_) );
NAND2X1 NAND2X1_100 ( .gnd(gnd), .vdd(vdd), .A(asr2_en_bF_buf8), .B(_228_), .Y(_243_) );
OAI21X1 OAI21X1_100 ( .gnd(gnd), .vdd(vdd), .A(asr2_en_bF_buf8), .B(_242_), .C(_243_), .Y(_234__3_) );
INVX1 INVX1_114 ( .gnd(gnd), .vdd(vdd), .A(asr2_cables_5__4_), .Y(_244_) );
NAND2X1 NAND2X1_101 ( .gnd(gnd), .vdd(vdd), .A(asr2_en_bF_buf9), .B(_229_), .Y(_245_) );
OAI21X1 OAI21X1_101 ( .gnd(gnd), .vdd(vdd), .A(asr2_en_bF_buf9), .B(_244_), .C(_245_), .Y(_234__4_) );
INVX1 INVX1_115 ( .gnd(gnd), .vdd(vdd), .A(asr2_cables_5__5_), .Y(_246_) );
NAND2X1 NAND2X1_102 ( .gnd(gnd), .vdd(vdd), .A(asr2_en_bF_buf1), .B(_230_), .Y(_247_) );
OAI21X1 OAI21X1_102 ( .gnd(gnd), .vdd(vdd), .A(asr2_en_bF_buf1), .B(_246_), .C(_247_), .Y(_234__5_) );
INVX1 INVX1_116 ( .gnd(gnd), .vdd(vdd), .A(asr2_cables_5__6_), .Y(_248_) );
NAND2X1 NAND2X1_103 ( .gnd(gnd), .vdd(vdd), .A(asr2_en_bF_buf6), .B(_231_), .Y(_249_) );
OAI21X1 OAI21X1_103 ( .gnd(gnd), .vdd(vdd), .A(asr2_en_bF_buf6), .B(_248_), .C(_249_), .Y(_234__6_) );
INVX1 INVX1_117 ( .gnd(gnd), .vdd(vdd), .A(asr2_cables_5__7_), .Y(_250_) );
NAND2X1 NAND2X1_104 ( .gnd(gnd), .vdd(vdd), .A(asr2_en_bF_buf9), .B(_232_), .Y(_251_) );
OAI21X1 OAI21X1_104 ( .gnd(gnd), .vdd(vdd), .A(asr2_en_bF_buf1), .B(_250_), .C(_251_), .Y(_234__7_) );
INVX1 INVX1_118 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf3), .Y(_235_) );
DFFSR DFFSR_97 ( .gnd(gnd), .vdd(vdd), .CLK(asr2_clk_bF_buf6), .D(_234__0_), .Q(asr2_cables_5__0_), .R(_235_), .S(vdd) );
DFFSR DFFSR_98 ( .gnd(gnd), .vdd(vdd), .CLK(asr2_clk_bF_buf5), .D(_234__1_), .Q(asr2_cables_5__1_), .R(_235_), .S(vdd) );
DFFSR DFFSR_99 ( .gnd(gnd), .vdd(vdd), .CLK(asr2_clk_bF_buf2), .D(_234__2_), .Q(asr2_cables_5__2_), .R(_235_), .S(vdd) );
DFFSR DFFSR_100 ( .gnd(gnd), .vdd(vdd), .CLK(asr2_clk_bF_buf5), .D(_234__3_), .Q(asr2_cables_5__3_), .R(_235_), .S(vdd) );
DFFSR DFFSR_101 ( .gnd(gnd), .vdd(vdd), .CLK(asr2_clk_bF_buf2), .D(_234__4_), .Q(asr2_cables_5__4_), .R(_235_), .S(vdd) );
DFFSR DFFSR_102 ( .gnd(gnd), .vdd(vdd), .CLK(asr2_clk_bF_buf2), .D(_234__5_), .Q(asr2_cables_5__5_), .R(_235_), .S(vdd) );
DFFSR DFFSR_103 ( .gnd(gnd), .vdd(vdd), .CLK(asr2_clk_bF_buf1), .D(_234__6_), .Q(asr2_cables_5__6_), .R(_235_), .S(vdd) );
DFFSR DFFSR_104 ( .gnd(gnd), .vdd(vdd), .CLK(asr2_clk_bF_buf2), .D(_234__7_), .Q(asr2_cables_5__7_), .R(_235_), .S(vdd) );
INVX1 INVX1_119 ( .gnd(gnd), .vdd(vdd), .A(asr2_cables_6__0_), .Y(_254_) );
NAND2X1 NAND2X1_105 ( .gnd(gnd), .vdd(vdd), .A(asr2_cables_5__0_), .B(asr2_en_bF_buf0), .Y(_255_) );
OAI21X1 OAI21X1_105 ( .gnd(gnd), .vdd(vdd), .A(asr2_en_bF_buf0), .B(_254_), .C(_255_), .Y(_252__0_) );
INVX1 INVX1_120 ( .gnd(gnd), .vdd(vdd), .A(asr2_cables_6__1_), .Y(_256_) );
NAND2X1 NAND2X1_106 ( .gnd(gnd), .vdd(vdd), .A(asr2_en_bF_buf0), .B(asr2_cables_5__1_), .Y(_257_) );
OAI21X1 OAI21X1_106 ( .gnd(gnd), .vdd(vdd), .A(asr2_en_bF_buf8), .B(_256_), .C(_257_), .Y(_252__1_) );
INVX1 INVX1_121 ( .gnd(gnd), .vdd(vdd), .A(asr2_cables_6__2_), .Y(_258_) );
NAND2X1 NAND2X1_107 ( .gnd(gnd), .vdd(vdd), .A(asr2_en_bF_buf9), .B(asr2_cables_5__2_), .Y(_259_) );
OAI21X1 OAI21X1_107 ( .gnd(gnd), .vdd(vdd), .A(asr2_en_bF_buf9), .B(_258_), .C(_259_), .Y(_252__2_) );
INVX1 INVX1_122 ( .gnd(gnd), .vdd(vdd), .A(asr2_cables_6__3_), .Y(_260_) );
NAND2X1 NAND2X1_108 ( .gnd(gnd), .vdd(vdd), .A(asr2_en_bF_buf3), .B(asr2_cables_5__3_), .Y(_261_) );
OAI21X1 OAI21X1_108 ( .gnd(gnd), .vdd(vdd), .A(asr2_en_bF_buf3), .B(_260_), .C(_261_), .Y(_252__3_) );
INVX1 INVX1_123 ( .gnd(gnd), .vdd(vdd), .A(asr2_cables_6__4_), .Y(_262_) );
NAND2X1 NAND2X1_109 ( .gnd(gnd), .vdd(vdd), .A(asr2_en_bF_buf7), .B(asr2_cables_5__4_), .Y(_263_) );
OAI21X1 OAI21X1_109 ( .gnd(gnd), .vdd(vdd), .A(asr2_en_bF_buf7), .B(_262_), .C(_263_), .Y(_252__4_) );
INVX1 INVX1_124 ( .gnd(gnd), .vdd(vdd), .A(asr2_cables_6__5_), .Y(_264_) );
NAND2X1 NAND2X1_110 ( .gnd(gnd), .vdd(vdd), .A(asr2_en_bF_buf1), .B(asr2_cables_5__5_), .Y(_265_) );
OAI21X1 OAI21X1_110 ( .gnd(gnd), .vdd(vdd), .A(asr2_en_bF_buf1), .B(_264_), .C(_265_), .Y(_252__5_) );
INVX1 INVX1_125 ( .gnd(gnd), .vdd(vdd), .A(asr2_cables_6__6_), .Y(_266_) );
NAND2X1 NAND2X1_111 ( .gnd(gnd), .vdd(vdd), .A(asr2_en_bF_buf6), .B(asr2_cables_5__6_), .Y(_267_) );
OAI21X1 OAI21X1_111 ( .gnd(gnd), .vdd(vdd), .A(asr2_en_bF_buf6), .B(_266_), .C(_267_), .Y(_252__6_) );
INVX1 INVX1_126 ( .gnd(gnd), .vdd(vdd), .A(asr2_cables_6__7_), .Y(_268_) );
NAND2X1 NAND2X1_112 ( .gnd(gnd), .vdd(vdd), .A(asr2_en_bF_buf9), .B(asr2_cables_5__7_), .Y(_269_) );
OAI21X1 OAI21X1_112 ( .gnd(gnd), .vdd(vdd), .A(asr2_en_bF_buf7), .B(_268_), .C(_269_), .Y(_252__7_) );
INVX1 INVX1_127 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf3), .Y(_253_) );
DFFSR DFFSR_105 ( .gnd(gnd), .vdd(vdd), .CLK(asr2_clk_bF_buf5), .D(_252__0_), .Q(asr2_cables_6__0_), .R(_253_), .S(vdd) );
DFFSR DFFSR_106 ( .gnd(gnd), .vdd(vdd), .CLK(asr2_clk_bF_buf5), .D(_252__1_), .Q(asr2_cables_6__1_), .R(_253_), .S(vdd) );
DFFSR DFFSR_107 ( .gnd(gnd), .vdd(vdd), .CLK(asr2_clk_bF_buf2), .D(_252__2_), .Q(asr2_cables_6__2_), .R(_253_), .S(vdd) );
DFFSR DFFSR_108 ( .gnd(gnd), .vdd(vdd), .CLK(asr2_clk_bF_buf3), .D(_252__3_), .Q(asr2_cables_6__3_), .R(_253_), .S(vdd) );
DFFSR DFFSR_109 ( .gnd(gnd), .vdd(vdd), .CLK(asr2_clk_bF_buf1), .D(_252__4_), .Q(asr2_cables_6__4_), .R(_253_), .S(vdd) );
DFFSR DFFSR_110 ( .gnd(gnd), .vdd(vdd), .CLK(asr2_clk_bF_buf2), .D(_252__5_), .Q(asr2_cables_6__5_), .R(_253_), .S(vdd) );
DFFSR DFFSR_111 ( .gnd(gnd), .vdd(vdd), .CLK(asr2_clk_bF_buf6), .D(_252__6_), .Q(asr2_cables_6__6_), .R(_253_), .S(vdd) );
DFFSR DFFSR_112 ( .gnd(gnd), .vdd(vdd), .CLK(asr2_clk_bF_buf1), .D(_252__7_), .Q(asr2_cables_6__7_), .R(_253_), .S(vdd) );
INVX1 INVX1_128 ( .gnd(gnd), .vdd(vdd), .A(asr2_cables_7__0_), .Y(_272_) );
NAND2X1 NAND2X1_113 ( .gnd(gnd), .vdd(vdd), .A(asr2_cables_6__0_), .B(asr2_en_bF_buf0), .Y(_273_) );
OAI21X1 OAI21X1_113 ( .gnd(gnd), .vdd(vdd), .A(asr2_en_bF_buf0), .B(_272_), .C(_273_), .Y(_270__0_) );
INVX1 INVX1_129 ( .gnd(gnd), .vdd(vdd), .A(asr2_cables_7__1_), .Y(_274_) );
NAND2X1 NAND2X1_114 ( .gnd(gnd), .vdd(vdd), .A(asr2_en_bF_buf8), .B(asr2_cables_6__1_), .Y(_275_) );
OAI21X1 OAI21X1_114 ( .gnd(gnd), .vdd(vdd), .A(asr2_en_bF_buf8), .B(_274_), .C(_275_), .Y(_270__1_) );
INVX1 INVX1_130 ( .gnd(gnd), .vdd(vdd), .A(asr2_cables_7__2_), .Y(_276_) );
NAND2X1 NAND2X1_115 ( .gnd(gnd), .vdd(vdd), .A(asr2_en_bF_buf9), .B(asr2_cables_6__2_), .Y(_277_) );
OAI21X1 OAI21X1_115 ( .gnd(gnd), .vdd(vdd), .A(asr2_en_bF_buf0), .B(_276_), .C(_277_), .Y(_270__2_) );
INVX1 INVX1_131 ( .gnd(gnd), .vdd(vdd), .A(asr2_cables_7__3_), .Y(_278_) );
NAND2X1 NAND2X1_116 ( .gnd(gnd), .vdd(vdd), .A(asr2_en_bF_buf3), .B(asr2_cables_6__3_), .Y(_279_) );
OAI21X1 OAI21X1_116 ( .gnd(gnd), .vdd(vdd), .A(asr2_en_bF_buf3), .B(_278_), .C(_279_), .Y(_270__3_) );
INVX1 INVX1_132 ( .gnd(gnd), .vdd(vdd), .A(asr2_cables_7__4_), .Y(_280_) );
NAND2X1 NAND2X1_117 ( .gnd(gnd), .vdd(vdd), .A(asr2_en_bF_buf7), .B(asr2_cables_6__4_), .Y(_281_) );
OAI21X1 OAI21X1_117 ( .gnd(gnd), .vdd(vdd), .A(asr2_en_bF_buf7), .B(_280_), .C(_281_), .Y(_270__4_) );
INVX1 INVX1_133 ( .gnd(gnd), .vdd(vdd), .A(asr2_cables_7__5_), .Y(_282_) );
NAND2X1 NAND2X1_118 ( .gnd(gnd), .vdd(vdd), .A(asr2_en_bF_buf3), .B(asr2_cables_6__5_), .Y(_283_) );
OAI21X1 OAI21X1_118 ( .gnd(gnd), .vdd(vdd), .A(asr2_en_bF_buf3), .B(_282_), .C(_283_), .Y(_270__5_) );
INVX1 INVX1_134 ( .gnd(gnd), .vdd(vdd), .A(asr2_cables_7__6_), .Y(_284_) );
NAND2X1 NAND2X1_119 ( .gnd(gnd), .vdd(vdd), .A(asr2_en_bF_buf6), .B(asr2_cables_6__6_), .Y(_285_) );
OAI21X1 OAI21X1_119 ( .gnd(gnd), .vdd(vdd), .A(asr2_en_bF_buf6), .B(_284_), .C(_285_), .Y(_270__6_) );
INVX1 INVX1_135 ( .gnd(gnd), .vdd(vdd), .A(asr2_cables_7__7_), .Y(_286_) );
NAND2X1 NAND2X1_120 ( .gnd(gnd), .vdd(vdd), .A(asr2_en_bF_buf9), .B(asr2_cables_6__7_), .Y(_287_) );
OAI21X1 OAI21X1_120 ( .gnd(gnd), .vdd(vdd), .A(asr2_en_bF_buf9), .B(_286_), .C(_287_), .Y(_270__7_) );
INVX1 INVX1_136 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf3), .Y(_271_) );
DFFSR DFFSR_113 ( .gnd(gnd), .vdd(vdd), .CLK(asr2_clk_bF_buf0), .D(_270__0_), .Q(asr2_cables_7__0_), .R(_271_), .S(vdd) );
DFFSR DFFSR_114 ( .gnd(gnd), .vdd(vdd), .CLK(asr2_clk_bF_buf3), .D(_270__1_), .Q(asr2_cables_7__1_), .R(_271_), .S(vdd) );
DFFSR DFFSR_115 ( .gnd(gnd), .vdd(vdd), .CLK(asr2_clk_bF_buf6), .D(_270__2_), .Q(asr2_cables_7__2_), .R(_271_), .S(vdd) );
DFFSR DFFSR_116 ( .gnd(gnd), .vdd(vdd), .CLK(asr2_clk_bF_buf3), .D(_270__3_), .Q(asr2_cables_7__3_), .R(_271_), .S(vdd) );
DFFSR DFFSR_117 ( .gnd(gnd), .vdd(vdd), .CLK(asr2_clk_bF_buf1), .D(_270__4_), .Q(asr2_cables_7__4_), .R(_271_), .S(vdd) );
DFFSR DFFSR_118 ( .gnd(gnd), .vdd(vdd), .CLK(asr2_clk_bF_buf2), .D(_270__5_), .Q(asr2_cables_7__5_), .R(_271_), .S(vdd) );
DFFSR DFFSR_119 ( .gnd(gnd), .vdd(vdd), .CLK(asr2_clk_bF_buf6), .D(_270__6_), .Q(asr2_cables_7__6_), .R(_271_), .S(vdd) );
DFFSR DFFSR_120 ( .gnd(gnd), .vdd(vdd), .CLK(asr2_clk_bF_buf3), .D(_270__7_), .Q(asr2_cables_7__7_), .R(_271_), .S(vdd) );
INVX1 INVX1_137 ( .gnd(gnd), .vdd(vdd), .A(asr2_cables_8__0_), .Y(_290_) );
NAND2X1 NAND2X1_121 ( .gnd(gnd), .vdd(vdd), .A(asr2_cables_7__0_), .B(asr2_en_bF_buf0), .Y(_291_) );
OAI21X1 OAI21X1_121 ( .gnd(gnd), .vdd(vdd), .A(asr2_en_bF_buf0), .B(_290_), .C(_291_), .Y(_288__0_) );
INVX1 INVX1_138 ( .gnd(gnd), .vdd(vdd), .A(asr2_cables_8__1_), .Y(_292_) );
NAND2X1 NAND2X1_122 ( .gnd(gnd), .vdd(vdd), .A(asr2_en_bF_buf8), .B(asr2_cables_7__1_), .Y(_293_) );
OAI21X1 OAI21X1_122 ( .gnd(gnd), .vdd(vdd), .A(asr2_en_bF_buf8), .B(_292_), .C(_293_), .Y(_288__1_) );
INVX1 INVX1_139 ( .gnd(gnd), .vdd(vdd), .A(asr2_cables_8__2_), .Y(_294_) );
NAND2X1 NAND2X1_123 ( .gnd(gnd), .vdd(vdd), .A(asr2_en_bF_buf10), .B(asr2_cables_7__2_), .Y(_295_) );
OAI21X1 OAI21X1_123 ( .gnd(gnd), .vdd(vdd), .A(asr2_en_bF_buf10), .B(_294_), .C(_295_), .Y(_288__2_) );
INVX1 INVX1_140 ( .gnd(gnd), .vdd(vdd), .A(asr2_cables_8__3_), .Y(_296_) );
NAND2X1 NAND2X1_124 ( .gnd(gnd), .vdd(vdd), .A(asr2_en_bF_buf8), .B(asr2_cables_7__3_), .Y(_297_) );
OAI21X1 OAI21X1_124 ( .gnd(gnd), .vdd(vdd), .A(asr2_en_bF_buf8), .B(_296_), .C(_297_), .Y(_288__3_) );
INVX1 INVX1_141 ( .gnd(gnd), .vdd(vdd), .A(asr2_cables_8__4_), .Y(_298_) );
NAND2X1 NAND2X1_125 ( .gnd(gnd), .vdd(vdd), .A(asr2_en_bF_buf7), .B(asr2_cables_7__4_), .Y(_299_) );
OAI21X1 OAI21X1_125 ( .gnd(gnd), .vdd(vdd), .A(asr2_en_bF_buf7), .B(_298_), .C(_299_), .Y(_288__4_) );
INVX1 INVX1_142 ( .gnd(gnd), .vdd(vdd), .A(asr2_cables_8__5_), .Y(_300_) );
NAND2X1 NAND2X1_126 ( .gnd(gnd), .vdd(vdd), .A(asr2_en_bF_buf3), .B(asr2_cables_7__5_), .Y(_301_) );
OAI21X1 OAI21X1_126 ( .gnd(gnd), .vdd(vdd), .A(asr2_en_bF_buf3), .B(_300_), .C(_301_), .Y(_288__5_) );
INVX1 INVX1_143 ( .gnd(gnd), .vdd(vdd), .A(asr2_cables_8__6_), .Y(_302_) );
NAND2X1 NAND2X1_127 ( .gnd(gnd), .vdd(vdd), .A(asr2_en_bF_buf6), .B(asr2_cables_7__6_), .Y(_303_) );
OAI21X1 OAI21X1_127 ( .gnd(gnd), .vdd(vdd), .A(asr2_en_bF_buf6), .B(_302_), .C(_303_), .Y(_288__6_) );
INVX1 INVX1_144 ( .gnd(gnd), .vdd(vdd), .A(asr2_cables_8__7_), .Y(_304_) );
NAND2X1 NAND2X1_128 ( .gnd(gnd), .vdd(vdd), .A(asr2_en_bF_buf1), .B(asr2_cables_7__7_), .Y(_305_) );
OAI21X1 OAI21X1_128 ( .gnd(gnd), .vdd(vdd), .A(asr2_en_bF_buf1), .B(_304_), .C(_305_), .Y(_288__7_) );
INVX1 INVX1_145 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf3), .Y(_289_) );
DFFSR DFFSR_121 ( .gnd(gnd), .vdd(vdd), .CLK(asr2_clk_bF_buf6), .D(_288__0_), .Q(asr2_cables_8__0_), .R(_289_), .S(vdd) );
DFFSR DFFSR_122 ( .gnd(gnd), .vdd(vdd), .CLK(asr2_clk_bF_buf5), .D(_288__1_), .Q(asr2_cables_8__1_), .R(_289_), .S(vdd) );
DFFSR DFFSR_123 ( .gnd(gnd), .vdd(vdd), .CLK(asr2_clk_bF_buf0), .D(_288__2_), .Q(asr2_cables_8__2_), .R(_289_), .S(vdd) );
DFFSR DFFSR_124 ( .gnd(gnd), .vdd(vdd), .CLK(asr2_clk_bF_buf5), .D(_288__3_), .Q(asr2_cables_8__3_), .R(_289_), .S(vdd) );
DFFSR DFFSR_125 ( .gnd(gnd), .vdd(vdd), .CLK(asr2_clk_bF_buf1), .D(_288__4_), .Q(asr2_cables_8__4_), .R(_289_), .S(vdd) );
DFFSR DFFSR_126 ( .gnd(gnd), .vdd(vdd), .CLK(asr2_clk_bF_buf3), .D(_288__5_), .Q(asr2_cables_8__5_), .R(_289_), .S(vdd) );
DFFSR DFFSR_127 ( .gnd(gnd), .vdd(vdd), .CLK(asr2_clk_bF_buf0), .D(_288__6_), .Q(asr2_cables_8__6_), .R(_289_), .S(vdd) );
DFFSR DFFSR_128 ( .gnd(gnd), .vdd(vdd), .CLK(asr2_clk_bF_buf3), .D(_288__7_), .Q(asr2_cables_8__7_), .R(_289_), .S(vdd) );
INVX1 INVX1_146 ( .gnd(gnd), .vdd(vdd), .A(retardo_asr_1_connect_wire_1__0_), .Y(_308_) );
NAND2X1 NAND2X1_129 ( .gnd(gnd), .vdd(vdd), .A(asr1_q_0_), .B(vdd), .Y(_309_) );
OAI21X1 OAI21X1_129 ( .gnd(gnd), .vdd(vdd), .A(vdd), .B(_308_), .C(_309_), .Y(_306__0_) );
INVX1 INVX1_147 ( .gnd(gnd), .vdd(vdd), .A(retardo_asr_1_connect_wire_1__1_), .Y(_310_) );
NAND2X1 NAND2X1_130 ( .gnd(gnd), .vdd(vdd), .A(vdd), .B(asr1_q_1_), .Y(_311_) );
OAI21X1 OAI21X1_130 ( .gnd(gnd), .vdd(vdd), .A(vdd), .B(_310_), .C(_311_), .Y(_306__1_) );
INVX1 INVX1_148 ( .gnd(gnd), .vdd(vdd), .A(retardo_asr_1_connect_wire_1__2_), .Y(_312_) );
NAND2X1 NAND2X1_131 ( .gnd(gnd), .vdd(vdd), .A(vdd), .B(asr1_q_2_), .Y(_313_) );
OAI21X1 OAI21X1_131 ( .gnd(gnd), .vdd(vdd), .A(vdd), .B(_312_), .C(_313_), .Y(_306__2_) );
INVX1 INVX1_149 ( .gnd(gnd), .vdd(vdd), .A(retardo_asr_1_connect_wire_1__3_), .Y(_314_) );
NAND2X1 NAND2X1_132 ( .gnd(gnd), .vdd(vdd), .A(vdd), .B(asr1_q_3_), .Y(_315_) );
OAI21X1 OAI21X1_132 ( .gnd(gnd), .vdd(vdd), .A(vdd), .B(_314_), .C(_315_), .Y(_306__3_) );
INVX1 INVX1_150 ( .gnd(gnd), .vdd(vdd), .A(retardo_asr_1_connect_wire_1__4_), .Y(_316_) );
NAND2X1 NAND2X1_133 ( .gnd(gnd), .vdd(vdd), .A(vdd), .B(asr1_q_4_), .Y(_317_) );
OAI21X1 OAI21X1_133 ( .gnd(gnd), .vdd(vdd), .A(vdd), .B(_316_), .C(_317_), .Y(_306__4_) );
INVX1 INVX1_151 ( .gnd(gnd), .vdd(vdd), .A(retardo_asr_1_connect_wire_1__5_), .Y(_318_) );
NAND2X1 NAND2X1_134 ( .gnd(gnd), .vdd(vdd), .A(vdd), .B(asr1_q_5_), .Y(_319_) );
OAI21X1 OAI21X1_134 ( .gnd(gnd), .vdd(vdd), .A(vdd), .B(_318_), .C(_319_), .Y(_306__5_) );
INVX1 INVX1_152 ( .gnd(gnd), .vdd(vdd), .A(retardo_asr_1_connect_wire_1__6_), .Y(_320_) );
NAND2X1 NAND2X1_135 ( .gnd(gnd), .vdd(vdd), .A(vdd), .B(asr1_q_6_), .Y(_321_) );
OAI21X1 OAI21X1_135 ( .gnd(gnd), .vdd(vdd), .A(vdd), .B(_320_), .C(_321_), .Y(_306__6_) );
INVX1 INVX1_153 ( .gnd(gnd), .vdd(vdd), .A(retardo_asr_1_connect_wire_1__7_), .Y(_322_) );
NAND2X1 NAND2X1_136 ( .gnd(gnd), .vdd(vdd), .A(vdd), .B(asr1_q_7_), .Y(_323_) );
OAI21X1 OAI21X1_136 ( .gnd(gnd), .vdd(vdd), .A(vdd), .B(_322_), .C(_323_), .Y(_306__7_) );
INVX1 INVX1_154 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf4), .Y(_307_) );
DFFSR DFFSR_129 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf1), .D(_306__0_), .Q(retardo_asr_1_connect_wire_1__0_), .R(_307_), .S(vdd) );
DFFSR DFFSR_130 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf1), .D(_306__1_), .Q(retardo_asr_1_connect_wire_1__1_), .R(_307_), .S(vdd) );
DFFSR DFFSR_131 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf0), .D(_306__2_), .Q(retardo_asr_1_connect_wire_1__2_), .R(_307_), .S(vdd) );
DFFSR DFFSR_132 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf0), .D(_306__3_), .Q(retardo_asr_1_connect_wire_1__3_), .R(_307_), .S(vdd) );
DFFSR DFFSR_133 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf1), .D(_306__4_), .Q(retardo_asr_1_connect_wire_1__4_), .R(_307_), .S(vdd) );
DFFSR DFFSR_134 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf1), .D(_306__5_), .Q(retardo_asr_1_connect_wire_1__5_), .R(_307_), .S(vdd) );
DFFSR DFFSR_135 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf0), .D(_306__6_), .Q(retardo_asr_1_connect_wire_1__6_), .R(_307_), .S(vdd) );
DFFSR DFFSR_136 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf1), .D(_306__7_), .Q(retardo_asr_1_connect_wire_1__7_), .R(_307_), .S(vdd) );
INVX1 INVX1_155 ( .gnd(gnd), .vdd(vdd), .A(retardo_asr_2_connect_wire_1__0_), .Y(_326_) );
NAND2X1 NAND2X1_137 ( .gnd(gnd), .vdd(vdd), .A(asr2_q_0_), .B(vdd), .Y(_327_) );
OAI21X1 OAI21X1_137 ( .gnd(gnd), .vdd(vdd), .A(vdd), .B(_326_), .C(_327_), .Y(_324__0_) );
INVX1 INVX1_156 ( .gnd(gnd), .vdd(vdd), .A(retardo_asr_2_connect_wire_1__1_), .Y(_328_) );
NAND2X1 NAND2X1_138 ( .gnd(gnd), .vdd(vdd), .A(vdd), .B(asr2_q_1_), .Y(_329_) );
OAI21X1 OAI21X1_138 ( .gnd(gnd), .vdd(vdd), .A(vdd), .B(_328_), .C(_329_), .Y(_324__1_) );
INVX1 INVX1_157 ( .gnd(gnd), .vdd(vdd), .A(retardo_asr_2_connect_wire_1__2_), .Y(_330_) );
NAND2X1 NAND2X1_139 ( .gnd(gnd), .vdd(vdd), .A(vdd), .B(asr2_q_2_), .Y(_331_) );
OAI21X1 OAI21X1_139 ( .gnd(gnd), .vdd(vdd), .A(vdd), .B(_330_), .C(_331_), .Y(_324__2_) );
INVX1 INVX1_158 ( .gnd(gnd), .vdd(vdd), .A(retardo_asr_2_connect_wire_1__3_), .Y(_332_) );
NAND2X1 NAND2X1_140 ( .gnd(gnd), .vdd(vdd), .A(vdd), .B(asr2_q_3_), .Y(_333_) );
OAI21X1 OAI21X1_140 ( .gnd(gnd), .vdd(vdd), .A(vdd), .B(_332_), .C(_333_), .Y(_324__3_) );
INVX1 INVX1_159 ( .gnd(gnd), .vdd(vdd), .A(retardo_asr_2_connect_wire_1__4_), .Y(_334_) );
NAND2X1 NAND2X1_141 ( .gnd(gnd), .vdd(vdd), .A(vdd), .B(asr2_q_4_), .Y(_335_) );
OAI21X1 OAI21X1_141 ( .gnd(gnd), .vdd(vdd), .A(vdd), .B(_334_), .C(_335_), .Y(_324__4_) );
INVX1 INVX1_160 ( .gnd(gnd), .vdd(vdd), .A(retardo_asr_2_connect_wire_1__5_), .Y(_336_) );
NAND2X1 NAND2X1_142 ( .gnd(gnd), .vdd(vdd), .A(vdd), .B(asr2_q_5_), .Y(_337_) );
OAI21X1 OAI21X1_142 ( .gnd(gnd), .vdd(vdd), .A(vdd), .B(_336_), .C(_337_), .Y(_324__5_) );
INVX1 INVX1_161 ( .gnd(gnd), .vdd(vdd), .A(retardo_asr_2_connect_wire_1__6_), .Y(_338_) );
NAND2X1 NAND2X1_143 ( .gnd(gnd), .vdd(vdd), .A(vdd), .B(asr2_q_6_), .Y(_339_) );
OAI21X1 OAI21X1_143 ( .gnd(gnd), .vdd(vdd), .A(vdd), .B(_338_), .C(_339_), .Y(_324__6_) );
INVX1 INVX1_162 ( .gnd(gnd), .vdd(vdd), .A(retardo_asr_2_connect_wire_1__7_), .Y(_340_) );
NAND2X1 NAND2X1_144 ( .gnd(gnd), .vdd(vdd), .A(vdd), .B(asr2_q_7_), .Y(_341_) );
OAI21X1 OAI21X1_144 ( .gnd(gnd), .vdd(vdd), .A(vdd), .B(_340_), .C(_341_), .Y(_324__7_) );
INVX1 INVX1_163 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf4), .Y(_325_) );
DFFSR DFFSR_137 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf1), .D(_324__0_), .Q(retardo_asr_2_connect_wire_1__0_), .R(_325_), .S(vdd) );
DFFSR DFFSR_138 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf0), .D(_324__1_), .Q(retardo_asr_2_connect_wire_1__1_), .R(_325_), .S(vdd) );
DFFSR DFFSR_139 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf0), .D(_324__2_), .Q(retardo_asr_2_connect_wire_1__2_), .R(_325_), .S(vdd) );
DFFSR DFFSR_140 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf0), .D(_324__3_), .Q(retardo_asr_2_connect_wire_1__3_), .R(_325_), .S(vdd) );
DFFSR DFFSR_141 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf3), .D(_324__4_), .Q(retardo_asr_2_connect_wire_1__4_), .R(_325_), .S(vdd) );
DFFSR DFFSR_142 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf0), .D(_324__5_), .Q(retardo_asr_2_connect_wire_1__5_), .R(_325_), .S(vdd) );
DFFSR DFFSR_143 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf0), .D(_324__6_), .Q(retardo_asr_2_connect_wire_1__6_), .R(_325_), .S(vdd) );
DFFSR DFFSR_144 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf0), .D(_324__7_), .Q(retardo_asr_2_connect_wire_1__7_), .R(_325_), .S(vdd) );
INVX1 INVX1_164 ( .gnd(gnd), .vdd(vdd), .A(retardo_clock_chico_connect_wire_1_), .Y(_344_) );
NAND2X1 NAND2X1_145 ( .gnd(gnd), .vdd(vdd), .A(enable_asr), .B(vdd), .Y(_345_) );
OAI21X1 OAI21X1_145 ( .gnd(gnd), .vdd(vdd), .A(vdd), .B(_344_), .C(_345_), .Y(_342_) );
INVX1 INVX1_165 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf4), .Y(_343_) );
DFFSR DFFSR_145 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf2), .D(_342_), .Q(retardo_clock_chico_connect_wire_1_), .R(_343_), .S(vdd) );
INVX1 INVX1_166 ( .gnd(gnd), .vdd(vdd), .A(retardo_clock_chico_connect_wire_2_), .Y(_348_) );
NAND2X1 NAND2X1_146 ( .gnd(gnd), .vdd(vdd), .A(retardo_clock_chico_connect_wire_1_), .B(vdd), .Y(_349_) );
OAI21X1 OAI21X1_146 ( .gnd(gnd), .vdd(vdd), .A(vdd), .B(_348_), .C(_349_), .Y(_346_) );
INVX1 INVX1_167 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf1), .Y(_347_) );
DFFSR DFFSR_146 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf2), .D(_346_), .Q(retardo_clock_chico_connect_wire_2_), .R(_347_), .S(vdd) );
INVX1 INVX1_168 ( .gnd(gnd), .vdd(vdd), .A(retardo_clock_chico_connect_wire_3_), .Y(_352_) );
NAND2X1 NAND2X1_147 ( .gnd(gnd), .vdd(vdd), .A(retardo_clock_chico_connect_wire_2_), .B(vdd), .Y(_353_) );
OAI21X1 OAI21X1_147 ( .gnd(gnd), .vdd(vdd), .A(vdd), .B(_352_), .C(_353_), .Y(_350_) );
INVX1 INVX1_169 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf4), .Y(_351_) );
DFFSR DFFSR_147 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf1), .D(_350_), .Q(retardo_clock_chico_connect_wire_3_), .R(_351_), .S(vdd) );
INVX1 INVX1_170 ( .gnd(gnd), .vdd(vdd), .A(retardo_clock_chico_connect_wire_4_), .Y(_356_) );
NAND2X1 NAND2X1_148 ( .gnd(gnd), .vdd(vdd), .A(retardo_clock_chico_connect_wire_3_), .B(vdd), .Y(_357_) );
OAI21X1 OAI21X1_148 ( .gnd(gnd), .vdd(vdd), .A(vdd), .B(_356_), .C(_357_), .Y(_354_) );
INVX1 INVX1_171 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf4), .Y(_355_) );
DFFSR DFFSR_148 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf1), .D(_354_), .Q(retardo_clock_chico_connect_wire_4_), .R(_355_), .S(vdd) );
INVX1 INVX1_172 ( .gnd(gnd), .vdd(vdd), .A(asr2_clk_bF_buf4), .Y(_360_) );
NAND2X1 NAND2X1_149 ( .gnd(gnd), .vdd(vdd), .A(retardo_clock_chico_connect_wire_4_), .B(vdd), .Y(_361_) );
OAI21X1 OAI21X1_149 ( .gnd(gnd), .vdd(vdd), .A(vdd), .B(_360_), .C(_361_), .Y(_358_) );
INVX1 INVX1_173 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf5), .Y(_359_) );
DFFSR DFFSR_149 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf4), .D(_358_), .Q(asr2_clk), .R(_359_), .S(vdd) );
INVX1 INVX1_174 ( .gnd(gnd), .vdd(vdd), .A(retardo_clock_mac_connect_wire_1_), .Y(_364_) );
NAND2X1 NAND2X1_150 ( .gnd(gnd), .vdd(vdd), .A(enable_asr), .B(vdd), .Y(_365_) );
OAI21X1 OAI21X1_150 ( .gnd(gnd), .vdd(vdd), .A(vdd), .B(_364_), .C(_365_), .Y(_362_) );
INVX1 INVX1_175 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf1), .Y(_363_) );
DFFSR DFFSR_150 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf2), .D(_362_), .Q(retardo_clock_mac_connect_wire_1_), .R(_363_), .S(vdd) );
INVX1 INVX1_176 ( .gnd(gnd), .vdd(vdd), .A(retardo_clock_mac_connect_wire_2_), .Y(_368_) );
NAND2X1 NAND2X1_151 ( .gnd(gnd), .vdd(vdd), .A(retardo_clock_mac_connect_wire_1_), .B(vdd), .Y(_369_) );
OAI21X1 OAI21X1_151 ( .gnd(gnd), .vdd(vdd), .A(vdd), .B(_368_), .C(_369_), .Y(_366_) );
INVX1 INVX1_177 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf5), .Y(_367_) );
DFFSR DFFSR_151 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf4), .D(_366_), .Q(retardo_clock_mac_connect_wire_2_), .R(_367_), .S(vdd) );
INVX1 INVX1_178 ( .gnd(gnd), .vdd(vdd), .A(retardo_clock_mac_connect_wire_3_), .Y(_372_) );
NAND2X1 NAND2X1_152 ( .gnd(gnd), .vdd(vdd), .A(retardo_clock_mac_connect_wire_2_), .B(vdd), .Y(_373_) );
OAI21X1 OAI21X1_152 ( .gnd(gnd), .vdd(vdd), .A(vdd), .B(_372_), .C(_373_), .Y(_370_) );
INVX1 INVX1_179 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf1), .Y(_371_) );
DFFSR DFFSR_152 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf4), .D(_370_), .Q(retardo_clock_mac_connect_wire_3_), .R(_371_), .S(vdd) );
INVX1 INVX1_180 ( .gnd(gnd), .vdd(vdd), .A(retardo_clock_mac_connect_wire_4_), .Y(_376_) );
NAND2X1 NAND2X1_153 ( .gnd(gnd), .vdd(vdd), .A(retardo_clock_mac_connect_wire_3_), .B(vdd), .Y(_377_) );
OAI21X1 OAI21X1_153 ( .gnd(gnd), .vdd(vdd), .A(vdd), .B(_376_), .C(_377_), .Y(_374_) );
INVX1 INVX1_181 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf4), .Y(_375_) );
DFFSR DFFSR_153 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf3), .D(_374_), .Q(retardo_clock_mac_connect_wire_4_), .R(_375_), .S(vdd) );
INVX1 INVX1_182 ( .gnd(gnd), .vdd(vdd), .A(retardo_clock_mac_connect_wire_5_), .Y(_380_) );
NAND2X1 NAND2X1_154 ( .gnd(gnd), .vdd(vdd), .A(retardo_clock_mac_connect_wire_4_), .B(vdd), .Y(_381_) );
OAI21X1 OAI21X1_154 ( .gnd(gnd), .vdd(vdd), .A(vdd), .B(_380_), .C(_381_), .Y(_378_) );
INVX1 INVX1_183 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf4), .Y(_379_) );
DFFSR DFFSR_154 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf4), .D(_378_), .Q(retardo_clock_mac_connect_wire_5_), .R(_379_), .S(vdd) );
INVX1 INVX1_184 ( .gnd(gnd), .vdd(vdd), .A(retardo_clock_mac_connect_wire_6_), .Y(_384_) );
NAND2X1 NAND2X1_155 ( .gnd(gnd), .vdd(vdd), .A(retardo_clock_mac_connect_wire_5_), .B(vdd), .Y(_385_) );
OAI21X1 OAI21X1_155 ( .gnd(gnd), .vdd(vdd), .A(vdd), .B(_384_), .C(_385_), .Y(_382_) );
INVX1 INVX1_185 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf5), .Y(_383_) );
DFFSR DFFSR_155 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf4), .D(_382_), .Q(retardo_clock_mac_connect_wire_6_), .R(_383_), .S(vdd) );
INVX1 INVX1_186 ( .gnd(gnd), .vdd(vdd), .A(retardo_clock_mac_connect_wire_7_), .Y(_388_) );
NAND2X1 NAND2X1_156 ( .gnd(gnd), .vdd(vdd), .A(retardo_clock_mac_connect_wire_6_), .B(vdd), .Y(_389_) );
OAI21X1 OAI21X1_156 ( .gnd(gnd), .vdd(vdd), .A(vdd), .B(_388_), .C(_389_), .Y(_386_) );
INVX1 INVX1_187 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf5), .Y(_387_) );
DFFSR DFFSR_156 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf4), .D(_386_), .Q(retardo_clock_mac_connect_wire_7_), .R(_387_), .S(vdd) );
INVX1 INVX1_188 ( .gnd(gnd), .vdd(vdd), .A(retardo_clock_mac_connect_wire_8_), .Y(_392_) );
NAND2X1 NAND2X1_157 ( .gnd(gnd), .vdd(vdd), .A(retardo_clock_mac_connect_wire_7_), .B(vdd), .Y(_393_) );
OAI21X1 OAI21X1_157 ( .gnd(gnd), .vdd(vdd), .A(vdd), .B(_392_), .C(_393_), .Y(_390_) );
INVX1 INVX1_189 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf1), .Y(_391_) );
DFFSR DFFSR_157 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf2), .D(_390_), .Q(retardo_clock_mac_connect_wire_8_), .R(_391_), .S(vdd) );
INVX1 INVX1_190 ( .gnd(gnd), .vdd(vdd), .A(retardo_clock_mac_connect_wire_9_), .Y(_396_) );
NAND2X1 NAND2X1_158 ( .gnd(gnd), .vdd(vdd), .A(retardo_clock_mac_connect_wire_8_), .B(vdd), .Y(_397_) );
OAI21X1 OAI21X1_158 ( .gnd(gnd), .vdd(vdd), .A(vdd), .B(_396_), .C(_397_), .Y(_394_) );
INVX1 INVX1_191 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf0), .Y(_395_) );
DFFSR DFFSR_158 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf7), .D(_394_), .Q(retardo_clock_mac_connect_wire_9_), .R(_395_), .S(vdd) );
INVX1 INVX1_192 ( .gnd(gnd), .vdd(vdd), .A(MAC_clr_bF_buf3), .Y(_400_) );
NAND2X1 NAND2X1_159 ( .gnd(gnd), .vdd(vdd), .A(retardo_clock_mac_connect_wire_9_), .B(vdd), .Y(_401_) );
OAI21X1 OAI21X1_159 ( .gnd(gnd), .vdd(vdd), .A(vdd), .B(_400_), .C(_401_), .Y(_398_) );
INVX1 INVX1_193 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf0), .Y(_399_) );
DFFSR DFFSR_159 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf7), .D(_398_), .Q(MAC_clr), .R(_399_), .S(vdd) );
INVX1 INVX1_194 ( .gnd(gnd), .vdd(vdd), .A(registro_salida_d_0_), .Y(_404_) );
NAND2X1 NAND2X1_160 ( .gnd(gnd), .vdd(vdd), .A(MAC_salida_correcta_0_), .B(MAC_clr_bF_buf0), .Y(_405_) );
OAI21X1 OAI21X1_160 ( .gnd(gnd), .vdd(vdd), .A(MAC_clr_bF_buf2), .B(_404_), .C(_405_), .Y(_402__0_) );
INVX1 INVX1_195 ( .gnd(gnd), .vdd(vdd), .A(registro_salida_d_1_), .Y(_406_) );
NAND2X1 NAND2X1_161 ( .gnd(gnd), .vdd(vdd), .A(MAC_clr_bF_buf0), .B(MAC_salida_correcta_1_), .Y(_407_) );
OAI21X1 OAI21X1_161 ( .gnd(gnd), .vdd(vdd), .A(MAC_clr_bF_buf2), .B(_406_), .C(_407_), .Y(_402__1_) );
INVX1 INVX1_196 ( .gnd(gnd), .vdd(vdd), .A(registro_salida_d_2_), .Y(_408_) );
NAND2X1 NAND2X1_162 ( .gnd(gnd), .vdd(vdd), .A(MAC_clr_bF_buf3), .B(MAC_salida_correcta_2_), .Y(_409_) );
OAI21X1 OAI21X1_162 ( .gnd(gnd), .vdd(vdd), .A(MAC_clr_bF_buf0), .B(_408_), .C(_409_), .Y(_402__2_) );
INVX1 INVX1_197 ( .gnd(gnd), .vdd(vdd), .A(registro_salida_d_3_), .Y(_410_) );
NAND2X1 NAND2X1_163 ( .gnd(gnd), .vdd(vdd), .A(MAC_clr_bF_buf2), .B(MAC_salida_correcta_3_), .Y(_411_) );
OAI21X1 OAI21X1_163 ( .gnd(gnd), .vdd(vdd), .A(MAC_clr_bF_buf2), .B(_410_), .C(_411_), .Y(_402__3_) );
INVX1 INVX1_198 ( .gnd(gnd), .vdd(vdd), .A(registro_salida_d_4_), .Y(_412_) );
NAND2X1 NAND2X1_164 ( .gnd(gnd), .vdd(vdd), .A(MAC_clr_bF_buf3), .B(MAC_salida_correcta_4_), .Y(_413_) );
OAI21X1 OAI21X1_164 ( .gnd(gnd), .vdd(vdd), .A(MAC_clr_bF_buf2), .B(_412_), .C(_413_), .Y(_402__4_) );
INVX1 INVX1_199 ( .gnd(gnd), .vdd(vdd), .A(registro_salida_d_5_), .Y(_414_) );
NAND2X1 NAND2X1_165 ( .gnd(gnd), .vdd(vdd), .A(MAC_clr_bF_buf0), .B(MAC_salida_correcta_5_), .Y(_415_) );
OAI21X1 OAI21X1_165 ( .gnd(gnd), .vdd(vdd), .A(MAC_clr_bF_buf1), .B(_414_), .C(_415_), .Y(_402__5_) );
INVX1 INVX1_200 ( .gnd(gnd), .vdd(vdd), .A(registro_salida_d_6_), .Y(_416_) );
NAND2X1 NAND2X1_166 ( .gnd(gnd), .vdd(vdd), .A(MAC_clr_bF_buf1), .B(MAC_salida_correcta_6_), .Y(_417_) );
OAI21X1 OAI21X1_166 ( .gnd(gnd), .vdd(vdd), .A(MAC_clr_bF_buf1), .B(_416_), .C(_417_), .Y(_402__6_) );
INVX1 INVX1_201 ( .gnd(gnd), .vdd(vdd), .A(registro_salida_d_7_), .Y(_418_) );
NAND2X1 NAND2X1_167 ( .gnd(gnd), .vdd(vdd), .A(MAC_clr_bF_buf1), .B(MAC_salida_correcta_7_), .Y(_419_) );
OAI21X1 OAI21X1_167 ( .gnd(gnd), .vdd(vdd), .A(MAC_clr_bF_buf1), .B(_418_), .C(_419_), .Y(_402__7_) );
INVX1 INVX1_202 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf0), .Y(_403_) );
DFFSR DFFSR_160 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf5), .D(_402__0_), .Q(registro_salida_d_0_), .R(_403_), .S(vdd) );
DFFSR DFFSR_161 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf7), .D(_402__1_), .Q(registro_salida_d_1_), .R(_403_), .S(vdd) );
DFFSR DFFSR_162 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf7), .D(_402__2_), .Q(registro_salida_d_2_), .R(_403_), .S(vdd) );
DFFSR DFFSR_163 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf5), .D(_402__3_), .Q(registro_salida_d_3_), .R(_403_), .S(vdd) );
DFFSR DFFSR_164 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf7), .D(_402__4_), .Q(registro_salida_d_4_), .R(_403_), .S(vdd) );
DFFSR DFFSR_165 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf5), .D(_402__5_), .Q(registro_salida_d_5_), .R(_403_), .S(vdd) );
DFFSR DFFSR_166 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf5), .D(_402__6_), .Q(registro_salida_d_6_), .R(_403_), .S(vdd) );
DFFSR DFFSR_167 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf5), .D(_402__7_), .Q(registro_salida_d_7_), .R(_403_), .S(vdd) );
INVX1 INVX1_203 ( .gnd(gnd), .vdd(vdd), .A(MAC_ROM_0_bF_buf3_), .Y(_422_) );
NAND2X1 NAND2X1_168 ( .gnd(gnd), .vdd(vdd), .A(memoria_q_0_), .B(vdd), .Y(_423_) );
OAI21X1 OAI21X1_168 ( .gnd(gnd), .vdd(vdd), .A(vdd), .B(_422_), .C(_423_), .Y(_420__0_) );
INVX1 INVX1_204 ( .gnd(gnd), .vdd(vdd), .A(MAC_ROM_1_), .Y(_424_) );
NAND2X1 NAND2X1_169 ( .gnd(gnd), .vdd(vdd), .A(vdd), .B(memoria_q_1_), .Y(_425_) );
OAI21X1 OAI21X1_169 ( .gnd(gnd), .vdd(vdd), .A(vdd), .B(_424_), .C(_425_), .Y(_420__1_) );
INVX1 INVX1_205 ( .gnd(gnd), .vdd(vdd), .A(MAC_ROM_2_), .Y(_426_) );
NAND2X1 NAND2X1_170 ( .gnd(gnd), .vdd(vdd), .A(vdd), .B(memoria_q_2_), .Y(_427_) );
OAI21X1 OAI21X1_170 ( .gnd(gnd), .vdd(vdd), .A(vdd), .B(_426_), .C(_427_), .Y(_420__2_) );
INVX1 INVX1_206 ( .gnd(gnd), .vdd(vdd), .A(MAC_ROM_3_), .Y(_428_) );
NAND2X1 NAND2X1_171 ( .gnd(gnd), .vdd(vdd), .A(vdd), .B(memoria_q_3_), .Y(_429_) );
OAI21X1 OAI21X1_171 ( .gnd(gnd), .vdd(vdd), .A(vdd), .B(_428_), .C(_429_), .Y(_420__3_) );
INVX1 INVX1_207 ( .gnd(gnd), .vdd(vdd), .A(MAC_ROM_4_), .Y(_430_) );
NAND2X1 NAND2X1_172 ( .gnd(gnd), .vdd(vdd), .A(vdd), .B(gnd), .Y(_431_) );
OAI21X1 OAI21X1_172 ( .gnd(gnd), .vdd(vdd), .A(vdd), .B(_430_), .C(_431_), .Y(_420__4_) );
INVX1 INVX1_208 ( .gnd(gnd), .vdd(vdd), .A(MAC_ROM_5_), .Y(_432_) );
NAND2X1 NAND2X1_173 ( .gnd(gnd), .vdd(vdd), .A(vdd), .B(gnd), .Y(_433_) );
OAI21X1 OAI21X1_173 ( .gnd(gnd), .vdd(vdd), .A(vdd), .B(_432_), .C(_433_), .Y(_420__5_) );
INVX1 INVX1_209 ( .gnd(gnd), .vdd(vdd), .A(MAC_ROM_6_), .Y(_434_) );
NAND2X1 NAND2X1_174 ( .gnd(gnd), .vdd(vdd), .A(vdd), .B(gnd), .Y(_435_) );
OAI21X1 OAI21X1_174 ( .gnd(gnd), .vdd(vdd), .A(vdd), .B(_434_), .C(_435_), .Y(_420__6_) );
INVX1 INVX1_210 ( .gnd(gnd), .vdd(vdd), .A(MAC_ROM_7_), .Y(_436_) );
NAND2X1 NAND2X1_175 ( .gnd(gnd), .vdd(vdd), .A(vdd), .B(gnd), .Y(_437_) );
OAI21X1 OAI21X1_175 ( .gnd(gnd), .vdd(vdd), .A(vdd), .B(_436_), .C(_437_), .Y(_420__7_) );
INVX1 INVX1_211 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf4), .Y(_421_) );
DFFSR DFFSR_168 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf3), .D(_420__0_), .Q(MAC_ROM_0_), .R(_421_), .S(vdd) );
DFFSR DFFSR_169 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf3), .D(_420__1_), .Q(MAC_ROM_1_), .R(_421_), .S(vdd) );
DFFSR DFFSR_170 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf3), .D(_420__2_), .Q(MAC_ROM_2_), .R(_421_), .S(vdd) );
DFFSR DFFSR_171 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf6), .D(_420__3_), .Q(MAC_ROM_3_), .R(_421_), .S(vdd) );
DFFSR DFFSR_172 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf3), .D(_420__4_), .Q(MAC_ROM_4_), .R(_421_), .S(vdd) );
DFFSR DFFSR_173 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf6), .D(_420__5_), .Q(MAC_ROM_5_), .R(_421_), .S(vdd) );
DFFSR DFFSR_174 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf6), .D(_420__6_), .Q(MAC_ROM_6_), .R(_421_), .S(vdd) );
DFFSR DFFSR_175 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf6), .D(_420__7_), .Q(MAC_ROM_7_), .R(_421_), .S(vdd) );
NAND2X1 NAND2X1_176 ( .gnd(gnd), .vdd(vdd), .A(MAC_ROM_0_bF_buf2_), .B(MAC_Adder_0_), .Y(_685_) );
INVX1 INVX1_212 ( .gnd(gnd), .vdd(vdd), .A(MAC_clr_bF_buf3), .Y(_696_) );
NAND2X1 NAND2X1_177 ( .gnd(gnd), .vdd(vdd), .A(MAC_salida_correcta_0_), .B(_696_), .Y(_707_) );
XOR2X1 XOR2X1_1 ( .gnd(gnd), .vdd(vdd), .A(_707_), .B(_685_), .Y(_438__0_) );
INVX1 INVX1_213 ( .gnd(gnd), .vdd(vdd), .A(MAC_ROM_0_bF_buf1_), .Y(_728_) );
INVX1 INVX1_214 ( .gnd(gnd), .vdd(vdd), .A(MAC_Adder_0_), .Y(_739_) );
INVX1 INVX1_215 ( .gnd(gnd), .vdd(vdd), .A(MAC_Adder_1_), .Y(_746_) );
INVX1 INVX1_216 ( .gnd(gnd), .vdd(vdd), .A(MAC_ROM_1_), .Y(_747_) );
OAI22X1 OAI22X1_1 ( .gnd(gnd), .vdd(vdd), .A(_728_), .B(_746_), .C(_739_), .D(_747_), .Y(_748_) );
NAND2X1 NAND2X1_178 ( .gnd(gnd), .vdd(vdd), .A(MAC_Adder_1_), .B(MAC_ROM_1_), .Y(_749_) );
OAI21X1 OAI21X1_176 ( .gnd(gnd), .vdd(vdd), .A(_685_), .B(_749_), .C(_748_), .Y(_750_) );
NAND3X1 NAND3X1_1 ( .gnd(gnd), .vdd(vdd), .A(MAC_ROM_0_bF_buf0_), .B(MAC_Adder_0_), .C(MAC_salida_correcta_0_), .Y(_751_) );
INVX1 INVX1_217 ( .gnd(gnd), .vdd(vdd), .A(_751_), .Y(_752_) );
INVX1 INVX1_218 ( .gnd(gnd), .vdd(vdd), .A(MAC_salida_correcta_1_), .Y(_753_) );
XOR2X1 XOR2X1_2 ( .gnd(gnd), .vdd(vdd), .A(_750_), .B(_753_), .Y(_754_) );
NAND2X1 NAND2X1_179 ( .gnd(gnd), .vdd(vdd), .A(_752_), .B(_754_), .Y(_755_) );
OR2X2 OR2X2_1 ( .gnd(gnd), .vdd(vdd), .A(_754_), .B(_752_), .Y(_756_) );
NAND3X1 NAND3X1_2 ( .gnd(gnd), .vdd(vdd), .A(_696_), .B(_755_), .C(_756_), .Y(_757_) );
OAI21X1 OAI21X1_177 ( .gnd(gnd), .vdd(vdd), .A(_696_), .B(_750_), .C(_757_), .Y(_438__1_) );
NAND2X1 NAND2X1_180 ( .gnd(gnd), .vdd(vdd), .A(MAC_Adder_0_), .B(MAC_ROM_2_), .Y(_758_) );
INVX1 INVX1_219 ( .gnd(gnd), .vdd(vdd), .A(_758_), .Y(_759_) );
AND2X2 AND2X2_2 ( .gnd(gnd), .vdd(vdd), .A(MAC_ROM_0_bF_buf3_), .B(MAC_Adder_2_), .Y(_760_) );
NAND3X1 NAND3X1_3 ( .gnd(gnd), .vdd(vdd), .A(MAC_Adder_1_), .B(MAC_ROM_1_), .C(_760_), .Y(_761_) );
AOI22X1 AOI22X1_1 ( .gnd(gnd), .vdd(vdd), .A(MAC_ROM_0_bF_buf2_), .B(MAC_Adder_2_), .C(MAC_Adder_1_), .D(MAC_ROM_1_), .Y(_762_) );
INVX1 INVX1_220 ( .gnd(gnd), .vdd(vdd), .A(_762_), .Y(_763_) );
NAND3X1 NAND3X1_4 ( .gnd(gnd), .vdd(vdd), .A(_763_), .B(_759_), .C(_761_), .Y(_764_) );
NAND2X1 NAND2X1_181 ( .gnd(gnd), .vdd(vdd), .A(MAC_ROM_0_bF_buf1_), .B(MAC_Adder_2_), .Y(_765_) );
NOR2X1 NOR2X1_3 ( .gnd(gnd), .vdd(vdd), .A(_749_), .B(_765_), .Y(_766_) );
OAI21X1 OAI21X1_178 ( .gnd(gnd), .vdd(vdd), .A(_762_), .B(_766_), .C(_758_), .Y(_767_) );
NAND2X1 NAND2X1_182 ( .gnd(gnd), .vdd(vdd), .A(_764_), .B(_767_), .Y(_768_) );
OAI21X1 OAI21X1_179 ( .gnd(gnd), .vdd(vdd), .A(_685_), .B(_749_), .C(_768_), .Y(_769_) );
NOR2X1 NOR2X1_4 ( .gnd(gnd), .vdd(vdd), .A(_685_), .B(_749_), .Y(_770_) );
NAND3X1 NAND3X1_5 ( .gnd(gnd), .vdd(vdd), .A(_770_), .B(_764_), .C(_767_), .Y(_771_) );
NAND2X1 NAND2X1_183 ( .gnd(gnd), .vdd(vdd), .A(_771_), .B(_769_), .Y(_772_) );
OAI21X1 OAI21X1_180 ( .gnd(gnd), .vdd(vdd), .A(_753_), .B(_750_), .C(_755_), .Y(_773_) );
INVX1 INVX1_221 ( .gnd(gnd), .vdd(vdd), .A(_773_), .Y(_774_) );
NAND3X1 NAND3X1_6 ( .gnd(gnd), .vdd(vdd), .A(MAC_salida_correcta_2_), .B(_771_), .C(_769_), .Y(_775_) );
INVX1 INVX1_222 ( .gnd(gnd), .vdd(vdd), .A(_775_), .Y(_776_) );
AOI21X1 AOI21X1_1 ( .gnd(gnd), .vdd(vdd), .A(_769_), .B(_771_), .C(MAC_salida_correcta_2_), .Y(_777_) );
NOR2X1 NOR2X1_5 ( .gnd(gnd), .vdd(vdd), .A(_777_), .B(_776_), .Y(_778_) );
AND2X2 AND2X2_3 ( .gnd(gnd), .vdd(vdd), .A(_778_), .B(_774_), .Y(_779_) );
NOR2X1 NOR2X1_6 ( .gnd(gnd), .vdd(vdd), .A(_774_), .B(_778_), .Y(_780_) );
OAI21X1 OAI21X1_181 ( .gnd(gnd), .vdd(vdd), .A(_780_), .B(_779_), .C(_696_), .Y(_781_) );
OAI21X1 OAI21X1_182 ( .gnd(gnd), .vdd(vdd), .A(_696_), .B(_772_), .C(_781_), .Y(_438__2_) );
OAI21X1 OAI21X1_183 ( .gnd(gnd), .vdd(vdd), .A(_777_), .B(_774_), .C(_775_), .Y(_782_) );
INVX1 INVX1_223 ( .gnd(gnd), .vdd(vdd), .A(_771_), .Y(_783_) );
NAND2X1 NAND2X1_184 ( .gnd(gnd), .vdd(vdd), .A(MAC_Adder_0_), .B(MAC_ROM_3_), .Y(_784_) );
INVX1 INVX1_224 ( .gnd(gnd), .vdd(vdd), .A(_784_), .Y(_785_) );
OAI21X1 OAI21X1_184 ( .gnd(gnd), .vdd(vdd), .A(_758_), .B(_762_), .C(_761_), .Y(_786_) );
NAND2X1 NAND2X1_185 ( .gnd(gnd), .vdd(vdd), .A(MAC_Adder_1_), .B(MAC_ROM_2_), .Y(_787_) );
INVX1 INVX1_225 ( .gnd(gnd), .vdd(vdd), .A(_787_), .Y(_788_) );
AND2X2 AND2X2_4 ( .gnd(gnd), .vdd(vdd), .A(MAC_ROM_1_), .B(MAC_Adder_2_), .Y(_789_) );
AND2X2 AND2X2_5 ( .gnd(gnd), .vdd(vdd), .A(MAC_ROM_0_bF_buf0_), .B(MAC_Adder_3_), .Y(_790_) );
NAND2X1 NAND2X1_186 ( .gnd(gnd), .vdd(vdd), .A(_789_), .B(_790_), .Y(_791_) );
INVX1 INVX1_226 ( .gnd(gnd), .vdd(vdd), .A(MAC_Adder_2_), .Y(_792_) );
NAND2X1 NAND2X1_187 ( .gnd(gnd), .vdd(vdd), .A(MAC_ROM_0_bF_buf3_), .B(MAC_Adder_3_), .Y(_793_) );
OAI21X1 OAI21X1_185 ( .gnd(gnd), .vdd(vdd), .A(_747_), .B(_792_), .C(_793_), .Y(_794_) );
NAND3X1 NAND3X1_7 ( .gnd(gnd), .vdd(vdd), .A(_794_), .B(_788_), .C(_791_), .Y(_795_) );
OAI21X1 OAI21X1_186 ( .gnd(gnd), .vdd(vdd), .A(_747_), .B(_792_), .C(_790_), .Y(_796_) );
INVX1 INVX1_227 ( .gnd(gnd), .vdd(vdd), .A(MAC_Adder_3_), .Y(_797_) );
OAI21X1 OAI21X1_187 ( .gnd(gnd), .vdd(vdd), .A(_728_), .B(_797_), .C(_789_), .Y(_798_) );
NAND3X1 NAND3X1_8 ( .gnd(gnd), .vdd(vdd), .A(_787_), .B(_796_), .C(_798_), .Y(_799_) );
NAND3X1 NAND3X1_9 ( .gnd(gnd), .vdd(vdd), .A(_795_), .B(_786_), .C(_799_), .Y(_800_) );
AOI21X1 AOI21X1_2 ( .gnd(gnd), .vdd(vdd), .A(_759_), .B(_763_), .C(_766_), .Y(_801_) );
NAND3X1 NAND3X1_10 ( .gnd(gnd), .vdd(vdd), .A(_787_), .B(_794_), .C(_791_), .Y(_802_) );
NAND3X1 NAND3X1_11 ( .gnd(gnd), .vdd(vdd), .A(_788_), .B(_796_), .C(_798_), .Y(_803_) );
NAND3X1 NAND3X1_12 ( .gnd(gnd), .vdd(vdd), .A(_802_), .B(_803_), .C(_801_), .Y(_439_) );
NAND3X1 NAND3X1_13 ( .gnd(gnd), .vdd(vdd), .A(_785_), .B(_800_), .C(_439_), .Y(_440_) );
NAND3X1 NAND3X1_14 ( .gnd(gnd), .vdd(vdd), .A(_795_), .B(_799_), .C(_801_), .Y(_441_) );
NAND3X1 NAND3X1_15 ( .gnd(gnd), .vdd(vdd), .A(_802_), .B(_786_), .C(_803_), .Y(_442_) );
NAND3X1 NAND3X1_16 ( .gnd(gnd), .vdd(vdd), .A(_784_), .B(_442_), .C(_441_), .Y(_443_) );
AOI21X1 AOI21X1_3 ( .gnd(gnd), .vdd(vdd), .A(_440_), .B(_443_), .C(_783_), .Y(_444_) );
INVX1 INVX1_228 ( .gnd(gnd), .vdd(vdd), .A(_444_), .Y(_445_) );
NAND3X1 NAND3X1_17 ( .gnd(gnd), .vdd(vdd), .A(_783_), .B(_440_), .C(_443_), .Y(_446_) );
NAND3X1 NAND3X1_18 ( .gnd(gnd), .vdd(vdd), .A(MAC_salida_correcta_3_), .B(_446_), .C(_445_), .Y(_447_) );
INVX1 INVX1_229 ( .gnd(gnd), .vdd(vdd), .A(MAC_salida_correcta_3_), .Y(_448_) );
INVX1 INVX1_230 ( .gnd(gnd), .vdd(vdd), .A(_446_), .Y(_449_) );
OAI21X1 OAI21X1_188 ( .gnd(gnd), .vdd(vdd), .A(_444_), .B(_449_), .C(_448_), .Y(_450_) );
NAND2X1 NAND2X1_188 ( .gnd(gnd), .vdd(vdd), .A(_447_), .B(_450_), .Y(_451_) );
XOR2X1 XOR2X1_3 ( .gnd(gnd), .vdd(vdd), .A(_451_), .B(_782_), .Y(_452_) );
NAND3X1 NAND3X1_19 ( .gnd(gnd), .vdd(vdd), .A(MAC_clr_bF_buf3), .B(_446_), .C(_445_), .Y(_453_) );
OAI21X1 OAI21X1_189 ( .gnd(gnd), .vdd(vdd), .A(MAC_clr_bF_buf3), .B(_452_), .C(_453_), .Y(_438__3_) );
NAND2X1 NAND2X1_189 ( .gnd(gnd), .vdd(vdd), .A(MAC_Adder_1_), .B(MAC_ROM_4_), .Y(_454_) );
INVX1 INVX1_231 ( .gnd(gnd), .vdd(vdd), .A(MAC_ROM_4_), .Y(_455_) );
NAND2X1 NAND2X1_190 ( .gnd(gnd), .vdd(vdd), .A(MAC_Adder_1_), .B(MAC_ROM_3_), .Y(_456_) );
OAI21X1 OAI21X1_190 ( .gnd(gnd), .vdd(vdd), .A(_739_), .B(_455_), .C(_456_), .Y(_457_) );
OAI21X1 OAI21X1_191 ( .gnd(gnd), .vdd(vdd), .A(_784_), .B(_454_), .C(_457_), .Y(_458_) );
AOI22X1 AOI22X1_2 ( .gnd(gnd), .vdd(vdd), .A(MAC_ROM_0_bF_buf2_), .B(MAC_Adder_3_), .C(MAC_ROM_1_), .D(MAC_Adder_2_), .Y(_459_) );
OAI21X1 OAI21X1_192 ( .gnd(gnd), .vdd(vdd), .A(_787_), .B(_459_), .C(_791_), .Y(_460_) );
NAND2X1 NAND2X1_191 ( .gnd(gnd), .vdd(vdd), .A(MAC_Adder_2_), .B(MAC_ROM_2_), .Y(_461_) );
INVX1 INVX1_232 ( .gnd(gnd), .vdd(vdd), .A(_461_), .Y(_462_) );
AND2X2 AND2X2_6 ( .gnd(gnd), .vdd(vdd), .A(MAC_ROM_1_), .B(MAC_Adder_4_), .Y(_463_) );
NAND2X1 NAND2X1_192 ( .gnd(gnd), .vdd(vdd), .A(_790_), .B(_463_), .Y(_464_) );
NAND2X1 NAND2X1_193 ( .gnd(gnd), .vdd(vdd), .A(MAC_ROM_1_), .B(MAC_Adder_3_), .Y(_465_) );
NAND2X1 NAND2X1_194 ( .gnd(gnd), .vdd(vdd), .A(MAC_ROM_0_bF_buf1_), .B(MAC_Adder_4_), .Y(_466_) );
NAND2X1 NAND2X1_195 ( .gnd(gnd), .vdd(vdd), .A(_465_), .B(_466_), .Y(_467_) );
NAND3X1 NAND3X1_20 ( .gnd(gnd), .vdd(vdd), .A(_462_), .B(_467_), .C(_464_), .Y(_468_) );
NAND3X1 NAND3X1_21 ( .gnd(gnd), .vdd(vdd), .A(MAC_ROM_0_bF_buf0_), .B(MAC_Adder_4_), .C(_465_), .Y(_469_) );
AND2X2 AND2X2_7 ( .gnd(gnd), .vdd(vdd), .A(MAC_ROM_1_), .B(MAC_Adder_3_), .Y(_470_) );
NAND2X1 NAND2X1_196 ( .gnd(gnd), .vdd(vdd), .A(_466_), .B(_470_), .Y(_471_) );
NAND3X1 NAND3X1_22 ( .gnd(gnd), .vdd(vdd), .A(_461_), .B(_469_), .C(_471_), .Y(_472_) );
NAND3X1 NAND3X1_23 ( .gnd(gnd), .vdd(vdd), .A(_460_), .B(_468_), .C(_472_), .Y(_473_) );
AOI22X1 AOI22X1_3 ( .gnd(gnd), .vdd(vdd), .A(_760_), .B(_470_), .C(_794_), .D(_788_), .Y(_474_) );
NAND3X1 NAND3X1_24 ( .gnd(gnd), .vdd(vdd), .A(_461_), .B(_467_), .C(_464_), .Y(_475_) );
NAND3X1 NAND3X1_25 ( .gnd(gnd), .vdd(vdd), .A(_462_), .B(_469_), .C(_471_), .Y(_476_) );
NAND3X1 NAND3X1_26 ( .gnd(gnd), .vdd(vdd), .A(_476_), .B(_475_), .C(_474_), .Y(_477_) );
NAND3X1 NAND3X1_27 ( .gnd(gnd), .vdd(vdd), .A(_458_), .B(_473_), .C(_477_), .Y(_478_) );
INVX1 INVX1_233 ( .gnd(gnd), .vdd(vdd), .A(_458_), .Y(_479_) );
AOI21X1 AOI21X1_4 ( .gnd(gnd), .vdd(vdd), .A(_475_), .B(_476_), .C(_474_), .Y(_480_) );
AOI21X1 AOI21X1_5 ( .gnd(gnd), .vdd(vdd), .A(_468_), .B(_472_), .C(_460_), .Y(_481_) );
OAI21X1 OAI21X1_193 ( .gnd(gnd), .vdd(vdd), .A(_481_), .B(_480_), .C(_479_), .Y(_482_) );
AOI22X1 AOI22X1_4 ( .gnd(gnd), .vdd(vdd), .A(_800_), .B(_440_), .C(_482_), .D(_478_), .Y(_483_) );
AOI21X1 AOI21X1_6 ( .gnd(gnd), .vdd(vdd), .A(_799_), .B(_795_), .C(_786_), .Y(_484_) );
OAI21X1 OAI21X1_194 ( .gnd(gnd), .vdd(vdd), .A(_784_), .B(_484_), .C(_800_), .Y(_485_) );
NAND3X1 NAND3X1_28 ( .gnd(gnd), .vdd(vdd), .A(_479_), .B(_473_), .C(_477_), .Y(_486_) );
OAI21X1 OAI21X1_195 ( .gnd(gnd), .vdd(vdd), .A(_481_), .B(_480_), .C(_458_), .Y(_487_) );
AOI21X1 AOI21X1_7 ( .gnd(gnd), .vdd(vdd), .A(_486_), .B(_487_), .C(_485_), .Y(_488_) );
OAI21X1 OAI21X1_196 ( .gnd(gnd), .vdd(vdd), .A(_483_), .B(_488_), .C(_446_), .Y(_489_) );
NAND3X1 NAND3X1_29 ( .gnd(gnd), .vdd(vdd), .A(_486_), .B(_487_), .C(_485_), .Y(_490_) );
AOI21X1 AOI21X1_8 ( .gnd(gnd), .vdd(vdd), .A(_802_), .B(_803_), .C(_801_), .Y(_491_) );
AOI21X1 AOI21X1_9 ( .gnd(gnd), .vdd(vdd), .A(_785_), .B(_439_), .C(_491_), .Y(_492_) );
NAND3X1 NAND3X1_30 ( .gnd(gnd), .vdd(vdd), .A(_478_), .B(_482_), .C(_492_), .Y(_493_) );
NAND3X1 NAND3X1_31 ( .gnd(gnd), .vdd(vdd), .A(_490_), .B(_493_), .C(_449_), .Y(_494_) );
NAND2X1 NAND2X1_197 ( .gnd(gnd), .vdd(vdd), .A(_489_), .B(_494_), .Y(_495_) );
INVX1 INVX1_234 ( .gnd(gnd), .vdd(vdd), .A(_777_), .Y(_496_) );
AOI21X1 AOI21X1_10 ( .gnd(gnd), .vdd(vdd), .A(_496_), .B(_773_), .C(_776_), .Y(_497_) );
AOI21X1 AOI21X1_11 ( .gnd(gnd), .vdd(vdd), .A(_445_), .B(_446_), .C(MAC_salida_correcta_3_), .Y(_498_) );
OAI21X1 OAI21X1_197 ( .gnd(gnd), .vdd(vdd), .A(_497_), .B(_498_), .C(_447_), .Y(_499_) );
NAND3X1 NAND3X1_32 ( .gnd(gnd), .vdd(vdd), .A(MAC_salida_correcta_4_), .B(_489_), .C(_494_), .Y(_500_) );
INVX1 INVX1_235 ( .gnd(gnd), .vdd(vdd), .A(MAC_salida_correcta_4_), .Y(_501_) );
NAND2X1 NAND2X1_198 ( .gnd(gnd), .vdd(vdd), .A(_501_), .B(_495_), .Y(_502_) );
NAND3X1 NAND3X1_33 ( .gnd(gnd), .vdd(vdd), .A(_500_), .B(_499_), .C(_502_), .Y(_503_) );
INVX1 INVX1_236 ( .gnd(gnd), .vdd(vdd), .A(_447_), .Y(_504_) );
AOI21X1 AOI21X1_12 ( .gnd(gnd), .vdd(vdd), .A(_450_), .B(_782_), .C(_504_), .Y(_505_) );
INVX1 INVX1_237 ( .gnd(gnd), .vdd(vdd), .A(_500_), .Y(_506_) );
AOI21X1 AOI21X1_13 ( .gnd(gnd), .vdd(vdd), .A(_494_), .B(_489_), .C(MAC_salida_correcta_4_), .Y(_507_) );
OAI21X1 OAI21X1_198 ( .gnd(gnd), .vdd(vdd), .A(_507_), .B(_506_), .C(_505_), .Y(_508_) );
NAND3X1 NAND3X1_34 ( .gnd(gnd), .vdd(vdd), .A(_696_), .B(_503_), .C(_508_), .Y(_509_) );
OAI21X1 OAI21X1_199 ( .gnd(gnd), .vdd(vdd), .A(_696_), .B(_495_), .C(_509_), .Y(_438__4_) );
NOR3X1 NOR3X1_1 ( .gnd(gnd), .vdd(vdd), .A(_446_), .B(_483_), .C(_488_), .Y(_510_) );
AND2X2 AND2X2_8 ( .gnd(gnd), .vdd(vdd), .A(MAC_Adder_1_), .B(MAC_ROM_4_), .Y(_511_) );
NAND2X1 NAND2X1_199 ( .gnd(gnd), .vdd(vdd), .A(_511_), .B(_785_), .Y(_512_) );
INVX1 INVX1_238 ( .gnd(gnd), .vdd(vdd), .A(_512_), .Y(_513_) );
OAI21X1 OAI21X1_200 ( .gnd(gnd), .vdd(vdd), .A(_458_), .B(_481_), .C(_473_), .Y(_514_) );
NAND2X1 NAND2X1_200 ( .gnd(gnd), .vdd(vdd), .A(MAC_Adder_0_), .B(MAC_ROM_5_), .Y(_515_) );
INVX1 INVX1_239 ( .gnd(gnd), .vdd(vdd), .A(_515_), .Y(_516_) );
AND2X2 AND2X2_9 ( .gnd(gnd), .vdd(vdd), .A(MAC_Adder_2_), .B(MAC_ROM_3_), .Y(_517_) );
NAND2X1 NAND2X1_201 ( .gnd(gnd), .vdd(vdd), .A(_511_), .B(_517_), .Y(_518_) );
INVX1 INVX1_240 ( .gnd(gnd), .vdd(vdd), .A(MAC_ROM_3_), .Y(_519_) );
OAI21X1 OAI21X1_201 ( .gnd(gnd), .vdd(vdd), .A(_792_), .B(_519_), .C(_454_), .Y(_520_) );
NAND3X1 NAND3X1_35 ( .gnd(gnd), .vdd(vdd), .A(_520_), .B(_516_), .C(_518_), .Y(_521_) );
OAI21X1 OAI21X1_202 ( .gnd(gnd), .vdd(vdd), .A(_746_), .B(_455_), .C(_517_), .Y(_522_) );
OAI21X1 OAI21X1_203 ( .gnd(gnd), .vdd(vdd), .A(_792_), .B(_519_), .C(_511_), .Y(_523_) );
NAND3X1 NAND3X1_36 ( .gnd(gnd), .vdd(vdd), .A(_515_), .B(_522_), .C(_523_), .Y(_524_) );
AOI22X1 AOI22X1_5 ( .gnd(gnd), .vdd(vdd), .A(_790_), .B(_463_), .C(_467_), .D(_462_), .Y(_525_) );
NAND2X1 NAND2X1_202 ( .gnd(gnd), .vdd(vdd), .A(MAC_ROM_2_), .B(MAC_Adder_3_), .Y(_526_) );
INVX1 INVX1_241 ( .gnd(gnd), .vdd(vdd), .A(_526_), .Y(_527_) );
AND2X2 AND2X2_10 ( .gnd(gnd), .vdd(vdd), .A(MAC_ROM_0_bF_buf3_), .B(MAC_Adder_5_), .Y(_528_) );
NAND2X1 NAND2X1_203 ( .gnd(gnd), .vdd(vdd), .A(_463_), .B(_528_), .Y(_529_) );
INVX1 INVX1_242 ( .gnd(gnd), .vdd(vdd), .A(MAC_Adder_5_), .Y(_530_) );
NAND2X1 NAND2X1_204 ( .gnd(gnd), .vdd(vdd), .A(MAC_ROM_1_), .B(MAC_Adder_4_), .Y(_531_) );
OAI21X1 OAI21X1_204 ( .gnd(gnd), .vdd(vdd), .A(_728_), .B(_530_), .C(_531_), .Y(_532_) );
NAND3X1 NAND3X1_37 ( .gnd(gnd), .vdd(vdd), .A(_527_), .B(_532_), .C(_529_), .Y(_533_) );
NAND3X1 NAND3X1_38 ( .gnd(gnd), .vdd(vdd), .A(MAC_ROM_0_bF_buf2_), .B(MAC_Adder_5_), .C(_531_), .Y(_534_) );
NAND2X1 NAND2X1_205 ( .gnd(gnd), .vdd(vdd), .A(MAC_ROM_0_bF_buf1_), .B(MAC_Adder_5_), .Y(_535_) );
NAND3X1 NAND3X1_39 ( .gnd(gnd), .vdd(vdd), .A(MAC_ROM_1_), .B(MAC_Adder_4_), .C(_535_), .Y(_536_) );
NAND3X1 NAND3X1_40 ( .gnd(gnd), .vdd(vdd), .A(_526_), .B(_534_), .C(_536_), .Y(_537_) );
NAND3X1 NAND3X1_41 ( .gnd(gnd), .vdd(vdd), .A(_525_), .B(_537_), .C(_533_), .Y(_538_) );
AOI22X1 AOI22X1_6 ( .gnd(gnd), .vdd(vdd), .A(MAC_ROM_0_bF_buf0_), .B(MAC_Adder_4_), .C(MAC_ROM_1_), .D(MAC_Adder_3_), .Y(_539_) );
OAI22X1 OAI22X1_2 ( .gnd(gnd), .vdd(vdd), .A(_793_), .B(_531_), .C(_461_), .D(_539_), .Y(_540_) );
NAND3X1 NAND3X1_42 ( .gnd(gnd), .vdd(vdd), .A(_526_), .B(_532_), .C(_529_), .Y(_541_) );
NAND3X1 NAND3X1_43 ( .gnd(gnd), .vdd(vdd), .A(_527_), .B(_534_), .C(_536_), .Y(_542_) );
NAND3X1 NAND3X1_44 ( .gnd(gnd), .vdd(vdd), .A(_540_), .B(_542_), .C(_541_), .Y(_543_) );
AOI22X1 AOI22X1_7 ( .gnd(gnd), .vdd(vdd), .A(_521_), .B(_524_), .C(_538_), .D(_543_), .Y(_544_) );
NAND3X1 NAND3X1_45 ( .gnd(gnd), .vdd(vdd), .A(_515_), .B(_520_), .C(_518_), .Y(_545_) );
NAND3X1 NAND3X1_46 ( .gnd(gnd), .vdd(vdd), .A(_516_), .B(_522_), .C(_523_), .Y(_546_) );
NAND3X1 NAND3X1_47 ( .gnd(gnd), .vdd(vdd), .A(_540_), .B(_537_), .C(_533_), .Y(_547_) );
NAND3X1 NAND3X1_48 ( .gnd(gnd), .vdd(vdd), .A(_525_), .B(_542_), .C(_541_), .Y(_548_) );
AOI22X1 AOI22X1_8 ( .gnd(gnd), .vdd(vdd), .A(_545_), .B(_546_), .C(_547_), .D(_548_), .Y(_549_) );
OAI21X1 OAI21X1_205 ( .gnd(gnd), .vdd(vdd), .A(_544_), .B(_549_), .C(_514_), .Y(_550_) );
AOI21X1 AOI21X1_14 ( .gnd(gnd), .vdd(vdd), .A(_479_), .B(_477_), .C(_480_), .Y(_551_) );
NAND2X1 NAND2X1_206 ( .gnd(gnd), .vdd(vdd), .A(_521_), .B(_524_), .Y(_552_) );
AOI21X1 AOI21X1_15 ( .gnd(gnd), .vdd(vdd), .A(_538_), .B(_543_), .C(_552_), .Y(_553_) );
NAND2X1 NAND2X1_207 ( .gnd(gnd), .vdd(vdd), .A(_545_), .B(_546_), .Y(_554_) );
AOI21X1 AOI21X1_16 ( .gnd(gnd), .vdd(vdd), .A(_547_), .B(_548_), .C(_554_), .Y(_555_) );
OAI21X1 OAI21X1_206 ( .gnd(gnd), .vdd(vdd), .A(_555_), .B(_553_), .C(_551_), .Y(_556_) );
NAND3X1 NAND3X1_49 ( .gnd(gnd), .vdd(vdd), .A(_513_), .B(_550_), .C(_556_), .Y(_557_) );
OAI21X1 OAI21X1_207 ( .gnd(gnd), .vdd(vdd), .A(_544_), .B(_549_), .C(_551_), .Y(_558_) );
OAI21X1 OAI21X1_208 ( .gnd(gnd), .vdd(vdd), .A(_555_), .B(_553_), .C(_514_), .Y(_559_) );
NAND3X1 NAND3X1_50 ( .gnd(gnd), .vdd(vdd), .A(_512_), .B(_558_), .C(_559_), .Y(_560_) );
NAND3X1 NAND3X1_51 ( .gnd(gnd), .vdd(vdd), .A(_483_), .B(_557_), .C(_560_), .Y(_561_) );
NAND3X1 NAND3X1_52 ( .gnd(gnd), .vdd(vdd), .A(_512_), .B(_550_), .C(_556_), .Y(_562_) );
NAND3X1 NAND3X1_53 ( .gnd(gnd), .vdd(vdd), .A(_513_), .B(_558_), .C(_559_), .Y(_563_) );
NAND3X1 NAND3X1_54 ( .gnd(gnd), .vdd(vdd), .A(_490_), .B(_562_), .C(_563_), .Y(_564_) );
NAND3X1 NAND3X1_55 ( .gnd(gnd), .vdd(vdd), .A(_510_), .B(_561_), .C(_564_), .Y(_565_) );
NAND3X1 NAND3X1_56 ( .gnd(gnd), .vdd(vdd), .A(_490_), .B(_557_), .C(_560_), .Y(_566_) );
NAND3X1 NAND3X1_57 ( .gnd(gnd), .vdd(vdd), .A(_483_), .B(_562_), .C(_563_), .Y(_567_) );
NAND3X1 NAND3X1_58 ( .gnd(gnd), .vdd(vdd), .A(_494_), .B(_566_), .C(_567_), .Y(_568_) );
NAND2X1 NAND2X1_208 ( .gnd(gnd), .vdd(vdd), .A(_565_), .B(_568_), .Y(_569_) );
OAI21X1 OAI21X1_209 ( .gnd(gnd), .vdd(vdd), .A(_507_), .B(_505_), .C(_500_), .Y(_570_) );
NAND3X1 NAND3X1_59 ( .gnd(gnd), .vdd(vdd), .A(MAC_salida_correcta_5_), .B(_565_), .C(_568_), .Y(_571_) );
INVX1 INVX1_243 ( .gnd(gnd), .vdd(vdd), .A(MAC_salida_correcta_5_), .Y(_572_) );
NAND2X1 NAND2X1_209 ( .gnd(gnd), .vdd(vdd), .A(_572_), .B(_569_), .Y(_573_) );
NAND3X1 NAND3X1_60 ( .gnd(gnd), .vdd(vdd), .A(_571_), .B(_573_), .C(_570_), .Y(_574_) );
AOI21X1 AOI21X1_17 ( .gnd(gnd), .vdd(vdd), .A(_499_), .B(_502_), .C(_506_), .Y(_575_) );
INVX1 INVX1_244 ( .gnd(gnd), .vdd(vdd), .A(_571_), .Y(_576_) );
AOI21X1 AOI21X1_18 ( .gnd(gnd), .vdd(vdd), .A(_565_), .B(_568_), .C(MAC_salida_correcta_5_), .Y(_577_) );
OAI21X1 OAI21X1_210 ( .gnd(gnd), .vdd(vdd), .A(_577_), .B(_576_), .C(_575_), .Y(_578_) );
NAND3X1 NAND3X1_61 ( .gnd(gnd), .vdd(vdd), .A(_696_), .B(_574_), .C(_578_), .Y(_579_) );
OAI21X1 OAI21X1_211 ( .gnd(gnd), .vdd(vdd), .A(_696_), .B(_569_), .C(_579_), .Y(_438__5_) );
AOI21X1 AOI21X1_19 ( .gnd(gnd), .vdd(vdd), .A(_566_), .B(_567_), .C(_494_), .Y(_580_) );
AOI21X1 AOI21X1_20 ( .gnd(gnd), .vdd(vdd), .A(_563_), .B(_562_), .C(_490_), .Y(_581_) );
NAND3X1 NAND3X1_62 ( .gnd(gnd), .vdd(vdd), .A(_547_), .B(_548_), .C(_554_), .Y(_582_) );
AOI21X1 AOI21X1_21 ( .gnd(gnd), .vdd(vdd), .A(_541_), .B(_542_), .C(_525_), .Y(_583_) );
AOI21X1 AOI21X1_22 ( .gnd(gnd), .vdd(vdd), .A(_533_), .B(_537_), .C(_540_), .Y(_584_) );
OAI21X1 OAI21X1_212 ( .gnd(gnd), .vdd(vdd), .A(_583_), .B(_584_), .C(_552_), .Y(_585_) );
AOI21X1 AOI21X1_23 ( .gnd(gnd), .vdd(vdd), .A(_585_), .B(_582_), .C(_514_), .Y(_586_) );
OAI21X1 OAI21X1_213 ( .gnd(gnd), .vdd(vdd), .A(_512_), .B(_586_), .C(_550_), .Y(_587_) );
AND2X2 AND2X2_11 ( .gnd(gnd), .vdd(vdd), .A(MAC_Adder_0_), .B(MAC_ROM_6_), .Y(_588_) );
NAND2X1 NAND2X1_210 ( .gnd(gnd), .vdd(vdd), .A(MAC_Adder_2_), .B(MAC_ROM_4_), .Y(_589_) );
OAI21X1 OAI21X1_214 ( .gnd(gnd), .vdd(vdd), .A(_456_), .B(_589_), .C(_521_), .Y(_590_) );
XNOR2X1 XNOR2X1_1 ( .gnd(gnd), .vdd(vdd), .A(_590_), .B(_588_), .Y(_591_) );
INVX1 INVX1_245 ( .gnd(gnd), .vdd(vdd), .A(_591_), .Y(_592_) );
OAI21X1 OAI21X1_215 ( .gnd(gnd), .vdd(vdd), .A(_552_), .B(_584_), .C(_547_), .Y(_593_) );
INVX1 INVX1_246 ( .gnd(gnd), .vdd(vdd), .A(MAC_ROM_5_), .Y(_594_) );
NOR2X1 NOR2X1_7 ( .gnd(gnd), .vdd(vdd), .A(_746_), .B(_594_), .Y(_595_) );
NAND2X1 NAND2X1_211 ( .gnd(gnd), .vdd(vdd), .A(MAC_Adder_3_), .B(MAC_ROM_3_), .Y(_596_) );
XOR2X1 XOR2X1_4 ( .gnd(gnd), .vdd(vdd), .A(_589_), .B(_596_), .Y(_597_) );
NAND2X1 NAND2X1_212 ( .gnd(gnd), .vdd(vdd), .A(_595_), .B(_597_), .Y(_598_) );
INVX1 INVX1_247 ( .gnd(gnd), .vdd(vdd), .A(_517_), .Y(_599_) );
NAND2X1 NAND2X1_213 ( .gnd(gnd), .vdd(vdd), .A(MAC_Adder_3_), .B(MAC_ROM_4_), .Y(_600_) );
OAI21X1 OAI21X1_216 ( .gnd(gnd), .vdd(vdd), .A(_797_), .B(_519_), .C(_589_), .Y(_601_) );
OAI21X1 OAI21X1_217 ( .gnd(gnd), .vdd(vdd), .A(_600_), .B(_599_), .C(_601_), .Y(_602_) );
OAI21X1 OAI21X1_218 ( .gnd(gnd), .vdd(vdd), .A(_746_), .B(_594_), .C(_602_), .Y(_603_) );
NOR2X1 NOR2X1_8 ( .gnd(gnd), .vdd(vdd), .A(_531_), .B(_535_), .Y(_604_) );
AOI21X1 AOI21X1_24 ( .gnd(gnd), .vdd(vdd), .A(_527_), .B(_532_), .C(_604_), .Y(_605_) );
NAND2X1 NAND2X1_214 ( .gnd(gnd), .vdd(vdd), .A(MAC_ROM_2_), .B(MAC_Adder_4_), .Y(_606_) );
INVX1 INVX1_248 ( .gnd(gnd), .vdd(vdd), .A(_606_), .Y(_607_) );
NAND3X1 NAND3X1_63 ( .gnd(gnd), .vdd(vdd), .A(MAC_ROM_1_), .B(MAC_Adder_6_), .C(_528_), .Y(_608_) );
AOI22X1 AOI22X1_9 ( .gnd(gnd), .vdd(vdd), .A(MAC_ROM_0_bF_buf3_), .B(MAC_Adder_6_), .C(MAC_ROM_1_), .D(MAC_Adder_5_), .Y(_609_) );
INVX1 INVX1_249 ( .gnd(gnd), .vdd(vdd), .A(_609_), .Y(_610_) );
NAND3X1 NAND3X1_64 ( .gnd(gnd), .vdd(vdd), .A(_610_), .B(_607_), .C(_608_), .Y(_611_) );
NAND2X1 NAND2X1_215 ( .gnd(gnd), .vdd(vdd), .A(MAC_ROM_1_), .B(MAC_Adder_6_), .Y(_612_) );
NOR2X1 NOR2X1_9 ( .gnd(gnd), .vdd(vdd), .A(_535_), .B(_612_), .Y(_613_) );
OAI21X1 OAI21X1_219 ( .gnd(gnd), .vdd(vdd), .A(_609_), .B(_613_), .C(_606_), .Y(_614_) );
NAND3X1 NAND3X1_65 ( .gnd(gnd), .vdd(vdd), .A(_611_), .B(_614_), .C(_605_), .Y(_615_) );
AND2X2 AND2X2_12 ( .gnd(gnd), .vdd(vdd), .A(_531_), .B(_535_), .Y(_616_) );
OAI21X1 OAI21X1_220 ( .gnd(gnd), .vdd(vdd), .A(_526_), .B(_616_), .C(_529_), .Y(_617_) );
NAND3X1 NAND3X1_66 ( .gnd(gnd), .vdd(vdd), .A(_606_), .B(_610_), .C(_608_), .Y(_618_) );
OAI21X1 OAI21X1_221 ( .gnd(gnd), .vdd(vdd), .A(_609_), .B(_613_), .C(_607_), .Y(_619_) );
NAND3X1 NAND3X1_67 ( .gnd(gnd), .vdd(vdd), .A(_618_), .B(_619_), .C(_617_), .Y(_620_) );
AOI22X1 AOI22X1_10 ( .gnd(gnd), .vdd(vdd), .A(_598_), .B(_603_), .C(_615_), .D(_620_), .Y(_621_) );
OAI21X1 OAI21X1_222 ( .gnd(gnd), .vdd(vdd), .A(_746_), .B(_594_), .C(_597_), .Y(_622_) );
NAND2X1 NAND2X1_216 ( .gnd(gnd), .vdd(vdd), .A(_595_), .B(_602_), .Y(_623_) );
NAND3X1 NAND3X1_68 ( .gnd(gnd), .vdd(vdd), .A(_611_), .B(_614_), .C(_617_), .Y(_624_) );
NAND3X1 NAND3X1_69 ( .gnd(gnd), .vdd(vdd), .A(_618_), .B(_619_), .C(_605_), .Y(_625_) );
AOI22X1 AOI22X1_11 ( .gnd(gnd), .vdd(vdd), .A(_622_), .B(_623_), .C(_625_), .D(_624_), .Y(_626_) );
OAI21X1 OAI21X1_223 ( .gnd(gnd), .vdd(vdd), .A(_621_), .B(_626_), .C(_593_), .Y(_627_) );
AOI21X1 AOI21X1_25 ( .gnd(gnd), .vdd(vdd), .A(_554_), .B(_548_), .C(_583_), .Y(_628_) );
AOI22X1 AOI22X1_12 ( .gnd(gnd), .vdd(vdd), .A(_622_), .B(_623_), .C(_615_), .D(_620_), .Y(_629_) );
AOI22X1 AOI22X1_13 ( .gnd(gnd), .vdd(vdd), .A(_598_), .B(_603_), .C(_625_), .D(_624_), .Y(_630_) );
OAI21X1 OAI21X1_224 ( .gnd(gnd), .vdd(vdd), .A(_629_), .B(_630_), .C(_628_), .Y(_631_) );
NAND3X1 NAND3X1_70 ( .gnd(gnd), .vdd(vdd), .A(_627_), .B(_592_), .C(_631_), .Y(_632_) );
OAI21X1 OAI21X1_225 ( .gnd(gnd), .vdd(vdd), .A(_621_), .B(_626_), .C(_628_), .Y(_633_) );
OAI21X1 OAI21X1_226 ( .gnd(gnd), .vdd(vdd), .A(_629_), .B(_630_), .C(_593_), .Y(_634_) );
NAND3X1 NAND3X1_71 ( .gnd(gnd), .vdd(vdd), .A(_591_), .B(_633_), .C(_634_), .Y(_635_) );
NAND3X1 NAND3X1_72 ( .gnd(gnd), .vdd(vdd), .A(_635_), .B(_632_), .C(_587_), .Y(_636_) );
NAND3X1 NAND3X1_73 ( .gnd(gnd), .vdd(vdd), .A(_547_), .B(_552_), .C(_548_), .Y(_637_) );
OAI21X1 OAI21X1_227 ( .gnd(gnd), .vdd(vdd), .A(_583_), .B(_584_), .C(_554_), .Y(_638_) );
AOI21X1 AOI21X1_26 ( .gnd(gnd), .vdd(vdd), .A(_638_), .B(_637_), .C(_551_), .Y(_639_) );
AOI21X1 AOI21X1_27 ( .gnd(gnd), .vdd(vdd), .A(_513_), .B(_556_), .C(_639_), .Y(_640_) );
NAND3X1 NAND3X1_74 ( .gnd(gnd), .vdd(vdd), .A(_591_), .B(_627_), .C(_631_), .Y(_641_) );
NAND3X1 NAND3X1_75 ( .gnd(gnd), .vdd(vdd), .A(_633_), .B(_592_), .C(_634_), .Y(_642_) );
NAND3X1 NAND3X1_76 ( .gnd(gnd), .vdd(vdd), .A(_641_), .B(_642_), .C(_640_), .Y(_643_) );
NAND3X1 NAND3X1_77 ( .gnd(gnd), .vdd(vdd), .A(_581_), .B(_643_), .C(_636_), .Y(_644_) );
NAND3X1 NAND3X1_78 ( .gnd(gnd), .vdd(vdd), .A(_635_), .B(_632_), .C(_640_), .Y(_645_) );
NAND3X1 NAND3X1_79 ( .gnd(gnd), .vdd(vdd), .A(_641_), .B(_642_), .C(_587_), .Y(_646_) );
NAND3X1 NAND3X1_80 ( .gnd(gnd), .vdd(vdd), .A(_561_), .B(_645_), .C(_646_), .Y(_647_) );
NAND3X1 NAND3X1_81 ( .gnd(gnd), .vdd(vdd), .A(_580_), .B(_644_), .C(_647_), .Y(_648_) );
NAND3X1 NAND3X1_82 ( .gnd(gnd), .vdd(vdd), .A(_561_), .B(_643_), .C(_636_), .Y(_649_) );
NAND3X1 NAND3X1_83 ( .gnd(gnd), .vdd(vdd), .A(_581_), .B(_645_), .C(_646_), .Y(_650_) );
NAND3X1 NAND3X1_84 ( .gnd(gnd), .vdd(vdd), .A(_565_), .B(_649_), .C(_650_), .Y(_651_) );
NAND2X1 NAND2X1_217 ( .gnd(gnd), .vdd(vdd), .A(_648_), .B(_651_), .Y(_652_) );
OAI21X1 OAI21X1_228 ( .gnd(gnd), .vdd(vdd), .A(_577_), .B(_575_), .C(_571_), .Y(_653_) );
NAND3X1 NAND3X1_85 ( .gnd(gnd), .vdd(vdd), .A(MAC_salida_correcta_6_), .B(_648_), .C(_651_), .Y(_654_) );
INVX1 INVX1_250 ( .gnd(gnd), .vdd(vdd), .A(MAC_salida_correcta_6_), .Y(_655_) );
NAND3X1 NAND3X1_86 ( .gnd(gnd), .vdd(vdd), .A(_565_), .B(_644_), .C(_647_), .Y(_656_) );
NAND3X1 NAND3X1_87 ( .gnd(gnd), .vdd(vdd), .A(_580_), .B(_649_), .C(_650_), .Y(_657_) );
NAND3X1 NAND3X1_88 ( .gnd(gnd), .vdd(vdd), .A(_655_), .B(_656_), .C(_657_), .Y(_658_) );
AOI21X1 AOI21X1_28 ( .gnd(gnd), .vdd(vdd), .A(_654_), .B(_658_), .C(_653_), .Y(_659_) );
AOI21X1 AOI21X1_29 ( .gnd(gnd), .vdd(vdd), .A(_570_), .B(_573_), .C(_576_), .Y(_660_) );
NAND2X1 NAND2X1_218 ( .gnd(gnd), .vdd(vdd), .A(_654_), .B(_658_), .Y(_661_) );
OAI21X1 OAI21X1_229 ( .gnd(gnd), .vdd(vdd), .A(_660_), .B(_661_), .C(_696_), .Y(_662_) );
OAI22X1 OAI22X1_3 ( .gnd(gnd), .vdd(vdd), .A(_696_), .B(_652_), .C(_659_), .D(_662_), .Y(_438__6_) );
NAND2X1 NAND2X1_219 ( .gnd(gnd), .vdd(vdd), .A(_644_), .B(_648_), .Y(_663_) );
INVX1 INVX1_251 ( .gnd(gnd), .vdd(vdd), .A(_663_), .Y(_664_) );
INVX1 INVX1_252 ( .gnd(gnd), .vdd(vdd), .A(_636_), .Y(_665_) );
NAND2X1 NAND2X1_220 ( .gnd(gnd), .vdd(vdd), .A(_588_), .B(_590_), .Y(_666_) );
INVX1 INVX1_253 ( .gnd(gnd), .vdd(vdd), .A(_666_), .Y(_667_) );
NAND2X1 NAND2X1_221 ( .gnd(gnd), .vdd(vdd), .A(_627_), .B(_632_), .Y(_668_) );
OAI21X1 OAI21X1_230 ( .gnd(gnd), .vdd(vdd), .A(_599_), .B(_600_), .C(_598_), .Y(_669_) );
NAND2X1 NAND2X1_222 ( .gnd(gnd), .vdd(vdd), .A(MAC_Adder_0_), .B(MAC_ROM_7_), .Y(_670_) );
NAND2X1 NAND2X1_223 ( .gnd(gnd), .vdd(vdd), .A(MAC_Adder_1_), .B(MAC_ROM_6_), .Y(_671_) );
XOR2X1 XOR2X1_5 ( .gnd(gnd), .vdd(vdd), .A(_670_), .B(_671_), .Y(_672_) );
XOR2X1 XOR2X1_6 ( .gnd(gnd), .vdd(vdd), .A(_669_), .B(_672_), .Y(_673_) );
INVX1 INVX1_254 ( .gnd(gnd), .vdd(vdd), .A(_673_), .Y(_674_) );
INVX1 INVX1_255 ( .gnd(gnd), .vdd(vdd), .A(_624_), .Y(_675_) );
OR2X2 OR2X2_2 ( .gnd(gnd), .vdd(vdd), .A(_629_), .B(_675_), .Y(_676_) );
INVX1 INVX1_256 ( .gnd(gnd), .vdd(vdd), .A(MAC_ROM_2_), .Y(_677_) );
NOR2X1 NOR2X1_10 ( .gnd(gnd), .vdd(vdd), .A(_677_), .B(_530_), .Y(_678_) );
NAND2X1 NAND2X1_224 ( .gnd(gnd), .vdd(vdd), .A(MAC_ROM_0_bF_buf2_), .B(MAC_Adder_7_), .Y(_679_) );
XNOR2X1 XNOR2X1_2 ( .gnd(gnd), .vdd(vdd), .A(_612_), .B(_679_), .Y(_680_) );
INVX1 INVX1_257 ( .gnd(gnd), .vdd(vdd), .A(_680_), .Y(_681_) );
NAND2X1 NAND2X1_225 ( .gnd(gnd), .vdd(vdd), .A(_678_), .B(_681_), .Y(_682_) );
OAI21X1 OAI21X1_231 ( .gnd(gnd), .vdd(vdd), .A(_677_), .B(_530_), .C(_680_), .Y(_683_) );
OAI21X1 OAI21X1_232 ( .gnd(gnd), .vdd(vdd), .A(_606_), .B(_609_), .C(_608_), .Y(_684_) );
INVX1 INVX1_258 ( .gnd(gnd), .vdd(vdd), .A(_684_), .Y(_686_) );
NAND3X1 NAND3X1_89 ( .gnd(gnd), .vdd(vdd), .A(_683_), .B(_686_), .C(_682_), .Y(_687_) );
NAND2X1 NAND2X1_226 ( .gnd(gnd), .vdd(vdd), .A(_678_), .B(_680_), .Y(_688_) );
OAI21X1 OAI21X1_233 ( .gnd(gnd), .vdd(vdd), .A(_677_), .B(_530_), .C(_681_), .Y(_689_) );
NAND3X1 NAND3X1_90 ( .gnd(gnd), .vdd(vdd), .A(_684_), .B(_688_), .C(_689_), .Y(_690_) );
NAND2X1 NAND2X1_227 ( .gnd(gnd), .vdd(vdd), .A(MAC_ROM_3_), .B(MAC_Adder_4_), .Y(_691_) );
XNOR2X1 XNOR2X1_3 ( .gnd(gnd), .vdd(vdd), .A(_600_), .B(_691_), .Y(_692_) );
NAND2X1 NAND2X1_228 ( .gnd(gnd), .vdd(vdd), .A(MAC_Adder_2_), .B(MAC_ROM_5_), .Y(_693_) );
XOR2X1 XOR2X1_7 ( .gnd(gnd), .vdd(vdd), .A(_692_), .B(_693_), .Y(_694_) );
INVX1 INVX1_259 ( .gnd(gnd), .vdd(vdd), .A(_694_), .Y(_695_) );
NAND3X1 NAND3X1_91 ( .gnd(gnd), .vdd(vdd), .A(_687_), .B(_690_), .C(_695_), .Y(_697_) );
NAND3X1 NAND3X1_92 ( .gnd(gnd), .vdd(vdd), .A(_683_), .B(_684_), .C(_682_), .Y(_698_) );
NAND3X1 NAND3X1_93 ( .gnd(gnd), .vdd(vdd), .A(_686_), .B(_688_), .C(_689_), .Y(_699_) );
NAND3X1 NAND3X1_94 ( .gnd(gnd), .vdd(vdd), .A(_694_), .B(_698_), .C(_699_), .Y(_700_) );
NAND3X1 NAND3X1_95 ( .gnd(gnd), .vdd(vdd), .A(_700_), .B(_697_), .C(_676_), .Y(_701_) );
NOR2X1 NOR2X1_11 ( .gnd(gnd), .vdd(vdd), .A(_675_), .B(_629_), .Y(_702_) );
NAND3X1 NAND3X1_96 ( .gnd(gnd), .vdd(vdd), .A(_698_), .B(_699_), .C(_695_), .Y(_703_) );
NAND3X1 NAND3X1_97 ( .gnd(gnd), .vdd(vdd), .A(_694_), .B(_687_), .C(_690_), .Y(_704_) );
NAND3X1 NAND3X1_98 ( .gnd(gnd), .vdd(vdd), .A(_702_), .B(_704_), .C(_703_), .Y(_705_) );
AOI21X1 AOI21X1_30 ( .gnd(gnd), .vdd(vdd), .A(_701_), .B(_705_), .C(_674_), .Y(_706_) );
NAND3X1 NAND3X1_99 ( .gnd(gnd), .vdd(vdd), .A(_702_), .B(_700_), .C(_697_), .Y(_708_) );
NAND3X1 NAND3X1_100 ( .gnd(gnd), .vdd(vdd), .A(_704_), .B(_703_), .C(_676_), .Y(_709_) );
AOI21X1 AOI21X1_31 ( .gnd(gnd), .vdd(vdd), .A(_709_), .B(_708_), .C(_673_), .Y(_710_) );
OAI21X1 OAI21X1_234 ( .gnd(gnd), .vdd(vdd), .A(_706_), .B(_710_), .C(_668_), .Y(_711_) );
INVX1 INVX1_260 ( .gnd(gnd), .vdd(vdd), .A(_668_), .Y(_712_) );
NAND3X1 NAND3X1_101 ( .gnd(gnd), .vdd(vdd), .A(_673_), .B(_708_), .C(_709_), .Y(_713_) );
NAND3X1 NAND3X1_102 ( .gnd(gnd), .vdd(vdd), .A(_674_), .B(_705_), .C(_701_), .Y(_714_) );
NAND3X1 NAND3X1_103 ( .gnd(gnd), .vdd(vdd), .A(_713_), .B(_714_), .C(_712_), .Y(_715_) );
AOI21X1 AOI21X1_32 ( .gnd(gnd), .vdd(vdd), .A(_715_), .B(_711_), .C(_667_), .Y(_716_) );
NAND3X1 NAND3X1_104 ( .gnd(gnd), .vdd(vdd), .A(_668_), .B(_713_), .C(_714_), .Y(_717_) );
OAI21X1 OAI21X1_235 ( .gnd(gnd), .vdd(vdd), .A(_706_), .B(_710_), .C(_712_), .Y(_718_) );
AOI21X1 AOI21X1_33 ( .gnd(gnd), .vdd(vdd), .A(_718_), .B(_717_), .C(_666_), .Y(_719_) );
OAI21X1 OAI21X1_236 ( .gnd(gnd), .vdd(vdd), .A(_719_), .B(_716_), .C(_665_), .Y(_720_) );
NAND3X1 NAND3X1_105 ( .gnd(gnd), .vdd(vdd), .A(_666_), .B(_717_), .C(_718_), .Y(_721_) );
NAND3X1 NAND3X1_106 ( .gnd(gnd), .vdd(vdd), .A(_667_), .B(_711_), .C(_715_), .Y(_722_) );
NAND3X1 NAND3X1_107 ( .gnd(gnd), .vdd(vdd), .A(_636_), .B(_721_), .C(_722_), .Y(_723_) );
NAND3X1 NAND3X1_108 ( .gnd(gnd), .vdd(vdd), .A(_664_), .B(_723_), .C(_720_), .Y(_724_) );
NAND2X1 NAND2X1_229 ( .gnd(gnd), .vdd(vdd), .A(_711_), .B(_715_), .Y(_725_) );
XOR2X1 XOR2X1_8 ( .gnd(gnd), .vdd(vdd), .A(_636_), .B(_667_), .Y(_726_) );
OR2X2 OR2X2_3 ( .gnd(gnd), .vdd(vdd), .A(_725_), .B(_726_), .Y(_727_) );
NAND2X1 NAND2X1_230 ( .gnd(gnd), .vdd(vdd), .A(_726_), .B(_725_), .Y(_729_) );
NAND3X1 NAND3X1_109 ( .gnd(gnd), .vdd(vdd), .A(_663_), .B(_729_), .C(_727_), .Y(_730_) );
NAND2X1 NAND2X1_231 ( .gnd(gnd), .vdd(vdd), .A(_730_), .B(_724_), .Y(_731_) );
INVX1 INVX1_261 ( .gnd(gnd), .vdd(vdd), .A(MAC_salida_correcta_7_), .Y(_732_) );
AOI21X1 AOI21X1_34 ( .gnd(gnd), .vdd(vdd), .A(_656_), .B(_657_), .C(_655_), .Y(_733_) );
AOI21X1 AOI21X1_35 ( .gnd(gnd), .vdd(vdd), .A(_653_), .B(_658_), .C(_733_), .Y(_734_) );
NAND2X1 NAND2X1_232 ( .gnd(gnd), .vdd(vdd), .A(_732_), .B(_734_), .Y(_735_) );
AOI21X1 AOI21X1_36 ( .gnd(gnd), .vdd(vdd), .A(_648_), .B(_651_), .C(MAC_salida_correcta_6_), .Y(_736_) );
OAI21X1 OAI21X1_237 ( .gnd(gnd), .vdd(vdd), .A(_736_), .B(_660_), .C(_654_), .Y(_737_) );
AOI21X1 AOI21X1_37 ( .gnd(gnd), .vdd(vdd), .A(_737_), .B(MAC_salida_correcta_7_), .C(MAC_clr_bF_buf0), .Y(_738_) );
NAND3X1 NAND3X1_110 ( .gnd(gnd), .vdd(vdd), .A(_731_), .B(_735_), .C(_738_), .Y(_740_) );
AOI21X1 AOI21X1_38 ( .gnd(gnd), .vdd(vdd), .A(_727_), .B(_729_), .C(_664_), .Y(_741_) );
AOI21X1 AOI21X1_39 ( .gnd(gnd), .vdd(vdd), .A(_720_), .B(_723_), .C(_663_), .Y(_742_) );
AND2X2 AND2X2_13 ( .gnd(gnd), .vdd(vdd), .A(_734_), .B(_732_), .Y(_743_) );
OAI21X1 OAI21X1_238 ( .gnd(gnd), .vdd(vdd), .A(_732_), .B(_734_), .C(_696_), .Y(_744_) );
OAI22X1 OAI22X1_4 ( .gnd(gnd), .vdd(vdd), .A(_741_), .B(_742_), .C(_744_), .D(_743_), .Y(_745_) );
NAND2X1 NAND2X1_233 ( .gnd(gnd), .vdd(vdd), .A(_745_), .B(_740_), .Y(_438__7_) );
DFFPOSX1 DFFPOSX1_2 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf5), .D(_438__0_), .Q(MAC_salida_correcta_0_) );
DFFPOSX1 DFFPOSX1_3 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf5), .D(_438__1_), .Q(MAC_salida_correcta_1_) );
DFFPOSX1 DFFPOSX1_4 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf7), .D(_438__2_), .Q(MAC_salida_correcta_2_) );
DFFPOSX1 DFFPOSX1_5 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf3), .D(_438__3_), .Q(MAC_salida_correcta_3_) );
DFFPOSX1 DFFPOSX1_6 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf7), .D(_438__4_), .Q(MAC_salida_correcta_4_) );
DFFPOSX1 DFFPOSX1_7 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf5), .D(_438__5_), .Q(MAC_salida_correcta_5_) );
DFFPOSX1 DFFPOSX1_8 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf5), .D(_438__6_), .Q(MAC_salida_correcta_6_) );
DFFPOSX1 DFFPOSX1_9 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf5), .D(_438__7_), .Q(MAC_salida_correcta_7_) );
INVX1 INVX1_262 ( .gnd(gnd), .vdd(vdd), .A(asr1_cables_1__0_), .Y(_911_) );
INVX1 INVX1_263 ( .gnd(gnd), .vdd(vdd), .A(asr1_cables_2__0_), .Y(_912_) );
INVX1 INVX1_264 ( .gnd(gnd), .vdd(vdd), .A(up_counter_contador_1_), .Y(_913_) );
INVX1 INVX1_265 ( .gnd(gnd), .vdd(vdd), .A(up_counter_contador_2_), .Y(_914_) );
NAND3X1 NAND3X1_111 ( .gnd(gnd), .vdd(vdd), .A(up_counter_contador_0_), .B(_913_), .C(_914_), .Y(_915_) );
INVX1 INVX1_266 ( .gnd(gnd), .vdd(vdd), .A(up_counter_contador_0_), .Y(_916_) );
NAND3X1 NAND3X1_112 ( .gnd(gnd), .vdd(vdd), .A(_916_), .B(_913_), .C(_914_), .Y(_917_) );
OAI22X1 OAI22X1_5 ( .gnd(gnd), .vdd(vdd), .A(_912_), .B(_915_), .C(_911_), .D(_917_), .Y(_918_) );
INVX1 INVX1_267 ( .gnd(gnd), .vdd(vdd), .A(asr1_cables_7__0_), .Y(_919_) );
INVX1 INVX1_268 ( .gnd(gnd), .vdd(vdd), .A(asr1_cables_3__0_), .Y(_920_) );
NAND3X1 NAND3X1_113 ( .gnd(gnd), .vdd(vdd), .A(up_counter_contador_1_), .B(_916_), .C(_914_), .Y(_921_) );
NAND3X1 NAND3X1_114 ( .gnd(gnd), .vdd(vdd), .A(up_counter_contador_1_), .B(up_counter_contador_2_), .C(_916_), .Y(_922_) );
OAI22X1 OAI22X1_6 ( .gnd(gnd), .vdd(vdd), .A(_919_), .B(_922_), .C(_920_), .D(_921_), .Y(_923_) );
NOR2X1 NOR2X1_12 ( .gnd(gnd), .vdd(vdd), .A(_923_), .B(_918_), .Y(_924_) );
INVX1 INVX1_269 ( .gnd(gnd), .vdd(vdd), .A(asr1_cables_5__0_), .Y(_925_) );
INVX1 INVX1_270 ( .gnd(gnd), .vdd(vdd), .A(asr1_cables_4_), .Y(_926_) );
NAND3X1 NAND3X1_115 ( .gnd(gnd), .vdd(vdd), .A(up_counter_contador_0_), .B(up_counter_contador_1_), .C(_914_), .Y(_804_) );
NAND3X1 NAND3X1_116 ( .gnd(gnd), .vdd(vdd), .A(up_counter_contador_2_), .B(_916_), .C(_913_), .Y(_805_) );
OAI22X1 OAI22X1_7 ( .gnd(gnd), .vdd(vdd), .A(_926_), .B(_804_), .C(_925_), .D(_805_), .Y(_806_) );
INVX1 INVX1_271 ( .gnd(gnd), .vdd(vdd), .A(asr1_cables_8__0_), .Y(_807_) );
INVX1 INVX1_272 ( .gnd(gnd), .vdd(vdd), .A(asr1_cables_6__0_), .Y(_808_) );
NAND3X1 NAND3X1_117 ( .gnd(gnd), .vdd(vdd), .A(up_counter_contador_0_), .B(up_counter_contador_1_), .C(up_counter_contador_2_), .Y(_809_) );
NAND3X1 NAND3X1_118 ( .gnd(gnd), .vdd(vdd), .A(up_counter_contador_0_), .B(up_counter_contador_2_), .C(_913_), .Y(_810_) );
OAI22X1 OAI22X1_8 ( .gnd(gnd), .vdd(vdd), .A(_807_), .B(_809_), .C(_808_), .D(_810_), .Y(_811_) );
NOR2X1 NOR2X1_13 ( .gnd(gnd), .vdd(vdd), .A(_811_), .B(_806_), .Y(_812_) );
NAND2X1 NAND2X1_234 ( .gnd(gnd), .vdd(vdd), .A(_812_), .B(_924_), .Y(asr1_q_0_) );
INVX1 INVX1_273 ( .gnd(gnd), .vdd(vdd), .A(asr1_cables_1__1_), .Y(_813_) );
INVX1 INVX1_274 ( .gnd(gnd), .vdd(vdd), .A(asr1_cables_2__1_), .Y(_814_) );
OAI22X1 OAI22X1_9 ( .gnd(gnd), .vdd(vdd), .A(_814_), .B(_915_), .C(_813_), .D(_917_), .Y(_815_) );
INVX1 INVX1_275 ( .gnd(gnd), .vdd(vdd), .A(asr1_cables_6__1_), .Y(_816_) );
INVX1 INVX1_276 ( .gnd(gnd), .vdd(vdd), .A(asr1_cables_3__1_), .Y(_817_) );
OAI22X1 OAI22X1_10 ( .gnd(gnd), .vdd(vdd), .A(_816_), .B(_810_), .C(_817_), .D(_921_), .Y(_818_) );
NOR2X1 NOR2X1_14 ( .gnd(gnd), .vdd(vdd), .A(_818_), .B(_815_), .Y(_819_) );
INVX1 INVX1_277 ( .gnd(gnd), .vdd(vdd), .A(asr1_cables_7__1_), .Y(_820_) );
INVX1 INVX1_278 ( .gnd(gnd), .vdd(vdd), .A(asr1_cables_8__1_), .Y(_821_) );
OAI22X1 OAI22X1_11 ( .gnd(gnd), .vdd(vdd), .A(_821_), .B(_809_), .C(_820_), .D(_922_), .Y(_822_) );
INVX1 INVX1_279 ( .gnd(gnd), .vdd(vdd), .A(asr1_cables_5__1_), .Y(_823_) );
INVX1 INVX1_280 ( .gnd(gnd), .vdd(vdd), .A(_76_), .Y(_824_) );
OAI22X1 OAI22X1_12 ( .gnd(gnd), .vdd(vdd), .A(_824_), .B(_804_), .C(_823_), .D(_805_), .Y(_825_) );
NOR2X1 NOR2X1_15 ( .gnd(gnd), .vdd(vdd), .A(_822_), .B(_825_), .Y(_826_) );
NAND2X1 NAND2X1_235 ( .gnd(gnd), .vdd(vdd), .A(_826_), .B(_819_), .Y(asr1_q_1_) );
INVX1 INVX1_281 ( .gnd(gnd), .vdd(vdd), .A(asr1_cables_1__2_), .Y(_827_) );
INVX1 INVX1_282 ( .gnd(gnd), .vdd(vdd), .A(asr1_cables_2__2_), .Y(_828_) );
OAI22X1 OAI22X1_13 ( .gnd(gnd), .vdd(vdd), .A(_828_), .B(_915_), .C(_827_), .D(_917_), .Y(_829_) );
INVX1 INVX1_283 ( .gnd(gnd), .vdd(vdd), .A(asr1_cables_7__2_), .Y(_830_) );
INVX1 INVX1_284 ( .gnd(gnd), .vdd(vdd), .A(asr1_cables_3__2_), .Y(_831_) );
OAI22X1 OAI22X1_14 ( .gnd(gnd), .vdd(vdd), .A(_830_), .B(_922_), .C(_831_), .D(_921_), .Y(_832_) );
NOR2X1 NOR2X1_16 ( .gnd(gnd), .vdd(vdd), .A(_832_), .B(_829_), .Y(_833_) );
INVX1 INVX1_285 ( .gnd(gnd), .vdd(vdd), .A(asr1_cables_5__2_), .Y(_834_) );
INVX1 INVX1_286 ( .gnd(gnd), .vdd(vdd), .A(_82_), .Y(_835_) );
OAI22X1 OAI22X1_15 ( .gnd(gnd), .vdd(vdd), .A(_835_), .B(_804_), .C(_834_), .D(_805_), .Y(_836_) );
INVX1 INVX1_287 ( .gnd(gnd), .vdd(vdd), .A(asr1_cables_8__2_), .Y(_837_) );
INVX1 INVX1_288 ( .gnd(gnd), .vdd(vdd), .A(asr1_cables_6__2_), .Y(_838_) );
OAI22X1 OAI22X1_16 ( .gnd(gnd), .vdd(vdd), .A(_837_), .B(_809_), .C(_838_), .D(_810_), .Y(_839_) );
NOR2X1 NOR2X1_17 ( .gnd(gnd), .vdd(vdd), .A(_839_), .B(_836_), .Y(_840_) );
NAND2X1 NAND2X1_236 ( .gnd(gnd), .vdd(vdd), .A(_840_), .B(_833_), .Y(asr1_q_2_) );
INVX1 INVX1_289 ( .gnd(gnd), .vdd(vdd), .A(asr1_cables_3__3_), .Y(_841_) );
INVX1 INVX1_290 ( .gnd(gnd), .vdd(vdd), .A(asr1_cables_2__3_), .Y(_842_) );
OAI22X1 OAI22X1_17 ( .gnd(gnd), .vdd(vdd), .A(_841_), .B(_921_), .C(_842_), .D(_915_), .Y(_843_) );
INVX1 INVX1_291 ( .gnd(gnd), .vdd(vdd), .A(asr1_cables_7__3_), .Y(_844_) );
INVX1 INVX1_292 ( .gnd(gnd), .vdd(vdd), .A(asr1_cables_6__3_), .Y(_845_) );
OAI22X1 OAI22X1_18 ( .gnd(gnd), .vdd(vdd), .A(_844_), .B(_922_), .C(_845_), .D(_810_), .Y(_846_) );
NOR2X1 NOR2X1_18 ( .gnd(gnd), .vdd(vdd), .A(_846_), .B(_843_), .Y(_847_) );
INVX1 INVX1_293 ( .gnd(gnd), .vdd(vdd), .A(asr1_cables_5__3_), .Y(_848_) );
INVX1 INVX1_294 ( .gnd(gnd), .vdd(vdd), .A(_77_), .Y(_849_) );
OAI22X1 OAI22X1_19 ( .gnd(gnd), .vdd(vdd), .A(_849_), .B(_804_), .C(_848_), .D(_805_), .Y(_850_) );
INVX1 INVX1_295 ( .gnd(gnd), .vdd(vdd), .A(asr1_cables_8__3_), .Y(_851_) );
INVX1 INVX1_296 ( .gnd(gnd), .vdd(vdd), .A(asr1_cables_1__3_), .Y(_852_) );
OAI22X1 OAI22X1_20 ( .gnd(gnd), .vdd(vdd), .A(_851_), .B(_809_), .C(_852_), .D(_917_), .Y(_853_) );
NOR2X1 NOR2X1_19 ( .gnd(gnd), .vdd(vdd), .A(_850_), .B(_853_), .Y(_854_) );
NAND2X1 NAND2X1_237 ( .gnd(gnd), .vdd(vdd), .A(_847_), .B(_854_), .Y(asr1_q_3_) );
INVX1 INVX1_297 ( .gnd(gnd), .vdd(vdd), .A(asr1_cables_1__4_), .Y(_855_) );
INVX1 INVX1_298 ( .gnd(gnd), .vdd(vdd), .A(asr1_cables_2__4_), .Y(_856_) );
OAI22X1 OAI22X1_21 ( .gnd(gnd), .vdd(vdd), .A(_856_), .B(_915_), .C(_855_), .D(_917_), .Y(_857_) );
INVX1 INVX1_299 ( .gnd(gnd), .vdd(vdd), .A(asr1_cables_7__4_), .Y(_858_) );
INVX1 INVX1_300 ( .gnd(gnd), .vdd(vdd), .A(asr1_cables_3__4_), .Y(_859_) );
OAI22X1 OAI22X1_22 ( .gnd(gnd), .vdd(vdd), .A(_858_), .B(_922_), .C(_859_), .D(_921_), .Y(_860_) );
NOR2X1 NOR2X1_20 ( .gnd(gnd), .vdd(vdd), .A(_860_), .B(_857_), .Y(_861_) );
INVX1 INVX1_301 ( .gnd(gnd), .vdd(vdd), .A(asr1_cables_5__4_), .Y(_862_) );
INVX1 INVX1_302 ( .gnd(gnd), .vdd(vdd), .A(_78_), .Y(_863_) );
OAI22X1 OAI22X1_23 ( .gnd(gnd), .vdd(vdd), .A(_863_), .B(_804_), .C(_862_), .D(_805_), .Y(_864_) );
INVX1 INVX1_303 ( .gnd(gnd), .vdd(vdd), .A(asr1_cables_8__4_), .Y(_865_) );
INVX1 INVX1_304 ( .gnd(gnd), .vdd(vdd), .A(asr1_cables_6__4_), .Y(_866_) );
OAI22X1 OAI22X1_24 ( .gnd(gnd), .vdd(vdd), .A(_865_), .B(_809_), .C(_866_), .D(_810_), .Y(_867_) );
NOR2X1 NOR2X1_21 ( .gnd(gnd), .vdd(vdd), .A(_867_), .B(_864_), .Y(_868_) );
NAND2X1 NAND2X1_238 ( .gnd(gnd), .vdd(vdd), .A(_868_), .B(_861_), .Y(asr1_q_4_) );
INVX1 INVX1_305 ( .gnd(gnd), .vdd(vdd), .A(asr1_cables_3__5_), .Y(_869_) );
INVX1 INVX1_306 ( .gnd(gnd), .vdd(vdd), .A(asr1_cables_2__5_), .Y(_870_) );
OAI22X1 OAI22X1_25 ( .gnd(gnd), .vdd(vdd), .A(_869_), .B(_921_), .C(_870_), .D(_915_), .Y(_871_) );
INVX1 INVX1_307 ( .gnd(gnd), .vdd(vdd), .A(asr1_cables_7__5_), .Y(_872_) );
INVX1 INVX1_308 ( .gnd(gnd), .vdd(vdd), .A(asr1_cables_6__5_), .Y(_873_) );
OAI22X1 OAI22X1_26 ( .gnd(gnd), .vdd(vdd), .A(_872_), .B(_922_), .C(_873_), .D(_810_), .Y(_874_) );
NOR2X1 NOR2X1_22 ( .gnd(gnd), .vdd(vdd), .A(_874_), .B(_871_), .Y(_875_) );
INVX1 INVX1_309 ( .gnd(gnd), .vdd(vdd), .A(asr1_cables_5__5_), .Y(_876_) );
INVX1 INVX1_310 ( .gnd(gnd), .vdd(vdd), .A(_79_), .Y(_877_) );
OAI22X1 OAI22X1_27 ( .gnd(gnd), .vdd(vdd), .A(_877_), .B(_804_), .C(_876_), .D(_805_), .Y(_878_) );
INVX1 INVX1_311 ( .gnd(gnd), .vdd(vdd), .A(asr1_cables_8__5_), .Y(_879_) );
INVX1 INVX1_312 ( .gnd(gnd), .vdd(vdd), .A(asr1_cables_1__5_), .Y(_880_) );
OAI22X1 OAI22X1_28 ( .gnd(gnd), .vdd(vdd), .A(_879_), .B(_809_), .C(_880_), .D(_917_), .Y(_881_) );
NOR2X1 NOR2X1_23 ( .gnd(gnd), .vdd(vdd), .A(_878_), .B(_881_), .Y(_882_) );
NAND2X1 NAND2X1_239 ( .gnd(gnd), .vdd(vdd), .A(_875_), .B(_882_), .Y(asr1_q_5_) );
INVX1 INVX1_313 ( .gnd(gnd), .vdd(vdd), .A(asr1_cables_1__6_), .Y(_883_) );
INVX1 INVX1_314 ( .gnd(gnd), .vdd(vdd), .A(asr1_cables_2__6_), .Y(_884_) );
OAI22X1 OAI22X1_29 ( .gnd(gnd), .vdd(vdd), .A(_884_), .B(_915_), .C(_883_), .D(_917_), .Y(_885_) );
INVX1 INVX1_315 ( .gnd(gnd), .vdd(vdd), .A(asr1_cables_7__6_), .Y(_886_) );
INVX1 INVX1_316 ( .gnd(gnd), .vdd(vdd), .A(asr1_cables_3__6_), .Y(_887_) );
OAI22X1 OAI22X1_30 ( .gnd(gnd), .vdd(vdd), .A(_886_), .B(_922_), .C(_887_), .D(_921_), .Y(_888_) );
NOR2X1 NOR2X1_24 ( .gnd(gnd), .vdd(vdd), .A(_888_), .B(_885_), .Y(_889_) );
INVX1 INVX1_317 ( .gnd(gnd), .vdd(vdd), .A(asr1_cables_5__6_), .Y(_890_) );
INVX1 INVX1_318 ( .gnd(gnd), .vdd(vdd), .A(_80_), .Y(_891_) );
OAI22X1 OAI22X1_31 ( .gnd(gnd), .vdd(vdd), .A(_891_), .B(_804_), .C(_890_), .D(_805_), .Y(_892_) );
INVX1 INVX1_319 ( .gnd(gnd), .vdd(vdd), .A(asr1_cables_8__6_), .Y(_893_) );
INVX1 INVX1_320 ( .gnd(gnd), .vdd(vdd), .A(asr1_cables_6__6_), .Y(_894_) );
OAI22X1 OAI22X1_32 ( .gnd(gnd), .vdd(vdd), .A(_893_), .B(_809_), .C(_894_), .D(_810_), .Y(_895_) );
NOR2X1 NOR2X1_25 ( .gnd(gnd), .vdd(vdd), .A(_895_), .B(_892_), .Y(_896_) );
NAND2X1 NAND2X1_240 ( .gnd(gnd), .vdd(vdd), .A(_896_), .B(_889_), .Y(asr1_q_6_) );
INVX1 INVX1_321 ( .gnd(gnd), .vdd(vdd), .A(asr1_cables_3__7_), .Y(_897_) );
INVX1 INVX1_322 ( .gnd(gnd), .vdd(vdd), .A(asr1_cables_2__7_), .Y(_898_) );
OAI22X1 OAI22X1_33 ( .gnd(gnd), .vdd(vdd), .A(_897_), .B(_921_), .C(_898_), .D(_915_), .Y(_899_) );
INVX1 INVX1_323 ( .gnd(gnd), .vdd(vdd), .A(asr1_cables_7__7_), .Y(_900_) );
INVX1 INVX1_324 ( .gnd(gnd), .vdd(vdd), .A(asr1_cables_6__7_), .Y(_901_) );
OAI22X1 OAI22X1_34 ( .gnd(gnd), .vdd(vdd), .A(_900_), .B(_922_), .C(_901_), .D(_810_), .Y(_902_) );
NOR2X1 NOR2X1_26 ( .gnd(gnd), .vdd(vdd), .A(_902_), .B(_899_), .Y(_903_) );
INVX1 INVX1_325 ( .gnd(gnd), .vdd(vdd), .A(asr1_cables_5__7_), .Y(_904_) );
INVX1 INVX1_326 ( .gnd(gnd), .vdd(vdd), .A(_81_), .Y(_905_) );
OAI22X1 OAI22X1_35 ( .gnd(gnd), .vdd(vdd), .A(_905_), .B(_804_), .C(_904_), .D(_805_), .Y(_906_) );
INVX1 INVX1_327 ( .gnd(gnd), .vdd(vdd), .A(asr1_cables_8__7_), .Y(_907_) );
INVX1 INVX1_328 ( .gnd(gnd), .vdd(vdd), .A(asr1_cables_1__7_), .Y(_908_) );
OAI22X1 OAI22X1_36 ( .gnd(gnd), .vdd(vdd), .A(_907_), .B(_809_), .C(_908_), .D(_917_), .Y(_909_) );
NOR2X1 NOR2X1_27 ( .gnd(gnd), .vdd(vdd), .A(_906_), .B(_909_), .Y(_910_) );
NAND2X1 NAND2X1_241 ( .gnd(gnd), .vdd(vdd), .A(_903_), .B(_910_), .Y(asr1_q_7_) );
INVX1 INVX1_329 ( .gnd(gnd), .vdd(vdd), .A(asr2_cables_1__0_), .Y(_1034_) );
INVX1 INVX1_330 ( .gnd(gnd), .vdd(vdd), .A(asr2_cables_2__0_), .Y(_1035_) );
INVX1 INVX1_331 ( .gnd(gnd), .vdd(vdd), .A(down_counter_contador_1_), .Y(_1036_) );
INVX1 INVX1_332 ( .gnd(gnd), .vdd(vdd), .A(down_counter_contador_2_), .Y(_1037_) );
NAND3X1 NAND3X1_119 ( .gnd(gnd), .vdd(vdd), .A(down_counter_contador_0_), .B(_1036_), .C(_1037_), .Y(_1038_) );
INVX1 INVX1_333 ( .gnd(gnd), .vdd(vdd), .A(down_counter_contador_0_), .Y(_1039_) );
NAND3X1 NAND3X1_120 ( .gnd(gnd), .vdd(vdd), .A(_1039_), .B(_1036_), .C(_1037_), .Y(_1040_) );
OAI22X1 OAI22X1_37 ( .gnd(gnd), .vdd(vdd), .A(_1035_), .B(_1038_), .C(_1034_), .D(_1040_), .Y(_1041_) );
INVX1 INVX1_334 ( .gnd(gnd), .vdd(vdd), .A(asr2_cables_7__0_), .Y(_1042_) );
INVX1 INVX1_335 ( .gnd(gnd), .vdd(vdd), .A(asr2_cables_3__0_), .Y(_1043_) );
NAND3X1 NAND3X1_121 ( .gnd(gnd), .vdd(vdd), .A(down_counter_contador_1_), .B(_1039_), .C(_1037_), .Y(_1044_) );
NAND3X1 NAND3X1_122 ( .gnd(gnd), .vdd(vdd), .A(down_counter_contador_1_), .B(down_counter_contador_2_), .C(_1039_), .Y(_1045_) );
OAI22X1 OAI22X1_38 ( .gnd(gnd), .vdd(vdd), .A(_1042_), .B(_1045_), .C(_1043_), .D(_1044_), .Y(_1046_) );
NOR2X1 NOR2X1_28 ( .gnd(gnd), .vdd(vdd), .A(_1046_), .B(_1041_), .Y(_1047_) );
INVX1 INVX1_336 ( .gnd(gnd), .vdd(vdd), .A(asr2_cables_5__0_), .Y(_1048_) );
INVX1 INVX1_337 ( .gnd(gnd), .vdd(vdd), .A(asr2_cables_4_), .Y(_1049_) );
NAND3X1 NAND3X1_123 ( .gnd(gnd), .vdd(vdd), .A(down_counter_contador_0_), .B(down_counter_contador_1_), .C(_1037_), .Y(_927_) );
NAND3X1 NAND3X1_124 ( .gnd(gnd), .vdd(vdd), .A(down_counter_contador_2_), .B(_1039_), .C(_1036_), .Y(_928_) );
OAI22X1 OAI22X1_39 ( .gnd(gnd), .vdd(vdd), .A(_1049_), .B(_927_), .C(_1048_), .D(_928_), .Y(_929_) );
INVX1 INVX1_338 ( .gnd(gnd), .vdd(vdd), .A(asr2_cables_8__0_), .Y(_930_) );
INVX1 INVX1_339 ( .gnd(gnd), .vdd(vdd), .A(asr2_cables_6__0_), .Y(_931_) );
NAND3X1 NAND3X1_125 ( .gnd(gnd), .vdd(vdd), .A(down_counter_contador_0_), .B(down_counter_contador_1_), .C(down_counter_contador_2_), .Y(_932_) );
NAND3X1 NAND3X1_126 ( .gnd(gnd), .vdd(vdd), .A(down_counter_contador_0_), .B(down_counter_contador_2_), .C(_1036_), .Y(_933_) );
OAI22X1 OAI22X1_40 ( .gnd(gnd), .vdd(vdd), .A(_930_), .B(_932_), .C(_931_), .D(_933_), .Y(_934_) );
NOR2X1 NOR2X1_29 ( .gnd(gnd), .vdd(vdd), .A(_934_), .B(_929_), .Y(_935_) );
NAND2X1 NAND2X1_242 ( .gnd(gnd), .vdd(vdd), .A(_935_), .B(_1047_), .Y(asr2_q_0_) );
INVX1 INVX1_340 ( .gnd(gnd), .vdd(vdd), .A(asr2_cables_1__1_), .Y(_936_) );
INVX1 INVX1_341 ( .gnd(gnd), .vdd(vdd), .A(asr2_cables_2__1_), .Y(_937_) );
OAI22X1 OAI22X1_41 ( .gnd(gnd), .vdd(vdd), .A(_937_), .B(_1038_), .C(_936_), .D(_1040_), .Y(_938_) );
INVX1 INVX1_342 ( .gnd(gnd), .vdd(vdd), .A(asr2_cables_6__1_), .Y(_939_) );
INVX1 INVX1_343 ( .gnd(gnd), .vdd(vdd), .A(asr2_cables_3__1_), .Y(_940_) );
OAI22X1 OAI22X1_42 ( .gnd(gnd), .vdd(vdd), .A(_939_), .B(_933_), .C(_940_), .D(_1044_), .Y(_941_) );
NOR2X1 NOR2X1_30 ( .gnd(gnd), .vdd(vdd), .A(_941_), .B(_938_), .Y(_942_) );
INVX1 INVX1_344 ( .gnd(gnd), .vdd(vdd), .A(asr2_cables_7__1_), .Y(_943_) );
INVX1 INVX1_345 ( .gnd(gnd), .vdd(vdd), .A(asr2_cables_8__1_), .Y(_944_) );
OAI22X1 OAI22X1_43 ( .gnd(gnd), .vdd(vdd), .A(_944_), .B(_932_), .C(_943_), .D(_1045_), .Y(_945_) );
INVX1 INVX1_346 ( .gnd(gnd), .vdd(vdd), .A(asr2_cables_5__1_), .Y(_946_) );
INVX1 INVX1_347 ( .gnd(gnd), .vdd(vdd), .A(_227_), .Y(_947_) );
OAI22X1 OAI22X1_44 ( .gnd(gnd), .vdd(vdd), .A(_947_), .B(_927_), .C(_946_), .D(_928_), .Y(_948_) );
NOR2X1 NOR2X1_31 ( .gnd(gnd), .vdd(vdd), .A(_945_), .B(_948_), .Y(_949_) );
NAND2X1 NAND2X1_243 ( .gnd(gnd), .vdd(vdd), .A(_949_), .B(_942_), .Y(asr2_q_1_) );
INVX1 INVX1_348 ( .gnd(gnd), .vdd(vdd), .A(asr2_cables_1__2_), .Y(_950_) );
INVX1 INVX1_349 ( .gnd(gnd), .vdd(vdd), .A(asr2_cables_2__2_), .Y(_951_) );
OAI22X1 OAI22X1_45 ( .gnd(gnd), .vdd(vdd), .A(_951_), .B(_1038_), .C(_950_), .D(_1040_), .Y(_952_) );
INVX1 INVX1_350 ( .gnd(gnd), .vdd(vdd), .A(asr2_cables_7__2_), .Y(_953_) );
INVX1 INVX1_351 ( .gnd(gnd), .vdd(vdd), .A(asr2_cables_3__2_), .Y(_954_) );
OAI22X1 OAI22X1_46 ( .gnd(gnd), .vdd(vdd), .A(_953_), .B(_1045_), .C(_954_), .D(_1044_), .Y(_955_) );
NOR2X1 NOR2X1_32 ( .gnd(gnd), .vdd(vdd), .A(_955_), .B(_952_), .Y(_956_) );
INVX1 INVX1_352 ( .gnd(gnd), .vdd(vdd), .A(asr2_cables_5__2_), .Y(_957_) );
INVX1 INVX1_353 ( .gnd(gnd), .vdd(vdd), .A(_233_), .Y(_958_) );
OAI22X1 OAI22X1_47 ( .gnd(gnd), .vdd(vdd), .A(_958_), .B(_927_), .C(_957_), .D(_928_), .Y(_959_) );
INVX1 INVX1_354 ( .gnd(gnd), .vdd(vdd), .A(asr2_cables_8__2_), .Y(_960_) );
INVX1 INVX1_355 ( .gnd(gnd), .vdd(vdd), .A(asr2_cables_6__2_), .Y(_961_) );
OAI22X1 OAI22X1_48 ( .gnd(gnd), .vdd(vdd), .A(_960_), .B(_932_), .C(_961_), .D(_933_), .Y(_962_) );
NOR2X1 NOR2X1_33 ( .gnd(gnd), .vdd(vdd), .A(_962_), .B(_959_), .Y(_963_) );
NAND2X1 NAND2X1_244 ( .gnd(gnd), .vdd(vdd), .A(_963_), .B(_956_), .Y(asr2_q_2_) );
INVX1 INVX1_356 ( .gnd(gnd), .vdd(vdd), .A(asr2_cables_3__3_), .Y(_964_) );
INVX1 INVX1_357 ( .gnd(gnd), .vdd(vdd), .A(asr2_cables_2__3_), .Y(_965_) );
OAI22X1 OAI22X1_49 ( .gnd(gnd), .vdd(vdd), .A(_964_), .B(_1044_), .C(_965_), .D(_1038_), .Y(_966_) );
INVX1 INVX1_358 ( .gnd(gnd), .vdd(vdd), .A(asr2_cables_7__3_), .Y(_967_) );
INVX1 INVX1_359 ( .gnd(gnd), .vdd(vdd), .A(asr2_cables_6__3_), .Y(_968_) );
OAI22X1 OAI22X1_50 ( .gnd(gnd), .vdd(vdd), .A(_967_), .B(_1045_), .C(_968_), .D(_933_), .Y(_969_) );
NOR2X1 NOR2X1_34 ( .gnd(gnd), .vdd(vdd), .A(_969_), .B(_966_), .Y(_970_) );
INVX1 INVX1_360 ( .gnd(gnd), .vdd(vdd), .A(asr2_cables_5__3_), .Y(_971_) );
INVX1 INVX1_361 ( .gnd(gnd), .vdd(vdd), .A(_228_), .Y(_972_) );
OAI22X1 OAI22X1_51 ( .gnd(gnd), .vdd(vdd), .A(_972_), .B(_927_), .C(_971_), .D(_928_), .Y(_973_) );
INVX1 INVX1_362 ( .gnd(gnd), .vdd(vdd), .A(asr2_cables_8__3_), .Y(_974_) );
INVX1 INVX1_363 ( .gnd(gnd), .vdd(vdd), .A(asr2_cables_1__3_), .Y(_975_) );
OAI22X1 OAI22X1_52 ( .gnd(gnd), .vdd(vdd), .A(_974_), .B(_932_), .C(_975_), .D(_1040_), .Y(_976_) );
NOR2X1 NOR2X1_35 ( .gnd(gnd), .vdd(vdd), .A(_973_), .B(_976_), .Y(_977_) );
NAND2X1 NAND2X1_245 ( .gnd(gnd), .vdd(vdd), .A(_970_), .B(_977_), .Y(asr2_q_3_) );
INVX1 INVX1_364 ( .gnd(gnd), .vdd(vdd), .A(asr2_cables_1__4_), .Y(_978_) );
INVX1 INVX1_365 ( .gnd(gnd), .vdd(vdd), .A(asr2_cables_2__4_), .Y(_979_) );
OAI22X1 OAI22X1_53 ( .gnd(gnd), .vdd(vdd), .A(_979_), .B(_1038_), .C(_978_), .D(_1040_), .Y(_980_) );
INVX1 INVX1_366 ( .gnd(gnd), .vdd(vdd), .A(asr2_cables_7__4_), .Y(_981_) );
INVX1 INVX1_367 ( .gnd(gnd), .vdd(vdd), .A(asr2_cables_3__4_), .Y(_982_) );
OAI22X1 OAI22X1_54 ( .gnd(gnd), .vdd(vdd), .A(_981_), .B(_1045_), .C(_982_), .D(_1044_), .Y(_983_) );
NOR2X1 NOR2X1_36 ( .gnd(gnd), .vdd(vdd), .A(_983_), .B(_980_), .Y(_984_) );
INVX1 INVX1_368 ( .gnd(gnd), .vdd(vdd), .A(asr2_cables_5__4_), .Y(_985_) );
INVX1 INVX1_369 ( .gnd(gnd), .vdd(vdd), .A(_229_), .Y(_986_) );
OAI22X1 OAI22X1_55 ( .gnd(gnd), .vdd(vdd), .A(_986_), .B(_927_), .C(_985_), .D(_928_), .Y(_987_) );
INVX1 INVX1_370 ( .gnd(gnd), .vdd(vdd), .A(asr2_cables_8__4_), .Y(_988_) );
INVX1 INVX1_371 ( .gnd(gnd), .vdd(vdd), .A(asr2_cables_6__4_), .Y(_989_) );
OAI22X1 OAI22X1_56 ( .gnd(gnd), .vdd(vdd), .A(_988_), .B(_932_), .C(_989_), .D(_933_), .Y(_990_) );
NOR2X1 NOR2X1_37 ( .gnd(gnd), .vdd(vdd), .A(_990_), .B(_987_), .Y(_991_) );
NAND2X1 NAND2X1_246 ( .gnd(gnd), .vdd(vdd), .A(_991_), .B(_984_), .Y(asr2_q_4_) );
INVX1 INVX1_372 ( .gnd(gnd), .vdd(vdd), .A(asr2_cables_3__5_), .Y(_992_) );
INVX1 INVX1_373 ( .gnd(gnd), .vdd(vdd), .A(asr2_cables_2__5_), .Y(_993_) );
OAI22X1 OAI22X1_57 ( .gnd(gnd), .vdd(vdd), .A(_992_), .B(_1044_), .C(_993_), .D(_1038_), .Y(_994_) );
INVX1 INVX1_374 ( .gnd(gnd), .vdd(vdd), .A(asr2_cables_7__5_), .Y(_995_) );
INVX1 INVX1_375 ( .gnd(gnd), .vdd(vdd), .A(asr2_cables_6__5_), .Y(_996_) );
OAI22X1 OAI22X1_58 ( .gnd(gnd), .vdd(vdd), .A(_995_), .B(_1045_), .C(_996_), .D(_933_), .Y(_997_) );
NOR2X1 NOR2X1_38 ( .gnd(gnd), .vdd(vdd), .A(_997_), .B(_994_), .Y(_998_) );
INVX1 INVX1_376 ( .gnd(gnd), .vdd(vdd), .A(asr2_cables_5__5_), .Y(_999_) );
INVX1 INVX1_377 ( .gnd(gnd), .vdd(vdd), .A(_230_), .Y(_1000_) );
OAI22X1 OAI22X1_59 ( .gnd(gnd), .vdd(vdd), .A(_1000_), .B(_927_), .C(_999_), .D(_928_), .Y(_1001_) );
INVX1 INVX1_378 ( .gnd(gnd), .vdd(vdd), .A(asr2_cables_8__5_), .Y(_1002_) );
INVX1 INVX1_379 ( .gnd(gnd), .vdd(vdd), .A(asr2_cables_1__5_), .Y(_1003_) );
OAI22X1 OAI22X1_60 ( .gnd(gnd), .vdd(vdd), .A(_1002_), .B(_932_), .C(_1003_), .D(_1040_), .Y(_1004_) );
NOR2X1 NOR2X1_39 ( .gnd(gnd), .vdd(vdd), .A(_1001_), .B(_1004_), .Y(_1005_) );
NAND2X1 NAND2X1_247 ( .gnd(gnd), .vdd(vdd), .A(_998_), .B(_1005_), .Y(asr2_q_5_) );
INVX1 INVX1_380 ( .gnd(gnd), .vdd(vdd), .A(asr2_cables_1__6_), .Y(_1006_) );
INVX1 INVX1_381 ( .gnd(gnd), .vdd(vdd), .A(asr2_cables_2__6_), .Y(_1007_) );
OAI22X1 OAI22X1_61 ( .gnd(gnd), .vdd(vdd), .A(_1007_), .B(_1038_), .C(_1006_), .D(_1040_), .Y(_1008_) );
INVX1 INVX1_382 ( .gnd(gnd), .vdd(vdd), .A(asr2_cables_7__6_), .Y(_1009_) );
INVX1 INVX1_383 ( .gnd(gnd), .vdd(vdd), .A(asr2_cables_3__6_), .Y(_1010_) );
OAI22X1 OAI22X1_62 ( .gnd(gnd), .vdd(vdd), .A(_1009_), .B(_1045_), .C(_1010_), .D(_1044_), .Y(_1011_) );
NOR2X1 NOR2X1_40 ( .gnd(gnd), .vdd(vdd), .A(_1011_), .B(_1008_), .Y(_1012_) );
INVX1 INVX1_384 ( .gnd(gnd), .vdd(vdd), .A(asr2_cables_5__6_), .Y(_1013_) );
INVX1 INVX1_385 ( .gnd(gnd), .vdd(vdd), .A(_231_), .Y(_1014_) );
OAI22X1 OAI22X1_63 ( .gnd(gnd), .vdd(vdd), .A(_1014_), .B(_927_), .C(_1013_), .D(_928_), .Y(_1015_) );
INVX1 INVX1_386 ( .gnd(gnd), .vdd(vdd), .A(asr2_cables_8__6_), .Y(_1016_) );
INVX1 INVX1_387 ( .gnd(gnd), .vdd(vdd), .A(asr2_cables_6__6_), .Y(_1017_) );
OAI22X1 OAI22X1_64 ( .gnd(gnd), .vdd(vdd), .A(_1016_), .B(_932_), .C(_1017_), .D(_933_), .Y(_1018_) );
NOR2X1 NOR2X1_41 ( .gnd(gnd), .vdd(vdd), .A(_1018_), .B(_1015_), .Y(_1019_) );
NAND2X1 NAND2X1_248 ( .gnd(gnd), .vdd(vdd), .A(_1019_), .B(_1012_), .Y(asr2_q_6_) );
INVX1 INVX1_388 ( .gnd(gnd), .vdd(vdd), .A(asr2_cables_3__7_), .Y(_1020_) );
INVX1 INVX1_389 ( .gnd(gnd), .vdd(vdd), .A(asr2_cables_2__7_), .Y(_1021_) );
OAI22X1 OAI22X1_65 ( .gnd(gnd), .vdd(vdd), .A(_1020_), .B(_1044_), .C(_1021_), .D(_1038_), .Y(_1022_) );
INVX1 INVX1_390 ( .gnd(gnd), .vdd(vdd), .A(asr2_cables_7__7_), .Y(_1023_) );
INVX1 INVX1_391 ( .gnd(gnd), .vdd(vdd), .A(asr2_cables_6__7_), .Y(_1024_) );
OAI22X1 OAI22X1_66 ( .gnd(gnd), .vdd(vdd), .A(_1023_), .B(_1045_), .C(_1024_), .D(_933_), .Y(_1025_) );
NOR2X1 NOR2X1_42 ( .gnd(gnd), .vdd(vdd), .A(_1025_), .B(_1022_), .Y(_1026_) );
INVX1 INVX1_392 ( .gnd(gnd), .vdd(vdd), .A(asr2_cables_5__7_), .Y(_1027_) );
INVX1 INVX1_393 ( .gnd(gnd), .vdd(vdd), .A(_232_), .Y(_1028_) );
OAI22X1 OAI22X1_67 ( .gnd(gnd), .vdd(vdd), .A(_1028_), .B(_927_), .C(_1027_), .D(_928_), .Y(_1029_) );
INVX1 INVX1_394 ( .gnd(gnd), .vdd(vdd), .A(asr2_cables_8__7_), .Y(_1030_) );
INVX1 INVX1_395 ( .gnd(gnd), .vdd(vdd), .A(asr2_cables_1__7_), .Y(_1031_) );
OAI22X1 OAI22X1_68 ( .gnd(gnd), .vdd(vdd), .A(_1030_), .B(_932_), .C(_1031_), .D(_1040_), .Y(_1032_) );
NOR2X1 NOR2X1_43 ( .gnd(gnd), .vdd(vdd), .A(_1029_), .B(_1032_), .Y(_1033_) );
NAND2X1 NAND2X1_249 ( .gnd(gnd), .vdd(vdd), .A(_1026_), .B(_1033_), .Y(asr2_q_7_) );
INVX1 INVX1_396 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf3), .Y(_1057_) );
NAND2X1 NAND2X1_250 ( .gnd(gnd), .vdd(vdd), .A(down_counter_contador_0_), .B(_1057_), .Y(_1050__0_) );
AOI21X1 AOI21X1_40 ( .gnd(gnd), .vdd(vdd), .A(down_counter_contador_0_), .B(down_counter_contador_1_), .C(rst_bF_buf3), .Y(_1051_) );
OAI21X1 OAI21X1_239 ( .gnd(gnd), .vdd(vdd), .A(down_counter_contador_0_), .B(down_counter_contador_1_), .C(_1051_), .Y(_1050__1_) );
OAI21X1 OAI21X1_240 ( .gnd(gnd), .vdd(vdd), .A(down_counter_contador_0_), .B(down_counter_contador_1_), .C(down_counter_contador_2_), .Y(_1052_) );
INVX1 INVX1_397 ( .gnd(gnd), .vdd(vdd), .A(down_counter_contador_0_), .Y(_1053_) );
INVX1 INVX1_398 ( .gnd(gnd), .vdd(vdd), .A(down_counter_contador_1_), .Y(_1054_) );
INVX1 INVX1_399 ( .gnd(gnd), .vdd(vdd), .A(down_counter_contador_2_), .Y(_1055_) );
NAND3X1 NAND3X1_127 ( .gnd(gnd), .vdd(vdd), .A(_1053_), .B(_1054_), .C(_1055_), .Y(_1056_) );
NAND3X1 NAND3X1_128 ( .gnd(gnd), .vdd(vdd), .A(_1057_), .B(_1052_), .C(_1056_), .Y(_1050__2_) );
DFFPOSX1 DFFPOSX1_10 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf1), .D(_1050__0_), .Q(down_counter_contador_0_) );
DFFPOSX1 DFFPOSX1_11 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf4), .D(_1050__1_), .Q(down_counter_contador_1_) );
DFFPOSX1 DFFPOSX1_12 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf4), .D(_1050__2_), .Q(down_counter_contador_2_) );
NOR2X1 NOR2X1_44 ( .gnd(gnd), .vdd(vdd), .A(generador_clock_counter_0_), .B(rst_bF_buf1), .Y(_1058__0_) );
AND2X2 AND2X2_14 ( .gnd(gnd), .vdd(vdd), .A(generador_clock_counter_0_), .B(generador_clock_counter_1_), .Y(_1059_) );
INVX1 INVX1_400 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf0), .Y(_1060_) );
OAI21X1 OAI21X1_241 ( .gnd(gnd), .vdd(vdd), .A(generador_clock_counter_0_), .B(generador_clock_counter_1_), .C(_1060_), .Y(_1061_) );
NOR2X1 NOR2X1_45 ( .gnd(gnd), .vdd(vdd), .A(_1059_), .B(_1061_), .Y(_1058__1_) );
INVX1 INVX1_401 ( .gnd(gnd), .vdd(vdd), .A(generador_clock_counter_2_), .Y(_1062_) );
NAND2X1 NAND2X1_251 ( .gnd(gnd), .vdd(vdd), .A(generador_clock_counter_0_), .B(generador_clock_counter_1_), .Y(_1063_) );
OAI21X1 OAI21X1_242 ( .gnd(gnd), .vdd(vdd), .A(_1062_), .B(_1063_), .C(_1060_), .Y(_1064_) );
AOI21X1 AOI21X1_41 ( .gnd(gnd), .vdd(vdd), .A(_1062_), .B(_1063_), .C(_1064_), .Y(_1058__2_) );
OAI21X1 OAI21X1_243 ( .gnd(gnd), .vdd(vdd), .A(_1062_), .B(_1063_), .C(generador_clock_counter_3_), .Y(_1065_) );
INVX1 INVX1_402 ( .gnd(gnd), .vdd(vdd), .A(generador_clock_counter_3_), .Y(asr1_clk) );
NAND3X1 NAND3X1_129 ( .gnd(gnd), .vdd(vdd), .A(asr1_clk_bF_buf7), .B(generador_clock_counter_2_), .C(_1059_), .Y(_1066_) );
AOI21X1 AOI21X1_42 ( .gnd(gnd), .vdd(vdd), .A(_1066_), .B(_1065_), .C(rst_bF_buf0), .Y(_1058__3_) );
DFFPOSX1 DFFPOSX1_13 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf2), .D(_1058__0_), .Q(generador_clock_counter_0_) );
DFFPOSX1 DFFPOSX1_14 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf7), .D(_1058__1_), .Q(generador_clock_counter_1_) );
DFFPOSX1 DFFPOSX1_15 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf7), .D(_1058__2_), .Q(generador_clock_counter_2_) );
DFFPOSX1 DFFPOSX1_16 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf7), .D(_1058__3_), .Q(generador_clock_counter_3_) );
INVX1 INVX1_403 ( .gnd(gnd), .vdd(vdd), .A(up_counter_contador_0_), .Y(_1067_) );
INVX1 INVX1_404 ( .gnd(gnd), .vdd(vdd), .A(up_counter_contador_2_), .Y(_1075_) );
NAND3X1 NAND3X1_130 ( .gnd(gnd), .vdd(vdd), .A(up_counter_contador_0_), .B(up_counter_contador_1_), .C(_1075_), .Y(_1071_) );
NAND2X1 NAND2X1_252 ( .gnd(gnd), .vdd(vdd), .A(up_counter_contador_0_), .B(up_counter_contador_1_), .Y(_1072_) );
NAND2X1 NAND2X1_253 ( .gnd(gnd), .vdd(vdd), .A(up_counter_contador_2_), .B(_1072_), .Y(_1073_) );
NAND2X1 NAND2X1_254 ( .gnd(gnd), .vdd(vdd), .A(_1073_), .B(_1071_), .Y(_1069_) );
NAND3X1 NAND3X1_131 ( .gnd(gnd), .vdd(vdd), .A(up_counter_contador_0_), .B(up_counter_contador_1_), .C(up_counter_contador_2_), .Y(_1074_) );
INVX1 INVX1_405 ( .gnd(gnd), .vdd(vdd), .A(_1074_), .Y(_1070_) );
XOR2X1 XOR2X1_9 ( .gnd(gnd), .vdd(vdd), .A(up_counter_contador_0_), .B(up_counter_contador_1_), .Y(_1068_) );
DFFPOSX1 DFFPOSX1_17 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf3), .D(_1067_), .Q(memoria_q_0_) );
DFFPOSX1 DFFPOSX1_18 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf2), .D(_1068_), .Q(memoria_q_1_) );
DFFPOSX1 DFFPOSX1_19 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf2), .D(_1069_), .Q(memoria_q_2_) );
DFFPOSX1 DFFPOSX1_20 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf2), .D(_1070_), .Q(memoria_q_3_) );
INVX1 INVX1_406 ( .gnd(gnd), .vdd(vdd), .A(asr1_cables_0__0_), .Y(_1078_) );
NAND2X1 NAND2X1_255 ( .gnd(gnd), .vdd(vdd), .A(din[0]), .B(vdd), .Y(_1079_) );
OAI21X1 OAI21X1_244 ( .gnd(gnd), .vdd(vdd), .A(vdd), .B(_1078_), .C(_1079_), .Y(_1076__0_) );
INVX1 INVX1_407 ( .gnd(gnd), .vdd(vdd), .A(asr1_cables_0__1_), .Y(_1080_) );
NAND2X1 NAND2X1_256 ( .gnd(gnd), .vdd(vdd), .A(vdd), .B(din[1]), .Y(_1081_) );
OAI21X1 OAI21X1_245 ( .gnd(gnd), .vdd(vdd), .A(vdd), .B(_1080_), .C(_1081_), .Y(_1076__1_) );
INVX1 INVX1_408 ( .gnd(gnd), .vdd(vdd), .A(asr1_cables_0__2_), .Y(_1082_) );
NAND2X1 NAND2X1_257 ( .gnd(gnd), .vdd(vdd), .A(vdd), .B(din[2]), .Y(_1083_) );
OAI21X1 OAI21X1_246 ( .gnd(gnd), .vdd(vdd), .A(vdd), .B(_1082_), .C(_1083_), .Y(_1076__2_) );
INVX1 INVX1_409 ( .gnd(gnd), .vdd(vdd), .A(asr1_cables_0__3_), .Y(_1084_) );
NAND2X1 NAND2X1_258 ( .gnd(gnd), .vdd(vdd), .A(vdd), .B(din[3]), .Y(_1085_) );
OAI21X1 OAI21X1_247 ( .gnd(gnd), .vdd(vdd), .A(vdd), .B(_1084_), .C(_1085_), .Y(_1076__3_) );
INVX1 INVX1_410 ( .gnd(gnd), .vdd(vdd), .A(asr1_cables_0__4_), .Y(_1086_) );
NAND2X1 NAND2X1_259 ( .gnd(gnd), .vdd(vdd), .A(vdd), .B(din[4]), .Y(_1087_) );
OAI21X1 OAI21X1_248 ( .gnd(gnd), .vdd(vdd), .A(vdd), .B(_1086_), .C(_1087_), .Y(_1076__4_) );
INVX1 INVX1_411 ( .gnd(gnd), .vdd(vdd), .A(asr1_cables_0__5_), .Y(_1088_) );
NAND2X1 NAND2X1_260 ( .gnd(gnd), .vdd(vdd), .A(vdd), .B(din[5]), .Y(_1089_) );
OAI21X1 OAI21X1_249 ( .gnd(gnd), .vdd(vdd), .A(vdd), .B(_1088_), .C(_1089_), .Y(_1076__5_) );
INVX1 INVX1_412 ( .gnd(gnd), .vdd(vdd), .A(asr1_cables_0__6_), .Y(_1090_) );
NAND2X1 NAND2X1_261 ( .gnd(gnd), .vdd(vdd), .A(vdd), .B(din[6]), .Y(_1091_) );
OAI21X1 OAI21X1_250 ( .gnd(gnd), .vdd(vdd), .A(vdd), .B(_1090_), .C(_1091_), .Y(_1076__6_) );
INVX1 INVX1_413 ( .gnd(gnd), .vdd(vdd), .A(asr1_cables_0__7_), .Y(_1092_) );
NAND2X1 NAND2X1_262 ( .gnd(gnd), .vdd(vdd), .A(vdd), .B(din[7]), .Y(_1093_) );
OAI21X1 OAI21X1_251 ( .gnd(gnd), .vdd(vdd), .A(vdd), .B(_1092_), .C(_1093_), .Y(_1076__7_) );
INVX1 INVX1_414 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf0), .Y(_1077_) );
DFFSR DFFSR_176 ( .gnd(gnd), .vdd(vdd), .CLK(asr1_clk_bF_buf4), .D(_1076__0_), .Q(asr1_cables_0__0_), .R(_1077_), .S(vdd) );
DFFSR DFFSR_177 ( .gnd(gnd), .vdd(vdd), .CLK(asr1_clk_bF_buf0), .D(_1076__1_), .Q(asr1_cables_0__1_), .R(_1077_), .S(vdd) );
DFFSR DFFSR_178 ( .gnd(gnd), .vdd(vdd), .CLK(asr1_clk_bF_buf2), .D(_1076__2_), .Q(asr1_cables_0__2_), .R(_1077_), .S(vdd) );
DFFSR DFFSR_179 ( .gnd(gnd), .vdd(vdd), .CLK(asr1_clk_bF_buf8), .D(_1076__3_), .Q(asr1_cables_0__3_), .R(_1077_), .S(vdd) );
DFFSR DFFSR_180 ( .gnd(gnd), .vdd(vdd), .CLK(asr1_clk_bF_buf8), .D(_1076__4_), .Q(asr1_cables_0__4_), .R(_1077_), .S(vdd) );
DFFSR DFFSR_181 ( .gnd(gnd), .vdd(vdd), .CLK(asr1_clk_bF_buf8), .D(_1076__5_), .Q(asr1_cables_0__5_), .R(_1077_), .S(vdd) );
DFFSR DFFSR_182 ( .gnd(gnd), .vdd(vdd), .CLK(asr1_clk_bF_buf6), .D(_1076__6_), .Q(asr1_cables_0__6_), .R(_1077_), .S(vdd) );
DFFSR DFFSR_183 ( .gnd(gnd), .vdd(vdd), .CLK(asr1_clk_bF_buf4), .D(_1076__7_), .Q(asr1_cables_0__7_), .R(_1077_), .S(vdd) );
INVX1 INVX1_415 ( .gnd(gnd), .vdd(vdd), .A(_3__0_), .Y(_1096_) );
NAND2X1 NAND2X1_263 ( .gnd(gnd), .vdd(vdd), .A(registro_salida_d_0_), .B(vdd), .Y(_1097_) );
OAI21X1 OAI21X1_252 ( .gnd(gnd), .vdd(vdd), .A(vdd), .B(_1096_), .C(_1097_), .Y(_1094__0_) );
INVX1 INVX1_416 ( .gnd(gnd), .vdd(vdd), .A(_3__1_), .Y(_1098_) );
NAND2X1 NAND2X1_264 ( .gnd(gnd), .vdd(vdd), .A(vdd), .B(registro_salida_d_1_), .Y(_1099_) );
OAI21X1 OAI21X1_253 ( .gnd(gnd), .vdd(vdd), .A(vdd), .B(_1098_), .C(_1099_), .Y(_1094__1_) );
INVX1 INVX1_417 ( .gnd(gnd), .vdd(vdd), .A(_3__2_), .Y(_1100_) );
NAND2X1 NAND2X1_265 ( .gnd(gnd), .vdd(vdd), .A(vdd), .B(registro_salida_d_2_), .Y(_1101_) );
OAI21X1 OAI21X1_254 ( .gnd(gnd), .vdd(vdd), .A(vdd), .B(_1100_), .C(_1101_), .Y(_1094__2_) );
INVX1 INVX1_418 ( .gnd(gnd), .vdd(vdd), .A(_3__3_), .Y(_1102_) );
NAND2X1 NAND2X1_266 ( .gnd(gnd), .vdd(vdd), .A(vdd), .B(registro_salida_d_3_), .Y(_1103_) );
OAI21X1 OAI21X1_255 ( .gnd(gnd), .vdd(vdd), .A(vdd), .B(_1102_), .C(_1103_), .Y(_1094__3_) );
INVX1 INVX1_419 ( .gnd(gnd), .vdd(vdd), .A(_3__4_), .Y(_1104_) );
NAND2X1 NAND2X1_267 ( .gnd(gnd), .vdd(vdd), .A(vdd), .B(registro_salida_d_4_), .Y(_1105_) );
OAI21X1 OAI21X1_256 ( .gnd(gnd), .vdd(vdd), .A(vdd), .B(_1104_), .C(_1105_), .Y(_1094__4_) );
INVX1 INVX1_420 ( .gnd(gnd), .vdd(vdd), .A(_3__5_), .Y(_1106_) );
NAND2X1 NAND2X1_268 ( .gnd(gnd), .vdd(vdd), .A(vdd), .B(registro_salida_d_5_), .Y(_1107_) );
OAI21X1 OAI21X1_257 ( .gnd(gnd), .vdd(vdd), .A(vdd), .B(_1106_), .C(_1107_), .Y(_1094__5_) );
INVX1 INVX1_421 ( .gnd(gnd), .vdd(vdd), .A(_3__6_), .Y(_1108_) );
NAND2X1 NAND2X1_269 ( .gnd(gnd), .vdd(vdd), .A(vdd), .B(registro_salida_d_6_), .Y(_1109_) );
OAI21X1 OAI21X1_258 ( .gnd(gnd), .vdd(vdd), .A(vdd), .B(_1108_), .C(_1109_), .Y(_1094__6_) );
INVX1 INVX1_422 ( .gnd(gnd), .vdd(vdd), .A(_3__7_), .Y(_1110_) );
NAND2X1 NAND2X1_270 ( .gnd(gnd), .vdd(vdd), .A(vdd), .B(registro_salida_d_7_), .Y(_1111_) );
OAI21X1 OAI21X1_259 ( .gnd(gnd), .vdd(vdd), .A(vdd), .B(_1110_), .C(_1111_), .Y(_1094__7_) );
INVX1 INVX1_423 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf0), .Y(_1095_) );
DFFSR DFFSR_184 ( .gnd(gnd), .vdd(vdd), .CLK(asr1_clk_bF_buf0), .D(_1094__0_), .Q(_3__0_), .R(_1095_), .S(vdd) );
DFFSR DFFSR_185 ( .gnd(gnd), .vdd(vdd), .CLK(asr1_clk_bF_buf0), .D(_1094__1_), .Q(_3__1_), .R(_1095_), .S(vdd) );
DFFSR DFFSR_186 ( .gnd(gnd), .vdd(vdd), .CLK(asr1_clk_bF_buf0), .D(_1094__2_), .Q(_3__2_), .R(_1095_), .S(vdd) );
DFFSR DFFSR_187 ( .gnd(gnd), .vdd(vdd), .CLK(asr1_clk_bF_buf0), .D(_1094__3_), .Q(_3__3_), .R(_1095_), .S(vdd) );
DFFSR DFFSR_188 ( .gnd(gnd), .vdd(vdd), .CLK(asr1_clk_bF_buf0), .D(_1094__4_), .Q(_3__4_), .R(_1095_), .S(vdd) );
DFFSR DFFSR_189 ( .gnd(gnd), .vdd(vdd), .CLK(asr1_clk_bF_buf0), .D(_1094__5_), .Q(_3__5_), .R(_1095_), .S(vdd) );
DFFSR DFFSR_190 ( .gnd(gnd), .vdd(vdd), .CLK(asr1_clk_bF_buf0), .D(_1094__6_), .Q(_3__6_), .R(_1095_), .S(vdd) );
DFFSR DFFSR_191 ( .gnd(gnd), .vdd(vdd), .CLK(asr1_clk_bF_buf0), .D(_1094__7_), .Q(_3__7_), .R(_1095_), .S(vdd) );
NAND2X1 NAND2X1_271 ( .gnd(gnd), .vdd(vdd), .A(retardo_asr_1_connect_wire_1__0_), .B(retardo_asr_2_connect_wire_1__0_), .Y(_1112_) );
NOR2X1 NOR2X1_46 ( .gnd(gnd), .vdd(vdd), .A(retardo_asr_1_connect_wire_1__1_), .B(retardo_asr_2_connect_wire_1__1_), .Y(_1113_) );
INVX1 INVX1_424 ( .gnd(gnd), .vdd(vdd), .A(_1113_), .Y(_1114_) );
NAND2X1 NAND2X1_272 ( .gnd(gnd), .vdd(vdd), .A(retardo_asr_1_connect_wire_1__1_), .B(retardo_asr_2_connect_wire_1__1_), .Y(_1115_) );
NAND2X1 NAND2X1_273 ( .gnd(gnd), .vdd(vdd), .A(_1115_), .B(_1114_), .Y(_1116_) );
XOR2X1 XOR2X1_10 ( .gnd(gnd), .vdd(vdd), .A(_1116_), .B(_1112_), .Y(sumador_suma_previa_1_) );
OAI21X1 OAI21X1_260 ( .gnd(gnd), .vdd(vdd), .A(_1112_), .B(_1113_), .C(_1115_), .Y(_1117_) );
XOR2X1 XOR2X1_11 ( .gnd(gnd), .vdd(vdd), .A(retardo_asr_1_connect_wire_1__2_), .B(retardo_asr_2_connect_wire_1__2_), .Y(_1118_) );
XOR2X1 XOR2X1_12 ( .gnd(gnd), .vdd(vdd), .A(_1117_), .B(_1118_), .Y(sumador_suma_previa_2_) );
AND2X2 AND2X2_15 ( .gnd(gnd), .vdd(vdd), .A(retardo_asr_1_connect_wire_1__2_), .B(retardo_asr_2_connect_wire_1__2_), .Y(_1119_) );
AOI21X1 AOI21X1_43 ( .gnd(gnd), .vdd(vdd), .A(_1117_), .B(_1118_), .C(_1119_), .Y(_1120_) );
XOR2X1 XOR2X1_13 ( .gnd(gnd), .vdd(vdd), .A(retardo_asr_1_connect_wire_1__3_), .B(retardo_asr_2_connect_wire_1__3_), .Y(_1121_) );
XNOR2X1 XNOR2X1_4 ( .gnd(gnd), .vdd(vdd), .A(_1120_), .B(_1121_), .Y(sumador_suma_previa_3_) );
NAND3X1 NAND3X1_132 ( .gnd(gnd), .vdd(vdd), .A(_1118_), .B(_1121_), .C(_1117_), .Y(_1122_) );
INVX1 INVX1_425 ( .gnd(gnd), .vdd(vdd), .A(retardo_asr_1_connect_wire_1__3_), .Y(_1123_) );
INVX1 INVX1_426 ( .gnd(gnd), .vdd(vdd), .A(retardo_asr_2_connect_wire_1__3_), .Y(_1124_) );
NAND2X1 NAND2X1_274 ( .gnd(gnd), .vdd(vdd), .A(_1123_), .B(_1124_), .Y(_1125_) );
NOR2X1 NOR2X1_47 ( .gnd(gnd), .vdd(vdd), .A(_1123_), .B(_1124_), .Y(_1126_) );
AOI21X1 AOI21X1_44 ( .gnd(gnd), .vdd(vdd), .A(_1119_), .B(_1125_), .C(_1126_), .Y(_1127_) );
NAND2X1 NAND2X1_275 ( .gnd(gnd), .vdd(vdd), .A(_1127_), .B(_1122_), .Y(_1128_) );
INVX1 INVX1_427 ( .gnd(gnd), .vdd(vdd), .A(retardo_asr_1_connect_wire_1__4_), .Y(_1129_) );
INVX1 INVX1_428 ( .gnd(gnd), .vdd(vdd), .A(retardo_asr_2_connect_wire_1__4_), .Y(_1130_) );
NAND2X1 NAND2X1_276 ( .gnd(gnd), .vdd(vdd), .A(_1129_), .B(_1130_), .Y(_1131_) );
NAND2X1 NAND2X1_277 ( .gnd(gnd), .vdd(vdd), .A(retardo_asr_1_connect_wire_1__4_), .B(retardo_asr_2_connect_wire_1__4_), .Y(_1132_) );
AND2X2 AND2X2_16 ( .gnd(gnd), .vdd(vdd), .A(_1131_), .B(_1132_), .Y(_1133_) );
XOR2X1 XOR2X1_14 ( .gnd(gnd), .vdd(vdd), .A(_1128_), .B(_1133_), .Y(sumador_suma_previa_4_) );
AND2X2 AND2X2_17 ( .gnd(gnd), .vdd(vdd), .A(_1122_), .B(_1127_), .Y(_1134_) );
NAND2X1 NAND2X1_278 ( .gnd(gnd), .vdd(vdd), .A(_1132_), .B(_1131_), .Y(_1135_) );
OAI21X1 OAI21X1_261 ( .gnd(gnd), .vdd(vdd), .A(_1135_), .B(_1134_), .C(_1132_), .Y(_1136_) );
INVX1 INVX1_429 ( .gnd(gnd), .vdd(vdd), .A(retardo_asr_1_connect_wire_1__5_), .Y(_1137_) );
INVX1 INVX1_430 ( .gnd(gnd), .vdd(vdd), .A(retardo_asr_2_connect_wire_1__5_), .Y(_1138_) );
NOR2X1 NOR2X1_48 ( .gnd(gnd), .vdd(vdd), .A(_1137_), .B(_1138_), .Y(_1139_) );
NOR2X1 NOR2X1_49 ( .gnd(gnd), .vdd(vdd), .A(retardo_asr_1_connect_wire_1__5_), .B(retardo_asr_2_connect_wire_1__5_), .Y(_1140_) );
NOR2X1 NOR2X1_50 ( .gnd(gnd), .vdd(vdd), .A(_1140_), .B(_1139_), .Y(_1141_) );
XOR2X1 XOR2X1_15 ( .gnd(gnd), .vdd(vdd), .A(_1136_), .B(_1141_), .Y(sumador_suma_previa_5_) );
NOR3X1 NOR3X1_2 ( .gnd(gnd), .vdd(vdd), .A(_1139_), .B(_1140_), .C(_1135_), .Y(_1142_) );
NAND2X1 NAND2X1_279 ( .gnd(gnd), .vdd(vdd), .A(_1142_), .B(_1128_), .Y(_1143_) );
INVX1 INVX1_431 ( .gnd(gnd), .vdd(vdd), .A(_1132_), .Y(_1144_) );
AOI21X1 AOI21X1_45 ( .gnd(gnd), .vdd(vdd), .A(_1141_), .B(_1144_), .C(_1139_), .Y(_1145_) );
INVX1 INVX1_432 ( .gnd(gnd), .vdd(vdd), .A(retardo_asr_1_connect_wire_1__6_), .Y(_1146_) );
NAND2X1 NAND2X1_280 ( .gnd(gnd), .vdd(vdd), .A(retardo_asr_2_connect_wire_1__6_), .B(_1146_), .Y(_1147_) );
INVX1 INVX1_433 ( .gnd(gnd), .vdd(vdd), .A(retardo_asr_2_connect_wire_1__6_), .Y(_1148_) );
NAND2X1 NAND2X1_281 ( .gnd(gnd), .vdd(vdd), .A(retardo_asr_1_connect_wire_1__6_), .B(_1148_), .Y(_1149_) );
AOI22X1 AOI22X1_14 ( .gnd(gnd), .vdd(vdd), .A(_1147_), .B(_1149_), .C(_1143_), .D(_1145_), .Y(_1150_) );
NAND2X1 NAND2X1_282 ( .gnd(gnd), .vdd(vdd), .A(_1133_), .B(_1141_), .Y(_1151_) );
OAI21X1 OAI21X1_262 ( .gnd(gnd), .vdd(vdd), .A(_1151_), .B(_1134_), .C(_1145_), .Y(_1152_) );
NAND2X1 NAND2X1_283 ( .gnd(gnd), .vdd(vdd), .A(_1147_), .B(_1149_), .Y(_1153_) );
NOR2X1 NOR2X1_51 ( .gnd(gnd), .vdd(vdd), .A(_1153_), .B(_1152_), .Y(_1154_) );
NOR2X1 NOR2X1_52 ( .gnd(gnd), .vdd(vdd), .A(_1150_), .B(_1154_), .Y(sumador_suma_previa_6_) );
NOR2X1 NOR2X1_53 ( .gnd(gnd), .vdd(vdd), .A(_1146_), .B(_1148_), .Y(_1155_) );
XOR2X1 XOR2X1_16 ( .gnd(gnd), .vdd(vdd), .A(retardo_asr_1_connect_wire_1__7_), .B(retardo_asr_2_connect_wire_1__7_), .Y(_1156_) );
INVX1 INVX1_434 ( .gnd(gnd), .vdd(vdd), .A(_1156_), .Y(_1157_) );
OAI21X1 OAI21X1_263 ( .gnd(gnd), .vdd(vdd), .A(_1155_), .B(_1150_), .C(_1157_), .Y(_1158_) );
INVX1 INVX1_435 ( .gnd(gnd), .vdd(vdd), .A(_1155_), .Y(_1159_) );
AOI21X1 AOI21X1_46 ( .gnd(gnd), .vdd(vdd), .A(_1122_), .B(_1127_), .C(_1151_), .Y(_1160_) );
INVX1 INVX1_436 ( .gnd(gnd), .vdd(vdd), .A(_1145_), .Y(_1161_) );
OAI21X1 OAI21X1_264 ( .gnd(gnd), .vdd(vdd), .A(_1161_), .B(_1160_), .C(_1153_), .Y(_1162_) );
NAND3X1 NAND3X1_133 ( .gnd(gnd), .vdd(vdd), .A(_1159_), .B(_1156_), .C(_1162_), .Y(_1163_) );
NAND2X1 NAND2X1_284 ( .gnd(gnd), .vdd(vdd), .A(_1163_), .B(_1158_), .Y(sumador_suma_previa_7_) );
XOR2X1 XOR2X1_17 ( .gnd(gnd), .vdd(vdd), .A(retardo_asr_1_connect_wire_1__0_), .B(retardo_asr_2_connect_wire_1__0_), .Y(sumador_suma_previa_0_) );
DFFPOSX1 DFFPOSX1_21 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf3), .D(sumador_suma_previa_0_), .Q(MAC_Adder_0_) );
DFFPOSX1 DFFPOSX1_22 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf3), .D(sumador_suma_previa_1_), .Q(MAC_Adder_1_) );
DFFPOSX1 DFFPOSX1_23 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf6), .D(sumador_suma_previa_2_), .Q(MAC_Adder_2_) );
DFFPOSX1 DFFPOSX1_24 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf6), .D(sumador_suma_previa_3_), .Q(MAC_Adder_3_) );
DFFPOSX1 DFFPOSX1_25 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf6), .D(sumador_suma_previa_4_), .Q(MAC_Adder_4_) );
DFFPOSX1 DFFPOSX1_26 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf6), .D(sumador_suma_previa_5_), .Q(MAC_Adder_5_) );
DFFPOSX1 DFFPOSX1_27 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf6), .D(sumador_suma_previa_6_), .Q(MAC_Adder_6_) );
DFFPOSX1 DFFPOSX1_28 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf6), .D(sumador_suma_previa_7_), .Q(MAC_Adder_7_) );
NOR2X1 NOR2X1_54 ( .gnd(gnd), .vdd(vdd), .A(up_counter_contador_0_), .B(rst_bF_buf5), .Y(_1164__0_) );
INVX1 INVX1_437 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf1), .Y(_1170_) );
OAI21X1 OAI21X1_265 ( .gnd(gnd), .vdd(vdd), .A(up_counter_contador_0_), .B(up_counter_contador_1_), .C(_1170_), .Y(_1165_) );
AOI21X1 AOI21X1_47 ( .gnd(gnd), .vdd(vdd), .A(up_counter_contador_0_), .B(up_counter_contador_1_), .C(_1165_), .Y(_1164__1_) );
NAND2X1 NAND2X1_285 ( .gnd(gnd), .vdd(vdd), .A(up_counter_contador_0_), .B(up_counter_contador_1_), .Y(_1166_) );
NAND2X1 NAND2X1_286 ( .gnd(gnd), .vdd(vdd), .A(up_counter_contador_2_), .B(_1166_), .Y(_1167_) );
INVX1 INVX1_438 ( .gnd(gnd), .vdd(vdd), .A(up_counter_contador_2_), .Y(_1168_) );
NAND3X1 NAND3X1_134 ( .gnd(gnd), .vdd(vdd), .A(up_counter_contador_0_), .B(up_counter_contador_1_), .C(_1168_), .Y(_1169_) );
AOI21X1 AOI21X1_48 ( .gnd(gnd), .vdd(vdd), .A(_1169_), .B(_1167_), .C(rst_bF_buf2), .Y(_1164__2_) );
DFFPOSX1 DFFPOSX1_29 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf4), .D(_1164__0_), .Q(up_counter_contador_0_) );
DFFPOSX1 DFFPOSX1_30 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf2), .D(_1164__1_), .Q(up_counter_contador_1_) );
DFFPOSX1 DFFPOSX1_31 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf2), .D(_1164__2_), .Q(up_counter_contador_2_) );
BUFX2 BUFX2_34 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(MAC_salida_correcta_8_) );
BUFX2 BUFX2_35 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(MAC_salida_correcta_9_) );
BUFX2 BUFX2_36 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(MAC_salida_correcta_10_) );
BUFX2 BUFX2_37 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(MAC_salida_correcta_11_) );
BUFX2 BUFX2_38 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(MAC_salida_correcta_12_) );
BUFX2 BUFX2_39 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(MAC_salida_correcta_13_) );
BUFX2 BUFX2_40 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(MAC_salida_correcta_14_) );
BUFX2 BUFX2_41 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(MAC_salida_correcta_15_) );
BUFX2 BUFX2_42 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(MAC_salida_correcta_16_) );
BUFX2 BUFX2_43 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(MAC_salida_correcta_17_) );
FILL FILL_0_0_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_0_0_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_0_0_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_0_1_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_0_1_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_0_1_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_0_2_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_0_2_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_0_2_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_1_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_1_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_1_0_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_1_0_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_1_0_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_1_1_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_1_1_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_1_1_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_1_2_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_1_2_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_1_2_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_2_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_2_0_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_2_0_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_2_0_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_2_1_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_2_1_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_2_1_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_2_2_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_2_2_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_2_2_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_3_0_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_3_0_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_3_0_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_3_1_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_3_1_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_3_1_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_3_2_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_3_2_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_3_2_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_4_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_4_0_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_4_0_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_4_0_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_4_1_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_4_1_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_4_1_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_4_2_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_4_2_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_4_2_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_5_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_5_0_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_5_0_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_5_0_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_5_1_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_5_1_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_5_1_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_5_2_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_5_2_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_5_2_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_6_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_6_0_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_6_0_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_6_0_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_6_1_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_6_1_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_6_1_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_6_2_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_6_2_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_6_2_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_7_0_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_7_0_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_7_0_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_7_1_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_7_1_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_7_1_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_7_2_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_7_2_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_7_2_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_8_0_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_8_0_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_8_0_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_8_1_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_8_1_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_8_1_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_8_2_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_8_2_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_8_2_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_9_0_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_9_0_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_9_0_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_9_1_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_9_1_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_9_1_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_9_2_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_9_2_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_9_2_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_10_0_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_10_0_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_10_0_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_10_1_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_10_1_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_10_1_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_10_2_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_10_2_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_10_2_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_11_0_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_11_0_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_11_0_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_11_1_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_11_1_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_11_1_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_11_2_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_11_2_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_11_2_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_12_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_12_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_12_0_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_12_0_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_12_0_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_12_1_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_12_1_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_12_1_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_12_2_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_12_2_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_12_2_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_13_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_13_0_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_13_0_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_13_0_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_13_1_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_13_1_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_13_1_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_13_2_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_13_2_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_13_2_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_14_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_14_0_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_14_0_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_14_0_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_14_1_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_14_1_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_14_1_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_14_2_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_14_2_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_14_2_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_15_0_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_15_0_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_15_0_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_15_1_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_15_1_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_15_1_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_15_2_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_15_2_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_15_2_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_16_0_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_16_0_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_16_0_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_16_1_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_16_1_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_16_1_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_16_2_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_16_2_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_16_2_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_17_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_17_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_17_0_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_17_0_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_17_0_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_17_1_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_17_1_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_17_1_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_17_2_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_17_2_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_17_2_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_18_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_18_0_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_18_0_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_18_0_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_18_1_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_18_1_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_18_1_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_18_2_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_18_2_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_18_2_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_19_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_19_0_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_19_0_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_19_0_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_19_1_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_19_1_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_19_1_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_19_2_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_19_2_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_19_2_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_20_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_20_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_20_0_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_20_0_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_20_0_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_20_1_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_20_1_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_20_1_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_20_2_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_20_2_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_20_2_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_21_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_21_0_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_21_0_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_21_0_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_21_1_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_21_1_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_21_1_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_21_2_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_21_2_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_21_2_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_22_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_22_0_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_22_0_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_22_0_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_22_1_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_22_1_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_22_1_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_22_2_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_22_2_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_22_2_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_23_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_23_0_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_23_0_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_23_0_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_23_1_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_23_1_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_23_1_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_23_2_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_23_2_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_23_2_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_24_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_24_0_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_24_0_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_24_0_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_24_1_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_24_1_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_24_1_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_24_2_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_24_2_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_24_2_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_25_0_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_25_0_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_25_0_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_25_1_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_25_1_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_25_1_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_25_2_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_25_2_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_25_2_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_26_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_26_0_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_26_0_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_26_0_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_26_1_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_26_1_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_26_1_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_26_2_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_26_2_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_26_2_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_27_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_27_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_0_0_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_0_0_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_0_0_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_0_1_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_0_1_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_0_1_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_0_2_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_0_2_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_0_2_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_1_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_1_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_1_0_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_1_0_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_1_0_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_1_1_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_1_1_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_1_1_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_1_2_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_1_2_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_1_2_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_2_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_2_0_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_2_0_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_2_0_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_2_1_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_2_1_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_2_1_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_2_2_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_2_2_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_2_2_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_3_0_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_3_0_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_3_0_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_3_1_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_3_1_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_3_1_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_3_2_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_3_2_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_3_2_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_4_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_4_0_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_4_0_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_4_0_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_4_1_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_4_1_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_4_1_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_4_2_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_4_2_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_4_2_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_5_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_5_0_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_5_0_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_5_0_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_5_1_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_5_1_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_5_1_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_5_2_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_5_2_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_5_2_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_6_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_6_0_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_6_0_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_6_0_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_6_1_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_6_1_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_6_1_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_6_2_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_6_2_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_6_2_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_7_0_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_7_0_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_7_0_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_7_1_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_7_1_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_7_1_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_7_2_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_7_2_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_7_2_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_8_0_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_8_0_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_8_0_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_8_1_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_8_1_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_8_1_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_8_2_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_8_2_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_8_2_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_9_0_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_9_0_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_9_0_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_9_1_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_9_1_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_9_1_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_9_2_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_9_2_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_9_2_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_10_0_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_10_0_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_10_0_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_10_1_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_10_1_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_10_1_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_10_2_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_10_2_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_10_2_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_11_0_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_11_0_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_11_0_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_11_1_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_11_1_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_11_1_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_11_2_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_11_2_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_11_2_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_12_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_12_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_12_0_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_12_0_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_12_0_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_12_1_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_12_1_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_12_1_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_12_2_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_12_2_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_12_2_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_13_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_13_0_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_13_0_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_13_0_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_13_1_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_13_1_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_13_1_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_13_2_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_13_2_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_13_2_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_14_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_14_0_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_14_0_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_14_0_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_14_1_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_14_1_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_14_1_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_14_2_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_14_2_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_14_2_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_15_0_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_15_0_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_15_0_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_15_1_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_15_1_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_15_1_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_15_2_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_15_2_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_15_2_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_16_0_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_16_0_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_16_0_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_16_1_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_16_1_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_16_1_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_16_2_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_16_2_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_16_2_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_17_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_17_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_17_0_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_17_0_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_17_0_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_17_1_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_17_1_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_17_1_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_17_2_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_17_2_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_17_2_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_18_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_18_0_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_18_0_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_18_0_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_18_1_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_18_1_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_18_1_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_18_2_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_18_2_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_18_2_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_19_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_19_0_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_19_0_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_19_0_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_19_1_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_19_1_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_19_1_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_19_2_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_19_2_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_19_2_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_20_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_20_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_20_0_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_20_0_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_20_0_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_20_1_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_20_1_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_20_1_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_20_2_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_20_2_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_20_2_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_21_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_21_0_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_21_0_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_21_0_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_21_1_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_21_1_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_21_1_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_21_2_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_21_2_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_21_2_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_22_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_22_0_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_22_0_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_22_0_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_22_1_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_22_1_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_22_1_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_22_2_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_22_2_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_22_2_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_23_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_23_0_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_23_0_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_23_0_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_23_1_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_23_1_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_23_1_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_23_2_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_23_2_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_23_2_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_24_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_24_0_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_24_0_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_24_0_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_24_1_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_24_1_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_24_1_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_24_2_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_24_2_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_24_2_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_25_0_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_25_0_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_25_0_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_25_1_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_25_1_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_25_1_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_25_2_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_25_2_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_25_2_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_26_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_26_0_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_26_0_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_26_0_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_26_1_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_26_1_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_26_1_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_26_2_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_26_2_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_26_2_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_27_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_27_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_0_0_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_0_0_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_0_0_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_0_1_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_0_1_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_0_1_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_0_2_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_0_2_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_0_2_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_1_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_1_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_1_0_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_1_0_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_1_0_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_1_1_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_1_1_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_1_1_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_1_2_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_1_2_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_1_2_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_2_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_2_0_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_2_0_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_2_0_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_2_1_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_2_1_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_2_1_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_2_2_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_2_2_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_2_2_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_3_0_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_3_0_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_3_0_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_3_1_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_3_1_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_3_1_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_3_2_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_3_2_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_3_2_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_4_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_4_0_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_4_0_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_4_0_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_4_1_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_4_1_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_4_1_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_4_2_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_4_2_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_4_2_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_5_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_5_0_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_5_0_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_5_0_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_5_1_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_5_1_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_5_1_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_5_2_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_5_2_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_5_2_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_6_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_6_0_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_6_0_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_6_0_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_6_1_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_6_1_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_6_1_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_6_2_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_6_2_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_6_2_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_7_0_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_7_0_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_7_0_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_7_1_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_7_1_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_7_1_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_7_2_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_7_2_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_7_2_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_8_0_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_8_0_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_8_0_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_8_1_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_8_1_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_8_1_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_8_2_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_8_2_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_8_2_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_9_0_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_9_0_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_9_0_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_9_1_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_9_1_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_9_1_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_9_2_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_9_2_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_9_2_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_10_0_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_10_0_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_10_0_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_10_1_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_10_1_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_10_1_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_10_2_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_10_2_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_10_2_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_11_0_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_11_0_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_11_0_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_11_1_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_11_1_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_11_1_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_11_2_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_11_2_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_11_2_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_12_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_12_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_12_0_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_12_0_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_12_0_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_12_1_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_12_1_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_12_1_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_12_2_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_12_2_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_12_2_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_13_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_13_0_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_13_0_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_13_0_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_13_1_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_13_1_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_13_1_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_13_2_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_13_2_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_13_2_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_14_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_14_0_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_14_0_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_14_0_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_14_1_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_14_1_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_14_1_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_14_2_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_14_2_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_14_2_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_15_0_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_15_0_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_15_0_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_15_1_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_15_1_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_15_1_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_15_2_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_15_2_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_15_2_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_16_0_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_16_0_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_16_0_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_16_1_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_16_1_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_16_1_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_16_2_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_16_2_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_16_2_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_17_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_17_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_17_0_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_17_0_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_17_0_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_17_1_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_17_1_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_17_1_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_17_2_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_17_2_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_17_2_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_18_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_18_0_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_18_0_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_18_0_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_18_1_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_18_1_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_18_1_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_18_2_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_18_2_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_18_2_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_19_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_19_0_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_19_0_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_19_0_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_19_1_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_19_1_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_19_1_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_19_2_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_19_2_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_19_2_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_20_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_20_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_20_0_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_20_0_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_20_0_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_20_1_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_20_1_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_20_1_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_20_2_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_20_2_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_20_2_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_21_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_21_0_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_21_0_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_21_0_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_21_1_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_21_1_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_21_1_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_21_2_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_21_2_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_21_2_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_22_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_22_0_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_22_0_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_22_0_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_22_1_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_22_1_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_22_1_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_22_2_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_22_2_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_22_2_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_23_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_23_0_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_23_0_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_23_0_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_23_1_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_23_1_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_23_1_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_23_2_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_23_2_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_23_2_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_24_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_24_0_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_24_0_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_24_0_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_24_1_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_24_1_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_24_1_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_24_2_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_24_2_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_24_2_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_25_0_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_25_0_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_25_0_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_25_1_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_25_1_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_25_1_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_25_2_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_25_2_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_25_2_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_26_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_26_0_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_26_0_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_26_0_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_26_1_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_26_1_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_26_1_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_26_2_0 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_26_2_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_26_2_2 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_27_1 ( .vdd(vdd), .gnd(gnd) );
FILL FILL_27_2 ( .vdd(vdd), .gnd(gnd) );
endmodule
