module FIR (clk, rst, din, dout);

input clk;
input rst;
input [7:0] din;
output [7:0] dout;

wire vdd = 1'b1;
wire gnd = 1'b0;

CLKBUF1 CLKBUF1_1 ( .A(asr2_clk), .Y(asr2_clk_bF_buf7) );
CLKBUF1 CLKBUF1_2 ( .A(asr2_clk), .Y(asr2_clk_bF_buf6) );
CLKBUF1 CLKBUF1_3 ( .A(asr2_clk), .Y(asr2_clk_bF_buf5) );
CLKBUF1 CLKBUF1_4 ( .A(asr2_clk), .Y(asr2_clk_bF_buf4) );
CLKBUF1 CLKBUF1_5 ( .A(asr2_clk), .Y(asr2_clk_bF_buf3) );
CLKBUF1 CLKBUF1_6 ( .A(asr2_clk), .Y(asr2_clk_bF_buf2) );
CLKBUF1 CLKBUF1_7 ( .A(asr2_clk), .Y(asr2_clk_bF_buf1) );
CLKBUF1 CLKBUF1_8 ( .A(asr2_clk), .Y(asr2_clk_bF_buf0) );
CLKBUF1 CLKBUF1_9 ( .A(clk), .Y(clk_bF_buf7) );
CLKBUF1 CLKBUF1_10 ( .A(clk), .Y(clk_bF_buf6) );
CLKBUF1 CLKBUF1_11 ( .A(clk), .Y(clk_bF_buf5) );
CLKBUF1 CLKBUF1_12 ( .A(clk), .Y(clk_bF_buf4) );
CLKBUF1 CLKBUF1_13 ( .A(clk), .Y(clk_bF_buf3) );
CLKBUF1 CLKBUF1_14 ( .A(clk), .Y(clk_bF_buf2) );
CLKBUF1 CLKBUF1_15 ( .A(clk), .Y(clk_bF_buf1) );
CLKBUF1 CLKBUF1_16 ( .A(clk), .Y(clk_bF_buf0) );
BUFX2 BUFX2_1 ( .A(MAC_clr), .Y(MAC_clr_bF_buf3) );
BUFX2 BUFX2_2 ( .A(MAC_clr), .Y(MAC_clr_bF_buf2) );
BUFX2 BUFX2_3 ( .A(MAC_clr), .Y(MAC_clr_bF_buf1) );
BUFX2 BUFX2_4 ( .A(MAC_clr), .Y(MAC_clr_bF_buf0) );
CLKBUF1 CLKBUF1_17 ( .A(asr1_clk), .Y(asr1_clk_bF_buf8) );
CLKBUF1 CLKBUF1_18 ( .A(asr1_clk), .Y(asr1_clk_bF_buf7) );
CLKBUF1 CLKBUF1_19 ( .A(asr1_clk), .Y(asr1_clk_bF_buf6) );
CLKBUF1 CLKBUF1_20 ( .A(asr1_clk), .Y(asr1_clk_bF_buf5) );
CLKBUF1 CLKBUF1_21 ( .A(asr1_clk), .Y(asr1_clk_bF_buf4) );
CLKBUF1 CLKBUF1_22 ( .A(asr1_clk), .Y(asr1_clk_bF_buf3) );
CLKBUF1 CLKBUF1_23 ( .A(asr1_clk), .Y(asr1_clk_bF_buf2) );
CLKBUF1 CLKBUF1_24 ( .A(asr1_clk), .Y(asr1_clk_bF_buf1) );
CLKBUF1 CLKBUF1_25 ( .A(asr1_clk), .Y(asr1_clk_bF_buf0) );
BUFX2 BUFX2_5 ( .A(rst), .Y(rst_bF_buf5) );
BUFX2 BUFX2_6 ( .A(rst), .Y(rst_bF_buf4) );
BUFX2 BUFX2_7 ( .A(rst), .Y(rst_bF_buf3) );
BUFX2 BUFX2_8 ( .A(rst), .Y(rst_bF_buf2) );
BUFX2 BUFX2_9 ( .A(rst), .Y(rst_bF_buf1) );
BUFX2 BUFX2_10 ( .A(rst), .Y(rst_bF_buf0) );
BUFX2 BUFX2_11 ( .A(MAC_ROM_0_), .Y(MAC_ROM_0_bF_buf3_) );
BUFX2 BUFX2_12 ( .A(MAC_ROM_0_), .Y(MAC_ROM_0_bF_buf2_) );
BUFX2 BUFX2_13 ( .A(MAC_ROM_0_), .Y(MAC_ROM_0_bF_buf1_) );
BUFX2 BUFX2_14 ( .A(MAC_ROM_0_), .Y(MAC_ROM_0_bF_buf0_) );
BUFX2 BUFX2_15 ( .A(asr2_en), .Y(asr2_en_bF_buf10) );
BUFX2 BUFX2_16 ( .A(asr2_en), .Y(asr2_en_bF_buf9) );
BUFX2 BUFX2_17 ( .A(asr2_en), .Y(asr2_en_bF_buf8) );
BUFX2 BUFX2_18 ( .A(asr2_en), .Y(asr2_en_bF_buf7) );
BUFX2 BUFX2_19 ( .A(asr2_en), .Y(asr2_en_bF_buf6) );
BUFX2 BUFX2_20 ( .A(asr2_en), .Y(asr2_en_bF_buf5) );
BUFX2 BUFX2_21 ( .A(asr2_en), .Y(asr2_en_bF_buf4) );
BUFX2 BUFX2_22 ( .A(asr2_en), .Y(asr2_en_bF_buf3) );
BUFX2 BUFX2_23 ( .A(asr2_en), .Y(asr2_en_bF_buf2) );
BUFX2 BUFX2_24 ( .A(asr2_en), .Y(asr2_en_bF_buf1) );
BUFX2 BUFX2_25 ( .A(asr2_en), .Y(asr2_en_bF_buf0) );
NOR2X1 NOR2X1_1 ( .A(up_counter_contador_1_), .B(up_counter_contador_0_), .Y(_1_) );
NOR2X1 NOR2X1_2 ( .A(up_counter_contador_2_), .B(rst_bF_buf3), .Y(_2_) );
AND2X2 AND2X2_1 ( .A(_1_), .B(_2_), .Y(_0_) );
INVX1 INVX1_1 ( .A(asr1_clk_bF_buf0), .Y(asr2_en) );
BUFX2 BUFX2_26 ( .A(_3__0_), .Y(dout[0]) );
BUFX2 BUFX2_27 ( .A(_3__1_), .Y(dout[1]) );
BUFX2 BUFX2_28 ( .A(_3__2_), .Y(dout[2]) );
BUFX2 BUFX2_29 ( .A(_3__3_), .Y(dout[3]) );
BUFX2 BUFX2_30 ( .A(_3__4_), .Y(dout[4]) );
BUFX2 BUFX2_31 ( .A(_3__5_), .Y(dout[5]) );
BUFX2 BUFX2_32 ( .A(_3__6_), .Y(dout[6]) );
BUFX2 BUFX2_33 ( .A(_3__7_), .Y(dout[7]) );
DFFPOSX1 DFFPOSX1_1 ( .CLK(clk_bF_buf4), .D(_0_), .Q(enable_asr) );
INVX1 INVX1_2 ( .A(asr1_cables_1__0_), .Y(_6_) );
NAND2X1 NAND2X1_1 ( .A(asr1_cables_0__0_), .B(vdd), .Y(_7_) );
OAI21X1 OAI21X1_1 ( .A(vdd), .B(_6_), .C(_7_), .Y(_4__0_) );
INVX1 INVX1_3 ( .A(asr1_cables_1__1_), .Y(_8_) );
NAND2X1 NAND2X1_2 ( .A(vdd), .B(asr1_cables_0__1_), .Y(_9_) );
OAI21X1 OAI21X1_2 ( .A(vdd), .B(_8_), .C(_9_), .Y(_4__1_) );
INVX1 INVX1_4 ( .A(asr1_cables_1__2_), .Y(_10_) );
NAND2X1 NAND2X1_3 ( .A(vdd), .B(asr1_cables_0__2_), .Y(_11_) );
OAI21X1 OAI21X1_3 ( .A(vdd), .B(_10_), .C(_11_), .Y(_4__2_) );
INVX1 INVX1_5 ( .A(asr1_cables_1__3_), .Y(_12_) );
NAND2X1 NAND2X1_4 ( .A(vdd), .B(asr1_cables_0__3_), .Y(_13_) );
OAI21X1 OAI21X1_4 ( .A(vdd), .B(_12_), .C(_13_), .Y(_4__3_) );
INVX1 INVX1_6 ( .A(asr1_cables_1__4_), .Y(_14_) );
NAND2X1 NAND2X1_5 ( .A(vdd), .B(asr1_cables_0__4_), .Y(_15_) );
OAI21X1 OAI21X1_5 ( .A(vdd), .B(_14_), .C(_15_), .Y(_4__4_) );
INVX1 INVX1_7 ( .A(asr1_cables_1__5_), .Y(_16_) );
NAND2X1 NAND2X1_6 ( .A(vdd), .B(asr1_cables_0__5_), .Y(_17_) );
OAI21X1 OAI21X1_6 ( .A(vdd), .B(_16_), .C(_17_), .Y(_4__5_) );
INVX1 INVX1_8 ( .A(asr1_cables_1__6_), .Y(_18_) );
NAND2X1 NAND2X1_7 ( .A(vdd), .B(asr1_cables_0__6_), .Y(_19_) );
OAI21X1 OAI21X1_7 ( .A(vdd), .B(_18_), .C(_19_), .Y(_4__6_) );
INVX1 INVX1_9 ( .A(asr1_cables_1__7_), .Y(_20_) );
NAND2X1 NAND2X1_8 ( .A(vdd), .B(asr1_cables_0__7_), .Y(_21_) );
OAI21X1 OAI21X1_8 ( .A(vdd), .B(_20_), .C(_21_), .Y(_4__7_) );
INVX1 INVX1_10 ( .A(rst_bF_buf0), .Y(_5_) );
DFFSR DFFSR_1 ( .CLK(asr1_clk_bF_buf6), .D(_4__0_), .Q(asr1_cables_1__0_), .R(_5_), .S(vdd) );
DFFSR DFFSR_2 ( .CLK(asr1_clk_bF_buf2), .D(_4__1_), .Q(asr1_cables_1__1_), .R(_5_), .S(vdd) );
DFFSR DFFSR_3 ( .CLK(asr1_clk_bF_buf7), .D(_4__2_), .Q(asr1_cables_1__2_), .R(_5_), .S(vdd) );
DFFSR DFFSR_4 ( .CLK(asr1_clk_bF_buf7), .D(_4__3_), .Q(asr1_cables_1__3_), .R(_5_), .S(vdd) );
DFFSR DFFSR_5 ( .CLK(asr1_clk_bF_buf2), .D(_4__4_), .Q(asr1_cables_1__4_), .R(_5_), .S(vdd) );
DFFSR DFFSR_6 ( .CLK(asr1_clk_bF_buf0), .D(_4__5_), .Q(asr1_cables_1__5_), .R(_5_), .S(vdd) );
DFFSR DFFSR_7 ( .CLK(asr1_clk_bF_buf2), .D(_4__6_), .Q(asr1_cables_1__6_), .R(_5_), .S(vdd) );
DFFSR DFFSR_8 ( .CLK(asr1_clk_bF_buf0), .D(_4__7_), .Q(asr1_cables_1__7_), .R(_5_), .S(vdd) );
INVX1 INVX1_11 ( .A(asr1_cables_2__0_), .Y(_24_) );
NAND2X1 NAND2X1_9 ( .A(asr1_cables_1__0_), .B(vdd), .Y(_25_) );
OAI21X1 OAI21X1_9 ( .A(vdd), .B(_24_), .C(_25_), .Y(_22__0_) );
INVX1 INVX1_12 ( .A(asr1_cables_2__1_), .Y(_26_) );
NAND2X1 NAND2X1_10 ( .A(vdd), .B(asr1_cables_1__1_), .Y(_27_) );
OAI21X1 OAI21X1_10 ( .A(vdd), .B(_26_), .C(_27_), .Y(_22__1_) );
INVX1 INVX1_13 ( .A(asr1_cables_2__2_), .Y(_28_) );
NAND2X1 NAND2X1_11 ( .A(vdd), .B(asr1_cables_1__2_), .Y(_29_) );
OAI21X1 OAI21X1_11 ( .A(vdd), .B(_28_), .C(_29_), .Y(_22__2_) );
INVX1 INVX1_14 ( .A(asr1_cables_2__3_), .Y(_30_) );
NAND2X1 NAND2X1_12 ( .A(vdd), .B(asr1_cables_1__3_), .Y(_31_) );
OAI21X1 OAI21X1_12 ( .A(vdd), .B(_30_), .C(_31_), .Y(_22__3_) );
INVX1 INVX1_15 ( .A(asr1_cables_2__4_), .Y(_32_) );
NAND2X1 NAND2X1_13 ( .A(vdd), .B(asr1_cables_1__4_), .Y(_33_) );
OAI21X1 OAI21X1_13 ( .A(vdd), .B(_32_), .C(_33_), .Y(_22__4_) );
INVX1 INVX1_16 ( .A(asr1_cables_2__5_), .Y(_34_) );
NAND2X1 NAND2X1_14 ( .A(vdd), .B(asr1_cables_1__5_), .Y(_35_) );
OAI21X1 OAI21X1_14 ( .A(vdd), .B(_34_), .C(_35_), .Y(_22__5_) );
INVX1 INVX1_17 ( .A(asr1_cables_2__6_), .Y(_36_) );
NAND2X1 NAND2X1_15 ( .A(vdd), .B(asr1_cables_1__6_), .Y(_37_) );
OAI21X1 OAI21X1_15 ( .A(vdd), .B(_36_), .C(_37_), .Y(_22__6_) );
INVX1 INVX1_18 ( .A(asr1_cables_2__7_), .Y(_38_) );
NAND2X1 NAND2X1_16 ( .A(vdd), .B(asr1_cables_1__7_), .Y(_39_) );
OAI21X1 OAI21X1_16 ( .A(vdd), .B(_38_), .C(_39_), .Y(_22__7_) );
INVX1 INVX1_19 ( .A(rst_bF_buf2), .Y(_23_) );
DFFSR DFFSR_9 ( .CLK(asr1_clk_bF_buf6), .D(_22__0_), .Q(asr1_cables_2__0_), .R(_23_), .S(vdd) );
DFFSR DFFSR_10 ( .CLK(asr1_clk_bF_buf8), .D(_22__1_), .Q(asr1_cables_2__1_), .R(_23_), .S(vdd) );
DFFSR DFFSR_11 ( .CLK(asr1_clk_bF_buf7), .D(_22__2_), .Q(asr1_cables_2__2_), .R(_23_), .S(vdd) );
DFFSR DFFSR_12 ( .CLK(asr1_clk_bF_buf1), .D(_22__3_), .Q(asr1_cables_2__3_), .R(_23_), .S(vdd) );
DFFSR DFFSR_13 ( .CLK(asr1_clk_bF_buf7), .D(_22__4_), .Q(asr1_cables_2__4_), .R(_23_), .S(vdd) );
DFFSR DFFSR_14 ( .CLK(asr1_clk_bF_buf0), .D(_22__5_), .Q(asr1_cables_2__5_), .R(_23_), .S(vdd) );
DFFSR DFFSR_15 ( .CLK(asr1_clk_bF_buf4), .D(_22__6_), .Q(asr1_cables_2__6_), .R(_23_), .S(vdd) );
DFFSR DFFSR_16 ( .CLK(asr1_clk_bF_buf3), .D(_22__7_), .Q(asr1_cables_2__7_), .R(_23_), .S(vdd) );
INVX1 INVX1_20 ( .A(asr1_cables_3__0_), .Y(_42_) );
NAND2X1 NAND2X1_17 ( .A(asr1_cables_2__0_), .B(vdd), .Y(_43_) );
OAI21X1 OAI21X1_17 ( .A(vdd), .B(_42_), .C(_43_), .Y(_40__0_) );
INVX1 INVX1_21 ( .A(asr1_cables_3__1_), .Y(_44_) );
NAND2X1 NAND2X1_18 ( .A(vdd), .B(asr1_cables_2__1_), .Y(_45_) );
OAI21X1 OAI21X1_18 ( .A(vdd), .B(_44_), .C(_45_), .Y(_40__1_) );
INVX1 INVX1_22 ( .A(asr1_cables_3__2_), .Y(_46_) );
NAND2X1 NAND2X1_19 ( .A(vdd), .B(asr1_cables_2__2_), .Y(_47_) );
OAI21X1 OAI21X1_19 ( .A(vdd), .B(_46_), .C(_47_), .Y(_40__2_) );
INVX1 INVX1_23 ( .A(asr1_cables_3__3_), .Y(_48_) );
NAND2X1 NAND2X1_20 ( .A(vdd), .B(asr1_cables_2__3_), .Y(_49_) );
OAI21X1 OAI21X1_20 ( .A(vdd), .B(_48_), .C(_49_), .Y(_40__3_) );
INVX1 INVX1_24 ( .A(asr1_cables_3__4_), .Y(_50_) );
NAND2X1 NAND2X1_21 ( .A(vdd), .B(asr1_cables_2__4_), .Y(_51_) );
OAI21X1 OAI21X1_21 ( .A(vdd), .B(_50_), .C(_51_), .Y(_40__4_) );
INVX1 INVX1_25 ( .A(asr1_cables_3__5_), .Y(_52_) );
NAND2X1 NAND2X1_22 ( .A(vdd), .B(asr1_cables_2__5_), .Y(_53_) );
OAI21X1 OAI21X1_22 ( .A(vdd), .B(_52_), .C(_53_), .Y(_40__5_) );
INVX1 INVX1_26 ( .A(asr1_cables_3__6_), .Y(_54_) );
NAND2X1 NAND2X1_23 ( .A(vdd), .B(asr1_cables_2__6_), .Y(_55_) );
OAI21X1 OAI21X1_23 ( .A(vdd), .B(_54_), .C(_55_), .Y(_40__6_) );
INVX1 INVX1_27 ( .A(asr1_cables_3__7_), .Y(_56_) );
NAND2X1 NAND2X1_24 ( .A(vdd), .B(asr1_cables_2__7_), .Y(_57_) );
OAI21X1 OAI21X1_24 ( .A(vdd), .B(_56_), .C(_57_), .Y(_40__7_) );
INVX1 INVX1_28 ( .A(rst_bF_buf0), .Y(_41_) );
DFFSR DFFSR_17 ( .CLK(asr1_clk_bF_buf2), .D(_40__0_), .Q(asr1_cables_3__0_), .R(_41_), .S(vdd) );
DFFSR DFFSR_18 ( .CLK(asr1_clk_bF_buf5), .D(_40__1_), .Q(asr1_cables_3__1_), .R(_41_), .S(vdd) );
DFFSR DFFSR_19 ( .CLK(asr1_clk_bF_buf4), .D(_40__2_), .Q(asr1_cables_3__2_), .R(_41_), .S(vdd) );
DFFSR DFFSR_20 ( .CLK(asr1_clk_bF_buf1), .D(_40__3_), .Q(asr1_cables_3__3_), .R(_41_), .S(vdd) );
DFFSR DFFSR_21 ( .CLK(asr1_clk_bF_buf6), .D(_40__4_), .Q(asr1_cables_3__4_), .R(_41_), .S(vdd) );
DFFSR DFFSR_22 ( .CLK(asr1_clk_bF_buf3), .D(_40__5_), .Q(asr1_cables_3__5_), .R(_41_), .S(vdd) );
DFFSR DFFSR_23 ( .CLK(asr1_clk_bF_buf1), .D(_40__6_), .Q(asr1_cables_3__6_), .R(_41_), .S(vdd) );
DFFSR DFFSR_24 ( .CLK(asr1_clk_bF_buf5), .D(_40__7_), .Q(asr1_cables_3__7_), .R(_41_), .S(vdd) );
INVX1 INVX1_29 ( .A(asr1_cables_4_), .Y(_60_) );
NAND2X1 NAND2X1_25 ( .A(asr1_cables_3__0_), .B(vdd), .Y(_61_) );
OAI21X1 OAI21X1_25 ( .A(vdd), .B(_60_), .C(_61_), .Y(_58__0_) );
INVX1 INVX1_30 ( .A(_76_), .Y(_62_) );
NAND2X1 NAND2X1_26 ( .A(vdd), .B(asr1_cables_3__1_), .Y(_63_) );
OAI21X1 OAI21X1_26 ( .A(vdd), .B(_62_), .C(_63_), .Y(_58__1_) );
INVX1 INVX1_31 ( .A(_82_), .Y(_64_) );
NAND2X1 NAND2X1_27 ( .A(vdd), .B(asr1_cables_3__2_), .Y(_65_) );
OAI21X1 OAI21X1_27 ( .A(vdd), .B(_64_), .C(_65_), .Y(_58__2_) );
INVX1 INVX1_32 ( .A(_77_), .Y(_66_) );
NAND2X1 NAND2X1_28 ( .A(vdd), .B(asr1_cables_3__3_), .Y(_67_) );
OAI21X1 OAI21X1_28 ( .A(vdd), .B(_66_), .C(_67_), .Y(_58__3_) );
INVX1 INVX1_33 ( .A(_78_), .Y(_68_) );
NAND2X1 NAND2X1_29 ( .A(vdd), .B(asr1_cables_3__4_), .Y(_69_) );
OAI21X1 OAI21X1_29 ( .A(vdd), .B(_68_), .C(_69_), .Y(_58__4_) );
INVX1 INVX1_34 ( .A(_79_), .Y(_70_) );
NAND2X1 NAND2X1_30 ( .A(vdd), .B(asr1_cables_3__5_), .Y(_71_) );
OAI21X1 OAI21X1_30 ( .A(vdd), .B(_70_), .C(_71_), .Y(_58__5_) );
INVX1 INVX1_35 ( .A(_80_), .Y(_72_) );
NAND2X1 NAND2X1_31 ( .A(vdd), .B(asr1_cables_3__6_), .Y(_73_) );
OAI21X1 OAI21X1_31 ( .A(vdd), .B(_72_), .C(_73_), .Y(_58__6_) );
INVX1 INVX1_36 ( .A(_81_), .Y(_74_) );
NAND2X1 NAND2X1_32 ( .A(vdd), .B(asr1_cables_3__7_), .Y(_75_) );
OAI21X1 OAI21X1_32 ( .A(vdd), .B(_74_), .C(_75_), .Y(_58__7_) );
INVX1 INVX1_37 ( .A(rst_bF_buf0), .Y(_59_) );
DFFSR DFFSR_25 ( .CLK(asr1_clk_bF_buf8), .D(_58__0_), .Q(asr1_cables_4_), .R(_59_), .S(vdd) );
DFFSR DFFSR_26 ( .CLK(asr1_clk_bF_buf5), .D(_58__1_), .Q(_76_), .R(_59_), .S(vdd) );
DFFSR DFFSR_27 ( .CLK(asr1_clk_bF_buf5), .D(_58__2_), .Q(_82_), .R(_59_), .S(vdd) );
DFFSR DFFSR_28 ( .CLK(asr1_clk_bF_buf3), .D(_58__3_), .Q(_77_), .R(_59_), .S(vdd) );
DFFSR DFFSR_29 ( .CLK(asr1_clk_bF_buf4), .D(_58__4_), .Q(_78_), .R(_59_), .S(vdd) );
DFFSR DFFSR_30 ( .CLK(asr1_clk_bF_buf8), .D(_58__5_), .Q(_79_), .R(_59_), .S(vdd) );
DFFSR DFFSR_31 ( .CLK(asr1_clk_bF_buf1), .D(_58__6_), .Q(_80_), .R(_59_), .S(vdd) );
DFFSR DFFSR_32 ( .CLK(asr1_clk_bF_buf5), .D(_58__7_), .Q(_81_), .R(_59_), .S(vdd) );
INVX1 INVX1_38 ( .A(asr1_cables_5__0_), .Y(_85_) );
NAND2X1 NAND2X1_33 ( .A(asr1_cables_4_), .B(vdd), .Y(_86_) );
OAI21X1 OAI21X1_33 ( .A(vdd), .B(_85_), .C(_86_), .Y(_83__0_) );
INVX1 INVX1_39 ( .A(asr1_cables_5__1_), .Y(_87_) );
NAND2X1 NAND2X1_34 ( .A(vdd), .B(_76_), .Y(_88_) );
OAI21X1 OAI21X1_34 ( .A(vdd), .B(_87_), .C(_88_), .Y(_83__1_) );
INVX1 INVX1_40 ( .A(asr1_cables_5__2_), .Y(_89_) );
NAND2X1 NAND2X1_35 ( .A(vdd), .B(_82_), .Y(_90_) );
OAI21X1 OAI21X1_35 ( .A(vdd), .B(_89_), .C(_90_), .Y(_83__2_) );
INVX1 INVX1_41 ( .A(asr1_cables_5__3_), .Y(_91_) );
NAND2X1 NAND2X1_36 ( .A(vdd), .B(_77_), .Y(_92_) );
OAI21X1 OAI21X1_36 ( .A(vdd), .B(_91_), .C(_92_), .Y(_83__3_) );
INVX1 INVX1_42 ( .A(asr1_cables_5__4_), .Y(_93_) );
NAND2X1 NAND2X1_37 ( .A(vdd), .B(_78_), .Y(_94_) );
OAI21X1 OAI21X1_37 ( .A(vdd), .B(_93_), .C(_94_), .Y(_83__4_) );
INVX1 INVX1_43 ( .A(asr1_cables_5__5_), .Y(_95_) );
NAND2X1 NAND2X1_38 ( .A(vdd), .B(_79_), .Y(_96_) );
OAI21X1 OAI21X1_38 ( .A(vdd), .B(_95_), .C(_96_), .Y(_83__5_) );
INVX1 INVX1_44 ( .A(asr1_cables_5__6_), .Y(_97_) );
NAND2X1 NAND2X1_39 ( .A(vdd), .B(_80_), .Y(_98_) );
OAI21X1 OAI21X1_39 ( .A(vdd), .B(_97_), .C(_98_), .Y(_83__6_) );
INVX1 INVX1_45 ( .A(asr1_cables_5__7_), .Y(_99_) );
NAND2X1 NAND2X1_40 ( .A(vdd), .B(_81_), .Y(_100_) );
OAI21X1 OAI21X1_40 ( .A(vdd), .B(_99_), .C(_100_), .Y(_83__7_) );
INVX1 INVX1_46 ( .A(rst_bF_buf0), .Y(_84_) );
DFFSR DFFSR_33 ( .CLK(asr1_clk_bF_buf3), .D(_83__0_), .Q(asr1_cables_5__0_), .R(_84_), .S(vdd) );
DFFSR DFFSR_34 ( .CLK(asr1_clk_bF_buf5), .D(_83__1_), .Q(asr1_cables_5__1_), .R(_84_), .S(vdd) );
DFFSR DFFSR_35 ( .CLK(asr1_clk_bF_buf2), .D(_83__2_), .Q(asr1_cables_5__2_), .R(_84_), .S(vdd) );
DFFSR DFFSR_36 ( .CLK(asr1_clk_bF_buf8), .D(_83__3_), .Q(asr1_cables_5__3_), .R(_84_), .S(vdd) );
DFFSR DFFSR_37 ( .CLK(asr1_clk_bF_buf2), .D(_83__4_), .Q(asr1_cables_5__4_), .R(_84_), .S(vdd) );
DFFSR DFFSR_38 ( .CLK(asr1_clk_bF_buf4), .D(_83__5_), .Q(asr1_cables_5__5_), .R(_84_), .S(vdd) );
DFFSR DFFSR_39 ( .CLK(asr1_clk_bF_buf8), .D(_83__6_), .Q(asr1_cables_5__6_), .R(_84_), .S(vdd) );
DFFSR DFFSR_40 ( .CLK(asr1_clk_bF_buf3), .D(_83__7_), .Q(asr1_cables_5__7_), .R(_84_), .S(vdd) );
INVX1 INVX1_47 ( .A(asr1_cables_6__0_), .Y(_103_) );
NAND2X1 NAND2X1_41 ( .A(asr1_cables_5__0_), .B(vdd), .Y(_104_) );
OAI21X1 OAI21X1_41 ( .A(vdd), .B(_103_), .C(_104_), .Y(_101__0_) );
INVX1 INVX1_48 ( .A(asr1_cables_6__1_), .Y(_105_) );
NAND2X1 NAND2X1_42 ( .A(vdd), .B(asr1_cables_5__1_), .Y(_106_) );
OAI21X1 OAI21X1_42 ( .A(vdd), .B(_105_), .C(_106_), .Y(_101__1_) );
INVX1 INVX1_49 ( .A(asr1_cables_6__2_), .Y(_107_) );
NAND2X1 NAND2X1_43 ( .A(vdd), .B(asr1_cables_5__2_), .Y(_108_) );
OAI21X1 OAI21X1_43 ( .A(vdd), .B(_107_), .C(_108_), .Y(_101__2_) );
INVX1 INVX1_50 ( .A(asr1_cables_6__3_), .Y(_109_) );
NAND2X1 NAND2X1_44 ( .A(vdd), .B(asr1_cables_5__3_), .Y(_110_) );
OAI21X1 OAI21X1_44 ( .A(vdd), .B(_109_), .C(_110_), .Y(_101__3_) );
INVX1 INVX1_51 ( .A(asr1_cables_6__4_), .Y(_111_) );
NAND2X1 NAND2X1_45 ( .A(vdd), .B(asr1_cables_5__4_), .Y(_112_) );
OAI21X1 OAI21X1_45 ( .A(vdd), .B(_111_), .C(_112_), .Y(_101__4_) );
INVX1 INVX1_52 ( .A(asr1_cables_6__5_), .Y(_113_) );
NAND2X1 NAND2X1_46 ( .A(vdd), .B(asr1_cables_5__5_), .Y(_114_) );
OAI21X1 OAI21X1_46 ( .A(vdd), .B(_113_), .C(_114_), .Y(_101__5_) );
INVX1 INVX1_53 ( .A(asr1_cables_6__6_), .Y(_115_) );
NAND2X1 NAND2X1_47 ( .A(vdd), .B(asr1_cables_5__6_), .Y(_116_) );
OAI21X1 OAI21X1_47 ( .A(vdd), .B(_115_), .C(_116_), .Y(_101__6_) );
INVX1 INVX1_54 ( .A(asr1_cables_6__7_), .Y(_117_) );
NAND2X1 NAND2X1_48 ( .A(vdd), .B(asr1_cables_5__7_), .Y(_118_) );
OAI21X1 OAI21X1_48 ( .A(vdd), .B(_117_), .C(_118_), .Y(_101__7_) );
INVX1 INVX1_55 ( .A(rst_bF_buf3), .Y(_102_) );
DFFSR DFFSR_41 ( .CLK(asr1_clk_bF_buf2), .D(_101__0_), .Q(asr1_cables_6__0_), .R(_102_), .S(vdd) );
DFFSR DFFSR_42 ( .CLK(asr1_clk_bF_buf5), .D(_101__1_), .Q(asr1_cables_6__1_), .R(_102_), .S(vdd) );
DFFSR DFFSR_43 ( .CLK(asr1_clk_bF_buf8), .D(_101__2_), .Q(asr1_cables_6__2_), .R(_102_), .S(vdd) );
DFFSR DFFSR_44 ( .CLK(asr1_clk_bF_buf8), .D(_101__3_), .Q(asr1_cables_6__3_), .R(_102_), .S(vdd) );
DFFSR DFFSR_45 ( .CLK(asr1_clk_bF_buf8), .D(_101__4_), .Q(asr1_cables_6__4_), .R(_102_), .S(vdd) );
DFFSR DFFSR_46 ( .CLK(asr1_clk_bF_buf0), .D(_101__5_), .Q(asr1_cables_6__5_), .R(_102_), .S(vdd) );
DFFSR DFFSR_47 ( .CLK(asr1_clk_bF_buf3), .D(_101__6_), .Q(asr1_cables_6__6_), .R(_102_), .S(vdd) );
DFFSR DFFSR_48 ( .CLK(asr1_clk_bF_buf5), .D(_101__7_), .Q(asr1_cables_6__7_), .R(_102_), .S(vdd) );
INVX1 INVX1_56 ( .A(asr1_cables_7__0_), .Y(_121_) );
NAND2X1 NAND2X1_49 ( .A(asr1_cables_6__0_), .B(vdd), .Y(_122_) );
OAI21X1 OAI21X1_49 ( .A(vdd), .B(_121_), .C(_122_), .Y(_119__0_) );
INVX1 INVX1_57 ( .A(asr1_cables_7__1_), .Y(_123_) );
NAND2X1 NAND2X1_50 ( .A(vdd), .B(asr1_cables_6__1_), .Y(_124_) );
OAI21X1 OAI21X1_50 ( .A(vdd), .B(_123_), .C(_124_), .Y(_119__1_) );
INVX1 INVX1_58 ( .A(asr1_cables_7__2_), .Y(_125_) );
NAND2X1 NAND2X1_51 ( .A(vdd), .B(asr1_cables_6__2_), .Y(_126_) );
OAI21X1 OAI21X1_51 ( .A(vdd), .B(_125_), .C(_126_), .Y(_119__2_) );
INVX1 INVX1_59 ( .A(asr1_cables_7__3_), .Y(_127_) );
NAND2X1 NAND2X1_52 ( .A(vdd), .B(asr1_cables_6__3_), .Y(_128_) );
OAI21X1 OAI21X1_52 ( .A(vdd), .B(_127_), .C(_128_), .Y(_119__3_) );
INVX1 INVX1_60 ( .A(asr1_cables_7__4_), .Y(_129_) );
NAND2X1 NAND2X1_53 ( .A(vdd), .B(asr1_cables_6__4_), .Y(_130_) );
OAI21X1 OAI21X1_53 ( .A(vdd), .B(_129_), .C(_130_), .Y(_119__4_) );
INVX1 INVX1_61 ( .A(asr1_cables_7__5_), .Y(_131_) );
NAND2X1 NAND2X1_54 ( .A(vdd), .B(asr1_cables_6__5_), .Y(_132_) );
OAI21X1 OAI21X1_54 ( .A(vdd), .B(_131_), .C(_132_), .Y(_119__5_) );
INVX1 INVX1_62 ( .A(asr1_cables_7__6_), .Y(_133_) );
NAND2X1 NAND2X1_55 ( .A(vdd), .B(asr1_cables_6__6_), .Y(_134_) );
OAI21X1 OAI21X1_55 ( .A(vdd), .B(_133_), .C(_134_), .Y(_119__6_) );
INVX1 INVX1_63 ( .A(asr1_cables_7__7_), .Y(_135_) );
NAND2X1 NAND2X1_56 ( .A(vdd), .B(asr1_cables_6__7_), .Y(_136_) );
OAI21X1 OAI21X1_56 ( .A(vdd), .B(_135_), .C(_136_), .Y(_119__7_) );
INVX1 INVX1_64 ( .A(rst_bF_buf3), .Y(_120_) );
DFFSR DFFSR_49 ( .CLK(asr1_clk_bF_buf2), .D(_119__0_), .Q(asr1_cables_7__0_), .R(_120_), .S(vdd) );
DFFSR DFFSR_50 ( .CLK(asr1_clk_bF_buf4), .D(_119__1_), .Q(asr1_cables_7__1_), .R(_120_), .S(vdd) );
DFFSR DFFSR_51 ( .CLK(asr1_clk_bF_buf4), .D(_119__2_), .Q(asr1_cables_7__2_), .R(_120_), .S(vdd) );
DFFSR DFFSR_52 ( .CLK(asr1_clk_bF_buf8), .D(_119__3_), .Q(asr1_cables_7__3_), .R(_120_), .S(vdd) );
DFFSR DFFSR_53 ( .CLK(asr1_clk_bF_buf8), .D(_119__4_), .Q(asr1_cables_7__4_), .R(_120_), .S(vdd) );
DFFSR DFFSR_54 ( .CLK(asr1_clk_bF_buf0), .D(_119__5_), .Q(asr1_cables_7__5_), .R(_120_), .S(vdd) );
DFFSR DFFSR_55 ( .CLK(asr1_clk_bF_buf3), .D(_119__6_), .Q(asr1_cables_7__6_), .R(_120_), .S(vdd) );
DFFSR DFFSR_56 ( .CLK(asr1_clk_bF_buf5), .D(_119__7_), .Q(asr1_cables_7__7_), .R(_120_), .S(vdd) );
INVX1 INVX1_65 ( .A(asr1_cables_8__0_), .Y(_139_) );
NAND2X1 NAND2X1_57 ( .A(asr1_cables_7__0_), .B(vdd), .Y(_140_) );
OAI21X1 OAI21X1_57 ( .A(vdd), .B(_139_), .C(_140_), .Y(_137__0_) );
INVX1 INVX1_66 ( .A(asr1_cables_8__1_), .Y(_141_) );
NAND2X1 NAND2X1_58 ( .A(vdd), .B(asr1_cables_7__1_), .Y(_142_) );
OAI21X1 OAI21X1_58 ( .A(vdd), .B(_141_), .C(_142_), .Y(_137__1_) );
INVX1 INVX1_67 ( .A(asr1_cables_8__2_), .Y(_143_) );
NAND2X1 NAND2X1_59 ( .A(vdd), .B(asr1_cables_7__2_), .Y(_144_) );
OAI21X1 OAI21X1_59 ( .A(vdd), .B(_143_), .C(_144_), .Y(_137__2_) );
INVX1 INVX1_68 ( .A(asr1_cables_8__3_), .Y(_145_) );
NAND2X1 NAND2X1_60 ( .A(vdd), .B(asr1_cables_7__3_), .Y(_146_) );
OAI21X1 OAI21X1_60 ( .A(vdd), .B(_145_), .C(_146_), .Y(_137__3_) );
INVX1 INVX1_69 ( .A(asr1_cables_8__4_), .Y(_147_) );
NAND2X1 NAND2X1_61 ( .A(vdd), .B(asr1_cables_7__4_), .Y(_148_) );
OAI21X1 OAI21X1_61 ( .A(vdd), .B(_147_), .C(_148_), .Y(_137__4_) );
INVX1 INVX1_70 ( .A(asr1_cables_8__5_), .Y(_149_) );
NAND2X1 NAND2X1_62 ( .A(vdd), .B(asr1_cables_7__5_), .Y(_150_) );
OAI21X1 OAI21X1_62 ( .A(vdd), .B(_149_), .C(_150_), .Y(_137__5_) );
INVX1 INVX1_71 ( .A(asr1_cables_8__6_), .Y(_151_) );
NAND2X1 NAND2X1_63 ( .A(vdd), .B(asr1_cables_7__6_), .Y(_152_) );
OAI21X1 OAI21X1_63 ( .A(vdd), .B(_151_), .C(_152_), .Y(_137__6_) );
INVX1 INVX1_72 ( .A(asr1_cables_8__7_), .Y(_153_) );
NAND2X1 NAND2X1_64 ( .A(vdd), .B(asr1_cables_7__7_), .Y(_154_) );
OAI21X1 OAI21X1_64 ( .A(vdd), .B(_153_), .C(_154_), .Y(_137__7_) );
INVX1 INVX1_73 ( .A(rst_bF_buf0), .Y(_138_) );
DFFSR DFFSR_57 ( .CLK(asr1_clk_bF_buf2), .D(_137__0_), .Q(asr1_cables_8__0_), .R(_138_), .S(vdd) );
DFFSR DFFSR_58 ( .CLK(asr1_clk_bF_buf4), .D(_137__1_), .Q(asr1_cables_8__1_), .R(_138_), .S(vdd) );
DFFSR DFFSR_59 ( .CLK(asr1_clk_bF_buf4), .D(_137__2_), .Q(asr1_cables_8__2_), .R(_138_), .S(vdd) );
DFFSR DFFSR_60 ( .CLK(asr1_clk_bF_buf0), .D(_137__3_), .Q(asr1_cables_8__3_), .R(_138_), .S(vdd) );
DFFSR DFFSR_61 ( .CLK(asr1_clk_bF_buf1), .D(_137__4_), .Q(asr1_cables_8__4_), .R(_138_), .S(vdd) );
DFFSR DFFSR_62 ( .CLK(asr1_clk_bF_buf3), .D(_137__5_), .Q(asr1_cables_8__5_), .R(_138_), .S(vdd) );
DFFSR DFFSR_63 ( .CLK(asr1_clk_bF_buf3), .D(_137__6_), .Q(asr1_cables_8__6_), .R(_138_), .S(vdd) );
DFFSR DFFSR_64 ( .CLK(asr1_clk_bF_buf4), .D(_137__7_), .Q(asr1_cables_8__7_), .R(_138_), .S(vdd) );
INVX1 INVX1_74 ( .A(asr2_cables_1__0_), .Y(_157_) );
NAND2X1 NAND2X1_65 ( .A(asr1_q_0_), .B(asr2_en_bF_buf1), .Y(_158_) );
OAI21X1 OAI21X1_65 ( .A(asr2_en_bF_buf1), .B(_157_), .C(_158_), .Y(_155__0_) );
INVX1 INVX1_75 ( .A(asr2_cables_1__1_), .Y(_159_) );
NAND2X1 NAND2X1_66 ( .A(asr2_en_bF_buf1), .B(asr1_q_1_), .Y(_160_) );
OAI21X1 OAI21X1_66 ( .A(asr2_en_bF_buf10), .B(_159_), .C(_160_), .Y(_155__1_) );
INVX1 INVX1_76 ( .A(asr2_cables_1__2_), .Y(_161_) );
NAND2X1 NAND2X1_67 ( .A(asr2_en_bF_buf1), .B(asr1_q_2_), .Y(_162_) );
OAI21X1 OAI21X1_67 ( .A(asr2_en_bF_buf1), .B(_161_), .C(_162_), .Y(_155__2_) );
INVX1 INVX1_77 ( .A(asr2_cables_1__3_), .Y(_163_) );
NAND2X1 NAND2X1_68 ( .A(asr2_en_bF_buf2), .B(asr1_q_3_), .Y(_164_) );
OAI21X1 OAI21X1_68 ( .A(asr2_en_bF_buf2), .B(_163_), .C(_164_), .Y(_155__3_) );
INVX1 INVX1_78 ( .A(asr2_cables_1__4_), .Y(_165_) );
NAND2X1 NAND2X1_69 ( .A(asr2_en_bF_buf2), .B(asr1_q_4_), .Y(_166_) );
OAI21X1 OAI21X1_69 ( .A(asr2_en_bF_buf2), .B(_165_), .C(_166_), .Y(_155__4_) );
INVX1 INVX1_79 ( .A(asr2_cables_1__5_), .Y(_167_) );
NAND2X1 NAND2X1_70 ( .A(asr2_en_bF_buf8), .B(asr1_q_5_), .Y(_168_) );
OAI21X1 OAI21X1_70 ( .A(asr2_en_bF_buf8), .B(_167_), .C(_168_), .Y(_155__5_) );
INVX1 INVX1_80 ( .A(asr2_cables_1__6_), .Y(_169_) );
NAND2X1 NAND2X1_71 ( .A(asr2_en_bF_buf2), .B(asr1_q_6_), .Y(_170_) );
OAI21X1 OAI21X1_71 ( .A(asr2_en_bF_buf6), .B(_169_), .C(_170_), .Y(_155__6_) );
INVX1 INVX1_81 ( .A(asr2_cables_1__7_), .Y(_171_) );
NAND2X1 NAND2X1_72 ( .A(asr2_en_bF_buf8), .B(asr1_q_7_), .Y(_172_) );
OAI21X1 OAI21X1_72 ( .A(asr2_en_bF_buf8), .B(_171_), .C(_172_), .Y(_155__7_) );
INVX1 INVX1_82 ( .A(rst_bF_buf5), .Y(_156_) );
DFFSR DFFSR_65 ( .CLK(asr2_clk_bF_buf5), .D(_155__0_), .Q(asr2_cables_1__0_), .R(_156_), .S(vdd) );
DFFSR DFFSR_66 ( .CLK(asr2_clk_bF_buf3), .D(_155__1_), .Q(asr2_cables_1__1_), .R(_156_), .S(vdd) );
DFFSR DFFSR_67 ( .CLK(asr2_clk_bF_buf6), .D(_155__2_), .Q(asr2_cables_1__2_), .R(_156_), .S(vdd) );
DFFSR DFFSR_68 ( .CLK(asr2_clk_bF_buf0), .D(_155__3_), .Q(asr2_cables_1__3_), .R(_156_), .S(vdd) );
DFFSR DFFSR_69 ( .CLK(asr2_clk_bF_buf0), .D(_155__4_), .Q(asr2_cables_1__4_), .R(_156_), .S(vdd) );
DFFSR DFFSR_70 ( .CLK(asr2_clk_bF_buf5), .D(_155__5_), .Q(asr2_cables_1__5_), .R(_156_), .S(vdd) );
DFFSR DFFSR_71 ( .CLK(asr2_clk_bF_buf7), .D(_155__6_), .Q(asr2_cables_1__6_), .R(_156_), .S(vdd) );
DFFSR DFFSR_72 ( .CLK(asr2_clk_bF_buf5), .D(_155__7_), .Q(asr2_cables_1__7_), .R(_156_), .S(vdd) );
INVX1 INVX1_83 ( .A(asr2_cables_2__0_), .Y(_175_) );
NAND2X1 NAND2X1_73 ( .A(asr2_cables_1__0_), .B(asr2_en_bF_buf9), .Y(_176_) );
OAI21X1 OAI21X1_73 ( .A(asr2_en_bF_buf9), .B(_175_), .C(_176_), .Y(_173__0_) );
INVX1 INVX1_84 ( .A(asr2_cables_2__1_), .Y(_177_) );
NAND2X1 NAND2X1_74 ( .A(asr2_en_bF_buf7), .B(asr2_cables_1__1_), .Y(_178_) );
OAI21X1 OAI21X1_74 ( .A(asr2_en_bF_buf7), .B(_177_), .C(_178_), .Y(_173__1_) );
INVX1 INVX1_85 ( .A(asr2_cables_2__2_), .Y(_179_) );
NAND2X1 NAND2X1_75 ( .A(asr2_en_bF_buf1), .B(asr2_cables_1__2_), .Y(_180_) );
OAI21X1 OAI21X1_75 ( .A(asr2_en_bF_buf7), .B(_179_), .C(_180_), .Y(_173__2_) );
INVX1 INVX1_86 ( .A(asr2_cables_2__3_), .Y(_181_) );
NAND2X1 NAND2X1_76 ( .A(asr2_en_bF_buf6), .B(asr2_cables_1__3_), .Y(_182_) );
OAI21X1 OAI21X1_76 ( .A(asr2_en_bF_buf6), .B(_181_), .C(_182_), .Y(_173__3_) );
INVX1 INVX1_87 ( .A(asr2_cables_2__4_), .Y(_183_) );
NAND2X1 NAND2X1_77 ( .A(asr2_en_bF_buf2), .B(asr2_cables_1__4_), .Y(_184_) );
OAI21X1 OAI21X1_77 ( .A(asr2_en_bF_buf8), .B(_183_), .C(_184_), .Y(_173__4_) );
INVX1 INVX1_88 ( .A(asr2_cables_2__5_), .Y(_185_) );
NAND2X1 NAND2X1_78 ( .A(asr2_en_bF_buf9), .B(asr2_cables_1__5_), .Y(_186_) );
OAI21X1 OAI21X1_78 ( .A(asr2_en_bF_buf7), .B(_185_), .C(_186_), .Y(_173__5_) );
INVX1 INVX1_89 ( .A(asr2_cables_2__6_), .Y(_187_) );
NAND2X1 NAND2X1_79 ( .A(asr2_en_bF_buf3), .B(asr2_cables_1__6_), .Y(_188_) );
OAI21X1 OAI21X1_79 ( .A(asr2_en_bF_buf3), .B(_187_), .C(_188_), .Y(_173__6_) );
INVX1 INVX1_90 ( .A(asr2_cables_2__7_), .Y(_189_) );
NAND2X1 NAND2X1_80 ( .A(asr2_en_bF_buf9), .B(asr2_cables_1__7_), .Y(_190_) );
OAI21X1 OAI21X1_80 ( .A(asr2_en_bF_buf8), .B(_189_), .C(_190_), .Y(_173__7_) );
INVX1 INVX1_91 ( .A(rst_bF_buf1), .Y(_174_) );
DFFSR DFFSR_73 ( .CLK(asr2_clk_bF_buf4), .D(_173__0_), .Q(asr2_cables_2__0_), .R(_174_), .S(vdd) );
DFFSR DFFSR_74 ( .CLK(asr2_clk_bF_buf3), .D(_173__1_), .Q(asr2_cables_2__1_), .R(_174_), .S(vdd) );
DFFSR DFFSR_75 ( .CLK(asr2_clk_bF_buf6), .D(_173__2_), .Q(asr2_cables_2__2_), .R(_174_), .S(vdd) );
DFFSR DFFSR_76 ( .CLK(asr2_clk_bF_buf2), .D(_173__3_), .Q(asr2_cables_2__3_), .R(_174_), .S(vdd) );
DFFSR DFFSR_77 ( .CLK(asr2_clk_bF_buf5), .D(_173__4_), .Q(asr2_cables_2__4_), .R(_174_), .S(vdd) );
DFFSR DFFSR_78 ( .CLK(asr2_clk_bF_buf3), .D(_173__5_), .Q(asr2_cables_2__5_), .R(_174_), .S(vdd) );
DFFSR DFFSR_79 ( .CLK(asr2_clk_bF_buf7), .D(_173__6_), .Q(asr2_cables_2__6_), .R(_174_), .S(vdd) );
DFFSR DFFSR_80 ( .CLK(asr2_clk_bF_buf5), .D(_173__7_), .Q(asr2_cables_2__7_), .R(_174_), .S(vdd) );
INVX1 INVX1_92 ( .A(asr2_cables_3__0_), .Y(_193_) );
NAND2X1 NAND2X1_81 ( .A(asr2_cables_2__0_), .B(asr2_en_bF_buf6), .Y(_194_) );
OAI21X1 OAI21X1_81 ( .A(asr2_en_bF_buf6), .B(_193_), .C(_194_), .Y(_191__0_) );
INVX1 INVX1_93 ( .A(asr2_cables_3__1_), .Y(_195_) );
NAND2X1 NAND2X1_82 ( .A(asr2_en_bF_buf7), .B(asr2_cables_2__1_), .Y(_196_) );
OAI21X1 OAI21X1_82 ( .A(asr2_en_bF_buf7), .B(_195_), .C(_196_), .Y(_191__1_) );
INVX1 INVX1_94 ( .A(asr2_cables_3__2_), .Y(_197_) );
NAND2X1 NAND2X1_83 ( .A(asr2_en_bF_buf6), .B(asr2_cables_2__2_), .Y(_198_) );
OAI21X1 OAI21X1_83 ( .A(asr2_en_bF_buf6), .B(_197_), .C(_198_), .Y(_191__2_) );
INVX1 INVX1_95 ( .A(asr2_cables_3__3_), .Y(_199_) );
NAND2X1 NAND2X1_84 ( .A(asr2_en_bF_buf5), .B(asr2_cables_2__3_), .Y(_200_) );
OAI21X1 OAI21X1_84 ( .A(asr2_en_bF_buf5), .B(_199_), .C(_200_), .Y(_191__3_) );
INVX1 INVX1_96 ( .A(asr2_cables_3__4_), .Y(_201_) );
NAND2X1 NAND2X1_85 ( .A(asr2_en_bF_buf2), .B(asr2_cables_2__4_), .Y(_202_) );
OAI21X1 OAI21X1_85 ( .A(asr2_en_bF_buf2), .B(_201_), .C(_202_), .Y(_191__4_) );
INVX1 INVX1_97 ( .A(asr2_cables_3__5_), .Y(_203_) );
NAND2X1 NAND2X1_86 ( .A(asr2_en_bF_buf10), .B(asr2_cables_2__5_), .Y(_204_) );
OAI21X1 OAI21X1_86 ( .A(asr2_en_bF_buf10), .B(_203_), .C(_204_), .Y(_191__5_) );
INVX1 INVX1_98 ( .A(asr2_cables_3__6_), .Y(_205_) );
NAND2X1 NAND2X1_87 ( .A(asr2_en_bF_buf3), .B(asr2_cables_2__6_), .Y(_206_) );
OAI21X1 OAI21X1_87 ( .A(asr2_en_bF_buf10), .B(_205_), .C(_206_), .Y(_191__6_) );
INVX1 INVX1_99 ( .A(asr2_cables_3__7_), .Y(_207_) );
NAND2X1 NAND2X1_88 ( .A(asr2_en_bF_buf7), .B(asr2_cables_2__7_), .Y(_208_) );
OAI21X1 OAI21X1_88 ( .A(asr2_en_bF_buf7), .B(_207_), .C(_208_), .Y(_191__7_) );
INVX1 INVX1_100 ( .A(rst_bF_buf2), .Y(_192_) );
DFFSR DFFSR_81 ( .CLK(asr2_clk_bF_buf2), .D(_191__0_), .Q(asr2_cables_3__0_), .R(_192_), .S(vdd) );
DFFSR DFFSR_82 ( .CLK(asr2_clk_bF_buf6), .D(_191__1_), .Q(asr2_cables_3__1_), .R(_192_), .S(vdd) );
DFFSR DFFSR_83 ( .CLK(asr2_clk_bF_buf2), .D(_191__2_), .Q(asr2_cables_3__2_), .R(_192_), .S(vdd) );
DFFSR DFFSR_84 ( .CLK(asr2_clk_bF_buf2), .D(_191__3_), .Q(asr2_cables_3__3_), .R(_192_), .S(vdd) );
DFFSR DFFSR_85 ( .CLK(asr2_clk_bF_buf6), .D(_191__4_), .Q(asr2_cables_3__4_), .R(_192_), .S(vdd) );
DFFSR DFFSR_86 ( .CLK(asr2_clk_bF_buf3), .D(_191__5_), .Q(asr2_cables_3__5_), .R(_192_), .S(vdd) );
DFFSR DFFSR_87 ( .CLK(asr2_clk_bF_buf4), .D(_191__6_), .Q(asr2_cables_3__6_), .R(_192_), .S(vdd) );
DFFSR DFFSR_88 ( .CLK(asr2_clk_bF_buf6), .D(_191__7_), .Q(asr2_cables_3__7_), .R(_192_), .S(vdd) );
INVX1 INVX1_101 ( .A(asr2_cables_4_), .Y(_211_) );
NAND2X1 NAND2X1_89 ( .A(asr2_cables_3__0_), .B(asr2_en_bF_buf5), .Y(_212_) );
OAI21X1 OAI21X1_89 ( .A(asr2_en_bF_buf4), .B(_211_), .C(_212_), .Y(_209__0_) );
INVX1 INVX1_102 ( .A(_227_), .Y(_213_) );
NAND2X1 NAND2X1_90 ( .A(asr2_en_bF_buf7), .B(asr2_cables_3__1_), .Y(_214_) );
OAI21X1 OAI21X1_90 ( .A(asr2_en_bF_buf7), .B(_213_), .C(_214_), .Y(_209__1_) );
INVX1 INVX1_103 ( .A(_233_), .Y(_215_) );
NAND2X1 NAND2X1_91 ( .A(asr2_en_bF_buf0), .B(asr2_cables_3__2_), .Y(_216_) );
OAI21X1 OAI21X1_91 ( .A(asr2_en_bF_buf0), .B(_215_), .C(_216_), .Y(_209__2_) );
INVX1 INVX1_104 ( .A(_228_), .Y(_217_) );
NAND2X1 NAND2X1_92 ( .A(asr2_en_bF_buf5), .B(asr2_cables_3__3_), .Y(_218_) );
OAI21X1 OAI21X1_92 ( .A(asr2_en_bF_buf0), .B(_217_), .C(_218_), .Y(_209__3_) );
INVX1 INVX1_105 ( .A(_229_), .Y(_219_) );
NAND2X1 NAND2X1_93 ( .A(asr2_en_bF_buf7), .B(asr2_cables_3__4_), .Y(_220_) );
OAI21X1 OAI21X1_93 ( .A(asr2_en_bF_buf10), .B(_219_), .C(_220_), .Y(_209__4_) );
INVX1 INVX1_106 ( .A(_230_), .Y(_221_) );
NAND2X1 NAND2X1_94 ( .A(asr2_en_bF_buf9), .B(asr2_cables_3__5_), .Y(_222_) );
OAI21X1 OAI21X1_94 ( .A(asr2_en_bF_buf9), .B(_221_), .C(_222_), .Y(_209__5_) );
INVX1 INVX1_107 ( .A(_231_), .Y(_223_) );
NAND2X1 NAND2X1_95 ( .A(asr2_en_bF_buf3), .B(asr2_cables_3__6_), .Y(_224_) );
OAI21X1 OAI21X1_95 ( .A(asr2_en_bF_buf3), .B(_223_), .C(_224_), .Y(_209__6_) );
INVX1 INVX1_108 ( .A(_232_), .Y(_225_) );
NAND2X1 NAND2X1_96 ( .A(asr2_en_bF_buf10), .B(asr2_cables_3__7_), .Y(_226_) );
OAI21X1 OAI21X1_96 ( .A(asr2_en_bF_buf10), .B(_225_), .C(_226_), .Y(_209__7_) );
INVX1 INVX1_109 ( .A(rst_bF_buf5), .Y(_210_) );
DFFSR DFFSR_89 ( .CLK(asr2_clk_bF_buf1), .D(_209__0_), .Q(asr2_cables_4_), .R(_210_), .S(vdd) );
DFFSR DFFSR_90 ( .CLK(asr2_clk_bF_buf6), .D(_209__1_), .Q(_227_), .R(_210_), .S(vdd) );
DFFSR DFFSR_91 ( .CLK(asr2_clk_bF_buf0), .D(_209__2_), .Q(_233_), .R(_210_), .S(vdd) );
DFFSR DFFSR_92 ( .CLK(asr2_clk_bF_buf0), .D(_209__3_), .Q(_228_), .R(_210_), .S(vdd) );
DFFSR DFFSR_93 ( .CLK(asr2_clk_bF_buf3), .D(_209__4_), .Q(_229_), .R(_210_), .S(vdd) );
DFFSR DFFSR_94 ( .CLK(asr2_clk_bF_buf3), .D(_209__5_), .Q(_230_), .R(_210_), .S(vdd) );
DFFSR DFFSR_95 ( .CLK(asr2_clk_bF_buf7), .D(_209__6_), .Q(_231_), .R(_210_), .S(vdd) );
DFFSR DFFSR_96 ( .CLK(asr2_clk_bF_buf3), .D(_209__7_), .Q(_232_), .R(_210_), .S(vdd) );
INVX1 INVX1_110 ( .A(asr2_cables_5__0_), .Y(_236_) );
NAND2X1 NAND2X1_97 ( .A(asr2_cables_4_), .B(asr2_en_bF_buf5), .Y(_237_) );
OAI21X1 OAI21X1_97 ( .A(asr2_en_bF_buf5), .B(_236_), .C(_237_), .Y(_234__0_) );
INVX1 INVX1_111 ( .A(asr2_cables_5__1_), .Y(_238_) );
NAND2X1 NAND2X1_98 ( .A(asr2_en_bF_buf7), .B(_227_), .Y(_239_) );
OAI21X1 OAI21X1_98 ( .A(asr2_en_bF_buf1), .B(_238_), .C(_239_), .Y(_234__1_) );
INVX1 INVX1_112 ( .A(asr2_cables_5__2_), .Y(_240_) );
NAND2X1 NAND2X1_99 ( .A(asr2_en_bF_buf0), .B(_233_), .Y(_241_) );
OAI21X1 OAI21X1_99 ( .A(asr2_en_bF_buf0), .B(_240_), .C(_241_), .Y(_234__2_) );
INVX1 INVX1_113 ( .A(asr2_cables_5__3_), .Y(_242_) );
NAND2X1 NAND2X1_100 ( .A(asr2_en_bF_buf0), .B(_228_), .Y(_243_) );
OAI21X1 OAI21X1_100 ( .A(asr2_en_bF_buf4), .B(_242_), .C(_243_), .Y(_234__3_) );
INVX1 INVX1_114 ( .A(asr2_cables_5__4_), .Y(_244_) );
NAND2X1 NAND2X1_101 ( .A(asr2_en_bF_buf9), .B(_229_), .Y(_245_) );
OAI21X1 OAI21X1_101 ( .A(asr2_en_bF_buf9), .B(_244_), .C(_245_), .Y(_234__4_) );
INVX1 INVX1_115 ( .A(asr2_cables_5__5_), .Y(_246_) );
NAND2X1 NAND2X1_102 ( .A(asr2_en_bF_buf9), .B(_230_), .Y(_247_) );
OAI21X1 OAI21X1_102 ( .A(asr2_en_bF_buf8), .B(_246_), .C(_247_), .Y(_234__5_) );
INVX1 INVX1_116 ( .A(asr2_cables_5__6_), .Y(_248_) );
NAND2X1 NAND2X1_103 ( .A(asr2_en_bF_buf3), .B(_231_), .Y(_249_) );
OAI21X1 OAI21X1_103 ( .A(asr2_en_bF_buf3), .B(_248_), .C(_249_), .Y(_234__6_) );
INVX1 INVX1_117 ( .A(asr2_cables_5__7_), .Y(_250_) );
NAND2X1 NAND2X1_104 ( .A(asr2_en_bF_buf10), .B(_232_), .Y(_251_) );
OAI21X1 OAI21X1_104 ( .A(asr2_en_bF_buf10), .B(_250_), .C(_251_), .Y(_234__7_) );
INVX1 INVX1_118 ( .A(rst_bF_buf1), .Y(_235_) );
DFFSR DFFSR_97 ( .CLK(asr2_clk_bF_buf1), .D(_234__0_), .Q(asr2_cables_5__0_), .R(_235_), .S(vdd) );
DFFSR DFFSR_98 ( .CLK(asr2_clk_bF_buf6), .D(_234__1_), .Q(asr2_cables_5__1_), .R(_235_), .S(vdd) );
DFFSR DFFSR_99 ( .CLK(asr2_clk_bF_buf0), .D(_234__2_), .Q(asr2_cables_5__2_), .R(_235_), .S(vdd) );
DFFSR DFFSR_100 ( .CLK(asr2_clk_bF_buf0), .D(_234__3_), .Q(asr2_cables_5__3_), .R(_235_), .S(vdd) );
DFFSR DFFSR_101 ( .CLK(asr2_clk_bF_buf4), .D(_234__4_), .Q(asr2_cables_5__4_), .R(_235_), .S(vdd) );
DFFSR DFFSR_102 ( .CLK(asr2_clk_bF_buf5), .D(_234__5_), .Q(asr2_cables_5__5_), .R(_235_), .S(vdd) );
DFFSR DFFSR_103 ( .CLK(asr2_clk_bF_buf4), .D(_234__6_), .Q(asr2_cables_5__6_), .R(_235_), .S(vdd) );
DFFSR DFFSR_104 ( .CLK(asr2_clk_bF_buf3), .D(_234__7_), .Q(asr2_cables_5__7_), .R(_235_), .S(vdd) );
INVX1 INVX1_119 ( .A(asr2_cables_6__0_), .Y(_254_) );
NAND2X1 NAND2X1_105 ( .A(asr2_cables_5__0_), .B(asr2_en_bF_buf4), .Y(_255_) );
OAI21X1 OAI21X1_105 ( .A(asr2_en_bF_buf4), .B(_254_), .C(_255_), .Y(_252__0_) );
INVX1 INVX1_120 ( .A(asr2_cables_6__1_), .Y(_256_) );
NAND2X1 NAND2X1_106 ( .A(asr2_en_bF_buf1), .B(asr2_cables_5__1_), .Y(_257_) );
OAI21X1 OAI21X1_106 ( .A(asr2_en_bF_buf1), .B(_256_), .C(_257_), .Y(_252__1_) );
INVX1 INVX1_121 ( .A(asr2_cables_6__2_), .Y(_258_) );
NAND2X1 NAND2X1_107 ( .A(asr2_en_bF_buf0), .B(asr2_cables_5__2_), .Y(_259_) );
OAI21X1 OAI21X1_107 ( .A(asr2_en_bF_buf0), .B(_258_), .C(_259_), .Y(_252__2_) );
INVX1 INVX1_122 ( .A(asr2_cables_6__3_), .Y(_260_) );
NAND2X1 NAND2X1_108 ( .A(asr2_en_bF_buf2), .B(asr2_cables_5__3_), .Y(_261_) );
OAI21X1 OAI21X1_108 ( .A(asr2_en_bF_buf6), .B(_260_), .C(_261_), .Y(_252__3_) );
INVX1 INVX1_123 ( .A(asr2_cables_6__4_), .Y(_262_) );
NAND2X1 NAND2X1_109 ( .A(asr2_en_bF_buf6), .B(asr2_cables_5__4_), .Y(_263_) );
OAI21X1 OAI21X1_109 ( .A(asr2_en_bF_buf5), .B(_262_), .C(_263_), .Y(_252__4_) );
INVX1 INVX1_124 ( .A(asr2_cables_6__5_), .Y(_264_) );
NAND2X1 NAND2X1_110 ( .A(asr2_en_bF_buf8), .B(asr2_cables_5__5_), .Y(_265_) );
OAI21X1 OAI21X1_110 ( .A(asr2_en_bF_buf1), .B(_264_), .C(_265_), .Y(_252__5_) );
INVX1 INVX1_125 ( .A(asr2_cables_6__6_), .Y(_266_) );
NAND2X1 NAND2X1_111 ( .A(asr2_en_bF_buf3), .B(asr2_cables_5__6_), .Y(_267_) );
OAI21X1 OAI21X1_111 ( .A(asr2_en_bF_buf3), .B(_266_), .C(_267_), .Y(_252__6_) );
INVX1 INVX1_126 ( .A(asr2_cables_6__7_), .Y(_268_) );
NAND2X1 NAND2X1_112 ( .A(asr2_en_bF_buf10), .B(asr2_cables_5__7_), .Y(_269_) );
OAI21X1 OAI21X1_112 ( .A(asr2_en_bF_buf10), .B(_268_), .C(_269_), .Y(_252__7_) );
INVX1 INVX1_127 ( .A(rst_bF_buf2), .Y(_253_) );
DFFSR DFFSR_105 ( .CLK(asr2_clk_bF_buf1), .D(_252__0_), .Q(asr2_cables_6__0_), .R(_253_), .S(vdd) );
DFFSR DFFSR_106 ( .CLK(asr2_clk_bF_buf6), .D(_252__1_), .Q(asr2_cables_6__1_), .R(_253_), .S(vdd) );
DFFSR DFFSR_107 ( .CLK(asr2_clk_bF_buf2), .D(_252__2_), .Q(asr2_cables_6__2_), .R(_253_), .S(vdd) );
DFFSR DFFSR_108 ( .CLK(asr2_clk_bF_buf7), .D(_252__3_), .Q(asr2_cables_6__3_), .R(_253_), .S(vdd) );
DFFSR DFFSR_109 ( .CLK(asr2_clk_bF_buf1), .D(_252__4_), .Q(asr2_cables_6__4_), .R(_253_), .S(vdd) );
DFFSR DFFSR_110 ( .CLK(asr2_clk_bF_buf5), .D(_252__5_), .Q(asr2_cables_6__5_), .R(_253_), .S(vdd) );
DFFSR DFFSR_111 ( .CLK(asr2_clk_bF_buf4), .D(_252__6_), .Q(asr2_cables_6__6_), .R(_253_), .S(vdd) );
DFFSR DFFSR_112 ( .CLK(asr2_clk_bF_buf4), .D(_252__7_), .Q(asr2_cables_6__7_), .R(_253_), .S(vdd) );
INVX1 INVX1_128 ( .A(asr2_cables_7__0_), .Y(_272_) );
NAND2X1 NAND2X1_113 ( .A(asr2_cables_6__0_), .B(asr2_en_bF_buf4), .Y(_273_) );
OAI21X1 OAI21X1_113 ( .A(asr2_en_bF_buf4), .B(_272_), .C(_273_), .Y(_270__0_) );
INVX1 INVX1_129 ( .A(asr2_cables_7__1_), .Y(_274_) );
NAND2X1 NAND2X1_114 ( .A(asr2_en_bF_buf8), .B(asr2_cables_6__1_), .Y(_275_) );
OAI21X1 OAI21X1_114 ( .A(asr2_en_bF_buf3), .B(_274_), .C(_275_), .Y(_270__1_) );
INVX1 INVX1_130 ( .A(asr2_cables_7__2_), .Y(_276_) );
NAND2X1 NAND2X1_115 ( .A(asr2_en_bF_buf0), .B(asr2_cables_6__2_), .Y(_277_) );
OAI21X1 OAI21X1_115 ( .A(asr2_en_bF_buf0), .B(_276_), .C(_277_), .Y(_270__2_) );
INVX1 INVX1_131 ( .A(asr2_cables_7__3_), .Y(_278_) );
NAND2X1 NAND2X1_116 ( .A(asr2_en_bF_buf8), .B(asr2_cables_6__3_), .Y(_279_) );
OAI21X1 OAI21X1_116 ( .A(asr2_en_bF_buf8), .B(_278_), .C(_279_), .Y(_270__3_) );
INVX1 INVX1_132 ( .A(asr2_cables_7__4_), .Y(_280_) );
NAND2X1 NAND2X1_117 ( .A(asr2_en_bF_buf4), .B(asr2_cables_6__4_), .Y(_281_) );
OAI21X1 OAI21X1_117 ( .A(asr2_en_bF_buf4), .B(_280_), .C(_281_), .Y(_270__4_) );
INVX1 INVX1_133 ( .A(asr2_cables_7__5_), .Y(_282_) );
NAND2X1 NAND2X1_118 ( .A(asr2_en_bF_buf1), .B(asr2_cables_6__5_), .Y(_283_) );
OAI21X1 OAI21X1_118 ( .A(asr2_en_bF_buf8), .B(_282_), .C(_283_), .Y(_270__5_) );
INVX1 INVX1_134 ( .A(asr2_cables_7__6_), .Y(_284_) );
NAND2X1 NAND2X1_119 ( .A(asr2_en_bF_buf5), .B(asr2_cables_6__6_), .Y(_285_) );
OAI21X1 OAI21X1_119 ( .A(asr2_en_bF_buf5), .B(_284_), .C(_285_), .Y(_270__6_) );
INVX1 INVX1_135 ( .A(asr2_cables_7__7_), .Y(_286_) );
NAND2X1 NAND2X1_120 ( .A(asr2_en_bF_buf10), .B(asr2_cables_6__7_), .Y(_287_) );
OAI21X1 OAI21X1_120 ( .A(asr2_en_bF_buf9), .B(_286_), .C(_287_), .Y(_270__7_) );
INVX1 INVX1_136 ( .A(rst_bF_buf5), .Y(_271_) );
DFFSR DFFSR_113 ( .CLK(asr2_clk_bF_buf1), .D(_270__0_), .Q(asr2_cables_7__0_), .R(_271_), .S(vdd) );
DFFSR DFFSR_114 ( .CLK(asr2_clk_bF_buf7), .D(_270__1_), .Q(asr2_cables_7__1_), .R(_271_), .S(vdd) );
DFFSR DFFSR_115 ( .CLK(asr2_clk_bF_buf0), .D(_270__2_), .Q(asr2_cables_7__2_), .R(_271_), .S(vdd) );
DFFSR DFFSR_116 ( .CLK(asr2_clk_bF_buf7), .D(_270__3_), .Q(asr2_cables_7__3_), .R(_271_), .S(vdd) );
DFFSR DFFSR_117 ( .CLK(asr2_clk_bF_buf1), .D(_270__4_), .Q(asr2_cables_7__4_), .R(_271_), .S(vdd) );
DFFSR DFFSR_118 ( .CLK(asr2_clk_bF_buf5), .D(_270__5_), .Q(asr2_cables_7__5_), .R(_271_), .S(vdd) );
DFFSR DFFSR_119 ( .CLK(asr2_clk_bF_buf2), .D(_270__6_), .Q(asr2_cables_7__6_), .R(_271_), .S(vdd) );
DFFSR DFFSR_120 ( .CLK(asr2_clk_bF_buf4), .D(_270__7_), .Q(asr2_cables_7__7_), .R(_271_), .S(vdd) );
INVX1 INVX1_137 ( .A(asr2_cables_8__0_), .Y(_290_) );
NAND2X1 NAND2X1_121 ( .A(asr2_cables_7__0_), .B(asr2_en_bF_buf5), .Y(_291_) );
OAI21X1 OAI21X1_121 ( .A(asr2_en_bF_buf5), .B(_290_), .C(_291_), .Y(_288__0_) );
INVX1 INVX1_138 ( .A(asr2_cables_8__1_), .Y(_292_) );
NAND2X1 NAND2X1_122 ( .A(asr2_en_bF_buf6), .B(asr2_cables_7__1_), .Y(_293_) );
OAI21X1 OAI21X1_122 ( .A(asr2_en_bF_buf6), .B(_292_), .C(_293_), .Y(_288__1_) );
INVX1 INVX1_139 ( .A(asr2_cables_8__2_), .Y(_294_) );
NAND2X1 NAND2X1_123 ( .A(asr2_en_bF_buf0), .B(asr2_cables_7__2_), .Y(_295_) );
OAI21X1 OAI21X1_123 ( .A(asr2_en_bF_buf4), .B(_294_), .C(_295_), .Y(_288__2_) );
INVX1 INVX1_140 ( .A(asr2_cables_8__3_), .Y(_296_) );
NAND2X1 NAND2X1_124 ( .A(asr2_en_bF_buf2), .B(asr2_cables_7__3_), .Y(_297_) );
OAI21X1 OAI21X1_124 ( .A(asr2_en_bF_buf2), .B(_296_), .C(_297_), .Y(_288__3_) );
INVX1 INVX1_141 ( .A(asr2_cables_8__4_), .Y(_298_) );
NAND2X1 NAND2X1_125 ( .A(asr2_en_bF_buf4), .B(asr2_cables_7__4_), .Y(_299_) );
OAI21X1 OAI21X1_125 ( .A(asr2_en_bF_buf4), .B(_298_), .C(_299_), .Y(_288__4_) );
INVX1 INVX1_142 ( .A(asr2_cables_8__5_), .Y(_300_) );
NAND2X1 NAND2X1_126 ( .A(asr2_en_bF_buf9), .B(asr2_cables_7__5_), .Y(_301_) );
OAI21X1 OAI21X1_126 ( .A(asr2_en_bF_buf9), .B(_300_), .C(_301_), .Y(_288__5_) );
INVX1 INVX1_143 ( .A(asr2_cables_8__6_), .Y(_302_) );
NAND2X1 NAND2X1_127 ( .A(asr2_en_bF_buf5), .B(asr2_cables_7__6_), .Y(_303_) );
OAI21X1 OAI21X1_127 ( .A(asr2_en_bF_buf4), .B(_302_), .C(_303_), .Y(_288__6_) );
INVX1 INVX1_144 ( .A(asr2_cables_8__7_), .Y(_304_) );
NAND2X1 NAND2X1_128 ( .A(asr2_en_bF_buf3), .B(asr2_cables_7__7_), .Y(_305_) );
OAI21X1 OAI21X1_128 ( .A(asr2_en_bF_buf6), .B(_304_), .C(_305_), .Y(_288__7_) );
INVX1 INVX1_145 ( .A(rst_bF_buf5), .Y(_289_) );
DFFSR DFFSR_121 ( .CLK(asr2_clk_bF_buf2), .D(_288__0_), .Q(asr2_cables_8__0_), .R(_289_), .S(vdd) );
DFFSR DFFSR_122 ( .CLK(asr2_clk_bF_buf7), .D(_288__1_), .Q(asr2_cables_8__1_), .R(_289_), .S(vdd) );
DFFSR DFFSR_123 ( .CLK(asr2_clk_bF_buf1), .D(_288__2_), .Q(asr2_cables_8__2_), .R(_289_), .S(vdd) );
DFFSR DFFSR_124 ( .CLK(asr2_clk_bF_buf7), .D(_288__3_), .Q(asr2_cables_8__3_), .R(_289_), .S(vdd) );
DFFSR DFFSR_125 ( .CLK(asr2_clk_bF_buf1), .D(_288__4_), .Q(asr2_cables_8__4_), .R(_289_), .S(vdd) );
DFFSR DFFSR_126 ( .CLK(asr2_clk_bF_buf4), .D(_288__5_), .Q(asr2_cables_8__5_), .R(_289_), .S(vdd) );
DFFSR DFFSR_127 ( .CLK(asr2_clk_bF_buf2), .D(_288__6_), .Q(asr2_cables_8__6_), .R(_289_), .S(vdd) );
DFFSR DFFSR_128 ( .CLK(asr2_clk_bF_buf7), .D(_288__7_), .Q(asr2_cables_8__7_), .R(_289_), .S(vdd) );
INVX1 INVX1_146 ( .A(retardo_asr_1_connect_wire_1__0_), .Y(_308_) );
NAND2X1 NAND2X1_129 ( .A(asr1_q_0_), .B(vdd), .Y(_309_) );
OAI21X1 OAI21X1_129 ( .A(vdd), .B(_308_), .C(_309_), .Y(_306__0_) );
INVX1 INVX1_147 ( .A(retardo_asr_1_connect_wire_1__1_), .Y(_310_) );
NAND2X1 NAND2X1_130 ( .A(vdd), .B(asr1_q_1_), .Y(_311_) );
OAI21X1 OAI21X1_130 ( .A(vdd), .B(_310_), .C(_311_), .Y(_306__1_) );
INVX1 INVX1_148 ( .A(retardo_asr_1_connect_wire_1__2_), .Y(_312_) );
NAND2X1 NAND2X1_131 ( .A(vdd), .B(asr1_q_2_), .Y(_313_) );
OAI21X1 OAI21X1_131 ( .A(vdd), .B(_312_), .C(_313_), .Y(_306__2_) );
INVX1 INVX1_149 ( .A(retardo_asr_1_connect_wire_1__3_), .Y(_314_) );
NAND2X1 NAND2X1_132 ( .A(vdd), .B(asr1_q_3_), .Y(_315_) );
OAI21X1 OAI21X1_132 ( .A(vdd), .B(_314_), .C(_315_), .Y(_306__3_) );
INVX1 INVX1_150 ( .A(retardo_asr_1_connect_wire_1__4_), .Y(_316_) );
NAND2X1 NAND2X1_133 ( .A(vdd), .B(asr1_q_4_), .Y(_317_) );
OAI21X1 OAI21X1_133 ( .A(vdd), .B(_316_), .C(_317_), .Y(_306__4_) );
INVX1 INVX1_151 ( .A(retardo_asr_1_connect_wire_1__5_), .Y(_318_) );
NAND2X1 NAND2X1_134 ( .A(vdd), .B(asr1_q_5_), .Y(_319_) );
OAI21X1 OAI21X1_134 ( .A(vdd), .B(_318_), .C(_319_), .Y(_306__5_) );
INVX1 INVX1_152 ( .A(retardo_asr_1_connect_wire_1__6_), .Y(_320_) );
NAND2X1 NAND2X1_135 ( .A(vdd), .B(asr1_q_6_), .Y(_321_) );
OAI21X1 OAI21X1_135 ( .A(vdd), .B(_320_), .C(_321_), .Y(_306__6_) );
INVX1 INVX1_153 ( .A(retardo_asr_1_connect_wire_1__7_), .Y(_322_) );
NAND2X1 NAND2X1_136 ( .A(vdd), .B(asr1_q_7_), .Y(_323_) );
OAI21X1 OAI21X1_136 ( .A(vdd), .B(_322_), .C(_323_), .Y(_306__7_) );
INVX1 INVX1_154 ( .A(rst_bF_buf2), .Y(_307_) );
DFFSR DFFSR_129 ( .CLK(clk_bF_buf3), .D(_306__0_), .Q(retardo_asr_1_connect_wire_1__0_), .R(_307_), .S(vdd) );
DFFSR DFFSR_130 ( .CLK(clk_bF_buf3), .D(_306__1_), .Q(retardo_asr_1_connect_wire_1__1_), .R(_307_), .S(vdd) );
DFFSR DFFSR_131 ( .CLK(clk_bF_buf3), .D(_306__2_), .Q(retardo_asr_1_connect_wire_1__2_), .R(_307_), .S(vdd) );
DFFSR DFFSR_132 ( .CLK(clk_bF_buf3), .D(_306__3_), .Q(retardo_asr_1_connect_wire_1__3_), .R(_307_), .S(vdd) );
DFFSR DFFSR_133 ( .CLK(clk_bF_buf5), .D(_306__4_), .Q(retardo_asr_1_connect_wire_1__4_), .R(_307_), .S(vdd) );
DFFSR DFFSR_134 ( .CLK(clk_bF_buf7), .D(_306__5_), .Q(retardo_asr_1_connect_wire_1__5_), .R(_307_), .S(vdd) );
DFFSR DFFSR_135 ( .CLK(clk_bF_buf5), .D(_306__6_), .Q(retardo_asr_1_connect_wire_1__6_), .R(_307_), .S(vdd) );
DFFSR DFFSR_136 ( .CLK(clk_bF_buf7), .D(_306__7_), .Q(retardo_asr_1_connect_wire_1__7_), .R(_307_), .S(vdd) );
INVX1 INVX1_155 ( .A(retardo_asr_2_connect_wire_1__0_), .Y(_326_) );
NAND2X1 NAND2X1_137 ( .A(asr2_q_0_), .B(vdd), .Y(_327_) );
OAI21X1 OAI21X1_137 ( .A(vdd), .B(_326_), .C(_327_), .Y(_324__0_) );
INVX1 INVX1_156 ( .A(retardo_asr_2_connect_wire_1__1_), .Y(_328_) );
NAND2X1 NAND2X1_138 ( .A(vdd), .B(asr2_q_1_), .Y(_329_) );
OAI21X1 OAI21X1_138 ( .A(vdd), .B(_328_), .C(_329_), .Y(_324__1_) );
INVX1 INVX1_157 ( .A(retardo_asr_2_connect_wire_1__2_), .Y(_330_) );
NAND2X1 NAND2X1_139 ( .A(vdd), .B(asr2_q_2_), .Y(_331_) );
OAI21X1 OAI21X1_139 ( .A(vdd), .B(_330_), .C(_331_), .Y(_324__2_) );
INVX1 INVX1_158 ( .A(retardo_asr_2_connect_wire_1__3_), .Y(_332_) );
NAND2X1 NAND2X1_140 ( .A(vdd), .B(asr2_q_3_), .Y(_333_) );
OAI21X1 OAI21X1_140 ( .A(vdd), .B(_332_), .C(_333_), .Y(_324__3_) );
INVX1 INVX1_159 ( .A(retardo_asr_2_connect_wire_1__4_), .Y(_334_) );
NAND2X1 NAND2X1_141 ( .A(vdd), .B(asr2_q_4_), .Y(_335_) );
OAI21X1 OAI21X1_141 ( .A(vdd), .B(_334_), .C(_335_), .Y(_324__4_) );
INVX1 INVX1_160 ( .A(retardo_asr_2_connect_wire_1__5_), .Y(_336_) );
NAND2X1 NAND2X1_142 ( .A(vdd), .B(asr2_q_5_), .Y(_337_) );
OAI21X1 OAI21X1_142 ( .A(vdd), .B(_336_), .C(_337_), .Y(_324__5_) );
INVX1 INVX1_161 ( .A(retardo_asr_2_connect_wire_1__6_), .Y(_338_) );
NAND2X1 NAND2X1_143 ( .A(vdd), .B(asr2_q_6_), .Y(_339_) );
OAI21X1 OAI21X1_143 ( .A(vdd), .B(_338_), .C(_339_), .Y(_324__6_) );
INVX1 INVX1_162 ( .A(retardo_asr_2_connect_wire_1__7_), .Y(_340_) );
NAND2X1 NAND2X1_144 ( .A(vdd), .B(asr2_q_7_), .Y(_341_) );
OAI21X1 OAI21X1_144 ( .A(vdd), .B(_340_), .C(_341_), .Y(_324__7_) );
INVX1 INVX1_163 ( .A(rst_bF_buf0), .Y(_325_) );
DFFSR DFFSR_137 ( .CLK(clk_bF_buf5), .D(_324__0_), .Q(retardo_asr_2_connect_wire_1__0_), .R(_325_), .S(vdd) );
DFFSR DFFSR_138 ( .CLK(clk_bF_buf3), .D(_324__1_), .Q(retardo_asr_2_connect_wire_1__1_), .R(_325_), .S(vdd) );
DFFSR DFFSR_139 ( .CLK(clk_bF_buf3), .D(_324__2_), .Q(retardo_asr_2_connect_wire_1__2_), .R(_325_), .S(vdd) );
DFFSR DFFSR_140 ( .CLK(clk_bF_buf7), .D(_324__3_), .Q(retardo_asr_2_connect_wire_1__3_), .R(_325_), .S(vdd) );
DFFSR DFFSR_141 ( .CLK(clk_bF_buf7), .D(_324__4_), .Q(retardo_asr_2_connect_wire_1__4_), .R(_325_), .S(vdd) );
DFFSR DFFSR_142 ( .CLK(clk_bF_buf7), .D(_324__5_), .Q(retardo_asr_2_connect_wire_1__5_), .R(_325_), .S(vdd) );
DFFSR DFFSR_143 ( .CLK(clk_bF_buf7), .D(_324__6_), .Q(retardo_asr_2_connect_wire_1__6_), .R(_325_), .S(vdd) );
DFFSR DFFSR_144 ( .CLK(clk_bF_buf7), .D(_324__7_), .Q(retardo_asr_2_connect_wire_1__7_), .R(_325_), .S(vdd) );
INVX1 INVX1_164 ( .A(retardo_clock_chico_connect_wire_1_), .Y(_344_) );
NAND2X1 NAND2X1_145 ( .A(enable_asr), .B(vdd), .Y(_345_) );
OAI21X1 OAI21X1_145 ( .A(vdd), .B(_344_), .C(_345_), .Y(_342_) );
INVX1 INVX1_165 ( .A(rst_bF_buf4), .Y(_343_) );
DFFSR DFFSR_145 ( .CLK(clk_bF_buf4), .D(_342_), .Q(retardo_clock_chico_connect_wire_1_), .R(_343_), .S(vdd) );
INVX1 INVX1_166 ( .A(retardo_clock_chico_connect_wire_2_), .Y(_348_) );
NAND2X1 NAND2X1_146 ( .A(retardo_clock_chico_connect_wire_1_), .B(vdd), .Y(_349_) );
OAI21X1 OAI21X1_146 ( .A(vdd), .B(_348_), .C(_349_), .Y(_346_) );
INVX1 INVX1_167 ( .A(rst_bF_buf4), .Y(_347_) );
DFFSR DFFSR_146 ( .CLK(clk_bF_buf4), .D(_346_), .Q(retardo_clock_chico_connect_wire_2_), .R(_347_), .S(vdd) );
INVX1 INVX1_168 ( .A(retardo_clock_chico_connect_wire_3_), .Y(_352_) );
NAND2X1 NAND2X1_147 ( .A(retardo_clock_chico_connect_wire_2_), .B(vdd), .Y(_353_) );
OAI21X1 OAI21X1_147 ( .A(vdd), .B(_352_), .C(_353_), .Y(_350_) );
INVX1 INVX1_169 ( .A(rst_bF_buf4), .Y(_351_) );
DFFSR DFFSR_147 ( .CLK(clk_bF_buf4), .D(_350_), .Q(retardo_clock_chico_connect_wire_3_), .R(_351_), .S(vdd) );
INVX1 INVX1_170 ( .A(retardo_clock_chico_connect_wire_4_), .Y(_356_) );
NAND2X1 NAND2X1_148 ( .A(retardo_clock_chico_connect_wire_3_), .B(vdd), .Y(_357_) );
OAI21X1 OAI21X1_148 ( .A(vdd), .B(_356_), .C(_357_), .Y(_354_) );
INVX1 INVX1_171 ( .A(rst_bF_buf5), .Y(_355_) );
DFFSR DFFSR_148 ( .CLK(clk_bF_buf4), .D(_354_), .Q(retardo_clock_chico_connect_wire_4_), .R(_355_), .S(vdd) );
INVX1 INVX1_172 ( .A(asr2_clk_bF_buf0), .Y(_360_) );
NAND2X1 NAND2X1_149 ( .A(retardo_clock_chico_connect_wire_4_), .B(vdd), .Y(_361_) );
OAI21X1 OAI21X1_149 ( .A(vdd), .B(_360_), .C(_361_), .Y(_358_) );
INVX1 INVX1_173 ( .A(rst_bF_buf5), .Y(_359_) );
DFFSR DFFSR_149 ( .CLK(clk_bF_buf4), .D(_358_), .Q(asr2_clk), .R(_359_), .S(vdd) );
INVX1 INVX1_174 ( .A(retardo_clock_mac_connect_wire_1_), .Y(_364_) );
NAND2X1 NAND2X1_150 ( .A(enable_asr), .B(vdd), .Y(_365_) );
OAI21X1 OAI21X1_150 ( .A(vdd), .B(_364_), .C(_365_), .Y(_362_) );
INVX1 INVX1_175 ( .A(rst_bF_buf1), .Y(_363_) );
DFFSR DFFSR_150 ( .CLK(clk_bF_buf7), .D(_362_), .Q(retardo_clock_mac_connect_wire_1_), .R(_363_), .S(vdd) );
INVX1 INVX1_176 ( .A(retardo_clock_mac_connect_wire_2_), .Y(_368_) );
NAND2X1 NAND2X1_151 ( .A(retardo_clock_mac_connect_wire_1_), .B(vdd), .Y(_369_) );
OAI21X1 OAI21X1_151 ( .A(vdd), .B(_368_), .C(_369_), .Y(_366_) );
INVX1 INVX1_177 ( .A(rst_bF_buf1), .Y(_367_) );
DFFSR DFFSR_151 ( .CLK(clk_bF_buf5), .D(_366_), .Q(retardo_clock_mac_connect_wire_2_), .R(_367_), .S(vdd) );
INVX1 INVX1_178 ( .A(retardo_clock_mac_connect_wire_3_), .Y(_372_) );
NAND2X1 NAND2X1_152 ( .A(retardo_clock_mac_connect_wire_2_), .B(vdd), .Y(_373_) );
OAI21X1 OAI21X1_152 ( .A(vdd), .B(_372_), .C(_373_), .Y(_370_) );
INVX1 INVX1_179 ( .A(rst_bF_buf5), .Y(_371_) );
DFFSR DFFSR_152 ( .CLK(clk_bF_buf5), .D(_370_), .Q(retardo_clock_mac_connect_wire_3_), .R(_371_), .S(vdd) );
INVX1 INVX1_180 ( .A(retardo_clock_mac_connect_wire_4_), .Y(_376_) );
NAND2X1 NAND2X1_153 ( .A(retardo_clock_mac_connect_wire_3_), .B(vdd), .Y(_377_) );
OAI21X1 OAI21X1_153 ( .A(vdd), .B(_376_), .C(_377_), .Y(_374_) );
INVX1 INVX1_181 ( .A(rst_bF_buf1), .Y(_375_) );
DFFSR DFFSR_153 ( .CLK(clk_bF_buf5), .D(_374_), .Q(retardo_clock_mac_connect_wire_4_), .R(_375_), .S(vdd) );
INVX1 INVX1_182 ( .A(retardo_clock_mac_connect_wire_5_), .Y(_380_) );
NAND2X1 NAND2X1_154 ( .A(retardo_clock_mac_connect_wire_4_), .B(vdd), .Y(_381_) );
OAI21X1 OAI21X1_154 ( .A(vdd), .B(_380_), .C(_381_), .Y(_378_) );
INVX1 INVX1_183 ( .A(rst_bF_buf1), .Y(_379_) );
DFFSR DFFSR_154 ( .CLK(clk_bF_buf5), .D(_378_), .Q(retardo_clock_mac_connect_wire_5_), .R(_379_), .S(vdd) );
INVX1 INVX1_184 ( .A(retardo_clock_mac_connect_wire_6_), .Y(_384_) );
NAND2X1 NAND2X1_155 ( .A(retardo_clock_mac_connect_wire_5_), .B(vdd), .Y(_385_) );
OAI21X1 OAI21X1_155 ( .A(vdd), .B(_384_), .C(_385_), .Y(_382_) );
INVX1 INVX1_185 ( .A(rst_bF_buf1), .Y(_383_) );
DFFSR DFFSR_155 ( .CLK(clk_bF_buf5), .D(_382_), .Q(retardo_clock_mac_connect_wire_6_), .R(_383_), .S(vdd) );
INVX1 INVX1_186 ( .A(retardo_clock_mac_connect_wire_7_), .Y(_388_) );
NAND2X1 NAND2X1_156 ( .A(retardo_clock_mac_connect_wire_6_), .B(vdd), .Y(_389_) );
OAI21X1 OAI21X1_156 ( .A(vdd), .B(_388_), .C(_389_), .Y(_386_) );
INVX1 INVX1_187 ( .A(rst_bF_buf4), .Y(_387_) );
DFFSR DFFSR_156 ( .CLK(clk_bF_buf4), .D(_386_), .Q(retardo_clock_mac_connect_wire_7_), .R(_387_), .S(vdd) );
INVX1 INVX1_188 ( .A(retardo_clock_mac_connect_wire_8_), .Y(_392_) );
NAND2X1 NAND2X1_157 ( .A(retardo_clock_mac_connect_wire_7_), .B(vdd), .Y(_393_) );
OAI21X1 OAI21X1_157 ( .A(vdd), .B(_392_), .C(_393_), .Y(_390_) );
INVX1 INVX1_189 ( .A(rst_bF_buf5), .Y(_391_) );
DFFSR DFFSR_157 ( .CLK(clk_bF_buf4), .D(_390_), .Q(retardo_clock_mac_connect_wire_8_), .R(_391_), .S(vdd) );
INVX1 INVX1_190 ( .A(retardo_clock_mac_connect_wire_9_), .Y(_396_) );
NAND2X1 NAND2X1_158 ( .A(retardo_clock_mac_connect_wire_8_), .B(vdd), .Y(_397_) );
OAI21X1 OAI21X1_158 ( .A(vdd), .B(_396_), .C(_397_), .Y(_394_) );
INVX1 INVX1_191 ( .A(rst_bF_buf3), .Y(_395_) );
DFFSR DFFSR_158 ( .CLK(clk_bF_buf2), .D(_394_), .Q(retardo_clock_mac_connect_wire_9_), .R(_395_), .S(vdd) );
INVX1 INVX1_192 ( .A(MAC_clr_bF_buf2), .Y(_400_) );
NAND2X1 NAND2X1_159 ( .A(retardo_clock_mac_connect_wire_9_), .B(vdd), .Y(_401_) );
OAI21X1 OAI21X1_159 ( .A(vdd), .B(_400_), .C(_401_), .Y(_398_) );
INVX1 INVX1_193 ( .A(rst_bF_buf3), .Y(_399_) );
DFFSR DFFSR_159 ( .CLK(clk_bF_buf1), .D(_398_), .Q(MAC_clr), .R(_399_), .S(vdd) );
INVX1 INVX1_194 ( .A(registro_salida_d_0_), .Y(_404_) );
NAND2X1 NAND2X1_160 ( .A(MAC_salida_correcta_0_), .B(MAC_clr_bF_buf1), .Y(_405_) );
OAI21X1 OAI21X1_160 ( .A(MAC_clr_bF_buf3), .B(_404_), .C(_405_), .Y(_402__0_) );
INVX1 INVX1_195 ( .A(registro_salida_d_1_), .Y(_406_) );
NAND2X1 NAND2X1_161 ( .A(MAC_clr_bF_buf2), .B(MAC_salida_correcta_1_), .Y(_407_) );
OAI21X1 OAI21X1_161 ( .A(MAC_clr_bF_buf2), .B(_406_), .C(_407_), .Y(_402__1_) );
INVX1 INVX1_196 ( .A(registro_salida_d_2_), .Y(_408_) );
NAND2X1 NAND2X1_162 ( .A(MAC_clr_bF_buf0), .B(MAC_salida_correcta_2_), .Y(_409_) );
OAI21X1 OAI21X1_162 ( .A(MAC_clr_bF_buf2), .B(_408_), .C(_409_), .Y(_402__2_) );
INVX1 INVX1_197 ( .A(registro_salida_d_3_), .Y(_410_) );
NAND2X1 NAND2X1_163 ( .A(MAC_clr_bF_buf3), .B(MAC_salida_correcta_3_), .Y(_411_) );
OAI21X1 OAI21X1_163 ( .A(MAC_clr_bF_buf3), .B(_410_), .C(_411_), .Y(_402__3_) );
INVX1 INVX1_198 ( .A(registro_salida_d_4_), .Y(_412_) );
NAND2X1 NAND2X1_164 ( .A(MAC_clr_bF_buf1), .B(MAC_salida_correcta_4_), .Y(_413_) );
OAI21X1 OAI21X1_164 ( .A(MAC_clr_bF_buf1), .B(_412_), .C(_413_), .Y(_402__4_) );
INVX1 INVX1_199 ( .A(registro_salida_d_5_), .Y(_414_) );
NAND2X1 NAND2X1_165 ( .A(MAC_clr_bF_buf0), .B(MAC_salida_correcta_5_), .Y(_415_) );
OAI21X1 OAI21X1_165 ( .A(MAC_clr_bF_buf2), .B(_414_), .C(_415_), .Y(_402__5_) );
INVX1 INVX1_200 ( .A(registro_salida_d_6_), .Y(_416_) );
NAND2X1 NAND2X1_166 ( .A(MAC_clr_bF_buf3), .B(MAC_salida_correcta_6_), .Y(_417_) );
OAI21X1 OAI21X1_166 ( .A(MAC_clr_bF_buf3), .B(_416_), .C(_417_), .Y(_402__6_) );
INVX1 INVX1_201 ( .A(registro_salida_d_7_), .Y(_418_) );
NAND2X1 NAND2X1_167 ( .A(MAC_clr_bF_buf0), .B(MAC_salida_correcta_7_), .Y(_419_) );
OAI21X1 OAI21X1_167 ( .A(MAC_clr_bF_buf0), .B(_418_), .C(_419_), .Y(_402__7_) );
INVX1 INVX1_202 ( .A(rst_bF_buf3), .Y(_403_) );
DFFSR DFFSR_160 ( .CLK(clk_bF_buf6), .D(_402__0_), .Q(registro_salida_d_0_), .R(_403_), .S(vdd) );
DFFSR DFFSR_161 ( .CLK(clk_bF_buf2), .D(_402__1_), .Q(registro_salida_d_1_), .R(_403_), .S(vdd) );
DFFSR DFFSR_162 ( .CLK(clk_bF_buf2), .D(_402__2_), .Q(registro_salida_d_2_), .R(_403_), .S(vdd) );
DFFSR DFFSR_163 ( .CLK(clk_bF_buf6), .D(_402__3_), .Q(registro_salida_d_3_), .R(_403_), .S(vdd) );
DFFSR DFFSR_164 ( .CLK(clk_bF_buf6), .D(_402__4_), .Q(registro_salida_d_4_), .R(_403_), .S(vdd) );
DFFSR DFFSR_165 ( .CLK(clk_bF_buf2), .D(_402__5_), .Q(registro_salida_d_5_), .R(_403_), .S(vdd) );
DFFSR DFFSR_166 ( .CLK(clk_bF_buf6), .D(_402__6_), .Q(registro_salida_d_6_), .R(_403_), .S(vdd) );
DFFSR DFFSR_167 ( .CLK(clk_bF_buf1), .D(_402__7_), .Q(registro_salida_d_7_), .R(_403_), .S(vdd) );
INVX1 INVX1_203 ( .A(MAC_ROM_0_bF_buf3_), .Y(_422_) );
NAND2X1 NAND2X1_168 ( .A(memoria_q_0_), .B(vdd), .Y(_423_) );
OAI21X1 OAI21X1_168 ( .A(vdd), .B(_422_), .C(_423_), .Y(_420__0_) );
INVX1 INVX1_204 ( .A(MAC_ROM_1_), .Y(_424_) );
NAND2X1 NAND2X1_169 ( .A(vdd), .B(memoria_q_1_), .Y(_425_) );
OAI21X1 OAI21X1_169 ( .A(vdd), .B(_424_), .C(_425_), .Y(_420__1_) );
INVX1 INVX1_205 ( .A(MAC_ROM_2_), .Y(_426_) );
NAND2X1 NAND2X1_170 ( .A(vdd), .B(memoria_q_2_), .Y(_427_) );
OAI21X1 OAI21X1_170 ( .A(vdd), .B(_426_), .C(_427_), .Y(_420__2_) );
INVX1 INVX1_206 ( .A(MAC_ROM_3_), .Y(_428_) );
NAND2X1 NAND2X1_171 ( .A(vdd), .B(memoria_q_3_), .Y(_429_) );
OAI21X1 OAI21X1_171 ( .A(vdd), .B(_428_), .C(_429_), .Y(_420__3_) );
INVX1 INVX1_207 ( .A(MAC_ROM_4_), .Y(_430_) );
NAND2X1 NAND2X1_172 ( .A(vdd), .B(gnd), .Y(_431_) );
OAI21X1 OAI21X1_172 ( .A(vdd), .B(_430_), .C(_431_), .Y(_420__4_) );
INVX1 INVX1_208 ( .A(MAC_ROM_5_), .Y(_432_) );
NAND2X1 NAND2X1_173 ( .A(vdd), .B(gnd), .Y(_433_) );
OAI21X1 OAI21X1_173 ( .A(vdd), .B(_432_), .C(_433_), .Y(_420__5_) );
INVX1 INVX1_209 ( .A(MAC_ROM_6_), .Y(_434_) );
NAND2X1 NAND2X1_174 ( .A(vdd), .B(gnd), .Y(_435_) );
OAI21X1 OAI21X1_174 ( .A(vdd), .B(_434_), .C(_435_), .Y(_420__6_) );
INVX1 INVX1_210 ( .A(MAC_ROM_7_), .Y(_436_) );
NAND2X1 NAND2X1_175 ( .A(vdd), .B(gnd), .Y(_437_) );
OAI21X1 OAI21X1_175 ( .A(vdd), .B(_436_), .C(_437_), .Y(_420__7_) );
INVX1 INVX1_211 ( .A(rst_bF_buf3), .Y(_421_) );
DFFSR DFFSR_168 ( .CLK(clk_bF_buf0), .D(_420__0_), .Q(MAC_ROM_0_), .R(_421_), .S(vdd) );
DFFSR DFFSR_169 ( .CLK(clk_bF_buf0), .D(_420__1_), .Q(MAC_ROM_1_), .R(_421_), .S(vdd) );
DFFSR DFFSR_170 ( .CLK(clk_bF_buf0), .D(_420__2_), .Q(MAC_ROM_2_), .R(_421_), .S(vdd) );
DFFSR DFFSR_171 ( .CLK(clk_bF_buf1), .D(_420__3_), .Q(MAC_ROM_3_), .R(_421_), .S(vdd) );
DFFSR DFFSR_172 ( .CLK(clk_bF_buf1), .D(_420__4_), .Q(MAC_ROM_4_), .R(_421_), .S(vdd) );
DFFSR DFFSR_173 ( .CLK(clk_bF_buf2), .D(_420__5_), .Q(MAC_ROM_5_), .R(_421_), .S(vdd) );
DFFSR DFFSR_174 ( .CLK(clk_bF_buf2), .D(_420__6_), .Q(MAC_ROM_6_), .R(_421_), .S(vdd) );
DFFSR DFFSR_175 ( .CLK(clk_bF_buf2), .D(_420__7_), .Q(MAC_ROM_7_), .R(_421_), .S(vdd) );
NAND2X1 NAND2X1_176 ( .A(MAC_ROM_0_bF_buf2_), .B(MAC_Adder_0_), .Y(_685_) );
INVX1 INVX1_212 ( .A(MAC_clr_bF_buf1), .Y(_696_) );
NAND2X1 NAND2X1_177 ( .A(MAC_salida_correcta_0_), .B(_696_), .Y(_707_) );
XOR2X1 XOR2X1_1 ( .A(_707_), .B(_685_), .Y(_438__0_) );
INVX1 INVX1_213 ( .A(MAC_ROM_0_bF_buf1_), .Y(_728_) );
INVX1 INVX1_214 ( .A(MAC_Adder_0_), .Y(_739_) );
INVX1 INVX1_215 ( .A(MAC_Adder_1_), .Y(_746_) );
INVX1 INVX1_216 ( .A(MAC_ROM_1_), .Y(_747_) );
OAI22X1 OAI22X1_1 ( .A(_728_), .B(_746_), .C(_739_), .D(_747_), .Y(_748_) );
NAND2X1 NAND2X1_178 ( .A(MAC_Adder_1_), .B(MAC_ROM_1_), .Y(_749_) );
OAI21X1 OAI21X1_176 ( .A(_685_), .B(_749_), .C(_748_), .Y(_750_) );
NAND3X1 NAND3X1_1 ( .A(MAC_ROM_0_bF_buf0_), .B(MAC_Adder_0_), .C(MAC_salida_correcta_0_), .Y(_751_) );
INVX1 INVX1_217 ( .A(_751_), .Y(_752_) );
INVX1 INVX1_218 ( .A(MAC_salida_correcta_1_), .Y(_753_) );
XOR2X1 XOR2X1_2 ( .A(_750_), .B(_753_), .Y(_754_) );
NAND2X1 NAND2X1_179 ( .A(_752_), .B(_754_), .Y(_755_) );
OR2X2 OR2X2_1 ( .A(_754_), .B(_752_), .Y(_756_) );
NAND3X1 NAND3X1_2 ( .A(_696_), .B(_755_), .C(_756_), .Y(_757_) );
OAI21X1 OAI21X1_177 ( .A(_696_), .B(_750_), .C(_757_), .Y(_438__1_) );
NAND2X1 NAND2X1_180 ( .A(MAC_Adder_0_), .B(MAC_ROM_2_), .Y(_758_) );
INVX1 INVX1_219 ( .A(_758_), .Y(_759_) );
AND2X2 AND2X2_2 ( .A(MAC_ROM_0_bF_buf3_), .B(MAC_Adder_2_), .Y(_760_) );
NAND3X1 NAND3X1_3 ( .A(MAC_Adder_1_), .B(MAC_ROM_1_), .C(_760_), .Y(_761_) );
AOI22X1 AOI22X1_1 ( .A(MAC_ROM_0_bF_buf2_), .B(MAC_Adder_2_), .C(MAC_Adder_1_), .D(MAC_ROM_1_), .Y(_762_) );
INVX1 INVX1_220 ( .A(_762_), .Y(_763_) );
NAND3X1 NAND3X1_4 ( .A(_763_), .B(_759_), .C(_761_), .Y(_764_) );
NAND2X1 NAND2X1_181 ( .A(MAC_ROM_0_bF_buf1_), .B(MAC_Adder_2_), .Y(_765_) );
NOR2X1 NOR2X1_3 ( .A(_749_), .B(_765_), .Y(_766_) );
OAI21X1 OAI21X1_178 ( .A(_762_), .B(_766_), .C(_758_), .Y(_767_) );
NAND2X1 NAND2X1_182 ( .A(_764_), .B(_767_), .Y(_768_) );
OAI21X1 OAI21X1_179 ( .A(_685_), .B(_749_), .C(_768_), .Y(_769_) );
NOR2X1 NOR2X1_4 ( .A(_685_), .B(_749_), .Y(_770_) );
NAND3X1 NAND3X1_5 ( .A(_770_), .B(_764_), .C(_767_), .Y(_771_) );
NAND2X1 NAND2X1_183 ( .A(_771_), .B(_769_), .Y(_772_) );
OAI21X1 OAI21X1_180 ( .A(_753_), .B(_750_), .C(_755_), .Y(_773_) );
INVX1 INVX1_221 ( .A(_773_), .Y(_774_) );
NAND3X1 NAND3X1_6 ( .A(MAC_salida_correcta_2_), .B(_771_), .C(_769_), .Y(_775_) );
INVX1 INVX1_222 ( .A(_775_), .Y(_776_) );
AOI21X1 AOI21X1_1 ( .A(_769_), .B(_771_), .C(MAC_salida_correcta_2_), .Y(_777_) );
NOR2X1 NOR2X1_5 ( .A(_777_), .B(_776_), .Y(_778_) );
AND2X2 AND2X2_3 ( .A(_778_), .B(_774_), .Y(_779_) );
NOR2X1 NOR2X1_6 ( .A(_774_), .B(_778_), .Y(_780_) );
OAI21X1 OAI21X1_181 ( .A(_780_), .B(_779_), .C(_696_), .Y(_781_) );
OAI21X1 OAI21X1_182 ( .A(_696_), .B(_772_), .C(_781_), .Y(_438__2_) );
OAI21X1 OAI21X1_183 ( .A(_777_), .B(_774_), .C(_775_), .Y(_782_) );
INVX1 INVX1_223 ( .A(_771_), .Y(_783_) );
NAND2X1 NAND2X1_184 ( .A(MAC_Adder_0_), .B(MAC_ROM_3_), .Y(_784_) );
INVX1 INVX1_224 ( .A(_784_), .Y(_785_) );
OAI21X1 OAI21X1_184 ( .A(_758_), .B(_762_), .C(_761_), .Y(_786_) );
NAND2X1 NAND2X1_185 ( .A(MAC_Adder_1_), .B(MAC_ROM_2_), .Y(_787_) );
INVX1 INVX1_225 ( .A(_787_), .Y(_788_) );
AND2X2 AND2X2_4 ( .A(MAC_ROM_1_), .B(MAC_Adder_2_), .Y(_789_) );
AND2X2 AND2X2_5 ( .A(MAC_ROM_0_bF_buf0_), .B(MAC_Adder_3_), .Y(_790_) );
NAND2X1 NAND2X1_186 ( .A(_789_), .B(_790_), .Y(_791_) );
INVX1 INVX1_226 ( .A(MAC_Adder_2_), .Y(_792_) );
NAND2X1 NAND2X1_187 ( .A(MAC_ROM_0_bF_buf3_), .B(MAC_Adder_3_), .Y(_793_) );
OAI21X1 OAI21X1_185 ( .A(_747_), .B(_792_), .C(_793_), .Y(_794_) );
NAND3X1 NAND3X1_7 ( .A(_794_), .B(_788_), .C(_791_), .Y(_795_) );
OAI21X1 OAI21X1_186 ( .A(_747_), .B(_792_), .C(_790_), .Y(_796_) );
INVX1 INVX1_227 ( .A(MAC_Adder_3_), .Y(_797_) );
OAI21X1 OAI21X1_187 ( .A(_728_), .B(_797_), .C(_789_), .Y(_798_) );
NAND3X1 NAND3X1_8 ( .A(_787_), .B(_796_), .C(_798_), .Y(_799_) );
NAND3X1 NAND3X1_9 ( .A(_795_), .B(_786_), .C(_799_), .Y(_800_) );
AOI21X1 AOI21X1_2 ( .A(_759_), .B(_763_), .C(_766_), .Y(_801_) );
NAND3X1 NAND3X1_10 ( .A(_787_), .B(_794_), .C(_791_), .Y(_802_) );
NAND3X1 NAND3X1_11 ( .A(_788_), .B(_796_), .C(_798_), .Y(_803_) );
NAND3X1 NAND3X1_12 ( .A(_802_), .B(_803_), .C(_801_), .Y(_439_) );
NAND3X1 NAND3X1_13 ( .A(_785_), .B(_800_), .C(_439_), .Y(_440_) );
NAND3X1 NAND3X1_14 ( .A(_795_), .B(_799_), .C(_801_), .Y(_441_) );
NAND3X1 NAND3X1_15 ( .A(_802_), .B(_786_), .C(_803_), .Y(_442_) );
NAND3X1 NAND3X1_16 ( .A(_784_), .B(_442_), .C(_441_), .Y(_443_) );
AOI21X1 AOI21X1_3 ( .A(_440_), .B(_443_), .C(_783_), .Y(_444_) );
INVX1 INVX1_228 ( .A(_444_), .Y(_445_) );
NAND3X1 NAND3X1_17 ( .A(_783_), .B(_440_), .C(_443_), .Y(_446_) );
NAND3X1 NAND3X1_18 ( .A(MAC_salida_correcta_3_), .B(_446_), .C(_445_), .Y(_447_) );
INVX1 INVX1_229 ( .A(MAC_salida_correcta_3_), .Y(_448_) );
INVX1 INVX1_230 ( .A(_446_), .Y(_449_) );
OAI21X1 OAI21X1_188 ( .A(_444_), .B(_449_), .C(_448_), .Y(_450_) );
NAND2X1 NAND2X1_188 ( .A(_447_), .B(_450_), .Y(_451_) );
XOR2X1 XOR2X1_3 ( .A(_451_), .B(_782_), .Y(_452_) );
NAND3X1 NAND3X1_19 ( .A(MAC_clr_bF_buf1), .B(_446_), .C(_445_), .Y(_453_) );
OAI21X1 OAI21X1_189 ( .A(MAC_clr_bF_buf3), .B(_452_), .C(_453_), .Y(_438__3_) );
NAND2X1 NAND2X1_189 ( .A(MAC_Adder_1_), .B(MAC_ROM_4_), .Y(_454_) );
INVX1 INVX1_231 ( .A(MAC_ROM_4_), .Y(_455_) );
NAND2X1 NAND2X1_190 ( .A(MAC_Adder_1_), .B(MAC_ROM_3_), .Y(_456_) );
OAI21X1 OAI21X1_190 ( .A(_739_), .B(_455_), .C(_456_), .Y(_457_) );
OAI21X1 OAI21X1_191 ( .A(_784_), .B(_454_), .C(_457_), .Y(_458_) );
AOI22X1 AOI22X1_2 ( .A(MAC_ROM_0_bF_buf2_), .B(MAC_Adder_3_), .C(MAC_ROM_1_), .D(MAC_Adder_2_), .Y(_459_) );
OAI21X1 OAI21X1_192 ( .A(_787_), .B(_459_), .C(_791_), .Y(_460_) );
NAND2X1 NAND2X1_191 ( .A(MAC_Adder_2_), .B(MAC_ROM_2_), .Y(_461_) );
INVX1 INVX1_232 ( .A(_461_), .Y(_462_) );
AND2X2 AND2X2_6 ( .A(MAC_ROM_1_), .B(MAC_Adder_4_), .Y(_463_) );
NAND2X1 NAND2X1_192 ( .A(_790_), .B(_463_), .Y(_464_) );
NAND2X1 NAND2X1_193 ( .A(MAC_ROM_1_), .B(MAC_Adder_3_), .Y(_465_) );
NAND2X1 NAND2X1_194 ( .A(MAC_ROM_0_bF_buf1_), .B(MAC_Adder_4_), .Y(_466_) );
NAND2X1 NAND2X1_195 ( .A(_465_), .B(_466_), .Y(_467_) );
NAND3X1 NAND3X1_20 ( .A(_462_), .B(_467_), .C(_464_), .Y(_468_) );
NAND3X1 NAND3X1_21 ( .A(MAC_ROM_0_bF_buf0_), .B(MAC_Adder_4_), .C(_465_), .Y(_469_) );
AND2X2 AND2X2_7 ( .A(MAC_ROM_1_), .B(MAC_Adder_3_), .Y(_470_) );
NAND2X1 NAND2X1_196 ( .A(_466_), .B(_470_), .Y(_471_) );
NAND3X1 NAND3X1_22 ( .A(_461_), .B(_469_), .C(_471_), .Y(_472_) );
NAND3X1 NAND3X1_23 ( .A(_460_), .B(_468_), .C(_472_), .Y(_473_) );
AOI22X1 AOI22X1_3 ( .A(_760_), .B(_470_), .C(_794_), .D(_788_), .Y(_474_) );
NAND3X1 NAND3X1_24 ( .A(_461_), .B(_467_), .C(_464_), .Y(_475_) );
NAND3X1 NAND3X1_25 ( .A(_462_), .B(_469_), .C(_471_), .Y(_476_) );
NAND3X1 NAND3X1_26 ( .A(_476_), .B(_475_), .C(_474_), .Y(_477_) );
NAND3X1 NAND3X1_27 ( .A(_458_), .B(_473_), .C(_477_), .Y(_478_) );
INVX1 INVX1_233 ( .A(_458_), .Y(_479_) );
AOI21X1 AOI21X1_4 ( .A(_475_), .B(_476_), .C(_474_), .Y(_480_) );
AOI21X1 AOI21X1_5 ( .A(_468_), .B(_472_), .C(_460_), .Y(_481_) );
OAI21X1 OAI21X1_193 ( .A(_481_), .B(_480_), .C(_479_), .Y(_482_) );
AOI22X1 AOI22X1_4 ( .A(_800_), .B(_440_), .C(_482_), .D(_478_), .Y(_483_) );
AOI21X1 AOI21X1_6 ( .A(_799_), .B(_795_), .C(_786_), .Y(_484_) );
OAI21X1 OAI21X1_194 ( .A(_784_), .B(_484_), .C(_800_), .Y(_485_) );
NAND3X1 NAND3X1_28 ( .A(_479_), .B(_473_), .C(_477_), .Y(_486_) );
OAI21X1 OAI21X1_195 ( .A(_481_), .B(_480_), .C(_458_), .Y(_487_) );
AOI21X1 AOI21X1_7 ( .A(_486_), .B(_487_), .C(_485_), .Y(_488_) );
OAI21X1 OAI21X1_196 ( .A(_483_), .B(_488_), .C(_446_), .Y(_489_) );
NAND3X1 NAND3X1_29 ( .A(_486_), .B(_487_), .C(_485_), .Y(_490_) );
AOI21X1 AOI21X1_8 ( .A(_802_), .B(_803_), .C(_801_), .Y(_491_) );
AOI21X1 AOI21X1_9 ( .A(_785_), .B(_439_), .C(_491_), .Y(_492_) );
NAND3X1 NAND3X1_30 ( .A(_478_), .B(_482_), .C(_492_), .Y(_493_) );
NAND3X1 NAND3X1_31 ( .A(_490_), .B(_493_), .C(_449_), .Y(_494_) );
NAND2X1 NAND2X1_197 ( .A(_489_), .B(_494_), .Y(_495_) );
INVX1 INVX1_234 ( .A(_777_), .Y(_496_) );
AOI21X1 AOI21X1_10 ( .A(_496_), .B(_773_), .C(_776_), .Y(_497_) );
AOI21X1 AOI21X1_11 ( .A(_445_), .B(_446_), .C(MAC_salida_correcta_3_), .Y(_498_) );
OAI21X1 OAI21X1_197 ( .A(_497_), .B(_498_), .C(_447_), .Y(_499_) );
NAND3X1 NAND3X1_32 ( .A(MAC_salida_correcta_4_), .B(_489_), .C(_494_), .Y(_500_) );
INVX1 INVX1_235 ( .A(MAC_salida_correcta_4_), .Y(_501_) );
NAND2X1 NAND2X1_198 ( .A(_501_), .B(_495_), .Y(_502_) );
NAND3X1 NAND3X1_33 ( .A(_500_), .B(_499_), .C(_502_), .Y(_503_) );
INVX1 INVX1_236 ( .A(_447_), .Y(_504_) );
AOI21X1 AOI21X1_12 ( .A(_450_), .B(_782_), .C(_504_), .Y(_505_) );
INVX1 INVX1_237 ( .A(_500_), .Y(_506_) );
AOI21X1 AOI21X1_13 ( .A(_494_), .B(_489_), .C(MAC_salida_correcta_4_), .Y(_507_) );
OAI21X1 OAI21X1_198 ( .A(_507_), .B(_506_), .C(_505_), .Y(_508_) );
NAND3X1 NAND3X1_34 ( .A(_696_), .B(_503_), .C(_508_), .Y(_509_) );
OAI21X1 OAI21X1_199 ( .A(_696_), .B(_495_), .C(_509_), .Y(_438__4_) );
NOR3X1 NOR3X1_1 ( .A(_446_), .B(_483_), .C(_488_), .Y(_510_) );
AND2X2 AND2X2_8 ( .A(MAC_Adder_1_), .B(MAC_ROM_4_), .Y(_511_) );
NAND2X1 NAND2X1_199 ( .A(_511_), .B(_785_), .Y(_512_) );
INVX1 INVX1_238 ( .A(_512_), .Y(_513_) );
OAI21X1 OAI21X1_200 ( .A(_458_), .B(_481_), .C(_473_), .Y(_514_) );
NAND2X1 NAND2X1_200 ( .A(MAC_Adder_0_), .B(MAC_ROM_5_), .Y(_515_) );
INVX1 INVX1_239 ( .A(_515_), .Y(_516_) );
AND2X2 AND2X2_9 ( .A(MAC_Adder_2_), .B(MAC_ROM_3_), .Y(_517_) );
NAND2X1 NAND2X1_201 ( .A(_511_), .B(_517_), .Y(_518_) );
INVX1 INVX1_240 ( .A(MAC_ROM_3_), .Y(_519_) );
OAI21X1 OAI21X1_201 ( .A(_792_), .B(_519_), .C(_454_), .Y(_520_) );
NAND3X1 NAND3X1_35 ( .A(_520_), .B(_516_), .C(_518_), .Y(_521_) );
OAI21X1 OAI21X1_202 ( .A(_746_), .B(_455_), .C(_517_), .Y(_522_) );
OAI21X1 OAI21X1_203 ( .A(_792_), .B(_519_), .C(_511_), .Y(_523_) );
NAND3X1 NAND3X1_36 ( .A(_515_), .B(_522_), .C(_523_), .Y(_524_) );
AOI22X1 AOI22X1_5 ( .A(_790_), .B(_463_), .C(_467_), .D(_462_), .Y(_525_) );
NAND2X1 NAND2X1_202 ( .A(MAC_ROM_2_), .B(MAC_Adder_3_), .Y(_526_) );
INVX1 INVX1_241 ( .A(_526_), .Y(_527_) );
AND2X2 AND2X2_10 ( .A(MAC_ROM_0_bF_buf3_), .B(MAC_Adder_5_), .Y(_528_) );
NAND2X1 NAND2X1_203 ( .A(_463_), .B(_528_), .Y(_529_) );
INVX1 INVX1_242 ( .A(MAC_Adder_5_), .Y(_530_) );
NAND2X1 NAND2X1_204 ( .A(MAC_ROM_1_), .B(MAC_Adder_4_), .Y(_531_) );
OAI21X1 OAI21X1_204 ( .A(_728_), .B(_530_), .C(_531_), .Y(_532_) );
NAND3X1 NAND3X1_37 ( .A(_527_), .B(_532_), .C(_529_), .Y(_533_) );
NAND3X1 NAND3X1_38 ( .A(MAC_ROM_0_bF_buf2_), .B(MAC_Adder_5_), .C(_531_), .Y(_534_) );
NAND2X1 NAND2X1_205 ( .A(MAC_ROM_0_bF_buf1_), .B(MAC_Adder_5_), .Y(_535_) );
NAND3X1 NAND3X1_39 ( .A(MAC_ROM_1_), .B(MAC_Adder_4_), .C(_535_), .Y(_536_) );
NAND3X1 NAND3X1_40 ( .A(_526_), .B(_534_), .C(_536_), .Y(_537_) );
NAND3X1 NAND3X1_41 ( .A(_525_), .B(_537_), .C(_533_), .Y(_538_) );
AOI22X1 AOI22X1_6 ( .A(MAC_ROM_0_bF_buf0_), .B(MAC_Adder_4_), .C(MAC_ROM_1_), .D(MAC_Adder_3_), .Y(_539_) );
OAI22X1 OAI22X1_2 ( .A(_793_), .B(_531_), .C(_461_), .D(_539_), .Y(_540_) );
NAND3X1 NAND3X1_42 ( .A(_526_), .B(_532_), .C(_529_), .Y(_541_) );
NAND3X1 NAND3X1_43 ( .A(_527_), .B(_534_), .C(_536_), .Y(_542_) );
NAND3X1 NAND3X1_44 ( .A(_540_), .B(_542_), .C(_541_), .Y(_543_) );
AOI22X1 AOI22X1_7 ( .A(_521_), .B(_524_), .C(_538_), .D(_543_), .Y(_544_) );
NAND3X1 NAND3X1_45 ( .A(_515_), .B(_520_), .C(_518_), .Y(_545_) );
NAND3X1 NAND3X1_46 ( .A(_516_), .B(_522_), .C(_523_), .Y(_546_) );
NAND3X1 NAND3X1_47 ( .A(_540_), .B(_537_), .C(_533_), .Y(_547_) );
NAND3X1 NAND3X1_48 ( .A(_525_), .B(_542_), .C(_541_), .Y(_548_) );
AOI22X1 AOI22X1_8 ( .A(_545_), .B(_546_), .C(_547_), .D(_548_), .Y(_549_) );
OAI21X1 OAI21X1_205 ( .A(_544_), .B(_549_), .C(_514_), .Y(_550_) );
AOI21X1 AOI21X1_14 ( .A(_479_), .B(_477_), .C(_480_), .Y(_551_) );
NAND2X1 NAND2X1_206 ( .A(_521_), .B(_524_), .Y(_552_) );
AOI21X1 AOI21X1_15 ( .A(_538_), .B(_543_), .C(_552_), .Y(_553_) );
NAND2X1 NAND2X1_207 ( .A(_545_), .B(_546_), .Y(_554_) );
AOI21X1 AOI21X1_16 ( .A(_547_), .B(_548_), .C(_554_), .Y(_555_) );
OAI21X1 OAI21X1_206 ( .A(_555_), .B(_553_), .C(_551_), .Y(_556_) );
NAND3X1 NAND3X1_49 ( .A(_513_), .B(_550_), .C(_556_), .Y(_557_) );
OAI21X1 OAI21X1_207 ( .A(_544_), .B(_549_), .C(_551_), .Y(_558_) );
OAI21X1 OAI21X1_208 ( .A(_555_), .B(_553_), .C(_514_), .Y(_559_) );
NAND3X1 NAND3X1_50 ( .A(_512_), .B(_558_), .C(_559_), .Y(_560_) );
NAND3X1 NAND3X1_51 ( .A(_483_), .B(_557_), .C(_560_), .Y(_561_) );
NAND3X1 NAND3X1_52 ( .A(_512_), .B(_550_), .C(_556_), .Y(_562_) );
NAND3X1 NAND3X1_53 ( .A(_513_), .B(_558_), .C(_559_), .Y(_563_) );
NAND3X1 NAND3X1_54 ( .A(_490_), .B(_562_), .C(_563_), .Y(_564_) );
NAND3X1 NAND3X1_55 ( .A(_510_), .B(_561_), .C(_564_), .Y(_565_) );
NAND3X1 NAND3X1_56 ( .A(_490_), .B(_557_), .C(_560_), .Y(_566_) );
NAND3X1 NAND3X1_57 ( .A(_483_), .B(_562_), .C(_563_), .Y(_567_) );
NAND3X1 NAND3X1_58 ( .A(_494_), .B(_566_), .C(_567_), .Y(_568_) );
NAND2X1 NAND2X1_208 ( .A(_565_), .B(_568_), .Y(_569_) );
OAI21X1 OAI21X1_209 ( .A(_507_), .B(_505_), .C(_500_), .Y(_570_) );
NAND3X1 NAND3X1_59 ( .A(MAC_salida_correcta_5_), .B(_565_), .C(_568_), .Y(_571_) );
INVX1 INVX1_243 ( .A(MAC_salida_correcta_5_), .Y(_572_) );
NAND2X1 NAND2X1_209 ( .A(_572_), .B(_569_), .Y(_573_) );
NAND3X1 NAND3X1_60 ( .A(_571_), .B(_573_), .C(_570_), .Y(_574_) );
AOI21X1 AOI21X1_17 ( .A(_499_), .B(_502_), .C(_506_), .Y(_575_) );
INVX1 INVX1_244 ( .A(_571_), .Y(_576_) );
AOI21X1 AOI21X1_18 ( .A(_565_), .B(_568_), .C(MAC_salida_correcta_5_), .Y(_577_) );
OAI21X1 OAI21X1_210 ( .A(_577_), .B(_576_), .C(_575_), .Y(_578_) );
NAND3X1 NAND3X1_61 ( .A(_696_), .B(_574_), .C(_578_), .Y(_579_) );
OAI21X1 OAI21X1_211 ( .A(_696_), .B(_569_), .C(_579_), .Y(_438__5_) );
AOI21X1 AOI21X1_19 ( .A(_566_), .B(_567_), .C(_494_), .Y(_580_) );
AOI21X1 AOI21X1_20 ( .A(_563_), .B(_562_), .C(_490_), .Y(_581_) );
NAND3X1 NAND3X1_62 ( .A(_547_), .B(_548_), .C(_554_), .Y(_582_) );
AOI21X1 AOI21X1_21 ( .A(_541_), .B(_542_), .C(_525_), .Y(_583_) );
AOI21X1 AOI21X1_22 ( .A(_533_), .B(_537_), .C(_540_), .Y(_584_) );
OAI21X1 OAI21X1_212 ( .A(_583_), .B(_584_), .C(_552_), .Y(_585_) );
AOI21X1 AOI21X1_23 ( .A(_585_), .B(_582_), .C(_514_), .Y(_586_) );
OAI21X1 OAI21X1_213 ( .A(_512_), .B(_586_), .C(_550_), .Y(_587_) );
AND2X2 AND2X2_11 ( .A(MAC_Adder_0_), .B(MAC_ROM_6_), .Y(_588_) );
NAND2X1 NAND2X1_210 ( .A(MAC_Adder_2_), .B(MAC_ROM_4_), .Y(_589_) );
OAI21X1 OAI21X1_214 ( .A(_456_), .B(_589_), .C(_521_), .Y(_590_) );
XNOR2X1 XNOR2X1_1 ( .A(_590_), .B(_588_), .Y(_591_) );
INVX1 INVX1_245 ( .A(_591_), .Y(_592_) );
OAI21X1 OAI21X1_215 ( .A(_552_), .B(_584_), .C(_547_), .Y(_593_) );
INVX1 INVX1_246 ( .A(MAC_ROM_5_), .Y(_594_) );
NOR2X1 NOR2X1_7 ( .A(_746_), .B(_594_), .Y(_595_) );
NAND2X1 NAND2X1_211 ( .A(MAC_Adder_3_), .B(MAC_ROM_3_), .Y(_596_) );
XOR2X1 XOR2X1_4 ( .A(_589_), .B(_596_), .Y(_597_) );
NAND2X1 NAND2X1_212 ( .A(_595_), .B(_597_), .Y(_598_) );
INVX1 INVX1_247 ( .A(_517_), .Y(_599_) );
NAND2X1 NAND2X1_213 ( .A(MAC_Adder_3_), .B(MAC_ROM_4_), .Y(_600_) );
OAI21X1 OAI21X1_216 ( .A(_797_), .B(_519_), .C(_589_), .Y(_601_) );
OAI21X1 OAI21X1_217 ( .A(_600_), .B(_599_), .C(_601_), .Y(_602_) );
OAI21X1 OAI21X1_218 ( .A(_746_), .B(_594_), .C(_602_), .Y(_603_) );
NOR2X1 NOR2X1_8 ( .A(_531_), .B(_535_), .Y(_604_) );
AOI21X1 AOI21X1_24 ( .A(_527_), .B(_532_), .C(_604_), .Y(_605_) );
NAND2X1 NAND2X1_214 ( .A(MAC_ROM_2_), .B(MAC_Adder_4_), .Y(_606_) );
INVX1 INVX1_248 ( .A(_606_), .Y(_607_) );
NAND3X1 NAND3X1_63 ( .A(MAC_ROM_1_), .B(MAC_Adder_6_), .C(_528_), .Y(_608_) );
AOI22X1 AOI22X1_9 ( .A(MAC_ROM_0_bF_buf3_), .B(MAC_Adder_6_), .C(MAC_ROM_1_), .D(MAC_Adder_5_), .Y(_609_) );
INVX1 INVX1_249 ( .A(_609_), .Y(_610_) );
NAND3X1 NAND3X1_64 ( .A(_610_), .B(_607_), .C(_608_), .Y(_611_) );
NAND2X1 NAND2X1_215 ( .A(MAC_ROM_1_), .B(MAC_Adder_6_), .Y(_612_) );
NOR2X1 NOR2X1_9 ( .A(_535_), .B(_612_), .Y(_613_) );
OAI21X1 OAI21X1_219 ( .A(_609_), .B(_613_), .C(_606_), .Y(_614_) );
NAND3X1 NAND3X1_65 ( .A(_611_), .B(_614_), .C(_605_), .Y(_615_) );
AND2X2 AND2X2_12 ( .A(_531_), .B(_535_), .Y(_616_) );
OAI21X1 OAI21X1_220 ( .A(_526_), .B(_616_), .C(_529_), .Y(_617_) );
NAND3X1 NAND3X1_66 ( .A(_606_), .B(_610_), .C(_608_), .Y(_618_) );
OAI21X1 OAI21X1_221 ( .A(_609_), .B(_613_), .C(_607_), .Y(_619_) );
NAND3X1 NAND3X1_67 ( .A(_618_), .B(_619_), .C(_617_), .Y(_620_) );
AOI22X1 AOI22X1_10 ( .A(_598_), .B(_603_), .C(_615_), .D(_620_), .Y(_621_) );
OAI21X1 OAI21X1_222 ( .A(_746_), .B(_594_), .C(_597_), .Y(_622_) );
NAND2X1 NAND2X1_216 ( .A(_595_), .B(_602_), .Y(_623_) );
NAND3X1 NAND3X1_68 ( .A(_611_), .B(_614_), .C(_617_), .Y(_624_) );
NAND3X1 NAND3X1_69 ( .A(_618_), .B(_619_), .C(_605_), .Y(_625_) );
AOI22X1 AOI22X1_11 ( .A(_622_), .B(_623_), .C(_625_), .D(_624_), .Y(_626_) );
OAI21X1 OAI21X1_223 ( .A(_621_), .B(_626_), .C(_593_), .Y(_627_) );
AOI21X1 AOI21X1_25 ( .A(_554_), .B(_548_), .C(_583_), .Y(_628_) );
AOI22X1 AOI22X1_12 ( .A(_622_), .B(_623_), .C(_615_), .D(_620_), .Y(_629_) );
AOI22X1 AOI22X1_13 ( .A(_598_), .B(_603_), .C(_625_), .D(_624_), .Y(_630_) );
OAI21X1 OAI21X1_224 ( .A(_629_), .B(_630_), .C(_628_), .Y(_631_) );
NAND3X1 NAND3X1_70 ( .A(_627_), .B(_592_), .C(_631_), .Y(_632_) );
OAI21X1 OAI21X1_225 ( .A(_621_), .B(_626_), .C(_628_), .Y(_633_) );
OAI21X1 OAI21X1_226 ( .A(_629_), .B(_630_), .C(_593_), .Y(_634_) );
NAND3X1 NAND3X1_71 ( .A(_591_), .B(_633_), .C(_634_), .Y(_635_) );
NAND3X1 NAND3X1_72 ( .A(_635_), .B(_632_), .C(_587_), .Y(_636_) );
NAND3X1 NAND3X1_73 ( .A(_547_), .B(_552_), .C(_548_), .Y(_637_) );
OAI21X1 OAI21X1_227 ( .A(_583_), .B(_584_), .C(_554_), .Y(_638_) );
AOI21X1 AOI21X1_26 ( .A(_638_), .B(_637_), .C(_551_), .Y(_639_) );
AOI21X1 AOI21X1_27 ( .A(_513_), .B(_556_), .C(_639_), .Y(_640_) );
NAND3X1 NAND3X1_74 ( .A(_591_), .B(_627_), .C(_631_), .Y(_641_) );
NAND3X1 NAND3X1_75 ( .A(_633_), .B(_592_), .C(_634_), .Y(_642_) );
NAND3X1 NAND3X1_76 ( .A(_641_), .B(_642_), .C(_640_), .Y(_643_) );
NAND3X1 NAND3X1_77 ( .A(_581_), .B(_643_), .C(_636_), .Y(_644_) );
NAND3X1 NAND3X1_78 ( .A(_635_), .B(_632_), .C(_640_), .Y(_645_) );
NAND3X1 NAND3X1_79 ( .A(_641_), .B(_642_), .C(_587_), .Y(_646_) );
NAND3X1 NAND3X1_80 ( .A(_561_), .B(_645_), .C(_646_), .Y(_647_) );
NAND3X1 NAND3X1_81 ( .A(_580_), .B(_644_), .C(_647_), .Y(_648_) );
NAND3X1 NAND3X1_82 ( .A(_561_), .B(_643_), .C(_636_), .Y(_649_) );
NAND3X1 NAND3X1_83 ( .A(_581_), .B(_645_), .C(_646_), .Y(_650_) );
NAND3X1 NAND3X1_84 ( .A(_565_), .B(_649_), .C(_650_), .Y(_651_) );
NAND2X1 NAND2X1_217 ( .A(_648_), .B(_651_), .Y(_652_) );
OAI21X1 OAI21X1_228 ( .A(_577_), .B(_575_), .C(_571_), .Y(_653_) );
NAND3X1 NAND3X1_85 ( .A(MAC_salida_correcta_6_), .B(_648_), .C(_651_), .Y(_654_) );
INVX1 INVX1_250 ( .A(MAC_salida_correcta_6_), .Y(_655_) );
NAND3X1 NAND3X1_86 ( .A(_565_), .B(_644_), .C(_647_), .Y(_656_) );
NAND3X1 NAND3X1_87 ( .A(_580_), .B(_649_), .C(_650_), .Y(_657_) );
NAND3X1 NAND3X1_88 ( .A(_655_), .B(_656_), .C(_657_), .Y(_658_) );
AOI21X1 AOI21X1_28 ( .A(_654_), .B(_658_), .C(_653_), .Y(_659_) );
AOI21X1 AOI21X1_29 ( .A(_570_), .B(_573_), .C(_576_), .Y(_660_) );
NAND2X1 NAND2X1_218 ( .A(_654_), .B(_658_), .Y(_661_) );
OAI21X1 OAI21X1_229 ( .A(_660_), .B(_661_), .C(_696_), .Y(_662_) );
OAI22X1 OAI22X1_3 ( .A(_696_), .B(_652_), .C(_659_), .D(_662_), .Y(_438__6_) );
NAND2X1 NAND2X1_219 ( .A(_644_), .B(_648_), .Y(_663_) );
INVX1 INVX1_251 ( .A(_663_), .Y(_664_) );
INVX1 INVX1_252 ( .A(_636_), .Y(_665_) );
NAND2X1 NAND2X1_220 ( .A(_588_), .B(_590_), .Y(_666_) );
INVX1 INVX1_253 ( .A(_666_), .Y(_667_) );
NAND2X1 NAND2X1_221 ( .A(_627_), .B(_632_), .Y(_668_) );
OAI21X1 OAI21X1_230 ( .A(_599_), .B(_600_), .C(_598_), .Y(_669_) );
NAND2X1 NAND2X1_222 ( .A(MAC_Adder_0_), .B(MAC_ROM_7_), .Y(_670_) );
NAND2X1 NAND2X1_223 ( .A(MAC_Adder_1_), .B(MAC_ROM_6_), .Y(_671_) );
XOR2X1 XOR2X1_5 ( .A(_670_), .B(_671_), .Y(_672_) );
XOR2X1 XOR2X1_6 ( .A(_669_), .B(_672_), .Y(_673_) );
INVX1 INVX1_254 ( .A(_673_), .Y(_674_) );
INVX1 INVX1_255 ( .A(_624_), .Y(_675_) );
OR2X2 OR2X2_2 ( .A(_629_), .B(_675_), .Y(_676_) );
INVX1 INVX1_256 ( .A(MAC_ROM_2_), .Y(_677_) );
NOR2X1 NOR2X1_10 ( .A(_677_), .B(_530_), .Y(_678_) );
NAND2X1 NAND2X1_224 ( .A(MAC_ROM_0_bF_buf2_), .B(MAC_Adder_7_), .Y(_679_) );
XNOR2X1 XNOR2X1_2 ( .A(_612_), .B(_679_), .Y(_680_) );
INVX1 INVX1_257 ( .A(_680_), .Y(_681_) );
NAND2X1 NAND2X1_225 ( .A(_678_), .B(_681_), .Y(_682_) );
OAI21X1 OAI21X1_231 ( .A(_677_), .B(_530_), .C(_680_), .Y(_683_) );
OAI21X1 OAI21X1_232 ( .A(_606_), .B(_609_), .C(_608_), .Y(_684_) );
INVX1 INVX1_258 ( .A(_684_), .Y(_686_) );
NAND3X1 NAND3X1_89 ( .A(_683_), .B(_686_), .C(_682_), .Y(_687_) );
NAND2X1 NAND2X1_226 ( .A(_678_), .B(_680_), .Y(_688_) );
OAI21X1 OAI21X1_233 ( .A(_677_), .B(_530_), .C(_681_), .Y(_689_) );
NAND3X1 NAND3X1_90 ( .A(_684_), .B(_688_), .C(_689_), .Y(_690_) );
NAND2X1 NAND2X1_227 ( .A(MAC_ROM_3_), .B(MAC_Adder_4_), .Y(_691_) );
XNOR2X1 XNOR2X1_3 ( .A(_600_), .B(_691_), .Y(_692_) );
NAND2X1 NAND2X1_228 ( .A(MAC_Adder_2_), .B(MAC_ROM_5_), .Y(_693_) );
XOR2X1 XOR2X1_7 ( .A(_692_), .B(_693_), .Y(_694_) );
INVX1 INVX1_259 ( .A(_694_), .Y(_695_) );
NAND3X1 NAND3X1_91 ( .A(_687_), .B(_690_), .C(_695_), .Y(_697_) );
NAND3X1 NAND3X1_92 ( .A(_683_), .B(_684_), .C(_682_), .Y(_698_) );
NAND3X1 NAND3X1_93 ( .A(_686_), .B(_688_), .C(_689_), .Y(_699_) );
NAND3X1 NAND3X1_94 ( .A(_694_), .B(_698_), .C(_699_), .Y(_700_) );
NAND3X1 NAND3X1_95 ( .A(_700_), .B(_697_), .C(_676_), .Y(_701_) );
NOR2X1 NOR2X1_11 ( .A(_675_), .B(_629_), .Y(_702_) );
NAND3X1 NAND3X1_96 ( .A(_698_), .B(_699_), .C(_695_), .Y(_703_) );
NAND3X1 NAND3X1_97 ( .A(_694_), .B(_687_), .C(_690_), .Y(_704_) );
NAND3X1 NAND3X1_98 ( .A(_702_), .B(_704_), .C(_703_), .Y(_705_) );
AOI21X1 AOI21X1_30 ( .A(_701_), .B(_705_), .C(_674_), .Y(_706_) );
NAND3X1 NAND3X1_99 ( .A(_702_), .B(_700_), .C(_697_), .Y(_708_) );
NAND3X1 NAND3X1_100 ( .A(_704_), .B(_703_), .C(_676_), .Y(_709_) );
AOI21X1 AOI21X1_31 ( .A(_709_), .B(_708_), .C(_673_), .Y(_710_) );
OAI21X1 OAI21X1_234 ( .A(_706_), .B(_710_), .C(_668_), .Y(_711_) );
INVX1 INVX1_260 ( .A(_668_), .Y(_712_) );
NAND3X1 NAND3X1_101 ( .A(_673_), .B(_708_), .C(_709_), .Y(_713_) );
NAND3X1 NAND3X1_102 ( .A(_674_), .B(_705_), .C(_701_), .Y(_714_) );
NAND3X1 NAND3X1_103 ( .A(_713_), .B(_714_), .C(_712_), .Y(_715_) );
AOI21X1 AOI21X1_32 ( .A(_715_), .B(_711_), .C(_667_), .Y(_716_) );
NAND3X1 NAND3X1_104 ( .A(_668_), .B(_713_), .C(_714_), .Y(_717_) );
OAI21X1 OAI21X1_235 ( .A(_706_), .B(_710_), .C(_712_), .Y(_718_) );
AOI21X1 AOI21X1_33 ( .A(_718_), .B(_717_), .C(_666_), .Y(_719_) );
OAI21X1 OAI21X1_236 ( .A(_719_), .B(_716_), .C(_665_), .Y(_720_) );
NAND3X1 NAND3X1_105 ( .A(_666_), .B(_717_), .C(_718_), .Y(_721_) );
NAND3X1 NAND3X1_106 ( .A(_667_), .B(_711_), .C(_715_), .Y(_722_) );
NAND3X1 NAND3X1_107 ( .A(_636_), .B(_721_), .C(_722_), .Y(_723_) );
NAND3X1 NAND3X1_108 ( .A(_664_), .B(_723_), .C(_720_), .Y(_724_) );
NAND2X1 NAND2X1_229 ( .A(_711_), .B(_715_), .Y(_725_) );
XOR2X1 XOR2X1_8 ( .A(_636_), .B(_667_), .Y(_726_) );
OR2X2 OR2X2_3 ( .A(_725_), .B(_726_), .Y(_727_) );
NAND2X1 NAND2X1_230 ( .A(_726_), .B(_725_), .Y(_729_) );
NAND3X1 NAND3X1_109 ( .A(_663_), .B(_729_), .C(_727_), .Y(_730_) );
NAND2X1 NAND2X1_231 ( .A(_730_), .B(_724_), .Y(_731_) );
INVX1 INVX1_261 ( .A(MAC_salida_correcta_7_), .Y(_732_) );
AOI21X1 AOI21X1_34 ( .A(_656_), .B(_657_), .C(_655_), .Y(_733_) );
AOI21X1 AOI21X1_35 ( .A(_653_), .B(_658_), .C(_733_), .Y(_734_) );
NAND2X1 NAND2X1_232 ( .A(_732_), .B(_734_), .Y(_735_) );
AOI21X1 AOI21X1_36 ( .A(_648_), .B(_651_), .C(MAC_salida_correcta_6_), .Y(_736_) );
OAI21X1 OAI21X1_237 ( .A(_736_), .B(_660_), .C(_654_), .Y(_737_) );
AOI21X1 AOI21X1_37 ( .A(_737_), .B(MAC_salida_correcta_7_), .C(MAC_clr_bF_buf0), .Y(_738_) );
NAND3X1 NAND3X1_110 ( .A(_731_), .B(_735_), .C(_738_), .Y(_740_) );
AOI21X1 AOI21X1_38 ( .A(_727_), .B(_729_), .C(_664_), .Y(_741_) );
AOI21X1 AOI21X1_39 ( .A(_720_), .B(_723_), .C(_663_), .Y(_742_) );
AND2X2 AND2X2_13 ( .A(_734_), .B(_732_), .Y(_743_) );
OAI21X1 OAI21X1_238 ( .A(_732_), .B(_734_), .C(_696_), .Y(_744_) );
OAI22X1 OAI22X1_4 ( .A(_741_), .B(_742_), .C(_744_), .D(_743_), .Y(_745_) );
NAND2X1 NAND2X1_233 ( .A(_745_), .B(_740_), .Y(_438__7_) );
DFFPOSX1 DFFPOSX1_2 ( .CLK(clk_bF_buf6), .D(_438__0_), .Q(MAC_salida_correcta_0_) );
DFFPOSX1 DFFPOSX1_3 ( .CLK(clk_bF_buf1), .D(_438__1_), .Q(MAC_salida_correcta_1_) );
DFFPOSX1 DFFPOSX1_4 ( .CLK(clk_bF_buf6), .D(_438__2_), .Q(MAC_salida_correcta_2_) );
DFFPOSX1 DFFPOSX1_5 ( .CLK(clk_bF_buf6), .D(_438__3_), .Q(MAC_salida_correcta_3_) );
DFFPOSX1 DFFPOSX1_6 ( .CLK(clk_bF_buf6), .D(_438__4_), .Q(MAC_salida_correcta_4_) );
DFFPOSX1 DFFPOSX1_7 ( .CLK(clk_bF_buf1), .D(_438__5_), .Q(MAC_salida_correcta_5_) );
DFFPOSX1 DFFPOSX1_8 ( .CLK(clk_bF_buf1), .D(_438__6_), .Q(MAC_salida_correcta_6_) );
DFFPOSX1 DFFPOSX1_9 ( .CLK(clk_bF_buf1), .D(_438__7_), .Q(MAC_salida_correcta_7_) );
INVX1 INVX1_262 ( .A(asr1_cables_1__0_), .Y(_911_) );
INVX1 INVX1_263 ( .A(asr1_cables_2__0_), .Y(_912_) );
INVX1 INVX1_264 ( .A(up_counter_contador_1_), .Y(_913_) );
INVX1 INVX1_265 ( .A(up_counter_contador_2_), .Y(_914_) );
NAND3X1 NAND3X1_111 ( .A(up_counter_contador_0_), .B(_913_), .C(_914_), .Y(_915_) );
INVX1 INVX1_266 ( .A(up_counter_contador_0_), .Y(_916_) );
NAND3X1 NAND3X1_112 ( .A(_916_), .B(_913_), .C(_914_), .Y(_917_) );
OAI22X1 OAI22X1_5 ( .A(_912_), .B(_915_), .C(_911_), .D(_917_), .Y(_918_) );
INVX1 INVX1_267 ( .A(asr1_cables_7__0_), .Y(_919_) );
INVX1 INVX1_268 ( .A(asr1_cables_3__0_), .Y(_920_) );
NAND3X1 NAND3X1_113 ( .A(up_counter_contador_1_), .B(_916_), .C(_914_), .Y(_921_) );
NAND3X1 NAND3X1_114 ( .A(up_counter_contador_1_), .B(up_counter_contador_2_), .C(_916_), .Y(_922_) );
OAI22X1 OAI22X1_6 ( .A(_919_), .B(_922_), .C(_920_), .D(_921_), .Y(_923_) );
NOR2X1 NOR2X1_12 ( .A(_923_), .B(_918_), .Y(_924_) );
INVX1 INVX1_269 ( .A(asr1_cables_5__0_), .Y(_925_) );
INVX1 INVX1_270 ( .A(asr1_cables_4_), .Y(_926_) );
NAND3X1 NAND3X1_115 ( .A(up_counter_contador_0_), .B(up_counter_contador_1_), .C(_914_), .Y(_804_) );
NAND3X1 NAND3X1_116 ( .A(up_counter_contador_2_), .B(_916_), .C(_913_), .Y(_805_) );
OAI22X1 OAI22X1_7 ( .A(_926_), .B(_804_), .C(_925_), .D(_805_), .Y(_806_) );
INVX1 INVX1_271 ( .A(asr1_cables_8__0_), .Y(_807_) );
INVX1 INVX1_272 ( .A(asr1_cables_6__0_), .Y(_808_) );
NAND3X1 NAND3X1_117 ( .A(up_counter_contador_0_), .B(up_counter_contador_1_), .C(up_counter_contador_2_), .Y(_809_) );
NAND3X1 NAND3X1_118 ( .A(up_counter_contador_0_), .B(up_counter_contador_2_), .C(_913_), .Y(_810_) );
OAI22X1 OAI22X1_8 ( .A(_807_), .B(_809_), .C(_808_), .D(_810_), .Y(_811_) );
NOR2X1 NOR2X1_13 ( .A(_811_), .B(_806_), .Y(_812_) );
NAND2X1 NAND2X1_234 ( .A(_812_), .B(_924_), .Y(asr1_q_0_) );
INVX1 INVX1_273 ( .A(asr1_cables_1__1_), .Y(_813_) );
INVX1 INVX1_274 ( .A(asr1_cables_2__1_), .Y(_814_) );
OAI22X1 OAI22X1_9 ( .A(_814_), .B(_915_), .C(_813_), .D(_917_), .Y(_815_) );
INVX1 INVX1_275 ( .A(asr1_cables_6__1_), .Y(_816_) );
INVX1 INVX1_276 ( .A(asr1_cables_3__1_), .Y(_817_) );
OAI22X1 OAI22X1_10 ( .A(_816_), .B(_810_), .C(_817_), .D(_921_), .Y(_818_) );
NOR2X1 NOR2X1_14 ( .A(_818_), .B(_815_), .Y(_819_) );
INVX1 INVX1_277 ( .A(asr1_cables_7__1_), .Y(_820_) );
INVX1 INVX1_278 ( .A(asr1_cables_8__1_), .Y(_821_) );
OAI22X1 OAI22X1_11 ( .A(_821_), .B(_809_), .C(_820_), .D(_922_), .Y(_822_) );
INVX1 INVX1_279 ( .A(asr1_cables_5__1_), .Y(_823_) );
INVX1 INVX1_280 ( .A(_76_), .Y(_824_) );
OAI22X1 OAI22X1_12 ( .A(_824_), .B(_804_), .C(_823_), .D(_805_), .Y(_825_) );
NOR2X1 NOR2X1_15 ( .A(_822_), .B(_825_), .Y(_826_) );
NAND2X1 NAND2X1_235 ( .A(_826_), .B(_819_), .Y(asr1_q_1_) );
INVX1 INVX1_281 ( .A(asr1_cables_1__2_), .Y(_827_) );
INVX1 INVX1_282 ( .A(asr1_cables_2__2_), .Y(_828_) );
OAI22X1 OAI22X1_13 ( .A(_828_), .B(_915_), .C(_827_), .D(_917_), .Y(_829_) );
INVX1 INVX1_283 ( .A(asr1_cables_7__2_), .Y(_830_) );
INVX1 INVX1_284 ( .A(asr1_cables_3__2_), .Y(_831_) );
OAI22X1 OAI22X1_14 ( .A(_830_), .B(_922_), .C(_831_), .D(_921_), .Y(_832_) );
NOR2X1 NOR2X1_16 ( .A(_832_), .B(_829_), .Y(_833_) );
INVX1 INVX1_285 ( .A(asr1_cables_5__2_), .Y(_834_) );
INVX1 INVX1_286 ( .A(_82_), .Y(_835_) );
OAI22X1 OAI22X1_15 ( .A(_835_), .B(_804_), .C(_834_), .D(_805_), .Y(_836_) );
INVX1 INVX1_287 ( .A(asr1_cables_8__2_), .Y(_837_) );
INVX1 INVX1_288 ( .A(asr1_cables_6__2_), .Y(_838_) );
OAI22X1 OAI22X1_16 ( .A(_837_), .B(_809_), .C(_838_), .D(_810_), .Y(_839_) );
NOR2X1 NOR2X1_17 ( .A(_839_), .B(_836_), .Y(_840_) );
NAND2X1 NAND2X1_236 ( .A(_840_), .B(_833_), .Y(asr1_q_2_) );
INVX1 INVX1_289 ( .A(asr1_cables_3__3_), .Y(_841_) );
INVX1 INVX1_290 ( .A(asr1_cables_2__3_), .Y(_842_) );
OAI22X1 OAI22X1_17 ( .A(_841_), .B(_921_), .C(_842_), .D(_915_), .Y(_843_) );
INVX1 INVX1_291 ( .A(asr1_cables_7__3_), .Y(_844_) );
INVX1 INVX1_292 ( .A(asr1_cables_6__3_), .Y(_845_) );
OAI22X1 OAI22X1_18 ( .A(_844_), .B(_922_), .C(_845_), .D(_810_), .Y(_846_) );
NOR2X1 NOR2X1_18 ( .A(_846_), .B(_843_), .Y(_847_) );
INVX1 INVX1_293 ( .A(asr1_cables_5__3_), .Y(_848_) );
INVX1 INVX1_294 ( .A(_77_), .Y(_849_) );
OAI22X1 OAI22X1_19 ( .A(_849_), .B(_804_), .C(_848_), .D(_805_), .Y(_850_) );
INVX1 INVX1_295 ( .A(asr1_cables_8__3_), .Y(_851_) );
INVX1 INVX1_296 ( .A(asr1_cables_1__3_), .Y(_852_) );
OAI22X1 OAI22X1_20 ( .A(_851_), .B(_809_), .C(_852_), .D(_917_), .Y(_853_) );
NOR2X1 NOR2X1_19 ( .A(_850_), .B(_853_), .Y(_854_) );
NAND2X1 NAND2X1_237 ( .A(_847_), .B(_854_), .Y(asr1_q_3_) );
INVX1 INVX1_297 ( .A(asr1_cables_1__4_), .Y(_855_) );
INVX1 INVX1_298 ( .A(asr1_cables_2__4_), .Y(_856_) );
OAI22X1 OAI22X1_21 ( .A(_856_), .B(_915_), .C(_855_), .D(_917_), .Y(_857_) );
INVX1 INVX1_299 ( .A(asr1_cables_7__4_), .Y(_858_) );
INVX1 INVX1_300 ( .A(asr1_cables_3__4_), .Y(_859_) );
OAI22X1 OAI22X1_22 ( .A(_858_), .B(_922_), .C(_859_), .D(_921_), .Y(_860_) );
NOR2X1 NOR2X1_20 ( .A(_860_), .B(_857_), .Y(_861_) );
INVX1 INVX1_301 ( .A(asr1_cables_5__4_), .Y(_862_) );
INVX1 INVX1_302 ( .A(_78_), .Y(_863_) );
OAI22X1 OAI22X1_23 ( .A(_863_), .B(_804_), .C(_862_), .D(_805_), .Y(_864_) );
INVX1 INVX1_303 ( .A(asr1_cables_8__4_), .Y(_865_) );
INVX1 INVX1_304 ( .A(asr1_cables_6__4_), .Y(_866_) );
OAI22X1 OAI22X1_24 ( .A(_865_), .B(_809_), .C(_866_), .D(_810_), .Y(_867_) );
NOR2X1 NOR2X1_21 ( .A(_867_), .B(_864_), .Y(_868_) );
NAND2X1 NAND2X1_238 ( .A(_868_), .B(_861_), .Y(asr1_q_4_) );
INVX1 INVX1_305 ( .A(asr1_cables_3__5_), .Y(_869_) );
INVX1 INVX1_306 ( .A(asr1_cables_2__5_), .Y(_870_) );
OAI22X1 OAI22X1_25 ( .A(_869_), .B(_921_), .C(_870_), .D(_915_), .Y(_871_) );
INVX1 INVX1_307 ( .A(asr1_cables_7__5_), .Y(_872_) );
INVX1 INVX1_308 ( .A(asr1_cables_6__5_), .Y(_873_) );
OAI22X1 OAI22X1_26 ( .A(_872_), .B(_922_), .C(_873_), .D(_810_), .Y(_874_) );
NOR2X1 NOR2X1_22 ( .A(_874_), .B(_871_), .Y(_875_) );
INVX1 INVX1_309 ( .A(asr1_cables_5__5_), .Y(_876_) );
INVX1 INVX1_310 ( .A(_79_), .Y(_877_) );
OAI22X1 OAI22X1_27 ( .A(_877_), .B(_804_), .C(_876_), .D(_805_), .Y(_878_) );
INVX1 INVX1_311 ( .A(asr1_cables_8__5_), .Y(_879_) );
INVX1 INVX1_312 ( .A(asr1_cables_1__5_), .Y(_880_) );
OAI22X1 OAI22X1_28 ( .A(_879_), .B(_809_), .C(_880_), .D(_917_), .Y(_881_) );
NOR2X1 NOR2X1_23 ( .A(_878_), .B(_881_), .Y(_882_) );
NAND2X1 NAND2X1_239 ( .A(_875_), .B(_882_), .Y(asr1_q_5_) );
INVX1 INVX1_313 ( .A(asr1_cables_1__6_), .Y(_883_) );
INVX1 INVX1_314 ( .A(asr1_cables_2__6_), .Y(_884_) );
OAI22X1 OAI22X1_29 ( .A(_884_), .B(_915_), .C(_883_), .D(_917_), .Y(_885_) );
INVX1 INVX1_315 ( .A(asr1_cables_7__6_), .Y(_886_) );
INVX1 INVX1_316 ( .A(asr1_cables_3__6_), .Y(_887_) );
OAI22X1 OAI22X1_30 ( .A(_886_), .B(_922_), .C(_887_), .D(_921_), .Y(_888_) );
NOR2X1 NOR2X1_24 ( .A(_888_), .B(_885_), .Y(_889_) );
INVX1 INVX1_317 ( .A(asr1_cables_5__6_), .Y(_890_) );
INVX1 INVX1_318 ( .A(_80_), .Y(_891_) );
OAI22X1 OAI22X1_31 ( .A(_891_), .B(_804_), .C(_890_), .D(_805_), .Y(_892_) );
INVX1 INVX1_319 ( .A(asr1_cables_8__6_), .Y(_893_) );
INVX1 INVX1_320 ( .A(asr1_cables_6__6_), .Y(_894_) );
OAI22X1 OAI22X1_32 ( .A(_893_), .B(_809_), .C(_894_), .D(_810_), .Y(_895_) );
NOR2X1 NOR2X1_25 ( .A(_895_), .B(_892_), .Y(_896_) );
NAND2X1 NAND2X1_240 ( .A(_896_), .B(_889_), .Y(asr1_q_6_) );
INVX1 INVX1_321 ( .A(asr1_cables_3__7_), .Y(_897_) );
INVX1 INVX1_322 ( .A(asr1_cables_2__7_), .Y(_898_) );
OAI22X1 OAI22X1_33 ( .A(_897_), .B(_921_), .C(_898_), .D(_915_), .Y(_899_) );
INVX1 INVX1_323 ( .A(asr1_cables_7__7_), .Y(_900_) );
INVX1 INVX1_324 ( .A(asr1_cables_6__7_), .Y(_901_) );
OAI22X1 OAI22X1_34 ( .A(_900_), .B(_922_), .C(_901_), .D(_810_), .Y(_902_) );
NOR2X1 NOR2X1_26 ( .A(_902_), .B(_899_), .Y(_903_) );
INVX1 INVX1_325 ( .A(asr1_cables_5__7_), .Y(_904_) );
INVX1 INVX1_326 ( .A(_81_), .Y(_905_) );
OAI22X1 OAI22X1_35 ( .A(_905_), .B(_804_), .C(_904_), .D(_805_), .Y(_906_) );
INVX1 INVX1_327 ( .A(asr1_cables_8__7_), .Y(_907_) );
INVX1 INVX1_328 ( .A(asr1_cables_1__7_), .Y(_908_) );
OAI22X1 OAI22X1_36 ( .A(_907_), .B(_809_), .C(_908_), .D(_917_), .Y(_909_) );
NOR2X1 NOR2X1_27 ( .A(_906_), .B(_909_), .Y(_910_) );
NAND2X1 NAND2X1_241 ( .A(_903_), .B(_910_), .Y(asr1_q_7_) );
INVX1 INVX1_329 ( .A(asr2_cables_1__0_), .Y(_1034_) );
INVX1 INVX1_330 ( .A(asr2_cables_2__0_), .Y(_1035_) );
INVX1 INVX1_331 ( .A(down_counter_contador_1_), .Y(_1036_) );
INVX1 INVX1_332 ( .A(down_counter_contador_2_), .Y(_1037_) );
NAND3X1 NAND3X1_119 ( .A(down_counter_contador_0_), .B(_1036_), .C(_1037_), .Y(_1038_) );
INVX1 INVX1_333 ( .A(down_counter_contador_0_), .Y(_1039_) );
NAND3X1 NAND3X1_120 ( .A(_1039_), .B(_1036_), .C(_1037_), .Y(_1040_) );
OAI22X1 OAI22X1_37 ( .A(_1035_), .B(_1038_), .C(_1034_), .D(_1040_), .Y(_1041_) );
INVX1 INVX1_334 ( .A(asr2_cables_7__0_), .Y(_1042_) );
INVX1 INVX1_335 ( .A(asr2_cables_3__0_), .Y(_1043_) );
NAND3X1 NAND3X1_121 ( .A(down_counter_contador_1_), .B(_1039_), .C(_1037_), .Y(_1044_) );
NAND3X1 NAND3X1_122 ( .A(down_counter_contador_1_), .B(down_counter_contador_2_), .C(_1039_), .Y(_1045_) );
OAI22X1 OAI22X1_38 ( .A(_1042_), .B(_1045_), .C(_1043_), .D(_1044_), .Y(_1046_) );
NOR2X1 NOR2X1_28 ( .A(_1046_), .B(_1041_), .Y(_1047_) );
INVX1 INVX1_336 ( .A(asr2_cables_5__0_), .Y(_1048_) );
INVX1 INVX1_337 ( .A(asr2_cables_4_), .Y(_1049_) );
NAND3X1 NAND3X1_123 ( .A(down_counter_contador_0_), .B(down_counter_contador_1_), .C(_1037_), .Y(_927_) );
NAND3X1 NAND3X1_124 ( .A(down_counter_contador_2_), .B(_1039_), .C(_1036_), .Y(_928_) );
OAI22X1 OAI22X1_39 ( .A(_1049_), .B(_927_), .C(_1048_), .D(_928_), .Y(_929_) );
INVX1 INVX1_338 ( .A(asr2_cables_8__0_), .Y(_930_) );
INVX1 INVX1_339 ( .A(asr2_cables_6__0_), .Y(_931_) );
NAND3X1 NAND3X1_125 ( .A(down_counter_contador_0_), .B(down_counter_contador_1_), .C(down_counter_contador_2_), .Y(_932_) );
NAND3X1 NAND3X1_126 ( .A(down_counter_contador_0_), .B(down_counter_contador_2_), .C(_1036_), .Y(_933_) );
OAI22X1 OAI22X1_40 ( .A(_930_), .B(_932_), .C(_931_), .D(_933_), .Y(_934_) );
NOR2X1 NOR2X1_29 ( .A(_934_), .B(_929_), .Y(_935_) );
NAND2X1 NAND2X1_242 ( .A(_935_), .B(_1047_), .Y(asr2_q_0_) );
INVX1 INVX1_340 ( .A(asr2_cables_1__1_), .Y(_936_) );
INVX1 INVX1_341 ( .A(asr2_cables_2__1_), .Y(_937_) );
OAI22X1 OAI22X1_41 ( .A(_937_), .B(_1038_), .C(_936_), .D(_1040_), .Y(_938_) );
INVX1 INVX1_342 ( .A(asr2_cables_6__1_), .Y(_939_) );
INVX1 INVX1_343 ( .A(asr2_cables_3__1_), .Y(_940_) );
OAI22X1 OAI22X1_42 ( .A(_939_), .B(_933_), .C(_940_), .D(_1044_), .Y(_941_) );
NOR2X1 NOR2X1_30 ( .A(_941_), .B(_938_), .Y(_942_) );
INVX1 INVX1_344 ( .A(asr2_cables_7__1_), .Y(_943_) );
INVX1 INVX1_345 ( .A(asr2_cables_8__1_), .Y(_944_) );
OAI22X1 OAI22X1_43 ( .A(_944_), .B(_932_), .C(_943_), .D(_1045_), .Y(_945_) );
INVX1 INVX1_346 ( .A(asr2_cables_5__1_), .Y(_946_) );
INVX1 INVX1_347 ( .A(_227_), .Y(_947_) );
OAI22X1 OAI22X1_44 ( .A(_947_), .B(_927_), .C(_946_), .D(_928_), .Y(_948_) );
NOR2X1 NOR2X1_31 ( .A(_945_), .B(_948_), .Y(_949_) );
NAND2X1 NAND2X1_243 ( .A(_949_), .B(_942_), .Y(asr2_q_1_) );
INVX1 INVX1_348 ( .A(asr2_cables_1__2_), .Y(_950_) );
INVX1 INVX1_349 ( .A(asr2_cables_2__2_), .Y(_951_) );
OAI22X1 OAI22X1_45 ( .A(_951_), .B(_1038_), .C(_950_), .D(_1040_), .Y(_952_) );
INVX1 INVX1_350 ( .A(asr2_cables_7__2_), .Y(_953_) );
INVX1 INVX1_351 ( .A(asr2_cables_3__2_), .Y(_954_) );
OAI22X1 OAI22X1_46 ( .A(_953_), .B(_1045_), .C(_954_), .D(_1044_), .Y(_955_) );
NOR2X1 NOR2X1_32 ( .A(_955_), .B(_952_), .Y(_956_) );
INVX1 INVX1_352 ( .A(asr2_cables_5__2_), .Y(_957_) );
INVX1 INVX1_353 ( .A(_233_), .Y(_958_) );
OAI22X1 OAI22X1_47 ( .A(_958_), .B(_927_), .C(_957_), .D(_928_), .Y(_959_) );
INVX1 INVX1_354 ( .A(asr2_cables_8__2_), .Y(_960_) );
INVX1 INVX1_355 ( .A(asr2_cables_6__2_), .Y(_961_) );
OAI22X1 OAI22X1_48 ( .A(_960_), .B(_932_), .C(_961_), .D(_933_), .Y(_962_) );
NOR2X1 NOR2X1_33 ( .A(_962_), .B(_959_), .Y(_963_) );
NAND2X1 NAND2X1_244 ( .A(_963_), .B(_956_), .Y(asr2_q_2_) );
INVX1 INVX1_356 ( .A(asr2_cables_3__3_), .Y(_964_) );
INVX1 INVX1_357 ( .A(asr2_cables_2__3_), .Y(_965_) );
OAI22X1 OAI22X1_49 ( .A(_964_), .B(_1044_), .C(_965_), .D(_1038_), .Y(_966_) );
INVX1 INVX1_358 ( .A(asr2_cables_7__3_), .Y(_967_) );
INVX1 INVX1_359 ( .A(asr2_cables_6__3_), .Y(_968_) );
OAI22X1 OAI22X1_50 ( .A(_967_), .B(_1045_), .C(_968_), .D(_933_), .Y(_969_) );
NOR2X1 NOR2X1_34 ( .A(_969_), .B(_966_), .Y(_970_) );
INVX1 INVX1_360 ( .A(asr2_cables_5__3_), .Y(_971_) );
INVX1 INVX1_361 ( .A(_228_), .Y(_972_) );
OAI22X1 OAI22X1_51 ( .A(_972_), .B(_927_), .C(_971_), .D(_928_), .Y(_973_) );
INVX1 INVX1_362 ( .A(asr2_cables_8__3_), .Y(_974_) );
INVX1 INVX1_363 ( .A(asr2_cables_1__3_), .Y(_975_) );
OAI22X1 OAI22X1_52 ( .A(_974_), .B(_932_), .C(_975_), .D(_1040_), .Y(_976_) );
NOR2X1 NOR2X1_35 ( .A(_973_), .B(_976_), .Y(_977_) );
NAND2X1 NAND2X1_245 ( .A(_970_), .B(_977_), .Y(asr2_q_3_) );
INVX1 INVX1_364 ( .A(asr2_cables_1__4_), .Y(_978_) );
INVX1 INVX1_365 ( .A(asr2_cables_2__4_), .Y(_979_) );
OAI22X1 OAI22X1_53 ( .A(_979_), .B(_1038_), .C(_978_), .D(_1040_), .Y(_980_) );
INVX1 INVX1_366 ( .A(asr2_cables_7__4_), .Y(_981_) );
INVX1 INVX1_367 ( .A(asr2_cables_3__4_), .Y(_982_) );
OAI22X1 OAI22X1_54 ( .A(_981_), .B(_1045_), .C(_982_), .D(_1044_), .Y(_983_) );
NOR2X1 NOR2X1_36 ( .A(_983_), .B(_980_), .Y(_984_) );
INVX1 INVX1_368 ( .A(asr2_cables_5__4_), .Y(_985_) );
INVX1 INVX1_369 ( .A(_229_), .Y(_986_) );
OAI22X1 OAI22X1_55 ( .A(_986_), .B(_927_), .C(_985_), .D(_928_), .Y(_987_) );
INVX1 INVX1_370 ( .A(asr2_cables_8__4_), .Y(_988_) );
INVX1 INVX1_371 ( .A(asr2_cables_6__4_), .Y(_989_) );
OAI22X1 OAI22X1_56 ( .A(_988_), .B(_932_), .C(_989_), .D(_933_), .Y(_990_) );
NOR2X1 NOR2X1_37 ( .A(_990_), .B(_987_), .Y(_991_) );
NAND2X1 NAND2X1_246 ( .A(_991_), .B(_984_), .Y(asr2_q_4_) );
INVX1 INVX1_372 ( .A(asr2_cables_3__5_), .Y(_992_) );
INVX1 INVX1_373 ( .A(asr2_cables_2__5_), .Y(_993_) );
OAI22X1 OAI22X1_57 ( .A(_992_), .B(_1044_), .C(_993_), .D(_1038_), .Y(_994_) );
INVX1 INVX1_374 ( .A(asr2_cables_7__5_), .Y(_995_) );
INVX1 INVX1_375 ( .A(asr2_cables_6__5_), .Y(_996_) );
OAI22X1 OAI22X1_58 ( .A(_995_), .B(_1045_), .C(_996_), .D(_933_), .Y(_997_) );
NOR2X1 NOR2X1_38 ( .A(_997_), .B(_994_), .Y(_998_) );
INVX1 INVX1_376 ( .A(asr2_cables_5__5_), .Y(_999_) );
INVX1 INVX1_377 ( .A(_230_), .Y(_1000_) );
OAI22X1 OAI22X1_59 ( .A(_1000_), .B(_927_), .C(_999_), .D(_928_), .Y(_1001_) );
INVX1 INVX1_378 ( .A(asr2_cables_8__5_), .Y(_1002_) );
INVX1 INVX1_379 ( .A(asr2_cables_1__5_), .Y(_1003_) );
OAI22X1 OAI22X1_60 ( .A(_1002_), .B(_932_), .C(_1003_), .D(_1040_), .Y(_1004_) );
NOR2X1 NOR2X1_39 ( .A(_1001_), .B(_1004_), .Y(_1005_) );
NAND2X1 NAND2X1_247 ( .A(_998_), .B(_1005_), .Y(asr2_q_5_) );
INVX1 INVX1_380 ( .A(asr2_cables_1__6_), .Y(_1006_) );
INVX1 INVX1_381 ( .A(asr2_cables_2__6_), .Y(_1007_) );
OAI22X1 OAI22X1_61 ( .A(_1007_), .B(_1038_), .C(_1006_), .D(_1040_), .Y(_1008_) );
INVX1 INVX1_382 ( .A(asr2_cables_7__6_), .Y(_1009_) );
INVX1 INVX1_383 ( .A(asr2_cables_3__6_), .Y(_1010_) );
OAI22X1 OAI22X1_62 ( .A(_1009_), .B(_1045_), .C(_1010_), .D(_1044_), .Y(_1011_) );
NOR2X1 NOR2X1_40 ( .A(_1011_), .B(_1008_), .Y(_1012_) );
INVX1 INVX1_384 ( .A(asr2_cables_5__6_), .Y(_1013_) );
INVX1 INVX1_385 ( .A(_231_), .Y(_1014_) );
OAI22X1 OAI22X1_63 ( .A(_1014_), .B(_927_), .C(_1013_), .D(_928_), .Y(_1015_) );
INVX1 INVX1_386 ( .A(asr2_cables_8__6_), .Y(_1016_) );
INVX1 INVX1_387 ( .A(asr2_cables_6__6_), .Y(_1017_) );
OAI22X1 OAI22X1_64 ( .A(_1016_), .B(_932_), .C(_1017_), .D(_933_), .Y(_1018_) );
NOR2X1 NOR2X1_41 ( .A(_1018_), .B(_1015_), .Y(_1019_) );
NAND2X1 NAND2X1_248 ( .A(_1019_), .B(_1012_), .Y(asr2_q_6_) );
INVX1 INVX1_388 ( .A(asr2_cables_3__7_), .Y(_1020_) );
INVX1 INVX1_389 ( .A(asr2_cables_2__7_), .Y(_1021_) );
OAI22X1 OAI22X1_65 ( .A(_1020_), .B(_1044_), .C(_1021_), .D(_1038_), .Y(_1022_) );
INVX1 INVX1_390 ( .A(asr2_cables_7__7_), .Y(_1023_) );
INVX1 INVX1_391 ( .A(asr2_cables_6__7_), .Y(_1024_) );
OAI22X1 OAI22X1_66 ( .A(_1023_), .B(_1045_), .C(_1024_), .D(_933_), .Y(_1025_) );
NOR2X1 NOR2X1_42 ( .A(_1025_), .B(_1022_), .Y(_1026_) );
INVX1 INVX1_392 ( .A(asr2_cables_5__7_), .Y(_1027_) );
INVX1 INVX1_393 ( .A(_232_), .Y(_1028_) );
OAI22X1 OAI22X1_67 ( .A(_1028_), .B(_927_), .C(_1027_), .D(_928_), .Y(_1029_) );
INVX1 INVX1_394 ( .A(asr2_cables_8__7_), .Y(_1030_) );
INVX1 INVX1_395 ( .A(asr2_cables_1__7_), .Y(_1031_) );
OAI22X1 OAI22X1_68 ( .A(_1030_), .B(_932_), .C(_1031_), .D(_1040_), .Y(_1032_) );
NOR2X1 NOR2X1_43 ( .A(_1029_), .B(_1032_), .Y(_1033_) );
NAND2X1 NAND2X1_249 ( .A(_1026_), .B(_1033_), .Y(asr2_q_7_) );
INVX1 INVX1_396 ( .A(rst_bF_buf2), .Y(_1057_) );
NAND2X1 NAND2X1_250 ( .A(down_counter_contador_0_), .B(_1057_), .Y(_1050__0_) );
AOI21X1 AOI21X1_40 ( .A(down_counter_contador_0_), .B(down_counter_contador_1_), .C(rst_bF_buf2), .Y(_1051_) );
OAI21X1 OAI21X1_239 ( .A(down_counter_contador_0_), .B(down_counter_contador_1_), .C(_1051_), .Y(_1050__1_) );
OAI21X1 OAI21X1_240 ( .A(down_counter_contador_0_), .B(down_counter_contador_1_), .C(down_counter_contador_2_), .Y(_1052_) );
INVX1 INVX1_397 ( .A(down_counter_contador_0_), .Y(_1053_) );
INVX1 INVX1_398 ( .A(down_counter_contador_1_), .Y(_1054_) );
INVX1 INVX1_399 ( .A(down_counter_contador_2_), .Y(_1055_) );
NAND3X1 NAND3X1_127 ( .A(_1053_), .B(_1054_), .C(_1055_), .Y(_1056_) );
NAND3X1 NAND3X1_128 ( .A(_1057_), .B(_1052_), .C(_1056_), .Y(_1050__2_) );
DFFPOSX1 DFFPOSX1_10 ( .CLK(clk_bF_buf7), .D(_1050__0_), .Q(down_counter_contador_0_) );
DFFPOSX1 DFFPOSX1_11 ( .CLK(clk_bF_buf3), .D(_1050__1_), .Q(down_counter_contador_1_) );
DFFPOSX1 DFFPOSX1_12 ( .CLK(clk_bF_buf7), .D(_1050__2_), .Q(down_counter_contador_2_) );
NOR2X1 NOR2X1_44 ( .A(generador_clock_counter_0_), .B(rst_bF_buf4), .Y(_1058__0_) );
AND2X2 AND2X2_14 ( .A(generador_clock_counter_0_), .B(generador_clock_counter_1_), .Y(_1059_) );
INVX1 INVX1_400 ( .A(rst_bF_buf4), .Y(_1060_) );
OAI21X1 OAI21X1_241 ( .A(generador_clock_counter_0_), .B(generador_clock_counter_1_), .C(_1060_), .Y(_1061_) );
NOR2X1 NOR2X1_45 ( .A(_1059_), .B(_1061_), .Y(_1058__1_) );
INVX1 INVX1_401 ( .A(generador_clock_counter_2_), .Y(_1062_) );
NAND2X1 NAND2X1_251 ( .A(generador_clock_counter_0_), .B(generador_clock_counter_1_), .Y(_1063_) );
OAI21X1 OAI21X1_242 ( .A(_1062_), .B(_1063_), .C(_1060_), .Y(_1064_) );
AOI21X1 AOI21X1_41 ( .A(_1062_), .B(_1063_), .C(_1064_), .Y(_1058__2_) );
OAI21X1 OAI21X1_243 ( .A(_1062_), .B(_1063_), .C(generador_clock_counter_3_), .Y(_1065_) );
INVX1 INVX1_402 ( .A(generador_clock_counter_3_), .Y(asr1_clk) );
NAND3X1 NAND3X1_129 ( .A(asr1_clk_bF_buf0), .B(generador_clock_counter_2_), .C(_1059_), .Y(_1066_) );
AOI21X1 AOI21X1_42 ( .A(_1066_), .B(_1065_), .C(rst_bF_buf4), .Y(_1058__3_) );
DFFPOSX1 DFFPOSX1_13 ( .CLK(clk_bF_buf4), .D(_1058__0_), .Q(generador_clock_counter_0_) );
DFFPOSX1 DFFPOSX1_14 ( .CLK(clk_bF_buf4), .D(_1058__1_), .Q(generador_clock_counter_1_) );
DFFPOSX1 DFFPOSX1_15 ( .CLK(clk_bF_buf2), .D(_1058__2_), .Q(generador_clock_counter_2_) );
DFFPOSX1 DFFPOSX1_16 ( .CLK(clk_bF_buf2), .D(_1058__3_), .Q(generador_clock_counter_3_) );
INVX1 INVX1_403 ( .A(up_counter_contador_0_), .Y(_1067_) );
INVX1 INVX1_404 ( .A(up_counter_contador_2_), .Y(_1075_) );
NAND3X1 NAND3X1_130 ( .A(up_counter_contador_0_), .B(up_counter_contador_1_), .C(_1075_), .Y(_1071_) );
NAND2X1 NAND2X1_252 ( .A(up_counter_contador_0_), .B(up_counter_contador_1_), .Y(_1072_) );
NAND2X1 NAND2X1_253 ( .A(up_counter_contador_2_), .B(_1072_), .Y(_1073_) );
NAND2X1 NAND2X1_254 ( .A(_1073_), .B(_1071_), .Y(_1069_) );
NAND3X1 NAND3X1_131 ( .A(up_counter_contador_0_), .B(up_counter_contador_1_), .C(up_counter_contador_2_), .Y(_1074_) );
INVX1 INVX1_405 ( .A(_1074_), .Y(_1070_) );
XOR2X1 XOR2X1_9 ( .A(up_counter_contador_0_), .B(up_counter_contador_1_), .Y(_1068_) );
DFFPOSX1 DFFPOSX1_17 ( .CLK(clk_bF_buf0), .D(_1067_), .Q(memoria_q_0_) );
DFFPOSX1 DFFPOSX1_18 ( .CLK(clk_bF_buf0), .D(_1068_), .Q(memoria_q_1_) );
DFFPOSX1 DFFPOSX1_19 ( .CLK(clk_bF_buf6), .D(_1069_), .Q(memoria_q_2_) );
DFFPOSX1 DFFPOSX1_20 ( .CLK(clk_bF_buf0), .D(_1070_), .Q(memoria_q_3_) );
INVX1 INVX1_406 ( .A(asr1_cables_0__0_), .Y(_1078_) );
NAND2X1 NAND2X1_255 ( .A(din[0]), .B(vdd), .Y(_1079_) );
OAI21X1 OAI21X1_244 ( .A(vdd), .B(_1078_), .C(_1079_), .Y(_1076__0_) );
INVX1 INVX1_407 ( .A(asr1_cables_0__1_), .Y(_1080_) );
NAND2X1 NAND2X1_256 ( .A(vdd), .B(din[1]), .Y(_1081_) );
OAI21X1 OAI21X1_245 ( .A(vdd), .B(_1080_), .C(_1081_), .Y(_1076__1_) );
INVX1 INVX1_408 ( .A(asr1_cables_0__2_), .Y(_1082_) );
NAND2X1 NAND2X1_257 ( .A(vdd), .B(din[2]), .Y(_1083_) );
OAI21X1 OAI21X1_246 ( .A(vdd), .B(_1082_), .C(_1083_), .Y(_1076__2_) );
INVX1 INVX1_409 ( .A(asr1_cables_0__3_), .Y(_1084_) );
NAND2X1 NAND2X1_258 ( .A(vdd), .B(din[3]), .Y(_1085_) );
OAI21X1 OAI21X1_247 ( .A(vdd), .B(_1084_), .C(_1085_), .Y(_1076__3_) );
INVX1 INVX1_410 ( .A(asr1_cables_0__4_), .Y(_1086_) );
NAND2X1 NAND2X1_259 ( .A(vdd), .B(din[4]), .Y(_1087_) );
OAI21X1 OAI21X1_248 ( .A(vdd), .B(_1086_), .C(_1087_), .Y(_1076__4_) );
INVX1 INVX1_411 ( .A(asr1_cables_0__5_), .Y(_1088_) );
NAND2X1 NAND2X1_260 ( .A(vdd), .B(din[5]), .Y(_1089_) );
OAI21X1 OAI21X1_249 ( .A(vdd), .B(_1088_), .C(_1089_), .Y(_1076__5_) );
INVX1 INVX1_412 ( .A(asr1_cables_0__6_), .Y(_1090_) );
NAND2X1 NAND2X1_261 ( .A(vdd), .B(din[6]), .Y(_1091_) );
OAI21X1 OAI21X1_250 ( .A(vdd), .B(_1090_), .C(_1091_), .Y(_1076__6_) );
INVX1 INVX1_413 ( .A(asr1_cables_0__7_), .Y(_1092_) );
NAND2X1 NAND2X1_262 ( .A(vdd), .B(din[7]), .Y(_1093_) );
OAI21X1 OAI21X1_251 ( .A(vdd), .B(_1092_), .C(_1093_), .Y(_1076__7_) );
INVX1 INVX1_414 ( .A(rst_bF_buf2), .Y(_1077_) );
DFFSR DFFSR_176 ( .CLK(asr1_clk_bF_buf7), .D(_1076__0_), .Q(asr1_cables_0__0_), .R(_1077_), .S(vdd) );
DFFSR DFFSR_177 ( .CLK(asr1_clk_bF_buf7), .D(_1076__1_), .Q(asr1_cables_0__1_), .R(_1077_), .S(vdd) );
DFFSR DFFSR_178 ( .CLK(asr1_clk_bF_buf6), .D(_1076__2_), .Q(asr1_cables_0__2_), .R(_1077_), .S(vdd) );
DFFSR DFFSR_179 ( .CLK(asr1_clk_bF_buf6), .D(_1076__3_), .Q(asr1_cables_0__3_), .R(_1077_), .S(vdd) );
DFFSR DFFSR_180 ( .CLK(asr1_clk_bF_buf7), .D(_1076__4_), .Q(asr1_cables_0__4_), .R(_1077_), .S(vdd) );
DFFSR DFFSR_181 ( .CLK(asr1_clk_bF_buf0), .D(_1076__5_), .Q(asr1_cables_0__5_), .R(_1077_), .S(vdd) );
DFFSR DFFSR_182 ( .CLK(asr1_clk_bF_buf7), .D(_1076__6_), .Q(asr1_cables_0__6_), .R(_1077_), .S(vdd) );
DFFSR DFFSR_183 ( .CLK(asr1_clk_bF_buf1), .D(_1076__7_), .Q(asr1_cables_0__7_), .R(_1077_), .S(vdd) );
INVX1 INVX1_415 ( .A(_3__0_), .Y(_1096_) );
NAND2X1 NAND2X1_263 ( .A(registro_salida_d_0_), .B(vdd), .Y(_1097_) );
OAI21X1 OAI21X1_252 ( .A(vdd), .B(_1096_), .C(_1097_), .Y(_1094__0_) );
INVX1 INVX1_416 ( .A(_3__1_), .Y(_1098_) );
NAND2X1 NAND2X1_264 ( .A(vdd), .B(registro_salida_d_1_), .Y(_1099_) );
OAI21X1 OAI21X1_253 ( .A(vdd), .B(_1098_), .C(_1099_), .Y(_1094__1_) );
INVX1 INVX1_417 ( .A(_3__2_), .Y(_1100_) );
NAND2X1 NAND2X1_265 ( .A(vdd), .B(registro_salida_d_2_), .Y(_1101_) );
OAI21X1 OAI21X1_254 ( .A(vdd), .B(_1100_), .C(_1101_), .Y(_1094__2_) );
INVX1 INVX1_418 ( .A(_3__3_), .Y(_1102_) );
NAND2X1 NAND2X1_266 ( .A(vdd), .B(registro_salida_d_3_), .Y(_1103_) );
OAI21X1 OAI21X1_255 ( .A(vdd), .B(_1102_), .C(_1103_), .Y(_1094__3_) );
INVX1 INVX1_419 ( .A(_3__4_), .Y(_1104_) );
NAND2X1 NAND2X1_267 ( .A(vdd), .B(registro_salida_d_4_), .Y(_1105_) );
OAI21X1 OAI21X1_256 ( .A(vdd), .B(_1104_), .C(_1105_), .Y(_1094__4_) );
INVX1 INVX1_420 ( .A(_3__5_), .Y(_1106_) );
NAND2X1 NAND2X1_268 ( .A(vdd), .B(registro_salida_d_5_), .Y(_1107_) );
OAI21X1 OAI21X1_257 ( .A(vdd), .B(_1106_), .C(_1107_), .Y(_1094__5_) );
INVX1 INVX1_421 ( .A(_3__6_), .Y(_1108_) );
NAND2X1 NAND2X1_269 ( .A(vdd), .B(registro_salida_d_6_), .Y(_1109_) );
OAI21X1 OAI21X1_258 ( .A(vdd), .B(_1108_), .C(_1109_), .Y(_1094__6_) );
INVX1 INVX1_422 ( .A(_3__7_), .Y(_1110_) );
NAND2X1 NAND2X1_270 ( .A(vdd), .B(registro_salida_d_7_), .Y(_1111_) );
OAI21X1 OAI21X1_259 ( .A(vdd), .B(_1110_), .C(_1111_), .Y(_1094__7_) );
INVX1 INVX1_423 ( .A(rst_bF_buf3), .Y(_1095_) );
DFFSR DFFSR_184 ( .CLK(asr1_clk_bF_buf6), .D(_1094__0_), .Q(_3__0_), .R(_1095_), .S(vdd) );
DFFSR DFFSR_185 ( .CLK(asr1_clk_bF_buf1), .D(_1094__1_), .Q(_3__1_), .R(_1095_), .S(vdd) );
DFFSR DFFSR_186 ( .CLK(asr1_clk_bF_buf1), .D(_1094__2_), .Q(_3__2_), .R(_1095_), .S(vdd) );
DFFSR DFFSR_187 ( .CLK(asr1_clk_bF_buf7), .D(_1094__3_), .Q(_3__3_), .R(_1095_), .S(vdd) );
DFFSR DFFSR_188 ( .CLK(asr1_clk_bF_buf6), .D(_1094__4_), .Q(_3__4_), .R(_1095_), .S(vdd) );
DFFSR DFFSR_189 ( .CLK(asr1_clk_bF_buf6), .D(_1094__5_), .Q(_3__5_), .R(_1095_), .S(vdd) );
DFFSR DFFSR_190 ( .CLK(asr1_clk_bF_buf6), .D(_1094__6_), .Q(_3__6_), .R(_1095_), .S(vdd) );
DFFSR DFFSR_191 ( .CLK(asr1_clk_bF_buf1), .D(_1094__7_), .Q(_3__7_), .R(_1095_), .S(vdd) );
NAND2X1 NAND2X1_271 ( .A(retardo_asr_1_connect_wire_1__0_), .B(retardo_asr_2_connect_wire_1__0_), .Y(_1112_) );
NOR2X1 NOR2X1_46 ( .A(retardo_asr_1_connect_wire_1__1_), .B(retardo_asr_2_connect_wire_1__1_), .Y(_1113_) );
INVX1 INVX1_424 ( .A(_1113_), .Y(_1114_) );
NAND2X1 NAND2X1_272 ( .A(retardo_asr_1_connect_wire_1__1_), .B(retardo_asr_2_connect_wire_1__1_), .Y(_1115_) );
NAND2X1 NAND2X1_273 ( .A(_1115_), .B(_1114_), .Y(_1116_) );
XOR2X1 XOR2X1_10 ( .A(_1116_), .B(_1112_), .Y(sumador_suma_previa_1_) );
OAI21X1 OAI21X1_260 ( .A(_1112_), .B(_1113_), .C(_1115_), .Y(_1117_) );
XOR2X1 XOR2X1_11 ( .A(retardo_asr_1_connect_wire_1__2_), .B(retardo_asr_2_connect_wire_1__2_), .Y(_1118_) );
XOR2X1 XOR2X1_12 ( .A(_1117_), .B(_1118_), .Y(sumador_suma_previa_2_) );
AND2X2 AND2X2_15 ( .A(retardo_asr_1_connect_wire_1__2_), .B(retardo_asr_2_connect_wire_1__2_), .Y(_1119_) );
AOI21X1 AOI21X1_43 ( .A(_1117_), .B(_1118_), .C(_1119_), .Y(_1120_) );
XOR2X1 XOR2X1_13 ( .A(retardo_asr_1_connect_wire_1__3_), .B(retardo_asr_2_connect_wire_1__3_), .Y(_1121_) );
XNOR2X1 XNOR2X1_4 ( .A(_1120_), .B(_1121_), .Y(sumador_suma_previa_3_) );
NAND3X1 NAND3X1_132 ( .A(_1118_), .B(_1121_), .C(_1117_), .Y(_1122_) );
INVX1 INVX1_425 ( .A(retardo_asr_1_connect_wire_1__3_), .Y(_1123_) );
INVX1 INVX1_426 ( .A(retardo_asr_2_connect_wire_1__3_), .Y(_1124_) );
NAND2X1 NAND2X1_274 ( .A(_1123_), .B(_1124_), .Y(_1125_) );
NOR2X1 NOR2X1_47 ( .A(_1123_), .B(_1124_), .Y(_1126_) );
AOI21X1 AOI21X1_44 ( .A(_1119_), .B(_1125_), .C(_1126_), .Y(_1127_) );
NAND2X1 NAND2X1_275 ( .A(_1127_), .B(_1122_), .Y(_1128_) );
INVX1 INVX1_427 ( .A(retardo_asr_1_connect_wire_1__4_), .Y(_1129_) );
INVX1 INVX1_428 ( .A(retardo_asr_2_connect_wire_1__4_), .Y(_1130_) );
NAND2X1 NAND2X1_276 ( .A(_1129_), .B(_1130_), .Y(_1131_) );
NAND2X1 NAND2X1_277 ( .A(retardo_asr_1_connect_wire_1__4_), .B(retardo_asr_2_connect_wire_1__4_), .Y(_1132_) );
AND2X2 AND2X2_16 ( .A(_1131_), .B(_1132_), .Y(_1133_) );
XOR2X1 XOR2X1_14 ( .A(_1128_), .B(_1133_), .Y(sumador_suma_previa_4_) );
AND2X2 AND2X2_17 ( .A(_1122_), .B(_1127_), .Y(_1134_) );
NAND2X1 NAND2X1_278 ( .A(_1132_), .B(_1131_), .Y(_1135_) );
OAI21X1 OAI21X1_261 ( .A(_1135_), .B(_1134_), .C(_1132_), .Y(_1136_) );
INVX1 INVX1_429 ( .A(retardo_asr_1_connect_wire_1__5_), .Y(_1137_) );
INVX1 INVX1_430 ( .A(retardo_asr_2_connect_wire_1__5_), .Y(_1138_) );
NOR2X1 NOR2X1_48 ( .A(_1137_), .B(_1138_), .Y(_1139_) );
NOR2X1 NOR2X1_49 ( .A(retardo_asr_1_connect_wire_1__5_), .B(retardo_asr_2_connect_wire_1__5_), .Y(_1140_) );
NOR2X1 NOR2X1_50 ( .A(_1140_), .B(_1139_), .Y(_1141_) );
XOR2X1 XOR2X1_15 ( .A(_1136_), .B(_1141_), .Y(sumador_suma_previa_5_) );
NOR3X1 NOR3X1_2 ( .A(_1139_), .B(_1140_), .C(_1135_), .Y(_1142_) );
NAND2X1 NAND2X1_279 ( .A(_1142_), .B(_1128_), .Y(_1143_) );
INVX1 INVX1_431 ( .A(_1132_), .Y(_1144_) );
AOI21X1 AOI21X1_45 ( .A(_1141_), .B(_1144_), .C(_1139_), .Y(_1145_) );
INVX1 INVX1_432 ( .A(retardo_asr_1_connect_wire_1__6_), .Y(_1146_) );
NAND2X1 NAND2X1_280 ( .A(retardo_asr_2_connect_wire_1__6_), .B(_1146_), .Y(_1147_) );
INVX1 INVX1_433 ( .A(retardo_asr_2_connect_wire_1__6_), .Y(_1148_) );
NAND2X1 NAND2X1_281 ( .A(retardo_asr_1_connect_wire_1__6_), .B(_1148_), .Y(_1149_) );
AOI22X1 AOI22X1_14 ( .A(_1147_), .B(_1149_), .C(_1143_), .D(_1145_), .Y(_1150_) );
NAND2X1 NAND2X1_282 ( .A(_1133_), .B(_1141_), .Y(_1151_) );
OAI21X1 OAI21X1_262 ( .A(_1151_), .B(_1134_), .C(_1145_), .Y(_1152_) );
NAND2X1 NAND2X1_283 ( .A(_1147_), .B(_1149_), .Y(_1153_) );
NOR2X1 NOR2X1_51 ( .A(_1153_), .B(_1152_), .Y(_1154_) );
NOR2X1 NOR2X1_52 ( .A(_1150_), .B(_1154_), .Y(sumador_suma_previa_6_) );
NOR2X1 NOR2X1_53 ( .A(_1146_), .B(_1148_), .Y(_1155_) );
XOR2X1 XOR2X1_16 ( .A(retardo_asr_1_connect_wire_1__7_), .B(retardo_asr_2_connect_wire_1__7_), .Y(_1156_) );
INVX1 INVX1_434 ( .A(_1156_), .Y(_1157_) );
OAI21X1 OAI21X1_263 ( .A(_1155_), .B(_1150_), .C(_1157_), .Y(_1158_) );
INVX1 INVX1_435 ( .A(_1155_), .Y(_1159_) );
AOI21X1 AOI21X1_46 ( .A(_1122_), .B(_1127_), .C(_1151_), .Y(_1160_) );
INVX1 INVX1_436 ( .A(_1145_), .Y(_1161_) );
OAI21X1 OAI21X1_264 ( .A(_1161_), .B(_1160_), .C(_1153_), .Y(_1162_) );
NAND3X1 NAND3X1_133 ( .A(_1159_), .B(_1156_), .C(_1162_), .Y(_1163_) );
NAND2X1 NAND2X1_284 ( .A(_1163_), .B(_1158_), .Y(sumador_suma_previa_7_) );
XOR2X1 XOR2X1_17 ( .A(retardo_asr_1_connect_wire_1__0_), .B(retardo_asr_2_connect_wire_1__0_), .Y(sumador_suma_previa_0_) );
DFFPOSX1 DFFPOSX1_21 ( .CLK(clk_bF_buf5), .D(sumador_suma_previa_0_), .Q(MAC_Adder_0_) );
DFFPOSX1 DFFPOSX1_22 ( .CLK(clk_bF_buf3), .D(sumador_suma_previa_1_), .Q(MAC_Adder_1_) );
DFFPOSX1 DFFPOSX1_23 ( .CLK(clk_bF_buf2), .D(sumador_suma_previa_2_), .Q(MAC_Adder_2_) );
DFFPOSX1 DFFPOSX1_24 ( .CLK(clk_bF_buf0), .D(sumador_suma_previa_3_), .Q(MAC_Adder_3_) );
DFFPOSX1 DFFPOSX1_25 ( .CLK(clk_bF_buf0), .D(sumador_suma_previa_4_), .Q(MAC_Adder_4_) );
DFFPOSX1 DFFPOSX1_26 ( .CLK(clk_bF_buf0), .D(sumador_suma_previa_5_), .Q(MAC_Adder_5_) );
DFFPOSX1 DFFPOSX1_27 ( .CLK(clk_bF_buf1), .D(sumador_suma_previa_6_), .Q(MAC_Adder_6_) );
DFFPOSX1 DFFPOSX1_28 ( .CLK(clk_bF_buf6), .D(sumador_suma_previa_7_), .Q(MAC_Adder_7_) );
NOR2X1 NOR2X1_54 ( .A(up_counter_contador_0_), .B(rst_bF_buf2), .Y(_1164__0_) );
INVX1 INVX1_437 ( .A(rst_bF_buf4), .Y(_1170_) );
OAI21X1 OAI21X1_265 ( .A(up_counter_contador_0_), .B(up_counter_contador_1_), .C(_1170_), .Y(_1165_) );
AOI21X1 AOI21X1_47 ( .A(up_counter_contador_0_), .B(up_counter_contador_1_), .C(_1165_), .Y(_1164__1_) );
NAND2X1 NAND2X1_285 ( .A(up_counter_contador_0_), .B(up_counter_contador_1_), .Y(_1166_) );
NAND2X1 NAND2X1_286 ( .A(up_counter_contador_2_), .B(_1166_), .Y(_1167_) );
INVX1 INVX1_438 ( .A(up_counter_contador_2_), .Y(_1168_) );
NAND3X1 NAND3X1_134 ( .A(up_counter_contador_0_), .B(up_counter_contador_1_), .C(_1168_), .Y(_1169_) );
AOI21X1 AOI21X1_48 ( .A(_1169_), .B(_1167_), .C(rst_bF_buf0), .Y(_1164__2_) );
DFFPOSX1 DFFPOSX1_29 ( .CLK(clk_bF_buf3), .D(_1164__0_), .Q(up_counter_contador_0_) );
DFFPOSX1 DFFPOSX1_30 ( .CLK(clk_bF_buf5), .D(_1164__1_), .Q(up_counter_contador_1_) );
DFFPOSX1 DFFPOSX1_31 ( .CLK(clk_bF_buf3), .D(_1164__2_), .Q(up_counter_contador_2_) );
BUFX2 BUFX2_34 ( .A(gnd), .Y(MAC_salida_correcta_8_) );
BUFX2 BUFX2_35 ( .A(gnd), .Y(MAC_salida_correcta_9_) );
BUFX2 BUFX2_36 ( .A(gnd), .Y(MAC_salida_correcta_10_) );
BUFX2 BUFX2_37 ( .A(gnd), .Y(MAC_salida_correcta_11_) );
BUFX2 BUFX2_38 ( .A(gnd), .Y(MAC_salida_correcta_12_) );
BUFX2 BUFX2_39 ( .A(gnd), .Y(MAC_salida_correcta_13_) );
BUFX2 BUFX2_40 ( .A(gnd), .Y(MAC_salida_correcta_14_) );
BUFX2 BUFX2_41 ( .A(gnd), .Y(MAC_salida_correcta_15_) );
BUFX2 BUFX2_42 ( .A(gnd), .Y(MAC_salida_correcta_16_) );
BUFX2 BUFX2_43 ( .A(gnd), .Y(MAC_salida_correcta_17_) );
FILL FILL_0_DFFSR_89 ( );
FILL FILL_1_DFFSR_89 ( );
FILL FILL_2_DFFSR_89 ( );
FILL FILL_3_DFFSR_89 ( );
FILL FILL_4_DFFSR_89 ( );
FILL FILL_5_DFFSR_89 ( );
FILL FILL_6_DFFSR_89 ( );
FILL FILL_7_DFFSR_89 ( );
FILL FILL_8_DFFSR_89 ( );
FILL FILL_9_DFFSR_89 ( );
FILL FILL_10_DFFSR_89 ( );
FILL FILL_11_DFFSR_89 ( );
FILL FILL_12_DFFSR_89 ( );
FILL FILL_13_DFFSR_89 ( );
FILL FILL_14_DFFSR_89 ( );
FILL FILL_15_DFFSR_89 ( );
FILL FILL_16_DFFSR_89 ( );
FILL FILL_17_DFFSR_89 ( );
FILL FILL_18_DFFSR_89 ( );
FILL FILL_19_DFFSR_89 ( );
FILL FILL_20_DFFSR_89 ( );
FILL FILL_21_DFFSR_89 ( );
FILL FILL_22_DFFSR_89 ( );
FILL FILL_23_DFFSR_89 ( );
FILL FILL_24_DFFSR_89 ( );
FILL FILL_25_DFFSR_89 ( );
FILL FILL_26_DFFSR_89 ( );
FILL FILL_27_DFFSR_89 ( );
FILL FILL_28_DFFSR_89 ( );
FILL FILL_29_DFFSR_89 ( );
FILL FILL_30_DFFSR_89 ( );
FILL FILL_31_DFFSR_89 ( );
FILL FILL_32_DFFSR_89 ( );
FILL FILL_33_DFFSR_89 ( );
FILL FILL_34_DFFSR_89 ( );
FILL FILL_35_DFFSR_89 ( );
FILL FILL_36_DFFSR_89 ( );
FILL FILL_37_DFFSR_89 ( );
FILL FILL_38_DFFSR_89 ( );
FILL FILL_39_DFFSR_89 ( );
FILL FILL_40_DFFSR_89 ( );
FILL FILL_41_DFFSR_89 ( );
FILL FILL_42_DFFSR_89 ( );
FILL FILL_43_DFFSR_89 ( );
FILL FILL_44_DFFSR_89 ( );
FILL FILL_45_DFFSR_89 ( );
FILL FILL_46_DFFSR_89 ( );
FILL FILL_47_DFFSR_89 ( );
FILL FILL_48_DFFSR_89 ( );
FILL FILL_49_DFFSR_89 ( );
FILL FILL_50_DFFSR_89 ( );
FILL FILL_0_DFFSR_92 ( );
FILL FILL_1_DFFSR_92 ( );
FILL FILL_2_DFFSR_92 ( );
FILL FILL_3_DFFSR_92 ( );
FILL FILL_4_DFFSR_92 ( );
FILL FILL_5_DFFSR_92 ( );
FILL FILL_6_DFFSR_92 ( );
FILL FILL_7_DFFSR_92 ( );
FILL FILL_8_DFFSR_92 ( );
FILL FILL_9_DFFSR_92 ( );
FILL FILL_10_DFFSR_92 ( );
FILL FILL_11_DFFSR_92 ( );
FILL FILL_12_DFFSR_92 ( );
FILL FILL_13_DFFSR_92 ( );
FILL FILL_14_DFFSR_92 ( );
FILL FILL_15_DFFSR_92 ( );
FILL FILL_16_DFFSR_92 ( );
FILL FILL_17_DFFSR_92 ( );
FILL FILL_18_DFFSR_92 ( );
FILL FILL_19_DFFSR_92 ( );
FILL FILL_20_DFFSR_92 ( );
FILL FILL_21_DFFSR_92 ( );
FILL FILL_22_DFFSR_92 ( );
FILL FILL_23_DFFSR_92 ( );
FILL FILL_24_DFFSR_92 ( );
FILL FILL_25_DFFSR_92 ( );
FILL FILL_26_DFFSR_92 ( );
FILL FILL_27_DFFSR_92 ( );
FILL FILL_28_DFFSR_92 ( );
FILL FILL_29_DFFSR_92 ( );
FILL FILL_30_DFFSR_92 ( );
FILL FILL_31_DFFSR_92 ( );
FILL FILL_32_DFFSR_92 ( );
FILL FILL_33_DFFSR_92 ( );
FILL FILL_34_DFFSR_92 ( );
FILL FILL_35_DFFSR_92 ( );
FILL FILL_36_DFFSR_92 ( );
FILL FILL_37_DFFSR_92 ( );
FILL FILL_38_DFFSR_92 ( );
FILL FILL_39_DFFSR_92 ( );
FILL FILL_40_DFFSR_92 ( );
FILL FILL_41_DFFSR_92 ( );
FILL FILL_42_DFFSR_92 ( );
FILL FILL_43_DFFSR_92 ( );
FILL FILL_44_DFFSR_92 ( );
FILL FILL_45_DFFSR_92 ( );
FILL FILL_46_DFFSR_92 ( );
FILL FILL_47_DFFSR_92 ( );
FILL FILL_48_DFFSR_92 ( );
FILL FILL_49_DFFSR_92 ( );
FILL FILL_50_DFFSR_92 ( );
FILL FILL_0_DFFSR_148 ( );
FILL FILL_1_DFFSR_148 ( );
FILL FILL_2_DFFSR_148 ( );
FILL FILL_3_DFFSR_148 ( );
FILL FILL_4_DFFSR_148 ( );
FILL FILL_5_DFFSR_148 ( );
FILL FILL_6_DFFSR_148 ( );
FILL FILL_7_DFFSR_148 ( );
FILL FILL_8_DFFSR_148 ( );
FILL FILL_9_DFFSR_148 ( );
FILL FILL_10_DFFSR_148 ( );
FILL FILL_11_DFFSR_148 ( );
FILL FILL_12_DFFSR_148 ( );
FILL FILL_13_DFFSR_148 ( );
FILL FILL_14_DFFSR_148 ( );
FILL FILL_15_DFFSR_148 ( );
FILL FILL_16_DFFSR_148 ( );
FILL FILL_17_DFFSR_148 ( );
FILL FILL_18_DFFSR_148 ( );
FILL FILL_19_DFFSR_148 ( );
FILL FILL_20_DFFSR_148 ( );
FILL FILL_21_DFFSR_148 ( );
FILL FILL_22_DFFSR_148 ( );
FILL FILL_23_DFFSR_148 ( );
FILL FILL_24_DFFSR_148 ( );
FILL FILL_25_DFFSR_148 ( );
FILL FILL_26_DFFSR_148 ( );
FILL FILL_27_DFFSR_148 ( );
FILL FILL_28_DFFSR_148 ( );
FILL FILL_29_DFFSR_148 ( );
FILL FILL_30_DFFSR_148 ( );
FILL FILL_31_DFFSR_148 ( );
FILL FILL_32_DFFSR_148 ( );
FILL FILL_33_DFFSR_148 ( );
FILL FILL_34_DFFSR_148 ( );
FILL FILL_35_DFFSR_148 ( );
FILL FILL_36_DFFSR_148 ( );
FILL FILL_37_DFFSR_148 ( );
FILL FILL_38_DFFSR_148 ( );
FILL FILL_39_DFFSR_148 ( );
FILL FILL_40_DFFSR_148 ( );
FILL FILL_41_DFFSR_148 ( );
FILL FILL_42_DFFSR_148 ( );
FILL FILL_43_DFFSR_148 ( );
FILL FILL_44_DFFSR_148 ( );
FILL FILL_45_DFFSR_148 ( );
FILL FILL_46_DFFSR_148 ( );
FILL FILL_47_DFFSR_148 ( );
FILL FILL_48_DFFSR_148 ( );
FILL FILL_49_DFFSR_148 ( );
FILL FILL_50_DFFSR_148 ( );
FILL FILL_0_NAND2X1_148 ( );
FILL FILL_1_NAND2X1_148 ( );
FILL FILL_2_NAND2X1_148 ( );
FILL FILL_3_NAND2X1_148 ( );
FILL FILL_4_NAND2X1_148 ( );
FILL FILL_5_NAND2X1_148 ( );
FILL FILL_6_NAND2X1_148 ( );
FILL FILL_0_INVX1_167 ( );
FILL FILL_1_INVX1_167 ( );
FILL FILL_2_INVX1_167 ( );
FILL FILL_3_INVX1_167 ( );
FILL FILL_4_INVX1_167 ( );
FILL FILL_0_INVX1_168 ( );
FILL FILL_1_INVX1_168 ( );
FILL FILL_2_INVX1_168 ( );
FILL FILL_3_INVX1_168 ( );
FILL FILL_4_INVX1_168 ( );
FILL FILL_0_DFFSR_146 ( );
FILL FILL_1_DFFSR_146 ( );
FILL FILL_2_DFFSR_146 ( );
FILL FILL_3_DFFSR_146 ( );
FILL FILL_4_DFFSR_146 ( );
FILL FILL_5_DFFSR_146 ( );
FILL FILL_6_DFFSR_146 ( );
FILL FILL_7_DFFSR_146 ( );
FILL FILL_8_DFFSR_146 ( );
FILL FILL_9_DFFSR_146 ( );
FILL FILL_10_DFFSR_146 ( );
FILL FILL_11_DFFSR_146 ( );
FILL FILL_12_DFFSR_146 ( );
FILL FILL_13_DFFSR_146 ( );
FILL FILL_14_DFFSR_146 ( );
FILL FILL_15_DFFSR_146 ( );
FILL FILL_16_DFFSR_146 ( );
FILL FILL_17_DFFSR_146 ( );
FILL FILL_18_DFFSR_146 ( );
FILL FILL_19_DFFSR_146 ( );
FILL FILL_20_DFFSR_146 ( );
FILL FILL_21_DFFSR_146 ( );
FILL FILL_22_DFFSR_146 ( );
FILL FILL_23_DFFSR_146 ( );
FILL FILL_24_DFFSR_146 ( );
FILL FILL_25_DFFSR_146 ( );
FILL FILL_26_DFFSR_146 ( );
FILL FILL_27_DFFSR_146 ( );
FILL FILL_28_DFFSR_146 ( );
FILL FILL_29_DFFSR_146 ( );
FILL FILL_30_DFFSR_146 ( );
FILL FILL_31_DFFSR_146 ( );
FILL FILL_32_DFFSR_146 ( );
FILL FILL_33_DFFSR_146 ( );
FILL FILL_34_DFFSR_146 ( );
FILL FILL_35_DFFSR_146 ( );
FILL FILL_36_DFFSR_146 ( );
FILL FILL_37_DFFSR_146 ( );
FILL FILL_38_DFFSR_146 ( );
FILL FILL_39_DFFSR_146 ( );
FILL FILL_40_DFFSR_146 ( );
FILL FILL_41_DFFSR_146 ( );
FILL FILL_42_DFFSR_146 ( );
FILL FILL_43_DFFSR_146 ( );
FILL FILL_44_DFFSR_146 ( );
FILL FILL_45_DFFSR_146 ( );
FILL FILL_46_DFFSR_146 ( );
FILL FILL_47_DFFSR_146 ( );
FILL FILL_48_DFFSR_146 ( );
FILL FILL_49_DFFSR_146 ( );
FILL FILL_50_DFFSR_146 ( );
FILL FILL_0_INVX1_166 ( );
FILL FILL_1_INVX1_166 ( );
FILL FILL_2_INVX1_166 ( );
FILL FILL_3_INVX1_166 ( );
FILL FILL_4_INVX1_166 ( );
FILL FILL_0_NAND2X1_147 ( );
FILL FILL_1_NAND2X1_147 ( );
FILL FILL_2_NAND2X1_147 ( );
FILL FILL_3_NAND2X1_147 ( );
FILL FILL_4_NAND2X1_147 ( );
FILL FILL_5_NAND2X1_147 ( );
FILL FILL_6_NAND2X1_147 ( );
FILL FILL_0_NAND2X1_262 ( );
FILL FILL_1_NAND2X1_262 ( );
FILL FILL_2_NAND2X1_262 ( );
FILL FILL_3_NAND2X1_262 ( );
FILL FILL_4_NAND2X1_262 ( );
FILL FILL_5_NAND2X1_262 ( );
FILL FILL_6_NAND2X1_262 ( );
FILL FILL_0_INVX1_413 ( );
FILL FILL_1_INVX1_413 ( );
FILL FILL_2_INVX1_413 ( );
FILL FILL_3_INVX1_413 ( );
FILL FILL_0_OAI21X1_251 ( );
FILL FILL_1_OAI21X1_251 ( );
FILL FILL_2_OAI21X1_251 ( );
FILL FILL_3_OAI21X1_251 ( );
FILL FILL_4_OAI21X1_251 ( );
FILL FILL_5_OAI21X1_251 ( );
FILL FILL_6_OAI21X1_251 ( );
FILL FILL_7_OAI21X1_251 ( );
FILL FILL_8_OAI21X1_251 ( );
FILL FILL_9_OAI21X1_251 ( );
FILL FILL_0_DFFSR_20 ( );
FILL FILL_1_DFFSR_20 ( );
FILL FILL_2_DFFSR_20 ( );
FILL FILL_3_DFFSR_20 ( );
FILL FILL_4_DFFSR_20 ( );
FILL FILL_5_DFFSR_20 ( );
FILL FILL_6_DFFSR_20 ( );
FILL FILL_7_DFFSR_20 ( );
FILL FILL_8_DFFSR_20 ( );
FILL FILL_9_DFFSR_20 ( );
FILL FILL_10_DFFSR_20 ( );
FILL FILL_11_DFFSR_20 ( );
FILL FILL_12_DFFSR_20 ( );
FILL FILL_13_DFFSR_20 ( );
FILL FILL_14_DFFSR_20 ( );
FILL FILL_15_DFFSR_20 ( );
FILL FILL_16_DFFSR_20 ( );
FILL FILL_17_DFFSR_20 ( );
FILL FILL_18_DFFSR_20 ( );
FILL FILL_19_DFFSR_20 ( );
FILL FILL_20_DFFSR_20 ( );
FILL FILL_21_DFFSR_20 ( );
FILL FILL_22_DFFSR_20 ( );
FILL FILL_23_DFFSR_20 ( );
FILL FILL_24_DFFSR_20 ( );
FILL FILL_25_DFFSR_20 ( );
FILL FILL_26_DFFSR_20 ( );
FILL FILL_27_DFFSR_20 ( );
FILL FILL_28_DFFSR_20 ( );
FILL FILL_29_DFFSR_20 ( );
FILL FILL_30_DFFSR_20 ( );
FILL FILL_31_DFFSR_20 ( );
FILL FILL_32_DFFSR_20 ( );
FILL FILL_33_DFFSR_20 ( );
FILL FILL_34_DFFSR_20 ( );
FILL FILL_35_DFFSR_20 ( );
FILL FILL_36_DFFSR_20 ( );
FILL FILL_37_DFFSR_20 ( );
FILL FILL_38_DFFSR_20 ( );
FILL FILL_39_DFFSR_20 ( );
FILL FILL_40_DFFSR_20 ( );
FILL FILL_41_DFFSR_20 ( );
FILL FILL_42_DFFSR_20 ( );
FILL FILL_43_DFFSR_20 ( );
FILL FILL_44_DFFSR_20 ( );
FILL FILL_45_DFFSR_20 ( );
FILL FILL_46_DFFSR_20 ( );
FILL FILL_47_DFFSR_20 ( );
FILL FILL_48_DFFSR_20 ( );
FILL FILL_49_DFFSR_20 ( );
FILL FILL_50_DFFSR_20 ( );
FILL FILL_0_DFFSR_162 ( );
FILL FILL_1_DFFSR_162 ( );
FILL FILL_2_DFFSR_162 ( );
FILL FILL_3_DFFSR_162 ( );
FILL FILL_4_DFFSR_162 ( );
FILL FILL_5_DFFSR_162 ( );
FILL FILL_6_DFFSR_162 ( );
FILL FILL_7_DFFSR_162 ( );
FILL FILL_8_DFFSR_162 ( );
FILL FILL_9_DFFSR_162 ( );
FILL FILL_10_DFFSR_162 ( );
FILL FILL_11_DFFSR_162 ( );
FILL FILL_12_DFFSR_162 ( );
FILL FILL_13_DFFSR_162 ( );
FILL FILL_14_DFFSR_162 ( );
FILL FILL_15_DFFSR_162 ( );
FILL FILL_16_DFFSR_162 ( );
FILL FILL_17_DFFSR_162 ( );
FILL FILL_18_DFFSR_162 ( );
FILL FILL_19_DFFSR_162 ( );
FILL FILL_20_DFFSR_162 ( );
FILL FILL_21_DFFSR_162 ( );
FILL FILL_22_DFFSR_162 ( );
FILL FILL_23_DFFSR_162 ( );
FILL FILL_24_DFFSR_162 ( );
FILL FILL_25_DFFSR_162 ( );
FILL FILL_26_DFFSR_162 ( );
FILL FILL_27_DFFSR_162 ( );
FILL FILL_28_DFFSR_162 ( );
FILL FILL_29_DFFSR_162 ( );
FILL FILL_30_DFFSR_162 ( );
FILL FILL_31_DFFSR_162 ( );
FILL FILL_32_DFFSR_162 ( );
FILL FILL_33_DFFSR_162 ( );
FILL FILL_34_DFFSR_162 ( );
FILL FILL_35_DFFSR_162 ( );
FILL FILL_36_DFFSR_162 ( );
FILL FILL_37_DFFSR_162 ( );
FILL FILL_38_DFFSR_162 ( );
FILL FILL_39_DFFSR_162 ( );
FILL FILL_40_DFFSR_162 ( );
FILL FILL_41_DFFSR_162 ( );
FILL FILL_42_DFFSR_162 ( );
FILL FILL_43_DFFSR_162 ( );
FILL FILL_44_DFFSR_162 ( );
FILL FILL_45_DFFSR_162 ( );
FILL FILL_46_DFFSR_162 ( );
FILL FILL_47_DFFSR_162 ( );
FILL FILL_48_DFFSR_162 ( );
FILL FILL_49_DFFSR_162 ( );
FILL FILL_50_DFFSR_162 ( );
FILL FILL_0_INVX1_246 ( );
FILL FILL_1_INVX1_246 ( );
FILL FILL_2_INVX1_246 ( );
FILL FILL_3_INVX1_246 ( );
FILL FILL_4_INVX1_246 ( );
FILL FILL_0_OAI21X1_222 ( );
FILL FILL_1_OAI21X1_222 ( );
FILL FILL_2_OAI21X1_222 ( );
FILL FILL_3_OAI21X1_222 ( );
FILL FILL_4_OAI21X1_222 ( );
FILL FILL_5_OAI21X1_222 ( );
FILL FILL_6_OAI21X1_222 ( );
FILL FILL_7_OAI21X1_222 ( );
FILL FILL_8_OAI21X1_222 ( );
FILL FILL_0_NOR2X1_7 ( );
FILL FILL_1_NOR2X1_7 ( );
FILL FILL_2_NOR2X1_7 ( );
FILL FILL_3_NOR2X1_7 ( );
FILL FILL_4_NOR2X1_7 ( );
FILL FILL_5_NOR2X1_7 ( );
FILL FILL_6_NOR2X1_7 ( );
FILL FILL_0_DFFSR_185 ( );
FILL FILL_1_DFFSR_185 ( );
FILL FILL_2_DFFSR_185 ( );
FILL FILL_3_DFFSR_185 ( );
FILL FILL_4_DFFSR_185 ( );
FILL FILL_5_DFFSR_185 ( );
FILL FILL_6_DFFSR_185 ( );
FILL FILL_7_DFFSR_185 ( );
FILL FILL_8_DFFSR_185 ( );
FILL FILL_9_DFFSR_185 ( );
FILL FILL_10_DFFSR_185 ( );
FILL FILL_11_DFFSR_185 ( );
FILL FILL_12_DFFSR_185 ( );
FILL FILL_13_DFFSR_185 ( );
FILL FILL_14_DFFSR_185 ( );
FILL FILL_15_DFFSR_185 ( );
FILL FILL_16_DFFSR_185 ( );
FILL FILL_17_DFFSR_185 ( );
FILL FILL_18_DFFSR_185 ( );
FILL FILL_19_DFFSR_185 ( );
FILL FILL_20_DFFSR_185 ( );
FILL FILL_21_DFFSR_185 ( );
FILL FILL_22_DFFSR_185 ( );
FILL FILL_23_DFFSR_185 ( );
FILL FILL_24_DFFSR_185 ( );
FILL FILL_25_DFFSR_185 ( );
FILL FILL_26_DFFSR_185 ( );
FILL FILL_27_DFFSR_185 ( );
FILL FILL_28_DFFSR_185 ( );
FILL FILL_29_DFFSR_185 ( );
FILL FILL_30_DFFSR_185 ( );
FILL FILL_31_DFFSR_185 ( );
FILL FILL_32_DFFSR_185 ( );
FILL FILL_33_DFFSR_185 ( );
FILL FILL_34_DFFSR_185 ( );
FILL FILL_35_DFFSR_185 ( );
FILL FILL_36_DFFSR_185 ( );
FILL FILL_37_DFFSR_185 ( );
FILL FILL_38_DFFSR_185 ( );
FILL FILL_39_DFFSR_185 ( );
FILL FILL_40_DFFSR_185 ( );
FILL FILL_41_DFFSR_185 ( );
FILL FILL_42_DFFSR_185 ( );
FILL FILL_43_DFFSR_185 ( );
FILL FILL_44_DFFSR_185 ( );
FILL FILL_45_DFFSR_185 ( );
FILL FILL_46_DFFSR_185 ( );
FILL FILL_47_DFFSR_185 ( );
FILL FILL_48_DFFSR_185 ( );
FILL FILL_49_DFFSR_185 ( );
FILL FILL_50_DFFSR_185 ( );
FILL FILL_0_OAI21X1_253 ( );
FILL FILL_1_OAI21X1_253 ( );
FILL FILL_2_OAI21X1_253 ( );
FILL FILL_3_OAI21X1_253 ( );
FILL FILL_4_OAI21X1_253 ( );
FILL FILL_5_OAI21X1_253 ( );
FILL FILL_6_OAI21X1_253 ( );
FILL FILL_7_OAI21X1_253 ( );
FILL FILL_8_OAI21X1_253 ( );
FILL FILL_0_INVX1_416 ( );
FILL FILL_1_INVX1_416 ( );
FILL FILL_2_INVX1_416 ( );
FILL FILL_3_INVX1_416 ( );
FILL FILL_4_INVX1_416 ( );
FILL FILL_0_DFFSR_105 ( );
FILL FILL_1_DFFSR_105 ( );
FILL FILL_2_DFFSR_105 ( );
FILL FILL_3_DFFSR_105 ( );
FILL FILL_4_DFFSR_105 ( );
FILL FILL_5_DFFSR_105 ( );
FILL FILL_6_DFFSR_105 ( );
FILL FILL_7_DFFSR_105 ( );
FILL FILL_8_DFFSR_105 ( );
FILL FILL_9_DFFSR_105 ( );
FILL FILL_10_DFFSR_105 ( );
FILL FILL_11_DFFSR_105 ( );
FILL FILL_12_DFFSR_105 ( );
FILL FILL_13_DFFSR_105 ( );
FILL FILL_14_DFFSR_105 ( );
FILL FILL_15_DFFSR_105 ( );
FILL FILL_16_DFFSR_105 ( );
FILL FILL_17_DFFSR_105 ( );
FILL FILL_18_DFFSR_105 ( );
FILL FILL_19_DFFSR_105 ( );
FILL FILL_20_DFFSR_105 ( );
FILL FILL_21_DFFSR_105 ( );
FILL FILL_22_DFFSR_105 ( );
FILL FILL_23_DFFSR_105 ( );
FILL FILL_24_DFFSR_105 ( );
FILL FILL_25_DFFSR_105 ( );
FILL FILL_26_DFFSR_105 ( );
FILL FILL_27_DFFSR_105 ( );
FILL FILL_28_DFFSR_105 ( );
FILL FILL_29_DFFSR_105 ( );
FILL FILL_30_DFFSR_105 ( );
FILL FILL_31_DFFSR_105 ( );
FILL FILL_32_DFFSR_105 ( );
FILL FILL_33_DFFSR_105 ( );
FILL FILL_34_DFFSR_105 ( );
FILL FILL_35_DFFSR_105 ( );
FILL FILL_36_DFFSR_105 ( );
FILL FILL_37_DFFSR_105 ( );
FILL FILL_38_DFFSR_105 ( );
FILL FILL_39_DFFSR_105 ( );
FILL FILL_40_DFFSR_105 ( );
FILL FILL_41_DFFSR_105 ( );
FILL FILL_42_DFFSR_105 ( );
FILL FILL_43_DFFSR_105 ( );
FILL FILL_44_DFFSR_105 ( );
FILL FILL_45_DFFSR_105 ( );
FILL FILL_46_DFFSR_105 ( );
FILL FILL_47_DFFSR_105 ( );
FILL FILL_48_DFFSR_105 ( );
FILL FILL_49_DFFSR_105 ( );
FILL FILL_50_DFFSR_105 ( );
FILL FILL_0_DFFSR_123 ( );
FILL FILL_1_DFFSR_123 ( );
FILL FILL_2_DFFSR_123 ( );
FILL FILL_3_DFFSR_123 ( );
FILL FILL_4_DFFSR_123 ( );
FILL FILL_5_DFFSR_123 ( );
FILL FILL_6_DFFSR_123 ( );
FILL FILL_7_DFFSR_123 ( );
FILL FILL_8_DFFSR_123 ( );
FILL FILL_9_DFFSR_123 ( );
FILL FILL_10_DFFSR_123 ( );
FILL FILL_11_DFFSR_123 ( );
FILL FILL_12_DFFSR_123 ( );
FILL FILL_13_DFFSR_123 ( );
FILL FILL_14_DFFSR_123 ( );
FILL FILL_15_DFFSR_123 ( );
FILL FILL_16_DFFSR_123 ( );
FILL FILL_17_DFFSR_123 ( );
FILL FILL_18_DFFSR_123 ( );
FILL FILL_19_DFFSR_123 ( );
FILL FILL_20_DFFSR_123 ( );
FILL FILL_21_DFFSR_123 ( );
FILL FILL_22_DFFSR_123 ( );
FILL FILL_23_DFFSR_123 ( );
FILL FILL_24_DFFSR_123 ( );
FILL FILL_25_DFFSR_123 ( );
FILL FILL_26_DFFSR_123 ( );
FILL FILL_27_DFFSR_123 ( );
FILL FILL_28_DFFSR_123 ( );
FILL FILL_29_DFFSR_123 ( );
FILL FILL_30_DFFSR_123 ( );
FILL FILL_31_DFFSR_123 ( );
FILL FILL_32_DFFSR_123 ( );
FILL FILL_33_DFFSR_123 ( );
FILL FILL_34_DFFSR_123 ( );
FILL FILL_35_DFFSR_123 ( );
FILL FILL_36_DFFSR_123 ( );
FILL FILL_37_DFFSR_123 ( );
FILL FILL_38_DFFSR_123 ( );
FILL FILL_39_DFFSR_123 ( );
FILL FILL_40_DFFSR_123 ( );
FILL FILL_41_DFFSR_123 ( );
FILL FILL_42_DFFSR_123 ( );
FILL FILL_43_DFFSR_123 ( );
FILL FILL_44_DFFSR_123 ( );
FILL FILL_45_DFFSR_123 ( );
FILL FILL_46_DFFSR_123 ( );
FILL FILL_47_DFFSR_123 ( );
FILL FILL_48_DFFSR_123 ( );
FILL FILL_49_DFFSR_123 ( );
FILL FILL_50_DFFSR_123 ( );
FILL FILL_0_INVX1_172 ( );
FILL FILL_1_INVX1_172 ( );
FILL FILL_2_INVX1_172 ( );
FILL FILL_3_INVX1_172 ( );
FILL FILL_4_INVX1_172 ( );
FILL FILL_0_OAI21X1_149 ( );
FILL FILL_1_OAI21X1_149 ( );
FILL FILL_2_OAI21X1_149 ( );
FILL FILL_3_OAI21X1_149 ( );
FILL FILL_4_OAI21X1_149 ( );
FILL FILL_5_OAI21X1_149 ( );
FILL FILL_6_OAI21X1_149 ( );
FILL FILL_7_OAI21X1_149 ( );
FILL FILL_8_OAI21X1_149 ( );
FILL FILL_0_NAND2X1_149 ( );
FILL FILL_1_NAND2X1_149 ( );
FILL FILL_2_NAND2X1_149 ( );
FILL FILL_3_NAND2X1_149 ( );
FILL FILL_4_NAND2X1_149 ( );
FILL FILL_5_NAND2X1_149 ( );
FILL FILL_6_NAND2X1_149 ( );
FILL FILL_0_OAI21X1_148 ( );
FILL FILL_1_OAI21X1_148 ( );
FILL FILL_2_OAI21X1_148 ( );
FILL FILL_3_OAI21X1_148 ( );
FILL FILL_4_OAI21X1_148 ( );
FILL FILL_5_OAI21X1_148 ( );
FILL FILL_6_OAI21X1_148 ( );
FILL FILL_7_OAI21X1_148 ( );
FILL FILL_8_OAI21X1_148 ( );
FILL FILL_0_OAI21X1_249 ( );
FILL FILL_1_OAI21X1_249 ( );
FILL FILL_2_OAI21X1_249 ( );
FILL FILL_3_OAI21X1_249 ( );
FILL FILL_4_OAI21X1_249 ( );
FILL FILL_5_OAI21X1_249 ( );
FILL FILL_6_OAI21X1_249 ( );
FILL FILL_7_OAI21X1_249 ( );
FILL FILL_8_OAI21X1_249 ( );
FILL FILL_9_OAI21X1_249 ( );
FILL FILL_0_NAND2X1_260 ( );
FILL FILL_1_NAND2X1_260 ( );
FILL FILL_2_NAND2X1_260 ( );
FILL FILL_3_NAND2X1_260 ( );
FILL FILL_4_NAND2X1_260 ( );
FILL FILL_5_NAND2X1_260 ( );
FILL FILL_6_NAND2X1_260 ( );
FILL FILL_0_INVX1_411 ( );
FILL FILL_1_INVX1_411 ( );
FILL FILL_2_INVX1_411 ( );
FILL FILL_3_INVX1_411 ( );
FILL FILL_0_DFFSR_147 ( );
FILL FILL_1_DFFSR_147 ( );
FILL FILL_2_DFFSR_147 ( );
FILL FILL_3_DFFSR_147 ( );
FILL FILL_4_DFFSR_147 ( );
FILL FILL_5_DFFSR_147 ( );
FILL FILL_6_DFFSR_147 ( );
FILL FILL_7_DFFSR_147 ( );
FILL FILL_8_DFFSR_147 ( );
FILL FILL_9_DFFSR_147 ( );
FILL FILL_10_DFFSR_147 ( );
FILL FILL_11_DFFSR_147 ( );
FILL FILL_12_DFFSR_147 ( );
FILL FILL_13_DFFSR_147 ( );
FILL FILL_14_DFFSR_147 ( );
FILL FILL_15_DFFSR_147 ( );
FILL FILL_16_DFFSR_147 ( );
FILL FILL_17_DFFSR_147 ( );
FILL FILL_18_DFFSR_147 ( );
FILL FILL_19_DFFSR_147 ( );
FILL FILL_20_DFFSR_147 ( );
FILL FILL_21_DFFSR_147 ( );
FILL FILL_22_DFFSR_147 ( );
FILL FILL_23_DFFSR_147 ( );
FILL FILL_24_DFFSR_147 ( );
FILL FILL_25_DFFSR_147 ( );
FILL FILL_26_DFFSR_147 ( );
FILL FILL_27_DFFSR_147 ( );
FILL FILL_28_DFFSR_147 ( );
FILL FILL_29_DFFSR_147 ( );
FILL FILL_30_DFFSR_147 ( );
FILL FILL_31_DFFSR_147 ( );
FILL FILL_32_DFFSR_147 ( );
FILL FILL_33_DFFSR_147 ( );
FILL FILL_34_DFFSR_147 ( );
FILL FILL_35_DFFSR_147 ( );
FILL FILL_36_DFFSR_147 ( );
FILL FILL_37_DFFSR_147 ( );
FILL FILL_38_DFFSR_147 ( );
FILL FILL_39_DFFSR_147 ( );
FILL FILL_40_DFFSR_147 ( );
FILL FILL_41_DFFSR_147 ( );
FILL FILL_42_DFFSR_147 ( );
FILL FILL_43_DFFSR_147 ( );
FILL FILL_44_DFFSR_147 ( );
FILL FILL_45_DFFSR_147 ( );
FILL FILL_46_DFFSR_147 ( );
FILL FILL_47_DFFSR_147 ( );
FILL FILL_48_DFFSR_147 ( );
FILL FILL_49_DFFSR_147 ( );
FILL FILL_50_DFFSR_147 ( );
FILL FILL_0_INVX1_169 ( );
FILL FILL_1_INVX1_169 ( );
FILL FILL_2_INVX1_169 ( );
FILL FILL_3_INVX1_169 ( );
FILL FILL_4_INVX1_169 ( );
FILL FILL_0_OAI21X1_147 ( );
FILL FILL_1_OAI21X1_147 ( );
FILL FILL_2_OAI21X1_147 ( );
FILL FILL_3_OAI21X1_147 ( );
FILL FILL_4_OAI21X1_147 ( );
FILL FILL_5_OAI21X1_147 ( );
FILL FILL_6_OAI21X1_147 ( );
FILL FILL_7_OAI21X1_147 ( );
FILL FILL_8_OAI21X1_147 ( );
FILL FILL_0_OAI21X1_146 ( );
FILL FILL_1_OAI21X1_146 ( );
FILL FILL_2_OAI21X1_146 ( );
FILL FILL_3_OAI21X1_146 ( );
FILL FILL_4_OAI21X1_146 ( );
FILL FILL_5_OAI21X1_146 ( );
FILL FILL_6_OAI21X1_146 ( );
FILL FILL_7_OAI21X1_146 ( );
FILL FILL_8_OAI21X1_146 ( );
FILL FILL_0_DFFSR_183 ( );
FILL FILL_1_DFFSR_183 ( );
FILL FILL_2_DFFSR_183 ( );
FILL FILL_3_DFFSR_183 ( );
FILL FILL_4_DFFSR_183 ( );
FILL FILL_5_DFFSR_183 ( );
FILL FILL_6_DFFSR_183 ( );
FILL FILL_7_DFFSR_183 ( );
FILL FILL_8_DFFSR_183 ( );
FILL FILL_9_DFFSR_183 ( );
FILL FILL_10_DFFSR_183 ( );
FILL FILL_11_DFFSR_183 ( );
FILL FILL_12_DFFSR_183 ( );
FILL FILL_13_DFFSR_183 ( );
FILL FILL_14_DFFSR_183 ( );
FILL FILL_15_DFFSR_183 ( );
FILL FILL_16_DFFSR_183 ( );
FILL FILL_17_DFFSR_183 ( );
FILL FILL_18_DFFSR_183 ( );
FILL FILL_19_DFFSR_183 ( );
FILL FILL_20_DFFSR_183 ( );
FILL FILL_21_DFFSR_183 ( );
FILL FILL_22_DFFSR_183 ( );
FILL FILL_23_DFFSR_183 ( );
FILL FILL_24_DFFSR_183 ( );
FILL FILL_25_DFFSR_183 ( );
FILL FILL_26_DFFSR_183 ( );
FILL FILL_27_DFFSR_183 ( );
FILL FILL_28_DFFSR_183 ( );
FILL FILL_29_DFFSR_183 ( );
FILL FILL_30_DFFSR_183 ( );
FILL FILL_31_DFFSR_183 ( );
FILL FILL_32_DFFSR_183 ( );
FILL FILL_33_DFFSR_183 ( );
FILL FILL_34_DFFSR_183 ( );
FILL FILL_35_DFFSR_183 ( );
FILL FILL_36_DFFSR_183 ( );
FILL FILL_37_DFFSR_183 ( );
FILL FILL_38_DFFSR_183 ( );
FILL FILL_39_DFFSR_183 ( );
FILL FILL_40_DFFSR_183 ( );
FILL FILL_41_DFFSR_183 ( );
FILL FILL_42_DFFSR_183 ( );
FILL FILL_43_DFFSR_183 ( );
FILL FILL_44_DFFSR_183 ( );
FILL FILL_45_DFFSR_183 ( );
FILL FILL_46_DFFSR_183 ( );
FILL FILL_47_DFFSR_183 ( );
FILL FILL_48_DFFSR_183 ( );
FILL FILL_49_DFFSR_183 ( );
FILL FILL_50_DFFSR_183 ( );
FILL FILL_0_OAI21X1_20 ( );
FILL FILL_1_OAI21X1_20 ( );
FILL FILL_2_OAI21X1_20 ( );
FILL FILL_3_OAI21X1_20 ( );
FILL FILL_4_OAI21X1_20 ( );
FILL FILL_5_OAI21X1_20 ( );
FILL FILL_6_OAI21X1_20 ( );
FILL FILL_7_OAI21X1_20 ( );
FILL FILL_8_OAI21X1_20 ( );
FILL FILL_0_XOR2X1_5 ( );
FILL FILL_1_XOR2X1_5 ( );
FILL FILL_2_XOR2X1_5 ( );
FILL FILL_3_XOR2X1_5 ( );
FILL FILL_4_XOR2X1_5 ( );
FILL FILL_5_XOR2X1_5 ( );
FILL FILL_6_XOR2X1_5 ( );
FILL FILL_7_XOR2X1_5 ( );
FILL FILL_8_XOR2X1_5 ( );
FILL FILL_9_XOR2X1_5 ( );
FILL FILL_10_XOR2X1_5 ( );
FILL FILL_11_XOR2X1_5 ( );
FILL FILL_12_XOR2X1_5 ( );
FILL FILL_13_XOR2X1_5 ( );
FILL FILL_14_XOR2X1_5 ( );
FILL FILL_15_XOR2X1_5 ( );
FILL FILL_0_BUFX2_28 ( );
FILL FILL_1_BUFX2_28 ( );
FILL FILL_2_BUFX2_28 ( );
FILL FILL_3_BUFX2_28 ( );
FILL FILL_4_BUFX2_28 ( );
FILL FILL_5_BUFX2_28 ( );
FILL FILL_6_BUFX2_28 ( );
FILL FILL_0_XOR2X1_4 ( );
FILL FILL_1_XOR2X1_4 ( );
FILL FILL_2_XOR2X1_4 ( );
FILL FILL_3_XOR2X1_4 ( );
FILL FILL_4_XOR2X1_4 ( );
FILL FILL_5_XOR2X1_4 ( );
FILL FILL_6_XOR2X1_4 ( );
FILL FILL_7_XOR2X1_4 ( );
FILL FILL_8_XOR2X1_4 ( );
FILL FILL_9_XOR2X1_4 ( );
FILL FILL_10_XOR2X1_4 ( );
FILL FILL_11_XOR2X1_4 ( );
FILL FILL_12_XOR2X1_4 ( );
FILL FILL_13_XOR2X1_4 ( );
FILL FILL_14_XOR2X1_4 ( );
FILL FILL_15_XOR2X1_4 ( );
FILL FILL_0_NAND2X1_265 ( );
FILL FILL_1_NAND2X1_265 ( );
FILL FILL_2_NAND2X1_265 ( );
FILL FILL_3_NAND2X1_265 ( );
FILL FILL_4_NAND2X1_265 ( );
FILL FILL_5_NAND2X1_265 ( );
FILL FILL_6_NAND2X1_265 ( );
FILL FILL_0_INVX1_196 ( );
FILL FILL_1_INVX1_196 ( );
FILL FILL_2_INVX1_196 ( );
FILL FILL_3_INVX1_196 ( );
FILL FILL_4_INVX1_196 ( );
FILL FILL_0_XOR2X1_6 ( );
FILL FILL_1_XOR2X1_6 ( );
FILL FILL_2_XOR2X1_6 ( );
FILL FILL_3_XOR2X1_6 ( );
FILL FILL_4_XOR2X1_6 ( );
FILL FILL_5_XOR2X1_6 ( );
FILL FILL_6_XOR2X1_6 ( );
FILL FILL_7_XOR2X1_6 ( );
FILL FILL_8_XOR2X1_6 ( );
FILL FILL_9_XOR2X1_6 ( );
FILL FILL_10_XOR2X1_6 ( );
FILL FILL_11_XOR2X1_6 ( );
FILL FILL_12_XOR2X1_6 ( );
FILL FILL_13_XOR2X1_6 ( );
FILL FILL_14_XOR2X1_6 ( );
FILL FILL_15_XOR2X1_6 ( );
FILL FILL_0_DFFSR_161 ( );
FILL FILL_1_DFFSR_161 ( );
FILL FILL_2_DFFSR_161 ( );
FILL FILL_3_DFFSR_161 ( );
FILL FILL_4_DFFSR_161 ( );
FILL FILL_5_DFFSR_161 ( );
FILL FILL_6_DFFSR_161 ( );
FILL FILL_7_DFFSR_161 ( );
FILL FILL_8_DFFSR_161 ( );
FILL FILL_9_DFFSR_161 ( );
FILL FILL_10_DFFSR_161 ( );
FILL FILL_11_DFFSR_161 ( );
FILL FILL_12_DFFSR_161 ( );
FILL FILL_13_DFFSR_161 ( );
FILL FILL_14_DFFSR_161 ( );
FILL FILL_15_DFFSR_161 ( );
FILL FILL_16_DFFSR_161 ( );
FILL FILL_17_DFFSR_161 ( );
FILL FILL_18_DFFSR_161 ( );
FILL FILL_19_DFFSR_161 ( );
FILL FILL_20_DFFSR_161 ( );
FILL FILL_21_DFFSR_161 ( );
FILL FILL_22_DFFSR_161 ( );
FILL FILL_23_DFFSR_161 ( );
FILL FILL_24_DFFSR_161 ( );
FILL FILL_25_DFFSR_161 ( );
FILL FILL_26_DFFSR_161 ( );
FILL FILL_27_DFFSR_161 ( );
FILL FILL_28_DFFSR_161 ( );
FILL FILL_29_DFFSR_161 ( );
FILL FILL_30_DFFSR_161 ( );
FILL FILL_31_DFFSR_161 ( );
FILL FILL_32_DFFSR_161 ( );
FILL FILL_33_DFFSR_161 ( );
FILL FILL_34_DFFSR_161 ( );
FILL FILL_35_DFFSR_161 ( );
FILL FILL_36_DFFSR_161 ( );
FILL FILL_37_DFFSR_161 ( );
FILL FILL_38_DFFSR_161 ( );
FILL FILL_39_DFFSR_161 ( );
FILL FILL_40_DFFSR_161 ( );
FILL FILL_41_DFFSR_161 ( );
FILL FILL_42_DFFSR_161 ( );
FILL FILL_43_DFFSR_161 ( );
FILL FILL_44_DFFSR_161 ( );
FILL FILL_45_DFFSR_161 ( );
FILL FILL_46_DFFSR_161 ( );
FILL FILL_47_DFFSR_161 ( );
FILL FILL_48_DFFSR_161 ( );
FILL FILL_49_DFFSR_161 ( );
FILL FILL_50_DFFSR_161 ( );
FILL FILL_51_DFFSR_161 ( );
FILL FILL_0_BUFX2_33 ( );
FILL FILL_1_BUFX2_33 ( );
FILL FILL_2_BUFX2_33 ( );
FILL FILL_3_BUFX2_33 ( );
FILL FILL_4_BUFX2_33 ( );
FILL FILL_5_BUFX2_33 ( );
FILL FILL_6_BUFX2_33 ( );
FILL FILL_0_NAND3X1_101 ( );
FILL FILL_1_NAND3X1_101 ( );
FILL FILL_2_NAND3X1_101 ( );
FILL FILL_3_NAND3X1_101 ( );
FILL FILL_4_NAND3X1_101 ( );
FILL FILL_5_NAND3X1_101 ( );
FILL FILL_6_NAND3X1_101 ( );
FILL FILL_7_NAND3X1_101 ( );
FILL FILL_8_NAND3X1_101 ( );
FILL FILL_9_NAND3X1_101 ( );
FILL FILL_0_NAND2X1_264 ( );
FILL FILL_1_NAND2X1_264 ( );
FILL FILL_2_NAND2X1_264 ( );
FILL FILL_3_NAND2X1_264 ( );
FILL FILL_4_NAND2X1_264 ( );
FILL FILL_5_NAND2X1_264 ( );
FILL FILL_6_NAND2X1_264 ( );
FILL FILL_0_BUFX2_27 ( );
FILL FILL_1_BUFX2_27 ( );
FILL FILL_2_BUFX2_27 ( );
FILL FILL_3_BUFX2_27 ( );
FILL FILL_4_BUFX2_27 ( );
FILL FILL_5_BUFX2_27 ( );
FILL FILL_6_BUFX2_27 ( );
FILL FILL_0_INVX1_260 ( );
FILL FILL_1_INVX1_260 ( );
FILL FILL_2_INVX1_260 ( );
FILL FILL_3_INVX1_260 ( );
FILL FILL_0_DFFSR_113 ( );
FILL FILL_1_DFFSR_113 ( );
FILL FILL_2_DFFSR_113 ( );
FILL FILL_3_DFFSR_113 ( );
FILL FILL_4_DFFSR_113 ( );
FILL FILL_5_DFFSR_113 ( );
FILL FILL_6_DFFSR_113 ( );
FILL FILL_7_DFFSR_113 ( );
FILL FILL_8_DFFSR_113 ( );
FILL FILL_9_DFFSR_113 ( );
FILL FILL_10_DFFSR_113 ( );
FILL FILL_11_DFFSR_113 ( );
FILL FILL_12_DFFSR_113 ( );
FILL FILL_13_DFFSR_113 ( );
FILL FILL_14_DFFSR_113 ( );
FILL FILL_15_DFFSR_113 ( );
FILL FILL_16_DFFSR_113 ( );
FILL FILL_17_DFFSR_113 ( );
FILL FILL_18_DFFSR_113 ( );
FILL FILL_19_DFFSR_113 ( );
FILL FILL_20_DFFSR_113 ( );
FILL FILL_21_DFFSR_113 ( );
FILL FILL_22_DFFSR_113 ( );
FILL FILL_23_DFFSR_113 ( );
FILL FILL_24_DFFSR_113 ( );
FILL FILL_25_DFFSR_113 ( );
FILL FILL_26_DFFSR_113 ( );
FILL FILL_27_DFFSR_113 ( );
FILL FILL_28_DFFSR_113 ( );
FILL FILL_29_DFFSR_113 ( );
FILL FILL_30_DFFSR_113 ( );
FILL FILL_31_DFFSR_113 ( );
FILL FILL_32_DFFSR_113 ( );
FILL FILL_33_DFFSR_113 ( );
FILL FILL_34_DFFSR_113 ( );
FILL FILL_35_DFFSR_113 ( );
FILL FILL_36_DFFSR_113 ( );
FILL FILL_37_DFFSR_113 ( );
FILL FILL_38_DFFSR_113 ( );
FILL FILL_39_DFFSR_113 ( );
FILL FILL_40_DFFSR_113 ( );
FILL FILL_41_DFFSR_113 ( );
FILL FILL_42_DFFSR_113 ( );
FILL FILL_43_DFFSR_113 ( );
FILL FILL_44_DFFSR_113 ( );
FILL FILL_45_DFFSR_113 ( );
FILL FILL_46_DFFSR_113 ( );
FILL FILL_47_DFFSR_113 ( );
FILL FILL_48_DFFSR_113 ( );
FILL FILL_49_DFFSR_113 ( );
FILL FILL_50_DFFSR_113 ( );
FILL FILL_0_DFFSR_100 ( );
FILL FILL_1_DFFSR_100 ( );
FILL FILL_2_DFFSR_100 ( );
FILL FILL_3_DFFSR_100 ( );
FILL FILL_4_DFFSR_100 ( );
FILL FILL_5_DFFSR_100 ( );
FILL FILL_6_DFFSR_100 ( );
FILL FILL_7_DFFSR_100 ( );
FILL FILL_8_DFFSR_100 ( );
FILL FILL_9_DFFSR_100 ( );
FILL FILL_10_DFFSR_100 ( );
FILL FILL_11_DFFSR_100 ( );
FILL FILL_12_DFFSR_100 ( );
FILL FILL_13_DFFSR_100 ( );
FILL FILL_14_DFFSR_100 ( );
FILL FILL_15_DFFSR_100 ( );
FILL FILL_16_DFFSR_100 ( );
FILL FILL_17_DFFSR_100 ( );
FILL FILL_18_DFFSR_100 ( );
FILL FILL_19_DFFSR_100 ( );
FILL FILL_20_DFFSR_100 ( );
FILL FILL_21_DFFSR_100 ( );
FILL FILL_22_DFFSR_100 ( );
FILL FILL_23_DFFSR_100 ( );
FILL FILL_24_DFFSR_100 ( );
FILL FILL_25_DFFSR_100 ( );
FILL FILL_26_DFFSR_100 ( );
FILL FILL_27_DFFSR_100 ( );
FILL FILL_28_DFFSR_100 ( );
FILL FILL_29_DFFSR_100 ( );
FILL FILL_30_DFFSR_100 ( );
FILL FILL_31_DFFSR_100 ( );
FILL FILL_32_DFFSR_100 ( );
FILL FILL_33_DFFSR_100 ( );
FILL FILL_34_DFFSR_100 ( );
FILL FILL_35_DFFSR_100 ( );
FILL FILL_36_DFFSR_100 ( );
FILL FILL_37_DFFSR_100 ( );
FILL FILL_38_DFFSR_100 ( );
FILL FILL_39_DFFSR_100 ( );
FILL FILL_40_DFFSR_100 ( );
FILL FILL_41_DFFSR_100 ( );
FILL FILL_42_DFFSR_100 ( );
FILL FILL_43_DFFSR_100 ( );
FILL FILL_44_DFFSR_100 ( );
FILL FILL_45_DFFSR_100 ( );
FILL FILL_46_DFFSR_100 ( );
FILL FILL_47_DFFSR_100 ( );
FILL FILL_48_DFFSR_100 ( );
FILL FILL_49_DFFSR_100 ( );
FILL FILL_50_DFFSR_100 ( );
FILL FILL_51_DFFSR_100 ( );
FILL FILL_0_DFFSR_181 ( );
FILL FILL_1_DFFSR_181 ( );
FILL FILL_2_DFFSR_181 ( );
FILL FILL_3_DFFSR_181 ( );
FILL FILL_4_DFFSR_181 ( );
FILL FILL_5_DFFSR_181 ( );
FILL FILL_6_DFFSR_181 ( );
FILL FILL_7_DFFSR_181 ( );
FILL FILL_8_DFFSR_181 ( );
FILL FILL_9_DFFSR_181 ( );
FILL FILL_10_DFFSR_181 ( );
FILL FILL_11_DFFSR_181 ( );
FILL FILL_12_DFFSR_181 ( );
FILL FILL_13_DFFSR_181 ( );
FILL FILL_14_DFFSR_181 ( );
FILL FILL_15_DFFSR_181 ( );
FILL FILL_16_DFFSR_181 ( );
FILL FILL_17_DFFSR_181 ( );
FILL FILL_18_DFFSR_181 ( );
FILL FILL_19_DFFSR_181 ( );
FILL FILL_20_DFFSR_181 ( );
FILL FILL_21_DFFSR_181 ( );
FILL FILL_22_DFFSR_181 ( );
FILL FILL_23_DFFSR_181 ( );
FILL FILL_24_DFFSR_181 ( );
FILL FILL_25_DFFSR_181 ( );
FILL FILL_26_DFFSR_181 ( );
FILL FILL_27_DFFSR_181 ( );
FILL FILL_28_DFFSR_181 ( );
FILL FILL_29_DFFSR_181 ( );
FILL FILL_30_DFFSR_181 ( );
FILL FILL_31_DFFSR_181 ( );
FILL FILL_32_DFFSR_181 ( );
FILL FILL_33_DFFSR_181 ( );
FILL FILL_34_DFFSR_181 ( );
FILL FILL_35_DFFSR_181 ( );
FILL FILL_36_DFFSR_181 ( );
FILL FILL_37_DFFSR_181 ( );
FILL FILL_38_DFFSR_181 ( );
FILL FILL_39_DFFSR_181 ( );
FILL FILL_40_DFFSR_181 ( );
FILL FILL_41_DFFSR_181 ( );
FILL FILL_42_DFFSR_181 ( );
FILL FILL_43_DFFSR_181 ( );
FILL FILL_44_DFFSR_181 ( );
FILL FILL_45_DFFSR_181 ( );
FILL FILL_46_DFFSR_181 ( );
FILL FILL_47_DFFSR_181 ( );
FILL FILL_48_DFFSR_181 ( );
FILL FILL_49_DFFSR_181 ( );
FILL FILL_50_DFFSR_181 ( );
FILL FILL_0_NAND2X1_6 ( );
FILL FILL_1_NAND2X1_6 ( );
FILL FILL_2_NAND2X1_6 ( );
FILL FILL_3_NAND2X1_6 ( );
FILL FILL_4_NAND2X1_6 ( );
FILL FILL_5_NAND2X1_6 ( );
FILL FILL_6_NAND2X1_6 ( );
FILL FILL_0_INVX1_187 ( );
FILL FILL_1_INVX1_187 ( );
FILL FILL_2_INVX1_187 ( );
FILL FILL_3_INVX1_187 ( );
FILL FILL_4_INVX1_187 ( );
FILL FILL_0_INVX1_165 ( );
FILL FILL_1_INVX1_165 ( );
FILL FILL_2_INVX1_165 ( );
FILL FILL_3_INVX1_165 ( );
FILL FILL_4_INVX1_165 ( );
FILL FILL_0_DFFSR_145 ( );
FILL FILL_1_DFFSR_145 ( );
FILL FILL_2_DFFSR_145 ( );
FILL FILL_3_DFFSR_145 ( );
FILL FILL_4_DFFSR_145 ( );
FILL FILL_5_DFFSR_145 ( );
FILL FILL_6_DFFSR_145 ( );
FILL FILL_7_DFFSR_145 ( );
FILL FILL_8_DFFSR_145 ( );
FILL FILL_9_DFFSR_145 ( );
FILL FILL_10_DFFSR_145 ( );
FILL FILL_11_DFFSR_145 ( );
FILL FILL_12_DFFSR_145 ( );
FILL FILL_13_DFFSR_145 ( );
FILL FILL_14_DFFSR_145 ( );
FILL FILL_15_DFFSR_145 ( );
FILL FILL_16_DFFSR_145 ( );
FILL FILL_17_DFFSR_145 ( );
FILL FILL_18_DFFSR_145 ( );
FILL FILL_19_DFFSR_145 ( );
FILL FILL_20_DFFSR_145 ( );
FILL FILL_21_DFFSR_145 ( );
FILL FILL_22_DFFSR_145 ( );
FILL FILL_23_DFFSR_145 ( );
FILL FILL_24_DFFSR_145 ( );
FILL FILL_25_DFFSR_145 ( );
FILL FILL_26_DFFSR_145 ( );
FILL FILL_27_DFFSR_145 ( );
FILL FILL_28_DFFSR_145 ( );
FILL FILL_29_DFFSR_145 ( );
FILL FILL_30_DFFSR_145 ( );
FILL FILL_31_DFFSR_145 ( );
FILL FILL_32_DFFSR_145 ( );
FILL FILL_33_DFFSR_145 ( );
FILL FILL_34_DFFSR_145 ( );
FILL FILL_35_DFFSR_145 ( );
FILL FILL_36_DFFSR_145 ( );
FILL FILL_37_DFFSR_145 ( );
FILL FILL_38_DFFSR_145 ( );
FILL FILL_39_DFFSR_145 ( );
FILL FILL_40_DFFSR_145 ( );
FILL FILL_41_DFFSR_145 ( );
FILL FILL_42_DFFSR_145 ( );
FILL FILL_43_DFFSR_145 ( );
FILL FILL_44_DFFSR_145 ( );
FILL FILL_45_DFFSR_145 ( );
FILL FILL_46_DFFSR_145 ( );
FILL FILL_47_DFFSR_145 ( );
FILL FILL_48_DFFSR_145 ( );
FILL FILL_49_DFFSR_145 ( );
FILL FILL_50_DFFSR_145 ( );
FILL FILL_0_CLKBUF1_25 ( );
FILL FILL_1_CLKBUF1_25 ( );
FILL FILL_2_CLKBUF1_25 ( );
FILL FILL_3_CLKBUF1_25 ( );
FILL FILL_4_CLKBUF1_25 ( );
FILL FILL_5_CLKBUF1_25 ( );
FILL FILL_6_CLKBUF1_25 ( );
FILL FILL_7_CLKBUF1_25 ( );
FILL FILL_8_CLKBUF1_25 ( );
FILL FILL_9_CLKBUF1_25 ( );
FILL FILL_10_CLKBUF1_25 ( );
FILL FILL_11_CLKBUF1_25 ( );
FILL FILL_12_CLKBUF1_25 ( );
FILL FILL_13_CLKBUF1_25 ( );
FILL FILL_14_CLKBUF1_25 ( );
FILL FILL_15_CLKBUF1_25 ( );
FILL FILL_16_CLKBUF1_25 ( );
FILL FILL_17_CLKBUF1_25 ( );
FILL FILL_18_CLKBUF1_25 ( );
FILL FILL_19_CLKBUF1_25 ( );
FILL FILL_0_CLKBUF1_24 ( );
FILL FILL_1_CLKBUF1_24 ( );
FILL FILL_2_CLKBUF1_24 ( );
FILL FILL_3_CLKBUF1_24 ( );
FILL FILL_4_CLKBUF1_24 ( );
FILL FILL_5_CLKBUF1_24 ( );
FILL FILL_6_CLKBUF1_24 ( );
FILL FILL_7_CLKBUF1_24 ( );
FILL FILL_8_CLKBUF1_24 ( );
FILL FILL_9_CLKBUF1_24 ( );
FILL FILL_10_CLKBUF1_24 ( );
FILL FILL_11_CLKBUF1_24 ( );
FILL FILL_12_CLKBUF1_24 ( );
FILL FILL_13_CLKBUF1_24 ( );
FILL FILL_14_CLKBUF1_24 ( );
FILL FILL_15_CLKBUF1_24 ( );
FILL FILL_16_CLKBUF1_24 ( );
FILL FILL_17_CLKBUF1_24 ( );
FILL FILL_18_CLKBUF1_24 ( );
FILL FILL_19_CLKBUF1_24 ( );
FILL FILL_20_CLKBUF1_24 ( );
FILL FILL_0_NAND2X1_222 ( );
FILL FILL_1_NAND2X1_222 ( );
FILL FILL_2_NAND2X1_222 ( );
FILL FILL_3_NAND2X1_222 ( );
FILL FILL_4_NAND2X1_222 ( );
FILL FILL_5_NAND2X1_222 ( );
FILL FILL_6_NAND2X1_222 ( );
FILL FILL_0_NAND2X1_20 ( );
FILL FILL_1_NAND2X1_20 ( );
FILL FILL_2_NAND2X1_20 ( );
FILL FILL_3_NAND2X1_20 ( );
FILL FILL_4_NAND2X1_20 ( );
FILL FILL_5_NAND2X1_20 ( );
FILL FILL_6_NAND2X1_20 ( );
FILL FILL_0_INVX1_208 ( );
FILL FILL_1_INVX1_208 ( );
FILL FILL_2_INVX1_208 ( );
FILL FILL_3_INVX1_208 ( );
FILL FILL_0_DFFSR_186 ( );
FILL FILL_1_DFFSR_186 ( );
FILL FILL_2_DFFSR_186 ( );
FILL FILL_3_DFFSR_186 ( );
FILL FILL_4_DFFSR_186 ( );
FILL FILL_5_DFFSR_186 ( );
FILL FILL_6_DFFSR_186 ( );
FILL FILL_7_DFFSR_186 ( );
FILL FILL_8_DFFSR_186 ( );
FILL FILL_9_DFFSR_186 ( );
FILL FILL_10_DFFSR_186 ( );
FILL FILL_11_DFFSR_186 ( );
FILL FILL_12_DFFSR_186 ( );
FILL FILL_13_DFFSR_186 ( );
FILL FILL_14_DFFSR_186 ( );
FILL FILL_15_DFFSR_186 ( );
FILL FILL_16_DFFSR_186 ( );
FILL FILL_17_DFFSR_186 ( );
FILL FILL_18_DFFSR_186 ( );
FILL FILL_19_DFFSR_186 ( );
FILL FILL_20_DFFSR_186 ( );
FILL FILL_21_DFFSR_186 ( );
FILL FILL_22_DFFSR_186 ( );
FILL FILL_23_DFFSR_186 ( );
FILL FILL_24_DFFSR_186 ( );
FILL FILL_25_DFFSR_186 ( );
FILL FILL_26_DFFSR_186 ( );
FILL FILL_27_DFFSR_186 ( );
FILL FILL_28_DFFSR_186 ( );
FILL FILL_29_DFFSR_186 ( );
FILL FILL_30_DFFSR_186 ( );
FILL FILL_31_DFFSR_186 ( );
FILL FILL_32_DFFSR_186 ( );
FILL FILL_33_DFFSR_186 ( );
FILL FILL_34_DFFSR_186 ( );
FILL FILL_35_DFFSR_186 ( );
FILL FILL_36_DFFSR_186 ( );
FILL FILL_37_DFFSR_186 ( );
FILL FILL_38_DFFSR_186 ( );
FILL FILL_39_DFFSR_186 ( );
FILL FILL_40_DFFSR_186 ( );
FILL FILL_41_DFFSR_186 ( );
FILL FILL_42_DFFSR_186 ( );
FILL FILL_43_DFFSR_186 ( );
FILL FILL_44_DFFSR_186 ( );
FILL FILL_45_DFFSR_186 ( );
FILL FILL_46_DFFSR_186 ( );
FILL FILL_47_DFFSR_186 ( );
FILL FILL_48_DFFSR_186 ( );
FILL FILL_49_DFFSR_186 ( );
FILL FILL_50_DFFSR_186 ( );
FILL FILL_51_DFFSR_186 ( );
FILL FILL_0_OAI21X1_230 ( );
FILL FILL_1_OAI21X1_230 ( );
FILL FILL_2_OAI21X1_230 ( );
FILL FILL_3_OAI21X1_230 ( );
FILL FILL_4_OAI21X1_230 ( );
FILL FILL_5_OAI21X1_230 ( );
FILL FILL_6_OAI21X1_230 ( );
FILL FILL_7_OAI21X1_230 ( );
FILL FILL_8_OAI21X1_230 ( );
FILL FILL_9_OAI21X1_230 ( );
FILL FILL_0_AOI22X1_13 ( );
FILL FILL_1_AOI22X1_13 ( );
FILL FILL_2_AOI22X1_13 ( );
FILL FILL_3_AOI22X1_13 ( );
FILL FILL_4_AOI22X1_13 ( );
FILL FILL_5_AOI22X1_13 ( );
FILL FILL_6_AOI22X1_13 ( );
FILL FILL_7_AOI22X1_13 ( );
FILL FILL_8_AOI22X1_13 ( );
FILL FILL_9_AOI22X1_13 ( );
FILL FILL_10_AOI22X1_13 ( );
FILL FILL_0_OAI21X1_218 ( );
FILL FILL_1_OAI21X1_218 ( );
FILL FILL_2_OAI21X1_218 ( );
FILL FILL_3_OAI21X1_218 ( );
FILL FILL_4_OAI21X1_218 ( );
FILL FILL_5_OAI21X1_218 ( );
FILL FILL_6_OAI21X1_218 ( );
FILL FILL_7_OAI21X1_218 ( );
FILL FILL_8_OAI21X1_218 ( );
FILL FILL_9_OAI21X1_218 ( );
FILL FILL_0_NAND2X1_212 ( );
FILL FILL_1_NAND2X1_212 ( );
FILL FILL_2_NAND2X1_212 ( );
FILL FILL_3_NAND2X1_212 ( );
FILL FILL_4_NAND2X1_212 ( );
FILL FILL_5_NAND2X1_212 ( );
FILL FILL_6_NAND2X1_212 ( );
FILL FILL_0_NAND2X1_161 ( );
FILL FILL_1_NAND2X1_161 ( );
FILL FILL_2_NAND2X1_161 ( );
FILL FILL_3_NAND2X1_161 ( );
FILL FILL_4_NAND2X1_161 ( );
FILL FILL_5_NAND2X1_161 ( );
FILL FILL_6_NAND2X1_161 ( );
FILL FILL_0_OAI21X1_161 ( );
FILL FILL_1_OAI21X1_161 ( );
FILL FILL_2_OAI21X1_161 ( );
FILL FILL_3_OAI21X1_161 ( );
FILL FILL_4_OAI21X1_161 ( );
FILL FILL_5_OAI21X1_161 ( );
FILL FILL_6_OAI21X1_161 ( );
FILL FILL_7_OAI21X1_161 ( );
FILL FILL_8_OAI21X1_161 ( );
FILL FILL_0_INVX1_195 ( );
FILL FILL_1_INVX1_195 ( );
FILL FILL_2_INVX1_195 ( );
FILL FILL_3_INVX1_195 ( );
FILL FILL_4_INVX1_195 ( );
FILL FILL_0_INVX1_422 ( );
FILL FILL_1_INVX1_422 ( );
FILL FILL_2_INVX1_422 ( );
FILL FILL_3_INVX1_422 ( );
FILL FILL_4_INVX1_422 ( );
FILL FILL_0_OAI21X1_259 ( );
FILL FILL_1_OAI21X1_259 ( );
FILL FILL_2_OAI21X1_259 ( );
FILL FILL_3_OAI21X1_259 ( );
FILL FILL_4_OAI21X1_259 ( );
FILL FILL_5_OAI21X1_259 ( );
FILL FILL_6_OAI21X1_259 ( );
FILL FILL_7_OAI21X1_259 ( );
FILL FILL_8_OAI21X1_259 ( );
FILL FILL_0_AOI21X1_31 ( );
FILL FILL_1_AOI21X1_31 ( );
FILL FILL_2_AOI21X1_31 ( );
FILL FILL_3_AOI21X1_31 ( );
FILL FILL_4_AOI21X1_31 ( );
FILL FILL_5_AOI21X1_31 ( );
FILL FILL_6_AOI21X1_31 ( );
FILL FILL_7_AOI21X1_31 ( );
FILL FILL_8_AOI21X1_31 ( );
FILL FILL_0_NAND3X1_102 ( );
FILL FILL_1_NAND3X1_102 ( );
FILL FILL_2_NAND3X1_102 ( );
FILL FILL_3_NAND3X1_102 ( );
FILL FILL_4_NAND3X1_102 ( );
FILL FILL_5_NAND3X1_102 ( );
FILL FILL_6_NAND3X1_102 ( );
FILL FILL_7_NAND3X1_102 ( );
FILL FILL_8_NAND3X1_102 ( );
FILL FILL_0_NAND3X1_104 ( );
FILL FILL_1_NAND3X1_104 ( );
FILL FILL_2_NAND3X1_104 ( );
FILL FILL_3_NAND3X1_104 ( );
FILL FILL_4_NAND3X1_104 ( );
FILL FILL_5_NAND3X1_104 ( );
FILL FILL_6_NAND3X1_104 ( );
FILL FILL_7_NAND3X1_104 ( );
FILL FILL_8_NAND3X1_104 ( );
FILL FILL_0_NAND3X1_103 ( );
FILL FILL_1_NAND3X1_103 ( );
FILL FILL_2_NAND3X1_103 ( );
FILL FILL_3_NAND3X1_103 ( );
FILL FILL_4_NAND3X1_103 ( );
FILL FILL_5_NAND3X1_103 ( );
FILL FILL_6_NAND3X1_103 ( );
FILL FILL_7_NAND3X1_103 ( );
FILL FILL_8_NAND3X1_103 ( );
FILL FILL_0_NAND2X1_113 ( );
FILL FILL_1_NAND2X1_113 ( );
FILL FILL_2_NAND2X1_113 ( );
FILL FILL_3_NAND2X1_113 ( );
FILL FILL_4_NAND2X1_113 ( );
FILL FILL_5_NAND2X1_113 ( );
FILL FILL_6_NAND2X1_113 ( );
FILL FILL_0_OAI21X1_113 ( );
FILL FILL_1_OAI21X1_113 ( );
FILL FILL_2_OAI21X1_113 ( );
FILL FILL_3_OAI21X1_113 ( );
FILL FILL_4_OAI21X1_113 ( );
FILL FILL_5_OAI21X1_113 ( );
FILL FILL_6_OAI21X1_113 ( );
FILL FILL_7_OAI21X1_113 ( );
FILL FILL_8_OAI21X1_113 ( );
FILL FILL_0_INVX1_128 ( );
FILL FILL_1_INVX1_128 ( );
FILL FILL_2_INVX1_128 ( );
FILL FILL_3_INVX1_128 ( );
FILL FILL_4_INVX1_128 ( );
FILL FILL_0_DFFSR_117 ( );
FILL FILL_1_DFFSR_117 ( );
FILL FILL_2_DFFSR_117 ( );
FILL FILL_3_DFFSR_117 ( );
FILL FILL_4_DFFSR_117 ( );
FILL FILL_5_DFFSR_117 ( );
FILL FILL_6_DFFSR_117 ( );
FILL FILL_7_DFFSR_117 ( );
FILL FILL_8_DFFSR_117 ( );
FILL FILL_9_DFFSR_117 ( );
FILL FILL_10_DFFSR_117 ( );
FILL FILL_11_DFFSR_117 ( );
FILL FILL_12_DFFSR_117 ( );
FILL FILL_13_DFFSR_117 ( );
FILL FILL_14_DFFSR_117 ( );
FILL FILL_15_DFFSR_117 ( );
FILL FILL_16_DFFSR_117 ( );
FILL FILL_17_DFFSR_117 ( );
FILL FILL_18_DFFSR_117 ( );
FILL FILL_19_DFFSR_117 ( );
FILL FILL_20_DFFSR_117 ( );
FILL FILL_21_DFFSR_117 ( );
FILL FILL_22_DFFSR_117 ( );
FILL FILL_23_DFFSR_117 ( );
FILL FILL_24_DFFSR_117 ( );
FILL FILL_25_DFFSR_117 ( );
FILL FILL_26_DFFSR_117 ( );
FILL FILL_27_DFFSR_117 ( );
FILL FILL_28_DFFSR_117 ( );
FILL FILL_29_DFFSR_117 ( );
FILL FILL_30_DFFSR_117 ( );
FILL FILL_31_DFFSR_117 ( );
FILL FILL_32_DFFSR_117 ( );
FILL FILL_33_DFFSR_117 ( );
FILL FILL_34_DFFSR_117 ( );
FILL FILL_35_DFFSR_117 ( );
FILL FILL_36_DFFSR_117 ( );
FILL FILL_37_DFFSR_117 ( );
FILL FILL_38_DFFSR_117 ( );
FILL FILL_39_DFFSR_117 ( );
FILL FILL_40_DFFSR_117 ( );
FILL FILL_41_DFFSR_117 ( );
FILL FILL_42_DFFSR_117 ( );
FILL FILL_43_DFFSR_117 ( );
FILL FILL_44_DFFSR_117 ( );
FILL FILL_45_DFFSR_117 ( );
FILL FILL_46_DFFSR_117 ( );
FILL FILL_47_DFFSR_117 ( );
FILL FILL_48_DFFSR_117 ( );
FILL FILL_49_DFFSR_117 ( );
FILL FILL_50_DFFSR_117 ( );
FILL FILL_0_OAI21X1_123 ( );
FILL FILL_1_OAI21X1_123 ( );
FILL FILL_2_OAI21X1_123 ( );
FILL FILL_3_OAI21X1_123 ( );
FILL FILL_4_OAI21X1_123 ( );
FILL FILL_5_OAI21X1_123 ( );
FILL FILL_6_OAI21X1_123 ( );
FILL FILL_7_OAI21X1_123 ( );
FILL FILL_8_OAI21X1_123 ( );
FILL FILL_0_OAI21X1_100 ( );
FILL FILL_1_OAI21X1_100 ( );
FILL FILL_2_OAI21X1_100 ( );
FILL FILL_3_OAI21X1_100 ( );
FILL FILL_4_OAI21X1_100 ( );
FILL FILL_5_OAI21X1_100 ( );
FILL FILL_6_OAI21X1_100 ( );
FILL FILL_7_OAI21X1_100 ( );
FILL FILL_8_OAI21X1_100 ( );
FILL FILL_9_OAI21X1_100 ( );
FILL FILL_0_INVX1_113 ( );
FILL FILL_1_INVX1_113 ( );
FILL FILL_2_INVX1_113 ( );
FILL FILL_3_INVX1_113 ( );
FILL FILL_0_DFFSR_149 ( );
FILL FILL_1_DFFSR_149 ( );
FILL FILL_2_DFFSR_149 ( );
FILL FILL_3_DFFSR_149 ( );
FILL FILL_4_DFFSR_149 ( );
FILL FILL_5_DFFSR_149 ( );
FILL FILL_6_DFFSR_149 ( );
FILL FILL_7_DFFSR_149 ( );
FILL FILL_8_DFFSR_149 ( );
FILL FILL_9_DFFSR_149 ( );
FILL FILL_10_DFFSR_149 ( );
FILL FILL_11_DFFSR_149 ( );
FILL FILL_12_DFFSR_149 ( );
FILL FILL_13_DFFSR_149 ( );
FILL FILL_14_DFFSR_149 ( );
FILL FILL_15_DFFSR_149 ( );
FILL FILL_16_DFFSR_149 ( );
FILL FILL_17_DFFSR_149 ( );
FILL FILL_18_DFFSR_149 ( );
FILL FILL_19_DFFSR_149 ( );
FILL FILL_20_DFFSR_149 ( );
FILL FILL_21_DFFSR_149 ( );
FILL FILL_22_DFFSR_149 ( );
FILL FILL_23_DFFSR_149 ( );
FILL FILL_24_DFFSR_149 ( );
FILL FILL_25_DFFSR_149 ( );
FILL FILL_26_DFFSR_149 ( );
FILL FILL_27_DFFSR_149 ( );
FILL FILL_28_DFFSR_149 ( );
FILL FILL_29_DFFSR_149 ( );
FILL FILL_30_DFFSR_149 ( );
FILL FILL_31_DFFSR_149 ( );
FILL FILL_32_DFFSR_149 ( );
FILL FILL_33_DFFSR_149 ( );
FILL FILL_34_DFFSR_149 ( );
FILL FILL_35_DFFSR_149 ( );
FILL FILL_36_DFFSR_149 ( );
FILL FILL_37_DFFSR_149 ( );
FILL FILL_38_DFFSR_149 ( );
FILL FILL_39_DFFSR_149 ( );
FILL FILL_40_DFFSR_149 ( );
FILL FILL_41_DFFSR_149 ( );
FILL FILL_42_DFFSR_149 ( );
FILL FILL_43_DFFSR_149 ( );
FILL FILL_44_DFFSR_149 ( );
FILL FILL_45_DFFSR_149 ( );
FILL FILL_46_DFFSR_149 ( );
FILL FILL_47_DFFSR_149 ( );
FILL FILL_48_DFFSR_149 ( );
FILL FILL_49_DFFSR_149 ( );
FILL FILL_50_DFFSR_149 ( );
FILL FILL_0_DFFSR_156 ( );
FILL FILL_1_DFFSR_156 ( );
FILL FILL_2_DFFSR_156 ( );
FILL FILL_3_DFFSR_156 ( );
FILL FILL_4_DFFSR_156 ( );
FILL FILL_5_DFFSR_156 ( );
FILL FILL_6_DFFSR_156 ( );
FILL FILL_7_DFFSR_156 ( );
FILL FILL_8_DFFSR_156 ( );
FILL FILL_9_DFFSR_156 ( );
FILL FILL_10_DFFSR_156 ( );
FILL FILL_11_DFFSR_156 ( );
FILL FILL_12_DFFSR_156 ( );
FILL FILL_13_DFFSR_156 ( );
FILL FILL_14_DFFSR_156 ( );
FILL FILL_15_DFFSR_156 ( );
FILL FILL_16_DFFSR_156 ( );
FILL FILL_17_DFFSR_156 ( );
FILL FILL_18_DFFSR_156 ( );
FILL FILL_19_DFFSR_156 ( );
FILL FILL_20_DFFSR_156 ( );
FILL FILL_21_DFFSR_156 ( );
FILL FILL_22_DFFSR_156 ( );
FILL FILL_23_DFFSR_156 ( );
FILL FILL_24_DFFSR_156 ( );
FILL FILL_25_DFFSR_156 ( );
FILL FILL_26_DFFSR_156 ( );
FILL FILL_27_DFFSR_156 ( );
FILL FILL_28_DFFSR_156 ( );
FILL FILL_29_DFFSR_156 ( );
FILL FILL_30_DFFSR_156 ( );
FILL FILL_31_DFFSR_156 ( );
FILL FILL_32_DFFSR_156 ( );
FILL FILL_33_DFFSR_156 ( );
FILL FILL_34_DFFSR_156 ( );
FILL FILL_35_DFFSR_156 ( );
FILL FILL_36_DFFSR_156 ( );
FILL FILL_37_DFFSR_156 ( );
FILL FILL_38_DFFSR_156 ( );
FILL FILL_39_DFFSR_156 ( );
FILL FILL_40_DFFSR_156 ( );
FILL FILL_41_DFFSR_156 ( );
FILL FILL_42_DFFSR_156 ( );
FILL FILL_43_DFFSR_156 ( );
FILL FILL_44_DFFSR_156 ( );
FILL FILL_45_DFFSR_156 ( );
FILL FILL_46_DFFSR_156 ( );
FILL FILL_47_DFFSR_156 ( );
FILL FILL_48_DFFSR_156 ( );
FILL FILL_49_DFFSR_156 ( );
FILL FILL_50_DFFSR_156 ( );
FILL FILL_0_OAI21X1_145 ( );
FILL FILL_1_OAI21X1_145 ( );
FILL FILL_2_OAI21X1_145 ( );
FILL FILL_3_OAI21X1_145 ( );
FILL FILL_4_OAI21X1_145 ( );
FILL FILL_5_OAI21X1_145 ( );
FILL FILL_6_OAI21X1_145 ( );
FILL FILL_7_OAI21X1_145 ( );
FILL FILL_8_OAI21X1_145 ( );
FILL FILL_0_INVX1_164 ( );
FILL FILL_1_INVX1_164 ( );
FILL FILL_2_INVX1_164 ( );
FILL FILL_3_INVX1_164 ( );
FILL FILL_4_INVX1_164 ( );
FILL FILL_0_AOI21X1_42 ( );
FILL FILL_1_AOI21X1_42 ( );
FILL FILL_2_AOI21X1_42 ( );
FILL FILL_3_AOI21X1_42 ( );
FILL FILL_4_AOI21X1_42 ( );
FILL FILL_5_AOI21X1_42 ( );
FILL FILL_6_AOI21X1_42 ( );
FILL FILL_7_AOI21X1_42 ( );
FILL FILL_8_AOI21X1_42 ( );
FILL FILL_9_AOI21X1_42 ( );
FILL FILL_0_NAND2X1_146 ( );
FILL FILL_1_NAND2X1_146 ( );
FILL FILL_2_NAND2X1_146 ( );
FILL FILL_3_NAND2X1_146 ( );
FILL FILL_4_NAND2X1_146 ( );
FILL FILL_5_NAND2X1_146 ( );
FILL FILL_6_NAND2X1_146 ( );
FILL FILL_0_DFFSR_175 ( );
FILL FILL_1_DFFSR_175 ( );
FILL FILL_2_DFFSR_175 ( );
FILL FILL_3_DFFSR_175 ( );
FILL FILL_4_DFFSR_175 ( );
FILL FILL_5_DFFSR_175 ( );
FILL FILL_6_DFFSR_175 ( );
FILL FILL_7_DFFSR_175 ( );
FILL FILL_8_DFFSR_175 ( );
FILL FILL_9_DFFSR_175 ( );
FILL FILL_10_DFFSR_175 ( );
FILL FILL_11_DFFSR_175 ( );
FILL FILL_12_DFFSR_175 ( );
FILL FILL_13_DFFSR_175 ( );
FILL FILL_14_DFFSR_175 ( );
FILL FILL_15_DFFSR_175 ( );
FILL FILL_16_DFFSR_175 ( );
FILL FILL_17_DFFSR_175 ( );
FILL FILL_18_DFFSR_175 ( );
FILL FILL_19_DFFSR_175 ( );
FILL FILL_20_DFFSR_175 ( );
FILL FILL_21_DFFSR_175 ( );
FILL FILL_22_DFFSR_175 ( );
FILL FILL_23_DFFSR_175 ( );
FILL FILL_24_DFFSR_175 ( );
FILL FILL_25_DFFSR_175 ( );
FILL FILL_26_DFFSR_175 ( );
FILL FILL_27_DFFSR_175 ( );
FILL FILL_28_DFFSR_175 ( );
FILL FILL_29_DFFSR_175 ( );
FILL FILL_30_DFFSR_175 ( );
FILL FILL_31_DFFSR_175 ( );
FILL FILL_32_DFFSR_175 ( );
FILL FILL_33_DFFSR_175 ( );
FILL FILL_34_DFFSR_175 ( );
FILL FILL_35_DFFSR_175 ( );
FILL FILL_36_DFFSR_175 ( );
FILL FILL_37_DFFSR_175 ( );
FILL FILL_38_DFFSR_175 ( );
FILL FILL_39_DFFSR_175 ( );
FILL FILL_40_DFFSR_175 ( );
FILL FILL_41_DFFSR_175 ( );
FILL FILL_42_DFFSR_175 ( );
FILL FILL_43_DFFSR_175 ( );
FILL FILL_44_DFFSR_175 ( );
FILL FILL_45_DFFSR_175 ( );
FILL FILL_46_DFFSR_175 ( );
FILL FILL_47_DFFSR_175 ( );
FILL FILL_48_DFFSR_175 ( );
FILL FILL_49_DFFSR_175 ( );
FILL FILL_50_DFFSR_175 ( );
FILL FILL_0_INVX1_23 ( );
FILL FILL_1_INVX1_23 ( );
FILL FILL_2_INVX1_23 ( );
FILL FILL_3_INVX1_23 ( );
FILL FILL_4_INVX1_23 ( );
FILL FILL_0_DFFPOSX1_23 ( );
FILL FILL_1_DFFPOSX1_23 ( );
FILL FILL_2_DFFPOSX1_23 ( );
FILL FILL_3_DFFPOSX1_23 ( );
FILL FILL_4_DFFPOSX1_23 ( );
FILL FILL_5_DFFPOSX1_23 ( );
FILL FILL_6_DFFPOSX1_23 ( );
FILL FILL_7_DFFPOSX1_23 ( );
FILL FILL_8_DFFPOSX1_23 ( );
FILL FILL_9_DFFPOSX1_23 ( );
FILL FILL_10_DFFPOSX1_23 ( );
FILL FILL_11_DFFPOSX1_23 ( );
FILL FILL_12_DFFPOSX1_23 ( );
FILL FILL_13_DFFPOSX1_23 ( );
FILL FILL_14_DFFPOSX1_23 ( );
FILL FILL_15_DFFPOSX1_23 ( );
FILL FILL_16_DFFPOSX1_23 ( );
FILL FILL_17_DFFPOSX1_23 ( );
FILL FILL_18_DFFPOSX1_23 ( );
FILL FILL_19_DFFPOSX1_23 ( );
FILL FILL_20_DFFPOSX1_23 ( );
FILL FILL_21_DFFPOSX1_23 ( );
FILL FILL_22_DFFPOSX1_23 ( );
FILL FILL_23_DFFPOSX1_23 ( );
FILL FILL_24_DFFPOSX1_23 ( );
FILL FILL_25_DFFPOSX1_23 ( );
FILL FILL_26_DFFPOSX1_23 ( );
FILL FILL_27_DFFPOSX1_23 ( );
FILL FILL_0_INVX1_417 ( );
FILL FILL_1_INVX1_417 ( );
FILL FILL_2_INVX1_417 ( );
FILL FILL_3_INVX1_417 ( );
FILL FILL_4_INVX1_417 ( );
FILL FILL_0_OAI21X1_254 ( );
FILL FILL_1_OAI21X1_254 ( );
FILL FILL_2_OAI21X1_254 ( );
FILL FILL_3_OAI21X1_254 ( );
FILL FILL_4_OAI21X1_254 ( );
FILL FILL_5_OAI21X1_254 ( );
FILL FILL_6_OAI21X1_254 ( );
FILL FILL_7_OAI21X1_254 ( );
FILL FILL_8_OAI21X1_254 ( );
FILL FILL_0_OAI21X1_217 ( );
FILL FILL_1_OAI21X1_217 ( );
FILL FILL_2_OAI21X1_217 ( );
FILL FILL_3_OAI21X1_217 ( );
FILL FILL_4_OAI21X1_217 ( );
FILL FILL_5_OAI21X1_217 ( );
FILL FILL_6_OAI21X1_217 ( );
FILL FILL_7_OAI21X1_217 ( );
FILL FILL_8_OAI21X1_217 ( );
FILL FILL_0_OAI21X1_162 ( );
FILL FILL_1_OAI21X1_162 ( );
FILL FILL_2_OAI21X1_162 ( );
FILL FILL_3_OAI21X1_162 ( );
FILL FILL_4_OAI21X1_162 ( );
FILL FILL_5_OAI21X1_162 ( );
FILL FILL_6_OAI21X1_162 ( );
FILL FILL_7_OAI21X1_162 ( );
FILL FILL_8_OAI21X1_162 ( );
FILL FILL_0_NAND2X1_228 ( );
FILL FILL_1_NAND2X1_228 ( );
FILL FILL_2_NAND2X1_228 ( );
FILL FILL_3_NAND2X1_228 ( );
FILL FILL_4_NAND2X1_228 ( );
FILL FILL_5_NAND2X1_228 ( );
FILL FILL_6_NAND2X1_228 ( );
FILL FILL_0_AOI22X1_11 ( );
FILL FILL_1_AOI22X1_11 ( );
FILL FILL_2_AOI22X1_11 ( );
FILL FILL_3_AOI22X1_11 ( );
FILL FILL_4_AOI22X1_11 ( );
FILL FILL_5_AOI22X1_11 ( );
FILL FILL_6_AOI22X1_11 ( );
FILL FILL_7_AOI22X1_11 ( );
FILL FILL_8_AOI22X1_11 ( );
FILL FILL_9_AOI22X1_11 ( );
FILL FILL_10_AOI22X1_11 ( );
FILL FILL_0_XOR2X1_7 ( );
FILL FILL_1_XOR2X1_7 ( );
FILL FILL_2_XOR2X1_7 ( );
FILL FILL_3_XOR2X1_7 ( );
FILL FILL_4_XOR2X1_7 ( );
FILL FILL_5_XOR2X1_7 ( );
FILL FILL_6_XOR2X1_7 ( );
FILL FILL_7_XOR2X1_7 ( );
FILL FILL_8_XOR2X1_7 ( );
FILL FILL_9_XOR2X1_7 ( );
FILL FILL_10_XOR2X1_7 ( );
FILL FILL_11_XOR2X1_7 ( );
FILL FILL_12_XOR2X1_7 ( );
FILL FILL_13_XOR2X1_7 ( );
FILL FILL_14_XOR2X1_7 ( );
FILL FILL_15_XOR2X1_7 ( );
FILL FILL_16_XOR2X1_7 ( );
FILL FILL_0_DFFSR_191 ( );
FILL FILL_1_DFFSR_191 ( );
FILL FILL_2_DFFSR_191 ( );
FILL FILL_3_DFFSR_191 ( );
FILL FILL_4_DFFSR_191 ( );
FILL FILL_5_DFFSR_191 ( );
FILL FILL_6_DFFSR_191 ( );
FILL FILL_7_DFFSR_191 ( );
FILL FILL_8_DFFSR_191 ( );
FILL FILL_9_DFFSR_191 ( );
FILL FILL_10_DFFSR_191 ( );
FILL FILL_11_DFFSR_191 ( );
FILL FILL_12_DFFSR_191 ( );
FILL FILL_13_DFFSR_191 ( );
FILL FILL_14_DFFSR_191 ( );
FILL FILL_15_DFFSR_191 ( );
FILL FILL_16_DFFSR_191 ( );
FILL FILL_17_DFFSR_191 ( );
FILL FILL_18_DFFSR_191 ( );
FILL FILL_19_DFFSR_191 ( );
FILL FILL_20_DFFSR_191 ( );
FILL FILL_21_DFFSR_191 ( );
FILL FILL_22_DFFSR_191 ( );
FILL FILL_23_DFFSR_191 ( );
FILL FILL_24_DFFSR_191 ( );
FILL FILL_25_DFFSR_191 ( );
FILL FILL_26_DFFSR_191 ( );
FILL FILL_27_DFFSR_191 ( );
FILL FILL_28_DFFSR_191 ( );
FILL FILL_29_DFFSR_191 ( );
FILL FILL_30_DFFSR_191 ( );
FILL FILL_31_DFFSR_191 ( );
FILL FILL_32_DFFSR_191 ( );
FILL FILL_33_DFFSR_191 ( );
FILL FILL_34_DFFSR_191 ( );
FILL FILL_35_DFFSR_191 ( );
FILL FILL_36_DFFSR_191 ( );
FILL FILL_37_DFFSR_191 ( );
FILL FILL_38_DFFSR_191 ( );
FILL FILL_39_DFFSR_191 ( );
FILL FILL_40_DFFSR_191 ( );
FILL FILL_41_DFFSR_191 ( );
FILL FILL_42_DFFSR_191 ( );
FILL FILL_43_DFFSR_191 ( );
FILL FILL_44_DFFSR_191 ( );
FILL FILL_45_DFFSR_191 ( );
FILL FILL_46_DFFSR_191 ( );
FILL FILL_47_DFFSR_191 ( );
FILL FILL_48_DFFSR_191 ( );
FILL FILL_49_DFFSR_191 ( );
FILL FILL_50_DFFSR_191 ( );
FILL FILL_0_AOI21X1_30 ( );
FILL FILL_1_AOI21X1_30 ( );
FILL FILL_2_AOI21X1_30 ( );
FILL FILL_3_AOI21X1_30 ( );
FILL FILL_4_AOI21X1_30 ( );
FILL FILL_5_AOI21X1_30 ( );
FILL FILL_6_AOI21X1_30 ( );
FILL FILL_7_AOI21X1_30 ( );
FILL FILL_8_AOI21X1_30 ( );
FILL FILL_0_DFFSR_125 ( );
FILL FILL_1_DFFSR_125 ( );
FILL FILL_2_DFFSR_125 ( );
FILL FILL_3_DFFSR_125 ( );
FILL FILL_4_DFFSR_125 ( );
FILL FILL_5_DFFSR_125 ( );
FILL FILL_6_DFFSR_125 ( );
FILL FILL_7_DFFSR_125 ( );
FILL FILL_8_DFFSR_125 ( );
FILL FILL_9_DFFSR_125 ( );
FILL FILL_10_DFFSR_125 ( );
FILL FILL_11_DFFSR_125 ( );
FILL FILL_12_DFFSR_125 ( );
FILL FILL_13_DFFSR_125 ( );
FILL FILL_14_DFFSR_125 ( );
FILL FILL_15_DFFSR_125 ( );
FILL FILL_16_DFFSR_125 ( );
FILL FILL_17_DFFSR_125 ( );
FILL FILL_18_DFFSR_125 ( );
FILL FILL_19_DFFSR_125 ( );
FILL FILL_20_DFFSR_125 ( );
FILL FILL_21_DFFSR_125 ( );
FILL FILL_22_DFFSR_125 ( );
FILL FILL_23_DFFSR_125 ( );
FILL FILL_24_DFFSR_125 ( );
FILL FILL_25_DFFSR_125 ( );
FILL FILL_26_DFFSR_125 ( );
FILL FILL_27_DFFSR_125 ( );
FILL FILL_28_DFFSR_125 ( );
FILL FILL_29_DFFSR_125 ( );
FILL FILL_30_DFFSR_125 ( );
FILL FILL_31_DFFSR_125 ( );
FILL FILL_32_DFFSR_125 ( );
FILL FILL_33_DFFSR_125 ( );
FILL FILL_34_DFFSR_125 ( );
FILL FILL_35_DFFSR_125 ( );
FILL FILL_36_DFFSR_125 ( );
FILL FILL_37_DFFSR_125 ( );
FILL FILL_38_DFFSR_125 ( );
FILL FILL_39_DFFSR_125 ( );
FILL FILL_40_DFFSR_125 ( );
FILL FILL_41_DFFSR_125 ( );
FILL FILL_42_DFFSR_125 ( );
FILL FILL_43_DFFSR_125 ( );
FILL FILL_44_DFFSR_125 ( );
FILL FILL_45_DFFSR_125 ( );
FILL FILL_46_DFFSR_125 ( );
FILL FILL_47_DFFSR_125 ( );
FILL FILL_48_DFFSR_125 ( );
FILL FILL_49_DFFSR_125 ( );
FILL FILL_50_DFFSR_125 ( );
FILL FILL_51_DFFSR_125 ( );
FILL FILL_0_INVX1_139 ( );
FILL FILL_1_INVX1_139 ( );
FILL FILL_2_INVX1_139 ( );
FILL FILL_3_INVX1_139 ( );
FILL FILL_4_INVX1_139 ( );
FILL FILL_0_DFFSR_91 ( );
FILL FILL_1_DFFSR_91 ( );
FILL FILL_2_DFFSR_91 ( );
FILL FILL_3_DFFSR_91 ( );
FILL FILL_4_DFFSR_91 ( );
FILL FILL_5_DFFSR_91 ( );
FILL FILL_6_DFFSR_91 ( );
FILL FILL_7_DFFSR_91 ( );
FILL FILL_8_DFFSR_91 ( );
FILL FILL_9_DFFSR_91 ( );
FILL FILL_10_DFFSR_91 ( );
FILL FILL_11_DFFSR_91 ( );
FILL FILL_12_DFFSR_91 ( );
FILL FILL_13_DFFSR_91 ( );
FILL FILL_14_DFFSR_91 ( );
FILL FILL_15_DFFSR_91 ( );
FILL FILL_16_DFFSR_91 ( );
FILL FILL_17_DFFSR_91 ( );
FILL FILL_18_DFFSR_91 ( );
FILL FILL_19_DFFSR_91 ( );
FILL FILL_20_DFFSR_91 ( );
FILL FILL_21_DFFSR_91 ( );
FILL FILL_22_DFFSR_91 ( );
FILL FILL_23_DFFSR_91 ( );
FILL FILL_24_DFFSR_91 ( );
FILL FILL_25_DFFSR_91 ( );
FILL FILL_26_DFFSR_91 ( );
FILL FILL_27_DFFSR_91 ( );
FILL FILL_28_DFFSR_91 ( );
FILL FILL_29_DFFSR_91 ( );
FILL FILL_30_DFFSR_91 ( );
FILL FILL_31_DFFSR_91 ( );
FILL FILL_32_DFFSR_91 ( );
FILL FILL_33_DFFSR_91 ( );
FILL FILL_34_DFFSR_91 ( );
FILL FILL_35_DFFSR_91 ( );
FILL FILL_36_DFFSR_91 ( );
FILL FILL_37_DFFSR_91 ( );
FILL FILL_38_DFFSR_91 ( );
FILL FILL_39_DFFSR_91 ( );
FILL FILL_40_DFFSR_91 ( );
FILL FILL_41_DFFSR_91 ( );
FILL FILL_42_DFFSR_91 ( );
FILL FILL_43_DFFSR_91 ( );
FILL FILL_44_DFFSR_91 ( );
FILL FILL_45_DFFSR_91 ( );
FILL FILL_46_DFFSR_91 ( );
FILL FILL_47_DFFSR_91 ( );
FILL FILL_48_DFFSR_91 ( );
FILL FILL_49_DFFSR_91 ( );
FILL FILL_50_DFFSR_91 ( );
FILL FILL_51_DFFSR_91 ( );
FILL FILL_0_INVX1_170 ( );
FILL FILL_1_INVX1_170 ( );
FILL FILL_2_INVX1_170 ( );
FILL FILL_3_INVX1_170 ( );
FILL FILL_4_INVX1_170 ( );
FILL FILL_0_DFFSR_157 ( );
FILL FILL_1_DFFSR_157 ( );
FILL FILL_2_DFFSR_157 ( );
FILL FILL_3_DFFSR_157 ( );
FILL FILL_4_DFFSR_157 ( );
FILL FILL_5_DFFSR_157 ( );
FILL FILL_6_DFFSR_157 ( );
FILL FILL_7_DFFSR_157 ( );
FILL FILL_8_DFFSR_157 ( );
FILL FILL_9_DFFSR_157 ( );
FILL FILL_10_DFFSR_157 ( );
FILL FILL_11_DFFSR_157 ( );
FILL FILL_12_DFFSR_157 ( );
FILL FILL_13_DFFSR_157 ( );
FILL FILL_14_DFFSR_157 ( );
FILL FILL_15_DFFSR_157 ( );
FILL FILL_16_DFFSR_157 ( );
FILL FILL_17_DFFSR_157 ( );
FILL FILL_18_DFFSR_157 ( );
FILL FILL_19_DFFSR_157 ( );
FILL FILL_20_DFFSR_157 ( );
FILL FILL_21_DFFSR_157 ( );
FILL FILL_22_DFFSR_157 ( );
FILL FILL_23_DFFSR_157 ( );
FILL FILL_24_DFFSR_157 ( );
FILL FILL_25_DFFSR_157 ( );
FILL FILL_26_DFFSR_157 ( );
FILL FILL_27_DFFSR_157 ( );
FILL FILL_28_DFFSR_157 ( );
FILL FILL_29_DFFSR_157 ( );
FILL FILL_30_DFFSR_157 ( );
FILL FILL_31_DFFSR_157 ( );
FILL FILL_32_DFFSR_157 ( );
FILL FILL_33_DFFSR_157 ( );
FILL FILL_34_DFFSR_157 ( );
FILL FILL_35_DFFSR_157 ( );
FILL FILL_36_DFFSR_157 ( );
FILL FILL_37_DFFSR_157 ( );
FILL FILL_38_DFFSR_157 ( );
FILL FILL_39_DFFSR_157 ( );
FILL FILL_40_DFFSR_157 ( );
FILL FILL_41_DFFSR_157 ( );
FILL FILL_42_DFFSR_157 ( );
FILL FILL_43_DFFSR_157 ( );
FILL FILL_44_DFFSR_157 ( );
FILL FILL_45_DFFSR_157 ( );
FILL FILL_46_DFFSR_157 ( );
FILL FILL_47_DFFSR_157 ( );
FILL FILL_48_DFFSR_157 ( );
FILL FILL_49_DFFSR_157 ( );
FILL FILL_50_DFFSR_157 ( );
FILL FILL_0_NAND2X1_145 ( );
FILL FILL_1_NAND2X1_145 ( );
FILL FILL_2_NAND2X1_145 ( );
FILL FILL_3_NAND2X1_145 ( );
FILL FILL_4_NAND2X1_145 ( );
FILL FILL_5_NAND2X1_145 ( );
FILL FILL_6_NAND2X1_145 ( );
FILL FILL_0_NOR2X1_44 ( );
FILL FILL_1_NOR2X1_44 ( );
FILL FILL_2_NOR2X1_44 ( );
FILL FILL_3_NOR2X1_44 ( );
FILL FILL_4_NOR2X1_44 ( );
FILL FILL_5_NOR2X1_44 ( );
FILL FILL_6_NOR2X1_44 ( );
FILL FILL_0_DFFPOSX1_13 ( );
FILL FILL_1_DFFPOSX1_13 ( );
FILL FILL_2_DFFPOSX1_13 ( );
FILL FILL_3_DFFPOSX1_13 ( );
FILL FILL_4_DFFPOSX1_13 ( );
FILL FILL_5_DFFPOSX1_13 ( );
FILL FILL_6_DFFPOSX1_13 ( );
FILL FILL_7_DFFPOSX1_13 ( );
FILL FILL_8_DFFPOSX1_13 ( );
FILL FILL_9_DFFPOSX1_13 ( );
FILL FILL_10_DFFPOSX1_13 ( );
FILL FILL_11_DFFPOSX1_13 ( );
FILL FILL_12_DFFPOSX1_13 ( );
FILL FILL_13_DFFPOSX1_13 ( );
FILL FILL_14_DFFPOSX1_13 ( );
FILL FILL_15_DFFPOSX1_13 ( );
FILL FILL_16_DFFPOSX1_13 ( );
FILL FILL_17_DFFPOSX1_13 ( );
FILL FILL_18_DFFPOSX1_13 ( );
FILL FILL_19_DFFPOSX1_13 ( );
FILL FILL_20_DFFPOSX1_13 ( );
FILL FILL_21_DFFPOSX1_13 ( );
FILL FILL_22_DFFPOSX1_13 ( );
FILL FILL_23_DFFPOSX1_13 ( );
FILL FILL_24_DFFPOSX1_13 ( );
FILL FILL_25_DFFPOSX1_13 ( );
FILL FILL_26_DFFPOSX1_13 ( );
FILL FILL_27_DFFPOSX1_13 ( );
FILL FILL_0_DFFPOSX1_16 ( );
FILL FILL_1_DFFPOSX1_16 ( );
FILL FILL_2_DFFPOSX1_16 ( );
FILL FILL_3_DFFPOSX1_16 ( );
FILL FILL_4_DFFPOSX1_16 ( );
FILL FILL_5_DFFPOSX1_16 ( );
FILL FILL_6_DFFPOSX1_16 ( );
FILL FILL_7_DFFPOSX1_16 ( );
FILL FILL_8_DFFPOSX1_16 ( );
FILL FILL_9_DFFPOSX1_16 ( );
FILL FILL_10_DFFPOSX1_16 ( );
FILL FILL_11_DFFPOSX1_16 ( );
FILL FILL_12_DFFPOSX1_16 ( );
FILL FILL_13_DFFPOSX1_16 ( );
FILL FILL_14_DFFPOSX1_16 ( );
FILL FILL_15_DFFPOSX1_16 ( );
FILL FILL_16_DFFPOSX1_16 ( );
FILL FILL_17_DFFPOSX1_16 ( );
FILL FILL_18_DFFPOSX1_16 ( );
FILL FILL_19_DFFPOSX1_16 ( );
FILL FILL_20_DFFPOSX1_16 ( );
FILL FILL_21_DFFPOSX1_16 ( );
FILL FILL_22_DFFPOSX1_16 ( );
FILL FILL_23_DFFPOSX1_16 ( );
FILL FILL_24_DFFPOSX1_16 ( );
FILL FILL_25_DFFPOSX1_16 ( );
FILL FILL_26_DFFPOSX1_16 ( );
FILL FILL_27_DFFPOSX1_16 ( );
FILL FILL_0_OAI21X1_175 ( );
FILL FILL_1_OAI21X1_175 ( );
FILL FILL_2_OAI21X1_175 ( );
FILL FILL_3_OAI21X1_175 ( );
FILL FILL_4_OAI21X1_175 ( );
FILL FILL_5_OAI21X1_175 ( );
FILL FILL_6_OAI21X1_175 ( );
FILL FILL_7_OAI21X1_175 ( );
FILL FILL_8_OAI21X1_175 ( );
FILL FILL_9_OAI21X1_175 ( );
FILL FILL_0_INVX1_210 ( );
FILL FILL_1_INVX1_210 ( );
FILL FILL_2_INVX1_210 ( );
FILL FILL_3_INVX1_210 ( );
FILL FILL_0_DFFSR_173 ( );
FILL FILL_1_DFFSR_173 ( );
FILL FILL_2_DFFSR_173 ( );
FILL FILL_3_DFFSR_173 ( );
FILL FILL_4_DFFSR_173 ( );
FILL FILL_5_DFFSR_173 ( );
FILL FILL_6_DFFSR_173 ( );
FILL FILL_7_DFFSR_173 ( );
FILL FILL_8_DFFSR_173 ( );
FILL FILL_9_DFFSR_173 ( );
FILL FILL_10_DFFSR_173 ( );
FILL FILL_11_DFFSR_173 ( );
FILL FILL_12_DFFSR_173 ( );
FILL FILL_13_DFFSR_173 ( );
FILL FILL_14_DFFSR_173 ( );
FILL FILL_15_DFFSR_173 ( );
FILL FILL_16_DFFSR_173 ( );
FILL FILL_17_DFFSR_173 ( );
FILL FILL_18_DFFSR_173 ( );
FILL FILL_19_DFFSR_173 ( );
FILL FILL_20_DFFSR_173 ( );
FILL FILL_21_DFFSR_173 ( );
FILL FILL_22_DFFSR_173 ( );
FILL FILL_23_DFFSR_173 ( );
FILL FILL_24_DFFSR_173 ( );
FILL FILL_25_DFFSR_173 ( );
FILL FILL_26_DFFSR_173 ( );
FILL FILL_27_DFFSR_173 ( );
FILL FILL_28_DFFSR_173 ( );
FILL FILL_29_DFFSR_173 ( );
FILL FILL_30_DFFSR_173 ( );
FILL FILL_31_DFFSR_173 ( );
FILL FILL_32_DFFSR_173 ( );
FILL FILL_33_DFFSR_173 ( );
FILL FILL_34_DFFSR_173 ( );
FILL FILL_35_DFFSR_173 ( );
FILL FILL_36_DFFSR_173 ( );
FILL FILL_37_DFFSR_173 ( );
FILL FILL_38_DFFSR_173 ( );
FILL FILL_39_DFFSR_173 ( );
FILL FILL_40_DFFSR_173 ( );
FILL FILL_41_DFFSR_173 ( );
FILL FILL_42_DFFSR_173 ( );
FILL FILL_43_DFFSR_173 ( );
FILL FILL_44_DFFSR_173 ( );
FILL FILL_45_DFFSR_173 ( );
FILL FILL_46_DFFSR_173 ( );
FILL FILL_47_DFFSR_173 ( );
FILL FILL_48_DFFSR_173 ( );
FILL FILL_49_DFFSR_173 ( );
FILL FILL_50_DFFSR_173 ( );
FILL FILL_0_NAND2X1_211 ( );
FILL FILL_1_NAND2X1_211 ( );
FILL FILL_2_NAND2X1_211 ( );
FILL FILL_3_NAND2X1_211 ( );
FILL FILL_4_NAND2X1_211 ( );
FILL FILL_5_NAND2X1_211 ( );
FILL FILL_6_NAND2X1_211 ( );
FILL FILL_0_NAND2X1_227 ( );
FILL FILL_1_NAND2X1_227 ( );
FILL FILL_2_NAND2X1_227 ( );
FILL FILL_3_NAND2X1_227 ( );
FILL FILL_4_NAND2X1_227 ( );
FILL FILL_5_NAND2X1_227 ( );
FILL FILL_6_NAND2X1_227 ( );
FILL FILL_0_XNOR2X1_3 ( );
FILL FILL_1_XNOR2X1_3 ( );
FILL FILL_2_XNOR2X1_3 ( );
FILL FILL_3_XNOR2X1_3 ( );
FILL FILL_4_XNOR2X1_3 ( );
FILL FILL_5_XNOR2X1_3 ( );
FILL FILL_6_XNOR2X1_3 ( );
FILL FILL_7_XNOR2X1_3 ( );
FILL FILL_8_XNOR2X1_3 ( );
FILL FILL_9_XNOR2X1_3 ( );
FILL FILL_10_XNOR2X1_3 ( );
FILL FILL_11_XNOR2X1_3 ( );
FILL FILL_12_XNOR2X1_3 ( );
FILL FILL_13_XNOR2X1_3 ( );
FILL FILL_14_XNOR2X1_3 ( );
FILL FILL_15_XNOR2X1_3 ( );
FILL FILL_0_INVX1_247 ( );
FILL FILL_1_INVX1_247 ( );
FILL FILL_2_INVX1_247 ( );
FILL FILL_3_INVX1_247 ( );
FILL FILL_4_INVX1_247 ( );
FILL FILL_0_AOI22X1_10 ( );
FILL FILL_1_AOI22X1_10 ( );
FILL FILL_2_AOI22X1_10 ( );
FILL FILL_3_AOI22X1_10 ( );
FILL FILL_4_AOI22X1_10 ( );
FILL FILL_5_AOI22X1_10 ( );
FILL FILL_6_AOI22X1_10 ( );
FILL FILL_7_AOI22X1_10 ( );
FILL FILL_8_AOI22X1_10 ( );
FILL FILL_9_AOI22X1_10 ( );
FILL FILL_10_AOI22X1_10 ( );
FILL FILL_11_AOI22X1_10 ( );
FILL FILL_0_AOI22X1_12 ( );
FILL FILL_1_AOI22X1_12 ( );
FILL FILL_2_AOI22X1_12 ( );
FILL FILL_3_AOI22X1_12 ( );
FILL FILL_4_AOI22X1_12 ( );
FILL FILL_5_AOI22X1_12 ( );
FILL FILL_6_AOI22X1_12 ( );
FILL FILL_7_AOI22X1_12 ( );
FILL FILL_8_AOI22X1_12 ( );
FILL FILL_9_AOI22X1_12 ( );
FILL FILL_10_AOI22X1_12 ( );
FILL FILL_11_AOI22X1_12 ( );
FILL FILL_0_INVX1_255 ( );
FILL FILL_1_INVX1_255 ( );
FILL FILL_2_INVX1_255 ( );
FILL FILL_3_INVX1_255 ( );
FILL FILL_4_INVX1_255 ( );
FILL FILL_0_OAI21X1_223 ( );
FILL FILL_1_OAI21X1_223 ( );
FILL FILL_2_OAI21X1_223 ( );
FILL FILL_3_OAI21X1_223 ( );
FILL FILL_4_OAI21X1_223 ( );
FILL FILL_5_OAI21X1_223 ( );
FILL FILL_6_OAI21X1_223 ( );
FILL FILL_7_OAI21X1_223 ( );
FILL FILL_8_OAI21X1_223 ( );
FILL FILL_9_OAI21X1_223 ( );
FILL FILL_0_OAI21X1_225 ( );
FILL FILL_1_OAI21X1_225 ( );
FILL FILL_2_OAI21X1_225 ( );
FILL FILL_3_OAI21X1_225 ( );
FILL FILL_4_OAI21X1_225 ( );
FILL FILL_5_OAI21X1_225 ( );
FILL FILL_6_OAI21X1_225 ( );
FILL FILL_7_OAI21X1_225 ( );
FILL FILL_8_OAI21X1_225 ( );
FILL FILL_0_OAI21X1_226 ( );
FILL FILL_1_OAI21X1_226 ( );
FILL FILL_2_OAI21X1_226 ( );
FILL FILL_3_OAI21X1_226 ( );
FILL FILL_4_OAI21X1_226 ( );
FILL FILL_5_OAI21X1_226 ( );
FILL FILL_6_OAI21X1_226 ( );
FILL FILL_7_OAI21X1_226 ( );
FILL FILL_8_OAI21X1_226 ( );
FILL FILL_9_OAI21X1_226 ( );
FILL FILL_0_OAI21X1_224 ( );
FILL FILL_1_OAI21X1_224 ( );
FILL FILL_2_OAI21X1_224 ( );
FILL FILL_3_OAI21X1_224 ( );
FILL FILL_4_OAI21X1_224 ( );
FILL FILL_5_OAI21X1_224 ( );
FILL FILL_6_OAI21X1_224 ( );
FILL FILL_7_OAI21X1_224 ( );
FILL FILL_8_OAI21X1_224 ( );
FILL FILL_9_OAI21X1_224 ( );
FILL FILL_0_OR2X2_2 ( );
FILL FILL_1_OR2X2_2 ( );
FILL FILL_2_OR2X2_2 ( );
FILL FILL_3_OR2X2_2 ( );
FILL FILL_4_OR2X2_2 ( );
FILL FILL_5_OR2X2_2 ( );
FILL FILL_6_OR2X2_2 ( );
FILL FILL_7_OR2X2_2 ( );
FILL FILL_8_OR2X2_2 ( );
FILL FILL_0_NAND3X1_95 ( );
FILL FILL_1_NAND3X1_95 ( );
FILL FILL_2_NAND3X1_95 ( );
FILL FILL_3_NAND3X1_95 ( );
FILL FILL_4_NAND3X1_95 ( );
FILL FILL_5_NAND3X1_95 ( );
FILL FILL_6_NAND3X1_95 ( );
FILL FILL_7_NAND3X1_95 ( );
FILL FILL_8_NAND3X1_95 ( );
FILL FILL_0_OAI21X1_234 ( );
FILL FILL_1_OAI21X1_234 ( );
FILL FILL_2_OAI21X1_234 ( );
FILL FILL_3_OAI21X1_234 ( );
FILL FILL_4_OAI21X1_234 ( );
FILL FILL_5_OAI21X1_234 ( );
FILL FILL_6_OAI21X1_234 ( );
FILL FILL_7_OAI21X1_234 ( );
FILL FILL_8_OAI21X1_234 ( );
FILL FILL_9_OAI21X1_234 ( );
FILL FILL_0_OAI21X1_235 ( );
FILL FILL_1_OAI21X1_235 ( );
FILL FILL_2_OAI21X1_235 ( );
FILL FILL_3_OAI21X1_235 ( );
FILL FILL_4_OAI21X1_235 ( );
FILL FILL_5_OAI21X1_235 ( );
FILL FILL_6_OAI21X1_235 ( );
FILL FILL_7_OAI21X1_235 ( );
FILL FILL_8_OAI21X1_235 ( );
FILL FILL_0_INVX1_119 ( );
FILL FILL_1_INVX1_119 ( );
FILL FILL_2_INVX1_119 ( );
FILL FILL_3_INVX1_119 ( );
FILL FILL_4_INVX1_119 ( );
FILL FILL_0_OAI21X1_105 ( );
FILL FILL_1_OAI21X1_105 ( );
FILL FILL_2_OAI21X1_105 ( );
FILL FILL_3_OAI21X1_105 ( );
FILL FILL_4_OAI21X1_105 ( );
FILL FILL_5_OAI21X1_105 ( );
FILL FILL_6_OAI21X1_105 ( );
FILL FILL_7_OAI21X1_105 ( );
FILL FILL_8_OAI21X1_105 ( );
FILL FILL_0_DFFSR_109 ( );
FILL FILL_1_DFFSR_109 ( );
FILL FILL_2_DFFSR_109 ( );
FILL FILL_3_DFFSR_109 ( );
FILL FILL_4_DFFSR_109 ( );
FILL FILL_5_DFFSR_109 ( );
FILL FILL_6_DFFSR_109 ( );
FILL FILL_7_DFFSR_109 ( );
FILL FILL_8_DFFSR_109 ( );
FILL FILL_9_DFFSR_109 ( );
FILL FILL_10_DFFSR_109 ( );
FILL FILL_11_DFFSR_109 ( );
FILL FILL_12_DFFSR_109 ( );
FILL FILL_13_DFFSR_109 ( );
FILL FILL_14_DFFSR_109 ( );
FILL FILL_15_DFFSR_109 ( );
FILL FILL_16_DFFSR_109 ( );
FILL FILL_17_DFFSR_109 ( );
FILL FILL_18_DFFSR_109 ( );
FILL FILL_19_DFFSR_109 ( );
FILL FILL_20_DFFSR_109 ( );
FILL FILL_21_DFFSR_109 ( );
FILL FILL_22_DFFSR_109 ( );
FILL FILL_23_DFFSR_109 ( );
FILL FILL_24_DFFSR_109 ( );
FILL FILL_25_DFFSR_109 ( );
FILL FILL_26_DFFSR_109 ( );
FILL FILL_27_DFFSR_109 ( );
FILL FILL_28_DFFSR_109 ( );
FILL FILL_29_DFFSR_109 ( );
FILL FILL_30_DFFSR_109 ( );
FILL FILL_31_DFFSR_109 ( );
FILL FILL_32_DFFSR_109 ( );
FILL FILL_33_DFFSR_109 ( );
FILL FILL_34_DFFSR_109 ( );
FILL FILL_35_DFFSR_109 ( );
FILL FILL_36_DFFSR_109 ( );
FILL FILL_37_DFFSR_109 ( );
FILL FILL_38_DFFSR_109 ( );
FILL FILL_39_DFFSR_109 ( );
FILL FILL_40_DFFSR_109 ( );
FILL FILL_41_DFFSR_109 ( );
FILL FILL_42_DFFSR_109 ( );
FILL FILL_43_DFFSR_109 ( );
FILL FILL_44_DFFSR_109 ( );
FILL FILL_45_DFFSR_109 ( );
FILL FILL_46_DFFSR_109 ( );
FILL FILL_47_DFFSR_109 ( );
FILL FILL_48_DFFSR_109 ( );
FILL FILL_49_DFFSR_109 ( );
FILL FILL_50_DFFSR_109 ( );
FILL FILL_0_NAND2X1_100 ( );
FILL FILL_1_NAND2X1_100 ( );
FILL FILL_2_NAND2X1_100 ( );
FILL FILL_3_NAND2X1_100 ( );
FILL FILL_4_NAND2X1_100 ( );
FILL FILL_5_NAND2X1_100 ( );
FILL FILL_6_NAND2X1_100 ( );
FILL FILL_0_NAND2X1_123 ( );
FILL FILL_1_NAND2X1_123 ( );
FILL FILL_2_NAND2X1_123 ( );
FILL FILL_3_NAND2X1_123 ( );
FILL FILL_4_NAND2X1_123 ( );
FILL FILL_5_NAND2X1_123 ( );
FILL FILL_6_NAND2X1_123 ( );
FILL FILL_0_DFFSR_115 ( );
FILL FILL_1_DFFSR_115 ( );
FILL FILL_2_DFFSR_115 ( );
FILL FILL_3_DFFSR_115 ( );
FILL FILL_4_DFFSR_115 ( );
FILL FILL_5_DFFSR_115 ( );
FILL FILL_6_DFFSR_115 ( );
FILL FILL_7_DFFSR_115 ( );
FILL FILL_8_DFFSR_115 ( );
FILL FILL_9_DFFSR_115 ( );
FILL FILL_10_DFFSR_115 ( );
FILL FILL_11_DFFSR_115 ( );
FILL FILL_12_DFFSR_115 ( );
FILL FILL_13_DFFSR_115 ( );
FILL FILL_14_DFFSR_115 ( );
FILL FILL_15_DFFSR_115 ( );
FILL FILL_16_DFFSR_115 ( );
FILL FILL_17_DFFSR_115 ( );
FILL FILL_18_DFFSR_115 ( );
FILL FILL_19_DFFSR_115 ( );
FILL FILL_20_DFFSR_115 ( );
FILL FILL_21_DFFSR_115 ( );
FILL FILL_22_DFFSR_115 ( );
FILL FILL_23_DFFSR_115 ( );
FILL FILL_24_DFFSR_115 ( );
FILL FILL_25_DFFSR_115 ( );
FILL FILL_26_DFFSR_115 ( );
FILL FILL_27_DFFSR_115 ( );
FILL FILL_28_DFFSR_115 ( );
FILL FILL_29_DFFSR_115 ( );
FILL FILL_30_DFFSR_115 ( );
FILL FILL_31_DFFSR_115 ( );
FILL FILL_32_DFFSR_115 ( );
FILL FILL_33_DFFSR_115 ( );
FILL FILL_34_DFFSR_115 ( );
FILL FILL_35_DFFSR_115 ( );
FILL FILL_36_DFFSR_115 ( );
FILL FILL_37_DFFSR_115 ( );
FILL FILL_38_DFFSR_115 ( );
FILL FILL_39_DFFSR_115 ( );
FILL FILL_40_DFFSR_115 ( );
FILL FILL_41_DFFSR_115 ( );
FILL FILL_42_DFFSR_115 ( );
FILL FILL_43_DFFSR_115 ( );
FILL FILL_44_DFFSR_115 ( );
FILL FILL_45_DFFSR_115 ( );
FILL FILL_46_DFFSR_115 ( );
FILL FILL_47_DFFSR_115 ( );
FILL FILL_48_DFFSR_115 ( );
FILL FILL_49_DFFSR_115 ( );
FILL FILL_50_DFFSR_115 ( );
FILL FILL_51_DFFSR_115 ( );
FILL FILL_0_OAI21X1_156 ( );
FILL FILL_1_OAI21X1_156 ( );
FILL FILL_2_OAI21X1_156 ( );
FILL FILL_3_OAI21X1_156 ( );
FILL FILL_4_OAI21X1_156 ( );
FILL FILL_5_OAI21X1_156 ( );
FILL FILL_6_OAI21X1_156 ( );
FILL FILL_7_OAI21X1_156 ( );
FILL FILL_8_OAI21X1_156 ( );
FILL FILL_0_INVX1_186 ( );
FILL FILL_1_INVX1_186 ( );
FILL FILL_2_INVX1_186 ( );
FILL FILL_3_INVX1_186 ( );
FILL FILL_4_INVX1_186 ( );
FILL FILL_0_DFFPOSX1_1 ( );
FILL FILL_1_DFFPOSX1_1 ( );
FILL FILL_2_DFFPOSX1_1 ( );
FILL FILL_3_DFFPOSX1_1 ( );
FILL FILL_4_DFFPOSX1_1 ( );
FILL FILL_5_DFFPOSX1_1 ( );
FILL FILL_6_DFFPOSX1_1 ( );
FILL FILL_7_DFFPOSX1_1 ( );
FILL FILL_8_DFFPOSX1_1 ( );
FILL FILL_9_DFFPOSX1_1 ( );
FILL FILL_10_DFFPOSX1_1 ( );
FILL FILL_11_DFFPOSX1_1 ( );
FILL FILL_12_DFFPOSX1_1 ( );
FILL FILL_13_DFFPOSX1_1 ( );
FILL FILL_14_DFFPOSX1_1 ( );
FILL FILL_15_DFFPOSX1_1 ( );
FILL FILL_16_DFFPOSX1_1 ( );
FILL FILL_17_DFFPOSX1_1 ( );
FILL FILL_18_DFFPOSX1_1 ( );
FILL FILL_19_DFFPOSX1_1 ( );
FILL FILL_20_DFFPOSX1_1 ( );
FILL FILL_21_DFFPOSX1_1 ( );
FILL FILL_22_DFFPOSX1_1 ( );
FILL FILL_23_DFFPOSX1_1 ( );
FILL FILL_24_DFFPOSX1_1 ( );
FILL FILL_25_DFFPOSX1_1 ( );
FILL FILL_26_DFFPOSX1_1 ( );
FILL FILL_27_DFFPOSX1_1 ( );
FILL FILL_0_BUFX2_6 ( );
FILL FILL_1_BUFX2_6 ( );
FILL FILL_2_BUFX2_6 ( );
FILL FILL_3_BUFX2_6 ( );
FILL FILL_4_BUFX2_6 ( );
FILL FILL_5_BUFX2_6 ( );
FILL FILL_6_BUFX2_6 ( );
FILL FILL_0_DFFPOSX1_14 ( );
FILL FILL_1_DFFPOSX1_14 ( );
FILL FILL_2_DFFPOSX1_14 ( );
FILL FILL_3_DFFPOSX1_14 ( );
FILL FILL_4_DFFPOSX1_14 ( );
FILL FILL_5_DFFPOSX1_14 ( );
FILL FILL_6_DFFPOSX1_14 ( );
FILL FILL_7_DFFPOSX1_14 ( );
FILL FILL_8_DFFPOSX1_14 ( );
FILL FILL_9_DFFPOSX1_14 ( );
FILL FILL_10_DFFPOSX1_14 ( );
FILL FILL_11_DFFPOSX1_14 ( );
FILL FILL_12_DFFPOSX1_14 ( );
FILL FILL_13_DFFPOSX1_14 ( );
FILL FILL_14_DFFPOSX1_14 ( );
FILL FILL_15_DFFPOSX1_14 ( );
FILL FILL_16_DFFPOSX1_14 ( );
FILL FILL_17_DFFPOSX1_14 ( );
FILL FILL_18_DFFPOSX1_14 ( );
FILL FILL_19_DFFPOSX1_14 ( );
FILL FILL_20_DFFPOSX1_14 ( );
FILL FILL_21_DFFPOSX1_14 ( );
FILL FILL_22_DFFPOSX1_14 ( );
FILL FILL_23_DFFPOSX1_14 ( );
FILL FILL_24_DFFPOSX1_14 ( );
FILL FILL_25_DFFPOSX1_14 ( );
FILL FILL_26_DFFPOSX1_14 ( );
FILL FILL_27_DFFPOSX1_14 ( );
FILL FILL_0_OAI21X1_243 ( );
FILL FILL_1_OAI21X1_243 ( );
FILL FILL_2_OAI21X1_243 ( );
FILL FILL_3_OAI21X1_243 ( );
FILL FILL_4_OAI21X1_243 ( );
FILL FILL_5_OAI21X1_243 ( );
FILL FILL_6_OAI21X1_243 ( );
FILL FILL_7_OAI21X1_243 ( );
FILL FILL_8_OAI21X1_243 ( );
FILL FILL_0_INVX1_402 ( );
FILL FILL_1_INVX1_402 ( );
FILL FILL_2_INVX1_402 ( );
FILL FILL_3_INVX1_402 ( );
FILL FILL_4_INVX1_402 ( );
FILL FILL_0_DFFSR_12 ( );
FILL FILL_1_DFFSR_12 ( );
FILL FILL_2_DFFSR_12 ( );
FILL FILL_3_DFFSR_12 ( );
FILL FILL_4_DFFSR_12 ( );
FILL FILL_5_DFFSR_12 ( );
FILL FILL_6_DFFSR_12 ( );
FILL FILL_7_DFFSR_12 ( );
FILL FILL_8_DFFSR_12 ( );
FILL FILL_9_DFFSR_12 ( );
FILL FILL_10_DFFSR_12 ( );
FILL FILL_11_DFFSR_12 ( );
FILL FILL_12_DFFSR_12 ( );
FILL FILL_13_DFFSR_12 ( );
FILL FILL_14_DFFSR_12 ( );
FILL FILL_15_DFFSR_12 ( );
FILL FILL_16_DFFSR_12 ( );
FILL FILL_17_DFFSR_12 ( );
FILL FILL_18_DFFSR_12 ( );
FILL FILL_19_DFFSR_12 ( );
FILL FILL_20_DFFSR_12 ( );
FILL FILL_21_DFFSR_12 ( );
FILL FILL_22_DFFSR_12 ( );
FILL FILL_23_DFFSR_12 ( );
FILL FILL_24_DFFSR_12 ( );
FILL FILL_25_DFFSR_12 ( );
FILL FILL_26_DFFSR_12 ( );
FILL FILL_27_DFFSR_12 ( );
FILL FILL_28_DFFSR_12 ( );
FILL FILL_29_DFFSR_12 ( );
FILL FILL_30_DFFSR_12 ( );
FILL FILL_31_DFFSR_12 ( );
FILL FILL_32_DFFSR_12 ( );
FILL FILL_33_DFFSR_12 ( );
FILL FILL_34_DFFSR_12 ( );
FILL FILL_35_DFFSR_12 ( );
FILL FILL_36_DFFSR_12 ( );
FILL FILL_37_DFFSR_12 ( );
FILL FILL_38_DFFSR_12 ( );
FILL FILL_39_DFFSR_12 ( );
FILL FILL_40_DFFSR_12 ( );
FILL FILL_41_DFFSR_12 ( );
FILL FILL_42_DFFSR_12 ( );
FILL FILL_43_DFFSR_12 ( );
FILL FILL_44_DFFSR_12 ( );
FILL FILL_45_DFFSR_12 ( );
FILL FILL_46_DFFSR_12 ( );
FILL FILL_47_DFFSR_12 ( );
FILL FILL_48_DFFSR_12 ( );
FILL FILL_49_DFFSR_12 ( );
FILL FILL_50_DFFSR_12 ( );
FILL FILL_51_DFFSR_12 ( );
FILL FILL_0_OAI21X1_173 ( );
FILL FILL_1_OAI21X1_173 ( );
FILL FILL_2_OAI21X1_173 ( );
FILL FILL_3_OAI21X1_173 ( );
FILL FILL_4_OAI21X1_173 ( );
FILL FILL_5_OAI21X1_173 ( );
FILL FILL_6_OAI21X1_173 ( );
FILL FILL_7_OAI21X1_173 ( );
FILL FILL_8_OAI21X1_173 ( );
FILL FILL_9_OAI21X1_173 ( );
FILL FILL_0_INVX1_248 ( );
FILL FILL_1_INVX1_248 ( );
FILL FILL_2_INVX1_248 ( );
FILL FILL_3_INVX1_248 ( );
FILL FILL_4_INVX1_248 ( );
FILL FILL_0_NAND2X1_223 ( );
FILL FILL_1_NAND2X1_223 ( );
FILL FILL_2_NAND2X1_223 ( );
FILL FILL_3_NAND2X1_223 ( );
FILL FILL_4_NAND2X1_223 ( );
FILL FILL_5_NAND2X1_223 ( );
FILL FILL_6_NAND2X1_223 ( );
FILL FILL_0_NAND3X1_66 ( );
FILL FILL_1_NAND3X1_66 ( );
FILL FILL_2_NAND3X1_66 ( );
FILL FILL_3_NAND3X1_66 ( );
FILL FILL_4_NAND3X1_66 ( );
FILL FILL_5_NAND3X1_66 ( );
FILL FILL_6_NAND3X1_66 ( );
FILL FILL_7_NAND3X1_66 ( );
FILL FILL_8_NAND3X1_66 ( );
FILL FILL_0_NAND3X1_67 ( );
FILL FILL_1_NAND3X1_67 ( );
FILL FILL_2_NAND3X1_67 ( );
FILL FILL_3_NAND3X1_67 ( );
FILL FILL_4_NAND3X1_67 ( );
FILL FILL_5_NAND3X1_67 ( );
FILL FILL_6_NAND3X1_67 ( );
FILL FILL_7_NAND3X1_67 ( );
FILL FILL_8_NAND3X1_67 ( );
FILL FILL_0_NAND3X1_69 ( );
FILL FILL_1_NAND3X1_69 ( );
FILL FILL_2_NAND3X1_69 ( );
FILL FILL_3_NAND3X1_69 ( );
FILL FILL_4_NAND3X1_69 ( );
FILL FILL_5_NAND3X1_69 ( );
FILL FILL_6_NAND3X1_69 ( );
FILL FILL_7_NAND3X1_69 ( );
FILL FILL_8_NAND3X1_69 ( );
FILL FILL_9_NAND3X1_69 ( );
FILL FILL_0_AND2X2_9 ( );
FILL FILL_1_AND2X2_9 ( );
FILL FILL_2_AND2X2_9 ( );
FILL FILL_3_AND2X2_9 ( );
FILL FILL_4_AND2X2_9 ( );
FILL FILL_5_AND2X2_9 ( );
FILL FILL_6_AND2X2_9 ( );
FILL FILL_7_AND2X2_9 ( );
FILL FILL_8_AND2X2_9 ( );
FILL FILL_9_AND2X2_9 ( );
FILL FILL_0_NAND2X1_200 ( );
FILL FILL_1_NAND2X1_200 ( );
FILL FILL_2_NAND2X1_200 ( );
FILL FILL_3_NAND2X1_200 ( );
FILL FILL_4_NAND2X1_200 ( );
FILL FILL_5_NAND2X1_200 ( );
FILL FILL_6_NAND2X1_200 ( );
FILL FILL_0_INVX1_215 ( );
FILL FILL_1_INVX1_215 ( );
FILL FILL_2_INVX1_215 ( );
FILL FILL_3_INVX1_215 ( );
FILL FILL_4_INVX1_215 ( );
FILL FILL_0_DFFSR_165 ( );
FILL FILL_1_DFFSR_165 ( );
FILL FILL_2_DFFSR_165 ( );
FILL FILL_3_DFFSR_165 ( );
FILL FILL_4_DFFSR_165 ( );
FILL FILL_5_DFFSR_165 ( );
FILL FILL_6_DFFSR_165 ( );
FILL FILL_7_DFFSR_165 ( );
FILL FILL_8_DFFSR_165 ( );
FILL FILL_9_DFFSR_165 ( );
FILL FILL_10_DFFSR_165 ( );
FILL FILL_11_DFFSR_165 ( );
FILL FILL_12_DFFSR_165 ( );
FILL FILL_13_DFFSR_165 ( );
FILL FILL_14_DFFSR_165 ( );
FILL FILL_15_DFFSR_165 ( );
FILL FILL_16_DFFSR_165 ( );
FILL FILL_17_DFFSR_165 ( );
FILL FILL_18_DFFSR_165 ( );
FILL FILL_19_DFFSR_165 ( );
FILL FILL_20_DFFSR_165 ( );
FILL FILL_21_DFFSR_165 ( );
FILL FILL_22_DFFSR_165 ( );
FILL FILL_23_DFFSR_165 ( );
FILL FILL_24_DFFSR_165 ( );
FILL FILL_25_DFFSR_165 ( );
FILL FILL_26_DFFSR_165 ( );
FILL FILL_27_DFFSR_165 ( );
FILL FILL_28_DFFSR_165 ( );
FILL FILL_29_DFFSR_165 ( );
FILL FILL_30_DFFSR_165 ( );
FILL FILL_31_DFFSR_165 ( );
FILL FILL_32_DFFSR_165 ( );
FILL FILL_33_DFFSR_165 ( );
FILL FILL_34_DFFSR_165 ( );
FILL FILL_35_DFFSR_165 ( );
FILL FILL_36_DFFSR_165 ( );
FILL FILL_37_DFFSR_165 ( );
FILL FILL_38_DFFSR_165 ( );
FILL FILL_39_DFFSR_165 ( );
FILL FILL_40_DFFSR_165 ( );
FILL FILL_41_DFFSR_165 ( );
FILL FILL_42_DFFSR_165 ( );
FILL FILL_43_DFFSR_165 ( );
FILL FILL_44_DFFSR_165 ( );
FILL FILL_45_DFFSR_165 ( );
FILL FILL_46_DFFSR_165 ( );
FILL FILL_47_DFFSR_165 ( );
FILL FILL_48_DFFSR_165 ( );
FILL FILL_49_DFFSR_165 ( );
FILL FILL_50_DFFSR_165 ( );
FILL FILL_0_NOR2X1_11 ( );
FILL FILL_1_NOR2X1_11 ( );
FILL FILL_2_NOR2X1_11 ( );
FILL FILL_3_NOR2X1_11 ( );
FILL FILL_4_NOR2X1_11 ( );
FILL FILL_5_NOR2X1_11 ( );
FILL FILL_6_NOR2X1_11 ( );
FILL FILL_0_NAND2X1_221 ( );
FILL FILL_1_NAND2X1_221 ( );
FILL FILL_2_NAND2X1_221 ( );
FILL FILL_3_NAND2X1_221 ( );
FILL FILL_4_NAND2X1_221 ( );
FILL FILL_5_NAND2X1_221 ( );
FILL FILL_6_NAND2X1_221 ( );
FILL FILL_0_INVX1_254 ( );
FILL FILL_1_INVX1_254 ( );
FILL FILL_2_INVX1_254 ( );
FILL FILL_3_INVX1_254 ( );
FILL FILL_4_INVX1_254 ( );
FILL FILL_0_NAND3X1_99 ( );
FILL FILL_1_NAND3X1_99 ( );
FILL FILL_2_NAND3X1_99 ( );
FILL FILL_3_NAND3X1_99 ( );
FILL FILL_4_NAND3X1_99 ( );
FILL FILL_5_NAND3X1_99 ( );
FILL FILL_6_NAND3X1_99 ( );
FILL FILL_7_NAND3X1_99 ( );
FILL FILL_8_NAND3X1_99 ( );
FILL FILL_9_NAND3X1_99 ( );
FILL FILL_0_NAND3X1_100 ( );
FILL FILL_1_NAND3X1_100 ( );
FILL FILL_2_NAND3X1_100 ( );
FILL FILL_3_NAND3X1_100 ( );
FILL FILL_4_NAND3X1_100 ( );
FILL FILL_5_NAND3X1_100 ( );
FILL FILL_6_NAND3X1_100 ( );
FILL FILL_7_NAND3X1_100 ( );
FILL FILL_8_NAND3X1_100 ( );
FILL FILL_0_NAND3X1_105 ( );
FILL FILL_1_NAND3X1_105 ( );
FILL FILL_2_NAND3X1_105 ( );
FILL FILL_3_NAND3X1_105 ( );
FILL FILL_4_NAND3X1_105 ( );
FILL FILL_5_NAND3X1_105 ( );
FILL FILL_6_NAND3X1_105 ( );
FILL FILL_7_NAND3X1_105 ( );
FILL FILL_8_NAND3X1_105 ( );
FILL FILL_0_NAND2X1_105 ( );
FILL FILL_1_NAND2X1_105 ( );
FILL FILL_2_NAND2X1_105 ( );
FILL FILL_3_NAND2X1_105 ( );
FILL FILL_4_NAND2X1_105 ( );
FILL FILL_5_NAND2X1_105 ( );
FILL FILL_6_NAND2X1_105 ( );
FILL FILL_0_OAI21X1_89 ( );
FILL FILL_1_OAI21X1_89 ( );
FILL FILL_2_OAI21X1_89 ( );
FILL FILL_3_OAI21X1_89 ( );
FILL FILL_4_OAI21X1_89 ( );
FILL FILL_5_OAI21X1_89 ( );
FILL FILL_6_OAI21X1_89 ( );
FILL FILL_7_OAI21X1_89 ( );
FILL FILL_8_OAI21X1_89 ( );
FILL FILL_0_INVX1_101 ( );
FILL FILL_1_INVX1_101 ( );
FILL FILL_2_INVX1_101 ( );
FILL FILL_3_INVX1_101 ( );
FILL FILL_4_INVX1_101 ( );
FILL FILL_0_OAI21X1_125 ( );
FILL FILL_1_OAI21X1_125 ( );
FILL FILL_2_OAI21X1_125 ( );
FILL FILL_3_OAI21X1_125 ( );
FILL FILL_4_OAI21X1_125 ( );
FILL FILL_5_OAI21X1_125 ( );
FILL FILL_6_OAI21X1_125 ( );
FILL FILL_7_OAI21X1_125 ( );
FILL FILL_8_OAI21X1_125 ( );
FILL FILL_0_INVX1_141 ( );
FILL FILL_1_INVX1_141 ( );
FILL FILL_2_INVX1_141 ( );
FILL FILL_3_INVX1_141 ( );
FILL FILL_4_INVX1_141 ( );
FILL FILL_0_NAND2X1_125 ( );
FILL FILL_1_NAND2X1_125 ( );
FILL FILL_2_NAND2X1_125 ( );
FILL FILL_3_NAND2X1_125 ( );
FILL FILL_4_NAND2X1_125 ( );
FILL FILL_5_NAND2X1_125 ( );
FILL FILL_6_NAND2X1_125 ( );
FILL FILL_0_NAND2X1_117 ( );
FILL FILL_1_NAND2X1_117 ( );
FILL FILL_2_NAND2X1_117 ( );
FILL FILL_3_NAND2X1_117 ( );
FILL FILL_4_NAND2X1_117 ( );
FILL FILL_5_NAND2X1_117 ( );
FILL FILL_6_NAND2X1_117 ( );
FILL FILL_0_DFFSR_68 ( );
FILL FILL_1_DFFSR_68 ( );
FILL FILL_2_DFFSR_68 ( );
FILL FILL_3_DFFSR_68 ( );
FILL FILL_4_DFFSR_68 ( );
FILL FILL_5_DFFSR_68 ( );
FILL FILL_6_DFFSR_68 ( );
FILL FILL_7_DFFSR_68 ( );
FILL FILL_8_DFFSR_68 ( );
FILL FILL_9_DFFSR_68 ( );
FILL FILL_10_DFFSR_68 ( );
FILL FILL_11_DFFSR_68 ( );
FILL FILL_12_DFFSR_68 ( );
FILL FILL_13_DFFSR_68 ( );
FILL FILL_14_DFFSR_68 ( );
FILL FILL_15_DFFSR_68 ( );
FILL FILL_16_DFFSR_68 ( );
FILL FILL_17_DFFSR_68 ( );
FILL FILL_18_DFFSR_68 ( );
FILL FILL_19_DFFSR_68 ( );
FILL FILL_20_DFFSR_68 ( );
FILL FILL_21_DFFSR_68 ( );
FILL FILL_22_DFFSR_68 ( );
FILL FILL_23_DFFSR_68 ( );
FILL FILL_24_DFFSR_68 ( );
FILL FILL_25_DFFSR_68 ( );
FILL FILL_26_DFFSR_68 ( );
FILL FILL_27_DFFSR_68 ( );
FILL FILL_28_DFFSR_68 ( );
FILL FILL_29_DFFSR_68 ( );
FILL FILL_30_DFFSR_68 ( );
FILL FILL_31_DFFSR_68 ( );
FILL FILL_32_DFFSR_68 ( );
FILL FILL_33_DFFSR_68 ( );
FILL FILL_34_DFFSR_68 ( );
FILL FILL_35_DFFSR_68 ( );
FILL FILL_36_DFFSR_68 ( );
FILL FILL_37_DFFSR_68 ( );
FILL FILL_38_DFFSR_68 ( );
FILL FILL_39_DFFSR_68 ( );
FILL FILL_40_DFFSR_68 ( );
FILL FILL_41_DFFSR_68 ( );
FILL FILL_42_DFFSR_68 ( );
FILL FILL_43_DFFSR_68 ( );
FILL FILL_44_DFFSR_68 ( );
FILL FILL_45_DFFSR_68 ( );
FILL FILL_46_DFFSR_68 ( );
FILL FILL_47_DFFSR_68 ( );
FILL FILL_48_DFFSR_68 ( );
FILL FILL_49_DFFSR_68 ( );
FILL FILL_50_DFFSR_68 ( );
FILL FILL_0_INVX1_173 ( );
FILL FILL_1_INVX1_173 ( );
FILL FILL_2_INVX1_173 ( );
FILL FILL_3_INVX1_173 ( );
FILL FILL_4_INVX1_173 ( );
FILL FILL_0_INVX1_171 ( );
FILL FILL_1_INVX1_171 ( );
FILL FILL_2_INVX1_171 ( );
FILL FILL_3_INVX1_171 ( );
FILL FILL_4_INVX1_171 ( );
FILL FILL_0_INVX1_189 ( );
FILL FILL_1_INVX1_189 ( );
FILL FILL_2_INVX1_189 ( );
FILL FILL_3_INVX1_189 ( );
FILL FILL_4_INVX1_189 ( );
FILL FILL_0_DFFSR_14 ( );
FILL FILL_1_DFFSR_14 ( );
FILL FILL_2_DFFSR_14 ( );
FILL FILL_3_DFFSR_14 ( );
FILL FILL_4_DFFSR_14 ( );
FILL FILL_5_DFFSR_14 ( );
FILL FILL_6_DFFSR_14 ( );
FILL FILL_7_DFFSR_14 ( );
FILL FILL_8_DFFSR_14 ( );
FILL FILL_9_DFFSR_14 ( );
FILL FILL_10_DFFSR_14 ( );
FILL FILL_11_DFFSR_14 ( );
FILL FILL_12_DFFSR_14 ( );
FILL FILL_13_DFFSR_14 ( );
FILL FILL_14_DFFSR_14 ( );
FILL FILL_15_DFFSR_14 ( );
FILL FILL_16_DFFSR_14 ( );
FILL FILL_17_DFFSR_14 ( );
FILL FILL_18_DFFSR_14 ( );
FILL FILL_19_DFFSR_14 ( );
FILL FILL_20_DFFSR_14 ( );
FILL FILL_21_DFFSR_14 ( );
FILL FILL_22_DFFSR_14 ( );
FILL FILL_23_DFFSR_14 ( );
FILL FILL_24_DFFSR_14 ( );
FILL FILL_25_DFFSR_14 ( );
FILL FILL_26_DFFSR_14 ( );
FILL FILL_27_DFFSR_14 ( );
FILL FILL_28_DFFSR_14 ( );
FILL FILL_29_DFFSR_14 ( );
FILL FILL_30_DFFSR_14 ( );
FILL FILL_31_DFFSR_14 ( );
FILL FILL_32_DFFSR_14 ( );
FILL FILL_33_DFFSR_14 ( );
FILL FILL_34_DFFSR_14 ( );
FILL FILL_35_DFFSR_14 ( );
FILL FILL_36_DFFSR_14 ( );
FILL FILL_37_DFFSR_14 ( );
FILL FILL_38_DFFSR_14 ( );
FILL FILL_39_DFFSR_14 ( );
FILL FILL_40_DFFSR_14 ( );
FILL FILL_41_DFFSR_14 ( );
FILL FILL_42_DFFSR_14 ( );
FILL FILL_43_DFFSR_14 ( );
FILL FILL_44_DFFSR_14 ( );
FILL FILL_45_DFFSR_14 ( );
FILL FILL_46_DFFSR_14 ( );
FILL FILL_47_DFFSR_14 ( );
FILL FILL_48_DFFSR_14 ( );
FILL FILL_49_DFFSR_14 ( );
FILL FILL_50_DFFSR_14 ( );
FILL FILL_0_NAND3X1_129 ( );
FILL FILL_1_NAND3X1_129 ( );
FILL FILL_2_NAND3X1_129 ( );
FILL FILL_3_NAND3X1_129 ( );
FILL FILL_4_NAND3X1_129 ( );
FILL FILL_5_NAND3X1_129 ( );
FILL FILL_6_NAND3X1_129 ( );
FILL FILL_7_NAND3X1_129 ( );
FILL FILL_8_NAND3X1_129 ( );
FILL FILL_0_NOR2X1_45 ( );
FILL FILL_1_NOR2X1_45 ( );
FILL FILL_2_NOR2X1_45 ( );
FILL FILL_3_NOR2X1_45 ( );
FILL FILL_4_NOR2X1_45 ( );
FILL FILL_5_NOR2X1_45 ( );
FILL FILL_6_NOR2X1_45 ( );
FILL FILL_0_INVX1_401 ( );
FILL FILL_1_INVX1_401 ( );
FILL FILL_2_INVX1_401 ( );
FILL FILL_3_INVX1_401 ( );
FILL FILL_0_AOI21X1_41 ( );
FILL FILL_1_AOI21X1_41 ( );
FILL FILL_2_AOI21X1_41 ( );
FILL FILL_3_AOI21X1_41 ( );
FILL FILL_4_AOI21X1_41 ( );
FILL FILL_5_AOI21X1_41 ( );
FILL FILL_6_AOI21X1_41 ( );
FILL FILL_7_AOI21X1_41 ( );
FILL FILL_8_AOI21X1_41 ( );
FILL FILL_0_DFFPOSX1_15 ( );
FILL FILL_1_DFFPOSX1_15 ( );
FILL FILL_2_DFFPOSX1_15 ( );
FILL FILL_3_DFFPOSX1_15 ( );
FILL FILL_4_DFFPOSX1_15 ( );
FILL FILL_5_DFFPOSX1_15 ( );
FILL FILL_6_DFFPOSX1_15 ( );
FILL FILL_7_DFFPOSX1_15 ( );
FILL FILL_8_DFFPOSX1_15 ( );
FILL FILL_9_DFFPOSX1_15 ( );
FILL FILL_10_DFFPOSX1_15 ( );
FILL FILL_11_DFFPOSX1_15 ( );
FILL FILL_12_DFFPOSX1_15 ( );
FILL FILL_13_DFFPOSX1_15 ( );
FILL FILL_14_DFFPOSX1_15 ( );
FILL FILL_15_DFFPOSX1_15 ( );
FILL FILL_16_DFFPOSX1_15 ( );
FILL FILL_17_DFFPOSX1_15 ( );
FILL FILL_18_DFFPOSX1_15 ( );
FILL FILL_19_DFFPOSX1_15 ( );
FILL FILL_20_DFFPOSX1_15 ( );
FILL FILL_21_DFFPOSX1_15 ( );
FILL FILL_22_DFFPOSX1_15 ( );
FILL FILL_23_DFFPOSX1_15 ( );
FILL FILL_24_DFFPOSX1_15 ( );
FILL FILL_25_DFFPOSX1_15 ( );
FILL FILL_26_DFFPOSX1_15 ( );
FILL FILL_27_DFFPOSX1_15 ( );
FILL FILL_0_BUFX2_35 ( );
FILL FILL_1_BUFX2_35 ( );
FILL FILL_2_BUFX2_35 ( );
FILL FILL_3_BUFX2_35 ( );
FILL FILL_4_BUFX2_35 ( );
FILL FILL_5_BUFX2_35 ( );
FILL FILL_6_BUFX2_35 ( );
FILL FILL_0_BUFX2_40 ( );
FILL FILL_1_BUFX2_40 ( );
FILL FILL_2_BUFX2_40 ( );
FILL FILL_3_BUFX2_40 ( );
FILL FILL_4_BUFX2_40 ( );
FILL FILL_5_BUFX2_40 ( );
FILL FILL_6_BUFX2_40 ( );
FILL FILL_0_NAND2X1_175 ( );
FILL FILL_1_NAND2X1_175 ( );
FILL FILL_2_NAND2X1_175 ( );
FILL FILL_3_NAND2X1_175 ( );
FILL FILL_4_NAND2X1_175 ( );
FILL FILL_5_NAND2X1_175 ( );
FILL FILL_6_NAND2X1_175 ( );
FILL FILL_0_OAI21X1_12 ( );
FILL FILL_1_OAI21X1_12 ( );
FILL FILL_2_OAI21X1_12 ( );
FILL FILL_3_OAI21X1_12 ( );
FILL FILL_4_OAI21X1_12 ( );
FILL FILL_5_OAI21X1_12 ( );
FILL FILL_6_OAI21X1_12 ( );
FILL FILL_7_OAI21X1_12 ( );
FILL FILL_8_OAI21X1_12 ( );
FILL FILL_9_OAI21X1_12 ( );
FILL FILL_0_INVX1_14 ( );
FILL FILL_1_INVX1_14 ( );
FILL FILL_2_INVX1_14 ( );
FILL FILL_3_INVX1_14 ( );
FILL FILL_0_NAND2X1_173 ( );
FILL FILL_1_NAND2X1_173 ( );
FILL FILL_2_NAND2X1_173 ( );
FILL FILL_3_NAND2X1_173 ( );
FILL FILL_4_NAND2X1_173 ( );
FILL FILL_5_NAND2X1_173 ( );
FILL FILL_6_NAND2X1_173 ( );
FILL FILL_0_AND2X2_11 ( );
FILL FILL_1_AND2X2_11 ( );
FILL FILL_2_AND2X2_11 ( );
FILL FILL_3_AND2X2_11 ( );
FILL FILL_4_AND2X2_11 ( );
FILL FILL_5_AND2X2_11 ( );
FILL FILL_6_AND2X2_11 ( );
FILL FILL_7_AND2X2_11 ( );
FILL FILL_8_AND2X2_11 ( );
FILL FILL_0_OAI21X1_221 ( );
FILL FILL_1_OAI21X1_221 ( );
FILL FILL_2_OAI21X1_221 ( );
FILL FILL_3_OAI21X1_221 ( );
FILL FILL_4_OAI21X1_221 ( );
FILL FILL_5_OAI21X1_221 ( );
FILL FILL_6_OAI21X1_221 ( );
FILL FILL_7_OAI21X1_221 ( );
FILL FILL_8_OAI21X1_221 ( );
FILL FILL_9_OAI21X1_221 ( );
FILL FILL_0_INVX1_249 ( );
FILL FILL_1_INVX1_249 ( );
FILL FILL_2_INVX1_249 ( );
FILL FILL_3_INVX1_249 ( );
FILL FILL_0_NAND3X1_64 ( );
FILL FILL_1_NAND3X1_64 ( );
FILL FILL_2_NAND3X1_64 ( );
FILL FILL_3_NAND3X1_64 ( );
FILL FILL_4_NAND3X1_64 ( );
FILL FILL_5_NAND3X1_64 ( );
FILL FILL_6_NAND3X1_64 ( );
FILL FILL_7_NAND3X1_64 ( );
FILL FILL_8_NAND3X1_64 ( );
FILL FILL_9_NAND3X1_64 ( );
FILL FILL_0_NAND3X1_68 ( );
FILL FILL_1_NAND3X1_68 ( );
FILL FILL_2_NAND3X1_68 ( );
FILL FILL_3_NAND3X1_68 ( );
FILL FILL_4_NAND3X1_68 ( );
FILL FILL_5_NAND3X1_68 ( );
FILL FILL_6_NAND3X1_68 ( );
FILL FILL_7_NAND3X1_68 ( );
FILL FILL_8_NAND3X1_68 ( );
FILL FILL_0_NAND3X1_65 ( );
FILL FILL_1_NAND3X1_65 ( );
FILL FILL_2_NAND3X1_65 ( );
FILL FILL_3_NAND3X1_65 ( );
FILL FILL_4_NAND3X1_65 ( );
FILL FILL_5_NAND3X1_65 ( );
FILL FILL_6_NAND3X1_65 ( );
FILL FILL_7_NAND3X1_65 ( );
FILL FILL_8_NAND3X1_65 ( );
FILL FILL_0_INVX1_226 ( );
FILL FILL_1_INVX1_226 ( );
FILL FILL_2_INVX1_226 ( );
FILL FILL_3_INVX1_226 ( );
FILL FILL_4_INVX1_226 ( );
FILL FILL_0_OAI21X1_216 ( );
FILL FILL_1_OAI21X1_216 ( );
FILL FILL_2_OAI21X1_216 ( );
FILL FILL_3_OAI21X1_216 ( );
FILL FILL_4_OAI21X1_216 ( );
FILL FILL_5_OAI21X1_216 ( );
FILL FILL_6_OAI21X1_216 ( );
FILL FILL_7_OAI21X1_216 ( );
FILL FILL_8_OAI21X1_216 ( );
FILL FILL_0_INVX1_240 ( );
FILL FILL_1_INVX1_240 ( );
FILL FILL_2_INVX1_240 ( );
FILL FILL_3_INVX1_240 ( );
FILL FILL_0_OAI21X1_203 ( );
FILL FILL_1_OAI21X1_203 ( );
FILL FILL_2_OAI21X1_203 ( );
FILL FILL_3_OAI21X1_203 ( );
FILL FILL_4_OAI21X1_203 ( );
FILL FILL_5_OAI21X1_203 ( );
FILL FILL_6_OAI21X1_203 ( );
FILL FILL_7_OAI21X1_203 ( );
FILL FILL_8_OAI21X1_203 ( );
FILL FILL_9_OAI21X1_203 ( );
FILL FILL_0_INVX1_192 ( );
FILL FILL_1_INVX1_192 ( );
FILL FILL_2_INVX1_192 ( );
FILL FILL_3_INVX1_192 ( );
FILL FILL_4_INVX1_192 ( );
FILL FILL_0_NAND2X1_201 ( );
FILL FILL_1_NAND2X1_201 ( );
FILL FILL_2_NAND2X1_201 ( );
FILL FILL_3_NAND2X1_201 ( );
FILL FILL_4_NAND2X1_201 ( );
FILL FILL_5_NAND2X1_201 ( );
FILL FILL_6_NAND2X1_201 ( );
FILL FILL_0_OAI21X1_202 ( );
FILL FILL_1_OAI21X1_202 ( );
FILL FILL_2_OAI21X1_202 ( );
FILL FILL_3_OAI21X1_202 ( );
FILL FILL_4_OAI21X1_202 ( );
FILL FILL_5_OAI21X1_202 ( );
FILL FILL_6_OAI21X1_202 ( );
FILL FILL_7_OAI21X1_202 ( );
FILL FILL_8_OAI21X1_202 ( );
FILL FILL_0_NAND2X1_220 ( );
FILL FILL_1_NAND2X1_220 ( );
FILL FILL_2_NAND2X1_220 ( );
FILL FILL_3_NAND2X1_220 ( );
FILL FILL_4_NAND2X1_220 ( );
FILL FILL_5_NAND2X1_220 ( );
FILL FILL_6_NAND2X1_220 ( );
FILL FILL_0_XNOR2X1_1 ( );
FILL FILL_1_XNOR2X1_1 ( );
FILL FILL_2_XNOR2X1_1 ( );
FILL FILL_3_XNOR2X1_1 ( );
FILL FILL_4_XNOR2X1_1 ( );
FILL FILL_5_XNOR2X1_1 ( );
FILL FILL_6_XNOR2X1_1 ( );
FILL FILL_7_XNOR2X1_1 ( );
FILL FILL_8_XNOR2X1_1 ( );
FILL FILL_9_XNOR2X1_1 ( );
FILL FILL_10_XNOR2X1_1 ( );
FILL FILL_11_XNOR2X1_1 ( );
FILL FILL_12_XNOR2X1_1 ( );
FILL FILL_13_XNOR2X1_1 ( );
FILL FILL_14_XNOR2X1_1 ( );
FILL FILL_15_XNOR2X1_1 ( );
FILL FILL_0_NAND3X1_71 ( );
FILL FILL_1_NAND3X1_71 ( );
FILL FILL_2_NAND3X1_71 ( );
FILL FILL_3_NAND3X1_71 ( );
FILL FILL_4_NAND3X1_71 ( );
FILL FILL_5_NAND3X1_71 ( );
FILL FILL_6_NAND3X1_71 ( );
FILL FILL_7_NAND3X1_71 ( );
FILL FILL_8_NAND3X1_71 ( );
FILL FILL_0_INVX1_245 ( );
FILL FILL_1_INVX1_245 ( );
FILL FILL_2_INVX1_245 ( );
FILL FILL_3_INVX1_245 ( );
FILL FILL_4_INVX1_245 ( );
FILL FILL_0_NAND3X1_70 ( );
FILL FILL_1_NAND3X1_70 ( );
FILL FILL_2_NAND3X1_70 ( );
FILL FILL_3_NAND3X1_70 ( );
FILL FILL_4_NAND3X1_70 ( );
FILL FILL_5_NAND3X1_70 ( );
FILL FILL_6_NAND3X1_70 ( );
FILL FILL_7_NAND3X1_70 ( );
FILL FILL_8_NAND3X1_70 ( );
FILL FILL_0_NAND3X1_74 ( );
FILL FILL_1_NAND3X1_74 ( );
FILL FILL_2_NAND3X1_74 ( );
FILL FILL_3_NAND3X1_74 ( );
FILL FILL_4_NAND3X1_74 ( );
FILL FILL_5_NAND3X1_74 ( );
FILL FILL_6_NAND3X1_74 ( );
FILL FILL_7_NAND3X1_74 ( );
FILL FILL_8_NAND3X1_74 ( );
FILL FILL_0_NAND3X1_98 ( );
FILL FILL_1_NAND3X1_98 ( );
FILL FILL_2_NAND3X1_98 ( );
FILL FILL_3_NAND3X1_98 ( );
FILL FILL_4_NAND3X1_98 ( );
FILL FILL_5_NAND3X1_98 ( );
FILL FILL_6_NAND3X1_98 ( );
FILL FILL_7_NAND3X1_98 ( );
FILL FILL_8_NAND3X1_98 ( );
FILL FILL_0_AOI21X1_33 ( );
FILL FILL_1_AOI21X1_33 ( );
FILL FILL_2_AOI21X1_33 ( );
FILL FILL_3_AOI21X1_33 ( );
FILL FILL_4_AOI21X1_33 ( );
FILL FILL_5_AOI21X1_33 ( );
FILL FILL_6_AOI21X1_33 ( );
FILL FILL_7_AOI21X1_33 ( );
FILL FILL_8_AOI21X1_33 ( );
FILL FILL_9_AOI21X1_33 ( );
FILL FILL_0_DFFSR_97 ( );
FILL FILL_1_DFFSR_97 ( );
FILL FILL_2_DFFSR_97 ( );
FILL FILL_3_DFFSR_97 ( );
FILL FILL_4_DFFSR_97 ( );
FILL FILL_5_DFFSR_97 ( );
FILL FILL_6_DFFSR_97 ( );
FILL FILL_7_DFFSR_97 ( );
FILL FILL_8_DFFSR_97 ( );
FILL FILL_9_DFFSR_97 ( );
FILL FILL_10_DFFSR_97 ( );
FILL FILL_11_DFFSR_97 ( );
FILL FILL_12_DFFSR_97 ( );
FILL FILL_13_DFFSR_97 ( );
FILL FILL_14_DFFSR_97 ( );
FILL FILL_15_DFFSR_97 ( );
FILL FILL_16_DFFSR_97 ( );
FILL FILL_17_DFFSR_97 ( );
FILL FILL_18_DFFSR_97 ( );
FILL FILL_19_DFFSR_97 ( );
FILL FILL_20_DFFSR_97 ( );
FILL FILL_21_DFFSR_97 ( );
FILL FILL_22_DFFSR_97 ( );
FILL FILL_23_DFFSR_97 ( );
FILL FILL_24_DFFSR_97 ( );
FILL FILL_25_DFFSR_97 ( );
FILL FILL_26_DFFSR_97 ( );
FILL FILL_27_DFFSR_97 ( );
FILL FILL_28_DFFSR_97 ( );
FILL FILL_29_DFFSR_97 ( );
FILL FILL_30_DFFSR_97 ( );
FILL FILL_31_DFFSR_97 ( );
FILL FILL_32_DFFSR_97 ( );
FILL FILL_33_DFFSR_97 ( );
FILL FILL_34_DFFSR_97 ( );
FILL FILL_35_DFFSR_97 ( );
FILL FILL_36_DFFSR_97 ( );
FILL FILL_37_DFFSR_97 ( );
FILL FILL_38_DFFSR_97 ( );
FILL FILL_39_DFFSR_97 ( );
FILL FILL_40_DFFSR_97 ( );
FILL FILL_41_DFFSR_97 ( );
FILL FILL_42_DFFSR_97 ( );
FILL FILL_43_DFFSR_97 ( );
FILL FILL_44_DFFSR_97 ( );
FILL FILL_45_DFFSR_97 ( );
FILL FILL_46_DFFSR_97 ( );
FILL FILL_47_DFFSR_97 ( );
FILL FILL_48_DFFSR_97 ( );
FILL FILL_49_DFFSR_97 ( );
FILL FILL_50_DFFSR_97 ( );
FILL FILL_51_DFFSR_97 ( );
FILL FILL_0_OAI21X1_117 ( );
FILL FILL_1_OAI21X1_117 ( );
FILL FILL_2_OAI21X1_117 ( );
FILL FILL_3_OAI21X1_117 ( );
FILL FILL_4_OAI21X1_117 ( );
FILL FILL_5_OAI21X1_117 ( );
FILL FILL_6_OAI21X1_117 ( );
FILL FILL_7_OAI21X1_117 ( );
FILL FILL_8_OAI21X1_117 ( );
FILL FILL_0_INVX1_132 ( );
FILL FILL_1_INVX1_132 ( );
FILL FILL_2_INVX1_132 ( );
FILL FILL_3_INVX1_132 ( );
FILL FILL_4_INVX1_132 ( );
FILL FILL_0_INVX1_354 ( );
FILL FILL_1_INVX1_354 ( );
FILL FILL_2_INVX1_354 ( );
FILL FILL_3_INVX1_354 ( );
FILL FILL_4_INVX1_354 ( );
FILL FILL_0_INVX1_109 ( );
FILL FILL_1_INVX1_109 ( );
FILL FILL_2_INVX1_109 ( );
FILL FILL_3_INVX1_109 ( );
FILL FILL_4_INVX1_109 ( );
FILL FILL_0_DFFSR_99 ( );
FILL FILL_1_DFFSR_99 ( );
FILL FILL_2_DFFSR_99 ( );
FILL FILL_3_DFFSR_99 ( );
FILL FILL_4_DFFSR_99 ( );
FILL FILL_5_DFFSR_99 ( );
FILL FILL_6_DFFSR_99 ( );
FILL FILL_7_DFFSR_99 ( );
FILL FILL_8_DFFSR_99 ( );
FILL FILL_9_DFFSR_99 ( );
FILL FILL_10_DFFSR_99 ( );
FILL FILL_11_DFFSR_99 ( );
FILL FILL_12_DFFSR_99 ( );
FILL FILL_13_DFFSR_99 ( );
FILL FILL_14_DFFSR_99 ( );
FILL FILL_15_DFFSR_99 ( );
FILL FILL_16_DFFSR_99 ( );
FILL FILL_17_DFFSR_99 ( );
FILL FILL_18_DFFSR_99 ( );
FILL FILL_19_DFFSR_99 ( );
FILL FILL_20_DFFSR_99 ( );
FILL FILL_21_DFFSR_99 ( );
FILL FILL_22_DFFSR_99 ( );
FILL FILL_23_DFFSR_99 ( );
FILL FILL_24_DFFSR_99 ( );
FILL FILL_25_DFFSR_99 ( );
FILL FILL_26_DFFSR_99 ( );
FILL FILL_27_DFFSR_99 ( );
FILL FILL_28_DFFSR_99 ( );
FILL FILL_29_DFFSR_99 ( );
FILL FILL_30_DFFSR_99 ( );
FILL FILL_31_DFFSR_99 ( );
FILL FILL_32_DFFSR_99 ( );
FILL FILL_33_DFFSR_99 ( );
FILL FILL_34_DFFSR_99 ( );
FILL FILL_35_DFFSR_99 ( );
FILL FILL_36_DFFSR_99 ( );
FILL FILL_37_DFFSR_99 ( );
FILL FILL_38_DFFSR_99 ( );
FILL FILL_39_DFFSR_99 ( );
FILL FILL_40_DFFSR_99 ( );
FILL FILL_41_DFFSR_99 ( );
FILL FILL_42_DFFSR_99 ( );
FILL FILL_43_DFFSR_99 ( );
FILL FILL_44_DFFSR_99 ( );
FILL FILL_45_DFFSR_99 ( );
FILL FILL_46_DFFSR_99 ( );
FILL FILL_47_DFFSR_99 ( );
FILL FILL_48_DFFSR_99 ( );
FILL FILL_49_DFFSR_99 ( );
FILL FILL_50_DFFSR_99 ( );
FILL FILL_0_INVX1_82 ( );
FILL FILL_1_INVX1_82 ( );
FILL FILL_2_INVX1_82 ( );
FILL FILL_3_INVX1_82 ( );
FILL FILL_4_INVX1_82 ( );
FILL FILL_0_OAI21X1_157 ( );
FILL FILL_1_OAI21X1_157 ( );
FILL FILL_2_OAI21X1_157 ( );
FILL FILL_3_OAI21X1_157 ( );
FILL FILL_4_OAI21X1_157 ( );
FILL FILL_5_OAI21X1_157 ( );
FILL FILL_6_OAI21X1_157 ( );
FILL FILL_7_OAI21X1_157 ( );
FILL FILL_8_OAI21X1_157 ( );
FILL FILL_0_INVX1_188 ( );
FILL FILL_1_INVX1_188 ( );
FILL FILL_2_INVX1_188 ( );
FILL FILL_3_INVX1_188 ( );
FILL FILL_4_INVX1_188 ( );
FILL FILL_0_NAND2X1_157 ( );
FILL FILL_1_NAND2X1_157 ( );
FILL FILL_2_NAND2X1_157 ( );
FILL FILL_3_NAND2X1_157 ( );
FILL FILL_4_NAND2X1_157 ( );
FILL FILL_5_NAND2X1_157 ( );
FILL FILL_6_NAND2X1_157 ( );
FILL FILL_0_NAND2X1_158 ( );
FILL FILL_1_NAND2X1_158 ( );
FILL FILL_2_NAND2X1_158 ( );
FILL FILL_3_NAND2X1_158 ( );
FILL FILL_4_NAND2X1_158 ( );
FILL FILL_5_NAND2X1_158 ( );
FILL FILL_6_NAND2X1_158 ( );
FILL FILL_0_INVX1_437 ( );
FILL FILL_1_INVX1_437 ( );
FILL FILL_2_INVX1_437 ( );
FILL FILL_3_INVX1_437 ( );
FILL FILL_4_INVX1_437 ( );
FILL FILL_0_AND2X2_14 ( );
FILL FILL_1_AND2X2_14 ( );
FILL FILL_2_AND2X2_14 ( );
FILL FILL_3_AND2X2_14 ( );
FILL FILL_4_AND2X2_14 ( );
FILL FILL_5_AND2X2_14 ( );
FILL FILL_6_AND2X2_14 ( );
FILL FILL_7_AND2X2_14 ( );
FILL FILL_8_AND2X2_14 ( );
FILL FILL_9_AND2X2_14 ( );
FILL FILL_0_OAI21X1_241 ( );
FILL FILL_1_OAI21X1_241 ( );
FILL FILL_2_OAI21X1_241 ( );
FILL FILL_3_OAI21X1_241 ( );
FILL FILL_4_OAI21X1_241 ( );
FILL FILL_5_OAI21X1_241 ( );
FILL FILL_6_OAI21X1_241 ( );
FILL FILL_7_OAI21X1_241 ( );
FILL FILL_8_OAI21X1_241 ( );
FILL FILL_9_OAI21X1_241 ( );
FILL FILL_0_NAND2X1_251 ( );
FILL FILL_1_NAND2X1_251 ( );
FILL FILL_2_NAND2X1_251 ( );
FILL FILL_3_NAND2X1_251 ( );
FILL FILL_4_NAND2X1_251 ( );
FILL FILL_5_NAND2X1_251 ( );
FILL FILL_6_NAND2X1_251 ( );
FILL FILL_0_INVX1_400 ( );
FILL FILL_1_INVX1_400 ( );
FILL FILL_2_INVX1_400 ( );
FILL FILL_3_INVX1_400 ( );
FILL FILL_0_OAI21X1_242 ( );
FILL FILL_1_OAI21X1_242 ( );
FILL FILL_2_OAI21X1_242 ( );
FILL FILL_3_OAI21X1_242 ( );
FILL FILL_4_OAI21X1_242 ( );
FILL FILL_5_OAI21X1_242 ( );
FILL FILL_6_OAI21X1_242 ( );
FILL FILL_7_OAI21X1_242 ( );
FILL FILL_8_OAI21X1_242 ( );
FILL FILL_9_OAI21X1_242 ( );
FILL FILL_0_BUFX2_43 ( );
FILL FILL_1_BUFX2_43 ( );
FILL FILL_2_BUFX2_43 ( );
FILL FILL_3_BUFX2_43 ( );
FILL FILL_4_BUFX2_43 ( );
FILL FILL_5_BUFX2_43 ( );
FILL FILL_6_BUFX2_43 ( );
FILL FILL_0_INVX1_35 ( );
FILL FILL_1_INVX1_35 ( );
FILL FILL_2_INVX1_35 ( );
FILL FILL_3_INVX1_35 ( );
FILL FILL_4_INVX1_35 ( );
FILL FILL_0_OAI21X1_31 ( );
FILL FILL_1_OAI21X1_31 ( );
FILL FILL_2_OAI21X1_31 ( );
FILL FILL_3_OAI21X1_31 ( );
FILL FILL_4_OAI21X1_31 ( );
FILL FILL_5_OAI21X1_31 ( );
FILL FILL_6_OAI21X1_31 ( );
FILL FILL_7_OAI21X1_31 ( );
FILL FILL_8_OAI21X1_31 ( );
FILL FILL_0_DFFSR_31 ( );
FILL FILL_1_DFFSR_31 ( );
FILL FILL_2_DFFSR_31 ( );
FILL FILL_3_DFFSR_31 ( );
FILL FILL_4_DFFSR_31 ( );
FILL FILL_5_DFFSR_31 ( );
FILL FILL_6_DFFSR_31 ( );
FILL FILL_7_DFFSR_31 ( );
FILL FILL_8_DFFSR_31 ( );
FILL FILL_9_DFFSR_31 ( );
FILL FILL_10_DFFSR_31 ( );
FILL FILL_11_DFFSR_31 ( );
FILL FILL_12_DFFSR_31 ( );
FILL FILL_13_DFFSR_31 ( );
FILL FILL_14_DFFSR_31 ( );
FILL FILL_15_DFFSR_31 ( );
FILL FILL_16_DFFSR_31 ( );
FILL FILL_17_DFFSR_31 ( );
FILL FILL_18_DFFSR_31 ( );
FILL FILL_19_DFFSR_31 ( );
FILL FILL_20_DFFSR_31 ( );
FILL FILL_21_DFFSR_31 ( );
FILL FILL_22_DFFSR_31 ( );
FILL FILL_23_DFFSR_31 ( );
FILL FILL_24_DFFSR_31 ( );
FILL FILL_25_DFFSR_31 ( );
FILL FILL_26_DFFSR_31 ( );
FILL FILL_27_DFFSR_31 ( );
FILL FILL_28_DFFSR_31 ( );
FILL FILL_29_DFFSR_31 ( );
FILL FILL_30_DFFSR_31 ( );
FILL FILL_31_DFFSR_31 ( );
FILL FILL_32_DFFSR_31 ( );
FILL FILL_33_DFFSR_31 ( );
FILL FILL_34_DFFSR_31 ( );
FILL FILL_35_DFFSR_31 ( );
FILL FILL_36_DFFSR_31 ( );
FILL FILL_37_DFFSR_31 ( );
FILL FILL_38_DFFSR_31 ( );
FILL FILL_39_DFFSR_31 ( );
FILL FILL_40_DFFSR_31 ( );
FILL FILL_41_DFFSR_31 ( );
FILL FILL_42_DFFSR_31 ( );
FILL FILL_43_DFFSR_31 ( );
FILL FILL_44_DFFSR_31 ( );
FILL FILL_45_DFFSR_31 ( );
FILL FILL_46_DFFSR_31 ( );
FILL FILL_47_DFFSR_31 ( );
FILL FILL_48_DFFSR_31 ( );
FILL FILL_49_DFFSR_31 ( );
FILL FILL_50_DFFSR_31 ( );
FILL FILL_0_OAI21X1_219 ( );
FILL FILL_1_OAI21X1_219 ( );
FILL FILL_2_OAI21X1_219 ( );
FILL FILL_3_OAI21X1_219 ( );
FILL FILL_4_OAI21X1_219 ( );
FILL FILL_5_OAI21X1_219 ( );
FILL FILL_6_OAI21X1_219 ( );
FILL FILL_7_OAI21X1_219 ( );
FILL FILL_8_OAI21X1_219 ( );
FILL FILL_0_NAND2X1_214 ( );
FILL FILL_1_NAND2X1_214 ( );
FILL FILL_2_NAND2X1_214 ( );
FILL FILL_3_NAND2X1_214 ( );
FILL FILL_4_NAND2X1_214 ( );
FILL FILL_5_NAND2X1_214 ( );
FILL FILL_6_NAND2X1_214 ( );
FILL FILL_0_OAI21X1_232 ( );
FILL FILL_1_OAI21X1_232 ( );
FILL FILL_2_OAI21X1_232 ( );
FILL FILL_3_OAI21X1_232 ( );
FILL FILL_4_OAI21X1_232 ( );
FILL FILL_5_OAI21X1_232 ( );
FILL FILL_6_OAI21X1_232 ( );
FILL FILL_7_OAI21X1_232 ( );
FILL FILL_8_OAI21X1_232 ( );
FILL FILL_0_NAND2X1_202 ( );
FILL FILL_1_NAND2X1_202 ( );
FILL FILL_2_NAND2X1_202 ( );
FILL FILL_3_NAND2X1_202 ( );
FILL FILL_4_NAND2X1_202 ( );
FILL FILL_5_NAND2X1_202 ( );
FILL FILL_6_NAND2X1_202 ( );
FILL FILL_0_NAND2X1_213 ( );
FILL FILL_1_NAND2X1_213 ( );
FILL FILL_2_NAND2X1_213 ( );
FILL FILL_3_NAND2X1_213 ( );
FILL FILL_4_NAND2X1_213 ( );
FILL FILL_5_NAND2X1_213 ( );
FILL FILL_6_NAND2X1_213 ( );
FILL FILL_0_NAND2X1_210 ( );
FILL FILL_1_NAND2X1_210 ( );
FILL FILL_2_NAND2X1_210 ( );
FILL FILL_3_NAND2X1_210 ( );
FILL FILL_4_NAND2X1_210 ( );
FILL FILL_5_NAND2X1_210 ( );
FILL FILL_6_NAND2X1_210 ( );
FILL FILL_0_NAND2X1_190 ( );
FILL FILL_1_NAND2X1_190 ( );
FILL FILL_2_NAND2X1_190 ( );
FILL FILL_3_NAND2X1_190 ( );
FILL FILL_4_NAND2X1_190 ( );
FILL FILL_5_NAND2X1_190 ( );
FILL FILL_6_NAND2X1_190 ( );
FILL FILL_0_OAI21X1_214 ( );
FILL FILL_1_OAI21X1_214 ( );
FILL FILL_2_OAI21X1_214 ( );
FILL FILL_3_OAI21X1_214 ( );
FILL FILL_4_OAI21X1_214 ( );
FILL FILL_5_OAI21X1_214 ( );
FILL FILL_6_OAI21X1_214 ( );
FILL FILL_7_OAI21X1_214 ( );
FILL FILL_8_OAI21X1_214 ( );
FILL FILL_9_OAI21X1_214 ( );
FILL FILL_0_OAI21X1_201 ( );
FILL FILL_1_OAI21X1_201 ( );
FILL FILL_2_OAI21X1_201 ( );
FILL FILL_3_OAI21X1_201 ( );
FILL FILL_4_OAI21X1_201 ( );
FILL FILL_5_OAI21X1_201 ( );
FILL FILL_6_OAI21X1_201 ( );
FILL FILL_7_OAI21X1_201 ( );
FILL FILL_8_OAI21X1_201 ( );
FILL FILL_9_OAI21X1_201 ( );
FILL FILL_0_NAND3X1_36 ( );
FILL FILL_1_NAND3X1_36 ( );
FILL FILL_2_NAND3X1_36 ( );
FILL FILL_3_NAND3X1_36 ( );
FILL FILL_4_NAND3X1_36 ( );
FILL FILL_5_NAND3X1_36 ( );
FILL FILL_6_NAND3X1_36 ( );
FILL FILL_7_NAND3X1_36 ( );
FILL FILL_8_NAND3X1_36 ( );
FILL FILL_0_NAND3X1_46 ( );
FILL FILL_1_NAND3X1_46 ( );
FILL FILL_2_NAND3X1_46 ( );
FILL FILL_3_NAND3X1_46 ( );
FILL FILL_4_NAND3X1_46 ( );
FILL FILL_5_NAND3X1_46 ( );
FILL FILL_6_NAND3X1_46 ( );
FILL FILL_7_NAND3X1_46 ( );
FILL FILL_8_NAND3X1_46 ( );
FILL FILL_0_INVX1_239 ( );
FILL FILL_1_INVX1_239 ( );
FILL FILL_2_INVX1_239 ( );
FILL FILL_3_INVX1_239 ( );
FILL FILL_0_NAND3X1_35 ( );
FILL FILL_1_NAND3X1_35 ( );
FILL FILL_2_NAND3X1_35 ( );
FILL FILL_3_NAND3X1_35 ( );
FILL FILL_4_NAND3X1_35 ( );
FILL FILL_5_NAND3X1_35 ( );
FILL FILL_6_NAND3X1_35 ( );
FILL FILL_7_NAND3X1_35 ( );
FILL FILL_8_NAND3X1_35 ( );
FILL FILL_0_NAND3X1_45 ( );
FILL FILL_1_NAND3X1_45 ( );
FILL FILL_2_NAND3X1_45 ( );
FILL FILL_3_NAND3X1_45 ( );
FILL FILL_4_NAND3X1_45 ( );
FILL FILL_5_NAND3X1_45 ( );
FILL FILL_6_NAND3X1_45 ( );
FILL FILL_7_NAND3X1_45 ( );
FILL FILL_8_NAND3X1_45 ( );
FILL FILL_9_NAND3X1_45 ( );
FILL FILL_0_OAI21X1_165 ( );
FILL FILL_1_OAI21X1_165 ( );
FILL FILL_2_OAI21X1_165 ( );
FILL FILL_3_OAI21X1_165 ( );
FILL FILL_4_OAI21X1_165 ( );
FILL FILL_5_OAI21X1_165 ( );
FILL FILL_6_OAI21X1_165 ( );
FILL FILL_7_OAI21X1_165 ( );
FILL FILL_8_OAI21X1_165 ( );
FILL FILL_0_INVX1_223 ( );
FILL FILL_1_INVX1_223 ( );
FILL FILL_2_INVX1_223 ( );
FILL FILL_3_INVX1_223 ( );
FILL FILL_4_INVX1_223 ( );
FILL FILL_0_INVX1_199 ( );
FILL FILL_1_INVX1_199 ( );
FILL FILL_2_INVX1_199 ( );
FILL FILL_3_INVX1_199 ( );
FILL FILL_4_INVX1_199 ( );
FILL FILL_0_NAND3X1_75 ( );
FILL FILL_1_NAND3X1_75 ( );
FILL FILL_2_NAND3X1_75 ( );
FILL FILL_3_NAND3X1_75 ( );
FILL FILL_4_NAND3X1_75 ( );
FILL FILL_5_NAND3X1_75 ( );
FILL FILL_6_NAND3X1_75 ( );
FILL FILL_7_NAND3X1_75 ( );
FILL FILL_8_NAND3X1_75 ( );
FILL FILL_0_NAND3X1_94 ( );
FILL FILL_1_NAND3X1_94 ( );
FILL FILL_2_NAND3X1_94 ( );
FILL FILL_3_NAND3X1_94 ( );
FILL FILL_4_NAND3X1_94 ( );
FILL FILL_5_NAND3X1_94 ( );
FILL FILL_6_NAND3X1_94 ( );
FILL FILL_7_NAND3X1_94 ( );
FILL FILL_8_NAND3X1_94 ( );
FILL FILL_9_NAND3X1_94 ( );
FILL FILL_0_NAND3X1_97 ( );
FILL FILL_1_NAND3X1_97 ( );
FILL FILL_2_NAND3X1_97 ( );
FILL FILL_3_NAND3X1_97 ( );
FILL FILL_4_NAND3X1_97 ( );
FILL FILL_5_NAND3X1_97 ( );
FILL FILL_6_NAND3X1_97 ( );
FILL FILL_7_NAND3X1_97 ( );
FILL FILL_8_NAND3X1_97 ( );
FILL FILL_9_NAND3X1_97 ( );
FILL FILL_0_INVX1_253 ( );
FILL FILL_1_INVX1_253 ( );
FILL FILL_2_INVX1_253 ( );
FILL FILL_3_INVX1_253 ( );
FILL FILL_0_DFFSR_127 ( );
FILL FILL_1_DFFSR_127 ( );
FILL FILL_2_DFFSR_127 ( );
FILL FILL_3_DFFSR_127 ( );
FILL FILL_4_DFFSR_127 ( );
FILL FILL_5_DFFSR_127 ( );
FILL FILL_6_DFFSR_127 ( );
FILL FILL_7_DFFSR_127 ( );
FILL FILL_8_DFFSR_127 ( );
FILL FILL_9_DFFSR_127 ( );
FILL FILL_10_DFFSR_127 ( );
FILL FILL_11_DFFSR_127 ( );
FILL FILL_12_DFFSR_127 ( );
FILL FILL_13_DFFSR_127 ( );
FILL FILL_14_DFFSR_127 ( );
FILL FILL_15_DFFSR_127 ( );
FILL FILL_16_DFFSR_127 ( );
FILL FILL_17_DFFSR_127 ( );
FILL FILL_18_DFFSR_127 ( );
FILL FILL_19_DFFSR_127 ( );
FILL FILL_20_DFFSR_127 ( );
FILL FILL_21_DFFSR_127 ( );
FILL FILL_22_DFFSR_127 ( );
FILL FILL_23_DFFSR_127 ( );
FILL FILL_24_DFFSR_127 ( );
FILL FILL_25_DFFSR_127 ( );
FILL FILL_26_DFFSR_127 ( );
FILL FILL_27_DFFSR_127 ( );
FILL FILL_28_DFFSR_127 ( );
FILL FILL_29_DFFSR_127 ( );
FILL FILL_30_DFFSR_127 ( );
FILL FILL_31_DFFSR_127 ( );
FILL FILL_32_DFFSR_127 ( );
FILL FILL_33_DFFSR_127 ( );
FILL FILL_34_DFFSR_127 ( );
FILL FILL_35_DFFSR_127 ( );
FILL FILL_36_DFFSR_127 ( );
FILL FILL_37_DFFSR_127 ( );
FILL FILL_38_DFFSR_127 ( );
FILL FILL_39_DFFSR_127 ( );
FILL FILL_40_DFFSR_127 ( );
FILL FILL_41_DFFSR_127 ( );
FILL FILL_42_DFFSR_127 ( );
FILL FILL_43_DFFSR_127 ( );
FILL FILL_44_DFFSR_127 ( );
FILL FILL_45_DFFSR_127 ( );
FILL FILL_46_DFFSR_127 ( );
FILL FILL_47_DFFSR_127 ( );
FILL FILL_48_DFFSR_127 ( );
FILL FILL_49_DFFSR_127 ( );
FILL FILL_50_DFFSR_127 ( );
FILL FILL_0_CLKBUF1_7 ( );
FILL FILL_1_CLKBUF1_7 ( );
FILL FILL_2_CLKBUF1_7 ( );
FILL FILL_3_CLKBUF1_7 ( );
FILL FILL_4_CLKBUF1_7 ( );
FILL FILL_5_CLKBUF1_7 ( );
FILL FILL_6_CLKBUF1_7 ( );
FILL FILL_7_CLKBUF1_7 ( );
FILL FILL_8_CLKBUF1_7 ( );
FILL FILL_9_CLKBUF1_7 ( );
FILL FILL_10_CLKBUF1_7 ( );
FILL FILL_11_CLKBUF1_7 ( );
FILL FILL_12_CLKBUF1_7 ( );
FILL FILL_13_CLKBUF1_7 ( );
FILL FILL_14_CLKBUF1_7 ( );
FILL FILL_15_CLKBUF1_7 ( );
FILL FILL_16_CLKBUF1_7 ( );
FILL FILL_17_CLKBUF1_7 ( );
FILL FILL_18_CLKBUF1_7 ( );
FILL FILL_19_CLKBUF1_7 ( );
FILL FILL_0_INVX1_145 ( );
FILL FILL_1_INVX1_145 ( );
FILL FILL_2_INVX1_145 ( );
FILL FILL_3_INVX1_145 ( );
FILL FILL_4_INVX1_145 ( );
FILL FILL_0_OAI21X1_91 ( );
FILL FILL_1_OAI21X1_91 ( );
FILL FILL_2_OAI21X1_91 ( );
FILL FILL_3_OAI21X1_91 ( );
FILL FILL_4_OAI21X1_91 ( );
FILL FILL_5_OAI21X1_91 ( );
FILL FILL_6_OAI21X1_91 ( );
FILL FILL_7_OAI21X1_91 ( );
FILL FILL_8_OAI21X1_91 ( );
FILL FILL_0_INVX1_103 ( );
FILL FILL_1_INVX1_103 ( );
FILL FILL_2_INVX1_103 ( );
FILL FILL_3_INVX1_103 ( );
FILL FILL_4_INVX1_103 ( );
FILL FILL_0_NAND2X1_99 ( );
FILL FILL_1_NAND2X1_99 ( );
FILL FILL_2_NAND2X1_99 ( );
FILL FILL_3_NAND2X1_99 ( );
FILL FILL_4_NAND2X1_99 ( );
FILL FILL_5_NAND2X1_99 ( );
FILL FILL_6_NAND2X1_99 ( );
FILL FILL_0_OAI21X1_99 ( );
FILL FILL_1_OAI21X1_99 ( );
FILL FILL_2_OAI21X1_99 ( );
FILL FILL_3_OAI21X1_99 ( );
FILL FILL_4_OAI21X1_99 ( );
FILL FILL_5_OAI21X1_99 ( );
FILL FILL_6_OAI21X1_99 ( );
FILL FILL_7_OAI21X1_99 ( );
FILL FILL_8_OAI21X1_99 ( );
FILL FILL_9_OAI21X1_99 ( );
FILL FILL_0_INVX1_112 ( );
FILL FILL_1_INVX1_112 ( );
FILL FILL_2_INVX1_112 ( );
FILL FILL_3_INVX1_112 ( );
FILL FILL_0_INVX1_136 ( );
FILL FILL_1_INVX1_136 ( );
FILL FILL_2_INVX1_136 ( );
FILL FILL_3_INVX1_136 ( );
FILL FILL_4_INVX1_136 ( );
FILL FILL_0_DFFSR_135 ( );
FILL FILL_1_DFFSR_135 ( );
FILL FILL_2_DFFSR_135 ( );
FILL FILL_3_DFFSR_135 ( );
FILL FILL_4_DFFSR_135 ( );
FILL FILL_5_DFFSR_135 ( );
FILL FILL_6_DFFSR_135 ( );
FILL FILL_7_DFFSR_135 ( );
FILL FILL_8_DFFSR_135 ( );
FILL FILL_9_DFFSR_135 ( );
FILL FILL_10_DFFSR_135 ( );
FILL FILL_11_DFFSR_135 ( );
FILL FILL_12_DFFSR_135 ( );
FILL FILL_13_DFFSR_135 ( );
FILL FILL_14_DFFSR_135 ( );
FILL FILL_15_DFFSR_135 ( );
FILL FILL_16_DFFSR_135 ( );
FILL FILL_17_DFFSR_135 ( );
FILL FILL_18_DFFSR_135 ( );
FILL FILL_19_DFFSR_135 ( );
FILL FILL_20_DFFSR_135 ( );
FILL FILL_21_DFFSR_135 ( );
FILL FILL_22_DFFSR_135 ( );
FILL FILL_23_DFFSR_135 ( );
FILL FILL_24_DFFSR_135 ( );
FILL FILL_25_DFFSR_135 ( );
FILL FILL_26_DFFSR_135 ( );
FILL FILL_27_DFFSR_135 ( );
FILL FILL_28_DFFSR_135 ( );
FILL FILL_29_DFFSR_135 ( );
FILL FILL_30_DFFSR_135 ( );
FILL FILL_31_DFFSR_135 ( );
FILL FILL_32_DFFSR_135 ( );
FILL FILL_33_DFFSR_135 ( );
FILL FILL_34_DFFSR_135 ( );
FILL FILL_35_DFFSR_135 ( );
FILL FILL_36_DFFSR_135 ( );
FILL FILL_37_DFFSR_135 ( );
FILL FILL_38_DFFSR_135 ( );
FILL FILL_39_DFFSR_135 ( );
FILL FILL_40_DFFSR_135 ( );
FILL FILL_41_DFFSR_135 ( );
FILL FILL_42_DFFSR_135 ( );
FILL FILL_43_DFFSR_135 ( );
FILL FILL_44_DFFSR_135 ( );
FILL FILL_45_DFFSR_135 ( );
FILL FILL_46_DFFSR_135 ( );
FILL FILL_47_DFFSR_135 ( );
FILL FILL_48_DFFSR_135 ( );
FILL FILL_49_DFFSR_135 ( );
FILL FILL_50_DFFSR_135 ( );
FILL FILL_51_DFFSR_135 ( );
FILL FILL_0_OAI21X1_265 ( );
FILL FILL_1_OAI21X1_265 ( );
FILL FILL_2_OAI21X1_265 ( );
FILL FILL_3_OAI21X1_265 ( );
FILL FILL_4_OAI21X1_265 ( );
FILL FILL_5_OAI21X1_265 ( );
FILL FILL_6_OAI21X1_265 ( );
FILL FILL_7_OAI21X1_265 ( );
FILL FILL_8_OAI21X1_265 ( );
FILL FILL_0_DFFPOSX1_30 ( );
FILL FILL_1_DFFPOSX1_30 ( );
FILL FILL_2_DFFPOSX1_30 ( );
FILL FILL_3_DFFPOSX1_30 ( );
FILL FILL_4_DFFPOSX1_30 ( );
FILL FILL_5_DFFPOSX1_30 ( );
FILL FILL_6_DFFPOSX1_30 ( );
FILL FILL_7_DFFPOSX1_30 ( );
FILL FILL_8_DFFPOSX1_30 ( );
FILL FILL_9_DFFPOSX1_30 ( );
FILL FILL_10_DFFPOSX1_30 ( );
FILL FILL_11_DFFPOSX1_30 ( );
FILL FILL_12_DFFPOSX1_30 ( );
FILL FILL_13_DFFPOSX1_30 ( );
FILL FILL_14_DFFPOSX1_30 ( );
FILL FILL_15_DFFPOSX1_30 ( );
FILL FILL_16_DFFPOSX1_30 ( );
FILL FILL_17_DFFPOSX1_30 ( );
FILL FILL_18_DFFPOSX1_30 ( );
FILL FILL_19_DFFPOSX1_30 ( );
FILL FILL_20_DFFPOSX1_30 ( );
FILL FILL_21_DFFPOSX1_30 ( );
FILL FILL_22_DFFPOSX1_30 ( );
FILL FILL_23_DFFPOSX1_30 ( );
FILL FILL_24_DFFPOSX1_30 ( );
FILL FILL_25_DFFPOSX1_30 ( );
FILL FILL_26_DFFPOSX1_30 ( );
FILL FILL_27_DFFPOSX1_30 ( );
FILL FILL_0_OAI21X1_158 ( );
FILL FILL_1_OAI21X1_158 ( );
FILL FILL_2_OAI21X1_158 ( );
FILL FILL_3_OAI21X1_158 ( );
FILL FILL_4_OAI21X1_158 ( );
FILL FILL_5_OAI21X1_158 ( );
FILL FILL_6_OAI21X1_158 ( );
FILL FILL_7_OAI21X1_158 ( );
FILL FILL_8_OAI21X1_158 ( );
FILL FILL_0_INVX1_190 ( );
FILL FILL_1_INVX1_190 ( );
FILL FILL_2_INVX1_190 ( );
FILL FILL_3_INVX1_190 ( );
FILL FILL_4_INVX1_190 ( );
FILL FILL_0_NAND2X1_31 ( );
FILL FILL_1_NAND2X1_31 ( );
FILL FILL_2_NAND2X1_31 ( );
FILL FILL_3_NAND2X1_31 ( );
FILL FILL_4_NAND2X1_31 ( );
FILL FILL_5_NAND2X1_31 ( );
FILL FILL_6_NAND2X1_31 ( );
FILL FILL_0_NAND2X1_159 ( );
FILL FILL_1_NAND2X1_159 ( );
FILL FILL_2_NAND2X1_159 ( );
FILL FILL_3_NAND2X1_159 ( );
FILL FILL_4_NAND2X1_159 ( );
FILL FILL_5_NAND2X1_159 ( );
FILL FILL_6_NAND2X1_159 ( );
FILL FILL_0_BUFX2_39 ( );
FILL FILL_1_BUFX2_39 ( );
FILL FILL_2_BUFX2_39 ( );
FILL FILL_3_BUFX2_39 ( );
FILL FILL_4_BUFX2_39 ( );
FILL FILL_5_BUFX2_39 ( );
FILL FILL_6_BUFX2_39 ( );
FILL FILL_0_NAND2X1_174 ( );
FILL FILL_1_NAND2X1_174 ( );
FILL FILL_2_NAND2X1_174 ( );
FILL FILL_3_NAND2X1_174 ( );
FILL FILL_4_NAND2X1_174 ( );
FILL FILL_5_NAND2X1_174 ( );
FILL FILL_6_NAND2X1_174 ( );
FILL FILL_0_DFFSR_174 ( );
FILL FILL_1_DFFSR_174 ( );
FILL FILL_2_DFFSR_174 ( );
FILL FILL_3_DFFSR_174 ( );
FILL FILL_4_DFFSR_174 ( );
FILL FILL_5_DFFSR_174 ( );
FILL FILL_6_DFFSR_174 ( );
FILL FILL_7_DFFSR_174 ( );
FILL FILL_8_DFFSR_174 ( );
FILL FILL_9_DFFSR_174 ( );
FILL FILL_10_DFFSR_174 ( );
FILL FILL_11_DFFSR_174 ( );
FILL FILL_12_DFFSR_174 ( );
FILL FILL_13_DFFSR_174 ( );
FILL FILL_14_DFFSR_174 ( );
FILL FILL_15_DFFSR_174 ( );
FILL FILL_16_DFFSR_174 ( );
FILL FILL_17_DFFSR_174 ( );
FILL FILL_18_DFFSR_174 ( );
FILL FILL_19_DFFSR_174 ( );
FILL FILL_20_DFFSR_174 ( );
FILL FILL_21_DFFSR_174 ( );
FILL FILL_22_DFFSR_174 ( );
FILL FILL_23_DFFSR_174 ( );
FILL FILL_24_DFFSR_174 ( );
FILL FILL_25_DFFSR_174 ( );
FILL FILL_26_DFFSR_174 ( );
FILL FILL_27_DFFSR_174 ( );
FILL FILL_28_DFFSR_174 ( );
FILL FILL_29_DFFSR_174 ( );
FILL FILL_30_DFFSR_174 ( );
FILL FILL_31_DFFSR_174 ( );
FILL FILL_32_DFFSR_174 ( );
FILL FILL_33_DFFSR_174 ( );
FILL FILL_34_DFFSR_174 ( );
FILL FILL_35_DFFSR_174 ( );
FILL FILL_36_DFFSR_174 ( );
FILL FILL_37_DFFSR_174 ( );
FILL FILL_38_DFFSR_174 ( );
FILL FILL_39_DFFSR_174 ( );
FILL FILL_40_DFFSR_174 ( );
FILL FILL_41_DFFSR_174 ( );
FILL FILL_42_DFFSR_174 ( );
FILL FILL_43_DFFSR_174 ( );
FILL FILL_44_DFFSR_174 ( );
FILL FILL_45_DFFSR_174 ( );
FILL FILL_46_DFFSR_174 ( );
FILL FILL_47_DFFSR_174 ( );
FILL FILL_48_DFFSR_174 ( );
FILL FILL_49_DFFSR_174 ( );
FILL FILL_50_DFFSR_174 ( );
FILL FILL_51_DFFSR_174 ( );
FILL FILL_0_NOR2X1_9 ( );
FILL FILL_1_NOR2X1_9 ( );
FILL FILL_2_NOR2X1_9 ( );
FILL FILL_3_NOR2X1_9 ( );
FILL FILL_4_NOR2X1_9 ( );
FILL FILL_5_NOR2X1_9 ( );
FILL FILL_6_NOR2X1_9 ( );
FILL FILL_0_AND2X2_12 ( );
FILL FILL_1_AND2X2_12 ( );
FILL FILL_2_AND2X2_12 ( );
FILL FILL_3_AND2X2_12 ( );
FILL FILL_4_AND2X2_12 ( );
FILL FILL_5_AND2X2_12 ( );
FILL FILL_6_AND2X2_12 ( );
FILL FILL_7_AND2X2_12 ( );
FILL FILL_8_AND2X2_12 ( );
FILL FILL_9_AND2X2_12 ( );
FILL FILL_0_OAI21X1_220 ( );
FILL FILL_1_OAI21X1_220 ( );
FILL FILL_2_OAI21X1_220 ( );
FILL FILL_3_OAI21X1_220 ( );
FILL FILL_4_OAI21X1_220 ( );
FILL FILL_5_OAI21X1_220 ( );
FILL FILL_6_OAI21X1_220 ( );
FILL FILL_7_OAI21X1_220 ( );
FILL FILL_8_OAI21X1_220 ( );
FILL FILL_0_AOI21X1_24 ( );
FILL FILL_1_AOI21X1_24 ( );
FILL FILL_2_AOI21X1_24 ( );
FILL FILL_3_AOI21X1_24 ( );
FILL FILL_4_AOI21X1_24 ( );
FILL FILL_5_AOI21X1_24 ( );
FILL FILL_6_AOI21X1_24 ( );
FILL FILL_7_AOI21X1_24 ( );
FILL FILL_8_AOI21X1_24 ( );
FILL FILL_0_NAND3X1_37 ( );
FILL FILL_1_NAND3X1_37 ( );
FILL FILL_2_NAND3X1_37 ( );
FILL FILL_3_NAND3X1_37 ( );
FILL FILL_4_NAND3X1_37 ( );
FILL FILL_5_NAND3X1_37 ( );
FILL FILL_6_NAND3X1_37 ( );
FILL FILL_7_NAND3X1_37 ( );
FILL FILL_8_NAND3X1_37 ( );
FILL FILL_0_OAI21X1_159 ( );
FILL FILL_1_OAI21X1_159 ( );
FILL FILL_2_OAI21X1_159 ( );
FILL FILL_3_OAI21X1_159 ( );
FILL FILL_4_OAI21X1_159 ( );
FILL FILL_5_OAI21X1_159 ( );
FILL FILL_6_OAI21X1_159 ( );
FILL FILL_7_OAI21X1_159 ( );
FILL FILL_8_OAI21X1_159 ( );
FILL FILL_0_AOI21X1_22 ( );
FILL FILL_1_AOI21X1_22 ( );
FILL FILL_2_AOI21X1_22 ( );
FILL FILL_3_AOI21X1_22 ( );
FILL FILL_4_AOI21X1_22 ( );
FILL FILL_5_AOI21X1_22 ( );
FILL FILL_6_AOI21X1_22 ( );
FILL FILL_7_AOI21X1_22 ( );
FILL FILL_8_AOI21X1_22 ( );
FILL FILL_0_NAND3X1_47 ( );
FILL FILL_1_NAND3X1_47 ( );
FILL FILL_2_NAND3X1_47 ( );
FILL FILL_3_NAND3X1_47 ( );
FILL FILL_4_NAND3X1_47 ( );
FILL FILL_5_NAND3X1_47 ( );
FILL FILL_6_NAND3X1_47 ( );
FILL FILL_7_NAND3X1_47 ( );
FILL FILL_8_NAND3X1_47 ( );
FILL FILL_0_NAND2X1_206 ( );
FILL FILL_1_NAND2X1_206 ( );
FILL FILL_2_NAND2X1_206 ( );
FILL FILL_3_NAND2X1_206 ( );
FILL FILL_4_NAND2X1_206 ( );
FILL FILL_5_NAND2X1_206 ( );
FILL FILL_6_NAND2X1_206 ( );
FILL FILL_0_OAI21X1_215 ( );
FILL FILL_1_OAI21X1_215 ( );
FILL FILL_2_OAI21X1_215 ( );
FILL FILL_3_OAI21X1_215 ( );
FILL FILL_4_OAI21X1_215 ( );
FILL FILL_5_OAI21X1_215 ( );
FILL FILL_6_OAI21X1_215 ( );
FILL FILL_7_OAI21X1_215 ( );
FILL FILL_8_OAI21X1_215 ( );
FILL FILL_0_AOI21X1_25 ( );
FILL FILL_1_AOI21X1_25 ( );
FILL FILL_2_AOI21X1_25 ( );
FILL FILL_3_AOI21X1_25 ( );
FILL FILL_4_AOI21X1_25 ( );
FILL FILL_5_AOI21X1_25 ( );
FILL FILL_6_AOI21X1_25 ( );
FILL FILL_7_AOI21X1_25 ( );
FILL FILL_8_AOI21X1_25 ( );
FILL FILL_0_AOI22X1_8 ( );
FILL FILL_1_AOI22X1_8 ( );
FILL FILL_2_AOI22X1_8 ( );
FILL FILL_3_AOI22X1_8 ( );
FILL FILL_4_AOI22X1_8 ( );
FILL FILL_5_AOI22X1_8 ( );
FILL FILL_6_AOI22X1_8 ( );
FILL FILL_7_AOI22X1_8 ( );
FILL FILL_8_AOI22X1_8 ( );
FILL FILL_9_AOI22X1_8 ( );
FILL FILL_10_AOI22X1_8 ( );
FILL FILL_0_NAND2X1_207 ( );
FILL FILL_1_NAND2X1_207 ( );
FILL FILL_2_NAND2X1_207 ( );
FILL FILL_3_NAND2X1_207 ( );
FILL FILL_4_NAND2X1_207 ( );
FILL FILL_5_NAND2X1_207 ( );
FILL FILL_6_NAND2X1_207 ( );
FILL FILL_0_NAND3X1_96 ( );
FILL FILL_1_NAND3X1_96 ( );
FILL FILL_2_NAND3X1_96 ( );
FILL FILL_3_NAND3X1_96 ( );
FILL FILL_4_NAND3X1_96 ( );
FILL FILL_5_NAND3X1_96 ( );
FILL FILL_6_NAND3X1_96 ( );
FILL FILL_7_NAND3X1_96 ( );
FILL FILL_8_NAND3X1_96 ( );
FILL FILL_0_NAND3X1_91 ( );
FILL FILL_1_NAND3X1_91 ( );
FILL FILL_2_NAND3X1_91 ( );
FILL FILL_3_NAND3X1_91 ( );
FILL FILL_4_NAND3X1_91 ( );
FILL FILL_5_NAND3X1_91 ( );
FILL FILL_6_NAND3X1_91 ( );
FILL FILL_7_NAND3X1_91 ( );
FILL FILL_8_NAND3X1_91 ( );
FILL FILL_9_NAND3X1_91 ( );
FILL FILL_0_NAND3X1_107 ( );
FILL FILL_1_NAND3X1_107 ( );
FILL FILL_2_NAND3X1_107 ( );
FILL FILL_3_NAND3X1_107 ( );
FILL FILL_4_NAND3X1_107 ( );
FILL FILL_5_NAND3X1_107 ( );
FILL FILL_6_NAND3X1_107 ( );
FILL FILL_7_NAND3X1_107 ( );
FILL FILL_8_NAND3X1_107 ( );
FILL FILL_0_OAI21X1_127 ( );
FILL FILL_1_OAI21X1_127 ( );
FILL FILL_2_OAI21X1_127 ( );
FILL FILL_3_OAI21X1_127 ( );
FILL FILL_4_OAI21X1_127 ( );
FILL FILL_5_OAI21X1_127 ( );
FILL FILL_6_OAI21X1_127 ( );
FILL FILL_7_OAI21X1_127 ( );
FILL FILL_8_OAI21X1_127 ( );
FILL FILL_0_DFFSR_84 ( );
FILL FILL_1_DFFSR_84 ( );
FILL FILL_2_DFFSR_84 ( );
FILL FILL_3_DFFSR_84 ( );
FILL FILL_4_DFFSR_84 ( );
FILL FILL_5_DFFSR_84 ( );
FILL FILL_6_DFFSR_84 ( );
FILL FILL_7_DFFSR_84 ( );
FILL FILL_8_DFFSR_84 ( );
FILL FILL_9_DFFSR_84 ( );
FILL FILL_10_DFFSR_84 ( );
FILL FILL_11_DFFSR_84 ( );
FILL FILL_12_DFFSR_84 ( );
FILL FILL_13_DFFSR_84 ( );
FILL FILL_14_DFFSR_84 ( );
FILL FILL_15_DFFSR_84 ( );
FILL FILL_16_DFFSR_84 ( );
FILL FILL_17_DFFSR_84 ( );
FILL FILL_18_DFFSR_84 ( );
FILL FILL_19_DFFSR_84 ( );
FILL FILL_20_DFFSR_84 ( );
FILL FILL_21_DFFSR_84 ( );
FILL FILL_22_DFFSR_84 ( );
FILL FILL_23_DFFSR_84 ( );
FILL FILL_24_DFFSR_84 ( );
FILL FILL_25_DFFSR_84 ( );
FILL FILL_26_DFFSR_84 ( );
FILL FILL_27_DFFSR_84 ( );
FILL FILL_28_DFFSR_84 ( );
FILL FILL_29_DFFSR_84 ( );
FILL FILL_30_DFFSR_84 ( );
FILL FILL_31_DFFSR_84 ( );
FILL FILL_32_DFFSR_84 ( );
FILL FILL_33_DFFSR_84 ( );
FILL FILL_34_DFFSR_84 ( );
FILL FILL_35_DFFSR_84 ( );
FILL FILL_36_DFFSR_84 ( );
FILL FILL_37_DFFSR_84 ( );
FILL FILL_38_DFFSR_84 ( );
FILL FILL_39_DFFSR_84 ( );
FILL FILL_40_DFFSR_84 ( );
FILL FILL_41_DFFSR_84 ( );
FILL FILL_42_DFFSR_84 ( );
FILL FILL_43_DFFSR_84 ( );
FILL FILL_44_DFFSR_84 ( );
FILL FILL_45_DFFSR_84 ( );
FILL FILL_46_DFFSR_84 ( );
FILL FILL_47_DFFSR_84 ( );
FILL FILL_48_DFFSR_84 ( );
FILL FILL_49_DFFSR_84 ( );
FILL FILL_50_DFFSR_84 ( );
FILL FILL_51_DFFSR_84 ( );
FILL FILL_0_DFFSR_69 ( );
FILL FILL_1_DFFSR_69 ( );
FILL FILL_2_DFFSR_69 ( );
FILL FILL_3_DFFSR_69 ( );
FILL FILL_4_DFFSR_69 ( );
FILL FILL_5_DFFSR_69 ( );
FILL FILL_6_DFFSR_69 ( );
FILL FILL_7_DFFSR_69 ( );
FILL FILL_8_DFFSR_69 ( );
FILL FILL_9_DFFSR_69 ( );
FILL FILL_10_DFFSR_69 ( );
FILL FILL_11_DFFSR_69 ( );
FILL FILL_12_DFFSR_69 ( );
FILL FILL_13_DFFSR_69 ( );
FILL FILL_14_DFFSR_69 ( );
FILL FILL_15_DFFSR_69 ( );
FILL FILL_16_DFFSR_69 ( );
FILL FILL_17_DFFSR_69 ( );
FILL FILL_18_DFFSR_69 ( );
FILL FILL_19_DFFSR_69 ( );
FILL FILL_20_DFFSR_69 ( );
FILL FILL_21_DFFSR_69 ( );
FILL FILL_22_DFFSR_69 ( );
FILL FILL_23_DFFSR_69 ( );
FILL FILL_24_DFFSR_69 ( );
FILL FILL_25_DFFSR_69 ( );
FILL FILL_26_DFFSR_69 ( );
FILL FILL_27_DFFSR_69 ( );
FILL FILL_28_DFFSR_69 ( );
FILL FILL_29_DFFSR_69 ( );
FILL FILL_30_DFFSR_69 ( );
FILL FILL_31_DFFSR_69 ( );
FILL FILL_32_DFFSR_69 ( );
FILL FILL_33_DFFSR_69 ( );
FILL FILL_34_DFFSR_69 ( );
FILL FILL_35_DFFSR_69 ( );
FILL FILL_36_DFFSR_69 ( );
FILL FILL_37_DFFSR_69 ( );
FILL FILL_38_DFFSR_69 ( );
FILL FILL_39_DFFSR_69 ( );
FILL FILL_40_DFFSR_69 ( );
FILL FILL_41_DFFSR_69 ( );
FILL FILL_42_DFFSR_69 ( );
FILL FILL_43_DFFSR_69 ( );
FILL FILL_44_DFFSR_69 ( );
FILL FILL_45_DFFSR_69 ( );
FILL FILL_46_DFFSR_69 ( );
FILL FILL_47_DFFSR_69 ( );
FILL FILL_48_DFFSR_69 ( );
FILL FILL_49_DFFSR_69 ( );
FILL FILL_50_DFFSR_69 ( );
FILL FILL_0_CLKBUF1_12 ( );
FILL FILL_1_CLKBUF1_12 ( );
FILL FILL_2_CLKBUF1_12 ( );
FILL FILL_3_CLKBUF1_12 ( );
FILL FILL_4_CLKBUF1_12 ( );
FILL FILL_5_CLKBUF1_12 ( );
FILL FILL_6_CLKBUF1_12 ( );
FILL FILL_7_CLKBUF1_12 ( );
FILL FILL_8_CLKBUF1_12 ( );
FILL FILL_9_CLKBUF1_12 ( );
FILL FILL_10_CLKBUF1_12 ( );
FILL FILL_11_CLKBUF1_12 ( );
FILL FILL_12_CLKBUF1_12 ( );
FILL FILL_13_CLKBUF1_12 ( );
FILL FILL_14_CLKBUF1_12 ( );
FILL FILL_15_CLKBUF1_12 ( );
FILL FILL_16_CLKBUF1_12 ( );
FILL FILL_17_CLKBUF1_12 ( );
FILL FILL_18_CLKBUF1_12 ( );
FILL FILL_19_CLKBUF1_12 ( );
FILL FILL_20_CLKBUF1_12 ( );
FILL FILL_21_CLKBUF1_12 ( );
FILL FILL_0_INVX1_16 ( );
FILL FILL_1_INVX1_16 ( );
FILL FILL_2_INVX1_16 ( );
FILL FILL_3_INVX1_16 ( );
FILL FILL_0_OAI21X1_14 ( );
FILL FILL_1_OAI21X1_14 ( );
FILL FILL_2_OAI21X1_14 ( );
FILL FILL_3_OAI21X1_14 ( );
FILL FILL_4_OAI21X1_14 ( );
FILL FILL_5_OAI21X1_14 ( );
FILL FILL_6_OAI21X1_14 ( );
FILL FILL_7_OAI21X1_14 ( );
FILL FILL_8_OAI21X1_14 ( );
FILL FILL_9_OAI21X1_14 ( );
FILL FILL_0_NAND2X1_14 ( );
FILL FILL_1_NAND2X1_14 ( );
FILL FILL_2_NAND2X1_14 ( );
FILL FILL_3_NAND2X1_14 ( );
FILL FILL_4_NAND2X1_14 ( );
FILL FILL_5_NAND2X1_14 ( );
FILL FILL_6_NAND2X1_14 ( );
FILL FILL_0_AOI21X1_47 ( );
FILL FILL_1_AOI21X1_47 ( );
FILL FILL_2_AOI21X1_47 ( );
FILL FILL_3_AOI21X1_47 ( );
FILL FILL_4_AOI21X1_47 ( );
FILL FILL_5_AOI21X1_47 ( );
FILL FILL_6_AOI21X1_47 ( );
FILL FILL_7_AOI21X1_47 ( );
FILL FILL_8_AOI21X1_47 ( );
FILL FILL_0_DFFSR_158 ( );
FILL FILL_1_DFFSR_158 ( );
FILL FILL_2_DFFSR_158 ( );
FILL FILL_3_DFFSR_158 ( );
FILL FILL_4_DFFSR_158 ( );
FILL FILL_5_DFFSR_158 ( );
FILL FILL_6_DFFSR_158 ( );
FILL FILL_7_DFFSR_158 ( );
FILL FILL_8_DFFSR_158 ( );
FILL FILL_9_DFFSR_158 ( );
FILL FILL_10_DFFSR_158 ( );
FILL FILL_11_DFFSR_158 ( );
FILL FILL_12_DFFSR_158 ( );
FILL FILL_13_DFFSR_158 ( );
FILL FILL_14_DFFSR_158 ( );
FILL FILL_15_DFFSR_158 ( );
FILL FILL_16_DFFSR_158 ( );
FILL FILL_17_DFFSR_158 ( );
FILL FILL_18_DFFSR_158 ( );
FILL FILL_19_DFFSR_158 ( );
FILL FILL_20_DFFSR_158 ( );
FILL FILL_21_DFFSR_158 ( );
FILL FILL_22_DFFSR_158 ( );
FILL FILL_23_DFFSR_158 ( );
FILL FILL_24_DFFSR_158 ( );
FILL FILL_25_DFFSR_158 ( );
FILL FILL_26_DFFSR_158 ( );
FILL FILL_27_DFFSR_158 ( );
FILL FILL_28_DFFSR_158 ( );
FILL FILL_29_DFFSR_158 ( );
FILL FILL_30_DFFSR_158 ( );
FILL FILL_31_DFFSR_158 ( );
FILL FILL_32_DFFSR_158 ( );
FILL FILL_33_DFFSR_158 ( );
FILL FILL_34_DFFSR_158 ( );
FILL FILL_35_DFFSR_158 ( );
FILL FILL_36_DFFSR_158 ( );
FILL FILL_37_DFFSR_158 ( );
FILL FILL_38_DFFSR_158 ( );
FILL FILL_39_DFFSR_158 ( );
FILL FILL_40_DFFSR_158 ( );
FILL FILL_41_DFFSR_158 ( );
FILL FILL_42_DFFSR_158 ( );
FILL FILL_43_DFFSR_158 ( );
FILL FILL_44_DFFSR_158 ( );
FILL FILL_45_DFFSR_158 ( );
FILL FILL_46_DFFSR_158 ( );
FILL FILL_47_DFFSR_158 ( );
FILL FILL_48_DFFSR_158 ( );
FILL FILL_49_DFFSR_158 ( );
FILL FILL_50_DFFSR_158 ( );
FILL FILL_0_INVX1_26 ( );
FILL FILL_1_INVX1_26 ( );
FILL FILL_2_INVX1_26 ( );
FILL FILL_3_INVX1_26 ( );
FILL FILL_4_INVX1_26 ( );
FILL FILL_0_CLKBUF1_14 ( );
FILL FILL_1_CLKBUF1_14 ( );
FILL FILL_2_CLKBUF1_14 ( );
FILL FILL_3_CLKBUF1_14 ( );
FILL FILL_4_CLKBUF1_14 ( );
FILL FILL_5_CLKBUF1_14 ( );
FILL FILL_6_CLKBUF1_14 ( );
FILL FILL_7_CLKBUF1_14 ( );
FILL FILL_8_CLKBUF1_14 ( );
FILL FILL_9_CLKBUF1_14 ( );
FILL FILL_10_CLKBUF1_14 ( );
FILL FILL_11_CLKBUF1_14 ( );
FILL FILL_12_CLKBUF1_14 ( );
FILL FILL_13_CLKBUF1_14 ( );
FILL FILL_14_CLKBUF1_14 ( );
FILL FILL_15_CLKBUF1_14 ( );
FILL FILL_16_CLKBUF1_14 ( );
FILL FILL_17_CLKBUF1_14 ( );
FILL FILL_18_CLKBUF1_14 ( );
FILL FILL_19_CLKBUF1_14 ( );
FILL FILL_0_OAI21X1_174 ( );
FILL FILL_1_OAI21X1_174 ( );
FILL FILL_2_OAI21X1_174 ( );
FILL FILL_3_OAI21X1_174 ( );
FILL FILL_4_OAI21X1_174 ( );
FILL FILL_5_OAI21X1_174 ( );
FILL FILL_6_OAI21X1_174 ( );
FILL FILL_7_OAI21X1_174 ( );
FILL FILL_8_OAI21X1_174 ( );
FILL FILL_9_OAI21X1_174 ( );
FILL FILL_0_INVX1_209 ( );
FILL FILL_1_INVX1_209 ( );
FILL FILL_2_INVX1_209 ( );
FILL FILL_3_INVX1_209 ( );
FILL FILL_0_DFFPOSX1_24 ( );
FILL FILL_1_DFFPOSX1_24 ( );
FILL FILL_2_DFFPOSX1_24 ( );
FILL FILL_3_DFFPOSX1_24 ( );
FILL FILL_4_DFFPOSX1_24 ( );
FILL FILL_5_DFFPOSX1_24 ( );
FILL FILL_6_DFFPOSX1_24 ( );
FILL FILL_7_DFFPOSX1_24 ( );
FILL FILL_8_DFFPOSX1_24 ( );
FILL FILL_9_DFFPOSX1_24 ( );
FILL FILL_10_DFFPOSX1_24 ( );
FILL FILL_11_DFFPOSX1_24 ( );
FILL FILL_12_DFFPOSX1_24 ( );
FILL FILL_13_DFFPOSX1_24 ( );
FILL FILL_14_DFFPOSX1_24 ( );
FILL FILL_15_DFFPOSX1_24 ( );
FILL FILL_16_DFFPOSX1_24 ( );
FILL FILL_17_DFFPOSX1_24 ( );
FILL FILL_18_DFFPOSX1_24 ( );
FILL FILL_19_DFFPOSX1_24 ( );
FILL FILL_20_DFFPOSX1_24 ( );
FILL FILL_21_DFFPOSX1_24 ( );
FILL FILL_22_DFFPOSX1_24 ( );
FILL FILL_23_DFFPOSX1_24 ( );
FILL FILL_24_DFFPOSX1_24 ( );
FILL FILL_25_DFFPOSX1_24 ( );
FILL FILL_26_DFFPOSX1_24 ( );
FILL FILL_27_DFFPOSX1_24 ( );
FILL FILL_0_NAND2X1_215 ( );
FILL FILL_1_NAND2X1_215 ( );
FILL FILL_2_NAND2X1_215 ( );
FILL FILL_3_NAND2X1_215 ( );
FILL FILL_4_NAND2X1_215 ( );
FILL FILL_5_NAND2X1_215 ( );
FILL FILL_6_NAND2X1_215 ( );
FILL FILL_0_NAND3X1_63 ( );
FILL FILL_1_NAND3X1_63 ( );
FILL FILL_2_NAND3X1_63 ( );
FILL FILL_3_NAND3X1_63 ( );
FILL FILL_4_NAND3X1_63 ( );
FILL FILL_5_NAND3X1_63 ( );
FILL FILL_6_NAND3X1_63 ( );
FILL FILL_7_NAND3X1_63 ( );
FILL FILL_8_NAND3X1_63 ( );
FILL FILL_0_NOR2X1_8 ( );
FILL FILL_1_NOR2X1_8 ( );
FILL FILL_2_NOR2X1_8 ( );
FILL FILL_3_NOR2X1_8 ( );
FILL FILL_4_NOR2X1_8 ( );
FILL FILL_5_NOR2X1_8 ( );
FILL FILL_6_NOR2X1_8 ( );
FILL FILL_0_NAND3X1_40 ( );
FILL FILL_1_NAND3X1_40 ( );
FILL FILL_2_NAND3X1_40 ( );
FILL FILL_3_NAND3X1_40 ( );
FILL FILL_4_NAND3X1_40 ( );
FILL FILL_5_NAND3X1_40 ( );
FILL FILL_6_NAND3X1_40 ( );
FILL FILL_7_NAND3X1_40 ( );
FILL FILL_8_NAND3X1_40 ( );
FILL FILL_0_INVX1_241 ( );
FILL FILL_1_INVX1_241 ( );
FILL FILL_2_INVX1_241 ( );
FILL FILL_3_INVX1_241 ( );
FILL FILL_0_NAND3X1_42 ( );
FILL FILL_1_NAND3X1_42 ( );
FILL FILL_2_NAND3X1_42 ( );
FILL FILL_3_NAND3X1_42 ( );
FILL FILL_4_NAND3X1_42 ( );
FILL FILL_5_NAND3X1_42 ( );
FILL FILL_6_NAND3X1_42 ( );
FILL FILL_7_NAND3X1_42 ( );
FILL FILL_8_NAND3X1_42 ( );
FILL FILL_0_NAND3X1_48 ( );
FILL FILL_1_NAND3X1_48 ( );
FILL FILL_2_NAND3X1_48 ( );
FILL FILL_3_NAND3X1_48 ( );
FILL FILL_4_NAND3X1_48 ( );
FILL FILL_5_NAND3X1_48 ( );
FILL FILL_6_NAND3X1_48 ( );
FILL FILL_7_NAND3X1_48 ( );
FILL FILL_8_NAND3X1_48 ( );
FILL FILL_9_NAND3X1_48 ( );
FILL FILL_0_NAND3X1_41 ( );
FILL FILL_1_NAND3X1_41 ( );
FILL FILL_2_NAND3X1_41 ( );
FILL FILL_3_NAND3X1_41 ( );
FILL FILL_4_NAND3X1_41 ( );
FILL FILL_5_NAND3X1_41 ( );
FILL FILL_6_NAND3X1_41 ( );
FILL FILL_7_NAND3X1_41 ( );
FILL FILL_8_NAND3X1_41 ( );
FILL FILL_0_AOI22X1_7 ( );
FILL FILL_1_AOI22X1_7 ( );
FILL FILL_2_AOI22X1_7 ( );
FILL FILL_3_AOI22X1_7 ( );
FILL FILL_4_AOI22X1_7 ( );
FILL FILL_5_AOI22X1_7 ( );
FILL FILL_6_AOI22X1_7 ( );
FILL FILL_7_AOI22X1_7 ( );
FILL FILL_8_AOI22X1_7 ( );
FILL FILL_9_AOI22X1_7 ( );
FILL FILL_10_AOI22X1_7 ( );
FILL FILL_0_INVX1_231 ( );
FILL FILL_1_INVX1_231 ( );
FILL FILL_2_INVX1_231 ( );
FILL FILL_3_INVX1_231 ( );
FILL FILL_0_BUFX2_2 ( );
FILL FILL_1_BUFX2_2 ( );
FILL FILL_2_BUFX2_2 ( );
FILL FILL_3_BUFX2_2 ( );
FILL FILL_4_BUFX2_2 ( );
FILL FILL_5_BUFX2_2 ( );
FILL FILL_6_BUFX2_2 ( );
FILL FILL_0_NAND3X1_62 ( );
FILL FILL_1_NAND3X1_62 ( );
FILL FILL_2_NAND3X1_62 ( );
FILL FILL_3_NAND3X1_62 ( );
FILL FILL_4_NAND3X1_62 ( );
FILL FILL_5_NAND3X1_62 ( );
FILL FILL_6_NAND3X1_62 ( );
FILL FILL_7_NAND3X1_62 ( );
FILL FILL_8_NAND3X1_62 ( );
FILL FILL_0_NAND3X1_73 ( );
FILL FILL_1_NAND3X1_73 ( );
FILL FILL_2_NAND3X1_73 ( );
FILL FILL_3_NAND3X1_73 ( );
FILL FILL_4_NAND3X1_73 ( );
FILL FILL_5_NAND3X1_73 ( );
FILL FILL_6_NAND3X1_73 ( );
FILL FILL_7_NAND3X1_73 ( );
FILL FILL_8_NAND3X1_73 ( );
FILL FILL_9_NAND3X1_73 ( );
FILL FILL_0_AOI21X1_16 ( );
FILL FILL_1_AOI21X1_16 ( );
FILL FILL_2_AOI21X1_16 ( );
FILL FILL_3_AOI21X1_16 ( );
FILL FILL_4_AOI21X1_16 ( );
FILL FILL_5_AOI21X1_16 ( );
FILL FILL_6_AOI21X1_16 ( );
FILL FILL_7_AOI21X1_16 ( );
FILL FILL_8_AOI21X1_16 ( );
FILL FILL_9_AOI21X1_16 ( );
FILL FILL_0_INVX1_258 ( );
FILL FILL_1_INVX1_258 ( );
FILL FILL_2_INVX1_258 ( );
FILL FILL_3_INVX1_258 ( );
FILL FILL_4_INVX1_258 ( );
FILL FILL_0_NAND3X1_92 ( );
FILL FILL_1_NAND3X1_92 ( );
FILL FILL_2_NAND3X1_92 ( );
FILL FILL_3_NAND3X1_92 ( );
FILL FILL_4_NAND3X1_92 ( );
FILL FILL_5_NAND3X1_92 ( );
FILL FILL_6_NAND3X1_92 ( );
FILL FILL_7_NAND3X1_92 ( );
FILL FILL_8_NAND3X1_92 ( );
FILL FILL_0_NAND3X1_89 ( );
FILL FILL_1_NAND3X1_89 ( );
FILL FILL_2_NAND3X1_89 ( );
FILL FILL_3_NAND3X1_89 ( );
FILL FILL_4_NAND3X1_89 ( );
FILL FILL_5_NAND3X1_89 ( );
FILL FILL_6_NAND3X1_89 ( );
FILL FILL_7_NAND3X1_89 ( );
FILL FILL_8_NAND3X1_89 ( );
FILL FILL_0_AOI21X1_32 ( );
FILL FILL_1_AOI21X1_32 ( );
FILL FILL_2_AOI21X1_32 ( );
FILL FILL_3_AOI21X1_32 ( );
FILL FILL_4_AOI21X1_32 ( );
FILL FILL_5_AOI21X1_32 ( );
FILL FILL_6_AOI21X1_32 ( );
FILL FILL_7_AOI21X1_32 ( );
FILL FILL_8_AOI21X1_32 ( );
FILL FILL_9_AOI21X1_32 ( );
FILL FILL_0_OR2X2_3 ( );
FILL FILL_1_OR2X2_3 ( );
FILL FILL_2_OR2X2_3 ( );
FILL FILL_3_OR2X2_3 ( );
FILL FILL_4_OR2X2_3 ( );
FILL FILL_5_OR2X2_3 ( );
FILL FILL_6_OR2X2_3 ( );
FILL FILL_7_OR2X2_3 ( );
FILL FILL_8_OR2X2_3 ( );
FILL FILL_0_OAI21X1_97 ( );
FILL FILL_1_OAI21X1_97 ( );
FILL FILL_2_OAI21X1_97 ( );
FILL FILL_3_OAI21X1_97 ( );
FILL FILL_4_OAI21X1_97 ( );
FILL FILL_5_OAI21X1_97 ( );
FILL FILL_6_OAI21X1_97 ( );
FILL FILL_7_OAI21X1_97 ( );
FILL FILL_8_OAI21X1_97 ( );
FILL FILL_9_OAI21X1_97 ( );
FILL FILL_0_INVX1_110 ( );
FILL FILL_1_INVX1_110 ( );
FILL FILL_2_INVX1_110 ( );
FILL FILL_3_INVX1_110 ( );
FILL FILL_0_NAND2X1_97 ( );
FILL FILL_1_NAND2X1_97 ( );
FILL FILL_2_NAND2X1_97 ( );
FILL FILL_3_NAND2X1_97 ( );
FILL FILL_4_NAND2X1_97 ( );
FILL FILL_5_NAND2X1_97 ( );
FILL FILL_6_NAND2X1_97 ( );
FILL FILL_0_INVX1_143 ( );
FILL FILL_1_INVX1_143 ( );
FILL FILL_2_INVX1_143 ( );
FILL FILL_3_INVX1_143 ( );
FILL FILL_4_INVX1_143 ( );
FILL FILL_0_CLKBUF1_6 ( );
FILL FILL_1_CLKBUF1_6 ( );
FILL FILL_2_CLKBUF1_6 ( );
FILL FILL_3_CLKBUF1_6 ( );
FILL FILL_4_CLKBUF1_6 ( );
FILL FILL_5_CLKBUF1_6 ( );
FILL FILL_6_CLKBUF1_6 ( );
FILL FILL_7_CLKBUF1_6 ( );
FILL FILL_8_CLKBUF1_6 ( );
FILL FILL_9_CLKBUF1_6 ( );
FILL FILL_10_CLKBUF1_6 ( );
FILL FILL_11_CLKBUF1_6 ( );
FILL FILL_12_CLKBUF1_6 ( );
FILL FILL_13_CLKBUF1_6 ( );
FILL FILL_14_CLKBUF1_6 ( );
FILL FILL_15_CLKBUF1_6 ( );
FILL FILL_16_CLKBUF1_6 ( );
FILL FILL_17_CLKBUF1_6 ( );
FILL FILL_18_CLKBUF1_6 ( );
FILL FILL_19_CLKBUF1_6 ( );
FILL FILL_20_CLKBUF1_6 ( );
FILL FILL_21_CLKBUF1_6 ( );
FILL FILL_0_INVX1_371 ( );
FILL FILL_1_INVX1_371 ( );
FILL FILL_2_INVX1_371 ( );
FILL FILL_3_INVX1_371 ( );
FILL FILL_0_NAND2X1_92 ( );
FILL FILL_1_NAND2X1_92 ( );
FILL FILL_2_NAND2X1_92 ( );
FILL FILL_3_NAND2X1_92 ( );
FILL FILL_4_NAND2X1_92 ( );
FILL FILL_5_NAND2X1_92 ( );
FILL FILL_6_NAND2X1_92 ( );
FILL FILL_0_OAI21X1_92 ( );
FILL FILL_1_OAI21X1_92 ( );
FILL FILL_2_OAI21X1_92 ( );
FILL FILL_3_OAI21X1_92 ( );
FILL FILL_4_OAI21X1_92 ( );
FILL FILL_5_OAI21X1_92 ( );
FILL FILL_6_OAI21X1_92 ( );
FILL FILL_7_OAI21X1_92 ( );
FILL FILL_8_OAI21X1_92 ( );
FILL FILL_0_INVX1_104 ( );
FILL FILL_1_INVX1_104 ( );
FILL FILL_2_INVX1_104 ( );
FILL FILL_3_INVX1_104 ( );
FILL FILL_4_INVX1_104 ( );
FILL FILL_0_NAND2X1_91 ( );
FILL FILL_1_NAND2X1_91 ( );
FILL FILL_2_NAND2X1_91 ( );
FILL FILL_3_NAND2X1_91 ( );
FILL FILL_4_NAND2X1_91 ( );
FILL FILL_5_NAND2X1_91 ( );
FILL FILL_6_NAND2X1_91 ( );
FILL FILL_0_DFFSR_152 ( );
FILL FILL_1_DFFSR_152 ( );
FILL FILL_2_DFFSR_152 ( );
FILL FILL_3_DFFSR_152 ( );
FILL FILL_4_DFFSR_152 ( );
FILL FILL_5_DFFSR_152 ( );
FILL FILL_6_DFFSR_152 ( );
FILL FILL_7_DFFSR_152 ( );
FILL FILL_8_DFFSR_152 ( );
FILL FILL_9_DFFSR_152 ( );
FILL FILL_10_DFFSR_152 ( );
FILL FILL_11_DFFSR_152 ( );
FILL FILL_12_DFFSR_152 ( );
FILL FILL_13_DFFSR_152 ( );
FILL FILL_14_DFFSR_152 ( );
FILL FILL_15_DFFSR_152 ( );
FILL FILL_16_DFFSR_152 ( );
FILL FILL_17_DFFSR_152 ( );
FILL FILL_18_DFFSR_152 ( );
FILL FILL_19_DFFSR_152 ( );
FILL FILL_20_DFFSR_152 ( );
FILL FILL_21_DFFSR_152 ( );
FILL FILL_22_DFFSR_152 ( );
FILL FILL_23_DFFSR_152 ( );
FILL FILL_24_DFFSR_152 ( );
FILL FILL_25_DFFSR_152 ( );
FILL FILL_26_DFFSR_152 ( );
FILL FILL_27_DFFSR_152 ( );
FILL FILL_28_DFFSR_152 ( );
FILL FILL_29_DFFSR_152 ( );
FILL FILL_30_DFFSR_152 ( );
FILL FILL_31_DFFSR_152 ( );
FILL FILL_32_DFFSR_152 ( );
FILL FILL_33_DFFSR_152 ( );
FILL FILL_34_DFFSR_152 ( );
FILL FILL_35_DFFSR_152 ( );
FILL FILL_36_DFFSR_152 ( );
FILL FILL_37_DFFSR_152 ( );
FILL FILL_38_DFFSR_152 ( );
FILL FILL_39_DFFSR_152 ( );
FILL FILL_40_DFFSR_152 ( );
FILL FILL_41_DFFSR_152 ( );
FILL FILL_42_DFFSR_152 ( );
FILL FILL_43_DFFSR_152 ( );
FILL FILL_44_DFFSR_152 ( );
FILL FILL_45_DFFSR_152 ( );
FILL FILL_46_DFFSR_152 ( );
FILL FILL_47_DFFSR_152 ( );
FILL FILL_48_DFFSR_152 ( );
FILL FILL_49_DFFSR_152 ( );
FILL FILL_50_DFFSR_152 ( );
FILL FILL_0_INVX1_179 ( );
FILL FILL_1_INVX1_179 ( );
FILL FILL_2_INVX1_179 ( );
FILL FILL_3_INVX1_179 ( );
FILL FILL_4_INVX1_179 ( );
FILL FILL_0_BUFX2_5 ( );
FILL FILL_1_BUFX2_5 ( );
FILL FILL_2_BUFX2_5 ( );
FILL FILL_3_BUFX2_5 ( );
FILL FILL_4_BUFX2_5 ( );
FILL FILL_5_BUFX2_5 ( );
FILL FILL_6_BUFX2_5 ( );
FILL FILL_0_OAI21X1_135 ( );
FILL FILL_1_OAI21X1_135 ( );
FILL FILL_2_OAI21X1_135 ( );
FILL FILL_3_OAI21X1_135 ( );
FILL FILL_4_OAI21X1_135 ( );
FILL FILL_5_OAI21X1_135 ( );
FILL FILL_6_OAI21X1_135 ( );
FILL FILL_7_OAI21X1_135 ( );
FILL FILL_8_OAI21X1_135 ( );
FILL FILL_9_OAI21X1_135 ( );
FILL FILL_0_INVX1_152 ( );
FILL FILL_1_INVX1_152 ( );
FILL FILL_2_INVX1_152 ( );
FILL FILL_3_INVX1_152 ( );
FILL FILL_0_AND2X2_1 ( );
FILL FILL_1_AND2X2_1 ( );
FILL FILL_2_AND2X2_1 ( );
FILL FILL_3_AND2X2_1 ( );
FILL FILL_4_AND2X2_1 ( );
FILL FILL_5_AND2X2_1 ( );
FILL FILL_6_AND2X2_1 ( );
FILL FILL_7_AND2X2_1 ( );
FILL FILL_8_AND2X2_1 ( );
FILL FILL_9_AND2X2_1 ( );
FILL FILL_0_DFFPOSX1_21 ( );
FILL FILL_1_DFFPOSX1_21 ( );
FILL FILL_2_DFFPOSX1_21 ( );
FILL FILL_3_DFFPOSX1_21 ( );
FILL FILL_4_DFFPOSX1_21 ( );
FILL FILL_5_DFFPOSX1_21 ( );
FILL FILL_6_DFFPOSX1_21 ( );
FILL FILL_7_DFFPOSX1_21 ( );
FILL FILL_8_DFFPOSX1_21 ( );
FILL FILL_9_DFFPOSX1_21 ( );
FILL FILL_10_DFFPOSX1_21 ( );
FILL FILL_11_DFFPOSX1_21 ( );
FILL FILL_12_DFFPOSX1_21 ( );
FILL FILL_13_DFFPOSX1_21 ( );
FILL FILL_14_DFFPOSX1_21 ( );
FILL FILL_15_DFFPOSX1_21 ( );
FILL FILL_16_DFFPOSX1_21 ( );
FILL FILL_17_DFFPOSX1_21 ( );
FILL FILL_18_DFFPOSX1_21 ( );
FILL FILL_19_DFFPOSX1_21 ( );
FILL FILL_20_DFFPOSX1_21 ( );
FILL FILL_21_DFFPOSX1_21 ( );
FILL FILL_22_DFFPOSX1_21 ( );
FILL FILL_23_DFFPOSX1_21 ( );
FILL FILL_24_DFFPOSX1_21 ( );
FILL FILL_25_DFFPOSX1_21 ( );
FILL FILL_26_DFFPOSX1_21 ( );
FILL FILL_27_DFFPOSX1_21 ( );
FILL FILL_0_INVX1_191 ( );
FILL FILL_1_INVX1_191 ( );
FILL FILL_2_INVX1_191 ( );
FILL FILL_3_INVX1_191 ( );
FILL FILL_4_INVX1_191 ( );
FILL FILL_0_BUFX2_36 ( );
FILL FILL_1_BUFX2_36 ( );
FILL FILL_2_BUFX2_36 ( );
FILL FILL_3_BUFX2_36 ( );
FILL FILL_4_BUFX2_36 ( );
FILL FILL_5_BUFX2_36 ( );
FILL FILL_6_BUFX2_36 ( );
FILL FILL_0_BUFX2_42 ( );
FILL FILL_1_BUFX2_42 ( );
FILL FILL_2_BUFX2_42 ( );
FILL FILL_3_BUFX2_42 ( );
FILL FILL_4_BUFX2_42 ( );
FILL FILL_5_BUFX2_42 ( );
FILL FILL_6_BUFX2_42 ( );
FILL FILL_0_OAI21X1_23 ( );
FILL FILL_1_OAI21X1_23 ( );
FILL FILL_2_OAI21X1_23 ( );
FILL FILL_3_OAI21X1_23 ( );
FILL FILL_4_OAI21X1_23 ( );
FILL FILL_5_OAI21X1_23 ( );
FILL FILL_6_OAI21X1_23 ( );
FILL FILL_7_OAI21X1_23 ( );
FILL FILL_8_OAI21X1_23 ( );
FILL FILL_0_DFFSR_23 ( );
FILL FILL_1_DFFSR_23 ( );
FILL FILL_2_DFFSR_23 ( );
FILL FILL_3_DFFSR_23 ( );
FILL FILL_4_DFFSR_23 ( );
FILL FILL_5_DFFSR_23 ( );
FILL FILL_6_DFFSR_23 ( );
FILL FILL_7_DFFSR_23 ( );
FILL FILL_8_DFFSR_23 ( );
FILL FILL_9_DFFSR_23 ( );
FILL FILL_10_DFFSR_23 ( );
FILL FILL_11_DFFSR_23 ( );
FILL FILL_12_DFFSR_23 ( );
FILL FILL_13_DFFSR_23 ( );
FILL FILL_14_DFFSR_23 ( );
FILL FILL_15_DFFSR_23 ( );
FILL FILL_16_DFFSR_23 ( );
FILL FILL_17_DFFSR_23 ( );
FILL FILL_18_DFFSR_23 ( );
FILL FILL_19_DFFSR_23 ( );
FILL FILL_20_DFFSR_23 ( );
FILL FILL_21_DFFSR_23 ( );
FILL FILL_22_DFFSR_23 ( );
FILL FILL_23_DFFSR_23 ( );
FILL FILL_24_DFFSR_23 ( );
FILL FILL_25_DFFSR_23 ( );
FILL FILL_26_DFFSR_23 ( );
FILL FILL_27_DFFSR_23 ( );
FILL FILL_28_DFFSR_23 ( );
FILL FILL_29_DFFSR_23 ( );
FILL FILL_30_DFFSR_23 ( );
FILL FILL_31_DFFSR_23 ( );
FILL FILL_32_DFFSR_23 ( );
FILL FILL_33_DFFSR_23 ( );
FILL FILL_34_DFFSR_23 ( );
FILL FILL_35_DFFSR_23 ( );
FILL FILL_36_DFFSR_23 ( );
FILL FILL_37_DFFSR_23 ( );
FILL FILL_38_DFFSR_23 ( );
FILL FILL_39_DFFSR_23 ( );
FILL FILL_40_DFFSR_23 ( );
FILL FILL_41_DFFSR_23 ( );
FILL FILL_42_DFFSR_23 ( );
FILL FILL_43_DFFSR_23 ( );
FILL FILL_44_DFFSR_23 ( );
FILL FILL_45_DFFSR_23 ( );
FILL FILL_46_DFFSR_23 ( );
FILL FILL_47_DFFSR_23 ( );
FILL FILL_48_DFFSR_23 ( );
FILL FILL_49_DFFSR_23 ( );
FILL FILL_50_DFFSR_23 ( );
FILL FILL_0_AOI22X1_9 ( );
FILL FILL_1_AOI22X1_9 ( );
FILL FILL_2_AOI22X1_9 ( );
FILL FILL_3_AOI22X1_9 ( );
FILL FILL_4_AOI22X1_9 ( );
FILL FILL_5_AOI22X1_9 ( );
FILL FILL_6_AOI22X1_9 ( );
FILL FILL_7_AOI22X1_9 ( );
FILL FILL_8_AOI22X1_9 ( );
FILL FILL_9_AOI22X1_9 ( );
FILL FILL_10_AOI22X1_9 ( );
FILL FILL_11_AOI22X1_9 ( );
FILL FILL_0_AND2X2_10 ( );
FILL FILL_1_AND2X2_10 ( );
FILL FILL_2_AND2X2_10 ( );
FILL FILL_3_AND2X2_10 ( );
FILL FILL_4_AND2X2_10 ( );
FILL FILL_5_AND2X2_10 ( );
FILL FILL_6_AND2X2_10 ( );
FILL FILL_7_AND2X2_10 ( );
FILL FILL_8_AND2X2_10 ( );
FILL FILL_9_AND2X2_10 ( );
FILL FILL_0_NAND3X1_39 ( );
FILL FILL_1_NAND3X1_39 ( );
FILL FILL_2_NAND3X1_39 ( );
FILL FILL_3_NAND3X1_39 ( );
FILL FILL_4_NAND3X1_39 ( );
FILL FILL_5_NAND3X1_39 ( );
FILL FILL_6_NAND3X1_39 ( );
FILL FILL_7_NAND3X1_39 ( );
FILL FILL_8_NAND3X1_39 ( );
FILL FILL_9_NAND3X1_39 ( );
FILL FILL_0_NAND3X1_43 ( );
FILL FILL_1_NAND3X1_43 ( );
FILL FILL_2_NAND3X1_43 ( );
FILL FILL_3_NAND3X1_43 ( );
FILL FILL_4_NAND3X1_43 ( );
FILL FILL_5_NAND3X1_43 ( );
FILL FILL_6_NAND3X1_43 ( );
FILL FILL_7_NAND3X1_43 ( );
FILL FILL_8_NAND3X1_43 ( );
FILL FILL_0_NAND2X1_203 ( );
FILL FILL_1_NAND2X1_203 ( );
FILL FILL_2_NAND2X1_203 ( );
FILL FILL_3_NAND2X1_203 ( );
FILL FILL_4_NAND2X1_203 ( );
FILL FILL_5_NAND2X1_203 ( );
FILL FILL_6_NAND2X1_203 ( );
FILL FILL_0_NAND3X1_44 ( );
FILL FILL_1_NAND3X1_44 ( );
FILL FILL_2_NAND3X1_44 ( );
FILL FILL_3_NAND3X1_44 ( );
FILL FILL_4_NAND3X1_44 ( );
FILL FILL_5_NAND3X1_44 ( );
FILL FILL_6_NAND3X1_44 ( );
FILL FILL_7_NAND3X1_44 ( );
FILL FILL_8_NAND3X1_44 ( );
FILL FILL_9_NAND3X1_44 ( );
FILL FILL_0_AOI21X1_21 ( );
FILL FILL_1_AOI21X1_21 ( );
FILL FILL_2_AOI21X1_21 ( );
FILL FILL_3_AOI21X1_21 ( );
FILL FILL_4_AOI21X1_21 ( );
FILL FILL_5_AOI21X1_21 ( );
FILL FILL_6_AOI21X1_21 ( );
FILL FILL_7_AOI21X1_21 ( );
FILL FILL_8_AOI21X1_21 ( );
FILL FILL_9_AOI21X1_21 ( );
FILL FILL_0_AND2X2_8 ( );
FILL FILL_1_AND2X2_8 ( );
FILL FILL_2_AND2X2_8 ( );
FILL FILL_3_AND2X2_8 ( );
FILL FILL_4_AND2X2_8 ( );
FILL FILL_5_AND2X2_8 ( );
FILL FILL_6_AND2X2_8 ( );
FILL FILL_7_AND2X2_8 ( );
FILL FILL_8_AND2X2_8 ( );
FILL FILL_9_AND2X2_8 ( );
FILL FILL_0_AOI21X1_15 ( );
FILL FILL_1_AOI21X1_15 ( );
FILL FILL_2_AOI21X1_15 ( );
FILL FILL_3_AOI21X1_15 ( );
FILL FILL_4_AOI21X1_15 ( );
FILL FILL_5_AOI21X1_15 ( );
FILL FILL_6_AOI21X1_15 ( );
FILL FILL_7_AOI21X1_15 ( );
FILL FILL_8_AOI21X1_15 ( );
FILL FILL_0_OAI21X1_212 ( );
FILL FILL_1_OAI21X1_212 ( );
FILL FILL_2_OAI21X1_212 ( );
FILL FILL_3_OAI21X1_212 ( );
FILL FILL_4_OAI21X1_212 ( );
FILL FILL_5_OAI21X1_212 ( );
FILL FILL_6_OAI21X1_212 ( );
FILL FILL_7_OAI21X1_212 ( );
FILL FILL_8_OAI21X1_212 ( );
FILL FILL_0_OAI21X1_227 ( );
FILL FILL_1_OAI21X1_227 ( );
FILL FILL_2_OAI21X1_227 ( );
FILL FILL_3_OAI21X1_227 ( );
FILL FILL_4_OAI21X1_227 ( );
FILL FILL_5_OAI21X1_227 ( );
FILL FILL_6_OAI21X1_227 ( );
FILL FILL_7_OAI21X1_227 ( );
FILL FILL_8_OAI21X1_227 ( );
FILL FILL_0_AOI21X1_26 ( );
FILL FILL_1_AOI21X1_26 ( );
FILL FILL_2_AOI21X1_26 ( );
FILL FILL_3_AOI21X1_26 ( );
FILL FILL_4_AOI21X1_26 ( );
FILL FILL_5_AOI21X1_26 ( );
FILL FILL_6_AOI21X1_26 ( );
FILL FILL_7_AOI21X1_26 ( );
FILL FILL_8_AOI21X1_26 ( );
FILL FILL_0_OAI21X1_206 ( );
FILL FILL_1_OAI21X1_206 ( );
FILL FILL_2_OAI21X1_206 ( );
FILL FILL_3_OAI21X1_206 ( );
FILL FILL_4_OAI21X1_206 ( );
FILL FILL_5_OAI21X1_206 ( );
FILL FILL_6_OAI21X1_206 ( );
FILL FILL_7_OAI21X1_206 ( );
FILL FILL_8_OAI21X1_206 ( );
FILL FILL_0_NAND3X1_90 ( );
FILL FILL_1_NAND3X1_90 ( );
FILL FILL_2_NAND3X1_90 ( );
FILL FILL_3_NAND3X1_90 ( );
FILL FILL_4_NAND3X1_90 ( );
FILL FILL_5_NAND3X1_90 ( );
FILL FILL_6_NAND3X1_90 ( );
FILL FILL_7_NAND3X1_90 ( );
FILL FILL_8_NAND3X1_90 ( );
FILL FILL_0_NAND3X1_93 ( );
FILL FILL_1_NAND3X1_93 ( );
FILL FILL_2_NAND3X1_93 ( );
FILL FILL_3_NAND3X1_93 ( );
FILL FILL_4_NAND3X1_93 ( );
FILL FILL_5_NAND3X1_93 ( );
FILL FILL_6_NAND3X1_93 ( );
FILL FILL_7_NAND3X1_93 ( );
FILL FILL_8_NAND3X1_93 ( );
FILL FILL_0_NAND3X1_72 ( );
FILL FILL_1_NAND3X1_72 ( );
FILL FILL_2_NAND3X1_72 ( );
FILL FILL_3_NAND3X1_72 ( );
FILL FILL_4_NAND3X1_72 ( );
FILL FILL_5_NAND3X1_72 ( );
FILL FILL_6_NAND3X1_72 ( );
FILL FILL_7_NAND3X1_72 ( );
FILL FILL_8_NAND3X1_72 ( );
FILL FILL_0_NAND2X1_229 ( );
FILL FILL_1_NAND2X1_229 ( );
FILL FILL_2_NAND2X1_229 ( );
FILL FILL_3_NAND2X1_229 ( );
FILL FILL_4_NAND2X1_229 ( );
FILL FILL_5_NAND2X1_229 ( );
FILL FILL_6_NAND2X1_229 ( );
FILL FILL_0_OAI21X1_236 ( );
FILL FILL_1_OAI21X1_236 ( );
FILL FILL_2_OAI21X1_236 ( );
FILL FILL_3_OAI21X1_236 ( );
FILL FILL_4_OAI21X1_236 ( );
FILL FILL_5_OAI21X1_236 ( );
FILL FILL_6_OAI21X1_236 ( );
FILL FILL_7_OAI21X1_236 ( );
FILL FILL_8_OAI21X1_236 ( );
FILL FILL_0_BUFX2_21 ( );
FILL FILL_1_BUFX2_21 ( );
FILL FILL_2_BUFX2_21 ( );
FILL FILL_3_BUFX2_21 ( );
FILL FILL_4_BUFX2_21 ( );
FILL FILL_5_BUFX2_21 ( );
FILL FILL_6_BUFX2_21 ( );
FILL FILL_0_NAND2X1_127 ( );
FILL FILL_1_NAND2X1_127 ( );
FILL FILL_2_NAND2X1_127 ( );
FILL FILL_3_NAND2X1_127 ( );
FILL FILL_4_NAND2X1_127 ( );
FILL FILL_5_NAND2X1_127 ( );
FILL FILL_6_NAND2X1_127 ( );
FILL FILL_0_BUFX2_20 ( );
FILL FILL_1_BUFX2_20 ( );
FILL FILL_2_BUFX2_20 ( );
FILL FILL_3_BUFX2_20 ( );
FILL FILL_4_BUFX2_20 ( );
FILL FILL_5_BUFX2_20 ( );
FILL FILL_6_BUFX2_20 ( );
FILL FILL_0_INVX1_336 ( );
FILL FILL_1_INVX1_336 ( );
FILL FILL_2_INVX1_336 ( );
FILL FILL_3_INVX1_336 ( );
FILL FILL_0_OAI21X1_109 ( );
FILL FILL_1_OAI21X1_109 ( );
FILL FILL_2_OAI21X1_109 ( );
FILL FILL_3_OAI21X1_109 ( );
FILL FILL_4_OAI21X1_109 ( );
FILL FILL_5_OAI21X1_109 ( );
FILL FILL_6_OAI21X1_109 ( );
FILL FILL_7_OAI21X1_109 ( );
FILL FILL_8_OAI21X1_109 ( );
FILL FILL_0_INVX1_123 ( );
FILL FILL_1_INVX1_123 ( );
FILL FILL_2_INVX1_123 ( );
FILL FILL_3_INVX1_123 ( );
FILL FILL_4_INVX1_123 ( );
FILL FILL_0_OAI21X1_84 ( );
FILL FILL_1_OAI21X1_84 ( );
FILL FILL_2_OAI21X1_84 ( );
FILL FILL_3_OAI21X1_84 ( );
FILL FILL_4_OAI21X1_84 ( );
FILL FILL_5_OAI21X1_84 ( );
FILL FILL_6_OAI21X1_84 ( );
FILL FILL_7_OAI21X1_84 ( );
FILL FILL_8_OAI21X1_84 ( );
FILL FILL_9_OAI21X1_84 ( );
FILL FILL_0_INVX1_95 ( );
FILL FILL_1_INVX1_95 ( );
FILL FILL_2_INVX1_95 ( );
FILL FILL_3_INVX1_95 ( );
FILL FILL_0_INVX1_356 ( );
FILL FILL_1_INVX1_356 ( );
FILL FILL_2_INVX1_356 ( );
FILL FILL_3_INVX1_356 ( );
FILL FILL_4_INVX1_356 ( );
FILL FILL_0_CLKBUF1_8 ( );
FILL FILL_1_CLKBUF1_8 ( );
FILL FILL_2_CLKBUF1_8 ( );
FILL FILL_3_CLKBUF1_8 ( );
FILL FILL_4_CLKBUF1_8 ( );
FILL FILL_5_CLKBUF1_8 ( );
FILL FILL_6_CLKBUF1_8 ( );
FILL FILL_7_CLKBUF1_8 ( );
FILL FILL_8_CLKBUF1_8 ( );
FILL FILL_9_CLKBUF1_8 ( );
FILL FILL_10_CLKBUF1_8 ( );
FILL FILL_11_CLKBUF1_8 ( );
FILL FILL_12_CLKBUF1_8 ( );
FILL FILL_13_CLKBUF1_8 ( );
FILL FILL_14_CLKBUF1_8 ( );
FILL FILL_15_CLKBUF1_8 ( );
FILL FILL_16_CLKBUF1_8 ( );
FILL FILL_17_CLKBUF1_8 ( );
FILL FILL_18_CLKBUF1_8 ( );
FILL FILL_19_CLKBUF1_8 ( );
FILL FILL_20_CLKBUF1_8 ( );
FILL FILL_0_INVX1_352 ( );
FILL FILL_1_INVX1_352 ( );
FILL FILL_2_INVX1_352 ( );
FILL FILL_3_INVX1_352 ( );
FILL FILL_4_INVX1_352 ( );
FILL FILL_0_BUFX2_25 ( );
FILL FILL_1_BUFX2_25 ( );
FILL FILL_2_BUFX2_25 ( );
FILL FILL_3_BUFX2_25 ( );
FILL FILL_4_BUFX2_25 ( );
FILL FILL_5_BUFX2_25 ( );
FILL FILL_6_BUFX2_25 ( );
FILL FILL_0_NAND2X1_156 ( );
FILL FILL_1_NAND2X1_156 ( );
FILL FILL_2_NAND2X1_156 ( );
FILL FILL_3_NAND2X1_156 ( );
FILL FILL_4_NAND2X1_156 ( );
FILL FILL_5_NAND2X1_156 ( );
FILL FILL_6_NAND2X1_156 ( );
FILL FILL_0_INVX1_178 ( );
FILL FILL_1_INVX1_178 ( );
FILL FILL_2_INVX1_178 ( );
FILL FILL_3_INVX1_178 ( );
FILL FILL_4_INVX1_178 ( );
FILL FILL_0_OAI21X1_152 ( );
FILL FILL_1_OAI21X1_152 ( );
FILL FILL_2_OAI21X1_152 ( );
FILL FILL_3_OAI21X1_152 ( );
FILL FILL_4_OAI21X1_152 ( );
FILL FILL_5_OAI21X1_152 ( );
FILL FILL_6_OAI21X1_152 ( );
FILL FILL_7_OAI21X1_152 ( );
FILL FILL_8_OAI21X1_152 ( );
FILL FILL_0_NAND2X1_152 ( );
FILL FILL_1_NAND2X1_152 ( );
FILL FILL_2_NAND2X1_152 ( );
FILL FILL_3_NAND2X1_152 ( );
FILL FILL_4_NAND2X1_152 ( );
FILL FILL_5_NAND2X1_152 ( );
FILL FILL_6_NAND2X1_152 ( );
FILL FILL_0_NAND2X1_153 ( );
FILL FILL_1_NAND2X1_153 ( );
FILL FILL_2_NAND2X1_153 ( );
FILL FILL_3_NAND2X1_153 ( );
FILL FILL_4_NAND2X1_153 ( );
FILL FILL_5_NAND2X1_153 ( );
FILL FILL_6_NAND2X1_153 ( );
FILL FILL_0_OAI21X1_153 ( );
FILL FILL_1_OAI21X1_153 ( );
FILL FILL_2_OAI21X1_153 ( );
FILL FILL_3_OAI21X1_153 ( );
FILL FILL_4_OAI21X1_153 ( );
FILL FILL_5_OAI21X1_153 ( );
FILL FILL_6_OAI21X1_153 ( );
FILL FILL_7_OAI21X1_153 ( );
FILL FILL_8_OAI21X1_153 ( );
FILL FILL_0_DFFSR_6 ( );
FILL FILL_1_DFFSR_6 ( );
FILL FILL_2_DFFSR_6 ( );
FILL FILL_3_DFFSR_6 ( );
FILL FILL_4_DFFSR_6 ( );
FILL FILL_5_DFFSR_6 ( );
FILL FILL_6_DFFSR_6 ( );
FILL FILL_7_DFFSR_6 ( );
FILL FILL_8_DFFSR_6 ( );
FILL FILL_9_DFFSR_6 ( );
FILL FILL_10_DFFSR_6 ( );
FILL FILL_11_DFFSR_6 ( );
FILL FILL_12_DFFSR_6 ( );
FILL FILL_13_DFFSR_6 ( );
FILL FILL_14_DFFSR_6 ( );
FILL FILL_15_DFFSR_6 ( );
FILL FILL_16_DFFSR_6 ( );
FILL FILL_17_DFFSR_6 ( );
FILL FILL_18_DFFSR_6 ( );
FILL FILL_19_DFFSR_6 ( );
FILL FILL_20_DFFSR_6 ( );
FILL FILL_21_DFFSR_6 ( );
FILL FILL_22_DFFSR_6 ( );
FILL FILL_23_DFFSR_6 ( );
FILL FILL_24_DFFSR_6 ( );
FILL FILL_25_DFFSR_6 ( );
FILL FILL_26_DFFSR_6 ( );
FILL FILL_27_DFFSR_6 ( );
FILL FILL_28_DFFSR_6 ( );
FILL FILL_29_DFFSR_6 ( );
FILL FILL_30_DFFSR_6 ( );
FILL FILL_31_DFFSR_6 ( );
FILL FILL_32_DFFSR_6 ( );
FILL FILL_33_DFFSR_6 ( );
FILL FILL_34_DFFSR_6 ( );
FILL FILL_35_DFFSR_6 ( );
FILL FILL_36_DFFSR_6 ( );
FILL FILL_37_DFFSR_6 ( );
FILL FILL_38_DFFSR_6 ( );
FILL FILL_39_DFFSR_6 ( );
FILL FILL_40_DFFSR_6 ( );
FILL FILL_41_DFFSR_6 ( );
FILL FILL_42_DFFSR_6 ( );
FILL FILL_43_DFFSR_6 ( );
FILL FILL_44_DFFSR_6 ( );
FILL FILL_45_DFFSR_6 ( );
FILL FILL_46_DFFSR_6 ( );
FILL FILL_47_DFFSR_6 ( );
FILL FILL_48_DFFSR_6 ( );
FILL FILL_49_DFFSR_6 ( );
FILL FILL_50_DFFSR_6 ( );
FILL FILL_0_NAND2X1_8 ( );
FILL FILL_1_NAND2X1_8 ( );
FILL FILL_2_NAND2X1_8 ( );
FILL FILL_3_NAND2X1_8 ( );
FILL FILL_4_NAND2X1_8 ( );
FILL FILL_5_NAND2X1_8 ( );
FILL FILL_6_NAND2X1_8 ( );
FILL FILL_0_DFFSR_61 ( );
FILL FILL_1_DFFSR_61 ( );
FILL FILL_2_DFFSR_61 ( );
FILL FILL_3_DFFSR_61 ( );
FILL FILL_4_DFFSR_61 ( );
FILL FILL_5_DFFSR_61 ( );
FILL FILL_6_DFFSR_61 ( );
FILL FILL_7_DFFSR_61 ( );
FILL FILL_8_DFFSR_61 ( );
FILL FILL_9_DFFSR_61 ( );
FILL FILL_10_DFFSR_61 ( );
FILL FILL_11_DFFSR_61 ( );
FILL FILL_12_DFFSR_61 ( );
FILL FILL_13_DFFSR_61 ( );
FILL FILL_14_DFFSR_61 ( );
FILL FILL_15_DFFSR_61 ( );
FILL FILL_16_DFFSR_61 ( );
FILL FILL_17_DFFSR_61 ( );
FILL FILL_18_DFFSR_61 ( );
FILL FILL_19_DFFSR_61 ( );
FILL FILL_20_DFFSR_61 ( );
FILL FILL_21_DFFSR_61 ( );
FILL FILL_22_DFFSR_61 ( );
FILL FILL_23_DFFSR_61 ( );
FILL FILL_24_DFFSR_61 ( );
FILL FILL_25_DFFSR_61 ( );
FILL FILL_26_DFFSR_61 ( );
FILL FILL_27_DFFSR_61 ( );
FILL FILL_28_DFFSR_61 ( );
FILL FILL_29_DFFSR_61 ( );
FILL FILL_30_DFFSR_61 ( );
FILL FILL_31_DFFSR_61 ( );
FILL FILL_32_DFFSR_61 ( );
FILL FILL_33_DFFSR_61 ( );
FILL FILL_34_DFFSR_61 ( );
FILL FILL_35_DFFSR_61 ( );
FILL FILL_36_DFFSR_61 ( );
FILL FILL_37_DFFSR_61 ( );
FILL FILL_38_DFFSR_61 ( );
FILL FILL_39_DFFSR_61 ( );
FILL FILL_40_DFFSR_61 ( );
FILL FILL_41_DFFSR_61 ( );
FILL FILL_42_DFFSR_61 ( );
FILL FILL_43_DFFSR_61 ( );
FILL FILL_44_DFFSR_61 ( );
FILL FILL_45_DFFSR_61 ( );
FILL FILL_46_DFFSR_61 ( );
FILL FILL_47_DFFSR_61 ( );
FILL FILL_48_DFFSR_61 ( );
FILL FILL_49_DFFSR_61 ( );
FILL FILL_50_DFFSR_61 ( );
FILL FILL_0_NAND2X1_23 ( );
FILL FILL_1_NAND2X1_23 ( );
FILL FILL_2_NAND2X1_23 ( );
FILL FILL_3_NAND2X1_23 ( );
FILL FILL_4_NAND2X1_23 ( );
FILL FILL_5_NAND2X1_23 ( );
FILL FILL_6_NAND2X1_23 ( );
FILL FILL_0_DFFSR_169 ( );
FILL FILL_1_DFFSR_169 ( );
FILL FILL_2_DFFSR_169 ( );
FILL FILL_3_DFFSR_169 ( );
FILL FILL_4_DFFSR_169 ( );
FILL FILL_5_DFFSR_169 ( );
FILL FILL_6_DFFSR_169 ( );
FILL FILL_7_DFFSR_169 ( );
FILL FILL_8_DFFSR_169 ( );
FILL FILL_9_DFFSR_169 ( );
FILL FILL_10_DFFSR_169 ( );
FILL FILL_11_DFFSR_169 ( );
FILL FILL_12_DFFSR_169 ( );
FILL FILL_13_DFFSR_169 ( );
FILL FILL_14_DFFSR_169 ( );
FILL FILL_15_DFFSR_169 ( );
FILL FILL_16_DFFSR_169 ( );
FILL FILL_17_DFFSR_169 ( );
FILL FILL_18_DFFSR_169 ( );
FILL FILL_19_DFFSR_169 ( );
FILL FILL_20_DFFSR_169 ( );
FILL FILL_21_DFFSR_169 ( );
FILL FILL_22_DFFSR_169 ( );
FILL FILL_23_DFFSR_169 ( );
FILL FILL_24_DFFSR_169 ( );
FILL FILL_25_DFFSR_169 ( );
FILL FILL_26_DFFSR_169 ( );
FILL FILL_27_DFFSR_169 ( );
FILL FILL_28_DFFSR_169 ( );
FILL FILL_29_DFFSR_169 ( );
FILL FILL_30_DFFSR_169 ( );
FILL FILL_31_DFFSR_169 ( );
FILL FILL_32_DFFSR_169 ( );
FILL FILL_33_DFFSR_169 ( );
FILL FILL_34_DFFSR_169 ( );
FILL FILL_35_DFFSR_169 ( );
FILL FILL_36_DFFSR_169 ( );
FILL FILL_37_DFFSR_169 ( );
FILL FILL_38_DFFSR_169 ( );
FILL FILL_39_DFFSR_169 ( );
FILL FILL_40_DFFSR_169 ( );
FILL FILL_41_DFFSR_169 ( );
FILL FILL_42_DFFSR_169 ( );
FILL FILL_43_DFFSR_169 ( );
FILL FILL_44_DFFSR_169 ( );
FILL FILL_45_DFFSR_169 ( );
FILL FILL_46_DFFSR_169 ( );
FILL FILL_47_DFFSR_169 ( );
FILL FILL_48_DFFSR_169 ( );
FILL FILL_49_DFFSR_169 ( );
FILL FILL_50_DFFSR_169 ( );
FILL FILL_0_NAND3X1_38 ( );
FILL FILL_1_NAND3X1_38 ( );
FILL FILL_2_NAND3X1_38 ( );
FILL FILL_3_NAND3X1_38 ( );
FILL FILL_4_NAND3X1_38 ( );
FILL FILL_5_NAND3X1_38 ( );
FILL FILL_6_NAND3X1_38 ( );
FILL FILL_7_NAND3X1_38 ( );
FILL FILL_8_NAND3X1_38 ( );
FILL FILL_0_NAND2X1_204 ( );
FILL FILL_1_NAND2X1_204 ( );
FILL FILL_2_NAND2X1_204 ( );
FILL FILL_3_NAND2X1_204 ( );
FILL FILL_4_NAND2X1_204 ( );
FILL FILL_5_NAND2X1_204 ( );
FILL FILL_6_NAND2X1_204 ( );
FILL FILL_0_AND2X2_6 ( );
FILL FILL_1_AND2X2_6 ( );
FILL FILL_2_AND2X2_6 ( );
FILL FILL_3_AND2X2_6 ( );
FILL FILL_4_AND2X2_6 ( );
FILL FILL_5_AND2X2_6 ( );
FILL FILL_6_AND2X2_6 ( );
FILL FILL_7_AND2X2_6 ( );
FILL FILL_8_AND2X2_6 ( );
FILL FILL_0_INVX1_227 ( );
FILL FILL_1_INVX1_227 ( );
FILL FILL_2_INVX1_227 ( );
FILL FILL_3_INVX1_227 ( );
FILL FILL_4_INVX1_227 ( );
FILL FILL_0_AOI22X1_5 ( );
FILL FILL_1_AOI22X1_5 ( );
FILL FILL_2_AOI22X1_5 ( );
FILL FILL_3_AOI22X1_5 ( );
FILL FILL_4_AOI22X1_5 ( );
FILL FILL_5_AOI22X1_5 ( );
FILL FILL_6_AOI22X1_5 ( );
FILL FILL_7_AOI22X1_5 ( );
FILL FILL_8_AOI22X1_5 ( );
FILL FILL_9_AOI22X1_5 ( );
FILL FILL_10_AOI22X1_5 ( );
FILL FILL_11_AOI22X1_5 ( );
FILL FILL_0_NAND2X1_192 ( );
FILL FILL_1_NAND2X1_192 ( );
FILL FILL_2_NAND2X1_192 ( );
FILL FILL_3_NAND2X1_192 ( );
FILL FILL_4_NAND2X1_192 ( );
FILL FILL_5_NAND2X1_192 ( );
FILL FILL_6_NAND2X1_192 ( );
FILL FILL_0_NAND2X1_189 ( );
FILL FILL_1_NAND2X1_189 ( );
FILL FILL_2_NAND2X1_189 ( );
FILL FILL_3_NAND2X1_189 ( );
FILL FILL_4_NAND2X1_189 ( );
FILL FILL_5_NAND2X1_189 ( );
FILL FILL_6_NAND2X1_189 ( );
FILL FILL_0_INVX1_214 ( );
FILL FILL_1_INVX1_214 ( );
FILL FILL_2_INVX1_214 ( );
FILL FILL_3_INVX1_214 ( );
FILL FILL_0_NAND2X1_216 ( );
FILL FILL_1_NAND2X1_216 ( );
FILL FILL_2_NAND2X1_216 ( );
FILL FILL_3_NAND2X1_216 ( );
FILL FILL_4_NAND2X1_216 ( );
FILL FILL_5_NAND2X1_216 ( );
FILL FILL_6_NAND2X1_216 ( );
FILL FILL_0_OAI21X1_190 ( );
FILL FILL_1_OAI21X1_190 ( );
FILL FILL_2_OAI21X1_190 ( );
FILL FILL_3_OAI21X1_190 ( );
FILL FILL_4_OAI21X1_190 ( );
FILL FILL_5_OAI21X1_190 ( );
FILL FILL_6_OAI21X1_190 ( );
FILL FILL_7_OAI21X1_190 ( );
FILL FILL_8_OAI21X1_190 ( );
FILL FILL_9_OAI21X1_190 ( );
FILL FILL_0_AOI21X1_23 ( );
FILL FILL_1_AOI21X1_23 ( );
FILL FILL_2_AOI21X1_23 ( );
FILL FILL_3_AOI21X1_23 ( );
FILL FILL_4_AOI21X1_23 ( );
FILL FILL_5_AOI21X1_23 ( );
FILL FILL_6_AOI21X1_23 ( );
FILL FILL_7_AOI21X1_23 ( );
FILL FILL_8_AOI21X1_23 ( );
FILL FILL_9_AOI21X1_23 ( );
FILL FILL_0_OAI21X1_208 ( );
FILL FILL_1_OAI21X1_208 ( );
FILL FILL_2_OAI21X1_208 ( );
FILL FILL_3_OAI21X1_208 ( );
FILL FILL_4_OAI21X1_208 ( );
FILL FILL_5_OAI21X1_208 ( );
FILL FILL_6_OAI21X1_208 ( );
FILL FILL_7_OAI21X1_208 ( );
FILL FILL_8_OAI21X1_208 ( );
FILL FILL_0_AOI21X1_27 ( );
FILL FILL_1_AOI21X1_27 ( );
FILL FILL_2_AOI21X1_27 ( );
FILL FILL_3_AOI21X1_27 ( );
FILL FILL_4_AOI21X1_27 ( );
FILL FILL_5_AOI21X1_27 ( );
FILL FILL_6_AOI21X1_27 ( );
FILL FILL_7_AOI21X1_27 ( );
FILL FILL_8_AOI21X1_27 ( );
FILL FILL_9_AOI21X1_27 ( );
FILL FILL_0_NAND3X1_76 ( );
FILL FILL_1_NAND3X1_76 ( );
FILL FILL_2_NAND3X1_76 ( );
FILL FILL_3_NAND3X1_76 ( );
FILL FILL_4_NAND3X1_76 ( );
FILL FILL_5_NAND3X1_76 ( );
FILL FILL_6_NAND3X1_76 ( );
FILL FILL_7_NAND3X1_76 ( );
FILL FILL_8_NAND3X1_76 ( );
FILL FILL_9_NAND3X1_76 ( );
FILL FILL_0_XOR2X1_8 ( );
FILL FILL_1_XOR2X1_8 ( );
FILL FILL_2_XOR2X1_8 ( );
FILL FILL_3_XOR2X1_8 ( );
FILL FILL_4_XOR2X1_8 ( );
FILL FILL_5_XOR2X1_8 ( );
FILL FILL_6_XOR2X1_8 ( );
FILL FILL_7_XOR2X1_8 ( );
FILL FILL_8_XOR2X1_8 ( );
FILL FILL_9_XOR2X1_8 ( );
FILL FILL_10_XOR2X1_8 ( );
FILL FILL_11_XOR2X1_8 ( );
FILL FILL_12_XOR2X1_8 ( );
FILL FILL_13_XOR2X1_8 ( );
FILL FILL_14_XOR2X1_8 ( );
FILL FILL_15_XOR2X1_8 ( );
FILL FILL_16_XOR2X1_8 ( );
FILL FILL_0_NAND3X1_106 ( );
FILL FILL_1_NAND3X1_106 ( );
FILL FILL_2_NAND3X1_106 ( );
FILL FILL_3_NAND3X1_106 ( );
FILL FILL_4_NAND3X1_106 ( );
FILL FILL_5_NAND3X1_106 ( );
FILL FILL_6_NAND3X1_106 ( );
FILL FILL_7_NAND3X1_106 ( );
FILL FILL_8_NAND3X1_106 ( );
FILL FILL_9_NAND3X1_106 ( );
FILL FILL_0_DFFSR_121 ( );
FILL FILL_1_DFFSR_121 ( );
FILL FILL_2_DFFSR_121 ( );
FILL FILL_3_DFFSR_121 ( );
FILL FILL_4_DFFSR_121 ( );
FILL FILL_5_DFFSR_121 ( );
FILL FILL_6_DFFSR_121 ( );
FILL FILL_7_DFFSR_121 ( );
FILL FILL_8_DFFSR_121 ( );
FILL FILL_9_DFFSR_121 ( );
FILL FILL_10_DFFSR_121 ( );
FILL FILL_11_DFFSR_121 ( );
FILL FILL_12_DFFSR_121 ( );
FILL FILL_13_DFFSR_121 ( );
FILL FILL_14_DFFSR_121 ( );
FILL FILL_15_DFFSR_121 ( );
FILL FILL_16_DFFSR_121 ( );
FILL FILL_17_DFFSR_121 ( );
FILL FILL_18_DFFSR_121 ( );
FILL FILL_19_DFFSR_121 ( );
FILL FILL_20_DFFSR_121 ( );
FILL FILL_21_DFFSR_121 ( );
FILL FILL_22_DFFSR_121 ( );
FILL FILL_23_DFFSR_121 ( );
FILL FILL_24_DFFSR_121 ( );
FILL FILL_25_DFFSR_121 ( );
FILL FILL_26_DFFSR_121 ( );
FILL FILL_27_DFFSR_121 ( );
FILL FILL_28_DFFSR_121 ( );
FILL FILL_29_DFFSR_121 ( );
FILL FILL_30_DFFSR_121 ( );
FILL FILL_31_DFFSR_121 ( );
FILL FILL_32_DFFSR_121 ( );
FILL FILL_33_DFFSR_121 ( );
FILL FILL_34_DFFSR_121 ( );
FILL FILL_35_DFFSR_121 ( );
FILL FILL_36_DFFSR_121 ( );
FILL FILL_37_DFFSR_121 ( );
FILL FILL_38_DFFSR_121 ( );
FILL FILL_39_DFFSR_121 ( );
FILL FILL_40_DFFSR_121 ( );
FILL FILL_41_DFFSR_121 ( );
FILL FILL_42_DFFSR_121 ( );
FILL FILL_43_DFFSR_121 ( );
FILL FILL_44_DFFSR_121 ( );
FILL FILL_45_DFFSR_121 ( );
FILL FILL_46_DFFSR_121 ( );
FILL FILL_47_DFFSR_121 ( );
FILL FILL_48_DFFSR_121 ( );
FILL FILL_49_DFFSR_121 ( );
FILL FILL_50_DFFSR_121 ( );
FILL FILL_0_NAND2X1_84 ( );
FILL FILL_1_NAND2X1_84 ( );
FILL FILL_2_NAND2X1_84 ( );
FILL FILL_3_NAND2X1_84 ( );
FILL FILL_4_NAND2X1_84 ( );
FILL FILL_5_NAND2X1_84 ( );
FILL FILL_6_NAND2X1_84 ( );
FILL FILL_0_INVX1_121 ( );
FILL FILL_1_INVX1_121 ( );
FILL FILL_2_INVX1_121 ( );
FILL FILL_3_INVX1_121 ( );
FILL FILL_4_INVX1_121 ( );
FILL FILL_0_OAI21X1_107 ( );
FILL FILL_1_OAI21X1_107 ( );
FILL FILL_2_OAI21X1_107 ( );
FILL FILL_3_OAI21X1_107 ( );
FILL FILL_4_OAI21X1_107 ( );
FILL FILL_5_OAI21X1_107 ( );
FILL FILL_6_OAI21X1_107 ( );
FILL FILL_7_OAI21X1_107 ( );
FILL FILL_8_OAI21X1_107 ( );
FILL FILL_0_NAND2X1_107 ( );
FILL FILL_1_NAND2X1_107 ( );
FILL FILL_2_NAND2X1_107 ( );
FILL FILL_3_NAND2X1_107 ( );
FILL FILL_4_NAND2X1_107 ( );
FILL FILL_5_NAND2X1_107 ( );
FILL FILL_6_NAND2X1_107 ( );
FILL FILL_0_NAND2X1_115 ( );
FILL FILL_1_NAND2X1_115 ( );
FILL FILL_2_NAND2X1_115 ( );
FILL FILL_3_NAND2X1_115 ( );
FILL FILL_4_NAND2X1_115 ( );
FILL FILL_5_NAND2X1_115 ( );
FILL FILL_6_NAND2X1_115 ( );
FILL FILL_0_INVX1_130 ( );
FILL FILL_1_INVX1_130 ( );
FILL FILL_2_INVX1_130 ( );
FILL FILL_3_INVX1_130 ( );
FILL FILL_4_INVX1_130 ( );
FILL FILL_0_OAI21X1_115 ( );
FILL FILL_1_OAI21X1_115 ( );
FILL FILL_2_OAI21X1_115 ( );
FILL FILL_3_OAI21X1_115 ( );
FILL FILL_4_OAI21X1_115 ( );
FILL FILL_5_OAI21X1_115 ( );
FILL FILL_6_OAI21X1_115 ( );
FILL FILL_7_OAI21X1_115 ( );
FILL FILL_8_OAI21X1_115 ( );
FILL FILL_0_DFFSR_154 ( );
FILL FILL_1_DFFSR_154 ( );
FILL FILL_2_DFFSR_154 ( );
FILL FILL_3_DFFSR_154 ( );
FILL FILL_4_DFFSR_154 ( );
FILL FILL_5_DFFSR_154 ( );
FILL FILL_6_DFFSR_154 ( );
FILL FILL_7_DFFSR_154 ( );
FILL FILL_8_DFFSR_154 ( );
FILL FILL_9_DFFSR_154 ( );
FILL FILL_10_DFFSR_154 ( );
FILL FILL_11_DFFSR_154 ( );
FILL FILL_12_DFFSR_154 ( );
FILL FILL_13_DFFSR_154 ( );
FILL FILL_14_DFFSR_154 ( );
FILL FILL_15_DFFSR_154 ( );
FILL FILL_16_DFFSR_154 ( );
FILL FILL_17_DFFSR_154 ( );
FILL FILL_18_DFFSR_154 ( );
FILL FILL_19_DFFSR_154 ( );
FILL FILL_20_DFFSR_154 ( );
FILL FILL_21_DFFSR_154 ( );
FILL FILL_22_DFFSR_154 ( );
FILL FILL_23_DFFSR_154 ( );
FILL FILL_24_DFFSR_154 ( );
FILL FILL_25_DFFSR_154 ( );
FILL FILL_26_DFFSR_154 ( );
FILL FILL_27_DFFSR_154 ( );
FILL FILL_28_DFFSR_154 ( );
FILL FILL_29_DFFSR_154 ( );
FILL FILL_30_DFFSR_154 ( );
FILL FILL_31_DFFSR_154 ( );
FILL FILL_32_DFFSR_154 ( );
FILL FILL_33_DFFSR_154 ( );
FILL FILL_34_DFFSR_154 ( );
FILL FILL_35_DFFSR_154 ( );
FILL FILL_36_DFFSR_154 ( );
FILL FILL_37_DFFSR_154 ( );
FILL FILL_38_DFFSR_154 ( );
FILL FILL_39_DFFSR_154 ( );
FILL FILL_40_DFFSR_154 ( );
FILL FILL_41_DFFSR_154 ( );
FILL FILL_42_DFFSR_154 ( );
FILL FILL_43_DFFSR_154 ( );
FILL FILL_44_DFFSR_154 ( );
FILL FILL_45_DFFSR_154 ( );
FILL FILL_46_DFFSR_154 ( );
FILL FILL_47_DFFSR_154 ( );
FILL FILL_48_DFFSR_154 ( );
FILL FILL_49_DFFSR_154 ( );
FILL FILL_50_DFFSR_154 ( );
FILL FILL_0_NAND2X1_135 ( );
FILL FILL_1_NAND2X1_135 ( );
FILL FILL_2_NAND2X1_135 ( );
FILL FILL_3_NAND2X1_135 ( );
FILL FILL_4_NAND2X1_135 ( );
FILL FILL_5_NAND2X1_135 ( );
FILL FILL_6_NAND2X1_135 ( );
FILL FILL_0_OAI21X1_6 ( );
FILL FILL_1_OAI21X1_6 ( );
FILL FILL_2_OAI21X1_6 ( );
FILL FILL_3_OAI21X1_6 ( );
FILL FILL_4_OAI21X1_6 ( );
FILL FILL_5_OAI21X1_6 ( );
FILL FILL_6_OAI21X1_6 ( );
FILL FILL_7_OAI21X1_6 ( );
FILL FILL_8_OAI21X1_6 ( );
FILL FILL_0_NOR2X1_1 ( );
FILL FILL_1_NOR2X1_1 ( );
FILL FILL_2_NOR2X1_1 ( );
FILL FILL_3_NOR2X1_1 ( );
FILL FILL_4_NOR2X1_1 ( );
FILL FILL_5_NOR2X1_1 ( );
FILL FILL_6_NOR2X1_1 ( );
FILL FILL_0_INVX1_9 ( );
FILL FILL_1_INVX1_9 ( );
FILL FILL_2_INVX1_9 ( );
FILL FILL_3_INVX1_9 ( );
FILL FILL_0_OAI21X1_8 ( );
FILL FILL_1_OAI21X1_8 ( );
FILL FILL_2_OAI21X1_8 ( );
FILL FILL_3_OAI21X1_8 ( );
FILL FILL_4_OAI21X1_8 ( );
FILL FILL_5_OAI21X1_8 ( );
FILL FILL_6_OAI21X1_8 ( );
FILL FILL_7_OAI21X1_8 ( );
FILL FILL_8_OAI21X1_8 ( );
FILL FILL_9_OAI21X1_8 ( );
FILL FILL_0_INVX1_312 ( );
FILL FILL_1_INVX1_312 ( );
FILL FILL_2_INVX1_312 ( );
FILL FILL_3_INVX1_312 ( );
FILL FILL_4_INVX1_312 ( );
FILL FILL_0_DFFSR_46 ( );
FILL FILL_1_DFFSR_46 ( );
FILL FILL_2_DFFSR_46 ( );
FILL FILL_3_DFFSR_46 ( );
FILL FILL_4_DFFSR_46 ( );
FILL FILL_5_DFFSR_46 ( );
FILL FILL_6_DFFSR_46 ( );
FILL FILL_7_DFFSR_46 ( );
FILL FILL_8_DFFSR_46 ( );
FILL FILL_9_DFFSR_46 ( );
FILL FILL_10_DFFSR_46 ( );
FILL FILL_11_DFFSR_46 ( );
FILL FILL_12_DFFSR_46 ( );
FILL FILL_13_DFFSR_46 ( );
FILL FILL_14_DFFSR_46 ( );
FILL FILL_15_DFFSR_46 ( );
FILL FILL_16_DFFSR_46 ( );
FILL FILL_17_DFFSR_46 ( );
FILL FILL_18_DFFSR_46 ( );
FILL FILL_19_DFFSR_46 ( );
FILL FILL_20_DFFSR_46 ( );
FILL FILL_21_DFFSR_46 ( );
FILL FILL_22_DFFSR_46 ( );
FILL FILL_23_DFFSR_46 ( );
FILL FILL_24_DFFSR_46 ( );
FILL FILL_25_DFFSR_46 ( );
FILL FILL_26_DFFSR_46 ( );
FILL FILL_27_DFFSR_46 ( );
FILL FILL_28_DFFSR_46 ( );
FILL FILL_29_DFFSR_46 ( );
FILL FILL_30_DFFSR_46 ( );
FILL FILL_31_DFFSR_46 ( );
FILL FILL_32_DFFSR_46 ( );
FILL FILL_33_DFFSR_46 ( );
FILL FILL_34_DFFSR_46 ( );
FILL FILL_35_DFFSR_46 ( );
FILL FILL_36_DFFSR_46 ( );
FILL FILL_37_DFFSR_46 ( );
FILL FILL_38_DFFSR_46 ( );
FILL FILL_39_DFFSR_46 ( );
FILL FILL_40_DFFSR_46 ( );
FILL FILL_41_DFFSR_46 ( );
FILL FILL_42_DFFSR_46 ( );
FILL FILL_43_DFFSR_46 ( );
FILL FILL_44_DFFSR_46 ( );
FILL FILL_45_DFFSR_46 ( );
FILL FILL_46_DFFSR_46 ( );
FILL FILL_47_DFFSR_46 ( );
FILL FILL_48_DFFSR_46 ( );
FILL FILL_49_DFFSR_46 ( );
FILL FILL_50_DFFSR_46 ( );
FILL FILL_0_NAND2X1_168 ( );
FILL FILL_1_NAND2X1_168 ( );
FILL FILL_2_NAND2X1_168 ( );
FILL FILL_3_NAND2X1_168 ( );
FILL FILL_4_NAND2X1_168 ( );
FILL FILL_5_NAND2X1_168 ( );
FILL FILL_6_NAND2X1_168 ( );
FILL FILL_0_OAI21X1_168 ( );
FILL FILL_1_OAI21X1_168 ( );
FILL FILL_2_OAI21X1_168 ( );
FILL FILL_3_OAI21X1_168 ( );
FILL FILL_4_OAI21X1_168 ( );
FILL FILL_5_OAI21X1_168 ( );
FILL FILL_6_OAI21X1_168 ( );
FILL FILL_7_OAI21X1_168 ( );
FILL FILL_8_OAI21X1_168 ( );
FILL FILL_9_OAI21X1_168 ( );
FILL FILL_0_INVX1_203 ( );
FILL FILL_1_INVX1_203 ( );
FILL FILL_2_INVX1_203 ( );
FILL FILL_3_INVX1_203 ( );
FILL FILL_0_CLKBUF1_16 ( );
FILL FILL_1_CLKBUF1_16 ( );
FILL FILL_2_CLKBUF1_16 ( );
FILL FILL_3_CLKBUF1_16 ( );
FILL FILL_4_CLKBUF1_16 ( );
FILL FILL_5_CLKBUF1_16 ( );
FILL FILL_6_CLKBUF1_16 ( );
FILL FILL_7_CLKBUF1_16 ( );
FILL FILL_8_CLKBUF1_16 ( );
FILL FILL_9_CLKBUF1_16 ( );
FILL FILL_10_CLKBUF1_16 ( );
FILL FILL_11_CLKBUF1_16 ( );
FILL FILL_12_CLKBUF1_16 ( );
FILL FILL_13_CLKBUF1_16 ( );
FILL FILL_14_CLKBUF1_16 ( );
FILL FILL_15_CLKBUF1_16 ( );
FILL FILL_16_CLKBUF1_16 ( );
FILL FILL_17_CLKBUF1_16 ( );
FILL FILL_18_CLKBUF1_16 ( );
FILL FILL_19_CLKBUF1_16 ( );
FILL FILL_20_CLKBUF1_16 ( );
FILL FILL_0_NAND2X1_172 ( );
FILL FILL_1_NAND2X1_172 ( );
FILL FILL_2_NAND2X1_172 ( );
FILL FILL_3_NAND2X1_172 ( );
FILL FILL_4_NAND2X1_172 ( );
FILL FILL_5_NAND2X1_172 ( );
FILL FILL_6_NAND2X1_172 ( );
FILL FILL_0_OAI21X1_172 ( );
FILL FILL_1_OAI21X1_172 ( );
FILL FILL_2_OAI21X1_172 ( );
FILL FILL_3_OAI21X1_172 ( );
FILL FILL_4_OAI21X1_172 ( );
FILL FILL_5_OAI21X1_172 ( );
FILL FILL_6_OAI21X1_172 ( );
FILL FILL_7_OAI21X1_172 ( );
FILL FILL_8_OAI21X1_172 ( );
FILL FILL_9_OAI21X1_172 ( );
FILL FILL_0_INVX1_207 ( );
FILL FILL_1_INVX1_207 ( );
FILL FILL_2_INVX1_207 ( );
FILL FILL_3_INVX1_207 ( );
FILL FILL_0_NAND2X1_205 ( );
FILL FILL_1_NAND2X1_205 ( );
FILL FILL_2_NAND2X1_205 ( );
FILL FILL_3_NAND2X1_205 ( );
FILL FILL_4_NAND2X1_205 ( );
FILL FILL_5_NAND2X1_205 ( );
FILL FILL_6_NAND2X1_205 ( );
FILL FILL_0_INVX1_242 ( );
FILL FILL_1_INVX1_242 ( );
FILL FILL_2_INVX1_242 ( );
FILL FILL_3_INVX1_242 ( );
FILL FILL_0_OAI21X1_204 ( );
FILL FILL_1_OAI21X1_204 ( );
FILL FILL_2_OAI21X1_204 ( );
FILL FILL_3_OAI21X1_204 ( );
FILL FILL_4_OAI21X1_204 ( );
FILL FILL_5_OAI21X1_204 ( );
FILL FILL_6_OAI21X1_204 ( );
FILL FILL_7_OAI21X1_204 ( );
FILL FILL_8_OAI21X1_204 ( );
FILL FILL_9_OAI21X1_204 ( );
FILL FILL_0_INVX1_216 ( );
FILL FILL_1_INVX1_216 ( );
FILL FILL_2_INVX1_216 ( );
FILL FILL_3_INVX1_216 ( );
FILL FILL_4_INVX1_216 ( );
FILL FILL_0_INVX1_193 ( );
FILL FILL_1_INVX1_193 ( );
FILL FILL_2_INVX1_193 ( );
FILL FILL_3_INVX1_193 ( );
FILL FILL_4_INVX1_193 ( );
FILL FILL_0_DFFSR_159 ( );
FILL FILL_1_DFFSR_159 ( );
FILL FILL_2_DFFSR_159 ( );
FILL FILL_3_DFFSR_159 ( );
FILL FILL_4_DFFSR_159 ( );
FILL FILL_5_DFFSR_159 ( );
FILL FILL_6_DFFSR_159 ( );
FILL FILL_7_DFFSR_159 ( );
FILL FILL_8_DFFSR_159 ( );
FILL FILL_9_DFFSR_159 ( );
FILL FILL_10_DFFSR_159 ( );
FILL FILL_11_DFFSR_159 ( );
FILL FILL_12_DFFSR_159 ( );
FILL FILL_13_DFFSR_159 ( );
FILL FILL_14_DFFSR_159 ( );
FILL FILL_15_DFFSR_159 ( );
FILL FILL_16_DFFSR_159 ( );
FILL FILL_17_DFFSR_159 ( );
FILL FILL_18_DFFSR_159 ( );
FILL FILL_19_DFFSR_159 ( );
FILL FILL_20_DFFSR_159 ( );
FILL FILL_21_DFFSR_159 ( );
FILL FILL_22_DFFSR_159 ( );
FILL FILL_23_DFFSR_159 ( );
FILL FILL_24_DFFSR_159 ( );
FILL FILL_25_DFFSR_159 ( );
FILL FILL_26_DFFSR_159 ( );
FILL FILL_27_DFFSR_159 ( );
FILL FILL_28_DFFSR_159 ( );
FILL FILL_29_DFFSR_159 ( );
FILL FILL_30_DFFSR_159 ( );
FILL FILL_31_DFFSR_159 ( );
FILL FILL_32_DFFSR_159 ( );
FILL FILL_33_DFFSR_159 ( );
FILL FILL_34_DFFSR_159 ( );
FILL FILL_35_DFFSR_159 ( );
FILL FILL_36_DFFSR_159 ( );
FILL FILL_37_DFFSR_159 ( );
FILL FILL_38_DFFSR_159 ( );
FILL FILL_39_DFFSR_159 ( );
FILL FILL_40_DFFSR_159 ( );
FILL FILL_41_DFFSR_159 ( );
FILL FILL_42_DFFSR_159 ( );
FILL FILL_43_DFFSR_159 ( );
FILL FILL_44_DFFSR_159 ( );
FILL FILL_45_DFFSR_159 ( );
FILL FILL_46_DFFSR_159 ( );
FILL FILL_47_DFFSR_159 ( );
FILL FILL_48_DFFSR_159 ( );
FILL FILL_49_DFFSR_159 ( );
FILL FILL_50_DFFSR_159 ( );
FILL FILL_0_OAI21X1_213 ( );
FILL FILL_1_OAI21X1_213 ( );
FILL FILL_2_OAI21X1_213 ( );
FILL FILL_3_OAI21X1_213 ( );
FILL FILL_4_OAI21X1_213 ( );
FILL FILL_5_OAI21X1_213 ( );
FILL FILL_6_OAI21X1_213 ( );
FILL FILL_7_OAI21X1_213 ( );
FILL FILL_8_OAI21X1_213 ( );
FILL FILL_0_OAI21X1_231 ( );
FILL FILL_1_OAI21X1_231 ( );
FILL FILL_2_OAI21X1_231 ( );
FILL FILL_3_OAI21X1_231 ( );
FILL FILL_4_OAI21X1_231 ( );
FILL FILL_5_OAI21X1_231 ( );
FILL FILL_6_OAI21X1_231 ( );
FILL FILL_7_OAI21X1_231 ( );
FILL FILL_8_OAI21X1_231 ( );
FILL FILL_0_NAND2X1_226 ( );
FILL FILL_1_NAND2X1_226 ( );
FILL FILL_2_NAND2X1_226 ( );
FILL FILL_3_NAND2X1_226 ( );
FILL FILL_4_NAND2X1_226 ( );
FILL FILL_5_NAND2X1_226 ( );
FILL FILL_6_NAND2X1_226 ( );
FILL FILL_0_NOR2X1_10 ( );
FILL FILL_1_NOR2X1_10 ( );
FILL FILL_2_NOR2X1_10 ( );
FILL FILL_3_NOR2X1_10 ( );
FILL FILL_4_NOR2X1_10 ( );
FILL FILL_5_NOR2X1_10 ( );
FILL FILL_6_NOR2X1_10 ( );
FILL FILL_0_INVX1_252 ( );
FILL FILL_1_INVX1_252 ( );
FILL FILL_2_INVX1_252 ( );
FILL FILL_3_INVX1_252 ( );
FILL FILL_4_INVX1_252 ( );
FILL FILL_0_NAND3X1_79 ( );
FILL FILL_1_NAND3X1_79 ( );
FILL FILL_2_NAND3X1_79 ( );
FILL FILL_3_NAND3X1_79 ( );
FILL FILL_4_NAND3X1_79 ( );
FILL FILL_5_NAND3X1_79 ( );
FILL FILL_6_NAND3X1_79 ( );
FILL FILL_7_NAND3X1_79 ( );
FILL FILL_8_NAND3X1_79 ( );
FILL FILL_9_NAND3X1_79 ( );
FILL FILL_0_NAND2X1_230 ( );
FILL FILL_1_NAND2X1_230 ( );
FILL FILL_2_NAND2X1_230 ( );
FILL FILL_3_NAND2X1_230 ( );
FILL FILL_4_NAND2X1_230 ( );
FILL FILL_5_NAND2X1_230 ( );
FILL FILL_6_NAND2X1_230 ( );
FILL FILL_0_INVX1_339 ( );
FILL FILL_1_INVX1_339 ( );
FILL FILL_2_INVX1_339 ( );
FILL FILL_3_INVX1_339 ( );
FILL FILL_4_INVX1_339 ( );
FILL FILL_0_NAND2X1_121 ( );
FILL FILL_1_NAND2X1_121 ( );
FILL FILL_2_NAND2X1_121 ( );
FILL FILL_3_NAND2X1_121 ( );
FILL FILL_4_NAND2X1_121 ( );
FILL FILL_5_NAND2X1_121 ( );
FILL FILL_6_NAND2X1_121 ( );
FILL FILL_0_OAI21X1_121 ( );
FILL FILL_1_OAI21X1_121 ( );
FILL FILL_2_OAI21X1_121 ( );
FILL FILL_3_OAI21X1_121 ( );
FILL FILL_4_OAI21X1_121 ( );
FILL FILL_5_OAI21X1_121 ( );
FILL FILL_6_OAI21X1_121 ( );
FILL FILL_7_OAI21X1_121 ( );
FILL FILL_8_OAI21X1_121 ( );
FILL FILL_0_INVX1_137 ( );
FILL FILL_1_INVX1_137 ( );
FILL FILL_2_INVX1_137 ( );
FILL FILL_3_INVX1_137 ( );
FILL FILL_4_INVX1_137 ( );
FILL FILL_0_INVX1_337 ( );
FILL FILL_1_INVX1_337 ( );
FILL FILL_2_INVX1_337 ( );
FILL FILL_3_INVX1_337 ( );
FILL FILL_4_INVX1_337 ( );
FILL FILL_0_INVX1_338 ( );
FILL FILL_1_INVX1_338 ( );
FILL FILL_2_INVX1_338 ( );
FILL FILL_3_INVX1_338 ( );
FILL FILL_4_INVX1_338 ( );
FILL FILL_0_INVX1_370 ( );
FILL FILL_1_INVX1_370 ( );
FILL FILL_2_INVX1_370 ( );
FILL FILL_3_INVX1_370 ( );
FILL FILL_4_INVX1_370 ( );
FILL FILL_0_DFFSR_107 ( );
FILL FILL_1_DFFSR_107 ( );
FILL FILL_2_DFFSR_107 ( );
FILL FILL_3_DFFSR_107 ( );
FILL FILL_4_DFFSR_107 ( );
FILL FILL_5_DFFSR_107 ( );
FILL FILL_6_DFFSR_107 ( );
FILL FILL_7_DFFSR_107 ( );
FILL FILL_8_DFFSR_107 ( );
FILL FILL_9_DFFSR_107 ( );
FILL FILL_10_DFFSR_107 ( );
FILL FILL_11_DFFSR_107 ( );
FILL FILL_12_DFFSR_107 ( );
FILL FILL_13_DFFSR_107 ( );
FILL FILL_14_DFFSR_107 ( );
FILL FILL_15_DFFSR_107 ( );
FILL FILL_16_DFFSR_107 ( );
FILL FILL_17_DFFSR_107 ( );
FILL FILL_18_DFFSR_107 ( );
FILL FILL_19_DFFSR_107 ( );
FILL FILL_20_DFFSR_107 ( );
FILL FILL_21_DFFSR_107 ( );
FILL FILL_22_DFFSR_107 ( );
FILL FILL_23_DFFSR_107 ( );
FILL FILL_24_DFFSR_107 ( );
FILL FILL_25_DFFSR_107 ( );
FILL FILL_26_DFFSR_107 ( );
FILL FILL_27_DFFSR_107 ( );
FILL FILL_28_DFFSR_107 ( );
FILL FILL_29_DFFSR_107 ( );
FILL FILL_30_DFFSR_107 ( );
FILL FILL_31_DFFSR_107 ( );
FILL FILL_32_DFFSR_107 ( );
FILL FILL_33_DFFSR_107 ( );
FILL FILL_34_DFFSR_107 ( );
FILL FILL_35_DFFSR_107 ( );
FILL FILL_36_DFFSR_107 ( );
FILL FILL_37_DFFSR_107 ( );
FILL FILL_38_DFFSR_107 ( );
FILL FILL_39_DFFSR_107 ( );
FILL FILL_40_DFFSR_107 ( );
FILL FILL_41_DFFSR_107 ( );
FILL FILL_42_DFFSR_107 ( );
FILL FILL_43_DFFSR_107 ( );
FILL FILL_44_DFFSR_107 ( );
FILL FILL_45_DFFSR_107 ( );
FILL FILL_46_DFFSR_107 ( );
FILL FILL_47_DFFSR_107 ( );
FILL FILL_48_DFFSR_107 ( );
FILL FILL_49_DFFSR_107 ( );
FILL FILL_50_DFFSR_107 ( );
FILL FILL_51_DFFSR_107 ( );
FILL FILL_0_INVX1_78 ( );
FILL FILL_1_INVX1_78 ( );
FILL FILL_2_INVX1_78 ( );
FILL FILL_3_INVX1_78 ( );
FILL FILL_4_INVX1_78 ( );
FILL FILL_0_DFFSR_153 ( );
FILL FILL_1_DFFSR_153 ( );
FILL FILL_2_DFFSR_153 ( );
FILL FILL_3_DFFSR_153 ( );
FILL FILL_4_DFFSR_153 ( );
FILL FILL_5_DFFSR_153 ( );
FILL FILL_6_DFFSR_153 ( );
FILL FILL_7_DFFSR_153 ( );
FILL FILL_8_DFFSR_153 ( );
FILL FILL_9_DFFSR_153 ( );
FILL FILL_10_DFFSR_153 ( );
FILL FILL_11_DFFSR_153 ( );
FILL FILL_12_DFFSR_153 ( );
FILL FILL_13_DFFSR_153 ( );
FILL FILL_14_DFFSR_153 ( );
FILL FILL_15_DFFSR_153 ( );
FILL FILL_16_DFFSR_153 ( );
FILL FILL_17_DFFSR_153 ( );
FILL FILL_18_DFFSR_153 ( );
FILL FILL_19_DFFSR_153 ( );
FILL FILL_20_DFFSR_153 ( );
FILL FILL_21_DFFSR_153 ( );
FILL FILL_22_DFFSR_153 ( );
FILL FILL_23_DFFSR_153 ( );
FILL FILL_24_DFFSR_153 ( );
FILL FILL_25_DFFSR_153 ( );
FILL FILL_26_DFFSR_153 ( );
FILL FILL_27_DFFSR_153 ( );
FILL FILL_28_DFFSR_153 ( );
FILL FILL_29_DFFSR_153 ( );
FILL FILL_30_DFFSR_153 ( );
FILL FILL_31_DFFSR_153 ( );
FILL FILL_32_DFFSR_153 ( );
FILL FILL_33_DFFSR_153 ( );
FILL FILL_34_DFFSR_153 ( );
FILL FILL_35_DFFSR_153 ( );
FILL FILL_36_DFFSR_153 ( );
FILL FILL_37_DFFSR_153 ( );
FILL FILL_38_DFFSR_153 ( );
FILL FILL_39_DFFSR_153 ( );
FILL FILL_40_DFFSR_153 ( );
FILL FILL_41_DFFSR_153 ( );
FILL FILL_42_DFFSR_153 ( );
FILL FILL_43_DFFSR_153 ( );
FILL FILL_44_DFFSR_153 ( );
FILL FILL_45_DFFSR_153 ( );
FILL FILL_46_DFFSR_153 ( );
FILL FILL_47_DFFSR_153 ( );
FILL FILL_48_DFFSR_153 ( );
FILL FILL_49_DFFSR_153 ( );
FILL FILL_50_DFFSR_153 ( );
FILL FILL_0_INVX1_7 ( );
FILL FILL_1_INVX1_7 ( );
FILL FILL_2_INVX1_7 ( );
FILL FILL_3_INVX1_7 ( );
FILL FILL_4_INVX1_7 ( );
FILL FILL_0_DFFSR_8 ( );
FILL FILL_1_DFFSR_8 ( );
FILL FILL_2_DFFSR_8 ( );
FILL FILL_3_DFFSR_8 ( );
FILL FILL_4_DFFSR_8 ( );
FILL FILL_5_DFFSR_8 ( );
FILL FILL_6_DFFSR_8 ( );
FILL FILL_7_DFFSR_8 ( );
FILL FILL_8_DFFSR_8 ( );
FILL FILL_9_DFFSR_8 ( );
FILL FILL_10_DFFSR_8 ( );
FILL FILL_11_DFFSR_8 ( );
FILL FILL_12_DFFSR_8 ( );
FILL FILL_13_DFFSR_8 ( );
FILL FILL_14_DFFSR_8 ( );
FILL FILL_15_DFFSR_8 ( );
FILL FILL_16_DFFSR_8 ( );
FILL FILL_17_DFFSR_8 ( );
FILL FILL_18_DFFSR_8 ( );
FILL FILL_19_DFFSR_8 ( );
FILL FILL_20_DFFSR_8 ( );
FILL FILL_21_DFFSR_8 ( );
FILL FILL_22_DFFSR_8 ( );
FILL FILL_23_DFFSR_8 ( );
FILL FILL_24_DFFSR_8 ( );
FILL FILL_25_DFFSR_8 ( );
FILL FILL_26_DFFSR_8 ( );
FILL FILL_27_DFFSR_8 ( );
FILL FILL_28_DFFSR_8 ( );
FILL FILL_29_DFFSR_8 ( );
FILL FILL_30_DFFSR_8 ( );
FILL FILL_31_DFFSR_8 ( );
FILL FILL_32_DFFSR_8 ( );
FILL FILL_33_DFFSR_8 ( );
FILL FILL_34_DFFSR_8 ( );
FILL FILL_35_DFFSR_8 ( );
FILL FILL_36_DFFSR_8 ( );
FILL FILL_37_DFFSR_8 ( );
FILL FILL_38_DFFSR_8 ( );
FILL FILL_39_DFFSR_8 ( );
FILL FILL_40_DFFSR_8 ( );
FILL FILL_41_DFFSR_8 ( );
FILL FILL_42_DFFSR_8 ( );
FILL FILL_43_DFFSR_8 ( );
FILL FILL_44_DFFSR_8 ( );
FILL FILL_45_DFFSR_8 ( );
FILL FILL_46_DFFSR_8 ( );
FILL FILL_47_DFFSR_8 ( );
FILL FILL_48_DFFSR_8 ( );
FILL FILL_49_DFFSR_8 ( );
FILL FILL_50_DFFSR_8 ( );
FILL FILL_51_DFFSR_8 ( );
FILL FILL_0_INVX1_55 ( );
FILL FILL_1_INVX1_55 ( );
FILL FILL_2_INVX1_55 ( );
FILL FILL_3_INVX1_55 ( );
FILL FILL_4_INVX1_55 ( );
FILL FILL_0_OAI21X1_61 ( );
FILL FILL_1_OAI21X1_61 ( );
FILL FILL_2_OAI21X1_61 ( );
FILL FILL_3_OAI21X1_61 ( );
FILL FILL_4_OAI21X1_61 ( );
FILL FILL_5_OAI21X1_61 ( );
FILL FILL_6_OAI21X1_61 ( );
FILL FILL_7_OAI21X1_61 ( );
FILL FILL_8_OAI21X1_61 ( );
FILL FILL_9_OAI21X1_61 ( );
FILL FILL_0_INVX1_69 ( );
FILL FILL_1_INVX1_69 ( );
FILL FILL_2_INVX1_69 ( );
FILL FILL_3_INVX1_69 ( );
FILL FILL_0_NAND2X1_169 ( );
FILL FILL_1_NAND2X1_169 ( );
FILL FILL_2_NAND2X1_169 ( );
FILL FILL_3_NAND2X1_169 ( );
FILL FILL_4_NAND2X1_169 ( );
FILL FILL_5_NAND2X1_169 ( );
FILL FILL_6_NAND2X1_169 ( );
FILL FILL_0_DFFSR_168 ( );
FILL FILL_1_DFFSR_168 ( );
FILL FILL_2_DFFSR_168 ( );
FILL FILL_3_DFFSR_168 ( );
FILL FILL_4_DFFSR_168 ( );
FILL FILL_5_DFFSR_168 ( );
FILL FILL_6_DFFSR_168 ( );
FILL FILL_7_DFFSR_168 ( );
FILL FILL_8_DFFSR_168 ( );
FILL FILL_9_DFFSR_168 ( );
FILL FILL_10_DFFSR_168 ( );
FILL FILL_11_DFFSR_168 ( );
FILL FILL_12_DFFSR_168 ( );
FILL FILL_13_DFFSR_168 ( );
FILL FILL_14_DFFSR_168 ( );
FILL FILL_15_DFFSR_168 ( );
FILL FILL_16_DFFSR_168 ( );
FILL FILL_17_DFFSR_168 ( );
FILL FILL_18_DFFSR_168 ( );
FILL FILL_19_DFFSR_168 ( );
FILL FILL_20_DFFSR_168 ( );
FILL FILL_21_DFFSR_168 ( );
FILL FILL_22_DFFSR_168 ( );
FILL FILL_23_DFFSR_168 ( );
FILL FILL_24_DFFSR_168 ( );
FILL FILL_25_DFFSR_168 ( );
FILL FILL_26_DFFSR_168 ( );
FILL FILL_27_DFFSR_168 ( );
FILL FILL_28_DFFSR_168 ( );
FILL FILL_29_DFFSR_168 ( );
FILL FILL_30_DFFSR_168 ( );
FILL FILL_31_DFFSR_168 ( );
FILL FILL_32_DFFSR_168 ( );
FILL FILL_33_DFFSR_168 ( );
FILL FILL_34_DFFSR_168 ( );
FILL FILL_35_DFFSR_168 ( );
FILL FILL_36_DFFSR_168 ( );
FILL FILL_37_DFFSR_168 ( );
FILL FILL_38_DFFSR_168 ( );
FILL FILL_39_DFFSR_168 ( );
FILL FILL_40_DFFSR_168 ( );
FILL FILL_41_DFFSR_168 ( );
FILL FILL_42_DFFSR_168 ( );
FILL FILL_43_DFFSR_168 ( );
FILL FILL_44_DFFSR_168 ( );
FILL FILL_45_DFFSR_168 ( );
FILL FILL_46_DFFSR_168 ( );
FILL FILL_47_DFFSR_168 ( );
FILL FILL_48_DFFSR_168 ( );
FILL FILL_49_DFFSR_168 ( );
FILL FILL_50_DFFSR_168 ( );
FILL FILL_51_DFFSR_168 ( );
FILL FILL_0_INVX1_290 ( );
FILL FILL_1_INVX1_290 ( );
FILL FILL_2_INVX1_290 ( );
FILL FILL_3_INVX1_290 ( );
FILL FILL_4_INVX1_290 ( );
FILL FILL_0_OAI21X1_169 ( );
FILL FILL_1_OAI21X1_169 ( );
FILL FILL_2_OAI21X1_169 ( );
FILL FILL_3_OAI21X1_169 ( );
FILL FILL_4_OAI21X1_169 ( );
FILL FILL_5_OAI21X1_169 ( );
FILL FILL_6_OAI21X1_169 ( );
FILL FILL_7_OAI21X1_169 ( );
FILL FILL_8_OAI21X1_169 ( );
FILL FILL_9_OAI21X1_169 ( );
FILL FILL_0_INVX1_204 ( );
FILL FILL_1_INVX1_204 ( );
FILL FILL_2_INVX1_204 ( );
FILL FILL_3_INVX1_204 ( );
FILL FILL_0_XNOR2X1_2 ( );
FILL FILL_1_XNOR2X1_2 ( );
FILL FILL_2_XNOR2X1_2 ( );
FILL FILL_3_XNOR2X1_2 ( );
FILL FILL_4_XNOR2X1_2 ( );
FILL FILL_5_XNOR2X1_2 ( );
FILL FILL_6_XNOR2X1_2 ( );
FILL FILL_7_XNOR2X1_2 ( );
FILL FILL_8_XNOR2X1_2 ( );
FILL FILL_9_XNOR2X1_2 ( );
FILL FILL_10_XNOR2X1_2 ( );
FILL FILL_11_XNOR2X1_2 ( );
FILL FILL_12_XNOR2X1_2 ( );
FILL FILL_13_XNOR2X1_2 ( );
FILL FILL_14_XNOR2X1_2 ( );
FILL FILL_15_XNOR2X1_2 ( );
FILL FILL_0_OAI22X1_2 ( );
FILL FILL_1_OAI22X1_2 ( );
FILL FILL_2_OAI22X1_2 ( );
FILL FILL_3_OAI22X1_2 ( );
FILL FILL_4_OAI22X1_2 ( );
FILL FILL_5_OAI22X1_2 ( );
FILL FILL_6_OAI22X1_2 ( );
FILL FILL_7_OAI22X1_2 ( );
FILL FILL_8_OAI22X1_2 ( );
FILL FILL_9_OAI22X1_2 ( );
FILL FILL_10_OAI22X1_2 ( );
FILL FILL_11_OAI22X1_2 ( );
FILL FILL_0_OAI21X1_185 ( );
FILL FILL_1_OAI21X1_185 ( );
FILL FILL_2_OAI21X1_185 ( );
FILL FILL_3_OAI21X1_185 ( );
FILL FILL_4_OAI21X1_185 ( );
FILL FILL_5_OAI21X1_185 ( );
FILL FILL_6_OAI21X1_185 ( );
FILL FILL_7_OAI21X1_185 ( );
FILL FILL_8_OAI21X1_185 ( );
FILL FILL_0_INVX1_213 ( );
FILL FILL_1_INVX1_213 ( );
FILL FILL_2_INVX1_213 ( );
FILL FILL_3_INVX1_213 ( );
FILL FILL_4_INVX1_213 ( );
FILL FILL_0_OAI21X1_186 ( );
FILL FILL_1_OAI21X1_186 ( );
FILL FILL_2_OAI21X1_186 ( );
FILL FILL_3_OAI21X1_186 ( );
FILL FILL_4_OAI21X1_186 ( );
FILL FILL_5_OAI21X1_186 ( );
FILL FILL_6_OAI21X1_186 ( );
FILL FILL_7_OAI21X1_186 ( );
FILL FILL_8_OAI21X1_186 ( );
FILL FILL_0_OAI22X1_1 ( );
FILL FILL_1_OAI22X1_1 ( );
FILL FILL_2_OAI22X1_1 ( );
FILL FILL_3_OAI22X1_1 ( );
FILL FILL_4_OAI22X1_1 ( );
FILL FILL_5_OAI22X1_1 ( );
FILL FILL_6_OAI22X1_1 ( );
FILL FILL_7_OAI22X1_1 ( );
FILL FILL_8_OAI22X1_1 ( );
FILL FILL_9_OAI22X1_1 ( );
FILL FILL_10_OAI22X1_1 ( );
FILL FILL_0_INVX1_256 ( );
FILL FILL_1_INVX1_256 ( );
FILL FILL_2_INVX1_256 ( );
FILL FILL_3_INVX1_256 ( );
FILL FILL_4_INVX1_256 ( );
FILL FILL_0_NAND2X1_199 ( );
FILL FILL_1_NAND2X1_199 ( );
FILL FILL_2_NAND2X1_199 ( );
FILL FILL_3_NAND2X1_199 ( );
FILL FILL_4_NAND2X1_199 ( );
FILL FILL_5_NAND2X1_199 ( );
FILL FILL_6_NAND2X1_199 ( );
FILL FILL_0_OAI21X1_205 ( );
FILL FILL_1_OAI21X1_205 ( );
FILL FILL_2_OAI21X1_205 ( );
FILL FILL_3_OAI21X1_205 ( );
FILL FILL_4_OAI21X1_205 ( );
FILL FILL_5_OAI21X1_205 ( );
FILL FILL_6_OAI21X1_205 ( );
FILL FILL_7_OAI21X1_205 ( );
FILL FILL_8_OAI21X1_205 ( );
FILL FILL_9_OAI21X1_205 ( );
FILL FILL_0_NAND3X1_52 ( );
FILL FILL_1_NAND3X1_52 ( );
FILL FILL_2_NAND3X1_52 ( );
FILL FILL_3_NAND3X1_52 ( );
FILL FILL_4_NAND3X1_52 ( );
FILL FILL_5_NAND3X1_52 ( );
FILL FILL_6_NAND3X1_52 ( );
FILL FILL_7_NAND3X1_52 ( );
FILL FILL_8_NAND3X1_52 ( );
FILL FILL_0_OAI21X1_233 ( );
FILL FILL_1_OAI21X1_233 ( );
FILL FILL_2_OAI21X1_233 ( );
FILL FILL_3_OAI21X1_233 ( );
FILL FILL_4_OAI21X1_233 ( );
FILL FILL_5_OAI21X1_233 ( );
FILL FILL_6_OAI21X1_233 ( );
FILL FILL_7_OAI21X1_233 ( );
FILL FILL_8_OAI21X1_233 ( );
FILL FILL_9_OAI21X1_233 ( );
FILL FILL_0_INVX1_257 ( );
FILL FILL_1_INVX1_257 ( );
FILL FILL_2_INVX1_257 ( );
FILL FILL_3_INVX1_257 ( );
FILL FILL_4_INVX1_257 ( );
FILL FILL_0_NAND2X1_225 ( );
FILL FILL_1_NAND2X1_225 ( );
FILL FILL_2_NAND2X1_225 ( );
FILL FILL_3_NAND2X1_225 ( );
FILL FILL_4_NAND2X1_225 ( );
FILL FILL_5_NAND2X1_225 ( );
FILL FILL_6_NAND2X1_225 ( );
FILL FILL_0_INVX1_251 ( );
FILL FILL_1_INVX1_251 ( );
FILL FILL_2_INVX1_251 ( );
FILL FILL_3_INVX1_251 ( );
FILL FILL_4_INVX1_251 ( );
FILL FILL_0_NAND3X1_109 ( );
FILL FILL_1_NAND3X1_109 ( );
FILL FILL_2_NAND3X1_109 ( );
FILL FILL_3_NAND3X1_109 ( );
FILL FILL_4_NAND3X1_109 ( );
FILL FILL_5_NAND3X1_109 ( );
FILL FILL_6_NAND3X1_109 ( );
FILL FILL_7_NAND3X1_109 ( );
FILL FILL_8_NAND3X1_109 ( );
FILL FILL_0_AOI21X1_38 ( );
FILL FILL_1_AOI21X1_38 ( );
FILL FILL_2_AOI21X1_38 ( );
FILL FILL_3_AOI21X1_38 ( );
FILL FILL_4_AOI21X1_38 ( );
FILL FILL_5_AOI21X1_38 ( );
FILL FILL_6_AOI21X1_38 ( );
FILL FILL_7_AOI21X1_38 ( );
FILL FILL_8_AOI21X1_38 ( );
FILL FILL_0_INVX1_134 ( );
FILL FILL_1_INVX1_134 ( );
FILL FILL_2_INVX1_134 ( );
FILL FILL_3_INVX1_134 ( );
FILL FILL_4_INVX1_134 ( );
FILL FILL_0_NAND2X1_89 ( );
FILL FILL_1_NAND2X1_89 ( );
FILL FILL_2_NAND2X1_89 ( );
FILL FILL_3_NAND2X1_89 ( );
FILL FILL_4_NAND2X1_89 ( );
FILL FILL_5_NAND2X1_89 ( );
FILL FILL_6_NAND2X1_89 ( );
FILL FILL_0_OAI21X1_119 ( );
FILL FILL_1_OAI21X1_119 ( );
FILL FILL_2_OAI21X1_119 ( );
FILL FILL_3_OAI21X1_119 ( );
FILL FILL_4_OAI21X1_119 ( );
FILL FILL_5_OAI21X1_119 ( );
FILL FILL_6_OAI21X1_119 ( );
FILL FILL_7_OAI21X1_119 ( );
FILL FILL_8_OAI21X1_119 ( );
FILL FILL_0_NAND2X1_119 ( );
FILL FILL_1_NAND2X1_119 ( );
FILL FILL_2_NAND2X1_119 ( );
FILL FILL_3_NAND2X1_119 ( );
FILL FILL_4_NAND2X1_119 ( );
FILL FILL_5_NAND2X1_119 ( );
FILL FILL_6_NAND2X1_119 ( );
FILL FILL_0_OAI22X1_40 ( );
FILL FILL_1_OAI22X1_40 ( );
FILL FILL_2_OAI22X1_40 ( );
FILL FILL_3_OAI22X1_40 ( );
FILL FILL_4_OAI22X1_40 ( );
FILL FILL_5_OAI22X1_40 ( );
FILL FILL_6_OAI22X1_40 ( );
FILL FILL_7_OAI22X1_40 ( );
FILL FILL_8_OAI22X1_40 ( );
FILL FILL_9_OAI22X1_40 ( );
FILL FILL_10_OAI22X1_40 ( );
FILL FILL_11_OAI22X1_40 ( );
FILL FILL_0_OAI22X1_39 ( );
FILL FILL_1_OAI22X1_39 ( );
FILL FILL_2_OAI22X1_39 ( );
FILL FILL_3_OAI22X1_39 ( );
FILL FILL_4_OAI22X1_39 ( );
FILL FILL_5_OAI22X1_39 ( );
FILL FILL_6_OAI22X1_39 ( );
FILL FILL_7_OAI22X1_39 ( );
FILL FILL_8_OAI22X1_39 ( );
FILL FILL_9_OAI22X1_39 ( );
FILL FILL_10_OAI22X1_39 ( );
FILL FILL_0_OAI22X1_56 ( );
FILL FILL_1_OAI22X1_56 ( );
FILL FILL_2_OAI22X1_56 ( );
FILL FILL_3_OAI22X1_56 ( );
FILL FILL_4_OAI22X1_56 ( );
FILL FILL_5_OAI22X1_56 ( );
FILL FILL_6_OAI22X1_56 ( );
FILL FILL_7_OAI22X1_56 ( );
FILL FILL_8_OAI22X1_56 ( );
FILL FILL_9_OAI22X1_56 ( );
FILL FILL_10_OAI22X1_56 ( );
FILL FILL_11_OAI22X1_56 ( );
FILL FILL_0_INVX1_355 ( );
FILL FILL_1_INVX1_355 ( );
FILL FILL_2_INVX1_355 ( );
FILL FILL_3_INVX1_355 ( );
FILL FILL_0_OAI22X1_47 ( );
FILL FILL_1_OAI22X1_47 ( );
FILL FILL_2_OAI22X1_47 ( );
FILL FILL_3_OAI22X1_47 ( );
FILL FILL_4_OAI22X1_47 ( );
FILL FILL_5_OAI22X1_47 ( );
FILL FILL_6_OAI22X1_47 ( );
FILL FILL_7_OAI22X1_47 ( );
FILL FILL_8_OAI22X1_47 ( );
FILL FILL_9_OAI22X1_47 ( );
FILL FILL_10_OAI22X1_47 ( );
FILL FILL_11_OAI22X1_47 ( );
FILL FILL_0_INVX1_353 ( );
FILL FILL_1_INVX1_353 ( );
FILL FILL_2_INVX1_353 ( );
FILL FILL_3_INVX1_353 ( );
FILL FILL_0_OAI21X1_69 ( );
FILL FILL_1_OAI21X1_69 ( );
FILL FILL_2_OAI21X1_69 ( );
FILL FILL_3_OAI21X1_69 ( );
FILL FILL_4_OAI21X1_69 ( );
FILL FILL_5_OAI21X1_69 ( );
FILL FILL_6_OAI21X1_69 ( );
FILL FILL_7_OAI21X1_69 ( );
FILL FILL_8_OAI21X1_69 ( );
FILL FILL_0_INVX1_118 ( );
FILL FILL_1_INVX1_118 ( );
FILL FILL_2_INVX1_118 ( );
FILL FILL_3_INVX1_118 ( );
FILL FILL_0_INVX1_182 ( );
FILL FILL_1_INVX1_182 ( );
FILL FILL_2_INVX1_182 ( );
FILL FILL_3_INVX1_182 ( );
FILL FILL_4_INVX1_182 ( );
FILL FILL_0_OAI21X1_154 ( );
FILL FILL_1_OAI21X1_154 ( );
FILL FILL_2_OAI21X1_154 ( );
FILL FILL_3_OAI21X1_154 ( );
FILL FILL_4_OAI21X1_154 ( );
FILL FILL_5_OAI21X1_154 ( );
FILL FILL_6_OAI21X1_154 ( );
FILL FILL_7_OAI21X1_154 ( );
FILL FILL_8_OAI21X1_154 ( );
FILL FILL_0_NAND2X1_154 ( );
FILL FILL_1_NAND2X1_154 ( );
FILL FILL_2_NAND2X1_154 ( );
FILL FILL_3_NAND2X1_154 ( );
FILL FILL_4_NAND2X1_154 ( );
FILL FILL_5_NAND2X1_154 ( );
FILL FILL_6_NAND2X1_154 ( );
FILL FILL_0_INVX1_180 ( );
FILL FILL_1_INVX1_180 ( );
FILL FILL_2_INVX1_180 ( );
FILL FILL_3_INVX1_180 ( );
FILL FILL_4_INVX1_180 ( );
FILL FILL_0_INVX1_181 ( );
FILL FILL_1_INVX1_181 ( );
FILL FILL_2_INVX1_181 ( );
FILL FILL_3_INVX1_181 ( );
FILL FILL_4_INVX1_181 ( );
FILL FILL_0_BUFX2_9 ( );
FILL FILL_1_BUFX2_9 ( );
FILL FILL_2_BUFX2_9 ( );
FILL FILL_3_BUFX2_9 ( );
FILL FILL_4_BUFX2_9 ( );
FILL FILL_5_BUFX2_9 ( );
FILL FILL_6_BUFX2_9 ( );
FILL FILL_0_INVX1_183 ( );
FILL FILL_1_INVX1_183 ( );
FILL FILL_2_INVX1_183 ( );
FILL FILL_3_INVX1_183 ( );
FILL FILL_4_INVX1_183 ( );
FILL FILL_0_DFFSR_60 ( );
FILL FILL_1_DFFSR_60 ( );
FILL FILL_2_DFFSR_60 ( );
FILL FILL_3_DFFSR_60 ( );
FILL FILL_4_DFFSR_60 ( );
FILL FILL_5_DFFSR_60 ( );
FILL FILL_6_DFFSR_60 ( );
FILL FILL_7_DFFSR_60 ( );
FILL FILL_8_DFFSR_60 ( );
FILL FILL_9_DFFSR_60 ( );
FILL FILL_10_DFFSR_60 ( );
FILL FILL_11_DFFSR_60 ( );
FILL FILL_12_DFFSR_60 ( );
FILL FILL_13_DFFSR_60 ( );
FILL FILL_14_DFFSR_60 ( );
FILL FILL_15_DFFSR_60 ( );
FILL FILL_16_DFFSR_60 ( );
FILL FILL_17_DFFSR_60 ( );
FILL FILL_18_DFFSR_60 ( );
FILL FILL_19_DFFSR_60 ( );
FILL FILL_20_DFFSR_60 ( );
FILL FILL_21_DFFSR_60 ( );
FILL FILL_22_DFFSR_60 ( );
FILL FILL_23_DFFSR_60 ( );
FILL FILL_24_DFFSR_60 ( );
FILL FILL_25_DFFSR_60 ( );
FILL FILL_26_DFFSR_60 ( );
FILL FILL_27_DFFSR_60 ( );
FILL FILL_28_DFFSR_60 ( );
FILL FILL_29_DFFSR_60 ( );
FILL FILL_30_DFFSR_60 ( );
FILL FILL_31_DFFSR_60 ( );
FILL FILL_32_DFFSR_60 ( );
FILL FILL_33_DFFSR_60 ( );
FILL FILL_34_DFFSR_60 ( );
FILL FILL_35_DFFSR_60 ( );
FILL FILL_36_DFFSR_60 ( );
FILL FILL_37_DFFSR_60 ( );
FILL FILL_38_DFFSR_60 ( );
FILL FILL_39_DFFSR_60 ( );
FILL FILL_40_DFFSR_60 ( );
FILL FILL_41_DFFSR_60 ( );
FILL FILL_42_DFFSR_60 ( );
FILL FILL_43_DFFSR_60 ( );
FILL FILL_44_DFFSR_60 ( );
FILL FILL_45_DFFSR_60 ( );
FILL FILL_46_DFFSR_60 ( );
FILL FILL_47_DFFSR_60 ( );
FILL FILL_48_DFFSR_60 ( );
FILL FILL_49_DFFSR_60 ( );
FILL FILL_50_DFFSR_60 ( );
FILL FILL_51_DFFSR_60 ( );
FILL FILL_0_DFFPOSX1_18 ( );
FILL FILL_1_DFFPOSX1_18 ( );
FILL FILL_2_DFFPOSX1_18 ( );
FILL FILL_3_DFFPOSX1_18 ( );
FILL FILL_4_DFFPOSX1_18 ( );
FILL FILL_5_DFFPOSX1_18 ( );
FILL FILL_6_DFFPOSX1_18 ( );
FILL FILL_7_DFFPOSX1_18 ( );
FILL FILL_8_DFFPOSX1_18 ( );
FILL FILL_9_DFFPOSX1_18 ( );
FILL FILL_10_DFFPOSX1_18 ( );
FILL FILL_11_DFFPOSX1_18 ( );
FILL FILL_12_DFFPOSX1_18 ( );
FILL FILL_13_DFFPOSX1_18 ( );
FILL FILL_14_DFFPOSX1_18 ( );
FILL FILL_15_DFFPOSX1_18 ( );
FILL FILL_16_DFFPOSX1_18 ( );
FILL FILL_17_DFFPOSX1_18 ( );
FILL FILL_18_DFFPOSX1_18 ( );
FILL FILL_19_DFFPOSX1_18 ( );
FILL FILL_20_DFFPOSX1_18 ( );
FILL FILL_21_DFFPOSX1_18 ( );
FILL FILL_22_DFFPOSX1_18 ( );
FILL FILL_23_DFFPOSX1_18 ( );
FILL FILL_24_DFFPOSX1_18 ( );
FILL FILL_25_DFFPOSX1_18 ( );
FILL FILL_26_DFFPOSX1_18 ( );
FILL FILL_27_DFFPOSX1_18 ( );
FILL FILL_0_INVX1_316 ( );
FILL FILL_1_INVX1_316 ( );
FILL FILL_2_INVX1_316 ( );
FILL FILL_3_INVX1_316 ( );
FILL FILL_4_INVX1_316 ( );
FILL FILL_0_INVX1_403 ( );
FILL FILL_1_INVX1_403 ( );
FILL FILL_2_INVX1_403 ( );
FILL FILL_3_INVX1_403 ( );
FILL FILL_0_DFFPOSX1_17 ( );
FILL FILL_1_DFFPOSX1_17 ( );
FILL FILL_2_DFFPOSX1_17 ( );
FILL FILL_3_DFFPOSX1_17 ( );
FILL FILL_4_DFFPOSX1_17 ( );
FILL FILL_5_DFFPOSX1_17 ( );
FILL FILL_6_DFFPOSX1_17 ( );
FILL FILL_7_DFFPOSX1_17 ( );
FILL FILL_8_DFFPOSX1_17 ( );
FILL FILL_9_DFFPOSX1_17 ( );
FILL FILL_10_DFFPOSX1_17 ( );
FILL FILL_11_DFFPOSX1_17 ( );
FILL FILL_12_DFFPOSX1_17 ( );
FILL FILL_13_DFFPOSX1_17 ( );
FILL FILL_14_DFFPOSX1_17 ( );
FILL FILL_15_DFFPOSX1_17 ( );
FILL FILL_16_DFFPOSX1_17 ( );
FILL FILL_17_DFFPOSX1_17 ( );
FILL FILL_18_DFFPOSX1_17 ( );
FILL FILL_19_DFFPOSX1_17 ( );
FILL FILL_20_DFFPOSX1_17 ( );
FILL FILL_21_DFFPOSX1_17 ( );
FILL FILL_22_DFFPOSX1_17 ( );
FILL FILL_23_DFFPOSX1_17 ( );
FILL FILL_24_DFFPOSX1_17 ( );
FILL FILL_25_DFFPOSX1_17 ( );
FILL FILL_26_DFFPOSX1_17 ( );
FILL FILL_27_DFFPOSX1_17 ( );
FILL FILL_0_INVX1_211 ( );
FILL FILL_1_INVX1_211 ( );
FILL FILL_2_INVX1_211 ( );
FILL FILL_3_INVX1_211 ( );
FILL FILL_0_DFFSR_172 ( );
FILL FILL_1_DFFSR_172 ( );
FILL FILL_2_DFFSR_172 ( );
FILL FILL_3_DFFSR_172 ( );
FILL FILL_4_DFFSR_172 ( );
FILL FILL_5_DFFSR_172 ( );
FILL FILL_6_DFFSR_172 ( );
FILL FILL_7_DFFSR_172 ( );
FILL FILL_8_DFFSR_172 ( );
FILL FILL_9_DFFSR_172 ( );
FILL FILL_10_DFFSR_172 ( );
FILL FILL_11_DFFSR_172 ( );
FILL FILL_12_DFFSR_172 ( );
FILL FILL_13_DFFSR_172 ( );
FILL FILL_14_DFFSR_172 ( );
FILL FILL_15_DFFSR_172 ( );
FILL FILL_16_DFFSR_172 ( );
FILL FILL_17_DFFSR_172 ( );
FILL FILL_18_DFFSR_172 ( );
FILL FILL_19_DFFSR_172 ( );
FILL FILL_20_DFFSR_172 ( );
FILL FILL_21_DFFSR_172 ( );
FILL FILL_22_DFFSR_172 ( );
FILL FILL_23_DFFSR_172 ( );
FILL FILL_24_DFFSR_172 ( );
FILL FILL_25_DFFSR_172 ( );
FILL FILL_26_DFFSR_172 ( );
FILL FILL_27_DFFSR_172 ( );
FILL FILL_28_DFFSR_172 ( );
FILL FILL_29_DFFSR_172 ( );
FILL FILL_30_DFFSR_172 ( );
FILL FILL_31_DFFSR_172 ( );
FILL FILL_32_DFFSR_172 ( );
FILL FILL_33_DFFSR_172 ( );
FILL FILL_34_DFFSR_172 ( );
FILL FILL_35_DFFSR_172 ( );
FILL FILL_36_DFFSR_172 ( );
FILL FILL_37_DFFSR_172 ( );
FILL FILL_38_DFFSR_172 ( );
FILL FILL_39_DFFSR_172 ( );
FILL FILL_40_DFFSR_172 ( );
FILL FILL_41_DFFSR_172 ( );
FILL FILL_42_DFFSR_172 ( );
FILL FILL_43_DFFSR_172 ( );
FILL FILL_44_DFFSR_172 ( );
FILL FILL_45_DFFSR_172 ( );
FILL FILL_46_DFFSR_172 ( );
FILL FILL_47_DFFSR_172 ( );
FILL FILL_48_DFFSR_172 ( );
FILL FILL_49_DFFSR_172 ( );
FILL FILL_50_DFFSR_172 ( );
FILL FILL_0_NAND2X1_187 ( );
FILL FILL_1_NAND2X1_187 ( );
FILL FILL_2_NAND2X1_187 ( );
FILL FILL_3_NAND2X1_187 ( );
FILL FILL_4_NAND2X1_187 ( );
FILL FILL_5_NAND2X1_187 ( );
FILL FILL_6_NAND2X1_187 ( );
FILL FILL_0_INVX1_423 ( );
FILL FILL_1_INVX1_423 ( );
FILL FILL_2_INVX1_423 ( );
FILL FILL_3_INVX1_423 ( );
FILL FILL_4_INVX1_423 ( );
FILL FILL_0_NAND2X1_191 ( );
FILL FILL_1_NAND2X1_191 ( );
FILL FILL_2_NAND2X1_191 ( );
FILL FILL_3_NAND2X1_191 ( );
FILL FILL_4_NAND2X1_191 ( );
FILL FILL_5_NAND2X1_191 ( );
FILL FILL_6_NAND2X1_191 ( );
FILL FILL_0_OAI21X1_187 ( );
FILL FILL_1_OAI21X1_187 ( );
FILL FILL_2_OAI21X1_187 ( );
FILL FILL_3_OAI21X1_187 ( );
FILL FILL_4_OAI21X1_187 ( );
FILL FILL_5_OAI21X1_187 ( );
FILL FILL_6_OAI21X1_187 ( );
FILL FILL_7_OAI21X1_187 ( );
FILL FILL_8_OAI21X1_187 ( );
FILL FILL_0_INVX1_232 ( );
FILL FILL_1_INVX1_232 ( );
FILL FILL_2_INVX1_232 ( );
FILL FILL_3_INVX1_232 ( );
FILL FILL_4_INVX1_232 ( );
FILL FILL_0_NAND3X1_24 ( );
FILL FILL_1_NAND3X1_24 ( );
FILL FILL_2_NAND3X1_24 ( );
FILL FILL_3_NAND3X1_24 ( );
FILL FILL_4_NAND3X1_24 ( );
FILL FILL_5_NAND3X1_24 ( );
FILL FILL_6_NAND3X1_24 ( );
FILL FILL_7_NAND3X1_24 ( );
FILL FILL_8_NAND3X1_24 ( );
FILL FILL_9_NAND3X1_24 ( );
FILL FILL_0_NAND3X1_20 ( );
FILL FILL_1_NAND3X1_20 ( );
FILL FILL_2_NAND3X1_20 ( );
FILL FILL_3_NAND3X1_20 ( );
FILL FILL_4_NAND3X1_20 ( );
FILL FILL_5_NAND3X1_20 ( );
FILL FILL_6_NAND3X1_20 ( );
FILL FILL_7_NAND3X1_20 ( );
FILL FILL_8_NAND3X1_20 ( );
FILL FILL_0_NAND2X1_184 ( );
FILL FILL_1_NAND2X1_184 ( );
FILL FILL_2_NAND2X1_184 ( );
FILL FILL_3_NAND2X1_184 ( );
FILL FILL_4_NAND2X1_184 ( );
FILL FILL_5_NAND2X1_184 ( );
FILL FILL_6_NAND2X1_184 ( );
FILL FILL_0_OAI21X1_191 ( );
FILL FILL_1_OAI21X1_191 ( );
FILL FILL_2_OAI21X1_191 ( );
FILL FILL_3_OAI21X1_191 ( );
FILL FILL_4_OAI21X1_191 ( );
FILL FILL_5_OAI21X1_191 ( );
FILL FILL_6_OAI21X1_191 ( );
FILL FILL_7_OAI21X1_191 ( );
FILL FILL_8_OAI21X1_191 ( );
FILL FILL_0_OAI21X1_200 ( );
FILL FILL_1_OAI21X1_200 ( );
FILL FILL_2_OAI21X1_200 ( );
FILL FILL_3_OAI21X1_200 ( );
FILL FILL_4_OAI21X1_200 ( );
FILL FILL_5_OAI21X1_200 ( );
FILL FILL_6_OAI21X1_200 ( );
FILL FILL_7_OAI21X1_200 ( );
FILL FILL_8_OAI21X1_200 ( );
FILL FILL_9_OAI21X1_200 ( );
FILL FILL_0_OAI21X1_207 ( );
FILL FILL_1_OAI21X1_207 ( );
FILL FILL_2_OAI21X1_207 ( );
FILL FILL_3_OAI21X1_207 ( );
FILL FILL_4_OAI21X1_207 ( );
FILL FILL_5_OAI21X1_207 ( );
FILL FILL_6_OAI21X1_207 ( );
FILL FILL_7_OAI21X1_207 ( );
FILL FILL_8_OAI21X1_207 ( );
FILL FILL_9_OAI21X1_207 ( );
FILL FILL_0_NAND3X1_49 ( );
FILL FILL_1_NAND3X1_49 ( );
FILL FILL_2_NAND3X1_49 ( );
FILL FILL_3_NAND3X1_49 ( );
FILL FILL_4_NAND3X1_49 ( );
FILL FILL_5_NAND3X1_49 ( );
FILL FILL_6_NAND3X1_49 ( );
FILL FILL_7_NAND3X1_49 ( );
FILL FILL_8_NAND3X1_49 ( );
FILL FILL_0_NAND2X1_268 ( );
FILL FILL_1_NAND2X1_268 ( );
FILL FILL_2_NAND2X1_268 ( );
FILL FILL_3_NAND2X1_268 ( );
FILL FILL_4_NAND2X1_268 ( );
FILL FILL_5_NAND2X1_268 ( );
FILL FILL_6_NAND2X1_268 ( );
FILL FILL_0_DFFPOSX1_9 ( );
FILL FILL_1_DFFPOSX1_9 ( );
FILL FILL_2_DFFPOSX1_9 ( );
FILL FILL_3_DFFPOSX1_9 ( );
FILL FILL_4_DFFPOSX1_9 ( );
FILL FILL_5_DFFPOSX1_9 ( );
FILL FILL_6_DFFPOSX1_9 ( );
FILL FILL_7_DFFPOSX1_9 ( );
FILL FILL_8_DFFPOSX1_9 ( );
FILL FILL_9_DFFPOSX1_9 ( );
FILL FILL_10_DFFPOSX1_9 ( );
FILL FILL_11_DFFPOSX1_9 ( );
FILL FILL_12_DFFPOSX1_9 ( );
FILL FILL_13_DFFPOSX1_9 ( );
FILL FILL_14_DFFPOSX1_9 ( );
FILL FILL_15_DFFPOSX1_9 ( );
FILL FILL_16_DFFPOSX1_9 ( );
FILL FILL_17_DFFPOSX1_9 ( );
FILL FILL_18_DFFPOSX1_9 ( );
FILL FILL_19_DFFPOSX1_9 ( );
FILL FILL_20_DFFPOSX1_9 ( );
FILL FILL_21_DFFPOSX1_9 ( );
FILL FILL_22_DFFPOSX1_9 ( );
FILL FILL_23_DFFPOSX1_9 ( );
FILL FILL_24_DFFPOSX1_9 ( );
FILL FILL_25_DFFPOSX1_9 ( );
FILL FILL_26_DFFPOSX1_9 ( );
FILL FILL_27_DFFPOSX1_9 ( );
FILL FILL_0_DFFSR_119 ( );
FILL FILL_1_DFFSR_119 ( );
FILL FILL_2_DFFSR_119 ( );
FILL FILL_3_DFFSR_119 ( );
FILL FILL_4_DFFSR_119 ( );
FILL FILL_5_DFFSR_119 ( );
FILL FILL_6_DFFSR_119 ( );
FILL FILL_7_DFFSR_119 ( );
FILL FILL_8_DFFSR_119 ( );
FILL FILL_9_DFFSR_119 ( );
FILL FILL_10_DFFSR_119 ( );
FILL FILL_11_DFFSR_119 ( );
FILL FILL_12_DFFSR_119 ( );
FILL FILL_13_DFFSR_119 ( );
FILL FILL_14_DFFSR_119 ( );
FILL FILL_15_DFFSR_119 ( );
FILL FILL_16_DFFSR_119 ( );
FILL FILL_17_DFFSR_119 ( );
FILL FILL_18_DFFSR_119 ( );
FILL FILL_19_DFFSR_119 ( );
FILL FILL_20_DFFSR_119 ( );
FILL FILL_21_DFFSR_119 ( );
FILL FILL_22_DFFSR_119 ( );
FILL FILL_23_DFFSR_119 ( );
FILL FILL_24_DFFSR_119 ( );
FILL FILL_25_DFFSR_119 ( );
FILL FILL_26_DFFSR_119 ( );
FILL FILL_27_DFFSR_119 ( );
FILL FILL_28_DFFSR_119 ( );
FILL FILL_29_DFFSR_119 ( );
FILL FILL_30_DFFSR_119 ( );
FILL FILL_31_DFFSR_119 ( );
FILL FILL_32_DFFSR_119 ( );
FILL FILL_33_DFFSR_119 ( );
FILL FILL_34_DFFSR_119 ( );
FILL FILL_35_DFFSR_119 ( );
FILL FILL_36_DFFSR_119 ( );
FILL FILL_37_DFFSR_119 ( );
FILL FILL_38_DFFSR_119 ( );
FILL FILL_39_DFFSR_119 ( );
FILL FILL_40_DFFSR_119 ( );
FILL FILL_41_DFFSR_119 ( );
FILL FILL_42_DFFSR_119 ( );
FILL FILL_43_DFFSR_119 ( );
FILL FILL_44_DFFSR_119 ( );
FILL FILL_45_DFFSR_119 ( );
FILL FILL_46_DFFSR_119 ( );
FILL FILL_47_DFFSR_119 ( );
FILL FILL_48_DFFSR_119 ( );
FILL FILL_49_DFFSR_119 ( );
FILL FILL_50_DFFSR_119 ( );
FILL FILL_0_NOR2X1_29 ( );
FILL FILL_1_NOR2X1_29 ( );
FILL FILL_2_NOR2X1_29 ( );
FILL FILL_3_NOR2X1_29 ( );
FILL FILL_4_NOR2X1_29 ( );
FILL FILL_5_NOR2X1_29 ( );
FILL FILL_6_NOR2X1_29 ( );
FILL FILL_0_INVX1_366 ( );
FILL FILL_1_INVX1_366 ( );
FILL FILL_2_INVX1_366 ( );
FILL FILL_3_INVX1_366 ( );
FILL FILL_4_INVX1_366 ( );
FILL FILL_0_OAI22X1_48 ( );
FILL FILL_1_OAI22X1_48 ( );
FILL FILL_2_OAI22X1_48 ( );
FILL FILL_3_OAI22X1_48 ( );
FILL FILL_4_OAI22X1_48 ( );
FILL FILL_5_OAI22X1_48 ( );
FILL FILL_6_OAI22X1_48 ( );
FILL FILL_7_OAI22X1_48 ( );
FILL FILL_8_OAI22X1_48 ( );
FILL FILL_9_OAI22X1_48 ( );
FILL FILL_10_OAI22X1_48 ( );
FILL FILL_11_OAI22X1_48 ( );
FILL FILL_0_NOR2X1_33 ( );
FILL FILL_1_NOR2X1_33 ( );
FILL FILL_2_NOR2X1_33 ( );
FILL FILL_3_NOR2X1_33 ( );
FILL FILL_4_NOR2X1_33 ( );
FILL FILL_5_NOR2X1_33 ( );
FILL FILL_6_NOR2X1_33 ( );
FILL FILL_0_INVX1_77 ( );
FILL FILL_1_INVX1_77 ( );
FILL FILL_2_INVX1_77 ( );
FILL FILL_3_INVX1_77 ( );
FILL FILL_4_INVX1_77 ( );
FILL FILL_0_OAI21X1_68 ( );
FILL FILL_1_OAI21X1_68 ( );
FILL FILL_2_OAI21X1_68 ( );
FILL FILL_3_OAI21X1_68 ( );
FILL FILL_4_OAI21X1_68 ( );
FILL FILL_5_OAI21X1_68 ( );
FILL FILL_6_OAI21X1_68 ( );
FILL FILL_7_OAI21X1_68 ( );
FILL FILL_8_OAI21X1_68 ( );
FILL FILL_0_NAND2X1_155 ( );
FILL FILL_1_NAND2X1_155 ( );
FILL FILL_2_NAND2X1_155 ( );
FILL FILL_3_NAND2X1_155 ( );
FILL FILL_4_NAND2X1_155 ( );
FILL FILL_5_NAND2X1_155 ( );
FILL FILL_6_NAND2X1_155 ( );
FILL FILL_0_INVX1_176 ( );
FILL FILL_1_INVX1_176 ( );
FILL FILL_2_INVX1_176 ( );
FILL FILL_3_INVX1_176 ( );
FILL FILL_4_INVX1_176 ( );
FILL FILL_0_NAND2X1_150 ( );
FILL FILL_1_NAND2X1_150 ( );
FILL FILL_2_NAND2X1_150 ( );
FILL FILL_3_NAND2X1_150 ( );
FILL FILL_4_NAND2X1_150 ( );
FILL FILL_5_NAND2X1_150 ( );
FILL FILL_6_NAND2X1_150 ( );
FILL FILL_0_OAI21X1_151 ( );
FILL FILL_1_OAI21X1_151 ( );
FILL FILL_2_OAI21X1_151 ( );
FILL FILL_3_OAI21X1_151 ( );
FILL FILL_4_OAI21X1_151 ( );
FILL FILL_5_OAI21X1_151 ( );
FILL FILL_6_OAI21X1_151 ( );
FILL FILL_7_OAI21X1_151 ( );
FILL FILL_8_OAI21X1_151 ( );
FILL FILL_0_INVX1_177 ( );
FILL FILL_1_INVX1_177 ( );
FILL FILL_2_INVX1_177 ( );
FILL FILL_3_INVX1_177 ( );
FILL FILL_4_INVX1_177 ( );
FILL FILL_0_INVX1_1 ( );
FILL FILL_1_INVX1_1 ( );
FILL FILL_2_INVX1_1 ( );
FILL FILL_3_INVX1_1 ( );
FILL FILL_0_DFFSR_133 ( );
FILL FILL_1_DFFSR_133 ( );
FILL FILL_2_DFFSR_133 ( );
FILL FILL_3_DFFSR_133 ( );
FILL FILL_4_DFFSR_133 ( );
FILL FILL_5_DFFSR_133 ( );
FILL FILL_6_DFFSR_133 ( );
FILL FILL_7_DFFSR_133 ( );
FILL FILL_8_DFFSR_133 ( );
FILL FILL_9_DFFSR_133 ( );
FILL FILL_10_DFFSR_133 ( );
FILL FILL_11_DFFSR_133 ( );
FILL FILL_12_DFFSR_133 ( );
FILL FILL_13_DFFSR_133 ( );
FILL FILL_14_DFFSR_133 ( );
FILL FILL_15_DFFSR_133 ( );
FILL FILL_16_DFFSR_133 ( );
FILL FILL_17_DFFSR_133 ( );
FILL FILL_18_DFFSR_133 ( );
FILL FILL_19_DFFSR_133 ( );
FILL FILL_20_DFFSR_133 ( );
FILL FILL_21_DFFSR_133 ( );
FILL FILL_22_DFFSR_133 ( );
FILL FILL_23_DFFSR_133 ( );
FILL FILL_24_DFFSR_133 ( );
FILL FILL_25_DFFSR_133 ( );
FILL FILL_26_DFFSR_133 ( );
FILL FILL_27_DFFSR_133 ( );
FILL FILL_28_DFFSR_133 ( );
FILL FILL_29_DFFSR_133 ( );
FILL FILL_30_DFFSR_133 ( );
FILL FILL_31_DFFSR_133 ( );
FILL FILL_32_DFFSR_133 ( );
FILL FILL_33_DFFSR_133 ( );
FILL FILL_34_DFFSR_133 ( );
FILL FILL_35_DFFSR_133 ( );
FILL FILL_36_DFFSR_133 ( );
FILL FILL_37_DFFSR_133 ( );
FILL FILL_38_DFFSR_133 ( );
FILL FILL_39_DFFSR_133 ( );
FILL FILL_40_DFFSR_133 ( );
FILL FILL_41_DFFSR_133 ( );
FILL FILL_42_DFFSR_133 ( );
FILL FILL_43_DFFSR_133 ( );
FILL FILL_44_DFFSR_133 ( );
FILL FILL_45_DFFSR_133 ( );
FILL FILL_46_DFFSR_133 ( );
FILL FILL_47_DFFSR_133 ( );
FILL FILL_48_DFFSR_133 ( );
FILL FILL_49_DFFSR_133 ( );
FILL FILL_50_DFFSR_133 ( );
FILL FILL_0_INVX1_68 ( );
FILL FILL_1_INVX1_68 ( );
FILL FILL_2_INVX1_68 ( );
FILL FILL_3_INVX1_68 ( );
FILL FILL_0_OAI21X1_60 ( );
FILL FILL_1_OAI21X1_60 ( );
FILL FILL_2_OAI21X1_60 ( );
FILL FILL_3_OAI21X1_60 ( );
FILL FILL_4_OAI21X1_60 ( );
FILL FILL_5_OAI21X1_60 ( );
FILL FILL_6_OAI21X1_60 ( );
FILL FILL_7_OAI21X1_60 ( );
FILL FILL_8_OAI21X1_60 ( );
FILL FILL_9_OAI21X1_60 ( );
FILL FILL_0_BUFX2_37 ( );
FILL FILL_1_BUFX2_37 ( );
FILL FILL_2_BUFX2_37 ( );
FILL FILL_3_BUFX2_37 ( );
FILL FILL_4_BUFX2_37 ( );
FILL FILL_5_BUFX2_37 ( );
FILL FILL_6_BUFX2_37 ( );
FILL FILL_0_BUFX2_41 ( );
FILL FILL_1_BUFX2_41 ( );
FILL FILL_2_BUFX2_41 ( );
FILL FILL_3_BUFX2_41 ( );
FILL FILL_4_BUFX2_41 ( );
FILL FILL_5_BUFX2_41 ( );
FILL FILL_6_BUFX2_41 ( );
FILL FILL_0_INVX1_52 ( );
FILL FILL_1_INVX1_52 ( );
FILL FILL_2_INVX1_52 ( );
FILL FILL_3_INVX1_52 ( );
FILL FILL_4_INVX1_52 ( );
FILL FILL_0_OAI21X1_46 ( );
FILL FILL_1_OAI21X1_46 ( );
FILL FILL_2_OAI21X1_46 ( );
FILL FILL_3_OAI21X1_46 ( );
FILL FILL_4_OAI21X1_46 ( );
FILL FILL_5_OAI21X1_46 ( );
FILL FILL_6_OAI21X1_46 ( );
FILL FILL_7_OAI21X1_46 ( );
FILL FILL_8_OAI21X1_46 ( );
FILL FILL_0_BUFX2_38 ( );
FILL FILL_1_BUFX2_38 ( );
FILL FILL_2_BUFX2_38 ( );
FILL FILL_3_BUFX2_38 ( );
FILL FILL_4_BUFX2_38 ( );
FILL FILL_5_BUFX2_38 ( );
FILL FILL_6_BUFX2_38 ( );
FILL FILL_0_NAND2X1_61 ( );
FILL FILL_1_NAND2X1_61 ( );
FILL FILL_2_NAND2X1_61 ( );
FILL FILL_3_NAND2X1_61 ( );
FILL FILL_4_NAND2X1_61 ( );
FILL FILL_5_NAND2X1_61 ( );
FILL FILL_6_NAND2X1_61 ( );
FILL FILL_0_BUFX2_34 ( );
FILL FILL_1_BUFX2_34 ( );
FILL FILL_2_BUFX2_34 ( );
FILL FILL_3_BUFX2_34 ( );
FILL FILL_4_BUFX2_34 ( );
FILL FILL_5_BUFX2_34 ( );
FILL FILL_6_BUFX2_34 ( );
FILL FILL_0_DFFPOSX1_26 ( );
FILL FILL_1_DFFPOSX1_26 ( );
FILL FILL_2_DFFPOSX1_26 ( );
FILL FILL_3_DFFPOSX1_26 ( );
FILL FILL_4_DFFPOSX1_26 ( );
FILL FILL_5_DFFPOSX1_26 ( );
FILL FILL_6_DFFPOSX1_26 ( );
FILL FILL_7_DFFPOSX1_26 ( );
FILL FILL_8_DFFPOSX1_26 ( );
FILL FILL_9_DFFPOSX1_26 ( );
FILL FILL_10_DFFPOSX1_26 ( );
FILL FILL_11_DFFPOSX1_26 ( );
FILL FILL_12_DFFPOSX1_26 ( );
FILL FILL_13_DFFPOSX1_26 ( );
FILL FILL_14_DFFPOSX1_26 ( );
FILL FILL_15_DFFPOSX1_26 ( );
FILL FILL_16_DFFPOSX1_26 ( );
FILL FILL_17_DFFPOSX1_26 ( );
FILL FILL_18_DFFPOSX1_26 ( );
FILL FILL_19_DFFPOSX1_26 ( );
FILL FILL_20_DFFPOSX1_26 ( );
FILL FILL_21_DFFPOSX1_26 ( );
FILL FILL_22_DFFPOSX1_26 ( );
FILL FILL_23_DFFPOSX1_26 ( );
FILL FILL_24_DFFPOSX1_26 ( );
FILL FILL_25_DFFPOSX1_26 ( );
FILL FILL_26_DFFPOSX1_26 ( );
FILL FILL_27_DFFPOSX1_26 ( );
FILL FILL_0_BUFX2_14 ( );
FILL FILL_1_BUFX2_14 ( );
FILL FILL_2_BUFX2_14 ( );
FILL FILL_3_BUFX2_14 ( );
FILL FILL_4_BUFX2_14 ( );
FILL FILL_5_BUFX2_14 ( );
FILL FILL_6_BUFX2_14 ( );
FILL FILL_0_AOI22X1_6 ( );
FILL FILL_1_AOI22X1_6 ( );
FILL FILL_2_AOI22X1_6 ( );
FILL FILL_3_AOI22X1_6 ( );
FILL FILL_4_AOI22X1_6 ( );
FILL FILL_5_AOI22X1_6 ( );
FILL FILL_6_AOI22X1_6 ( );
FILL FILL_7_AOI22X1_6 ( );
FILL FILL_8_AOI22X1_6 ( );
FILL FILL_9_AOI22X1_6 ( );
FILL FILL_10_AOI22X1_6 ( );
FILL FILL_11_AOI22X1_6 ( );
FILL FILL_0_BUFX2_12 ( );
FILL FILL_1_BUFX2_12 ( );
FILL FILL_2_BUFX2_12 ( );
FILL FILL_3_BUFX2_12 ( );
FILL FILL_4_BUFX2_12 ( );
FILL FILL_5_BUFX2_12 ( );
FILL FILL_6_BUFX2_12 ( );
FILL FILL_0_AOI22X1_2 ( );
FILL FILL_1_AOI22X1_2 ( );
FILL FILL_2_AOI22X1_2 ( );
FILL FILL_3_AOI22X1_2 ( );
FILL FILL_4_AOI22X1_2 ( );
FILL FILL_5_AOI22X1_2 ( );
FILL FILL_6_AOI22X1_2 ( );
FILL FILL_7_AOI22X1_2 ( );
FILL FILL_8_AOI22X1_2 ( );
FILL FILL_9_AOI22X1_2 ( );
FILL FILL_10_AOI22X1_2 ( );
FILL FILL_11_AOI22X1_2 ( );
FILL FILL_0_AND2X2_5 ( );
FILL FILL_1_AND2X2_5 ( );
FILL FILL_2_AND2X2_5 ( );
FILL FILL_3_AND2X2_5 ( );
FILL FILL_4_AND2X2_5 ( );
FILL FILL_5_AND2X2_5 ( );
FILL FILL_6_AND2X2_5 ( );
FILL FILL_7_AND2X2_5 ( );
FILL FILL_8_AND2X2_5 ( );
FILL FILL_0_INVX1_202 ( );
FILL FILL_1_INVX1_202 ( );
FILL FILL_2_INVX1_202 ( );
FILL FILL_3_INVX1_202 ( );
FILL FILL_4_INVX1_202 ( );
FILL FILL_0_NAND3X1_22 ( );
FILL FILL_1_NAND3X1_22 ( );
FILL FILL_2_NAND3X1_22 ( );
FILL FILL_3_NAND3X1_22 ( );
FILL FILL_4_NAND3X1_22 ( );
FILL FILL_5_NAND3X1_22 ( );
FILL FILL_6_NAND3X1_22 ( );
FILL FILL_7_NAND3X1_22 ( );
FILL FILL_8_NAND3X1_22 ( );
FILL FILL_0_NAND2X1_186 ( );
FILL FILL_1_NAND2X1_186 ( );
FILL FILL_2_NAND2X1_186 ( );
FILL FILL_3_NAND2X1_186 ( );
FILL FILL_4_NAND2X1_186 ( );
FILL FILL_5_NAND2X1_186 ( );
FILL FILL_6_NAND2X1_186 ( );
FILL FILL_0_OAI21X1_192 ( );
FILL FILL_1_OAI21X1_192 ( );
FILL FILL_2_OAI21X1_192 ( );
FILL FILL_3_OAI21X1_192 ( );
FILL FILL_4_OAI21X1_192 ( );
FILL FILL_5_OAI21X1_192 ( );
FILL FILL_6_OAI21X1_192 ( );
FILL FILL_7_OAI21X1_192 ( );
FILL FILL_8_OAI21X1_192 ( );
FILL FILL_0_AOI21X1_5 ( );
FILL FILL_1_AOI21X1_5 ( );
FILL FILL_2_AOI21X1_5 ( );
FILL FILL_3_AOI21X1_5 ( );
FILL FILL_4_AOI21X1_5 ( );
FILL FILL_5_AOI21X1_5 ( );
FILL FILL_6_AOI21X1_5 ( );
FILL FILL_7_AOI21X1_5 ( );
FILL FILL_8_AOI21X1_5 ( );
FILL FILL_0_NAND3X1_23 ( );
FILL FILL_1_NAND3X1_23 ( );
FILL FILL_2_NAND3X1_23 ( );
FILL FILL_3_NAND3X1_23 ( );
FILL FILL_4_NAND3X1_23 ( );
FILL FILL_5_NAND3X1_23 ( );
FILL FILL_6_NAND3X1_23 ( );
FILL FILL_7_NAND3X1_23 ( );
FILL FILL_8_NAND3X1_23 ( );
FILL FILL_9_NAND3X1_23 ( );
FILL FILL_0_NAND3X1_27 ( );
FILL FILL_1_NAND3X1_27 ( );
FILL FILL_2_NAND3X1_27 ( );
FILL FILL_3_NAND3X1_27 ( );
FILL FILL_4_NAND3X1_27 ( );
FILL FILL_5_NAND3X1_27 ( );
FILL FILL_6_NAND3X1_27 ( );
FILL FILL_7_NAND3X1_27 ( );
FILL FILL_8_NAND3X1_27 ( );
FILL FILL_9_NAND3X1_27 ( );
FILL FILL_0_INVX1_238 ( );
FILL FILL_1_INVX1_238 ( );
FILL FILL_2_INVX1_238 ( );
FILL FILL_3_INVX1_238 ( );
FILL FILL_0_NAND3X1_53 ( );
FILL FILL_1_NAND3X1_53 ( );
FILL FILL_2_NAND3X1_53 ( );
FILL FILL_3_NAND3X1_53 ( );
FILL FILL_4_NAND3X1_53 ( );
FILL FILL_5_NAND3X1_53 ( );
FILL FILL_6_NAND3X1_53 ( );
FILL FILL_7_NAND3X1_53 ( );
FILL FILL_8_NAND3X1_53 ( );
FILL FILL_0_NAND3X1_50 ( );
FILL FILL_1_NAND3X1_50 ( );
FILL FILL_2_NAND3X1_50 ( );
FILL FILL_3_NAND3X1_50 ( );
FILL FILL_4_NAND3X1_50 ( );
FILL FILL_5_NAND3X1_50 ( );
FILL FILL_6_NAND3X1_50 ( );
FILL FILL_7_NAND3X1_50 ( );
FILL FILL_8_NAND3X1_50 ( );
FILL FILL_0_NAND3X1_83 ( );
FILL FILL_1_NAND3X1_83 ( );
FILL FILL_2_NAND3X1_83 ( );
FILL FILL_3_NAND3X1_83 ( );
FILL FILL_4_NAND3X1_83 ( );
FILL FILL_5_NAND3X1_83 ( );
FILL FILL_6_NAND3X1_83 ( );
FILL FILL_7_NAND3X1_83 ( );
FILL FILL_8_NAND3X1_83 ( );
FILL FILL_0_NAND3X1_77 ( );
FILL FILL_1_NAND3X1_77 ( );
FILL FILL_2_NAND3X1_77 ( );
FILL FILL_3_NAND3X1_77 ( );
FILL FILL_4_NAND3X1_77 ( );
FILL FILL_5_NAND3X1_77 ( );
FILL FILL_6_NAND3X1_77 ( );
FILL FILL_7_NAND3X1_77 ( );
FILL FILL_8_NAND3X1_77 ( );
FILL FILL_0_NAND2X1_231 ( );
FILL FILL_1_NAND2X1_231 ( );
FILL FILL_2_NAND2X1_231 ( );
FILL FILL_3_NAND2X1_231 ( );
FILL FILL_4_NAND2X1_231 ( );
FILL FILL_5_NAND2X1_231 ( );
FILL FILL_6_NAND2X1_231 ( );
FILL FILL_0_NAND3X1_108 ( );
FILL FILL_1_NAND3X1_108 ( );
FILL FILL_2_NAND3X1_108 ( );
FILL FILL_3_NAND3X1_108 ( );
FILL FILL_4_NAND3X1_108 ( );
FILL FILL_5_NAND3X1_108 ( );
FILL FILL_6_NAND3X1_108 ( );
FILL FILL_7_NAND3X1_108 ( );
FILL FILL_8_NAND3X1_108 ( );
FILL FILL_0_INVX1_259 ( );
FILL FILL_1_INVX1_259 ( );
FILL FILL_2_INVX1_259 ( );
FILL FILL_3_INVX1_259 ( );
FILL FILL_0_DFFSR_81 ( );
FILL FILL_1_DFFSR_81 ( );
FILL FILL_2_DFFSR_81 ( );
FILL FILL_3_DFFSR_81 ( );
FILL FILL_4_DFFSR_81 ( );
FILL FILL_5_DFFSR_81 ( );
FILL FILL_6_DFFSR_81 ( );
FILL FILL_7_DFFSR_81 ( );
FILL FILL_8_DFFSR_81 ( );
FILL FILL_9_DFFSR_81 ( );
FILL FILL_10_DFFSR_81 ( );
FILL FILL_11_DFFSR_81 ( );
FILL FILL_12_DFFSR_81 ( );
FILL FILL_13_DFFSR_81 ( );
FILL FILL_14_DFFSR_81 ( );
FILL FILL_15_DFFSR_81 ( );
FILL FILL_16_DFFSR_81 ( );
FILL FILL_17_DFFSR_81 ( );
FILL FILL_18_DFFSR_81 ( );
FILL FILL_19_DFFSR_81 ( );
FILL FILL_20_DFFSR_81 ( );
FILL FILL_21_DFFSR_81 ( );
FILL FILL_22_DFFSR_81 ( );
FILL FILL_23_DFFSR_81 ( );
FILL FILL_24_DFFSR_81 ( );
FILL FILL_25_DFFSR_81 ( );
FILL FILL_26_DFFSR_81 ( );
FILL FILL_27_DFFSR_81 ( );
FILL FILL_28_DFFSR_81 ( );
FILL FILL_29_DFFSR_81 ( );
FILL FILL_30_DFFSR_81 ( );
FILL FILL_31_DFFSR_81 ( );
FILL FILL_32_DFFSR_81 ( );
FILL FILL_33_DFFSR_81 ( );
FILL FILL_34_DFFSR_81 ( );
FILL FILL_35_DFFSR_81 ( );
FILL FILL_36_DFFSR_81 ( );
FILL FILL_37_DFFSR_81 ( );
FILL FILL_38_DFFSR_81 ( );
FILL FILL_39_DFFSR_81 ( );
FILL FILL_40_DFFSR_81 ( );
FILL FILL_41_DFFSR_81 ( );
FILL FILL_42_DFFSR_81 ( );
FILL FILL_43_DFFSR_81 ( );
FILL FILL_44_DFFSR_81 ( );
FILL FILL_45_DFFSR_81 ( );
FILL FILL_46_DFFSR_81 ( );
FILL FILL_47_DFFSR_81 ( );
FILL FILL_48_DFFSR_81 ( );
FILL FILL_49_DFFSR_81 ( );
FILL FILL_50_DFFSR_81 ( );
FILL FILL_51_DFFSR_81 ( );
FILL FILL_0_INVX1_334 ( );
FILL FILL_1_INVX1_334 ( );
FILL FILL_2_INVX1_334 ( );
FILL FILL_3_INVX1_334 ( );
FILL FILL_4_INVX1_334 ( );
FILL FILL_0_INVX1_360 ( );
FILL FILL_1_INVX1_360 ( );
FILL FILL_2_INVX1_360 ( );
FILL FILL_3_INVX1_360 ( );
FILL FILL_4_INVX1_360 ( );
FILL FILL_0_INVX1_361 ( );
FILL FILL_1_INVX1_361 ( );
FILL FILL_2_INVX1_361 ( );
FILL FILL_3_INVX1_361 ( );
FILL FILL_0_OAI22X1_51 ( );
FILL FILL_1_OAI22X1_51 ( );
FILL FILL_2_OAI22X1_51 ( );
FILL FILL_3_OAI22X1_51 ( );
FILL FILL_4_OAI22X1_51 ( );
FILL FILL_5_OAI22X1_51 ( );
FILL FILL_6_OAI22X1_51 ( );
FILL FILL_7_OAI22X1_51 ( );
FILL FILL_8_OAI22X1_51 ( );
FILL FILL_9_OAI22X1_51 ( );
FILL FILL_10_OAI22X1_51 ( );
FILL FILL_11_OAI22X1_51 ( );
FILL FILL_0_OAI21X1_155 ( );
FILL FILL_1_OAI21X1_155 ( );
FILL FILL_2_OAI21X1_155 ( );
FILL FILL_3_OAI21X1_155 ( );
FILL FILL_4_OAI21X1_155 ( );
FILL FILL_5_OAI21X1_155 ( );
FILL FILL_6_OAI21X1_155 ( );
FILL FILL_7_OAI21X1_155 ( );
FILL FILL_8_OAI21X1_155 ( );
FILL FILL_0_INVX1_184 ( );
FILL FILL_1_INVX1_184 ( );
FILL FILL_2_INVX1_184 ( );
FILL FILL_3_INVX1_184 ( );
FILL FILL_4_INVX1_184 ( );
FILL FILL_0_INVX1_350 ( );
FILL FILL_1_INVX1_350 ( );
FILL FILL_2_INVX1_350 ( );
FILL FILL_3_INVX1_350 ( );
FILL FILL_4_INVX1_350 ( );
FILL FILL_0_DFFSR_151 ( );
FILL FILL_1_DFFSR_151 ( );
FILL FILL_2_DFFSR_151 ( );
FILL FILL_3_DFFSR_151 ( );
FILL FILL_4_DFFSR_151 ( );
FILL FILL_5_DFFSR_151 ( );
FILL FILL_6_DFFSR_151 ( );
FILL FILL_7_DFFSR_151 ( );
FILL FILL_8_DFFSR_151 ( );
FILL FILL_9_DFFSR_151 ( );
FILL FILL_10_DFFSR_151 ( );
FILL FILL_11_DFFSR_151 ( );
FILL FILL_12_DFFSR_151 ( );
FILL FILL_13_DFFSR_151 ( );
FILL FILL_14_DFFSR_151 ( );
FILL FILL_15_DFFSR_151 ( );
FILL FILL_16_DFFSR_151 ( );
FILL FILL_17_DFFSR_151 ( );
FILL FILL_18_DFFSR_151 ( );
FILL FILL_19_DFFSR_151 ( );
FILL FILL_20_DFFSR_151 ( );
FILL FILL_21_DFFSR_151 ( );
FILL FILL_22_DFFSR_151 ( );
FILL FILL_23_DFFSR_151 ( );
FILL FILL_24_DFFSR_151 ( );
FILL FILL_25_DFFSR_151 ( );
FILL FILL_26_DFFSR_151 ( );
FILL FILL_27_DFFSR_151 ( );
FILL FILL_28_DFFSR_151 ( );
FILL FILL_29_DFFSR_151 ( );
FILL FILL_30_DFFSR_151 ( );
FILL FILL_31_DFFSR_151 ( );
FILL FILL_32_DFFSR_151 ( );
FILL FILL_33_DFFSR_151 ( );
FILL FILL_34_DFFSR_151 ( );
FILL FILL_35_DFFSR_151 ( );
FILL FILL_36_DFFSR_151 ( );
FILL FILL_37_DFFSR_151 ( );
FILL FILL_38_DFFSR_151 ( );
FILL FILL_39_DFFSR_151 ( );
FILL FILL_40_DFFSR_151 ( );
FILL FILL_41_DFFSR_151 ( );
FILL FILL_42_DFFSR_151 ( );
FILL FILL_43_DFFSR_151 ( );
FILL FILL_44_DFFSR_151 ( );
FILL FILL_45_DFFSR_151 ( );
FILL FILL_46_DFFSR_151 ( );
FILL FILL_47_DFFSR_151 ( );
FILL FILL_48_DFFSR_151 ( );
FILL FILL_49_DFFSR_151 ( );
FILL FILL_50_DFFSR_151 ( );
FILL FILL_0_BUFX2_10 ( );
FILL FILL_1_BUFX2_10 ( );
FILL FILL_2_BUFX2_10 ( );
FILL FILL_3_BUFX2_10 ( );
FILL FILL_4_BUFX2_10 ( );
FILL FILL_5_BUFX2_10 ( );
FILL FILL_6_BUFX2_10 ( );
FILL FILL_0_OAI21X1_133 ( );
FILL FILL_1_OAI21X1_133 ( );
FILL FILL_2_OAI21X1_133 ( );
FILL FILL_3_OAI21X1_133 ( );
FILL FILL_4_OAI21X1_133 ( );
FILL FILL_5_OAI21X1_133 ( );
FILL FILL_6_OAI21X1_133 ( );
FILL FILL_7_OAI21X1_133 ( );
FILL FILL_8_OAI21X1_133 ( );
FILL FILL_9_OAI21X1_133 ( );
FILL FILL_0_BUFX2_7 ( );
FILL FILL_1_BUFX2_7 ( );
FILL FILL_2_BUFX2_7 ( );
FILL FILL_3_BUFX2_7 ( );
FILL FILL_4_BUFX2_7 ( );
FILL FILL_5_BUFX2_7 ( );
FILL FILL_6_BUFX2_7 ( );
FILL FILL_0_INVX1_10 ( );
FILL FILL_1_INVX1_10 ( );
FILL FILL_2_INVX1_10 ( );
FILL FILL_3_INVX1_10 ( );
FILL FILL_0_NOR2X1_2 ( );
FILL FILL_1_NOR2X1_2 ( );
FILL FILL_2_NOR2X1_2 ( );
FILL FILL_3_NOR2X1_2 ( );
FILL FILL_4_NOR2X1_2 ( );
FILL FILL_5_NOR2X1_2 ( );
FILL FILL_6_NOR2X1_2 ( );
FILL FILL_0_DFFSR_54 ( );
FILL FILL_1_DFFSR_54 ( );
FILL FILL_2_DFFSR_54 ( );
FILL FILL_3_DFFSR_54 ( );
FILL FILL_4_DFFSR_54 ( );
FILL FILL_5_DFFSR_54 ( );
FILL FILL_6_DFFSR_54 ( );
FILL FILL_7_DFFSR_54 ( );
FILL FILL_8_DFFSR_54 ( );
FILL FILL_9_DFFSR_54 ( );
FILL FILL_10_DFFSR_54 ( );
FILL FILL_11_DFFSR_54 ( );
FILL FILL_12_DFFSR_54 ( );
FILL FILL_13_DFFSR_54 ( );
FILL FILL_14_DFFSR_54 ( );
FILL FILL_15_DFFSR_54 ( );
FILL FILL_16_DFFSR_54 ( );
FILL FILL_17_DFFSR_54 ( );
FILL FILL_18_DFFSR_54 ( );
FILL FILL_19_DFFSR_54 ( );
FILL FILL_20_DFFSR_54 ( );
FILL FILL_21_DFFSR_54 ( );
FILL FILL_22_DFFSR_54 ( );
FILL FILL_23_DFFSR_54 ( );
FILL FILL_24_DFFSR_54 ( );
FILL FILL_25_DFFSR_54 ( );
FILL FILL_26_DFFSR_54 ( );
FILL FILL_27_DFFSR_54 ( );
FILL FILL_28_DFFSR_54 ( );
FILL FILL_29_DFFSR_54 ( );
FILL FILL_30_DFFSR_54 ( );
FILL FILL_31_DFFSR_54 ( );
FILL FILL_32_DFFSR_54 ( );
FILL FILL_33_DFFSR_54 ( );
FILL FILL_34_DFFSR_54 ( );
FILL FILL_35_DFFSR_54 ( );
FILL FILL_36_DFFSR_54 ( );
FILL FILL_37_DFFSR_54 ( );
FILL FILL_38_DFFSR_54 ( );
FILL FILL_39_DFFSR_54 ( );
FILL FILL_40_DFFSR_54 ( );
FILL FILL_41_DFFSR_54 ( );
FILL FILL_42_DFFSR_54 ( );
FILL FILL_43_DFFSR_54 ( );
FILL FILL_44_DFFSR_54 ( );
FILL FILL_45_DFFSR_54 ( );
FILL FILL_46_DFFSR_54 ( );
FILL FILL_47_DFFSR_54 ( );
FILL FILL_48_DFFSR_54 ( );
FILL FILL_49_DFFSR_54 ( );
FILL FILL_50_DFFSR_54 ( );
FILL FILL_0_INVX1_64 ( );
FILL FILL_1_INVX1_64 ( );
FILL FILL_2_INVX1_64 ( );
FILL FILL_3_INVX1_64 ( );
FILL FILL_4_INVX1_64 ( );
FILL FILL_0_OAI21X1_28 ( );
FILL FILL_1_OAI21X1_28 ( );
FILL FILL_2_OAI21X1_28 ( );
FILL FILL_3_OAI21X1_28 ( );
FILL FILL_4_OAI21X1_28 ( );
FILL FILL_5_OAI21X1_28 ( );
FILL FILL_6_OAI21X1_28 ( );
FILL FILL_7_OAI21X1_28 ( );
FILL FILL_8_OAI21X1_28 ( );
FILL FILL_0_NAND2X1_28 ( );
FILL FILL_1_NAND2X1_28 ( );
FILL FILL_2_NAND2X1_28 ( );
FILL FILL_3_NAND2X1_28 ( );
FILL FILL_4_NAND2X1_28 ( );
FILL FILL_5_NAND2X1_28 ( );
FILL FILL_6_NAND2X1_28 ( );
FILL FILL_0_DFFSR_170 ( );
FILL FILL_1_DFFSR_170 ( );
FILL FILL_2_DFFSR_170 ( );
FILL FILL_3_DFFSR_170 ( );
FILL FILL_4_DFFSR_170 ( );
FILL FILL_5_DFFSR_170 ( );
FILL FILL_6_DFFSR_170 ( );
FILL FILL_7_DFFSR_170 ( );
FILL FILL_8_DFFSR_170 ( );
FILL FILL_9_DFFSR_170 ( );
FILL FILL_10_DFFSR_170 ( );
FILL FILL_11_DFFSR_170 ( );
FILL FILL_12_DFFSR_170 ( );
FILL FILL_13_DFFSR_170 ( );
FILL FILL_14_DFFSR_170 ( );
FILL FILL_15_DFFSR_170 ( );
FILL FILL_16_DFFSR_170 ( );
FILL FILL_17_DFFSR_170 ( );
FILL FILL_18_DFFSR_170 ( );
FILL FILL_19_DFFSR_170 ( );
FILL FILL_20_DFFSR_170 ( );
FILL FILL_21_DFFSR_170 ( );
FILL FILL_22_DFFSR_170 ( );
FILL FILL_23_DFFSR_170 ( );
FILL FILL_24_DFFSR_170 ( );
FILL FILL_25_DFFSR_170 ( );
FILL FILL_26_DFFSR_170 ( );
FILL FILL_27_DFFSR_170 ( );
FILL FILL_28_DFFSR_170 ( );
FILL FILL_29_DFFSR_170 ( );
FILL FILL_30_DFFSR_170 ( );
FILL FILL_31_DFFSR_170 ( );
FILL FILL_32_DFFSR_170 ( );
FILL FILL_33_DFFSR_170 ( );
FILL FILL_34_DFFSR_170 ( );
FILL FILL_35_DFFSR_170 ( );
FILL FILL_36_DFFSR_170 ( );
FILL FILL_37_DFFSR_170 ( );
FILL FILL_38_DFFSR_170 ( );
FILL FILL_39_DFFSR_170 ( );
FILL FILL_40_DFFSR_170 ( );
FILL FILL_41_DFFSR_170 ( );
FILL FILL_42_DFFSR_170 ( );
FILL FILL_43_DFFSR_170 ( );
FILL FILL_44_DFFSR_170 ( );
FILL FILL_45_DFFSR_170 ( );
FILL FILL_46_DFFSR_170 ( );
FILL FILL_47_DFFSR_170 ( );
FILL FILL_48_DFFSR_170 ( );
FILL FILL_49_DFFSR_170 ( );
FILL FILL_50_DFFSR_170 ( );
FILL FILL_0_NAND2X1_193 ( );
FILL FILL_1_NAND2X1_193 ( );
FILL FILL_2_NAND2X1_193 ( );
FILL FILL_3_NAND2X1_193 ( );
FILL FILL_4_NAND2X1_193 ( );
FILL FILL_5_NAND2X1_193 ( );
FILL FILL_6_NAND2X1_193 ( );
FILL FILL_0_NAND3X1_21 ( );
FILL FILL_1_NAND3X1_21 ( );
FILL FILL_2_NAND3X1_21 ( );
FILL FILL_3_NAND3X1_21 ( );
FILL FILL_4_NAND3X1_21 ( );
FILL FILL_5_NAND3X1_21 ( );
FILL FILL_6_NAND3X1_21 ( );
FILL FILL_7_NAND3X1_21 ( );
FILL FILL_8_NAND3X1_21 ( );
FILL FILL_9_NAND3X1_21 ( );
FILL FILL_0_NAND2X1_195 ( );
FILL FILL_1_NAND2X1_195 ( );
FILL FILL_2_NAND2X1_195 ( );
FILL FILL_3_NAND2X1_195 ( );
FILL FILL_4_NAND2X1_195 ( );
FILL FILL_5_NAND2X1_195 ( );
FILL FILL_6_NAND2X1_195 ( );
FILL FILL_0_NAND3X1_25 ( );
FILL FILL_1_NAND3X1_25 ( );
FILL FILL_2_NAND3X1_25 ( );
FILL FILL_3_NAND3X1_25 ( );
FILL FILL_4_NAND3X1_25 ( );
FILL FILL_5_NAND3X1_25 ( );
FILL FILL_6_NAND3X1_25 ( );
FILL FILL_7_NAND3X1_25 ( );
FILL FILL_8_NAND3X1_25 ( );
FILL FILL_0_NAND3X1_26 ( );
FILL FILL_1_NAND3X1_26 ( );
FILL FILL_2_NAND3X1_26 ( );
FILL FILL_3_NAND3X1_26 ( );
FILL FILL_4_NAND3X1_26 ( );
FILL FILL_5_NAND3X1_26 ( );
FILL FILL_6_NAND3X1_26 ( );
FILL FILL_7_NAND3X1_26 ( );
FILL FILL_8_NAND3X1_26 ( );
FILL FILL_0_AOI21X1_4 ( );
FILL FILL_1_AOI21X1_4 ( );
FILL FILL_2_AOI21X1_4 ( );
FILL FILL_3_AOI21X1_4 ( );
FILL FILL_4_AOI21X1_4 ( );
FILL FILL_5_AOI21X1_4 ( );
FILL FILL_6_AOI21X1_4 ( );
FILL FILL_7_AOI21X1_4 ( );
FILL FILL_8_AOI21X1_4 ( );
FILL FILL_9_AOI21X1_4 ( );
FILL FILL_0_OAI21X1_195 ( );
FILL FILL_1_OAI21X1_195 ( );
FILL FILL_2_OAI21X1_195 ( );
FILL FILL_3_OAI21X1_195 ( );
FILL FILL_4_OAI21X1_195 ( );
FILL FILL_5_OAI21X1_195 ( );
FILL FILL_6_OAI21X1_195 ( );
FILL FILL_7_OAI21X1_195 ( );
FILL FILL_8_OAI21X1_195 ( );
FILL FILL_0_AOI21X1_14 ( );
FILL FILL_1_AOI21X1_14 ( );
FILL FILL_2_AOI21X1_14 ( );
FILL FILL_3_AOI21X1_14 ( );
FILL FILL_4_AOI21X1_14 ( );
FILL FILL_5_AOI21X1_14 ( );
FILL FILL_6_AOI21X1_14 ( );
FILL FILL_7_AOI21X1_14 ( );
FILL FILL_8_AOI21X1_14 ( );
FILL FILL_0_NAND3X1_28 ( );
FILL FILL_1_NAND3X1_28 ( );
FILL FILL_2_NAND3X1_28 ( );
FILL FILL_3_NAND3X1_28 ( );
FILL FILL_4_NAND3X1_28 ( );
FILL FILL_5_NAND3X1_28 ( );
FILL FILL_6_NAND3X1_28 ( );
FILL FILL_7_NAND3X1_28 ( );
FILL FILL_8_NAND3X1_28 ( );
FILL FILL_0_AOI21X1_20 ( );
FILL FILL_1_AOI21X1_20 ( );
FILL FILL_2_AOI21X1_20 ( );
FILL FILL_3_AOI21X1_20 ( );
FILL FILL_4_AOI21X1_20 ( );
FILL FILL_5_AOI21X1_20 ( );
FILL FILL_6_AOI21X1_20 ( );
FILL FILL_7_AOI21X1_20 ( );
FILL FILL_8_AOI21X1_20 ( );
FILL FILL_0_NAND3X1_56 ( );
FILL FILL_1_NAND3X1_56 ( );
FILL FILL_2_NAND3X1_56 ( );
FILL FILL_3_NAND3X1_56 ( );
FILL FILL_4_NAND3X1_56 ( );
FILL FILL_5_NAND3X1_56 ( );
FILL FILL_6_NAND3X1_56 ( );
FILL FILL_7_NAND3X1_56 ( );
FILL FILL_8_NAND3X1_56 ( );
FILL FILL_0_NAND3X1_51 ( );
FILL FILL_1_NAND3X1_51 ( );
FILL FILL_2_NAND3X1_51 ( );
FILL FILL_3_NAND3X1_51 ( );
FILL FILL_4_NAND3X1_51 ( );
FILL FILL_5_NAND3X1_51 ( );
FILL FILL_6_NAND3X1_51 ( );
FILL FILL_7_NAND3X1_51 ( );
FILL FILL_8_NAND3X1_51 ( );
FILL FILL_9_NAND3X1_51 ( );
FILL FILL_0_NAND3X1_82 ( );
FILL FILL_1_NAND3X1_82 ( );
FILL FILL_2_NAND3X1_82 ( );
FILL FILL_3_NAND3X1_82 ( );
FILL FILL_4_NAND3X1_82 ( );
FILL FILL_5_NAND3X1_82 ( );
FILL FILL_6_NAND3X1_82 ( );
FILL FILL_7_NAND3X1_82 ( );
FILL FILL_8_NAND3X1_82 ( );
FILL FILL_9_NAND3X1_82 ( );
FILL FILL_0_NAND2X1_233 ( );
FILL FILL_1_NAND2X1_233 ( );
FILL FILL_2_NAND2X1_233 ( );
FILL FILL_3_NAND2X1_233 ( );
FILL FILL_4_NAND2X1_233 ( );
FILL FILL_5_NAND2X1_233 ( );
FILL FILL_6_NAND2X1_233 ( );
FILL FILL_0_AOI21X1_39 ( );
FILL FILL_1_AOI21X1_39 ( );
FILL FILL_2_AOI21X1_39 ( );
FILL FILL_3_AOI21X1_39 ( );
FILL FILL_4_AOI21X1_39 ( );
FILL FILL_5_AOI21X1_39 ( );
FILL FILL_6_AOI21X1_39 ( );
FILL FILL_7_AOI21X1_39 ( );
FILL FILL_8_AOI21X1_39 ( );
FILL FILL_9_AOI21X1_39 ( );
FILL FILL_0_DFFSR_76 ( );
FILL FILL_1_DFFSR_76 ( );
FILL FILL_2_DFFSR_76 ( );
FILL FILL_3_DFFSR_76 ( );
FILL FILL_4_DFFSR_76 ( );
FILL FILL_5_DFFSR_76 ( );
FILL FILL_6_DFFSR_76 ( );
FILL FILL_7_DFFSR_76 ( );
FILL FILL_8_DFFSR_76 ( );
FILL FILL_9_DFFSR_76 ( );
FILL FILL_10_DFFSR_76 ( );
FILL FILL_11_DFFSR_76 ( );
FILL FILL_12_DFFSR_76 ( );
FILL FILL_13_DFFSR_76 ( );
FILL FILL_14_DFFSR_76 ( );
FILL FILL_15_DFFSR_76 ( );
FILL FILL_16_DFFSR_76 ( );
FILL FILL_17_DFFSR_76 ( );
FILL FILL_18_DFFSR_76 ( );
FILL FILL_19_DFFSR_76 ( );
FILL FILL_20_DFFSR_76 ( );
FILL FILL_21_DFFSR_76 ( );
FILL FILL_22_DFFSR_76 ( );
FILL FILL_23_DFFSR_76 ( );
FILL FILL_24_DFFSR_76 ( );
FILL FILL_25_DFFSR_76 ( );
FILL FILL_26_DFFSR_76 ( );
FILL FILL_27_DFFSR_76 ( );
FILL FILL_28_DFFSR_76 ( );
FILL FILL_29_DFFSR_76 ( );
FILL FILL_30_DFFSR_76 ( );
FILL FILL_31_DFFSR_76 ( );
FILL FILL_32_DFFSR_76 ( );
FILL FILL_33_DFFSR_76 ( );
FILL FILL_34_DFFSR_76 ( );
FILL FILL_35_DFFSR_76 ( );
FILL FILL_36_DFFSR_76 ( );
FILL FILL_37_DFFSR_76 ( );
FILL FILL_38_DFFSR_76 ( );
FILL FILL_39_DFFSR_76 ( );
FILL FILL_40_DFFSR_76 ( );
FILL FILL_41_DFFSR_76 ( );
FILL FILL_42_DFFSR_76 ( );
FILL FILL_43_DFFSR_76 ( );
FILL FILL_44_DFFSR_76 ( );
FILL FILL_45_DFFSR_76 ( );
FILL FILL_46_DFFSR_76 ( );
FILL FILL_47_DFFSR_76 ( );
FILL FILL_48_DFFSR_76 ( );
FILL FILL_49_DFFSR_76 ( );
FILL FILL_50_DFFSR_76 ( );
FILL FILL_0_NAND2X1_108 ( );
FILL FILL_1_NAND2X1_108 ( );
FILL FILL_2_NAND2X1_108 ( );
FILL FILL_3_NAND2X1_108 ( );
FILL FILL_4_NAND2X1_108 ( );
FILL FILL_5_NAND2X1_108 ( );
FILL FILL_6_NAND2X1_108 ( );
FILL FILL_0_DFFSR_155 ( );
FILL FILL_1_DFFSR_155 ( );
FILL FILL_2_DFFSR_155 ( );
FILL FILL_3_DFFSR_155 ( );
FILL FILL_4_DFFSR_155 ( );
FILL FILL_5_DFFSR_155 ( );
FILL FILL_6_DFFSR_155 ( );
FILL FILL_7_DFFSR_155 ( );
FILL FILL_8_DFFSR_155 ( );
FILL FILL_9_DFFSR_155 ( );
FILL FILL_10_DFFSR_155 ( );
FILL FILL_11_DFFSR_155 ( );
FILL FILL_12_DFFSR_155 ( );
FILL FILL_13_DFFSR_155 ( );
FILL FILL_14_DFFSR_155 ( );
FILL FILL_15_DFFSR_155 ( );
FILL FILL_16_DFFSR_155 ( );
FILL FILL_17_DFFSR_155 ( );
FILL FILL_18_DFFSR_155 ( );
FILL FILL_19_DFFSR_155 ( );
FILL FILL_20_DFFSR_155 ( );
FILL FILL_21_DFFSR_155 ( );
FILL FILL_22_DFFSR_155 ( );
FILL FILL_23_DFFSR_155 ( );
FILL FILL_24_DFFSR_155 ( );
FILL FILL_25_DFFSR_155 ( );
FILL FILL_26_DFFSR_155 ( );
FILL FILL_27_DFFSR_155 ( );
FILL FILL_28_DFFSR_155 ( );
FILL FILL_29_DFFSR_155 ( );
FILL FILL_30_DFFSR_155 ( );
FILL FILL_31_DFFSR_155 ( );
FILL FILL_32_DFFSR_155 ( );
FILL FILL_33_DFFSR_155 ( );
FILL FILL_34_DFFSR_155 ( );
FILL FILL_35_DFFSR_155 ( );
FILL FILL_36_DFFSR_155 ( );
FILL FILL_37_DFFSR_155 ( );
FILL FILL_38_DFFSR_155 ( );
FILL FILL_39_DFFSR_155 ( );
FILL FILL_40_DFFSR_155 ( );
FILL FILL_41_DFFSR_155 ( );
FILL FILL_42_DFFSR_155 ( );
FILL FILL_43_DFFSR_155 ( );
FILL FILL_44_DFFSR_155 ( );
FILL FILL_45_DFFSR_155 ( );
FILL FILL_46_DFFSR_155 ( );
FILL FILL_47_DFFSR_155 ( );
FILL FILL_48_DFFSR_155 ( );
FILL FILL_49_DFFSR_155 ( );
FILL FILL_50_DFFSR_155 ( );
FILL FILL_0_DFFSR_137 ( );
FILL FILL_1_DFFSR_137 ( );
FILL FILL_2_DFFSR_137 ( );
FILL FILL_3_DFFSR_137 ( );
FILL FILL_4_DFFSR_137 ( );
FILL FILL_5_DFFSR_137 ( );
FILL FILL_6_DFFSR_137 ( );
FILL FILL_7_DFFSR_137 ( );
FILL FILL_8_DFFSR_137 ( );
FILL FILL_9_DFFSR_137 ( );
FILL FILL_10_DFFSR_137 ( );
FILL FILL_11_DFFSR_137 ( );
FILL FILL_12_DFFSR_137 ( );
FILL FILL_13_DFFSR_137 ( );
FILL FILL_14_DFFSR_137 ( );
FILL FILL_15_DFFSR_137 ( );
FILL FILL_16_DFFSR_137 ( );
FILL FILL_17_DFFSR_137 ( );
FILL FILL_18_DFFSR_137 ( );
FILL FILL_19_DFFSR_137 ( );
FILL FILL_20_DFFSR_137 ( );
FILL FILL_21_DFFSR_137 ( );
FILL FILL_22_DFFSR_137 ( );
FILL FILL_23_DFFSR_137 ( );
FILL FILL_24_DFFSR_137 ( );
FILL FILL_25_DFFSR_137 ( );
FILL FILL_26_DFFSR_137 ( );
FILL FILL_27_DFFSR_137 ( );
FILL FILL_28_DFFSR_137 ( );
FILL FILL_29_DFFSR_137 ( );
FILL FILL_30_DFFSR_137 ( );
FILL FILL_31_DFFSR_137 ( );
FILL FILL_32_DFFSR_137 ( );
FILL FILL_33_DFFSR_137 ( );
FILL FILL_34_DFFSR_137 ( );
FILL FILL_35_DFFSR_137 ( );
FILL FILL_36_DFFSR_137 ( );
FILL FILL_37_DFFSR_137 ( );
FILL FILL_38_DFFSR_137 ( );
FILL FILL_39_DFFSR_137 ( );
FILL FILL_40_DFFSR_137 ( );
FILL FILL_41_DFFSR_137 ( );
FILL FILL_42_DFFSR_137 ( );
FILL FILL_43_DFFSR_137 ( );
FILL FILL_44_DFFSR_137 ( );
FILL FILL_45_DFFSR_137 ( );
FILL FILL_46_DFFSR_137 ( );
FILL FILL_47_DFFSR_137 ( );
FILL FILL_48_DFFSR_137 ( );
FILL FILL_49_DFFSR_137 ( );
FILL FILL_50_DFFSR_137 ( );
FILL FILL_0_INVX1_150 ( );
FILL FILL_1_INVX1_150 ( );
FILL FILL_2_INVX1_150 ( );
FILL FILL_3_INVX1_150 ( );
FILL FILL_0_CLKBUF1_11 ( );
FILL FILL_1_CLKBUF1_11 ( );
FILL FILL_2_CLKBUF1_11 ( );
FILL FILL_3_CLKBUF1_11 ( );
FILL FILL_4_CLKBUF1_11 ( );
FILL FILL_5_CLKBUF1_11 ( );
FILL FILL_6_CLKBUF1_11 ( );
FILL FILL_7_CLKBUF1_11 ( );
FILL FILL_8_CLKBUF1_11 ( );
FILL FILL_9_CLKBUF1_11 ( );
FILL FILL_10_CLKBUF1_11 ( );
FILL FILL_11_CLKBUF1_11 ( );
FILL FILL_12_CLKBUF1_11 ( );
FILL FILL_13_CLKBUF1_11 ( );
FILL FILL_14_CLKBUF1_11 ( );
FILL FILL_15_CLKBUF1_11 ( );
FILL FILL_16_CLKBUF1_11 ( );
FILL FILL_17_CLKBUF1_11 ( );
FILL FILL_18_CLKBUF1_11 ( );
FILL FILL_19_CLKBUF1_11 ( );
FILL FILL_20_CLKBUF1_11 ( );
FILL FILL_0_INVX1_61 ( );
FILL FILL_1_INVX1_61 ( );
FILL FILL_2_INVX1_61 ( );
FILL FILL_3_INVX1_61 ( );
FILL FILL_4_INVX1_61 ( );
FILL FILL_0_OAI21X1_54 ( );
FILL FILL_1_OAI21X1_54 ( );
FILL FILL_2_OAI21X1_54 ( );
FILL FILL_3_OAI21X1_54 ( );
FILL FILL_4_OAI21X1_54 ( );
FILL FILL_5_OAI21X1_54 ( );
FILL FILL_6_OAI21X1_54 ( );
FILL FILL_7_OAI21X1_54 ( );
FILL FILL_8_OAI21X1_54 ( );
FILL FILL_0_NAND2X1_54 ( );
FILL FILL_1_NAND2X1_54 ( );
FILL FILL_2_NAND2X1_54 ( );
FILL FILL_3_NAND2X1_54 ( );
FILL FILL_4_NAND2X1_54 ( );
FILL FILL_5_NAND2X1_54 ( );
FILL FILL_6_NAND2X1_54 ( );
FILL FILL_0_INVX1_308 ( );
FILL FILL_1_INVX1_308 ( );
FILL FILL_2_INVX1_308 ( );
FILL FILL_3_INVX1_308 ( );
FILL FILL_4_INVX1_308 ( );
FILL FILL_0_INVX1_295 ( );
FILL FILL_1_INVX1_295 ( );
FILL FILL_2_INVX1_295 ( );
FILL FILL_3_INVX1_295 ( );
FILL FILL_4_INVX1_295 ( );
FILL FILL_0_NAND2X1_252 ( );
FILL FILL_1_NAND2X1_252 ( );
FILL FILL_2_NAND2X1_252 ( );
FILL FILL_3_NAND2X1_252 ( );
FILL FILL_4_NAND2X1_252 ( );
FILL FILL_5_NAND2X1_252 ( );
FILL FILL_6_NAND2X1_252 ( );
FILL FILL_0_NAND2X1_253 ( );
FILL FILL_1_NAND2X1_253 ( );
FILL FILL_2_NAND2X1_253 ( );
FILL FILL_3_NAND2X1_253 ( );
FILL FILL_4_NAND2X1_253 ( );
FILL FILL_5_NAND2X1_253 ( );
FILL FILL_6_NAND2X1_253 ( );
FILL FILL_0_NAND3X1_131 ( );
FILL FILL_1_NAND3X1_131 ( );
FILL FILL_2_NAND3X1_131 ( );
FILL FILL_3_NAND3X1_131 ( );
FILL FILL_4_NAND3X1_131 ( );
FILL FILL_5_NAND3X1_131 ( );
FILL FILL_6_NAND3X1_131 ( );
FILL FILL_7_NAND3X1_131 ( );
FILL FILL_8_NAND3X1_131 ( );
FILL FILL_9_NAND3X1_131 ( );
FILL FILL_0_INVX1_32 ( );
FILL FILL_1_INVX1_32 ( );
FILL FILL_2_INVX1_32 ( );
FILL FILL_3_INVX1_32 ( );
FILL FILL_4_INVX1_32 ( );
FILL FILL_0_NAND2X1_60 ( );
FILL FILL_1_NAND2X1_60 ( );
FILL FILL_2_NAND2X1_60 ( );
FILL FILL_3_NAND2X1_60 ( );
FILL FILL_4_NAND2X1_60 ( );
FILL FILL_5_NAND2X1_60 ( );
FILL FILL_6_NAND2X1_60 ( );
FILL FILL_0_INVX1_405 ( );
FILL FILL_1_INVX1_405 ( );
FILL FILL_2_INVX1_405 ( );
FILL FILL_3_INVX1_405 ( );
FILL FILL_0_DFFPOSX1_20 ( );
FILL FILL_1_DFFPOSX1_20 ( );
FILL FILL_2_DFFPOSX1_20 ( );
FILL FILL_3_DFFPOSX1_20 ( );
FILL FILL_4_DFFPOSX1_20 ( );
FILL FILL_5_DFFPOSX1_20 ( );
FILL FILL_6_DFFPOSX1_20 ( );
FILL FILL_7_DFFPOSX1_20 ( );
FILL FILL_8_DFFPOSX1_20 ( );
FILL FILL_9_DFFPOSX1_20 ( );
FILL FILL_10_DFFPOSX1_20 ( );
FILL FILL_11_DFFPOSX1_20 ( );
FILL FILL_12_DFFPOSX1_20 ( );
FILL FILL_13_DFFPOSX1_20 ( );
FILL FILL_14_DFFPOSX1_20 ( );
FILL FILL_15_DFFPOSX1_20 ( );
FILL FILL_16_DFFPOSX1_20 ( );
FILL FILL_17_DFFPOSX1_20 ( );
FILL FILL_18_DFFPOSX1_20 ( );
FILL FILL_19_DFFPOSX1_20 ( );
FILL FILL_20_DFFPOSX1_20 ( );
FILL FILL_21_DFFPOSX1_20 ( );
FILL FILL_22_DFFPOSX1_20 ( );
FILL FILL_23_DFFPOSX1_20 ( );
FILL FILL_24_DFFPOSX1_20 ( );
FILL FILL_25_DFFPOSX1_20 ( );
FILL FILL_26_DFFPOSX1_20 ( );
FILL FILL_27_DFFPOSX1_20 ( );
FILL FILL_0_BUFX2_11 ( );
FILL FILL_1_BUFX2_11 ( );
FILL FILL_2_BUFX2_11 ( );
FILL FILL_3_BUFX2_11 ( );
FILL FILL_4_BUFX2_11 ( );
FILL FILL_5_BUFX2_11 ( );
FILL FILL_6_BUFX2_11 ( );
FILL FILL_0_BUFX2_13 ( );
FILL FILL_1_BUFX2_13 ( );
FILL FILL_2_BUFX2_13 ( );
FILL FILL_3_BUFX2_13 ( );
FILL FILL_4_BUFX2_13 ( );
FILL FILL_5_BUFX2_13 ( );
FILL FILL_6_BUFX2_13 ( );
FILL FILL_0_AND2X2_2 ( );
FILL FILL_1_AND2X2_2 ( );
FILL FILL_2_AND2X2_2 ( );
FILL FILL_3_AND2X2_2 ( );
FILL FILL_4_AND2X2_2 ( );
FILL FILL_5_AND2X2_2 ( );
FILL FILL_6_AND2X2_2 ( );
FILL FILL_7_AND2X2_2 ( );
FILL FILL_8_AND2X2_2 ( );
FILL FILL_9_AND2X2_2 ( );
FILL FILL_0_AND2X2_7 ( );
FILL FILL_1_AND2X2_7 ( );
FILL FILL_2_AND2X2_7 ( );
FILL FILL_3_AND2X2_7 ( );
FILL FILL_4_AND2X2_7 ( );
FILL FILL_5_AND2X2_7 ( );
FILL FILL_6_AND2X2_7 ( );
FILL FILL_7_AND2X2_7 ( );
FILL FILL_8_AND2X2_7 ( );
FILL FILL_0_NAND2X1_194 ( );
FILL FILL_1_NAND2X1_194 ( );
FILL FILL_2_NAND2X1_194 ( );
FILL FILL_3_NAND2X1_194 ( );
FILL FILL_4_NAND2X1_194 ( );
FILL FILL_5_NAND2X1_194 ( );
FILL FILL_6_NAND2X1_194 ( );
FILL FILL_0_NAND2X1_196 ( );
FILL FILL_1_NAND2X1_196 ( );
FILL FILL_2_NAND2X1_196 ( );
FILL FILL_3_NAND2X1_196 ( );
FILL FILL_4_NAND2X1_196 ( );
FILL FILL_5_NAND2X1_196 ( );
FILL FILL_6_NAND2X1_196 ( );
FILL FILL_0_AOI22X1_3 ( );
FILL FILL_1_AOI22X1_3 ( );
FILL FILL_2_AOI22X1_3 ( );
FILL FILL_3_AOI22X1_3 ( );
FILL FILL_4_AOI22X1_3 ( );
FILL FILL_5_AOI22X1_3 ( );
FILL FILL_6_AOI22X1_3 ( );
FILL FILL_7_AOI22X1_3 ( );
FILL FILL_8_AOI22X1_3 ( );
FILL FILL_9_AOI22X1_3 ( );
FILL FILL_10_AOI22X1_3 ( );
FILL FILL_0_NAND3X1_7 ( );
FILL FILL_1_NAND3X1_7 ( );
FILL FILL_2_NAND3X1_7 ( );
FILL FILL_3_NAND3X1_7 ( );
FILL FILL_4_NAND3X1_7 ( );
FILL FILL_5_NAND3X1_7 ( );
FILL FILL_6_NAND3X1_7 ( );
FILL FILL_7_NAND3X1_7 ( );
FILL FILL_8_NAND3X1_7 ( );
FILL FILL_9_NAND3X1_7 ( );
FILL FILL_0_NAND3X1_10 ( );
FILL FILL_1_NAND3X1_10 ( );
FILL FILL_2_NAND3X1_10 ( );
FILL FILL_3_NAND3X1_10 ( );
FILL FILL_4_NAND3X1_10 ( );
FILL FILL_5_NAND3X1_10 ( );
FILL FILL_6_NAND3X1_10 ( );
FILL FILL_7_NAND3X1_10 ( );
FILL FILL_8_NAND3X1_10 ( );
FILL FILL_0_INVX1_233 ( );
FILL FILL_1_INVX1_233 ( );
FILL FILL_2_INVX1_233 ( );
FILL FILL_3_INVX1_233 ( );
FILL FILL_0_OAI21X1_193 ( );
FILL FILL_1_OAI21X1_193 ( );
FILL FILL_2_OAI21X1_193 ( );
FILL FILL_3_OAI21X1_193 ( );
FILL FILL_4_OAI21X1_193 ( );
FILL FILL_5_OAI21X1_193 ( );
FILL FILL_6_OAI21X1_193 ( );
FILL FILL_7_OAI21X1_193 ( );
FILL FILL_8_OAI21X1_193 ( );
FILL FILL_0_INVX1_224 ( );
FILL FILL_1_INVX1_224 ( );
FILL FILL_2_INVX1_224 ( );
FILL FILL_3_INVX1_224 ( );
FILL FILL_4_INVX1_224 ( );
FILL FILL_0_NAND3X1_29 ( );
FILL FILL_1_NAND3X1_29 ( );
FILL FILL_2_NAND3X1_29 ( );
FILL FILL_3_NAND3X1_29 ( );
FILL FILL_4_NAND3X1_29 ( );
FILL FILL_5_NAND3X1_29 ( );
FILL FILL_6_NAND3X1_29 ( );
FILL FILL_7_NAND3X1_29 ( );
FILL FILL_8_NAND3X1_29 ( );
FILL FILL_0_NAND3X1_54 ( );
FILL FILL_1_NAND3X1_54 ( );
FILL FILL_2_NAND3X1_54 ( );
FILL FILL_3_NAND3X1_54 ( );
FILL FILL_4_NAND3X1_54 ( );
FILL FILL_5_NAND3X1_54 ( );
FILL FILL_6_NAND3X1_54 ( );
FILL FILL_7_NAND3X1_54 ( );
FILL FILL_8_NAND3X1_54 ( );
FILL FILL_9_NAND3X1_54 ( );
FILL FILL_0_NAND3X1_55 ( );
FILL FILL_1_NAND3X1_55 ( );
FILL FILL_2_NAND3X1_55 ( );
FILL FILL_3_NAND3X1_55 ( );
FILL FILL_4_NAND3X1_55 ( );
FILL FILL_5_NAND3X1_55 ( );
FILL FILL_6_NAND3X1_55 ( );
FILL FILL_7_NAND3X1_55 ( );
FILL FILL_8_NAND3X1_55 ( );
FILL FILL_0_NAND3X1_80 ( );
FILL FILL_1_NAND3X1_80 ( );
FILL FILL_2_NAND3X1_80 ( );
FILL FILL_3_NAND3X1_80 ( );
FILL FILL_4_NAND3X1_80 ( );
FILL FILL_5_NAND3X1_80 ( );
FILL FILL_6_NAND3X1_80 ( );
FILL FILL_7_NAND3X1_80 ( );
FILL FILL_8_NAND3X1_80 ( );
FILL FILL_0_NAND3X1_110 ( );
FILL FILL_1_NAND3X1_110 ( );
FILL FILL_2_NAND3X1_110 ( );
FILL FILL_3_NAND3X1_110 ( );
FILL FILL_4_NAND3X1_110 ( );
FILL FILL_5_NAND3X1_110 ( );
FILL FILL_6_NAND3X1_110 ( );
FILL FILL_7_NAND3X1_110 ( );
FILL FILL_8_NAND3X1_110 ( );
FILL FILL_0_NAND2X1_232 ( );
FILL FILL_1_NAND2X1_232 ( );
FILL FILL_2_NAND2X1_232 ( );
FILL FILL_3_NAND2X1_232 ( );
FILL FILL_4_NAND2X1_232 ( );
FILL FILL_5_NAND2X1_232 ( );
FILL FILL_6_NAND2X1_232 ( );
FILL FILL_0_OAI22X1_4 ( );
FILL FILL_1_OAI22X1_4 ( );
FILL FILL_2_OAI22X1_4 ( );
FILL FILL_3_OAI22X1_4 ( );
FILL FILL_4_OAI22X1_4 ( );
FILL FILL_5_OAI22X1_4 ( );
FILL FILL_6_OAI22X1_4 ( );
FILL FILL_7_OAI22X1_4 ( );
FILL FILL_8_OAI22X1_4 ( );
FILL FILL_9_OAI22X1_4 ( );
FILL FILL_10_OAI22X1_4 ( );
FILL FILL_11_OAI22X1_4 ( );
FILL FILL_0_BUFX2_19 ( );
FILL FILL_1_BUFX2_19 ( );
FILL FILL_2_BUFX2_19 ( );
FILL FILL_3_BUFX2_19 ( );
FILL FILL_4_BUFX2_19 ( );
FILL FILL_5_BUFX2_19 ( );
FILL FILL_6_BUFX2_19 ( );
FILL FILL_0_OAI21X1_81 ( );
FILL FILL_1_OAI21X1_81 ( );
FILL FILL_2_OAI21X1_81 ( );
FILL FILL_3_OAI21X1_81 ( );
FILL FILL_4_OAI21X1_81 ( );
FILL FILL_5_OAI21X1_81 ( );
FILL FILL_6_OAI21X1_81 ( );
FILL FILL_7_OAI21X1_81 ( );
FILL FILL_8_OAI21X1_81 ( );
FILL FILL_9_OAI21X1_81 ( );
FILL FILL_0_INVX1_92 ( );
FILL FILL_1_INVX1_92 ( );
FILL FILL_2_INVX1_92 ( );
FILL FILL_3_INVX1_92 ( );
FILL FILL_0_OAI21X1_76 ( );
FILL FILL_1_OAI21X1_76 ( );
FILL FILL_2_OAI21X1_76 ( );
FILL FILL_3_OAI21X1_76 ( );
FILL FILL_4_OAI21X1_76 ( );
FILL FILL_5_OAI21X1_76 ( );
FILL FILL_6_OAI21X1_76 ( );
FILL FILL_7_OAI21X1_76 ( );
FILL FILL_8_OAI21X1_76 ( );
FILL FILL_0_INVX1_382 ( );
FILL FILL_1_INVX1_382 ( );
FILL FILL_2_INVX1_382 ( );
FILL FILL_3_INVX1_382 ( );
FILL FILL_4_INVX1_382 ( );
FILL FILL_0_INVX1_335 ( );
FILL FILL_1_INVX1_335 ( );
FILL FILL_2_INVX1_335 ( );
FILL FILL_3_INVX1_335 ( );
FILL FILL_0_DFFSR_83 ( );
FILL FILL_1_DFFSR_83 ( );
FILL FILL_2_DFFSR_83 ( );
FILL FILL_3_DFFSR_83 ( );
FILL FILL_4_DFFSR_83 ( );
FILL FILL_5_DFFSR_83 ( );
FILL FILL_6_DFFSR_83 ( );
FILL FILL_7_DFFSR_83 ( );
FILL FILL_8_DFFSR_83 ( );
FILL FILL_9_DFFSR_83 ( );
FILL FILL_10_DFFSR_83 ( );
FILL FILL_11_DFFSR_83 ( );
FILL FILL_12_DFFSR_83 ( );
FILL FILL_13_DFFSR_83 ( );
FILL FILL_14_DFFSR_83 ( );
FILL FILL_15_DFFSR_83 ( );
FILL FILL_16_DFFSR_83 ( );
FILL FILL_17_DFFSR_83 ( );
FILL FILL_18_DFFSR_83 ( );
FILL FILL_19_DFFSR_83 ( );
FILL FILL_20_DFFSR_83 ( );
FILL FILL_21_DFFSR_83 ( );
FILL FILL_22_DFFSR_83 ( );
FILL FILL_23_DFFSR_83 ( );
FILL FILL_24_DFFSR_83 ( );
FILL FILL_25_DFFSR_83 ( );
FILL FILL_26_DFFSR_83 ( );
FILL FILL_27_DFFSR_83 ( );
FILL FILL_28_DFFSR_83 ( );
FILL FILL_29_DFFSR_83 ( );
FILL FILL_30_DFFSR_83 ( );
FILL FILL_31_DFFSR_83 ( );
FILL FILL_32_DFFSR_83 ( );
FILL FILL_33_DFFSR_83 ( );
FILL FILL_34_DFFSR_83 ( );
FILL FILL_35_DFFSR_83 ( );
FILL FILL_36_DFFSR_83 ( );
FILL FILL_37_DFFSR_83 ( );
FILL FILL_38_DFFSR_83 ( );
FILL FILL_39_DFFSR_83 ( );
FILL FILL_40_DFFSR_83 ( );
FILL FILL_41_DFFSR_83 ( );
FILL FILL_42_DFFSR_83 ( );
FILL FILL_43_DFFSR_83 ( );
FILL FILL_44_DFFSR_83 ( );
FILL FILL_45_DFFSR_83 ( );
FILL FILL_46_DFFSR_83 ( );
FILL FILL_47_DFFSR_83 ( );
FILL FILL_48_DFFSR_83 ( );
FILL FILL_49_DFFSR_83 ( );
FILL FILL_50_DFFSR_83 ( );
FILL FILL_0_INVX1_351 ( );
FILL FILL_1_INVX1_351 ( );
FILL FILL_2_INVX1_351 ( );
FILL FILL_3_INVX1_351 ( );
FILL FILL_0_BUFX2_23 ( );
FILL FILL_1_BUFX2_23 ( );
FILL FILL_2_BUFX2_23 ( );
FILL FILL_3_BUFX2_23 ( );
FILL FILL_4_BUFX2_23 ( );
FILL FILL_5_BUFX2_23 ( );
FILL FILL_6_BUFX2_23 ( );
FILL FILL_0_NAND2X1_69 ( );
FILL FILL_1_NAND2X1_69 ( );
FILL FILL_2_NAND2X1_69 ( );
FILL FILL_3_NAND2X1_69 ( );
FILL FILL_4_NAND2X1_69 ( );
FILL FILL_5_NAND2X1_69 ( );
FILL FILL_6_NAND2X1_69 ( );
FILL FILL_0_DFFSR_142 ( );
FILL FILL_1_DFFSR_142 ( );
FILL FILL_2_DFFSR_142 ( );
FILL FILL_3_DFFSR_142 ( );
FILL FILL_4_DFFSR_142 ( );
FILL FILL_5_DFFSR_142 ( );
FILL FILL_6_DFFSR_142 ( );
FILL FILL_7_DFFSR_142 ( );
FILL FILL_8_DFFSR_142 ( );
FILL FILL_9_DFFSR_142 ( );
FILL FILL_10_DFFSR_142 ( );
FILL FILL_11_DFFSR_142 ( );
FILL FILL_12_DFFSR_142 ( );
FILL FILL_13_DFFSR_142 ( );
FILL FILL_14_DFFSR_142 ( );
FILL FILL_15_DFFSR_142 ( );
FILL FILL_16_DFFSR_142 ( );
FILL FILL_17_DFFSR_142 ( );
FILL FILL_18_DFFSR_142 ( );
FILL FILL_19_DFFSR_142 ( );
FILL FILL_20_DFFSR_142 ( );
FILL FILL_21_DFFSR_142 ( );
FILL FILL_22_DFFSR_142 ( );
FILL FILL_23_DFFSR_142 ( );
FILL FILL_24_DFFSR_142 ( );
FILL FILL_25_DFFSR_142 ( );
FILL FILL_26_DFFSR_142 ( );
FILL FILL_27_DFFSR_142 ( );
FILL FILL_28_DFFSR_142 ( );
FILL FILL_29_DFFSR_142 ( );
FILL FILL_30_DFFSR_142 ( );
FILL FILL_31_DFFSR_142 ( );
FILL FILL_32_DFFSR_142 ( );
FILL FILL_33_DFFSR_142 ( );
FILL FILL_34_DFFSR_142 ( );
FILL FILL_35_DFFSR_142 ( );
FILL FILL_36_DFFSR_142 ( );
FILL FILL_37_DFFSR_142 ( );
FILL FILL_38_DFFSR_142 ( );
FILL FILL_39_DFFSR_142 ( );
FILL FILL_40_DFFSR_142 ( );
FILL FILL_41_DFFSR_142 ( );
FILL FILL_42_DFFSR_142 ( );
FILL FILL_43_DFFSR_142 ( );
FILL FILL_44_DFFSR_142 ( );
FILL FILL_45_DFFSR_142 ( );
FILL FILL_46_DFFSR_142 ( );
FILL FILL_47_DFFSR_142 ( );
FILL FILL_48_DFFSR_142 ( );
FILL FILL_49_DFFSR_142 ( );
FILL FILL_50_DFFSR_142 ( );
FILL FILL_51_DFFSR_142 ( );
FILL FILL_0_NAND2X1_133 ( );
FILL FILL_1_NAND2X1_133 ( );
FILL FILL_2_NAND2X1_133 ( );
FILL FILL_3_NAND2X1_133 ( );
FILL FILL_4_NAND2X1_133 ( );
FILL FILL_5_NAND2X1_133 ( );
FILL FILL_6_NAND2X1_133 ( );
FILL FILL_0_INVX1_28 ( );
FILL FILL_1_INVX1_28 ( );
FILL FILL_2_INVX1_28 ( );
FILL FILL_3_INVX1_28 ( );
FILL FILL_4_INVX1_28 ( );
FILL FILL_0_INVX1_73 ( );
FILL FILL_1_INVX1_73 ( );
FILL FILL_2_INVX1_73 ( );
FILL FILL_3_INVX1_73 ( );
FILL FILL_0_NAND2X1_62 ( );
FILL FILL_1_NAND2X1_62 ( );
FILL FILL_2_NAND2X1_62 ( );
FILL FILL_3_NAND2X1_62 ( );
FILL FILL_4_NAND2X1_62 ( );
FILL FILL_5_NAND2X1_62 ( );
FILL FILL_6_NAND2X1_62 ( );
FILL FILL_0_OAI21X1_62 ( );
FILL FILL_1_OAI21X1_62 ( );
FILL FILL_2_OAI21X1_62 ( );
FILL FILL_3_OAI21X1_62 ( );
FILL FILL_4_OAI21X1_62 ( );
FILL FILL_5_OAI21X1_62 ( );
FILL FILL_6_OAI21X1_62 ( );
FILL FILL_7_OAI21X1_62 ( );
FILL FILL_8_OAI21X1_62 ( );
FILL FILL_9_OAI21X1_62 ( );
FILL FILL_0_INVX1_70 ( );
FILL FILL_1_INVX1_70 ( );
FILL FILL_2_INVX1_70 ( );
FILL FILL_3_INVX1_70 ( );
FILL FILL_0_INVX1_307 ( );
FILL FILL_1_INVX1_307 ( );
FILL FILL_2_INVX1_307 ( );
FILL FILL_3_INVX1_307 ( );
FILL FILL_4_INVX1_307 ( );
FILL FILL_0_DFFSR_28 ( );
FILL FILL_1_DFFSR_28 ( );
FILL FILL_2_DFFSR_28 ( );
FILL FILL_3_DFFSR_28 ( );
FILL FILL_4_DFFSR_28 ( );
FILL FILL_5_DFFSR_28 ( );
FILL FILL_6_DFFSR_28 ( );
FILL FILL_7_DFFSR_28 ( );
FILL FILL_8_DFFSR_28 ( );
FILL FILL_9_DFFSR_28 ( );
FILL FILL_10_DFFSR_28 ( );
FILL FILL_11_DFFSR_28 ( );
FILL FILL_12_DFFSR_28 ( );
FILL FILL_13_DFFSR_28 ( );
FILL FILL_14_DFFSR_28 ( );
FILL FILL_15_DFFSR_28 ( );
FILL FILL_16_DFFSR_28 ( );
FILL FILL_17_DFFSR_28 ( );
FILL FILL_18_DFFSR_28 ( );
FILL FILL_19_DFFSR_28 ( );
FILL FILL_20_DFFSR_28 ( );
FILL FILL_21_DFFSR_28 ( );
FILL FILL_22_DFFSR_28 ( );
FILL FILL_23_DFFSR_28 ( );
FILL FILL_24_DFFSR_28 ( );
FILL FILL_25_DFFSR_28 ( );
FILL FILL_26_DFFSR_28 ( );
FILL FILL_27_DFFSR_28 ( );
FILL FILL_28_DFFSR_28 ( );
FILL FILL_29_DFFSR_28 ( );
FILL FILL_30_DFFSR_28 ( );
FILL FILL_31_DFFSR_28 ( );
FILL FILL_32_DFFSR_28 ( );
FILL FILL_33_DFFSR_28 ( );
FILL FILL_34_DFFSR_28 ( );
FILL FILL_35_DFFSR_28 ( );
FILL FILL_36_DFFSR_28 ( );
FILL FILL_37_DFFSR_28 ( );
FILL FILL_38_DFFSR_28 ( );
FILL FILL_39_DFFSR_28 ( );
FILL FILL_40_DFFSR_28 ( );
FILL FILL_41_DFFSR_28 ( );
FILL FILL_42_DFFSR_28 ( );
FILL FILL_43_DFFSR_28 ( );
FILL FILL_44_DFFSR_28 ( );
FILL FILL_45_DFFSR_28 ( );
FILL FILL_46_DFFSR_28 ( );
FILL FILL_47_DFFSR_28 ( );
FILL FILL_48_DFFSR_28 ( );
FILL FILL_49_DFFSR_28 ( );
FILL FILL_50_DFFSR_28 ( );
FILL FILL_0_DFFPOSX1_25 ( );
FILL FILL_1_DFFPOSX1_25 ( );
FILL FILL_2_DFFPOSX1_25 ( );
FILL FILL_3_DFFPOSX1_25 ( );
FILL FILL_4_DFFPOSX1_25 ( );
FILL FILL_5_DFFPOSX1_25 ( );
FILL FILL_6_DFFPOSX1_25 ( );
FILL FILL_7_DFFPOSX1_25 ( );
FILL FILL_8_DFFPOSX1_25 ( );
FILL FILL_9_DFFPOSX1_25 ( );
FILL FILL_10_DFFPOSX1_25 ( );
FILL FILL_11_DFFPOSX1_25 ( );
FILL FILL_12_DFFPOSX1_25 ( );
FILL FILL_13_DFFPOSX1_25 ( );
FILL FILL_14_DFFPOSX1_25 ( );
FILL FILL_15_DFFPOSX1_25 ( );
FILL FILL_16_DFFPOSX1_25 ( );
FILL FILL_17_DFFPOSX1_25 ( );
FILL FILL_18_DFFPOSX1_25 ( );
FILL FILL_19_DFFPOSX1_25 ( );
FILL FILL_20_DFFPOSX1_25 ( );
FILL FILL_21_DFFPOSX1_25 ( );
FILL FILL_22_DFFPOSX1_25 ( );
FILL FILL_23_DFFPOSX1_25 ( );
FILL FILL_24_DFFPOSX1_25 ( );
FILL FILL_25_DFFPOSX1_25 ( );
FILL FILL_26_DFFPOSX1_25 ( );
FILL FILL_27_DFFPOSX1_25 ( );
FILL FILL_0_NAND2X1_171 ( );
FILL FILL_1_NAND2X1_171 ( );
FILL FILL_2_NAND2X1_171 ( );
FILL FILL_3_NAND2X1_171 ( );
FILL FILL_4_NAND2X1_171 ( );
FILL FILL_5_NAND2X1_171 ( );
FILL FILL_6_NAND2X1_171 ( );
FILL FILL_0_OAI21X1_171 ( );
FILL FILL_1_OAI21X1_171 ( );
FILL FILL_2_OAI21X1_171 ( );
FILL FILL_3_OAI21X1_171 ( );
FILL FILL_4_OAI21X1_171 ( );
FILL FILL_5_OAI21X1_171 ( );
FILL FILL_6_OAI21X1_171 ( );
FILL FILL_7_OAI21X1_171 ( );
FILL FILL_8_OAI21X1_171 ( );
FILL FILL_9_OAI21X1_171 ( );
FILL FILL_0_INVX1_206 ( );
FILL FILL_1_INVX1_206 ( );
FILL FILL_2_INVX1_206 ( );
FILL FILL_3_INVX1_206 ( );
FILL FILL_0_AOI22X1_1 ( );
FILL FILL_1_AOI22X1_1 ( );
FILL FILL_2_AOI22X1_1 ( );
FILL FILL_3_AOI22X1_1 ( );
FILL FILL_4_AOI22X1_1 ( );
FILL FILL_5_AOI22X1_1 ( );
FILL FILL_6_AOI22X1_1 ( );
FILL FILL_7_AOI22X1_1 ( );
FILL FILL_8_AOI22X1_1 ( );
FILL FILL_9_AOI22X1_1 ( );
FILL FILL_10_AOI22X1_1 ( );
FILL FILL_11_AOI22X1_1 ( );
FILL FILL_0_AND2X2_4 ( );
FILL FILL_1_AND2X2_4 ( );
FILL FILL_2_AND2X2_4 ( );
FILL FILL_3_AND2X2_4 ( );
FILL FILL_4_AND2X2_4 ( );
FILL FILL_5_AND2X2_4 ( );
FILL FILL_6_AND2X2_4 ( );
FILL FILL_7_AND2X2_4 ( );
FILL FILL_8_AND2X2_4 ( );
FILL FILL_0_NAND3X1_3 ( );
FILL FILL_1_NAND3X1_3 ( );
FILL FILL_2_NAND3X1_3 ( );
FILL FILL_3_NAND3X1_3 ( );
FILL FILL_4_NAND3X1_3 ( );
FILL FILL_5_NAND3X1_3 ( );
FILL FILL_6_NAND3X1_3 ( );
FILL FILL_7_NAND3X1_3 ( );
FILL FILL_8_NAND3X1_3 ( );
FILL FILL_0_NAND3X1_11 ( );
FILL FILL_1_NAND3X1_11 ( );
FILL FILL_2_NAND3X1_11 ( );
FILL FILL_3_NAND3X1_11 ( );
FILL FILL_4_NAND3X1_11 ( );
FILL FILL_5_NAND3X1_11 ( );
FILL FILL_6_NAND3X1_11 ( );
FILL FILL_7_NAND3X1_11 ( );
FILL FILL_8_NAND3X1_11 ( );
FILL FILL_9_NAND3X1_11 ( );
FILL FILL_0_INVX1_225 ( );
FILL FILL_1_INVX1_225 ( );
FILL FILL_2_INVX1_225 ( );
FILL FILL_3_INVX1_225 ( );
FILL FILL_4_INVX1_225 ( );
FILL FILL_0_NAND3X1_8 ( );
FILL FILL_1_NAND3X1_8 ( );
FILL FILL_2_NAND3X1_8 ( );
FILL FILL_3_NAND3X1_8 ( );
FILL FILL_4_NAND3X1_8 ( );
FILL FILL_5_NAND3X1_8 ( );
FILL FILL_6_NAND3X1_8 ( );
FILL FILL_7_NAND3X1_8 ( );
FILL FILL_8_NAND3X1_8 ( );
FILL FILL_0_AOI21X1_6 ( );
FILL FILL_1_AOI21X1_6 ( );
FILL FILL_2_AOI21X1_6 ( );
FILL FILL_3_AOI21X1_6 ( );
FILL FILL_4_AOI21X1_6 ( );
FILL FILL_5_AOI21X1_6 ( );
FILL FILL_6_AOI21X1_6 ( );
FILL FILL_7_AOI21X1_6 ( );
FILL FILL_8_AOI21X1_6 ( );
FILL FILL_0_OAI21X1_194 ( );
FILL FILL_1_OAI21X1_194 ( );
FILL FILL_2_OAI21X1_194 ( );
FILL FILL_3_OAI21X1_194 ( );
FILL FILL_4_OAI21X1_194 ( );
FILL FILL_5_OAI21X1_194 ( );
FILL FILL_6_OAI21X1_194 ( );
FILL FILL_7_OAI21X1_194 ( );
FILL FILL_8_OAI21X1_194 ( );
FILL FILL_9_OAI21X1_194 ( );
FILL FILL_0_AOI21X1_7 ( );
FILL FILL_1_AOI21X1_7 ( );
FILL FILL_2_AOI21X1_7 ( );
FILL FILL_3_AOI21X1_7 ( );
FILL FILL_4_AOI21X1_7 ( );
FILL FILL_5_AOI21X1_7 ( );
FILL FILL_6_AOI21X1_7 ( );
FILL FILL_7_AOI21X1_7 ( );
FILL FILL_8_AOI21X1_7 ( );
FILL FILL_9_AOI21X1_7 ( );
FILL FILL_0_NAND3X1_57 ( );
FILL FILL_1_NAND3X1_57 ( );
FILL FILL_2_NAND3X1_57 ( );
FILL FILL_3_NAND3X1_57 ( );
FILL FILL_4_NAND3X1_57 ( );
FILL FILL_5_NAND3X1_57 ( );
FILL FILL_6_NAND3X1_57 ( );
FILL FILL_7_NAND3X1_57 ( );
FILL FILL_8_NAND3X1_57 ( );
FILL FILL_9_NAND3X1_57 ( );
FILL FILL_0_NAND3X1_58 ( );
FILL FILL_1_NAND3X1_58 ( );
FILL FILL_2_NAND3X1_58 ( );
FILL FILL_3_NAND3X1_58 ( );
FILL FILL_4_NAND3X1_58 ( );
FILL FILL_5_NAND3X1_58 ( );
FILL FILL_6_NAND3X1_58 ( );
FILL FILL_7_NAND3X1_58 ( );
FILL FILL_8_NAND3X1_58 ( );
FILL FILL_0_NAND3X1_78 ( );
FILL FILL_1_NAND3X1_78 ( );
FILL FILL_2_NAND3X1_78 ( );
FILL FILL_3_NAND3X1_78 ( );
FILL FILL_4_NAND3X1_78 ( );
FILL FILL_5_NAND3X1_78 ( );
FILL FILL_6_NAND3X1_78 ( );
FILL FILL_7_NAND3X1_78 ( );
FILL FILL_8_NAND3X1_78 ( );
FILL FILL_0_AOI21X1_19 ( );
FILL FILL_1_AOI21X1_19 ( );
FILL FILL_2_AOI21X1_19 ( );
FILL FILL_3_AOI21X1_19 ( );
FILL FILL_4_AOI21X1_19 ( );
FILL FILL_5_AOI21X1_19 ( );
FILL FILL_6_AOI21X1_19 ( );
FILL FILL_7_AOI21X1_19 ( );
FILL FILL_8_AOI21X1_19 ( );
FILL FILL_9_AOI21X1_19 ( );
FILL FILL_0_NAND2X1_219 ( );
FILL FILL_1_NAND2X1_219 ( );
FILL FILL_2_NAND2X1_219 ( );
FILL FILL_3_NAND2X1_219 ( );
FILL FILL_4_NAND2X1_219 ( );
FILL FILL_5_NAND2X1_219 ( );
FILL FILL_6_NAND2X1_219 ( );
FILL FILL_0_AND2X2_13 ( );
FILL FILL_1_AND2X2_13 ( );
FILL FILL_2_AND2X2_13 ( );
FILL FILL_3_AND2X2_13 ( );
FILL FILL_4_AND2X2_13 ( );
FILL FILL_5_AND2X2_13 ( );
FILL FILL_6_AND2X2_13 ( );
FILL FILL_7_AND2X2_13 ( );
FILL FILL_8_AND2X2_13 ( );
FILL FILL_0_DFFSR_128 ( );
FILL FILL_1_DFFSR_128 ( );
FILL FILL_2_DFFSR_128 ( );
FILL FILL_3_DFFSR_128 ( );
FILL FILL_4_DFFSR_128 ( );
FILL FILL_5_DFFSR_128 ( );
FILL FILL_6_DFFSR_128 ( );
FILL FILL_7_DFFSR_128 ( );
FILL FILL_8_DFFSR_128 ( );
FILL FILL_9_DFFSR_128 ( );
FILL FILL_10_DFFSR_128 ( );
FILL FILL_11_DFFSR_128 ( );
FILL FILL_12_DFFSR_128 ( );
FILL FILL_13_DFFSR_128 ( );
FILL FILL_14_DFFSR_128 ( );
FILL FILL_15_DFFSR_128 ( );
FILL FILL_16_DFFSR_128 ( );
FILL FILL_17_DFFSR_128 ( );
FILL FILL_18_DFFSR_128 ( );
FILL FILL_19_DFFSR_128 ( );
FILL FILL_20_DFFSR_128 ( );
FILL FILL_21_DFFSR_128 ( );
FILL FILL_22_DFFSR_128 ( );
FILL FILL_23_DFFSR_128 ( );
FILL FILL_24_DFFSR_128 ( );
FILL FILL_25_DFFSR_128 ( );
FILL FILL_26_DFFSR_128 ( );
FILL FILL_27_DFFSR_128 ( );
FILL FILL_28_DFFSR_128 ( );
FILL FILL_29_DFFSR_128 ( );
FILL FILL_30_DFFSR_128 ( );
FILL FILL_31_DFFSR_128 ( );
FILL FILL_32_DFFSR_128 ( );
FILL FILL_33_DFFSR_128 ( );
FILL FILL_34_DFFSR_128 ( );
FILL FILL_35_DFFSR_128 ( );
FILL FILL_36_DFFSR_128 ( );
FILL FILL_37_DFFSR_128 ( );
FILL FILL_38_DFFSR_128 ( );
FILL FILL_39_DFFSR_128 ( );
FILL FILL_40_DFFSR_128 ( );
FILL FILL_41_DFFSR_128 ( );
FILL FILL_42_DFFSR_128 ( );
FILL FILL_43_DFFSR_128 ( );
FILL FILL_44_DFFSR_128 ( );
FILL FILL_45_DFFSR_128 ( );
FILL FILL_46_DFFSR_128 ( );
FILL FILL_47_DFFSR_128 ( );
FILL FILL_48_DFFSR_128 ( );
FILL FILL_49_DFFSR_128 ( );
FILL FILL_50_DFFSR_128 ( );
FILL FILL_51_DFFSR_128 ( );
FILL FILL_0_INVX1_86 ( );
FILL FILL_1_INVX1_86 ( );
FILL FILL_2_INVX1_86 ( );
FILL FILL_3_INVX1_86 ( );
FILL FILL_4_INVX1_86 ( );
FILL FILL_0_INVX1_357 ( );
FILL FILL_1_INVX1_357 ( );
FILL FILL_2_INVX1_357 ( );
FILL FILL_3_INVX1_357 ( );
FILL FILL_0_OAI22X1_38 ( );
FILL FILL_1_OAI22X1_38 ( );
FILL FILL_2_OAI22X1_38 ( );
FILL FILL_3_OAI22X1_38 ( );
FILL FILL_4_OAI22X1_38 ( );
FILL FILL_5_OAI22X1_38 ( );
FILL FILL_6_OAI22X1_38 ( );
FILL FILL_7_OAI22X1_38 ( );
FILL FILL_8_OAI22X1_38 ( );
FILL FILL_9_OAI22X1_38 ( );
FILL FILL_10_OAI22X1_38 ( );
FILL FILL_11_OAI22X1_38 ( );
FILL FILL_0_NAND2X1_242 ( );
FILL FILL_1_NAND2X1_242 ( );
FILL FILL_2_NAND2X1_242 ( );
FILL FILL_3_NAND2X1_242 ( );
FILL FILL_4_NAND2X1_242 ( );
FILL FILL_5_NAND2X1_242 ( );
FILL FILL_6_NAND2X1_242 ( );
FILL FILL_0_NAND2X1_76 ( );
FILL FILL_1_NAND2X1_76 ( );
FILL FILL_2_NAND2X1_76 ( );
FILL FILL_3_NAND2X1_76 ( );
FILL FILL_4_NAND2X1_76 ( );
FILL FILL_5_NAND2X1_76 ( );
FILL FILL_6_NAND2X1_76 ( );
FILL FILL_0_OAI22X1_46 ( );
FILL FILL_1_OAI22X1_46 ( );
FILL FILL_2_OAI22X1_46 ( );
FILL FILL_3_OAI22X1_46 ( );
FILL FILL_4_OAI22X1_46 ( );
FILL FILL_5_OAI22X1_46 ( );
FILL FILL_6_OAI22X1_46 ( );
FILL FILL_7_OAI22X1_46 ( );
FILL FILL_8_OAI22X1_46 ( );
FILL FILL_9_OAI22X1_46 ( );
FILL FILL_10_OAI22X1_46 ( );
FILL FILL_11_OAI22X1_46 ( );
FILL FILL_0_INVX1_185 ( );
FILL FILL_1_INVX1_185 ( );
FILL FILL_2_INVX1_185 ( );
FILL FILL_3_INVX1_185 ( );
FILL FILL_4_INVX1_185 ( );
FILL FILL_0_NAND2X1_151 ( );
FILL FILL_1_NAND2X1_151 ( );
FILL FILL_2_NAND2X1_151 ( );
FILL FILL_3_NAND2X1_151 ( );
FILL FILL_4_NAND2X1_151 ( );
FILL FILL_5_NAND2X1_151 ( );
FILL FILL_6_NAND2X1_151 ( );
FILL FILL_0_NAND2X1_137 ( );
FILL FILL_1_NAND2X1_137 ( );
FILL FILL_2_NAND2X1_137 ( );
FILL FILL_3_NAND2X1_137 ( );
FILL FILL_4_NAND2X1_137 ( );
FILL FILL_5_NAND2X1_137 ( );
FILL FILL_6_NAND2X1_137 ( );
FILL FILL_0_INVX1_91 ( );
FILL FILL_1_INVX1_91 ( );
FILL FILL_2_INVX1_91 ( );
FILL FILL_3_INVX1_91 ( );
FILL FILL_4_INVX1_91 ( );
FILL FILL_0_OAI21X1_137 ( );
FILL FILL_1_OAI21X1_137 ( );
FILL FILL_2_OAI21X1_137 ( );
FILL FILL_3_OAI21X1_137 ( );
FILL FILL_4_OAI21X1_137 ( );
FILL FILL_5_OAI21X1_137 ( );
FILL FILL_6_OAI21X1_137 ( );
FILL FILL_7_OAI21X1_137 ( );
FILL FILL_8_OAI21X1_137 ( );
FILL FILL_0_OAI21X1_142 ( );
FILL FILL_1_OAI21X1_142 ( );
FILL FILL_2_OAI21X1_142 ( );
FILL FILL_3_OAI21X1_142 ( );
FILL FILL_4_OAI21X1_142 ( );
FILL FILL_5_OAI21X1_142 ( );
FILL FILL_6_OAI21X1_142 ( );
FILL FILL_7_OAI21X1_142 ( );
FILL FILL_8_OAI21X1_142 ( );
FILL FILL_0_INVX1_160 ( );
FILL FILL_1_INVX1_160 ( );
FILL FILL_2_INVX1_160 ( );
FILL FILL_3_INVX1_160 ( );
FILL FILL_4_INVX1_160 ( );
FILL FILL_0_NAND2X1_22 ( );
FILL FILL_1_NAND2X1_22 ( );
FILL FILL_2_NAND2X1_22 ( );
FILL FILL_3_NAND2X1_22 ( );
FILL FILL_4_NAND2X1_22 ( );
FILL FILL_5_NAND2X1_22 ( );
FILL FILL_6_NAND2X1_22 ( );
FILL FILL_0_XOR2X1_17 ( );
FILL FILL_1_XOR2X1_17 ( );
FILL FILL_2_XOR2X1_17 ( );
FILL FILL_3_XOR2X1_17 ( );
FILL FILL_4_XOR2X1_17 ( );
FILL FILL_5_XOR2X1_17 ( );
FILL FILL_6_XOR2X1_17 ( );
FILL FILL_7_XOR2X1_17 ( );
FILL FILL_8_XOR2X1_17 ( );
FILL FILL_9_XOR2X1_17 ( );
FILL FILL_10_XOR2X1_17 ( );
FILL FILL_11_XOR2X1_17 ( );
FILL FILL_12_XOR2X1_17 ( );
FILL FILL_13_XOR2X1_17 ( );
FILL FILL_14_XOR2X1_17 ( );
FILL FILL_15_XOR2X1_17 ( );
FILL FILL_0_DFFSR_62 ( );
FILL FILL_1_DFFSR_62 ( );
FILL FILL_2_DFFSR_62 ( );
FILL FILL_3_DFFSR_62 ( );
FILL FILL_4_DFFSR_62 ( );
FILL FILL_5_DFFSR_62 ( );
FILL FILL_6_DFFSR_62 ( );
FILL FILL_7_DFFSR_62 ( );
FILL FILL_8_DFFSR_62 ( );
FILL FILL_9_DFFSR_62 ( );
FILL FILL_10_DFFSR_62 ( );
FILL FILL_11_DFFSR_62 ( );
FILL FILL_12_DFFSR_62 ( );
FILL FILL_13_DFFSR_62 ( );
FILL FILL_14_DFFSR_62 ( );
FILL FILL_15_DFFSR_62 ( );
FILL FILL_16_DFFSR_62 ( );
FILL FILL_17_DFFSR_62 ( );
FILL FILL_18_DFFSR_62 ( );
FILL FILL_19_DFFSR_62 ( );
FILL FILL_20_DFFSR_62 ( );
FILL FILL_21_DFFSR_62 ( );
FILL FILL_22_DFFSR_62 ( );
FILL FILL_23_DFFSR_62 ( );
FILL FILL_24_DFFSR_62 ( );
FILL FILL_25_DFFSR_62 ( );
FILL FILL_26_DFFSR_62 ( );
FILL FILL_27_DFFSR_62 ( );
FILL FILL_28_DFFSR_62 ( );
FILL FILL_29_DFFSR_62 ( );
FILL FILL_30_DFFSR_62 ( );
FILL FILL_31_DFFSR_62 ( );
FILL FILL_32_DFFSR_62 ( );
FILL FILL_33_DFFSR_62 ( );
FILL FILL_34_DFFSR_62 ( );
FILL FILL_35_DFFSR_62 ( );
FILL FILL_36_DFFSR_62 ( );
FILL FILL_37_DFFSR_62 ( );
FILL FILL_38_DFFSR_62 ( );
FILL FILL_39_DFFSR_62 ( );
FILL FILL_40_DFFSR_62 ( );
FILL FILL_41_DFFSR_62 ( );
FILL FILL_42_DFFSR_62 ( );
FILL FILL_43_DFFSR_62 ( );
FILL FILL_44_DFFSR_62 ( );
FILL FILL_45_DFFSR_62 ( );
FILL FILL_46_DFFSR_62 ( );
FILL FILL_47_DFFSR_62 ( );
FILL FILL_48_DFFSR_62 ( );
FILL FILL_49_DFFSR_62 ( );
FILL FILL_50_DFFSR_62 ( );
FILL FILL_0_XOR2X1_9 ( );
FILL FILL_1_XOR2X1_9 ( );
FILL FILL_2_XOR2X1_9 ( );
FILL FILL_3_XOR2X1_9 ( );
FILL FILL_4_XOR2X1_9 ( );
FILL FILL_5_XOR2X1_9 ( );
FILL FILL_6_XOR2X1_9 ( );
FILL FILL_7_XOR2X1_9 ( );
FILL FILL_8_XOR2X1_9 ( );
FILL FILL_9_XOR2X1_9 ( );
FILL FILL_10_XOR2X1_9 ( );
FILL FILL_11_XOR2X1_9 ( );
FILL FILL_12_XOR2X1_9 ( );
FILL FILL_13_XOR2X1_9 ( );
FILL FILL_14_XOR2X1_9 ( );
FILL FILL_15_XOR2X1_9 ( );
FILL FILL_16_XOR2X1_9 ( );
FILL FILL_0_INVX1_404 ( );
FILL FILL_1_INVX1_404 ( );
FILL FILL_2_INVX1_404 ( );
FILL FILL_3_INVX1_404 ( );
FILL FILL_4_INVX1_404 ( );
FILL FILL_0_NAND3X1_130 ( );
FILL FILL_1_NAND3X1_130 ( );
FILL FILL_2_NAND3X1_130 ( );
FILL FILL_3_NAND3X1_130 ( );
FILL FILL_4_NAND3X1_130 ( );
FILL FILL_5_NAND3X1_130 ( );
FILL FILL_6_NAND3X1_130 ( );
FILL FILL_7_NAND3X1_130 ( );
FILL FILL_8_NAND3X1_130 ( );
FILL FILL_0_NAND2X1_254 ( );
FILL FILL_1_NAND2X1_254 ( );
FILL FILL_2_NAND2X1_254 ( );
FILL FILL_3_NAND2X1_254 ( );
FILL FILL_4_NAND2X1_254 ( );
FILL FILL_5_NAND2X1_254 ( );
FILL FILL_6_NAND2X1_254 ( );
FILL FILL_0_INVX1_289 ( );
FILL FILL_1_INVX1_289 ( );
FILL FILL_2_INVX1_289 ( );
FILL FILL_3_INVX1_289 ( );
FILL FILL_4_INVX1_289 ( );
FILL FILL_0_OAI21X1_33 ( );
FILL FILL_1_OAI21X1_33 ( );
FILL FILL_2_OAI21X1_33 ( );
FILL FILL_3_OAI21X1_33 ( );
FILL FILL_4_OAI21X1_33 ( );
FILL FILL_5_OAI21X1_33 ( );
FILL FILL_6_OAI21X1_33 ( );
FILL FILL_7_OAI21X1_33 ( );
FILL FILL_8_OAI21X1_33 ( );
FILL FILL_9_OAI21X1_33 ( );
FILL FILL_0_NAND2X1_33 ( );
FILL FILL_1_NAND2X1_33 ( );
FILL FILL_2_NAND2X1_33 ( );
FILL FILL_3_NAND2X1_33 ( );
FILL FILL_4_NAND2X1_33 ( );
FILL FILL_5_NAND2X1_33 ( );
FILL FILL_6_NAND2X1_33 ( );
FILL FILL_0_DFFSR_171 ( );
FILL FILL_1_DFFSR_171 ( );
FILL FILL_2_DFFSR_171 ( );
FILL FILL_3_DFFSR_171 ( );
FILL FILL_4_DFFSR_171 ( );
FILL FILL_5_DFFSR_171 ( );
FILL FILL_6_DFFSR_171 ( );
FILL FILL_7_DFFSR_171 ( );
FILL FILL_8_DFFSR_171 ( );
FILL FILL_9_DFFSR_171 ( );
FILL FILL_10_DFFSR_171 ( );
FILL FILL_11_DFFSR_171 ( );
FILL FILL_12_DFFSR_171 ( );
FILL FILL_13_DFFSR_171 ( );
FILL FILL_14_DFFSR_171 ( );
FILL FILL_15_DFFSR_171 ( );
FILL FILL_16_DFFSR_171 ( );
FILL FILL_17_DFFSR_171 ( );
FILL FILL_18_DFFSR_171 ( );
FILL FILL_19_DFFSR_171 ( );
FILL FILL_20_DFFSR_171 ( );
FILL FILL_21_DFFSR_171 ( );
FILL FILL_22_DFFSR_171 ( );
FILL FILL_23_DFFSR_171 ( );
FILL FILL_24_DFFSR_171 ( );
FILL FILL_25_DFFSR_171 ( );
FILL FILL_26_DFFSR_171 ( );
FILL FILL_27_DFFSR_171 ( );
FILL FILL_28_DFFSR_171 ( );
FILL FILL_29_DFFSR_171 ( );
FILL FILL_30_DFFSR_171 ( );
FILL FILL_31_DFFSR_171 ( );
FILL FILL_32_DFFSR_171 ( );
FILL FILL_33_DFFSR_171 ( );
FILL FILL_34_DFFSR_171 ( );
FILL FILL_35_DFFSR_171 ( );
FILL FILL_36_DFFSR_171 ( );
FILL FILL_37_DFFSR_171 ( );
FILL FILL_38_DFFSR_171 ( );
FILL FILL_39_DFFSR_171 ( );
FILL FILL_40_DFFSR_171 ( );
FILL FILL_41_DFFSR_171 ( );
FILL FILL_42_DFFSR_171 ( );
FILL FILL_43_DFFSR_171 ( );
FILL FILL_44_DFFSR_171 ( );
FILL FILL_45_DFFSR_171 ( );
FILL FILL_46_DFFSR_171 ( );
FILL FILL_47_DFFSR_171 ( );
FILL FILL_48_DFFSR_171 ( );
FILL FILL_49_DFFSR_171 ( );
FILL FILL_50_DFFSR_171 ( );
FILL FILL_51_DFFSR_171 ( );
FILL FILL_0_NAND2X1_224 ( );
FILL FILL_1_NAND2X1_224 ( );
FILL FILL_2_NAND2X1_224 ( );
FILL FILL_3_NAND2X1_224 ( );
FILL FILL_4_NAND2X1_224 ( );
FILL FILL_5_NAND2X1_224 ( );
FILL FILL_6_NAND2X1_224 ( );
FILL FILL_0_NAND2X1_181 ( );
FILL FILL_1_NAND2X1_181 ( );
FILL FILL_2_NAND2X1_181 ( );
FILL FILL_3_NAND2X1_181 ( );
FILL FILL_4_NAND2X1_181 ( );
FILL FILL_5_NAND2X1_181 ( );
FILL FILL_6_NAND2X1_181 ( );
FILL FILL_0_OAI21X1_184 ( );
FILL FILL_1_OAI21X1_184 ( );
FILL FILL_2_OAI21X1_184 ( );
FILL FILL_3_OAI21X1_184 ( );
FILL FILL_4_OAI21X1_184 ( );
FILL FILL_5_OAI21X1_184 ( );
FILL FILL_6_OAI21X1_184 ( );
FILL FILL_7_OAI21X1_184 ( );
FILL FILL_8_OAI21X1_184 ( );
FILL FILL_0_NAND2X1_185 ( );
FILL FILL_1_NAND2X1_185 ( );
FILL FILL_2_NAND2X1_185 ( );
FILL FILL_3_NAND2X1_185 ( );
FILL FILL_4_NAND2X1_185 ( );
FILL FILL_5_NAND2X1_185 ( );
FILL FILL_6_NAND2X1_185 ( );
FILL FILL_0_NAND3X1_15 ( );
FILL FILL_1_NAND3X1_15 ( );
FILL FILL_2_NAND3X1_15 ( );
FILL FILL_3_NAND3X1_15 ( );
FILL FILL_4_NAND3X1_15 ( );
FILL FILL_5_NAND3X1_15 ( );
FILL FILL_6_NAND3X1_15 ( );
FILL FILL_7_NAND3X1_15 ( );
FILL FILL_8_NAND3X1_15 ( );
FILL FILL_0_NAND3X1_9 ( );
FILL FILL_1_NAND3X1_9 ( );
FILL FILL_2_NAND3X1_9 ( );
FILL FILL_3_NAND3X1_9 ( );
FILL FILL_4_NAND3X1_9 ( );
FILL FILL_5_NAND3X1_9 ( );
FILL FILL_6_NAND3X1_9 ( );
FILL FILL_7_NAND3X1_9 ( );
FILL FILL_8_NAND3X1_9 ( );
FILL FILL_9_NAND3X1_9 ( );
FILL FILL_0_NAND3X1_14 ( );
FILL FILL_1_NAND3X1_14 ( );
FILL FILL_2_NAND3X1_14 ( );
FILL FILL_3_NAND3X1_14 ( );
FILL FILL_4_NAND3X1_14 ( );
FILL FILL_5_NAND3X1_14 ( );
FILL FILL_6_NAND3X1_14 ( );
FILL FILL_7_NAND3X1_14 ( );
FILL FILL_8_NAND3X1_14 ( );
FILL FILL_9_NAND3X1_14 ( );
FILL FILL_0_NAND3X1_16 ( );
FILL FILL_1_NAND3X1_16 ( );
FILL FILL_2_NAND3X1_16 ( );
FILL FILL_3_NAND3X1_16 ( );
FILL FILL_4_NAND3X1_16 ( );
FILL FILL_5_NAND3X1_16 ( );
FILL FILL_6_NAND3X1_16 ( );
FILL FILL_7_NAND3X1_16 ( );
FILL FILL_8_NAND3X1_16 ( );
FILL FILL_0_NAND2X1_270 ( );
FILL FILL_1_NAND2X1_270 ( );
FILL FILL_2_NAND2X1_270 ( );
FILL FILL_3_NAND2X1_270 ( );
FILL FILL_4_NAND2X1_270 ( );
FILL FILL_5_NAND2X1_270 ( );
FILL FILL_6_NAND2X1_270 ( );
FILL FILL_0_NAND3X1_86 ( );
FILL FILL_1_NAND3X1_86 ( );
FILL FILL_2_NAND3X1_86 ( );
FILL FILL_3_NAND3X1_86 ( );
FILL FILL_4_NAND3X1_86 ( );
FILL FILL_5_NAND3X1_86 ( );
FILL FILL_6_NAND3X1_86 ( );
FILL FILL_7_NAND3X1_86 ( );
FILL FILL_8_NAND3X1_86 ( );
FILL FILL_0_NAND3X1_81 ( );
FILL FILL_1_NAND3X1_81 ( );
FILL FILL_2_NAND3X1_81 ( );
FILL FILL_3_NAND3X1_81 ( );
FILL FILL_4_NAND3X1_81 ( );
FILL FILL_5_NAND3X1_81 ( );
FILL FILL_6_NAND3X1_81 ( );
FILL FILL_7_NAND3X1_81 ( );
FILL FILL_8_NAND3X1_81 ( );
FILL FILL_0_OAI21X1_238 ( );
FILL FILL_1_OAI21X1_238 ( );
FILL FILL_2_OAI21X1_238 ( );
FILL FILL_3_OAI21X1_238 ( );
FILL FILL_4_OAI21X1_238 ( );
FILL FILL_5_OAI21X1_238 ( );
FILL FILL_6_OAI21X1_238 ( );
FILL FILL_7_OAI21X1_238 ( );
FILL FILL_8_OAI21X1_238 ( );
FILL FILL_0_INVX1_261 ( );
FILL FILL_1_INVX1_261 ( );
FILL FILL_2_INVX1_261 ( );
FILL FILL_3_INVX1_261 ( );
FILL FILL_4_INVX1_261 ( );
FILL FILL_0_DFFSR_122 ( );
FILL FILL_1_DFFSR_122 ( );
FILL FILL_2_DFFSR_122 ( );
FILL FILL_3_DFFSR_122 ( );
FILL FILL_4_DFFSR_122 ( );
FILL FILL_5_DFFSR_122 ( );
FILL FILL_6_DFFSR_122 ( );
FILL FILL_7_DFFSR_122 ( );
FILL FILL_8_DFFSR_122 ( );
FILL FILL_9_DFFSR_122 ( );
FILL FILL_10_DFFSR_122 ( );
FILL FILL_11_DFFSR_122 ( );
FILL FILL_12_DFFSR_122 ( );
FILL FILL_13_DFFSR_122 ( );
FILL FILL_14_DFFSR_122 ( );
FILL FILL_15_DFFSR_122 ( );
FILL FILL_16_DFFSR_122 ( );
FILL FILL_17_DFFSR_122 ( );
FILL FILL_18_DFFSR_122 ( );
FILL FILL_19_DFFSR_122 ( );
FILL FILL_20_DFFSR_122 ( );
FILL FILL_21_DFFSR_122 ( );
FILL FILL_22_DFFSR_122 ( );
FILL FILL_23_DFFSR_122 ( );
FILL FILL_24_DFFSR_122 ( );
FILL FILL_25_DFFSR_122 ( );
FILL FILL_26_DFFSR_122 ( );
FILL FILL_27_DFFSR_122 ( );
FILL FILL_28_DFFSR_122 ( );
FILL FILL_29_DFFSR_122 ( );
FILL FILL_30_DFFSR_122 ( );
FILL FILL_31_DFFSR_122 ( );
FILL FILL_32_DFFSR_122 ( );
FILL FILL_33_DFFSR_122 ( );
FILL FILL_34_DFFSR_122 ( );
FILL FILL_35_DFFSR_122 ( );
FILL FILL_36_DFFSR_122 ( );
FILL FILL_37_DFFSR_122 ( );
FILL FILL_38_DFFSR_122 ( );
FILL FILL_39_DFFSR_122 ( );
FILL FILL_40_DFFSR_122 ( );
FILL FILL_41_DFFSR_122 ( );
FILL FILL_42_DFFSR_122 ( );
FILL FILL_43_DFFSR_122 ( );
FILL FILL_44_DFFSR_122 ( );
FILL FILL_45_DFFSR_122 ( );
FILL FILL_46_DFFSR_122 ( );
FILL FILL_47_DFFSR_122 ( );
FILL FILL_48_DFFSR_122 ( );
FILL FILL_49_DFFSR_122 ( );
FILL FILL_50_DFFSR_122 ( );
FILL FILL_51_DFFSR_122 ( );
FILL FILL_0_INVX1_386 ( );
FILL FILL_1_INVX1_386 ( );
FILL FILL_2_INVX1_386 ( );
FILL FILL_3_INVX1_386 ( );
FILL FILL_4_INVX1_386 ( );
FILL FILL_0_INVX1_345 ( );
FILL FILL_1_INVX1_345 ( );
FILL FILL_2_INVX1_345 ( );
FILL FILL_3_INVX1_345 ( );
FILL FILL_0_NOR2X1_28 ( );
FILL FILL_1_NOR2X1_28 ( );
FILL FILL_2_NOR2X1_28 ( );
FILL FILL_3_NOR2X1_28 ( );
FILL FILL_4_NOR2X1_28 ( );
FILL FILL_5_NOR2X1_28 ( );
FILL FILL_6_NOR2X1_28 ( );
FILL FILL_0_NOR2X1_35 ( );
FILL FILL_1_NOR2X1_35 ( );
FILL FILL_2_NOR2X1_35 ( );
FILL FILL_3_NOR2X1_35 ( );
FILL FILL_4_NOR2X1_35 ( );
FILL FILL_5_NOR2X1_35 ( );
FILL FILL_6_NOR2X1_35 ( );
FILL FILL_0_OAI21X1_83 ( );
FILL FILL_1_OAI21X1_83 ( );
FILL FILL_2_OAI21X1_83 ( );
FILL FILL_3_OAI21X1_83 ( );
FILL FILL_4_OAI21X1_83 ( );
FILL FILL_5_OAI21X1_83 ( );
FILL FILL_6_OAI21X1_83 ( );
FILL FILL_7_OAI21X1_83 ( );
FILL FILL_8_OAI21X1_83 ( );
FILL FILL_9_OAI21X1_83 ( );
FILL FILL_0_INVX1_94 ( );
FILL FILL_1_INVX1_94 ( );
FILL FILL_2_INVX1_94 ( );
FILL FILL_3_INVX1_94 ( );
FILL FILL_0_NOR2X1_32 ( );
FILL FILL_1_NOR2X1_32 ( );
FILL FILL_2_NOR2X1_32 ( );
FILL FILL_3_NOR2X1_32 ( );
FILL FILL_4_NOR2X1_32 ( );
FILL FILL_5_NOR2X1_32 ( );
FILL FILL_6_NOR2X1_32 ( );
FILL FILL_0_OAI21X1_150 ( );
FILL FILL_1_OAI21X1_150 ( );
FILL FILL_2_OAI21X1_150 ( );
FILL FILL_3_OAI21X1_150 ( );
FILL FILL_4_OAI21X1_150 ( );
FILL FILL_5_OAI21X1_150 ( );
FILL FILL_6_OAI21X1_150 ( );
FILL FILL_7_OAI21X1_150 ( );
FILL FILL_8_OAI21X1_150 ( );
FILL FILL_0_NAND2X1_244 ( );
FILL FILL_1_NAND2X1_244 ( );
FILL FILL_2_NAND2X1_244 ( );
FILL FILL_3_NAND2X1_244 ( );
FILL FILL_4_NAND2X1_244 ( );
FILL FILL_5_NAND2X1_244 ( );
FILL FILL_6_NAND2X1_244 ( );
FILL FILL_0_INVX1_175 ( );
FILL FILL_1_INVX1_175 ( );
FILL FILL_2_INVX1_175 ( );
FILL FILL_3_INVX1_175 ( );
FILL FILL_4_INVX1_175 ( );
FILL FILL_0_OAI21X1_141 ( );
FILL FILL_1_OAI21X1_141 ( );
FILL FILL_2_OAI21X1_141 ( );
FILL FILL_3_OAI21X1_141 ( );
FILL FILL_4_OAI21X1_141 ( );
FILL FILL_5_OAI21X1_141 ( );
FILL FILL_6_OAI21X1_141 ( );
FILL FILL_7_OAI21X1_141 ( );
FILL FILL_8_OAI21X1_141 ( );
FILL FILL_0_INVX1_155 ( );
FILL FILL_1_INVX1_155 ( );
FILL FILL_2_INVX1_155 ( );
FILL FILL_3_INVX1_155 ( );
FILL FILL_4_INVX1_155 ( );
FILL FILL_0_INVX1_159 ( );
FILL FILL_1_INVX1_159 ( );
FILL FILL_2_INVX1_159 ( );
FILL FILL_3_INVX1_159 ( );
FILL FILL_4_INVX1_159 ( );
FILL FILL_0_INVX1_163 ( );
FILL FILL_1_INVX1_163 ( );
FILL FILL_2_INVX1_163 ( );
FILL FILL_3_INVX1_163 ( );
FILL FILL_4_INVX1_163 ( );
FILL FILL_0_DFFSR_63 ( );
FILL FILL_1_DFFSR_63 ( );
FILL FILL_2_DFFSR_63 ( );
FILL FILL_3_DFFSR_63 ( );
FILL FILL_4_DFFSR_63 ( );
FILL FILL_5_DFFSR_63 ( );
FILL FILL_6_DFFSR_63 ( );
FILL FILL_7_DFFSR_63 ( );
FILL FILL_8_DFFSR_63 ( );
FILL FILL_9_DFFSR_63 ( );
FILL FILL_10_DFFSR_63 ( );
FILL FILL_11_DFFSR_63 ( );
FILL FILL_12_DFFSR_63 ( );
FILL FILL_13_DFFSR_63 ( );
FILL FILL_14_DFFSR_63 ( );
FILL FILL_15_DFFSR_63 ( );
FILL FILL_16_DFFSR_63 ( );
FILL FILL_17_DFFSR_63 ( );
FILL FILL_18_DFFSR_63 ( );
FILL FILL_19_DFFSR_63 ( );
FILL FILL_20_DFFSR_63 ( );
FILL FILL_21_DFFSR_63 ( );
FILL FILL_22_DFFSR_63 ( );
FILL FILL_23_DFFSR_63 ( );
FILL FILL_24_DFFSR_63 ( );
FILL FILL_25_DFFSR_63 ( );
FILL FILL_26_DFFSR_63 ( );
FILL FILL_27_DFFSR_63 ( );
FILL FILL_28_DFFSR_63 ( );
FILL FILL_29_DFFSR_63 ( );
FILL FILL_30_DFFSR_63 ( );
FILL FILL_31_DFFSR_63 ( );
FILL FILL_32_DFFSR_63 ( );
FILL FILL_33_DFFSR_63 ( );
FILL FILL_34_DFFSR_63 ( );
FILL FILL_35_DFFSR_63 ( );
FILL FILL_36_DFFSR_63 ( );
FILL FILL_37_DFFSR_63 ( );
FILL FILL_38_DFFSR_63 ( );
FILL FILL_39_DFFSR_63 ( );
FILL FILL_40_DFFSR_63 ( );
FILL FILL_41_DFFSR_63 ( );
FILL FILL_42_DFFSR_63 ( );
FILL FILL_43_DFFSR_63 ( );
FILL FILL_44_DFFSR_63 ( );
FILL FILL_45_DFFSR_63 ( );
FILL FILL_46_DFFSR_63 ( );
FILL FILL_47_DFFSR_63 ( );
FILL FILL_48_DFFSR_63 ( );
FILL FILL_49_DFFSR_63 ( );
FILL FILL_50_DFFSR_63 ( );
FILL FILL_51_DFFSR_63 ( );
FILL FILL_0_INVX1_37 ( );
FILL FILL_1_INVX1_37 ( );
FILL FILL_2_INVX1_37 ( );
FILL FILL_3_INVX1_37 ( );
FILL FILL_4_INVX1_37 ( );
FILL FILL_0_INVX1_311 ( );
FILL FILL_1_INVX1_311 ( );
FILL FILL_2_INVX1_311 ( );
FILL FILL_3_INVX1_311 ( );
FILL FILL_4_INVX1_311 ( );
FILL FILL_0_OAI22X1_26 ( );
FILL FILL_1_OAI22X1_26 ( );
FILL FILL_2_OAI22X1_26 ( );
FILL FILL_3_OAI22X1_26 ( );
FILL FILL_4_OAI22X1_26 ( );
FILL FILL_5_OAI22X1_26 ( );
FILL FILL_6_OAI22X1_26 ( );
FILL FILL_7_OAI22X1_26 ( );
FILL FILL_8_OAI22X1_26 ( );
FILL FILL_9_OAI22X1_26 ( );
FILL FILL_10_OAI22X1_26 ( );
FILL FILL_0_DFFSR_33 ( );
FILL FILL_1_DFFSR_33 ( );
FILL FILL_2_DFFSR_33 ( );
FILL FILL_3_DFFSR_33 ( );
FILL FILL_4_DFFSR_33 ( );
FILL FILL_5_DFFSR_33 ( );
FILL FILL_6_DFFSR_33 ( );
FILL FILL_7_DFFSR_33 ( );
FILL FILL_8_DFFSR_33 ( );
FILL FILL_9_DFFSR_33 ( );
FILL FILL_10_DFFSR_33 ( );
FILL FILL_11_DFFSR_33 ( );
FILL FILL_12_DFFSR_33 ( );
FILL FILL_13_DFFSR_33 ( );
FILL FILL_14_DFFSR_33 ( );
FILL FILL_15_DFFSR_33 ( );
FILL FILL_16_DFFSR_33 ( );
FILL FILL_17_DFFSR_33 ( );
FILL FILL_18_DFFSR_33 ( );
FILL FILL_19_DFFSR_33 ( );
FILL FILL_20_DFFSR_33 ( );
FILL FILL_21_DFFSR_33 ( );
FILL FILL_22_DFFSR_33 ( );
FILL FILL_23_DFFSR_33 ( );
FILL FILL_24_DFFSR_33 ( );
FILL FILL_25_DFFSR_33 ( );
FILL FILL_26_DFFSR_33 ( );
FILL FILL_27_DFFSR_33 ( );
FILL FILL_28_DFFSR_33 ( );
FILL FILL_29_DFFSR_33 ( );
FILL FILL_30_DFFSR_33 ( );
FILL FILL_31_DFFSR_33 ( );
FILL FILL_32_DFFSR_33 ( );
FILL FILL_33_DFFSR_33 ( );
FILL FILL_34_DFFSR_33 ( );
FILL FILL_35_DFFSR_33 ( );
FILL FILL_36_DFFSR_33 ( );
FILL FILL_37_DFFSR_33 ( );
FILL FILL_38_DFFSR_33 ( );
FILL FILL_39_DFFSR_33 ( );
FILL FILL_40_DFFSR_33 ( );
FILL FILL_41_DFFSR_33 ( );
FILL FILL_42_DFFSR_33 ( );
FILL FILL_43_DFFSR_33 ( );
FILL FILL_44_DFFSR_33 ( );
FILL FILL_45_DFFSR_33 ( );
FILL FILL_46_DFFSR_33 ( );
FILL FILL_47_DFFSR_33 ( );
FILL FILL_48_DFFSR_33 ( );
FILL FILL_49_DFFSR_33 ( );
FILL FILL_50_DFFSR_33 ( );
FILL FILL_51_DFFSR_33 ( );
FILL FILL_0_INVX1_38 ( );
FILL FILL_1_INVX1_38 ( );
FILL FILL_2_INVX1_38 ( );
FILL FILL_3_INVX1_38 ( );
FILL FILL_0_DFFSR_52 ( );
FILL FILL_1_DFFSR_52 ( );
FILL FILL_2_DFFSR_52 ( );
FILL FILL_3_DFFSR_52 ( );
FILL FILL_4_DFFSR_52 ( );
FILL FILL_5_DFFSR_52 ( );
FILL FILL_6_DFFSR_52 ( );
FILL FILL_7_DFFSR_52 ( );
FILL FILL_8_DFFSR_52 ( );
FILL FILL_9_DFFSR_52 ( );
FILL FILL_10_DFFSR_52 ( );
FILL FILL_11_DFFSR_52 ( );
FILL FILL_12_DFFSR_52 ( );
FILL FILL_13_DFFSR_52 ( );
FILL FILL_14_DFFSR_52 ( );
FILL FILL_15_DFFSR_52 ( );
FILL FILL_16_DFFSR_52 ( );
FILL FILL_17_DFFSR_52 ( );
FILL FILL_18_DFFSR_52 ( );
FILL FILL_19_DFFSR_52 ( );
FILL FILL_20_DFFSR_52 ( );
FILL FILL_21_DFFSR_52 ( );
FILL FILL_22_DFFSR_52 ( );
FILL FILL_23_DFFSR_52 ( );
FILL FILL_24_DFFSR_52 ( );
FILL FILL_25_DFFSR_52 ( );
FILL FILL_26_DFFSR_52 ( );
FILL FILL_27_DFFSR_52 ( );
FILL FILL_28_DFFSR_52 ( );
FILL FILL_29_DFFSR_52 ( );
FILL FILL_30_DFFSR_52 ( );
FILL FILL_31_DFFSR_52 ( );
FILL FILL_32_DFFSR_52 ( );
FILL FILL_33_DFFSR_52 ( );
FILL FILL_34_DFFSR_52 ( );
FILL FILL_35_DFFSR_52 ( );
FILL FILL_36_DFFSR_52 ( );
FILL FILL_37_DFFSR_52 ( );
FILL FILL_38_DFFSR_52 ( );
FILL FILL_39_DFFSR_52 ( );
FILL FILL_40_DFFSR_52 ( );
FILL FILL_41_DFFSR_52 ( );
FILL FILL_42_DFFSR_52 ( );
FILL FILL_43_DFFSR_52 ( );
FILL FILL_44_DFFSR_52 ( );
FILL FILL_45_DFFSR_52 ( );
FILL FILL_46_DFFSR_52 ( );
FILL FILL_47_DFFSR_52 ( );
FILL FILL_48_DFFSR_52 ( );
FILL FILL_49_DFFSR_52 ( );
FILL FILL_50_DFFSR_52 ( );
FILL FILL_0_INVX1_220 ( );
FILL FILL_1_INVX1_220 ( );
FILL FILL_2_INVX1_220 ( );
FILL FILL_3_INVX1_220 ( );
FILL FILL_0_NAND3X1_4 ( );
FILL FILL_1_NAND3X1_4 ( );
FILL FILL_2_NAND3X1_4 ( );
FILL FILL_3_NAND3X1_4 ( );
FILL FILL_4_NAND3X1_4 ( );
FILL FILL_5_NAND3X1_4 ( );
FILL FILL_6_NAND3X1_4 ( );
FILL FILL_7_NAND3X1_4 ( );
FILL FILL_8_NAND3X1_4 ( );
FILL FILL_9_NAND3X1_4 ( );
FILL FILL_0_AOI21X1_2 ( );
FILL FILL_1_AOI21X1_2 ( );
FILL FILL_2_AOI21X1_2 ( );
FILL FILL_3_AOI21X1_2 ( );
FILL FILL_4_AOI21X1_2 ( );
FILL FILL_5_AOI21X1_2 ( );
FILL FILL_6_AOI21X1_2 ( );
FILL FILL_7_AOI21X1_2 ( );
FILL FILL_8_AOI21X1_2 ( );
FILL FILL_0_INVX1_219 ( );
FILL FILL_1_INVX1_219 ( );
FILL FILL_2_INVX1_219 ( );
FILL FILL_3_INVX1_219 ( );
FILL FILL_0_NAND2X1_180 ( );
FILL FILL_1_NAND2X1_180 ( );
FILL FILL_2_NAND2X1_180 ( );
FILL FILL_3_NAND2X1_180 ( );
FILL FILL_4_NAND2X1_180 ( );
FILL FILL_5_NAND2X1_180 ( );
FILL FILL_6_NAND2X1_180 ( );
FILL FILL_0_AOI21X1_8 ( );
FILL FILL_1_AOI21X1_8 ( );
FILL FILL_2_AOI21X1_8 ( );
FILL FILL_3_AOI21X1_8 ( );
FILL FILL_4_AOI21X1_8 ( );
FILL FILL_5_AOI21X1_8 ( );
FILL FILL_6_AOI21X1_8 ( );
FILL FILL_7_AOI21X1_8 ( );
FILL FILL_8_AOI21X1_8 ( );
FILL FILL_9_AOI21X1_8 ( );
FILL FILL_0_NAND3X1_12 ( );
FILL FILL_1_NAND3X1_12 ( );
FILL FILL_2_NAND3X1_12 ( );
FILL FILL_3_NAND3X1_12 ( );
FILL FILL_4_NAND3X1_12 ( );
FILL FILL_5_NAND3X1_12 ( );
FILL FILL_6_NAND3X1_12 ( );
FILL FILL_7_NAND3X1_12 ( );
FILL FILL_8_NAND3X1_12 ( );
FILL FILL_0_AOI21X1_9 ( );
FILL FILL_1_AOI21X1_9 ( );
FILL FILL_2_AOI21X1_9 ( );
FILL FILL_3_AOI21X1_9 ( );
FILL FILL_4_AOI21X1_9 ( );
FILL FILL_5_AOI21X1_9 ( );
FILL FILL_6_AOI21X1_9 ( );
FILL FILL_7_AOI21X1_9 ( );
FILL FILL_8_AOI21X1_9 ( );
FILL FILL_0_NAND3X1_30 ( );
FILL FILL_1_NAND3X1_30 ( );
FILL FILL_2_NAND3X1_30 ( );
FILL FILL_3_NAND3X1_30 ( );
FILL FILL_4_NAND3X1_30 ( );
FILL FILL_5_NAND3X1_30 ( );
FILL FILL_6_NAND3X1_30 ( );
FILL FILL_7_NAND3X1_30 ( );
FILL FILL_8_NAND3X1_30 ( );
FILL FILL_0_NAND3X1_31 ( );
FILL FILL_1_NAND3X1_31 ( );
FILL FILL_2_NAND3X1_31 ( );
FILL FILL_3_NAND3X1_31 ( );
FILL FILL_4_NAND3X1_31 ( );
FILL FILL_5_NAND3X1_31 ( );
FILL FILL_6_NAND3X1_31 ( );
FILL FILL_7_NAND3X1_31 ( );
FILL FILL_8_NAND3X1_31 ( );
FILL FILL_9_NAND3X1_31 ( );
FILL FILL_0_NOR3X1_1 ( );
FILL FILL_1_NOR3X1_1 ( );
FILL FILL_2_NOR3X1_1 ( );
FILL FILL_3_NOR3X1_1 ( );
FILL FILL_4_NOR3X1_1 ( );
FILL FILL_5_NOR3X1_1 ( );
FILL FILL_6_NOR3X1_1 ( );
FILL FILL_7_NOR3X1_1 ( );
FILL FILL_8_NOR3X1_1 ( );
FILL FILL_9_NOR3X1_1 ( );
FILL FILL_10_NOR3X1_1 ( );
FILL FILL_11_NOR3X1_1 ( );
FILL FILL_12_NOR3X1_1 ( );
FILL FILL_13_NOR3X1_1 ( );
FILL FILL_14_NOR3X1_1 ( );
FILL FILL_15_NOR3X1_1 ( );
FILL FILL_16_NOR3X1_1 ( );
FILL FILL_17_NOR3X1_1 ( );
FILL FILL_0_NAND3X1_87 ( );
FILL FILL_1_NAND3X1_87 ( );
FILL FILL_2_NAND3X1_87 ( );
FILL FILL_3_NAND3X1_87 ( );
FILL FILL_4_NAND3X1_87 ( );
FILL FILL_5_NAND3X1_87 ( );
FILL FILL_6_NAND3X1_87 ( );
FILL FILL_7_NAND3X1_87 ( );
FILL FILL_8_NAND3X1_87 ( );
FILL FILL_0_NAND3X1_88 ( );
FILL FILL_1_NAND3X1_88 ( );
FILL FILL_2_NAND3X1_88 ( );
FILL FILL_3_NAND3X1_88 ( );
FILL FILL_4_NAND3X1_88 ( );
FILL FILL_5_NAND3X1_88 ( );
FILL FILL_6_NAND3X1_88 ( );
FILL FILL_7_NAND3X1_88 ( );
FILL FILL_8_NAND3X1_88 ( );
FILL FILL_9_NAND3X1_88 ( );
FILL FILL_0_NAND2X1_122 ( );
FILL FILL_1_NAND2X1_122 ( );
FILL FILL_2_NAND2X1_122 ( );
FILL FILL_3_NAND2X1_122 ( );
FILL FILL_4_NAND2X1_122 ( );
FILL FILL_5_NAND2X1_122 ( );
FILL FILL_6_NAND2X1_122 ( );
FILL FILL_0_NAND2X1_81 ( );
FILL FILL_1_NAND2X1_81 ( );
FILL FILL_2_NAND2X1_81 ( );
FILL FILL_3_NAND2X1_81 ( );
FILL FILL_4_NAND2X1_81 ( );
FILL FILL_5_NAND2X1_81 ( );
FILL FILL_6_NAND2X1_81 ( );
FILL FILL_0_OAI21X1_122 ( );
FILL FILL_1_OAI21X1_122 ( );
FILL FILL_2_OAI21X1_122 ( );
FILL FILL_3_OAI21X1_122 ( );
FILL FILL_4_OAI21X1_122 ( );
FILL FILL_5_OAI21X1_122 ( );
FILL FILL_6_OAI21X1_122 ( );
FILL FILL_7_OAI21X1_122 ( );
FILL FILL_8_OAI21X1_122 ( );
FILL FILL_0_INVX1_138 ( );
FILL FILL_1_INVX1_138 ( );
FILL FILL_2_INVX1_138 ( );
FILL FILL_3_INVX1_138 ( );
FILL FILL_4_INVX1_138 ( );
FILL FILL_0_NAND2X1_109 ( );
FILL FILL_1_NAND2X1_109 ( );
FILL FILL_2_NAND2X1_109 ( );
FILL FILL_3_NAND2X1_109 ( );
FILL FILL_4_NAND2X1_109 ( );
FILL FILL_5_NAND2X1_109 ( );
FILL FILL_6_NAND2X1_109 ( );
FILL FILL_0_INVX1_387 ( );
FILL FILL_1_INVX1_387 ( );
FILL FILL_2_INVX1_387 ( );
FILL FILL_3_INVX1_387 ( );
FILL FILL_0_OAI22X1_64 ( );
FILL FILL_1_OAI22X1_64 ( );
FILL FILL_2_OAI22X1_64 ( );
FILL FILL_3_OAI22X1_64 ( );
FILL FILL_4_OAI22X1_64 ( );
FILL FILL_5_OAI22X1_64 ( );
FILL FILL_6_OAI22X1_64 ( );
FILL FILL_7_OAI22X1_64 ( );
FILL FILL_8_OAI22X1_64 ( );
FILL FILL_9_OAI22X1_64 ( );
FILL FILL_10_OAI22X1_64 ( );
FILL FILL_11_OAI22X1_64 ( );
FILL FILL_0_OAI22X1_49 ( );
FILL FILL_1_OAI22X1_49 ( );
FILL FILL_2_OAI22X1_49 ( );
FILL FILL_3_OAI22X1_49 ( );
FILL FILL_4_OAI22X1_49 ( );
FILL FILL_5_OAI22X1_49 ( );
FILL FILL_6_OAI22X1_49 ( );
FILL FILL_7_OAI22X1_49 ( );
FILL FILL_8_OAI22X1_49 ( );
FILL FILL_9_OAI22X1_49 ( );
FILL FILL_10_OAI22X1_49 ( );
FILL FILL_11_OAI22X1_49 ( );
FILL FILL_0_NOR2X1_37 ( );
FILL FILL_1_NOR2X1_37 ( );
FILL FILL_2_NOR2X1_37 ( );
FILL FILL_3_NOR2X1_37 ( );
FILL FILL_4_NOR2X1_37 ( );
FILL FILL_5_NOR2X1_37 ( );
FILL FILL_6_NOR2X1_37 ( );
FILL FILL_0_OAI22X1_52 ( );
FILL FILL_1_OAI22X1_52 ( );
FILL FILL_2_OAI22X1_52 ( );
FILL FILL_3_OAI22X1_52 ( );
FILL FILL_4_OAI22X1_52 ( );
FILL FILL_5_OAI22X1_52 ( );
FILL FILL_6_OAI22X1_52 ( );
FILL FILL_7_OAI22X1_52 ( );
FILL FILL_8_OAI22X1_52 ( );
FILL FILL_9_OAI22X1_52 ( );
FILL FILL_10_OAI22X1_52 ( );
FILL FILL_11_OAI22X1_52 ( );
FILL FILL_0_INVX1_363 ( );
FILL FILL_1_INVX1_363 ( );
FILL FILL_2_INVX1_363 ( );
FILL FILL_3_INVX1_363 ( );
FILL FILL_0_NAND2X1_246 ( );
FILL FILL_1_NAND2X1_246 ( );
FILL FILL_2_NAND2X1_246 ( );
FILL FILL_3_NAND2X1_246 ( );
FILL FILL_4_NAND2X1_246 ( );
FILL FILL_5_NAND2X1_246 ( );
FILL FILL_6_NAND2X1_246 ( );
FILL FILL_0_INVX1_174 ( );
FILL FILL_1_INVX1_174 ( );
FILL FILL_2_INVX1_174 ( );
FILL FILL_3_INVX1_174 ( );
FILL FILL_4_INVX1_174 ( );
FILL FILL_0_NAND2X1_141 ( );
FILL FILL_1_NAND2X1_141 ( );
FILL FILL_2_NAND2X1_141 ( );
FILL FILL_3_NAND2X1_141 ( );
FILL FILL_4_NAND2X1_141 ( );
FILL FILL_5_NAND2X1_141 ( );
FILL FILL_6_NAND2X1_141 ( );
FILL FILL_0_DFFSR_141 ( );
FILL FILL_1_DFFSR_141 ( );
FILL FILL_2_DFFSR_141 ( );
FILL FILL_3_DFFSR_141 ( );
FILL FILL_4_DFFSR_141 ( );
FILL FILL_5_DFFSR_141 ( );
FILL FILL_6_DFFSR_141 ( );
FILL FILL_7_DFFSR_141 ( );
FILL FILL_8_DFFSR_141 ( );
FILL FILL_9_DFFSR_141 ( );
FILL FILL_10_DFFSR_141 ( );
FILL FILL_11_DFFSR_141 ( );
FILL FILL_12_DFFSR_141 ( );
FILL FILL_13_DFFSR_141 ( );
FILL FILL_14_DFFSR_141 ( );
FILL FILL_15_DFFSR_141 ( );
FILL FILL_16_DFFSR_141 ( );
FILL FILL_17_DFFSR_141 ( );
FILL FILL_18_DFFSR_141 ( );
FILL FILL_19_DFFSR_141 ( );
FILL FILL_20_DFFSR_141 ( );
FILL FILL_21_DFFSR_141 ( );
FILL FILL_22_DFFSR_141 ( );
FILL FILL_23_DFFSR_141 ( );
FILL FILL_24_DFFSR_141 ( );
FILL FILL_25_DFFSR_141 ( );
FILL FILL_26_DFFSR_141 ( );
FILL FILL_27_DFFSR_141 ( );
FILL FILL_28_DFFSR_141 ( );
FILL FILL_29_DFFSR_141 ( );
FILL FILL_30_DFFSR_141 ( );
FILL FILL_31_DFFSR_141 ( );
FILL FILL_32_DFFSR_141 ( );
FILL FILL_33_DFFSR_141 ( );
FILL FILL_34_DFFSR_141 ( );
FILL FILL_35_DFFSR_141 ( );
FILL FILL_36_DFFSR_141 ( );
FILL FILL_37_DFFSR_141 ( );
FILL FILL_38_DFFSR_141 ( );
FILL FILL_39_DFFSR_141 ( );
FILL FILL_40_DFFSR_141 ( );
FILL FILL_41_DFFSR_141 ( );
FILL FILL_42_DFFSR_141 ( );
FILL FILL_43_DFFSR_141 ( );
FILL FILL_44_DFFSR_141 ( );
FILL FILL_45_DFFSR_141 ( );
FILL FILL_46_DFFSR_141 ( );
FILL FILL_47_DFFSR_141 ( );
FILL FILL_48_DFFSR_141 ( );
FILL FILL_49_DFFSR_141 ( );
FILL FILL_50_DFFSR_141 ( );
FILL FILL_0_INVX1_306 ( );
FILL FILL_1_INVX1_306 ( );
FILL FILL_2_INVX1_306 ( );
FILL FILL_3_INVX1_306 ( );
FILL FILL_4_INVX1_306 ( );
FILL FILL_0_OAI21X1_63 ( );
FILL FILL_1_OAI21X1_63 ( );
FILL FILL_2_OAI21X1_63 ( );
FILL FILL_3_OAI21X1_63 ( );
FILL FILL_4_OAI21X1_63 ( );
FILL FILL_5_OAI21X1_63 ( );
FILL FILL_6_OAI21X1_63 ( );
FILL FILL_7_OAI21X1_63 ( );
FILL FILL_8_OAI21X1_63 ( );
FILL FILL_9_OAI21X1_63 ( );
FILL FILL_0_INVX1_71 ( );
FILL FILL_1_INVX1_71 ( );
FILL FILL_2_INVX1_71 ( );
FILL FILL_3_INVX1_71 ( );
FILL FILL_0_INVX1_319 ( );
FILL FILL_1_INVX1_319 ( );
FILL FILL_2_INVX1_319 ( );
FILL FILL_3_INVX1_319 ( );
FILL FILL_4_INVX1_319 ( );
FILL FILL_0_NAND3X1_117 ( );
FILL FILL_1_NAND3X1_117 ( );
FILL FILL_2_NAND3X1_117 ( );
FILL FILL_3_NAND3X1_117 ( );
FILL FILL_4_NAND3X1_117 ( );
FILL FILL_5_NAND3X1_117 ( );
FILL FILL_6_NAND3X1_117 ( );
FILL FILL_7_NAND3X1_117 ( );
FILL FILL_8_NAND3X1_117 ( );
FILL FILL_9_NAND3X1_117 ( );
FILL FILL_0_OAI22X1_28 ( );
FILL FILL_1_OAI22X1_28 ( );
FILL FILL_2_OAI22X1_28 ( );
FILL FILL_3_OAI22X1_28 ( );
FILL FILL_4_OAI22X1_28 ( );
FILL FILL_5_OAI22X1_28 ( );
FILL FILL_6_OAI22X1_28 ( );
FILL FILL_7_OAI22X1_28 ( );
FILL FILL_8_OAI22X1_28 ( );
FILL FILL_9_OAI22X1_28 ( );
FILL FILL_10_OAI22X1_28 ( );
FILL FILL_0_CLKBUF1_22 ( );
FILL FILL_1_CLKBUF1_22 ( );
FILL FILL_2_CLKBUF1_22 ( );
FILL FILL_3_CLKBUF1_22 ( );
FILL FILL_4_CLKBUF1_22 ( );
FILL FILL_5_CLKBUF1_22 ( );
FILL FILL_6_CLKBUF1_22 ( );
FILL FILL_7_CLKBUF1_22 ( );
FILL FILL_8_CLKBUF1_22 ( );
FILL FILL_9_CLKBUF1_22 ( );
FILL FILL_10_CLKBUF1_22 ( );
FILL FILL_11_CLKBUF1_22 ( );
FILL FILL_12_CLKBUF1_22 ( );
FILL FILL_13_CLKBUF1_22 ( );
FILL FILL_14_CLKBUF1_22 ( );
FILL FILL_15_CLKBUF1_22 ( );
FILL FILL_16_CLKBUF1_22 ( );
FILL FILL_17_CLKBUF1_22 ( );
FILL FILL_18_CLKBUF1_22 ( );
FILL FILL_19_CLKBUF1_22 ( );
FILL FILL_20_CLKBUF1_22 ( );
FILL FILL_21_CLKBUF1_22 ( );
FILL FILL_0_OAI22X1_30 ( );
FILL FILL_1_OAI22X1_30 ( );
FILL FILL_2_OAI22X1_30 ( );
FILL FILL_3_OAI22X1_30 ( );
FILL FILL_4_OAI22X1_30 ( );
FILL FILL_5_OAI22X1_30 ( );
FILL FILL_6_OAI22X1_30 ( );
FILL FILL_7_OAI22X1_30 ( );
FILL FILL_8_OAI22X1_30 ( );
FILL FILL_9_OAI22X1_30 ( );
FILL FILL_10_OAI22X1_30 ( );
FILL FILL_0_INVX1_303 ( );
FILL FILL_1_INVX1_303 ( );
FILL FILL_2_INVX1_303 ( );
FILL FILL_3_INVX1_303 ( );
FILL FILL_4_INVX1_303 ( );
FILL FILL_0_DFFSR_43 ( );
FILL FILL_1_DFFSR_43 ( );
FILL FILL_2_DFFSR_43 ( );
FILL FILL_3_DFFSR_43 ( );
FILL FILL_4_DFFSR_43 ( );
FILL FILL_5_DFFSR_43 ( );
FILL FILL_6_DFFSR_43 ( );
FILL FILL_7_DFFSR_43 ( );
FILL FILL_8_DFFSR_43 ( );
FILL FILL_9_DFFSR_43 ( );
FILL FILL_10_DFFSR_43 ( );
FILL FILL_11_DFFSR_43 ( );
FILL FILL_12_DFFSR_43 ( );
FILL FILL_13_DFFSR_43 ( );
FILL FILL_14_DFFSR_43 ( );
FILL FILL_15_DFFSR_43 ( );
FILL FILL_16_DFFSR_43 ( );
FILL FILL_17_DFFSR_43 ( );
FILL FILL_18_DFFSR_43 ( );
FILL FILL_19_DFFSR_43 ( );
FILL FILL_20_DFFSR_43 ( );
FILL FILL_21_DFFSR_43 ( );
FILL FILL_22_DFFSR_43 ( );
FILL FILL_23_DFFSR_43 ( );
FILL FILL_24_DFFSR_43 ( );
FILL FILL_25_DFFSR_43 ( );
FILL FILL_26_DFFSR_43 ( );
FILL FILL_27_DFFSR_43 ( );
FILL FILL_28_DFFSR_43 ( );
FILL FILL_29_DFFSR_43 ( );
FILL FILL_30_DFFSR_43 ( );
FILL FILL_31_DFFSR_43 ( );
FILL FILL_32_DFFSR_43 ( );
FILL FILL_33_DFFSR_43 ( );
FILL FILL_34_DFFSR_43 ( );
FILL FILL_35_DFFSR_43 ( );
FILL FILL_36_DFFSR_43 ( );
FILL FILL_37_DFFSR_43 ( );
FILL FILL_38_DFFSR_43 ( );
FILL FILL_39_DFFSR_43 ( );
FILL FILL_40_DFFSR_43 ( );
FILL FILL_41_DFFSR_43 ( );
FILL FILL_42_DFFSR_43 ( );
FILL FILL_43_DFFSR_43 ( );
FILL FILL_44_DFFSR_43 ( );
FILL FILL_45_DFFSR_43 ( );
FILL FILL_46_DFFSR_43 ( );
FILL FILL_47_DFFSR_43 ( );
FILL FILL_48_DFFSR_43 ( );
FILL FILL_49_DFFSR_43 ( );
FILL FILL_50_DFFSR_43 ( );
FILL FILL_0_INVX1_59 ( );
FILL FILL_1_INVX1_59 ( );
FILL FILL_2_INVX1_59 ( );
FILL FILL_3_INVX1_59 ( );
FILL FILL_4_INVX1_59 ( );
FILL FILL_0_OAI21X1_52 ( );
FILL FILL_1_OAI21X1_52 ( );
FILL FILL_2_OAI21X1_52 ( );
FILL FILL_3_OAI21X1_52 ( );
FILL FILL_4_OAI21X1_52 ( );
FILL FILL_5_OAI21X1_52 ( );
FILL FILL_6_OAI21X1_52 ( );
FILL FILL_7_OAI21X1_52 ( );
FILL FILL_8_OAI21X1_52 ( );
FILL FILL_0_INVX1_205 ( );
FILL FILL_1_INVX1_205 ( );
FILL FILL_2_INVX1_205 ( );
FILL FILL_3_INVX1_205 ( );
FILL FILL_0_OAI21X1_170 ( );
FILL FILL_1_OAI21X1_170 ( );
FILL FILL_2_OAI21X1_170 ( );
FILL FILL_3_OAI21X1_170 ( );
FILL FILL_4_OAI21X1_170 ( );
FILL FILL_5_OAI21X1_170 ( );
FILL FILL_6_OAI21X1_170 ( );
FILL FILL_7_OAI21X1_170 ( );
FILL FILL_8_OAI21X1_170 ( );
FILL FILL_9_OAI21X1_170 ( );
FILL FILL_0_CLKBUF1_17 ( );
FILL FILL_1_CLKBUF1_17 ( );
FILL FILL_2_CLKBUF1_17 ( );
FILL FILL_3_CLKBUF1_17 ( );
FILL FILL_4_CLKBUF1_17 ( );
FILL FILL_5_CLKBUF1_17 ( );
FILL FILL_6_CLKBUF1_17 ( );
FILL FILL_7_CLKBUF1_17 ( );
FILL FILL_8_CLKBUF1_17 ( );
FILL FILL_9_CLKBUF1_17 ( );
FILL FILL_10_CLKBUF1_17 ( );
FILL FILL_11_CLKBUF1_17 ( );
FILL FILL_12_CLKBUF1_17 ( );
FILL FILL_13_CLKBUF1_17 ( );
FILL FILL_14_CLKBUF1_17 ( );
FILL FILL_15_CLKBUF1_17 ( );
FILL FILL_16_CLKBUF1_17 ( );
FILL FILL_17_CLKBUF1_17 ( );
FILL FILL_18_CLKBUF1_17 ( );
FILL FILL_19_CLKBUF1_17 ( );
FILL FILL_20_CLKBUF1_17 ( );
FILL FILL_0_NOR2X1_3 ( );
FILL FILL_1_NOR2X1_3 ( );
FILL FILL_2_NOR2X1_3 ( );
FILL FILL_3_NOR2X1_3 ( );
FILL FILL_4_NOR2X1_3 ( );
FILL FILL_5_NOR2X1_3 ( );
FILL FILL_6_NOR2X1_3 ( );
FILL FILL_0_OAI21X1_178 ( );
FILL FILL_1_OAI21X1_178 ( );
FILL FILL_2_OAI21X1_178 ( );
FILL FILL_3_OAI21X1_178 ( );
FILL FILL_4_OAI21X1_178 ( );
FILL FILL_5_OAI21X1_178 ( );
FILL FILL_6_OAI21X1_178 ( );
FILL FILL_7_OAI21X1_178 ( );
FILL FILL_8_OAI21X1_178 ( );
FILL FILL_0_NAND2X1_176 ( );
FILL FILL_1_NAND2X1_176 ( );
FILL FILL_2_NAND2X1_176 ( );
FILL FILL_3_NAND2X1_176 ( );
FILL FILL_4_NAND2X1_176 ( );
FILL FILL_5_NAND2X1_176 ( );
FILL FILL_6_NAND2X1_176 ( );
FILL FILL_0_NAND3X1_1 ( );
FILL FILL_1_NAND3X1_1 ( );
FILL FILL_2_NAND3X1_1 ( );
FILL FILL_3_NAND3X1_1 ( );
FILL FILL_4_NAND3X1_1 ( );
FILL FILL_5_NAND3X1_1 ( );
FILL FILL_6_NAND3X1_1 ( );
FILL FILL_7_NAND3X1_1 ( );
FILL FILL_8_NAND3X1_1 ( );
FILL FILL_0_INVX1_217 ( );
FILL FILL_1_INVX1_217 ( );
FILL FILL_2_INVX1_217 ( );
FILL FILL_3_INVX1_217 ( );
FILL FILL_4_INVX1_217 ( );
FILL FILL_0_NAND3X1_13 ( );
FILL FILL_1_NAND3X1_13 ( );
FILL FILL_2_NAND3X1_13 ( );
FILL FILL_3_NAND3X1_13 ( );
FILL FILL_4_NAND3X1_13 ( );
FILL FILL_5_NAND3X1_13 ( );
FILL FILL_6_NAND3X1_13 ( );
FILL FILL_7_NAND3X1_13 ( );
FILL FILL_8_NAND3X1_13 ( );
FILL FILL_0_AOI22X1_4 ( );
FILL FILL_1_AOI22X1_4 ( );
FILL FILL_2_AOI22X1_4 ( );
FILL FILL_3_AOI22X1_4 ( );
FILL FILL_4_AOI22X1_4 ( );
FILL FILL_5_AOI22X1_4 ( );
FILL FILL_6_AOI22X1_4 ( );
FILL FILL_7_AOI22X1_4 ( );
FILL FILL_8_AOI22X1_4 ( );
FILL FILL_9_AOI22X1_4 ( );
FILL FILL_10_AOI22X1_4 ( );
FILL FILL_11_AOI22X1_4 ( );
FILL FILL_0_OAI21X1_196 ( );
FILL FILL_1_OAI21X1_196 ( );
FILL FILL_2_OAI21X1_196 ( );
FILL FILL_3_OAI21X1_196 ( );
FILL FILL_4_OAI21X1_196 ( );
FILL FILL_5_OAI21X1_196 ( );
FILL FILL_6_OAI21X1_196 ( );
FILL FILL_7_OAI21X1_196 ( );
FILL FILL_8_OAI21X1_196 ( );
FILL FILL_0_NAND3X1_84 ( );
FILL FILL_1_NAND3X1_84 ( );
FILL FILL_2_NAND3X1_84 ( );
FILL FILL_3_NAND3X1_84 ( );
FILL FILL_4_NAND3X1_84 ( );
FILL FILL_5_NAND3X1_84 ( );
FILL FILL_6_NAND3X1_84 ( );
FILL FILL_7_NAND3X1_84 ( );
FILL FILL_8_NAND3X1_84 ( );
FILL FILL_0_AOI21X1_35 ( );
FILL FILL_1_AOI21X1_35 ( );
FILL FILL_2_AOI21X1_35 ( );
FILL FILL_3_AOI21X1_35 ( );
FILL FILL_4_AOI21X1_35 ( );
FILL FILL_5_AOI21X1_35 ( );
FILL FILL_6_AOI21X1_35 ( );
FILL FILL_7_AOI21X1_35 ( );
FILL FILL_8_AOI21X1_35 ( );
FILL FILL_9_AOI21X1_35 ( );
FILL FILL_0_AOI21X1_34 ( );
FILL FILL_1_AOI21X1_34 ( );
FILL FILL_2_AOI21X1_34 ( );
FILL FILL_3_AOI21X1_34 ( );
FILL FILL_4_AOI21X1_34 ( );
FILL FILL_5_AOI21X1_34 ( );
FILL FILL_6_AOI21X1_34 ( );
FILL FILL_7_AOI21X1_34 ( );
FILL FILL_8_AOI21X1_34 ( );
FILL FILL_0_INVX1_250 ( );
FILL FILL_1_INVX1_250 ( );
FILL FILL_2_INVX1_250 ( );
FILL FILL_3_INVX1_250 ( );
FILL FILL_4_INVX1_250 ( );
FILL FILL_0_CLKBUF1_1 ( );
FILL FILL_1_CLKBUF1_1 ( );
FILL FILL_2_CLKBUF1_1 ( );
FILL FILL_3_CLKBUF1_1 ( );
FILL FILL_4_CLKBUF1_1 ( );
FILL FILL_5_CLKBUF1_1 ( );
FILL FILL_6_CLKBUF1_1 ( );
FILL FILL_7_CLKBUF1_1 ( );
FILL FILL_8_CLKBUF1_1 ( );
FILL FILL_9_CLKBUF1_1 ( );
FILL FILL_10_CLKBUF1_1 ( );
FILL FILL_11_CLKBUF1_1 ( );
FILL FILL_12_CLKBUF1_1 ( );
FILL FILL_13_CLKBUF1_1 ( );
FILL FILL_14_CLKBUF1_1 ( );
FILL FILL_15_CLKBUF1_1 ( );
FILL FILL_16_CLKBUF1_1 ( );
FILL FILL_17_CLKBUF1_1 ( );
FILL FILL_18_CLKBUF1_1 ( );
FILL FILL_19_CLKBUF1_1 ( );
FILL FILL_20_CLKBUF1_1 ( );
FILL FILL_0_OAI21X1_128 ( );
FILL FILL_1_OAI21X1_128 ( );
FILL FILL_2_OAI21X1_128 ( );
FILL FILL_3_OAI21X1_128 ( );
FILL FILL_4_OAI21X1_128 ( );
FILL FILL_5_OAI21X1_128 ( );
FILL FILL_6_OAI21X1_128 ( );
FILL FILL_7_OAI21X1_128 ( );
FILL FILL_8_OAI21X1_128 ( );
FILL FILL_0_INVX1_144 ( );
FILL FILL_1_INVX1_144 ( );
FILL FILL_2_INVX1_144 ( );
FILL FILL_3_INVX1_144 ( );
FILL FILL_4_INVX1_144 ( );
FILL FILL_0_OAI22X1_62 ( );
FILL FILL_1_OAI22X1_62 ( );
FILL FILL_2_OAI22X1_62 ( );
FILL FILL_3_OAI22X1_62 ( );
FILL FILL_4_OAI22X1_62 ( );
FILL FILL_5_OAI22X1_62 ( );
FILL FILL_6_OAI22X1_62 ( );
FILL FILL_7_OAI22X1_62 ( );
FILL FILL_8_OAI22X1_62 ( );
FILL FILL_9_OAI22X1_62 ( );
FILL FILL_10_OAI22X1_62 ( );
FILL FILL_11_OAI22X1_62 ( );
FILL FILL_0_INVX1_344 ( );
FILL FILL_1_INVX1_344 ( );
FILL FILL_2_INVX1_344 ( );
FILL FILL_3_INVX1_344 ( );
FILL FILL_4_INVX1_344 ( );
FILL FILL_0_OAI22X1_43 ( );
FILL FILL_1_OAI22X1_43 ( );
FILL FILL_2_OAI22X1_43 ( );
FILL FILL_3_OAI22X1_43 ( );
FILL FILL_4_OAI22X1_43 ( );
FILL FILL_5_OAI22X1_43 ( );
FILL FILL_6_OAI22X1_43 ( );
FILL FILL_7_OAI22X1_43 ( );
FILL FILL_8_OAI22X1_43 ( );
FILL FILL_9_OAI22X1_43 ( );
FILL FILL_10_OAI22X1_43 ( );
FILL FILL_11_OAI22X1_43 ( );
FILL FILL_0_OAI21X1_108 ( );
FILL FILL_1_OAI21X1_108 ( );
FILL FILL_2_OAI21X1_108 ( );
FILL FILL_3_OAI21X1_108 ( );
FILL FILL_4_OAI21X1_108 ( );
FILL FILL_5_OAI21X1_108 ( );
FILL FILL_6_OAI21X1_108 ( );
FILL FILL_7_OAI21X1_108 ( );
FILL FILL_8_OAI21X1_108 ( );
FILL FILL_0_NAND2X1_83 ( );
FILL FILL_1_NAND2X1_83 ( );
FILL FILL_2_NAND2X1_83 ( );
FILL FILL_3_NAND2X1_83 ( );
FILL FILL_4_NAND2X1_83 ( );
FILL FILL_5_NAND2X1_83 ( );
FILL FILL_6_NAND2X1_83 ( );
FILL FILL_0_DFFSR_150 ( );
FILL FILL_1_DFFSR_150 ( );
FILL FILL_2_DFFSR_150 ( );
FILL FILL_3_DFFSR_150 ( );
FILL FILL_4_DFFSR_150 ( );
FILL FILL_5_DFFSR_150 ( );
FILL FILL_6_DFFSR_150 ( );
FILL FILL_7_DFFSR_150 ( );
FILL FILL_8_DFFSR_150 ( );
FILL FILL_9_DFFSR_150 ( );
FILL FILL_10_DFFSR_150 ( );
FILL FILL_11_DFFSR_150 ( );
FILL FILL_12_DFFSR_150 ( );
FILL FILL_13_DFFSR_150 ( );
FILL FILL_14_DFFSR_150 ( );
FILL FILL_15_DFFSR_150 ( );
FILL FILL_16_DFFSR_150 ( );
FILL FILL_17_DFFSR_150 ( );
FILL FILL_18_DFFSR_150 ( );
FILL FILL_19_DFFSR_150 ( );
FILL FILL_20_DFFSR_150 ( );
FILL FILL_21_DFFSR_150 ( );
FILL FILL_22_DFFSR_150 ( );
FILL FILL_23_DFFSR_150 ( );
FILL FILL_24_DFFSR_150 ( );
FILL FILL_25_DFFSR_150 ( );
FILL FILL_26_DFFSR_150 ( );
FILL FILL_27_DFFSR_150 ( );
FILL FILL_28_DFFSR_150 ( );
FILL FILL_29_DFFSR_150 ( );
FILL FILL_30_DFFSR_150 ( );
FILL FILL_31_DFFSR_150 ( );
FILL FILL_32_DFFSR_150 ( );
FILL FILL_33_DFFSR_150 ( );
FILL FILL_34_DFFSR_150 ( );
FILL FILL_35_DFFSR_150 ( );
FILL FILL_36_DFFSR_150 ( );
FILL FILL_37_DFFSR_150 ( );
FILL FILL_38_DFFSR_150 ( );
FILL FILL_39_DFFSR_150 ( );
FILL FILL_40_DFFSR_150 ( );
FILL FILL_41_DFFSR_150 ( );
FILL FILL_42_DFFSR_150 ( );
FILL FILL_43_DFFSR_150 ( );
FILL FILL_44_DFFSR_150 ( );
FILL FILL_45_DFFSR_150 ( );
FILL FILL_46_DFFSR_150 ( );
FILL FILL_47_DFFSR_150 ( );
FILL FILL_48_DFFSR_150 ( );
FILL FILL_49_DFFSR_150 ( );
FILL FILL_50_DFFSR_150 ( );
FILL FILL_0_DFFSR_143 ( );
FILL FILL_1_DFFSR_143 ( );
FILL FILL_2_DFFSR_143 ( );
FILL FILL_3_DFFSR_143 ( );
FILL FILL_4_DFFSR_143 ( );
FILL FILL_5_DFFSR_143 ( );
FILL FILL_6_DFFSR_143 ( );
FILL FILL_7_DFFSR_143 ( );
FILL FILL_8_DFFSR_143 ( );
FILL FILL_9_DFFSR_143 ( );
FILL FILL_10_DFFSR_143 ( );
FILL FILL_11_DFFSR_143 ( );
FILL FILL_12_DFFSR_143 ( );
FILL FILL_13_DFFSR_143 ( );
FILL FILL_14_DFFSR_143 ( );
FILL FILL_15_DFFSR_143 ( );
FILL FILL_16_DFFSR_143 ( );
FILL FILL_17_DFFSR_143 ( );
FILL FILL_18_DFFSR_143 ( );
FILL FILL_19_DFFSR_143 ( );
FILL FILL_20_DFFSR_143 ( );
FILL FILL_21_DFFSR_143 ( );
FILL FILL_22_DFFSR_143 ( );
FILL FILL_23_DFFSR_143 ( );
FILL FILL_24_DFFSR_143 ( );
FILL FILL_25_DFFSR_143 ( );
FILL FILL_26_DFFSR_143 ( );
FILL FILL_27_DFFSR_143 ( );
FILL FILL_28_DFFSR_143 ( );
FILL FILL_29_DFFSR_143 ( );
FILL FILL_30_DFFSR_143 ( );
FILL FILL_31_DFFSR_143 ( );
FILL FILL_32_DFFSR_143 ( );
FILL FILL_33_DFFSR_143 ( );
FILL FILL_34_DFFSR_143 ( );
FILL FILL_35_DFFSR_143 ( );
FILL FILL_36_DFFSR_143 ( );
FILL FILL_37_DFFSR_143 ( );
FILL FILL_38_DFFSR_143 ( );
FILL FILL_39_DFFSR_143 ( );
FILL FILL_40_DFFSR_143 ( );
FILL FILL_41_DFFSR_143 ( );
FILL FILL_42_DFFSR_143 ( );
FILL FILL_43_DFFSR_143 ( );
FILL FILL_44_DFFSR_143 ( );
FILL FILL_45_DFFSR_143 ( );
FILL FILL_46_DFFSR_143 ( );
FILL FILL_47_DFFSR_143 ( );
FILL FILL_48_DFFSR_143 ( );
FILL FILL_49_DFFSR_143 ( );
FILL FILL_50_DFFSR_143 ( );
FILL FILL_0_OAI21X1_22 ( );
FILL FILL_1_OAI21X1_22 ( );
FILL FILL_2_OAI21X1_22 ( );
FILL FILL_3_OAI21X1_22 ( );
FILL FILL_4_OAI21X1_22 ( );
FILL FILL_5_OAI21X1_22 ( );
FILL FILL_6_OAI21X1_22 ( );
FILL FILL_7_OAI21X1_22 ( );
FILL FILL_8_OAI21X1_22 ( );
FILL FILL_0_INVX1_25 ( );
FILL FILL_1_INVX1_25 ( );
FILL FILL_2_INVX1_25 ( );
FILL FILL_3_INVX1_25 ( );
FILL FILL_4_INVX1_25 ( );
FILL FILL_0_NAND2X1_63 ( );
FILL FILL_1_NAND2X1_63 ( );
FILL FILL_2_NAND2X1_63 ( );
FILL FILL_3_NAND2X1_63 ( );
FILL FILL_4_NAND2X1_63 ( );
FILL FILL_5_NAND2X1_63 ( );
FILL FILL_6_NAND2X1_63 ( );
FILL FILL_0_INVX1_305 ( );
FILL FILL_1_INVX1_305 ( );
FILL FILL_2_INVX1_305 ( );
FILL FILL_3_INVX1_305 ( );
FILL FILL_4_INVX1_305 ( );
FILL FILL_0_OAI22X1_25 ( );
FILL FILL_1_OAI22X1_25 ( );
FILL FILL_2_OAI22X1_25 ( );
FILL FILL_3_OAI22X1_25 ( );
FILL FILL_4_OAI22X1_25 ( );
FILL FILL_5_OAI22X1_25 ( );
FILL FILL_6_OAI22X1_25 ( );
FILL FILL_7_OAI22X1_25 ( );
FILL FILL_8_OAI22X1_25 ( );
FILL FILL_9_OAI22X1_25 ( );
FILL FILL_10_OAI22X1_25 ( );
FILL FILL_0_NOR2X1_22 ( );
FILL FILL_1_NOR2X1_22 ( );
FILL FILL_2_NOR2X1_22 ( );
FILL FILL_3_NOR2X1_22 ( );
FILL FILL_4_NOR2X1_22 ( );
FILL FILL_5_NOR2X1_22 ( );
FILL FILL_6_NOR2X1_22 ( );
FILL FILL_0_INVX1_315 ( );
FILL FILL_1_INVX1_315 ( );
FILL FILL_2_INVX1_315 ( );
FILL FILL_3_INVX1_315 ( );
FILL FILL_4_INVX1_315 ( );
FILL FILL_0_NAND2X1_46 ( );
FILL FILL_1_NAND2X1_46 ( );
FILL FILL_2_NAND2X1_46 ( );
FILL FILL_3_NAND2X1_46 ( );
FILL FILL_4_NAND2X1_46 ( );
FILL FILL_5_NAND2X1_46 ( );
FILL FILL_6_NAND2X1_46 ( );
FILL FILL_0_OAI22X1_20 ( );
FILL FILL_1_OAI22X1_20 ( );
FILL FILL_2_OAI22X1_20 ( );
FILL FILL_3_OAI22X1_20 ( );
FILL FILL_4_OAI22X1_20 ( );
FILL FILL_5_OAI22X1_20 ( );
FILL FILL_6_OAI22X1_20 ( );
FILL FILL_7_OAI22X1_20 ( );
FILL FILL_8_OAI22X1_20 ( );
FILL FILL_9_OAI22X1_20 ( );
FILL FILL_10_OAI22X1_20 ( );
FILL FILL_0_INVX1_296 ( );
FILL FILL_1_INVX1_296 ( );
FILL FILL_2_INVX1_296 ( );
FILL FILL_3_INVX1_296 ( );
FILL FILL_4_INVX1_296 ( );
FILL FILL_0_INVX1_291 ( );
FILL FILL_1_INVX1_291 ( );
FILL FILL_2_INVX1_291 ( );
FILL FILL_3_INVX1_291 ( );
FILL FILL_4_INVX1_291 ( );
FILL FILL_0_OAI22X1_17 ( );
FILL FILL_1_OAI22X1_17 ( );
FILL FILL_2_OAI22X1_17 ( );
FILL FILL_3_OAI22X1_17 ( );
FILL FILL_4_OAI22X1_17 ( );
FILL FILL_5_OAI22X1_17 ( );
FILL FILL_6_OAI22X1_17 ( );
FILL FILL_7_OAI22X1_17 ( );
FILL FILL_8_OAI22X1_17 ( );
FILL FILL_9_OAI22X1_17 ( );
FILL FILL_10_OAI22X1_17 ( );
FILL FILL_0_DFFSR_25 ( );
FILL FILL_1_DFFSR_25 ( );
FILL FILL_2_DFFSR_25 ( );
FILL FILL_3_DFFSR_25 ( );
FILL FILL_4_DFFSR_25 ( );
FILL FILL_5_DFFSR_25 ( );
FILL FILL_6_DFFSR_25 ( );
FILL FILL_7_DFFSR_25 ( );
FILL FILL_8_DFFSR_25 ( );
FILL FILL_9_DFFSR_25 ( );
FILL FILL_10_DFFSR_25 ( );
FILL FILL_11_DFFSR_25 ( );
FILL FILL_12_DFFSR_25 ( );
FILL FILL_13_DFFSR_25 ( );
FILL FILL_14_DFFSR_25 ( );
FILL FILL_15_DFFSR_25 ( );
FILL FILL_16_DFFSR_25 ( );
FILL FILL_17_DFFSR_25 ( );
FILL FILL_18_DFFSR_25 ( );
FILL FILL_19_DFFSR_25 ( );
FILL FILL_20_DFFSR_25 ( );
FILL FILL_21_DFFSR_25 ( );
FILL FILL_22_DFFSR_25 ( );
FILL FILL_23_DFFSR_25 ( );
FILL FILL_24_DFFSR_25 ( );
FILL FILL_25_DFFSR_25 ( );
FILL FILL_26_DFFSR_25 ( );
FILL FILL_27_DFFSR_25 ( );
FILL FILL_28_DFFSR_25 ( );
FILL FILL_29_DFFSR_25 ( );
FILL FILL_30_DFFSR_25 ( );
FILL FILL_31_DFFSR_25 ( );
FILL FILL_32_DFFSR_25 ( );
FILL FILL_33_DFFSR_25 ( );
FILL FILL_34_DFFSR_25 ( );
FILL FILL_35_DFFSR_25 ( );
FILL FILL_36_DFFSR_25 ( );
FILL FILL_37_DFFSR_25 ( );
FILL FILL_38_DFFSR_25 ( );
FILL FILL_39_DFFSR_25 ( );
FILL FILL_40_DFFSR_25 ( );
FILL FILL_41_DFFSR_25 ( );
FILL FILL_42_DFFSR_25 ( );
FILL FILL_43_DFFSR_25 ( );
FILL FILL_44_DFFSR_25 ( );
FILL FILL_45_DFFSR_25 ( );
FILL FILL_46_DFFSR_25 ( );
FILL FILL_47_DFFSR_25 ( );
FILL FILL_48_DFFSR_25 ( );
FILL FILL_49_DFFSR_25 ( );
FILL FILL_50_DFFSR_25 ( );
FILL FILL_0_INVX1_50 ( );
FILL FILL_1_INVX1_50 ( );
FILL FILL_2_INVX1_50 ( );
FILL FILL_3_INVX1_50 ( );
FILL FILL_4_INVX1_50 ( );
FILL FILL_0_NAND2X1_178 ( );
FILL FILL_1_NAND2X1_178 ( );
FILL FILL_2_NAND2X1_178 ( );
FILL FILL_3_NAND2X1_178 ( );
FILL FILL_4_NAND2X1_178 ( );
FILL FILL_5_NAND2X1_178 ( );
FILL FILL_6_NAND2X1_178 ( );
FILL FILL_0_CLKBUF1_18 ( );
FILL FILL_1_CLKBUF1_18 ( );
FILL FILL_2_CLKBUF1_18 ( );
FILL FILL_3_CLKBUF1_18 ( );
FILL FILL_4_CLKBUF1_18 ( );
FILL FILL_5_CLKBUF1_18 ( );
FILL FILL_6_CLKBUF1_18 ( );
FILL FILL_7_CLKBUF1_18 ( );
FILL FILL_8_CLKBUF1_18 ( );
FILL FILL_9_CLKBUF1_18 ( );
FILL FILL_10_CLKBUF1_18 ( );
FILL FILL_11_CLKBUF1_18 ( );
FILL FILL_12_CLKBUF1_18 ( );
FILL FILL_13_CLKBUF1_18 ( );
FILL FILL_14_CLKBUF1_18 ( );
FILL FILL_15_CLKBUF1_18 ( );
FILL FILL_16_CLKBUF1_18 ( );
FILL FILL_17_CLKBUF1_18 ( );
FILL FILL_18_CLKBUF1_18 ( );
FILL FILL_19_CLKBUF1_18 ( );
FILL FILL_20_CLKBUF1_18 ( );
FILL FILL_0_NAND2X1_182 ( );
FILL FILL_1_NAND2X1_182 ( );
FILL FILL_2_NAND2X1_182 ( );
FILL FILL_3_NAND2X1_182 ( );
FILL FILL_4_NAND2X1_182 ( );
FILL FILL_5_NAND2X1_182 ( );
FILL FILL_6_NAND2X1_182 ( );
FILL FILL_0_NAND2X1_162 ( );
FILL FILL_1_NAND2X1_162 ( );
FILL FILL_2_NAND2X1_162 ( );
FILL FILL_3_NAND2X1_162 ( );
FILL FILL_4_NAND2X1_162 ( );
FILL FILL_5_NAND2X1_162 ( );
FILL FILL_6_NAND2X1_162 ( );
FILL FILL_0_OAI21X1_176 ( );
FILL FILL_1_OAI21X1_176 ( );
FILL FILL_2_OAI21X1_176 ( );
FILL FILL_3_OAI21X1_176 ( );
FILL FILL_4_OAI21X1_176 ( );
FILL FILL_5_OAI21X1_176 ( );
FILL FILL_6_OAI21X1_176 ( );
FILL FILL_7_OAI21X1_176 ( );
FILL FILL_8_OAI21X1_176 ( );
FILL FILL_9_OAI21X1_176 ( );
FILL FILL_0_NAND2X1_179 ( );
FILL FILL_1_NAND2X1_179 ( );
FILL FILL_2_NAND2X1_179 ( );
FILL FILL_3_NAND2X1_179 ( );
FILL FILL_4_NAND2X1_179 ( );
FILL FILL_5_NAND2X1_179 ( );
FILL FILL_6_NAND2X1_179 ( );
FILL FILL_0_BUFX2_4 ( );
FILL FILL_1_BUFX2_4 ( );
FILL FILL_2_BUFX2_4 ( );
FILL FILL_3_BUFX2_4 ( );
FILL FILL_4_BUFX2_4 ( );
FILL FILL_5_BUFX2_4 ( );
FILL FILL_6_BUFX2_4 ( );
FILL FILL_0_NAND2X1_165 ( );
FILL FILL_1_NAND2X1_165 ( );
FILL FILL_2_NAND2X1_165 ( );
FILL FILL_3_NAND2X1_165 ( );
FILL FILL_4_NAND2X1_165 ( );
FILL FILL_5_NAND2X1_165 ( );
FILL FILL_6_NAND2X1_165 ( );
FILL FILL_0_INVX1_201 ( );
FILL FILL_1_INVX1_201 ( );
FILL FILL_2_INVX1_201 ( );
FILL FILL_3_INVX1_201 ( );
FILL FILL_4_INVX1_201 ( );
FILL FILL_0_NAND3X1_59 ( );
FILL FILL_1_NAND3X1_59 ( );
FILL FILL_2_NAND3X1_59 ( );
FILL FILL_3_NAND3X1_59 ( );
FILL FILL_4_NAND3X1_59 ( );
FILL FILL_5_NAND3X1_59 ( );
FILL FILL_6_NAND3X1_59 ( );
FILL FILL_7_NAND3X1_59 ( );
FILL FILL_8_NAND3X1_59 ( );
FILL FILL_0_OAI21X1_167 ( );
FILL FILL_1_OAI21X1_167 ( );
FILL FILL_2_OAI21X1_167 ( );
FILL FILL_3_OAI21X1_167 ( );
FILL FILL_4_OAI21X1_167 ( );
FILL FILL_5_OAI21X1_167 ( );
FILL FILL_6_OAI21X1_167 ( );
FILL FILL_7_OAI21X1_167 ( );
FILL FILL_8_OAI21X1_167 ( );
FILL FILL_0_AOI21X1_36 ( );
FILL FILL_1_AOI21X1_36 ( );
FILL FILL_2_AOI21X1_36 ( );
FILL FILL_3_AOI21X1_36 ( );
FILL FILL_4_AOI21X1_36 ( );
FILL FILL_5_AOI21X1_36 ( );
FILL FILL_6_AOI21X1_36 ( );
FILL FILL_7_AOI21X1_36 ( );
FILL FILL_8_AOI21X1_36 ( );
FILL FILL_0_AOI21X1_37 ( );
FILL FILL_1_AOI21X1_37 ( );
FILL FILL_2_AOI21X1_37 ( );
FILL FILL_3_AOI21X1_37 ( );
FILL FILL_4_AOI21X1_37 ( );
FILL FILL_5_AOI21X1_37 ( );
FILL FILL_6_AOI21X1_37 ( );
FILL FILL_7_AOI21X1_37 ( );
FILL FILL_8_AOI21X1_37 ( );
FILL FILL_9_AOI21X1_37 ( );
FILL FILL_0_CLKBUF1_4 ( );
FILL FILL_1_CLKBUF1_4 ( );
FILL FILL_2_CLKBUF1_4 ( );
FILL FILL_3_CLKBUF1_4 ( );
FILL FILL_4_CLKBUF1_4 ( );
FILL FILL_5_CLKBUF1_4 ( );
FILL FILL_6_CLKBUF1_4 ( );
FILL FILL_7_CLKBUF1_4 ( );
FILL FILL_8_CLKBUF1_4 ( );
FILL FILL_9_CLKBUF1_4 ( );
FILL FILL_10_CLKBUF1_4 ( );
FILL FILL_11_CLKBUF1_4 ( );
FILL FILL_12_CLKBUF1_4 ( );
FILL FILL_13_CLKBUF1_4 ( );
FILL FILL_14_CLKBUF1_4 ( );
FILL FILL_15_CLKBUF1_4 ( );
FILL FILL_16_CLKBUF1_4 ( );
FILL FILL_17_CLKBUF1_4 ( );
FILL FILL_18_CLKBUF1_4 ( );
FILL FILL_19_CLKBUF1_4 ( );
FILL FILL_0_INVX1_385 ( );
FILL FILL_1_INVX1_385 ( );
FILL FILL_2_INVX1_385 ( );
FILL FILL_3_INVX1_385 ( );
FILL FILL_0_INVX1_80 ( );
FILL FILL_1_INVX1_80 ( );
FILL FILL_2_INVX1_80 ( );
FILL FILL_3_INVX1_80 ( );
FILL FILL_4_INVX1_80 ( );
FILL FILL_0_OAI21X1_71 ( );
FILL FILL_1_OAI21X1_71 ( );
FILL FILL_2_OAI21X1_71 ( );
FILL FILL_3_OAI21X1_71 ( );
FILL FILL_4_OAI21X1_71 ( );
FILL FILL_5_OAI21X1_71 ( );
FILL FILL_6_OAI21X1_71 ( );
FILL FILL_7_OAI21X1_71 ( );
FILL FILL_8_OAI21X1_71 ( );
FILL FILL_0_OAI22X1_63 ( );
FILL FILL_1_OAI22X1_63 ( );
FILL FILL_2_OAI22X1_63 ( );
FILL FILL_3_OAI22X1_63 ( );
FILL FILL_4_OAI22X1_63 ( );
FILL FILL_5_OAI22X1_63 ( );
FILL FILL_6_OAI22X1_63 ( );
FILL FILL_7_OAI22X1_63 ( );
FILL FILL_8_OAI22X1_63 ( );
FILL FILL_9_OAI22X1_63 ( );
FILL FILL_10_OAI22X1_63 ( );
FILL FILL_11_OAI22X1_63 ( );
FILL FILL_0_NOR2X1_41 ( );
FILL FILL_1_NOR2X1_41 ( );
FILL FILL_2_NOR2X1_41 ( );
FILL FILL_3_NOR2X1_41 ( );
FILL FILL_4_NOR2X1_41 ( );
FILL FILL_5_NOR2X1_41 ( );
FILL FILL_6_NOR2X1_41 ( );
FILL FILL_0_NOR2X1_40 ( );
FILL FILL_1_NOR2X1_40 ( );
FILL FILL_2_NOR2X1_40 ( );
FILL FILL_3_NOR2X1_40 ( );
FILL FILL_4_NOR2X1_40 ( );
FILL FILL_5_NOR2X1_40 ( );
FILL FILL_6_NOR2X1_40 ( );
FILL FILL_0_NAND2X1_248 ( );
FILL FILL_1_NAND2X1_248 ( );
FILL FILL_2_NAND2X1_248 ( );
FILL FILL_3_NAND2X1_248 ( );
FILL FILL_4_NAND2X1_248 ( );
FILL FILL_5_NAND2X1_248 ( );
FILL FILL_6_NAND2X1_248 ( );
FILL FILL_0_NAND2X1_71 ( );
FILL FILL_1_NAND2X1_71 ( );
FILL FILL_2_NAND2X1_71 ( );
FILL FILL_3_NAND2X1_71 ( );
FILL FILL_4_NAND2X1_71 ( );
FILL FILL_5_NAND2X1_71 ( );
FILL FILL_6_NAND2X1_71 ( );
FILL FILL_0_OAI22X1_54 ( );
FILL FILL_1_OAI22X1_54 ( );
FILL FILL_2_OAI22X1_54 ( );
FILL FILL_3_OAI22X1_54 ( );
FILL FILL_4_OAI22X1_54 ( );
FILL FILL_5_OAI22X1_54 ( );
FILL FILL_6_OAI22X1_54 ( );
FILL FILL_7_OAI22X1_54 ( );
FILL FILL_8_OAI22X1_54 ( );
FILL FILL_9_OAI22X1_54 ( );
FILL FILL_10_OAI22X1_54 ( );
FILL FILL_11_OAI22X1_54 ( );
FILL FILL_0_NOR2X1_36 ( );
FILL FILL_1_NOR2X1_36 ( );
FILL FILL_2_NOR2X1_36 ( );
FILL FILL_3_NOR2X1_36 ( );
FILL FILL_4_NOR2X1_36 ( );
FILL FILL_5_NOR2X1_36 ( );
FILL FILL_6_NOR2X1_36 ( );
FILL FILL_0_NAND2X1_68 ( );
FILL FILL_1_NAND2X1_68 ( );
FILL FILL_2_NAND2X1_68 ( );
FILL FILL_3_NAND2X1_68 ( );
FILL FILL_4_NAND2X1_68 ( );
FILL FILL_5_NAND2X1_68 ( );
FILL FILL_6_NAND2X1_68 ( );
FILL FILL_0_NAND2X1_143 ( );
FILL FILL_1_NAND2X1_143 ( );
FILL FILL_2_NAND2X1_143 ( );
FILL FILL_3_NAND2X1_143 ( );
FILL FILL_4_NAND2X1_143 ( );
FILL FILL_5_NAND2X1_143 ( );
FILL FILL_6_NAND2X1_143 ( );
FILL FILL_0_OAI21X1_143 ( );
FILL FILL_1_OAI21X1_143 ( );
FILL FILL_2_OAI21X1_143 ( );
FILL FILL_3_OAI21X1_143 ( );
FILL FILL_4_OAI21X1_143 ( );
FILL FILL_5_OAI21X1_143 ( );
FILL FILL_6_OAI21X1_143 ( );
FILL FILL_7_OAI21X1_143 ( );
FILL FILL_8_OAI21X1_143 ( );
FILL FILL_0_INVX1_161 ( );
FILL FILL_1_INVX1_161 ( );
FILL FILL_2_INVX1_161 ( );
FILL FILL_3_INVX1_161 ( );
FILL FILL_4_INVX1_161 ( );
FILL FILL_0_BUFX2_8 ( );
FILL FILL_1_BUFX2_8 ( );
FILL FILL_2_BUFX2_8 ( );
FILL FILL_3_BUFX2_8 ( );
FILL FILL_4_BUFX2_8 ( );
FILL FILL_5_BUFX2_8 ( );
FILL FILL_6_BUFX2_8 ( );
FILL FILL_0_DFFSR_22 ( );
FILL FILL_1_DFFSR_22 ( );
FILL FILL_2_DFFSR_22 ( );
FILL FILL_3_DFFSR_22 ( );
FILL FILL_4_DFFSR_22 ( );
FILL FILL_5_DFFSR_22 ( );
FILL FILL_6_DFFSR_22 ( );
FILL FILL_7_DFFSR_22 ( );
FILL FILL_8_DFFSR_22 ( );
FILL FILL_9_DFFSR_22 ( );
FILL FILL_10_DFFSR_22 ( );
FILL FILL_11_DFFSR_22 ( );
FILL FILL_12_DFFSR_22 ( );
FILL FILL_13_DFFSR_22 ( );
FILL FILL_14_DFFSR_22 ( );
FILL FILL_15_DFFSR_22 ( );
FILL FILL_16_DFFSR_22 ( );
FILL FILL_17_DFFSR_22 ( );
FILL FILL_18_DFFSR_22 ( );
FILL FILL_19_DFFSR_22 ( );
FILL FILL_20_DFFSR_22 ( );
FILL FILL_21_DFFSR_22 ( );
FILL FILL_22_DFFSR_22 ( );
FILL FILL_23_DFFSR_22 ( );
FILL FILL_24_DFFSR_22 ( );
FILL FILL_25_DFFSR_22 ( );
FILL FILL_26_DFFSR_22 ( );
FILL FILL_27_DFFSR_22 ( );
FILL FILL_28_DFFSR_22 ( );
FILL FILL_29_DFFSR_22 ( );
FILL FILL_30_DFFSR_22 ( );
FILL FILL_31_DFFSR_22 ( );
FILL FILL_32_DFFSR_22 ( );
FILL FILL_33_DFFSR_22 ( );
FILL FILL_34_DFFSR_22 ( );
FILL FILL_35_DFFSR_22 ( );
FILL FILL_36_DFFSR_22 ( );
FILL FILL_37_DFFSR_22 ( );
FILL FILL_38_DFFSR_22 ( );
FILL FILL_39_DFFSR_22 ( );
FILL FILL_40_DFFSR_22 ( );
FILL FILL_41_DFFSR_22 ( );
FILL FILL_42_DFFSR_22 ( );
FILL FILL_43_DFFSR_22 ( );
FILL FILL_44_DFFSR_22 ( );
FILL FILL_45_DFFSR_22 ( );
FILL FILL_46_DFFSR_22 ( );
FILL FILL_47_DFFSR_22 ( );
FILL FILL_48_DFFSR_22 ( );
FILL FILL_49_DFFSR_22 ( );
FILL FILL_50_DFFSR_22 ( );
FILL FILL_51_DFFSR_22 ( );
FILL FILL_0_NAND2X1_240 ( );
FILL FILL_1_NAND2X1_240 ( );
FILL FILL_2_NAND2X1_240 ( );
FILL FILL_3_NAND2X1_240 ( );
FILL FILL_4_NAND2X1_240 ( );
FILL FILL_5_NAND2X1_240 ( );
FILL FILL_6_NAND2X1_240 ( );
FILL FILL_0_NOR2X1_24 ( );
FILL FILL_1_NOR2X1_24 ( );
FILL FILL_2_NOR2X1_24 ( );
FILL FILL_3_NOR2X1_24 ( );
FILL FILL_4_NOR2X1_24 ( );
FILL FILL_5_NOR2X1_24 ( );
FILL FILL_6_NOR2X1_24 ( );
FILL FILL_0_INVX1_266 ( );
FILL FILL_1_INVX1_266 ( );
FILL FILL_2_INVX1_266 ( );
FILL FILL_3_INVX1_266 ( );
FILL FILL_4_INVX1_266 ( );
FILL FILL_0_NAND3X1_113 ( );
FILL FILL_1_NAND3X1_113 ( );
FILL FILL_2_NAND3X1_113 ( );
FILL FILL_3_NAND3X1_113 ( );
FILL FILL_4_NAND3X1_113 ( );
FILL FILL_5_NAND3X1_113 ( );
FILL FILL_6_NAND3X1_113 ( );
FILL FILL_7_NAND3X1_113 ( );
FILL FILL_8_NAND3X1_113 ( );
FILL FILL_0_NAND3X1_115 ( );
FILL FILL_1_NAND3X1_115 ( );
FILL FILL_2_NAND3X1_115 ( );
FILL FILL_3_NAND3X1_115 ( );
FILL FILL_4_NAND3X1_115 ( );
FILL FILL_5_NAND3X1_115 ( );
FILL FILL_6_NAND3X1_115 ( );
FILL FILL_7_NAND3X1_115 ( );
FILL FILL_8_NAND3X1_115 ( );
FILL FILL_0_NAND2X1_237 ( );
FILL FILL_1_NAND2X1_237 ( );
FILL FILL_2_NAND2X1_237 ( );
FILL FILL_3_NAND2X1_237 ( );
FILL FILL_4_NAND2X1_237 ( );
FILL FILL_5_NAND2X1_237 ( );
FILL FILL_6_NAND2X1_237 ( );
FILL FILL_0_NOR2X1_18 ( );
FILL FILL_1_NOR2X1_18 ( );
FILL FILL_2_NOR2X1_18 ( );
FILL FILL_3_NOR2X1_18 ( );
FILL FILL_4_NOR2X1_18 ( );
FILL FILL_5_NOR2X1_18 ( );
FILL FILL_6_NOR2X1_18 ( );
FILL FILL_0_NOR2X1_19 ( );
FILL FILL_1_NOR2X1_19 ( );
FILL FILL_2_NOR2X1_19 ( );
FILL FILL_3_NOR2X1_19 ( );
FILL FILL_4_NOR2X1_19 ( );
FILL FILL_5_NOR2X1_19 ( );
FILL FILL_6_NOR2X1_19 ( );
FILL FILL_0_NAND2X1_12 ( );
FILL FILL_1_NAND2X1_12 ( );
FILL FILL_2_NAND2X1_12 ( );
FILL FILL_3_NAND2X1_12 ( );
FILL FILL_4_NAND2X1_12 ( );
FILL FILL_5_NAND2X1_12 ( );
FILL FILL_6_NAND2X1_12 ( );
FILL FILL_0_OAI22X1_18 ( );
FILL FILL_1_OAI22X1_18 ( );
FILL FILL_2_OAI22X1_18 ( );
FILL FILL_3_OAI22X1_18 ( );
FILL FILL_4_OAI22X1_18 ( );
FILL FILL_5_OAI22X1_18 ( );
FILL FILL_6_OAI22X1_18 ( );
FILL FILL_7_OAI22X1_18 ( );
FILL FILL_8_OAI22X1_18 ( );
FILL FILL_9_OAI22X1_18 ( );
FILL FILL_10_OAI22X1_18 ( );
FILL FILL_0_OAI21X1_43 ( );
FILL FILL_1_OAI21X1_43 ( );
FILL FILL_2_OAI21X1_43 ( );
FILL FILL_3_OAI21X1_43 ( );
FILL FILL_4_OAI21X1_43 ( );
FILL FILL_5_OAI21X1_43 ( );
FILL FILL_6_OAI21X1_43 ( );
FILL FILL_7_OAI21X1_43 ( );
FILL FILL_8_OAI21X1_43 ( );
FILL FILL_0_INVX1_49 ( );
FILL FILL_1_INVX1_49 ( );
FILL FILL_2_INVX1_49 ( );
FILL FILL_3_INVX1_49 ( );
FILL FILL_4_INVX1_49 ( );
FILL FILL_0_INVX1_292 ( );
FILL FILL_1_INVX1_292 ( );
FILL FILL_2_INVX1_292 ( );
FILL FILL_3_INVX1_292 ( );
FILL FILL_4_INVX1_292 ( );
FILL FILL_0_INVX1_29 ( );
FILL FILL_1_INVX1_29 ( );
FILL FILL_2_INVX1_29 ( );
FILL FILL_3_INVX1_29 ( );
FILL FILL_4_INVX1_29 ( );
FILL FILL_0_OAI21X1_25 ( );
FILL FILL_1_OAI21X1_25 ( );
FILL FILL_2_OAI21X1_25 ( );
FILL FILL_3_OAI21X1_25 ( );
FILL FILL_4_OAI21X1_25 ( );
FILL FILL_5_OAI21X1_25 ( );
FILL FILL_6_OAI21X1_25 ( );
FILL FILL_7_OAI21X1_25 ( );
FILL FILL_8_OAI21X1_25 ( );
FILL FILL_0_DFFSR_44 ( );
FILL FILL_1_DFFSR_44 ( );
FILL FILL_2_DFFSR_44 ( );
FILL FILL_3_DFFSR_44 ( );
FILL FILL_4_DFFSR_44 ( );
FILL FILL_5_DFFSR_44 ( );
FILL FILL_6_DFFSR_44 ( );
FILL FILL_7_DFFSR_44 ( );
FILL FILL_8_DFFSR_44 ( );
FILL FILL_9_DFFSR_44 ( );
FILL FILL_10_DFFSR_44 ( );
FILL FILL_11_DFFSR_44 ( );
FILL FILL_12_DFFSR_44 ( );
FILL FILL_13_DFFSR_44 ( );
FILL FILL_14_DFFSR_44 ( );
FILL FILL_15_DFFSR_44 ( );
FILL FILL_16_DFFSR_44 ( );
FILL FILL_17_DFFSR_44 ( );
FILL FILL_18_DFFSR_44 ( );
FILL FILL_19_DFFSR_44 ( );
FILL FILL_20_DFFSR_44 ( );
FILL FILL_21_DFFSR_44 ( );
FILL FILL_22_DFFSR_44 ( );
FILL FILL_23_DFFSR_44 ( );
FILL FILL_24_DFFSR_44 ( );
FILL FILL_25_DFFSR_44 ( );
FILL FILL_26_DFFSR_44 ( );
FILL FILL_27_DFFSR_44 ( );
FILL FILL_28_DFFSR_44 ( );
FILL FILL_29_DFFSR_44 ( );
FILL FILL_30_DFFSR_44 ( );
FILL FILL_31_DFFSR_44 ( );
FILL FILL_32_DFFSR_44 ( );
FILL FILL_33_DFFSR_44 ( );
FILL FILL_34_DFFSR_44 ( );
FILL FILL_35_DFFSR_44 ( );
FILL FILL_36_DFFSR_44 ( );
FILL FILL_37_DFFSR_44 ( );
FILL FILL_38_DFFSR_44 ( );
FILL FILL_39_DFFSR_44 ( );
FILL FILL_40_DFFSR_44 ( );
FILL FILL_41_DFFSR_44 ( );
FILL FILL_42_DFFSR_44 ( );
FILL FILL_43_DFFSR_44 ( );
FILL FILL_44_DFFSR_44 ( );
FILL FILL_45_DFFSR_44 ( );
FILL FILL_46_DFFSR_44 ( );
FILL FILL_47_DFFSR_44 ( );
FILL FILL_48_DFFSR_44 ( );
FILL FILL_49_DFFSR_44 ( );
FILL FILL_50_DFFSR_44 ( );
FILL FILL_0_NAND3X1_5 ( );
FILL FILL_1_NAND3X1_5 ( );
FILL FILL_2_NAND3X1_5 ( );
FILL FILL_3_NAND3X1_5 ( );
FILL FILL_4_NAND3X1_5 ( );
FILL FILL_5_NAND3X1_5 ( );
FILL FILL_6_NAND3X1_5 ( );
FILL FILL_7_NAND3X1_5 ( );
FILL FILL_8_NAND3X1_5 ( );
FILL FILL_9_NAND3X1_5 ( );
FILL FILL_0_NOR2X1_4 ( );
FILL FILL_1_NOR2X1_4 ( );
FILL FILL_2_NOR2X1_4 ( );
FILL FILL_3_NOR2X1_4 ( );
FILL FILL_4_NOR2X1_4 ( );
FILL FILL_5_NOR2X1_4 ( );
FILL FILL_6_NOR2X1_4 ( );
FILL FILL_0_NAND3X1_2 ( );
FILL FILL_1_NAND3X1_2 ( );
FILL FILL_2_NAND3X1_2 ( );
FILL FILL_3_NAND3X1_2 ( );
FILL FILL_4_NAND3X1_2 ( );
FILL FILL_5_NAND3X1_2 ( );
FILL FILL_6_NAND3X1_2 ( );
FILL FILL_7_NAND3X1_2 ( );
FILL FILL_8_NAND3X1_2 ( );
FILL FILL_0_OR2X2_1 ( );
FILL FILL_1_OR2X2_1 ( );
FILL FILL_2_OR2X2_1 ( );
FILL FILL_3_OR2X2_1 ( );
FILL FILL_4_OR2X2_1 ( );
FILL FILL_5_OR2X2_1 ( );
FILL FILL_6_OR2X2_1 ( );
FILL FILL_7_OR2X2_1 ( );
FILL FILL_8_OR2X2_1 ( );
FILL FILL_0_XOR2X1_2 ( );
FILL FILL_1_XOR2X1_2 ( );
FILL FILL_2_XOR2X1_2 ( );
FILL FILL_3_XOR2X1_2 ( );
FILL FILL_4_XOR2X1_2 ( );
FILL FILL_5_XOR2X1_2 ( );
FILL FILL_6_XOR2X1_2 ( );
FILL FILL_7_XOR2X1_2 ( );
FILL FILL_8_XOR2X1_2 ( );
FILL FILL_9_XOR2X1_2 ( );
FILL FILL_10_XOR2X1_2 ( );
FILL FILL_11_XOR2X1_2 ( );
FILL FILL_12_XOR2X1_2 ( );
FILL FILL_13_XOR2X1_2 ( );
FILL FILL_14_XOR2X1_2 ( );
FILL FILL_15_XOR2X1_2 ( );
FILL FILL_16_XOR2X1_2 ( );
FILL FILL_0_NAND2X1_208 ( );
FILL FILL_1_NAND2X1_208 ( );
FILL FILL_2_NAND2X1_208 ( );
FILL FILL_3_NAND2X1_208 ( );
FILL FILL_4_NAND2X1_208 ( );
FILL FILL_5_NAND2X1_208 ( );
FILL FILL_6_NAND2X1_208 ( );
FILL FILL_0_AOI21X1_18 ( );
FILL FILL_1_AOI21X1_18 ( );
FILL FILL_2_AOI21X1_18 ( );
FILL FILL_3_AOI21X1_18 ( );
FILL FILL_4_AOI21X1_18 ( );
FILL FILL_5_AOI21X1_18 ( );
FILL FILL_6_AOI21X1_18 ( );
FILL FILL_7_AOI21X1_18 ( );
FILL FILL_8_AOI21X1_18 ( );
FILL FILL_0_NAND3X1_85 ( );
FILL FILL_1_NAND3X1_85 ( );
FILL FILL_2_NAND3X1_85 ( );
FILL FILL_3_NAND3X1_85 ( );
FILL FILL_4_NAND3X1_85 ( );
FILL FILL_5_NAND3X1_85 ( );
FILL FILL_6_NAND3X1_85 ( );
FILL FILL_7_NAND3X1_85 ( );
FILL FILL_8_NAND3X1_85 ( );
FILL FILL_0_NAND2X1_217 ( );
FILL FILL_1_NAND2X1_217 ( );
FILL FILL_2_NAND2X1_217 ( );
FILL FILL_3_NAND2X1_217 ( );
FILL FILL_4_NAND2X1_217 ( );
FILL FILL_5_NAND2X1_217 ( );
FILL FILL_6_NAND2X1_217 ( );
FILL FILL_0_OAI21X1_237 ( );
FILL FILL_1_OAI21X1_237 ( );
FILL FILL_2_OAI21X1_237 ( );
FILL FILL_3_OAI21X1_237 ( );
FILL FILL_4_OAI21X1_237 ( );
FILL FILL_5_OAI21X1_237 ( );
FILL FILL_6_OAI21X1_237 ( );
FILL FILL_7_OAI21X1_237 ( );
FILL FILL_8_OAI21X1_237 ( );
FILL FILL_0_NAND2X1_261 ( );
FILL FILL_1_NAND2X1_261 ( );
FILL FILL_2_NAND2X1_261 ( );
FILL FILL_3_NAND2X1_261 ( );
FILL FILL_4_NAND2X1_261 ( );
FILL FILL_5_NAND2X1_261 ( );
FILL FILL_6_NAND2X1_261 ( );
FILL FILL_0_DFFSR_71 ( );
FILL FILL_1_DFFSR_71 ( );
FILL FILL_2_DFFSR_71 ( );
FILL FILL_3_DFFSR_71 ( );
FILL FILL_4_DFFSR_71 ( );
FILL FILL_5_DFFSR_71 ( );
FILL FILL_6_DFFSR_71 ( );
FILL FILL_7_DFFSR_71 ( );
FILL FILL_8_DFFSR_71 ( );
FILL FILL_9_DFFSR_71 ( );
FILL FILL_10_DFFSR_71 ( );
FILL FILL_11_DFFSR_71 ( );
FILL FILL_12_DFFSR_71 ( );
FILL FILL_13_DFFSR_71 ( );
FILL FILL_14_DFFSR_71 ( );
FILL FILL_15_DFFSR_71 ( );
FILL FILL_16_DFFSR_71 ( );
FILL FILL_17_DFFSR_71 ( );
FILL FILL_18_DFFSR_71 ( );
FILL FILL_19_DFFSR_71 ( );
FILL FILL_20_DFFSR_71 ( );
FILL FILL_21_DFFSR_71 ( );
FILL FILL_22_DFFSR_71 ( );
FILL FILL_23_DFFSR_71 ( );
FILL FILL_24_DFFSR_71 ( );
FILL FILL_25_DFFSR_71 ( );
FILL FILL_26_DFFSR_71 ( );
FILL FILL_27_DFFSR_71 ( );
FILL FILL_28_DFFSR_71 ( );
FILL FILL_29_DFFSR_71 ( );
FILL FILL_30_DFFSR_71 ( );
FILL FILL_31_DFFSR_71 ( );
FILL FILL_32_DFFSR_71 ( );
FILL FILL_33_DFFSR_71 ( );
FILL FILL_34_DFFSR_71 ( );
FILL FILL_35_DFFSR_71 ( );
FILL FILL_36_DFFSR_71 ( );
FILL FILL_37_DFFSR_71 ( );
FILL FILL_38_DFFSR_71 ( );
FILL FILL_39_DFFSR_71 ( );
FILL FILL_40_DFFSR_71 ( );
FILL FILL_41_DFFSR_71 ( );
FILL FILL_42_DFFSR_71 ( );
FILL FILL_43_DFFSR_71 ( );
FILL FILL_44_DFFSR_71 ( );
FILL FILL_45_DFFSR_71 ( );
FILL FILL_46_DFFSR_71 ( );
FILL FILL_47_DFFSR_71 ( );
FILL FILL_48_DFFSR_71 ( );
FILL FILL_49_DFFSR_71 ( );
FILL FILL_50_DFFSR_71 ( );
FILL FILL_0_NOR2X1_34 ( );
FILL FILL_1_NOR2X1_34 ( );
FILL FILL_2_NOR2X1_34 ( );
FILL FILL_3_NOR2X1_34 ( );
FILL FILL_4_NOR2X1_34 ( );
FILL FILL_5_NOR2X1_34 ( );
FILL FILL_6_NOR2X1_34 ( );
FILL FILL_0_NAND2X1_245 ( );
FILL FILL_1_NAND2X1_245 ( );
FILL FILL_2_NAND2X1_245 ( );
FILL FILL_3_NAND2X1_245 ( );
FILL FILL_4_NAND2X1_245 ( );
FILL FILL_5_NAND2X1_245 ( );
FILL FILL_6_NAND2X1_245 ( );
FILL FILL_0_INVX1_122 ( );
FILL FILL_1_INVX1_122 ( );
FILL FILL_2_INVX1_122 ( );
FILL FILL_3_INVX1_122 ( );
FILL FILL_4_INVX1_122 ( );
FILL FILL_0_NAND2X1_140 ( );
FILL FILL_1_NAND2X1_140 ( );
FILL FILL_2_NAND2X1_140 ( );
FILL FILL_3_NAND2X1_140 ( );
FILL FILL_4_NAND2X1_140 ( );
FILL FILL_5_NAND2X1_140 ( );
FILL FILL_6_NAND2X1_140 ( );
FILL FILL_0_INVX1_367 ( );
FILL FILL_1_INVX1_367 ( );
FILL FILL_2_INVX1_367 ( );
FILL FILL_3_INVX1_367 ( );
FILL FILL_0_INVX1_362 ( );
FILL FILL_1_INVX1_362 ( );
FILL FILL_2_INVX1_362 ( );
FILL FILL_3_INVX1_362 ( );
FILL FILL_4_INVX1_362 ( );
FILL FILL_0_INVX1_364 ( );
FILL FILL_1_INVX1_364 ( );
FILL FILL_2_INVX1_364 ( );
FILL FILL_3_INVX1_364 ( );
FILL FILL_4_INVX1_364 ( );
FILL FILL_0_OAI22X1_53 ( );
FILL FILL_1_OAI22X1_53 ( );
FILL FILL_2_OAI22X1_53 ( );
FILL FILL_3_OAI22X1_53 ( );
FILL FILL_4_OAI22X1_53 ( );
FILL FILL_5_OAI22X1_53 ( );
FILL FILL_6_OAI22X1_53 ( );
FILL FILL_7_OAI22X1_53 ( );
FILL FILL_8_OAI22X1_53 ( );
FILL FILL_9_OAI22X1_53 ( );
FILL FILL_10_OAI22X1_53 ( );
FILL FILL_11_OAI22X1_53 ( );
FILL FILL_0_DFFSR_140 ( );
FILL FILL_1_DFFSR_140 ( );
FILL FILL_2_DFFSR_140 ( );
FILL FILL_3_DFFSR_140 ( );
FILL FILL_4_DFFSR_140 ( );
FILL FILL_5_DFFSR_140 ( );
FILL FILL_6_DFFSR_140 ( );
FILL FILL_7_DFFSR_140 ( );
FILL FILL_8_DFFSR_140 ( );
FILL FILL_9_DFFSR_140 ( );
FILL FILL_10_DFFSR_140 ( );
FILL FILL_11_DFFSR_140 ( );
FILL FILL_12_DFFSR_140 ( );
FILL FILL_13_DFFSR_140 ( );
FILL FILL_14_DFFSR_140 ( );
FILL FILL_15_DFFSR_140 ( );
FILL FILL_16_DFFSR_140 ( );
FILL FILL_17_DFFSR_140 ( );
FILL FILL_18_DFFSR_140 ( );
FILL FILL_19_DFFSR_140 ( );
FILL FILL_20_DFFSR_140 ( );
FILL FILL_21_DFFSR_140 ( );
FILL FILL_22_DFFSR_140 ( );
FILL FILL_23_DFFSR_140 ( );
FILL FILL_24_DFFSR_140 ( );
FILL FILL_25_DFFSR_140 ( );
FILL FILL_26_DFFSR_140 ( );
FILL FILL_27_DFFSR_140 ( );
FILL FILL_28_DFFSR_140 ( );
FILL FILL_29_DFFSR_140 ( );
FILL FILL_30_DFFSR_140 ( );
FILL FILL_31_DFFSR_140 ( );
FILL FILL_32_DFFSR_140 ( );
FILL FILL_33_DFFSR_140 ( );
FILL FILL_34_DFFSR_140 ( );
FILL FILL_35_DFFSR_140 ( );
FILL FILL_36_DFFSR_140 ( );
FILL FILL_37_DFFSR_140 ( );
FILL FILL_38_DFFSR_140 ( );
FILL FILL_39_DFFSR_140 ( );
FILL FILL_40_DFFSR_140 ( );
FILL FILL_41_DFFSR_140 ( );
FILL FILL_42_DFFSR_140 ( );
FILL FILL_43_DFFSR_140 ( );
FILL FILL_44_DFFSR_140 ( );
FILL FILL_45_DFFSR_140 ( );
FILL FILL_46_DFFSR_140 ( );
FILL FILL_47_DFFSR_140 ( );
FILL FILL_48_DFFSR_140 ( );
FILL FILL_49_DFFSR_140 ( );
FILL FILL_50_DFFSR_140 ( );
FILL FILL_0_INVX1_428 ( );
FILL FILL_1_INVX1_428 ( );
FILL FILL_2_INVX1_428 ( );
FILL FILL_3_INVX1_428 ( );
FILL FILL_4_INVX1_428 ( );
FILL FILL_0_NAND2X1_277 ( );
FILL FILL_1_NAND2X1_277 ( );
FILL FILL_2_NAND2X1_277 ( );
FILL FILL_3_NAND2X1_277 ( );
FILL FILL_4_NAND2X1_277 ( );
FILL FILL_5_NAND2X1_277 ( );
FILL FILL_6_NAND2X1_277 ( );
FILL FILL_0_INVX1_427 ( );
FILL FILL_1_INVX1_427 ( );
FILL FILL_2_INVX1_427 ( );
FILL FILL_3_INVX1_427 ( );
FILL FILL_0_NAND2X1_276 ( );
FILL FILL_1_NAND2X1_276 ( );
FILL FILL_2_NAND2X1_276 ( );
FILL FILL_3_NAND2X1_276 ( );
FILL FILL_4_NAND2X1_276 ( );
FILL FILL_5_NAND2X1_276 ( );
FILL FILL_6_NAND2X1_276 ( );
FILL FILL_0_NAND3X1_134 ( );
FILL FILL_1_NAND3X1_134 ( );
FILL FILL_2_NAND3X1_134 ( );
FILL FILL_3_NAND3X1_134 ( );
FILL FILL_4_NAND3X1_134 ( );
FILL FILL_5_NAND3X1_134 ( );
FILL FILL_6_NAND3X1_134 ( );
FILL FILL_7_NAND3X1_134 ( );
FILL FILL_8_NAND3X1_134 ( );
FILL FILL_0_INVX1_438 ( );
FILL FILL_1_INVX1_438 ( );
FILL FILL_2_INVX1_438 ( );
FILL FILL_3_INVX1_438 ( );
FILL FILL_4_INVX1_438 ( );
FILL FILL_0_NAND2X1_285 ( );
FILL FILL_1_NAND2X1_285 ( );
FILL FILL_2_NAND2X1_285 ( );
FILL FILL_3_NAND2X1_285 ( );
FILL FILL_4_NAND2X1_285 ( );
FILL FILL_5_NAND2X1_285 ( );
FILL FILL_6_NAND2X1_285 ( );
FILL FILL_0_INVX1_264 ( );
FILL FILL_1_INVX1_264 ( );
FILL FILL_2_INVX1_264 ( );
FILL FILL_3_INVX1_264 ( );
FILL FILL_4_INVX1_264 ( );
FILL FILL_0_NAND3X1_112 ( );
FILL FILL_1_NAND3X1_112 ( );
FILL FILL_2_NAND3X1_112 ( );
FILL FILL_3_NAND3X1_112 ( );
FILL FILL_4_NAND3X1_112 ( );
FILL FILL_5_NAND3X1_112 ( );
FILL FILL_6_NAND3X1_112 ( );
FILL FILL_7_NAND3X1_112 ( );
FILL FILL_8_NAND3X1_112 ( );
FILL FILL_0_INVX1_265 ( );
FILL FILL_1_INVX1_265 ( );
FILL FILL_2_INVX1_265 ( );
FILL FILL_3_INVX1_265 ( );
FILL FILL_4_INVX1_265 ( );
FILL FILL_0_NAND3X1_114 ( );
FILL FILL_1_NAND3X1_114 ( );
FILL FILL_2_NAND3X1_114 ( );
FILL FILL_3_NAND3X1_114 ( );
FILL FILL_4_NAND3X1_114 ( );
FILL FILL_5_NAND3X1_114 ( );
FILL FILL_6_NAND3X1_114 ( );
FILL FILL_7_NAND3X1_114 ( );
FILL FILL_8_NAND3X1_114 ( );
FILL FILL_9_NAND3X1_114 ( );
FILL FILL_0_OAI22X1_32 ( );
FILL FILL_1_OAI22X1_32 ( );
FILL FILL_2_OAI22X1_32 ( );
FILL FILL_3_OAI22X1_32 ( );
FILL FILL_4_OAI22X1_32 ( );
FILL FILL_5_OAI22X1_32 ( );
FILL FILL_6_OAI22X1_32 ( );
FILL FILL_7_OAI22X1_32 ( );
FILL FILL_8_OAI22X1_32 ( );
FILL FILL_9_OAI22X1_32 ( );
FILL FILL_10_OAI22X1_32 ( );
FILL FILL_0_NAND2X1_39 ( );
FILL FILL_1_NAND2X1_39 ( );
FILL FILL_2_NAND2X1_39 ( );
FILL FILL_3_NAND2X1_39 ( );
FILL FILL_4_NAND2X1_39 ( );
FILL FILL_5_NAND2X1_39 ( );
FILL FILL_6_NAND2X1_39 ( );
FILL FILL_0_INVX1_294 ( );
FILL FILL_1_INVX1_294 ( );
FILL FILL_2_INVX1_294 ( );
FILL FILL_3_INVX1_294 ( );
FILL FILL_4_INVX1_294 ( );
FILL FILL_0_DFFSR_53 ( );
FILL FILL_1_DFFSR_53 ( );
FILL FILL_2_DFFSR_53 ( );
FILL FILL_3_DFFSR_53 ( );
FILL FILL_4_DFFSR_53 ( );
FILL FILL_5_DFFSR_53 ( );
FILL FILL_6_DFFSR_53 ( );
FILL FILL_7_DFFSR_53 ( );
FILL FILL_8_DFFSR_53 ( );
FILL FILL_9_DFFSR_53 ( );
FILL FILL_10_DFFSR_53 ( );
FILL FILL_11_DFFSR_53 ( );
FILL FILL_12_DFFSR_53 ( );
FILL FILL_13_DFFSR_53 ( );
FILL FILL_14_DFFSR_53 ( );
FILL FILL_15_DFFSR_53 ( );
FILL FILL_16_DFFSR_53 ( );
FILL FILL_17_DFFSR_53 ( );
FILL FILL_18_DFFSR_53 ( );
FILL FILL_19_DFFSR_53 ( );
FILL FILL_20_DFFSR_53 ( );
FILL FILL_21_DFFSR_53 ( );
FILL FILL_22_DFFSR_53 ( );
FILL FILL_23_DFFSR_53 ( );
FILL FILL_24_DFFSR_53 ( );
FILL FILL_25_DFFSR_53 ( );
FILL FILL_26_DFFSR_53 ( );
FILL FILL_27_DFFSR_53 ( );
FILL FILL_28_DFFSR_53 ( );
FILL FILL_29_DFFSR_53 ( );
FILL FILL_30_DFFSR_53 ( );
FILL FILL_31_DFFSR_53 ( );
FILL FILL_32_DFFSR_53 ( );
FILL FILL_33_DFFSR_53 ( );
FILL FILL_34_DFFSR_53 ( );
FILL FILL_35_DFFSR_53 ( );
FILL FILL_36_DFFSR_53 ( );
FILL FILL_37_DFFSR_53 ( );
FILL FILL_38_DFFSR_53 ( );
FILL FILL_39_DFFSR_53 ( );
FILL FILL_40_DFFSR_53 ( );
FILL FILL_41_DFFSR_53 ( );
FILL FILL_42_DFFSR_53 ( );
FILL FILL_43_DFFSR_53 ( );
FILL FILL_44_DFFSR_53 ( );
FILL FILL_45_DFFSR_53 ( );
FILL FILL_46_DFFSR_53 ( );
FILL FILL_47_DFFSR_53 ( );
FILL FILL_48_DFFSR_53 ( );
FILL FILL_49_DFFSR_53 ( );
FILL FILL_50_DFFSR_53 ( );
FILL FILL_51_DFFSR_53 ( );
FILL FILL_0_NAND2X1_52 ( );
FILL FILL_1_NAND2X1_52 ( );
FILL FILL_2_NAND2X1_52 ( );
FILL FILL_3_NAND2X1_52 ( );
FILL FILL_4_NAND2X1_52 ( );
FILL FILL_5_NAND2X1_52 ( );
FILL FILL_6_NAND2X1_52 ( );
FILL FILL_0_DFFSR_10 ( );
FILL FILL_1_DFFSR_10 ( );
FILL FILL_2_DFFSR_10 ( );
FILL FILL_3_DFFSR_10 ( );
FILL FILL_4_DFFSR_10 ( );
FILL FILL_5_DFFSR_10 ( );
FILL FILL_6_DFFSR_10 ( );
FILL FILL_7_DFFSR_10 ( );
FILL FILL_8_DFFSR_10 ( );
FILL FILL_9_DFFSR_10 ( );
FILL FILL_10_DFFSR_10 ( );
FILL FILL_11_DFFSR_10 ( );
FILL FILL_12_DFFSR_10 ( );
FILL FILL_13_DFFSR_10 ( );
FILL FILL_14_DFFSR_10 ( );
FILL FILL_15_DFFSR_10 ( );
FILL FILL_16_DFFSR_10 ( );
FILL FILL_17_DFFSR_10 ( );
FILL FILL_18_DFFSR_10 ( );
FILL FILL_19_DFFSR_10 ( );
FILL FILL_20_DFFSR_10 ( );
FILL FILL_21_DFFSR_10 ( );
FILL FILL_22_DFFSR_10 ( );
FILL FILL_23_DFFSR_10 ( );
FILL FILL_24_DFFSR_10 ( );
FILL FILL_25_DFFSR_10 ( );
FILL FILL_26_DFFSR_10 ( );
FILL FILL_27_DFFSR_10 ( );
FILL FILL_28_DFFSR_10 ( );
FILL FILL_29_DFFSR_10 ( );
FILL FILL_30_DFFSR_10 ( );
FILL FILL_31_DFFSR_10 ( );
FILL FILL_32_DFFSR_10 ( );
FILL FILL_33_DFFSR_10 ( );
FILL FILL_34_DFFSR_10 ( );
FILL FILL_35_DFFSR_10 ( );
FILL FILL_36_DFFSR_10 ( );
FILL FILL_37_DFFSR_10 ( );
FILL FILL_38_DFFSR_10 ( );
FILL FILL_39_DFFSR_10 ( );
FILL FILL_40_DFFSR_10 ( );
FILL FILL_41_DFFSR_10 ( );
FILL FILL_42_DFFSR_10 ( );
FILL FILL_43_DFFSR_10 ( );
FILL FILL_44_DFFSR_10 ( );
FILL FILL_45_DFFSR_10 ( );
FILL FILL_46_DFFSR_10 ( );
FILL FILL_47_DFFSR_10 ( );
FILL FILL_48_DFFSR_10 ( );
FILL FILL_49_DFFSR_10 ( );
FILL FILL_50_DFFSR_10 ( );
FILL FILL_0_OAI21X1_179 ( );
FILL FILL_1_OAI21X1_179 ( );
FILL FILL_2_OAI21X1_179 ( );
FILL FILL_3_OAI21X1_179 ( );
FILL FILL_4_OAI21X1_179 ( );
FILL FILL_5_OAI21X1_179 ( );
FILL FILL_6_OAI21X1_179 ( );
FILL FILL_7_OAI21X1_179 ( );
FILL FILL_8_OAI21X1_179 ( );
FILL FILL_0_OAI21X1_177 ( );
FILL FILL_1_OAI21X1_177 ( );
FILL FILL_2_OAI21X1_177 ( );
FILL FILL_3_OAI21X1_177 ( );
FILL FILL_4_OAI21X1_177 ( );
FILL FILL_5_OAI21X1_177 ( );
FILL FILL_6_OAI21X1_177 ( );
FILL FILL_7_OAI21X1_177 ( );
FILL FILL_8_OAI21X1_177 ( );
FILL FILL_9_OAI21X1_177 ( );
FILL FILL_0_OAI21X1_180 ( );
FILL FILL_1_OAI21X1_180 ( );
FILL FILL_2_OAI21X1_180 ( );
FILL FILL_3_OAI21X1_180 ( );
FILL FILL_4_OAI21X1_180 ( );
FILL FILL_5_OAI21X1_180 ( );
FILL FILL_6_OAI21X1_180 ( );
FILL FILL_7_OAI21X1_180 ( );
FILL FILL_8_OAI21X1_180 ( );
FILL FILL_0_INVX1_218 ( );
FILL FILL_1_INVX1_218 ( );
FILL FILL_2_INVX1_218 ( );
FILL FILL_3_INVX1_218 ( );
FILL FILL_0_OAI21X1_211 ( );
FILL FILL_1_OAI21X1_211 ( );
FILL FILL_2_OAI21X1_211 ( );
FILL FILL_3_OAI21X1_211 ( );
FILL FILL_4_OAI21X1_211 ( );
FILL FILL_5_OAI21X1_211 ( );
FILL FILL_6_OAI21X1_211 ( );
FILL FILL_7_OAI21X1_211 ( );
FILL FILL_8_OAI21X1_211 ( );
FILL FILL_0_INVX1_243 ( );
FILL FILL_1_INVX1_243 ( );
FILL FILL_2_INVX1_243 ( );
FILL FILL_3_INVX1_243 ( );
FILL FILL_4_INVX1_243 ( );
FILL FILL_0_NAND2X1_209 ( );
FILL FILL_1_NAND2X1_209 ( );
FILL FILL_2_NAND2X1_209 ( );
FILL FILL_3_NAND2X1_209 ( );
FILL FILL_4_NAND2X1_209 ( );
FILL FILL_5_NAND2X1_209 ( );
FILL FILL_6_NAND2X1_209 ( );
FILL FILL_0_OAI21X1_228 ( );
FILL FILL_1_OAI21X1_228 ( );
FILL FILL_2_OAI21X1_228 ( );
FILL FILL_3_OAI21X1_228 ( );
FILL FILL_4_OAI21X1_228 ( );
FILL FILL_5_OAI21X1_228 ( );
FILL FILL_6_OAI21X1_228 ( );
FILL FILL_7_OAI21X1_228 ( );
FILL FILL_8_OAI21X1_228 ( );
FILL FILL_9_OAI21X1_228 ( );
FILL FILL_0_AOI21X1_28 ( );
FILL FILL_1_AOI21X1_28 ( );
FILL FILL_2_AOI21X1_28 ( );
FILL FILL_3_AOI21X1_28 ( );
FILL FILL_4_AOI21X1_28 ( );
FILL FILL_5_AOI21X1_28 ( );
FILL FILL_6_AOI21X1_28 ( );
FILL FILL_7_AOI21X1_28 ( );
FILL FILL_8_AOI21X1_28 ( );
FILL FILL_0_NAND3X1_60 ( );
FILL FILL_1_NAND3X1_60 ( );
FILL FILL_2_NAND3X1_60 ( );
FILL FILL_3_NAND3X1_60 ( );
FILL FILL_4_NAND3X1_60 ( );
FILL FILL_5_NAND3X1_60 ( );
FILL FILL_6_NAND3X1_60 ( );
FILL FILL_7_NAND3X1_60 ( );
FILL FILL_8_NAND3X1_60 ( );
FILL FILL_0_DFFSR_114 ( );
FILL FILL_1_DFFSR_114 ( );
FILL FILL_2_DFFSR_114 ( );
FILL FILL_3_DFFSR_114 ( );
FILL FILL_4_DFFSR_114 ( );
FILL FILL_5_DFFSR_114 ( );
FILL FILL_6_DFFSR_114 ( );
FILL FILL_7_DFFSR_114 ( );
FILL FILL_8_DFFSR_114 ( );
FILL FILL_9_DFFSR_114 ( );
FILL FILL_10_DFFSR_114 ( );
FILL FILL_11_DFFSR_114 ( );
FILL FILL_12_DFFSR_114 ( );
FILL FILL_13_DFFSR_114 ( );
FILL FILL_14_DFFSR_114 ( );
FILL FILL_15_DFFSR_114 ( );
FILL FILL_16_DFFSR_114 ( );
FILL FILL_17_DFFSR_114 ( );
FILL FILL_18_DFFSR_114 ( );
FILL FILL_19_DFFSR_114 ( );
FILL FILL_20_DFFSR_114 ( );
FILL FILL_21_DFFSR_114 ( );
FILL FILL_22_DFFSR_114 ( );
FILL FILL_23_DFFSR_114 ( );
FILL FILL_24_DFFSR_114 ( );
FILL FILL_25_DFFSR_114 ( );
FILL FILL_26_DFFSR_114 ( );
FILL FILL_27_DFFSR_114 ( );
FILL FILL_28_DFFSR_114 ( );
FILL FILL_29_DFFSR_114 ( );
FILL FILL_30_DFFSR_114 ( );
FILL FILL_31_DFFSR_114 ( );
FILL FILL_32_DFFSR_114 ( );
FILL FILL_33_DFFSR_114 ( );
FILL FILL_34_DFFSR_114 ( );
FILL FILL_35_DFFSR_114 ( );
FILL FILL_36_DFFSR_114 ( );
FILL FILL_37_DFFSR_114 ( );
FILL FILL_38_DFFSR_114 ( );
FILL FILL_39_DFFSR_114 ( );
FILL FILL_40_DFFSR_114 ( );
FILL FILL_41_DFFSR_114 ( );
FILL FILL_42_DFFSR_114 ( );
FILL FILL_43_DFFSR_114 ( );
FILL FILL_44_DFFSR_114 ( );
FILL FILL_45_DFFSR_114 ( );
FILL FILL_46_DFFSR_114 ( );
FILL FILL_47_DFFSR_114 ( );
FILL FILL_48_DFFSR_114 ( );
FILL FILL_49_DFFSR_114 ( );
FILL FILL_50_DFFSR_114 ( );
FILL FILL_0_INVX1_330 ( );
FILL FILL_1_INVX1_330 ( );
FILL FILL_2_INVX1_330 ( );
FILL FILL_3_INVX1_330 ( );
FILL FILL_4_INVX1_330 ( );
FILL FILL_0_OAI22X1_37 ( );
FILL FILL_1_OAI22X1_37 ( );
FILL FILL_2_OAI22X1_37 ( );
FILL FILL_3_OAI22X1_37 ( );
FILL FILL_4_OAI22X1_37 ( );
FILL FILL_5_OAI22X1_37 ( );
FILL FILL_6_OAI22X1_37 ( );
FILL FILL_7_OAI22X1_37 ( );
FILL FILL_8_OAI22X1_37 ( );
FILL FILL_9_OAI22X1_37 ( );
FILL FILL_10_OAI22X1_37 ( );
FILL FILL_11_OAI22X1_37 ( );
FILL FILL_0_DFFSR_85 ( );
FILL FILL_1_DFFSR_85 ( );
FILL FILL_2_DFFSR_85 ( );
FILL FILL_3_DFFSR_85 ( );
FILL FILL_4_DFFSR_85 ( );
FILL FILL_5_DFFSR_85 ( );
FILL FILL_6_DFFSR_85 ( );
FILL FILL_7_DFFSR_85 ( );
FILL FILL_8_DFFSR_85 ( );
FILL FILL_9_DFFSR_85 ( );
FILL FILL_10_DFFSR_85 ( );
FILL FILL_11_DFFSR_85 ( );
FILL FILL_12_DFFSR_85 ( );
FILL FILL_13_DFFSR_85 ( );
FILL FILL_14_DFFSR_85 ( );
FILL FILL_15_DFFSR_85 ( );
FILL FILL_16_DFFSR_85 ( );
FILL FILL_17_DFFSR_85 ( );
FILL FILL_18_DFFSR_85 ( );
FILL FILL_19_DFFSR_85 ( );
FILL FILL_20_DFFSR_85 ( );
FILL FILL_21_DFFSR_85 ( );
FILL FILL_22_DFFSR_85 ( );
FILL FILL_23_DFFSR_85 ( );
FILL FILL_24_DFFSR_85 ( );
FILL FILL_25_DFFSR_85 ( );
FILL FILL_26_DFFSR_85 ( );
FILL FILL_27_DFFSR_85 ( );
FILL FILL_28_DFFSR_85 ( );
FILL FILL_29_DFFSR_85 ( );
FILL FILL_30_DFFSR_85 ( );
FILL FILL_31_DFFSR_85 ( );
FILL FILL_32_DFFSR_85 ( );
FILL FILL_33_DFFSR_85 ( );
FILL FILL_34_DFFSR_85 ( );
FILL FILL_35_DFFSR_85 ( );
FILL FILL_36_DFFSR_85 ( );
FILL FILL_37_DFFSR_85 ( );
FILL FILL_38_DFFSR_85 ( );
FILL FILL_39_DFFSR_85 ( );
FILL FILL_40_DFFSR_85 ( );
FILL FILL_41_DFFSR_85 ( );
FILL FILL_42_DFFSR_85 ( );
FILL FILL_43_DFFSR_85 ( );
FILL FILL_44_DFFSR_85 ( );
FILL FILL_45_DFFSR_85 ( );
FILL FILL_46_DFFSR_85 ( );
FILL FILL_47_DFFSR_85 ( );
FILL FILL_48_DFFSR_85 ( );
FILL FILL_49_DFFSR_85 ( );
FILL FILL_50_DFFSR_85 ( );
FILL FILL_0_OAI21X1_140 ( );
FILL FILL_1_OAI21X1_140 ( );
FILL FILL_2_OAI21X1_140 ( );
FILL FILL_3_OAI21X1_140 ( );
FILL FILL_4_OAI21X1_140 ( );
FILL FILL_5_OAI21X1_140 ( );
FILL FILL_6_OAI21X1_140 ( );
FILL FILL_7_OAI21X1_140 ( );
FILL FILL_8_OAI21X1_140 ( );
FILL FILL_0_DFFSR_16 ( );
FILL FILL_1_DFFSR_16 ( );
FILL FILL_2_DFFSR_16 ( );
FILL FILL_3_DFFSR_16 ( );
FILL FILL_4_DFFSR_16 ( );
FILL FILL_5_DFFSR_16 ( );
FILL FILL_6_DFFSR_16 ( );
FILL FILL_7_DFFSR_16 ( );
FILL FILL_8_DFFSR_16 ( );
FILL FILL_9_DFFSR_16 ( );
FILL FILL_10_DFFSR_16 ( );
FILL FILL_11_DFFSR_16 ( );
FILL FILL_12_DFFSR_16 ( );
FILL FILL_13_DFFSR_16 ( );
FILL FILL_14_DFFSR_16 ( );
FILL FILL_15_DFFSR_16 ( );
FILL FILL_16_DFFSR_16 ( );
FILL FILL_17_DFFSR_16 ( );
FILL FILL_18_DFFSR_16 ( );
FILL FILL_19_DFFSR_16 ( );
FILL FILL_20_DFFSR_16 ( );
FILL FILL_21_DFFSR_16 ( );
FILL FILL_22_DFFSR_16 ( );
FILL FILL_23_DFFSR_16 ( );
FILL FILL_24_DFFSR_16 ( );
FILL FILL_25_DFFSR_16 ( );
FILL FILL_26_DFFSR_16 ( );
FILL FILL_27_DFFSR_16 ( );
FILL FILL_28_DFFSR_16 ( );
FILL FILL_29_DFFSR_16 ( );
FILL FILL_30_DFFSR_16 ( );
FILL FILL_31_DFFSR_16 ( );
FILL FILL_32_DFFSR_16 ( );
FILL FILL_33_DFFSR_16 ( );
FILL FILL_34_DFFSR_16 ( );
FILL FILL_35_DFFSR_16 ( );
FILL FILL_36_DFFSR_16 ( );
FILL FILL_37_DFFSR_16 ( );
FILL FILL_38_DFFSR_16 ( );
FILL FILL_39_DFFSR_16 ( );
FILL FILL_40_DFFSR_16 ( );
FILL FILL_41_DFFSR_16 ( );
FILL FILL_42_DFFSR_16 ( );
FILL FILL_43_DFFSR_16 ( );
FILL FILL_44_DFFSR_16 ( );
FILL FILL_45_DFFSR_16 ( );
FILL FILL_46_DFFSR_16 ( );
FILL FILL_47_DFFSR_16 ( );
FILL FILL_48_DFFSR_16 ( );
FILL FILL_49_DFFSR_16 ( );
FILL FILL_50_DFFSR_16 ( );
FILL FILL_0_AOI21X1_48 ( );
FILL FILL_1_AOI21X1_48 ( );
FILL FILL_2_AOI21X1_48 ( );
FILL FILL_3_AOI21X1_48 ( );
FILL FILL_4_AOI21X1_48 ( );
FILL FILL_5_AOI21X1_48 ( );
FILL FILL_6_AOI21X1_48 ( );
FILL FILL_7_AOI21X1_48 ( );
FILL FILL_8_AOI21X1_48 ( );
FILL FILL_9_AOI21X1_48 ( );
FILL FILL_0_NAND2X1_286 ( );
FILL FILL_1_NAND2X1_286 ( );
FILL FILL_2_NAND2X1_286 ( );
FILL FILL_3_NAND2X1_286 ( );
FILL FILL_4_NAND2X1_286 ( );
FILL FILL_5_NAND2X1_286 ( );
FILL FILL_6_NAND2X1_286 ( );
FILL FILL_0_INVX1_46 ( );
FILL FILL_1_INVX1_46 ( );
FILL FILL_2_INVX1_46 ( );
FILL FILL_3_INVX1_46 ( );
FILL FILL_0_INVX1_432 ( );
FILL FILL_1_INVX1_432 ( );
FILL FILL_2_INVX1_432 ( );
FILL FILL_3_INVX1_432 ( );
FILL FILL_0_NAND3X1_111 ( );
FILL FILL_1_NAND3X1_111 ( );
FILL FILL_2_NAND3X1_111 ( );
FILL FILL_3_NAND3X1_111 ( );
FILL FILL_4_NAND3X1_111 ( );
FILL FILL_5_NAND3X1_111 ( );
FILL FILL_6_NAND3X1_111 ( );
FILL FILL_7_NAND3X1_111 ( );
FILL FILL_8_NAND3X1_111 ( );
FILL FILL_0_NAND3X1_116 ( );
FILL FILL_1_NAND3X1_116 ( );
FILL FILL_2_NAND3X1_116 ( );
FILL FILL_3_NAND3X1_116 ( );
FILL FILL_4_NAND3X1_116 ( );
FILL FILL_5_NAND3X1_116 ( );
FILL FILL_6_NAND3X1_116 ( );
FILL FILL_7_NAND3X1_116 ( );
FILL FILL_8_NAND3X1_116 ( );
FILL FILL_0_NOR2X1_25 ( );
FILL FILL_1_NOR2X1_25 ( );
FILL FILL_2_NOR2X1_25 ( );
FILL FILL_3_NOR2X1_25 ( );
FILL FILL_4_NOR2X1_25 ( );
FILL FILL_5_NOR2X1_25 ( );
FILL FILL_6_NOR2X1_25 ( );
FILL FILL_0_INVX1_318 ( );
FILL FILL_1_INVX1_318 ( );
FILL FILL_2_INVX1_318 ( );
FILL FILL_3_INVX1_318 ( );
FILL FILL_4_INVX1_318 ( );
FILL FILL_0_OAI22X1_31 ( );
FILL FILL_1_OAI22X1_31 ( );
FILL FILL_2_OAI22X1_31 ( );
FILL FILL_3_OAI22X1_31 ( );
FILL FILL_4_OAI22X1_31 ( );
FILL FILL_5_OAI22X1_31 ( );
FILL FILL_6_OAI22X1_31 ( );
FILL FILL_7_OAI22X1_31 ( );
FILL FILL_8_OAI22X1_31 ( );
FILL FILL_9_OAI22X1_31 ( );
FILL FILL_10_OAI22X1_31 ( );
FILL FILL_0_OAI22X1_19 ( );
FILL FILL_1_OAI22X1_19 ( );
FILL FILL_2_OAI22X1_19 ( );
FILL FILL_3_OAI22X1_19 ( );
FILL FILL_4_OAI22X1_19 ( );
FILL FILL_5_OAI22X1_19 ( );
FILL FILL_6_OAI22X1_19 ( );
FILL FILL_7_OAI22X1_19 ( );
FILL FILL_8_OAI22X1_19 ( );
FILL FILL_9_OAI22X1_19 ( );
FILL FILL_10_OAI22X1_19 ( );
FILL FILL_0_OAI21X1_39 ( );
FILL FILL_1_OAI21X1_39 ( );
FILL FILL_2_OAI21X1_39 ( );
FILL FILL_3_OAI21X1_39 ( );
FILL FILL_4_OAI21X1_39 ( );
FILL FILL_5_OAI21X1_39 ( );
FILL FILL_6_OAI21X1_39 ( );
FILL FILL_7_OAI21X1_39 ( );
FILL FILL_8_OAI21X1_39 ( );
FILL FILL_9_OAI21X1_39 ( );
FILL FILL_0_INVX1_293 ( );
FILL FILL_1_INVX1_293 ( );
FILL FILL_2_INVX1_293 ( );
FILL FILL_3_INVX1_293 ( );
FILL FILL_4_INVX1_293 ( );
FILL FILL_0_INVX1_60 ( );
FILL FILL_1_INVX1_60 ( );
FILL FILL_2_INVX1_60 ( );
FILL FILL_3_INVX1_60 ( );
FILL FILL_4_INVX1_60 ( );
FILL FILL_0_OAI21X1_53 ( );
FILL FILL_1_OAI21X1_53 ( );
FILL FILL_2_OAI21X1_53 ( );
FILL FILL_3_OAI21X1_53 ( );
FILL FILL_4_OAI21X1_53 ( );
FILL FILL_5_OAI21X1_53 ( );
FILL FILL_6_OAI21X1_53 ( );
FILL FILL_7_OAI21X1_53 ( );
FILL FILL_8_OAI21X1_53 ( );
FILL FILL_0_DFFPOSX1_27 ( );
FILL FILL_1_DFFPOSX1_27 ( );
FILL FILL_2_DFFPOSX1_27 ( );
FILL FILL_3_DFFPOSX1_27 ( );
FILL FILL_4_DFFPOSX1_27 ( );
FILL FILL_5_DFFPOSX1_27 ( );
FILL FILL_6_DFFPOSX1_27 ( );
FILL FILL_7_DFFPOSX1_27 ( );
FILL FILL_8_DFFPOSX1_27 ( );
FILL FILL_9_DFFPOSX1_27 ( );
FILL FILL_10_DFFPOSX1_27 ( );
FILL FILL_11_DFFPOSX1_27 ( );
FILL FILL_12_DFFPOSX1_27 ( );
FILL FILL_13_DFFPOSX1_27 ( );
FILL FILL_14_DFFPOSX1_27 ( );
FILL FILL_15_DFFPOSX1_27 ( );
FILL FILL_16_DFFPOSX1_27 ( );
FILL FILL_17_DFFPOSX1_27 ( );
FILL FILL_18_DFFPOSX1_27 ( );
FILL FILL_19_DFFPOSX1_27 ( );
FILL FILL_20_DFFPOSX1_27 ( );
FILL FILL_21_DFFPOSX1_27 ( );
FILL FILL_22_DFFPOSX1_27 ( );
FILL FILL_23_DFFPOSX1_27 ( );
FILL FILL_24_DFFPOSX1_27 ( );
FILL FILL_25_DFFPOSX1_27 ( );
FILL FILL_26_DFFPOSX1_27 ( );
FILL FILL_27_DFFPOSX1_27 ( );
FILL FILL_0_NAND2X1_36 ( );
FILL FILL_1_NAND2X1_36 ( );
FILL FILL_2_NAND2X1_36 ( );
FILL FILL_3_NAND2X1_36 ( );
FILL FILL_4_NAND2X1_36 ( );
FILL FILL_5_NAND2X1_36 ( );
FILL FILL_6_NAND2X1_36 ( );
FILL FILL_0_OAI21X1_44 ( );
FILL FILL_1_OAI21X1_44 ( );
FILL FILL_2_OAI21X1_44 ( );
FILL FILL_3_OAI21X1_44 ( );
FILL FILL_4_OAI21X1_44 ( );
FILL FILL_5_OAI21X1_44 ( );
FILL FILL_6_OAI21X1_44 ( );
FILL FILL_7_OAI21X1_44 ( );
FILL FILL_8_OAI21X1_44 ( );
FILL FILL_0_NAND2X1_44 ( );
FILL FILL_1_NAND2X1_44 ( );
FILL FILL_2_NAND2X1_44 ( );
FILL FILL_3_NAND2X1_44 ( );
FILL FILL_4_NAND2X1_44 ( );
FILL FILL_5_NAND2X1_44 ( );
FILL FILL_6_NAND2X1_44 ( );
FILL FILL_0_INVX1_12 ( );
FILL FILL_1_INVX1_12 ( );
FILL FILL_2_INVX1_12 ( );
FILL FILL_3_INVX1_12 ( );
FILL FILL_0_OAI21X1_10 ( );
FILL FILL_1_OAI21X1_10 ( );
FILL FILL_2_OAI21X1_10 ( );
FILL FILL_3_OAI21X1_10 ( );
FILL FILL_4_OAI21X1_10 ( );
FILL FILL_5_OAI21X1_10 ( );
FILL FILL_6_OAI21X1_10 ( );
FILL FILL_7_OAI21X1_10 ( );
FILL FILL_8_OAI21X1_10 ( );
FILL FILL_9_OAI21X1_10 ( );
FILL FILL_0_DFFPOSX1_3 ( );
FILL FILL_1_DFFPOSX1_3 ( );
FILL FILL_2_DFFPOSX1_3 ( );
FILL FILL_3_DFFPOSX1_3 ( );
FILL FILL_4_DFFPOSX1_3 ( );
FILL FILL_5_DFFPOSX1_3 ( );
FILL FILL_6_DFFPOSX1_3 ( );
FILL FILL_7_DFFPOSX1_3 ( );
FILL FILL_8_DFFPOSX1_3 ( );
FILL FILL_9_DFFPOSX1_3 ( );
FILL FILL_10_DFFPOSX1_3 ( );
FILL FILL_11_DFFPOSX1_3 ( );
FILL FILL_12_DFFPOSX1_3 ( );
FILL FILL_13_DFFPOSX1_3 ( );
FILL FILL_14_DFFPOSX1_3 ( );
FILL FILL_15_DFFPOSX1_3 ( );
FILL FILL_16_DFFPOSX1_3 ( );
FILL FILL_17_DFFPOSX1_3 ( );
FILL FILL_18_DFFPOSX1_3 ( );
FILL FILL_19_DFFPOSX1_3 ( );
FILL FILL_20_DFFPOSX1_3 ( );
FILL FILL_21_DFFPOSX1_3 ( );
FILL FILL_22_DFFPOSX1_3 ( );
FILL FILL_23_DFFPOSX1_3 ( );
FILL FILL_24_DFFPOSX1_3 ( );
FILL FILL_25_DFFPOSX1_3 ( );
FILL FILL_26_DFFPOSX1_3 ( );
FILL FILL_27_DFFPOSX1_3 ( );
FILL FILL_0_DFFPOSX1_7 ( );
FILL FILL_1_DFFPOSX1_7 ( );
FILL FILL_2_DFFPOSX1_7 ( );
FILL FILL_3_DFFPOSX1_7 ( );
FILL FILL_4_DFFPOSX1_7 ( );
FILL FILL_5_DFFPOSX1_7 ( );
FILL FILL_6_DFFPOSX1_7 ( );
FILL FILL_7_DFFPOSX1_7 ( );
FILL FILL_8_DFFPOSX1_7 ( );
FILL FILL_9_DFFPOSX1_7 ( );
FILL FILL_10_DFFPOSX1_7 ( );
FILL FILL_11_DFFPOSX1_7 ( );
FILL FILL_12_DFFPOSX1_7 ( );
FILL FILL_13_DFFPOSX1_7 ( );
FILL FILL_14_DFFPOSX1_7 ( );
FILL FILL_15_DFFPOSX1_7 ( );
FILL FILL_16_DFFPOSX1_7 ( );
FILL FILL_17_DFFPOSX1_7 ( );
FILL FILL_18_DFFPOSX1_7 ( );
FILL FILL_19_DFFPOSX1_7 ( );
FILL FILL_20_DFFPOSX1_7 ( );
FILL FILL_21_DFFPOSX1_7 ( );
FILL FILL_22_DFFPOSX1_7 ( );
FILL FILL_23_DFFPOSX1_7 ( );
FILL FILL_24_DFFPOSX1_7 ( );
FILL FILL_25_DFFPOSX1_7 ( );
FILL FILL_26_DFFPOSX1_7 ( );
FILL FILL_27_DFFPOSX1_7 ( );
FILL FILL_0_INVX1_244 ( );
FILL FILL_1_INVX1_244 ( );
FILL FILL_2_INVX1_244 ( );
FILL FILL_3_INVX1_244 ( );
FILL FILL_4_INVX1_244 ( );
FILL FILL_0_OAI21X1_210 ( );
FILL FILL_1_OAI21X1_210 ( );
FILL FILL_2_OAI21X1_210 ( );
FILL FILL_3_OAI21X1_210 ( );
FILL FILL_4_OAI21X1_210 ( );
FILL FILL_5_OAI21X1_210 ( );
FILL FILL_6_OAI21X1_210 ( );
FILL FILL_7_OAI21X1_210 ( );
FILL FILL_8_OAI21X1_210 ( );
FILL FILL_9_OAI21X1_210 ( );
FILL FILL_0_AOI21X1_29 ( );
FILL FILL_1_AOI21X1_29 ( );
FILL FILL_2_AOI21X1_29 ( );
FILL FILL_3_AOI21X1_29 ( );
FILL FILL_4_AOI21X1_29 ( );
FILL FILL_5_AOI21X1_29 ( );
FILL FILL_6_AOI21X1_29 ( );
FILL FILL_7_AOI21X1_29 ( );
FILL FILL_8_AOI21X1_29 ( );
FILL FILL_0_OAI21X1_229 ( );
FILL FILL_1_OAI21X1_229 ( );
FILL FILL_2_OAI21X1_229 ( );
FILL FILL_3_OAI21X1_229 ( );
FILL FILL_4_OAI21X1_229 ( );
FILL FILL_5_OAI21X1_229 ( );
FILL FILL_6_OAI21X1_229 ( );
FILL FILL_7_OAI21X1_229 ( );
FILL FILL_8_OAI21X1_229 ( );
FILL FILL_9_OAI21X1_229 ( );
FILL FILL_0_DFFSR_95 ( );
FILL FILL_1_DFFSR_95 ( );
FILL FILL_2_DFFSR_95 ( );
FILL FILL_3_DFFSR_95 ( );
FILL FILL_4_DFFSR_95 ( );
FILL FILL_5_DFFSR_95 ( );
FILL FILL_6_DFFSR_95 ( );
FILL FILL_7_DFFSR_95 ( );
FILL FILL_8_DFFSR_95 ( );
FILL FILL_9_DFFSR_95 ( );
FILL FILL_10_DFFSR_95 ( );
FILL FILL_11_DFFSR_95 ( );
FILL FILL_12_DFFSR_95 ( );
FILL FILL_13_DFFSR_95 ( );
FILL FILL_14_DFFSR_95 ( );
FILL FILL_15_DFFSR_95 ( );
FILL FILL_16_DFFSR_95 ( );
FILL FILL_17_DFFSR_95 ( );
FILL FILL_18_DFFSR_95 ( );
FILL FILL_19_DFFSR_95 ( );
FILL FILL_20_DFFSR_95 ( );
FILL FILL_21_DFFSR_95 ( );
FILL FILL_22_DFFSR_95 ( );
FILL FILL_23_DFFSR_95 ( );
FILL FILL_24_DFFSR_95 ( );
FILL FILL_25_DFFSR_95 ( );
FILL FILL_26_DFFSR_95 ( );
FILL FILL_27_DFFSR_95 ( );
FILL FILL_28_DFFSR_95 ( );
FILL FILL_29_DFFSR_95 ( );
FILL FILL_30_DFFSR_95 ( );
FILL FILL_31_DFFSR_95 ( );
FILL FILL_32_DFFSR_95 ( );
FILL FILL_33_DFFSR_95 ( );
FILL FILL_34_DFFSR_95 ( );
FILL FILL_35_DFFSR_95 ( );
FILL FILL_36_DFFSR_95 ( );
FILL FILL_37_DFFSR_95 ( );
FILL FILL_38_DFFSR_95 ( );
FILL FILL_39_DFFSR_95 ( );
FILL FILL_40_DFFSR_95 ( );
FILL FILL_41_DFFSR_95 ( );
FILL FILL_42_DFFSR_95 ( );
FILL FILL_43_DFFSR_95 ( );
FILL FILL_44_DFFSR_95 ( );
FILL FILL_45_DFFSR_95 ( );
FILL FILL_46_DFFSR_95 ( );
FILL FILL_47_DFFSR_95 ( );
FILL FILL_48_DFFSR_95 ( );
FILL FILL_49_DFFSR_95 ( );
FILL FILL_50_DFFSR_95 ( );
FILL FILL_0_INVX1_381 ( );
FILL FILL_1_INVX1_381 ( );
FILL FILL_2_INVX1_381 ( );
FILL FILL_3_INVX1_381 ( );
FILL FILL_0_INVX1_380 ( );
FILL FILL_1_INVX1_380 ( );
FILL FILL_2_INVX1_380 ( );
FILL FILL_3_INVX1_380 ( );
FILL FILL_4_INVX1_380 ( );
FILL FILL_0_OAI22X1_61 ( );
FILL FILL_1_OAI22X1_61 ( );
FILL FILL_2_OAI22X1_61 ( );
FILL FILL_3_OAI22X1_61 ( );
FILL FILL_4_OAI22X1_61 ( );
FILL FILL_5_OAI22X1_61 ( );
FILL FILL_6_OAI22X1_61 ( );
FILL FILL_7_OAI22X1_61 ( );
FILL FILL_8_OAI22X1_61 ( );
FILL FILL_9_OAI22X1_61 ( );
FILL FILL_10_OAI22X1_61 ( );
FILL FILL_11_OAI22X1_61 ( );
FILL FILL_0_INVX1_329 ( );
FILL FILL_1_INVX1_329 ( );
FILL FILL_2_INVX1_329 ( );
FILL FILL_3_INVX1_329 ( );
FILL FILL_4_INVX1_329 ( );
FILL FILL_0_CLKBUF1_2 ( );
FILL FILL_1_CLKBUF1_2 ( );
FILL FILL_2_CLKBUF1_2 ( );
FILL FILL_3_CLKBUF1_2 ( );
FILL FILL_4_CLKBUF1_2 ( );
FILL FILL_5_CLKBUF1_2 ( );
FILL FILL_6_CLKBUF1_2 ( );
FILL FILL_7_CLKBUF1_2 ( );
FILL FILL_8_CLKBUF1_2 ( );
FILL FILL_9_CLKBUF1_2 ( );
FILL FILL_10_CLKBUF1_2 ( );
FILL FILL_11_CLKBUF1_2 ( );
FILL FILL_12_CLKBUF1_2 ( );
FILL FILL_13_CLKBUF1_2 ( );
FILL FILL_14_CLKBUF1_2 ( );
FILL FILL_15_CLKBUF1_2 ( );
FILL FILL_16_CLKBUF1_2 ( );
FILL FILL_17_CLKBUF1_2 ( );
FILL FILL_18_CLKBUF1_2 ( );
FILL FILL_19_CLKBUF1_2 ( );
FILL FILL_20_CLKBUF1_2 ( );
FILL FILL_0_INVX1_140 ( );
FILL FILL_1_INVX1_140 ( );
FILL FILL_2_INVX1_140 ( );
FILL FILL_3_INVX1_140 ( );
FILL FILL_4_INVX1_140 ( );
FILL FILL_0_OAI21X1_85 ( );
FILL FILL_1_OAI21X1_85 ( );
FILL FILL_2_OAI21X1_85 ( );
FILL FILL_3_OAI21X1_85 ( );
FILL FILL_4_OAI21X1_85 ( );
FILL FILL_5_OAI21X1_85 ( );
FILL FILL_6_OAI21X1_85 ( );
FILL FILL_7_OAI21X1_85 ( );
FILL FILL_8_OAI21X1_85 ( );
FILL FILL_9_OAI21X1_85 ( );
FILL FILL_0_NAND2X1_85 ( );
FILL FILL_1_NAND2X1_85 ( );
FILL FILL_2_NAND2X1_85 ( );
FILL FILL_3_NAND2X1_85 ( );
FILL FILL_4_NAND2X1_85 ( );
FILL FILL_5_NAND2X1_85 ( );
FILL FILL_6_NAND2X1_85 ( );
FILL FILL_0_INVX1_365 ( );
FILL FILL_1_INVX1_365 ( );
FILL FILL_2_INVX1_365 ( );
FILL FILL_3_INVX1_365 ( );
FILL FILL_0_DFFSR_134 ( );
FILL FILL_1_DFFSR_134 ( );
FILL FILL_2_DFFSR_134 ( );
FILL FILL_3_DFFSR_134 ( );
FILL FILL_4_DFFSR_134 ( );
FILL FILL_5_DFFSR_134 ( );
FILL FILL_6_DFFSR_134 ( );
FILL FILL_7_DFFSR_134 ( );
FILL FILL_8_DFFSR_134 ( );
FILL FILL_9_DFFSR_134 ( );
FILL FILL_10_DFFSR_134 ( );
FILL FILL_11_DFFSR_134 ( );
FILL FILL_12_DFFSR_134 ( );
FILL FILL_13_DFFSR_134 ( );
FILL FILL_14_DFFSR_134 ( );
FILL FILL_15_DFFSR_134 ( );
FILL FILL_16_DFFSR_134 ( );
FILL FILL_17_DFFSR_134 ( );
FILL FILL_18_DFFSR_134 ( );
FILL FILL_19_DFFSR_134 ( );
FILL FILL_20_DFFSR_134 ( );
FILL FILL_21_DFFSR_134 ( );
FILL FILL_22_DFFSR_134 ( );
FILL FILL_23_DFFSR_134 ( );
FILL FILL_24_DFFSR_134 ( );
FILL FILL_25_DFFSR_134 ( );
FILL FILL_26_DFFSR_134 ( );
FILL FILL_27_DFFSR_134 ( );
FILL FILL_28_DFFSR_134 ( );
FILL FILL_29_DFFSR_134 ( );
FILL FILL_30_DFFSR_134 ( );
FILL FILL_31_DFFSR_134 ( );
FILL FILL_32_DFFSR_134 ( );
FILL FILL_33_DFFSR_134 ( );
FILL FILL_34_DFFSR_134 ( );
FILL FILL_35_DFFSR_134 ( );
FILL FILL_36_DFFSR_134 ( );
FILL FILL_37_DFFSR_134 ( );
FILL FILL_38_DFFSR_134 ( );
FILL FILL_39_DFFSR_134 ( );
FILL FILL_40_DFFSR_134 ( );
FILL FILL_41_DFFSR_134 ( );
FILL FILL_42_DFFSR_134 ( );
FILL FILL_43_DFFSR_134 ( );
FILL FILL_44_DFFSR_134 ( );
FILL FILL_45_DFFSR_134 ( );
FILL FILL_46_DFFSR_134 ( );
FILL FILL_47_DFFSR_134 ( );
FILL FILL_48_DFFSR_134 ( );
FILL FILL_49_DFFSR_134 ( );
FILL FILL_50_DFFSR_134 ( );
FILL FILL_0_NAND2X1_278 ( );
FILL FILL_1_NAND2X1_278 ( );
FILL FILL_2_NAND2X1_278 ( );
FILL FILL_3_NAND2X1_278 ( );
FILL FILL_4_NAND2X1_278 ( );
FILL FILL_5_NAND2X1_278 ( );
FILL FILL_6_NAND2X1_278 ( );
FILL FILL_0_AND2X2_16 ( );
FILL FILL_1_AND2X2_16 ( );
FILL FILL_2_AND2X2_16 ( );
FILL FILL_3_AND2X2_16 ( );
FILL FILL_4_AND2X2_16 ( );
FILL FILL_5_AND2X2_16 ( );
FILL FILL_6_AND2X2_16 ( );
FILL FILL_7_AND2X2_16 ( );
FILL FILL_8_AND2X2_16 ( );
FILL FILL_0_INVX1_433 ( );
FILL FILL_1_INVX1_433 ( );
FILL FILL_2_INVX1_433 ( );
FILL FILL_3_INVX1_433 ( );
FILL FILL_4_INVX1_433 ( );
FILL FILL_0_NAND2X1_281 ( );
FILL FILL_1_NAND2X1_281 ( );
FILL FILL_2_NAND2X1_281 ( );
FILL FILL_3_NAND2X1_281 ( );
FILL FILL_4_NAND2X1_281 ( );
FILL FILL_5_NAND2X1_281 ( );
FILL FILL_6_NAND2X1_281 ( );
FILL FILL_0_NAND2X1_280 ( );
FILL FILL_1_NAND2X1_280 ( );
FILL FILL_2_NAND2X1_280 ( );
FILL FILL_3_NAND2X1_280 ( );
FILL FILL_4_NAND2X1_280 ( );
FILL FILL_5_NAND2X1_280 ( );
FILL FILL_6_NAND2X1_280 ( );
FILL FILL_0_NOR2X1_53 ( );
FILL FILL_1_NOR2X1_53 ( );
FILL FILL_2_NOR2X1_53 ( );
FILL FILL_3_NOR2X1_53 ( );
FILL FILL_4_NOR2X1_53 ( );
FILL FILL_5_NOR2X1_53 ( );
FILL FILL_6_NOR2X1_53 ( );
FILL FILL_0_NAND2X1_239 ( );
FILL FILL_1_NAND2X1_239 ( );
FILL FILL_2_NAND2X1_239 ( );
FILL FILL_3_NAND2X1_239 ( );
FILL FILL_4_NAND2X1_239 ( );
FILL FILL_5_NAND2X1_239 ( );
FILL FILL_6_NAND2X1_239 ( );
FILL FILL_0_NOR2X1_23 ( );
FILL FILL_1_NOR2X1_23 ( );
FILL FILL_2_NOR2X1_23 ( );
FILL FILL_3_NOR2X1_23 ( );
FILL FILL_4_NOR2X1_23 ( );
FILL FILL_5_NOR2X1_23 ( );
FILL FILL_6_NOR2X1_23 ( );
FILL FILL_0_NAND3X1_118 ( );
FILL FILL_1_NAND3X1_118 ( );
FILL FILL_2_NAND3X1_118 ( );
FILL FILL_3_NAND3X1_118 ( );
FILL FILL_4_NAND3X1_118 ( );
FILL FILL_5_NAND3X1_118 ( );
FILL FILL_6_NAND3X1_118 ( );
FILL FILL_7_NAND3X1_118 ( );
FILL FILL_8_NAND3X1_118 ( );
FILL FILL_0_INVX1_317 ( );
FILL FILL_1_INVX1_317 ( );
FILL FILL_2_INVX1_317 ( );
FILL FILL_3_INVX1_317 ( );
FILL FILL_4_INVX1_317 ( );
FILL FILL_0_NAND2X1_47 ( );
FILL FILL_1_NAND2X1_47 ( );
FILL FILL_2_NAND2X1_47 ( );
FILL FILL_3_NAND2X1_47 ( );
FILL FILL_4_NAND2X1_47 ( );
FILL FILL_5_NAND2X1_47 ( );
FILL FILL_6_NAND2X1_47 ( );
FILL FILL_0_DFFSR_39 ( );
FILL FILL_1_DFFSR_39 ( );
FILL FILL_2_DFFSR_39 ( );
FILL FILL_3_DFFSR_39 ( );
FILL FILL_4_DFFSR_39 ( );
FILL FILL_5_DFFSR_39 ( );
FILL FILL_6_DFFSR_39 ( );
FILL FILL_7_DFFSR_39 ( );
FILL FILL_8_DFFSR_39 ( );
FILL FILL_9_DFFSR_39 ( );
FILL FILL_10_DFFSR_39 ( );
FILL FILL_11_DFFSR_39 ( );
FILL FILL_12_DFFSR_39 ( );
FILL FILL_13_DFFSR_39 ( );
FILL FILL_14_DFFSR_39 ( );
FILL FILL_15_DFFSR_39 ( );
FILL FILL_16_DFFSR_39 ( );
FILL FILL_17_DFFSR_39 ( );
FILL FILL_18_DFFSR_39 ( );
FILL FILL_19_DFFSR_39 ( );
FILL FILL_20_DFFSR_39 ( );
FILL FILL_21_DFFSR_39 ( );
FILL FILL_22_DFFSR_39 ( );
FILL FILL_23_DFFSR_39 ( );
FILL FILL_24_DFFSR_39 ( );
FILL FILL_25_DFFSR_39 ( );
FILL FILL_26_DFFSR_39 ( );
FILL FILL_27_DFFSR_39 ( );
FILL FILL_28_DFFSR_39 ( );
FILL FILL_29_DFFSR_39 ( );
FILL FILL_30_DFFSR_39 ( );
FILL FILL_31_DFFSR_39 ( );
FILL FILL_32_DFFSR_39 ( );
FILL FILL_33_DFFSR_39 ( );
FILL FILL_34_DFFSR_39 ( );
FILL FILL_35_DFFSR_39 ( );
FILL FILL_36_DFFSR_39 ( );
FILL FILL_37_DFFSR_39 ( );
FILL FILL_38_DFFSR_39 ( );
FILL FILL_39_DFFSR_39 ( );
FILL FILL_40_DFFSR_39 ( );
FILL FILL_41_DFFSR_39 ( );
FILL FILL_42_DFFSR_39 ( );
FILL FILL_43_DFFSR_39 ( );
FILL FILL_44_DFFSR_39 ( );
FILL FILL_45_DFFSR_39 ( );
FILL FILL_46_DFFSR_39 ( );
FILL FILL_47_DFFSR_39 ( );
FILL FILL_48_DFFSR_39 ( );
FILL FILL_49_DFFSR_39 ( );
FILL FILL_50_DFFSR_39 ( );
FILL FILL_51_DFFSR_39 ( );
FILL FILL_0_NAND2X1_25 ( );
FILL FILL_1_NAND2X1_25 ( );
FILL FILL_2_NAND2X1_25 ( );
FILL FILL_3_NAND2X1_25 ( );
FILL FILL_4_NAND2X1_25 ( );
FILL FILL_5_NAND2X1_25 ( );
FILL FILL_6_NAND2X1_25 ( );
FILL FILL_0_NAND2X1_53 ( );
FILL FILL_1_NAND2X1_53 ( );
FILL FILL_2_NAND2X1_53 ( );
FILL FILL_3_NAND2X1_53 ( );
FILL FILL_4_NAND2X1_53 ( );
FILL FILL_5_NAND2X1_53 ( );
FILL FILL_6_NAND2X1_53 ( );
FILL FILL_0_OAI21X1_36 ( );
FILL FILL_1_OAI21X1_36 ( );
FILL FILL_2_OAI21X1_36 ( );
FILL FILL_3_OAI21X1_36 ( );
FILL FILL_4_OAI21X1_36 ( );
FILL FILL_5_OAI21X1_36 ( );
FILL FILL_6_OAI21X1_36 ( );
FILL FILL_7_OAI21X1_36 ( );
FILL FILL_8_OAI21X1_36 ( );
FILL FILL_9_OAI21X1_36 ( );
FILL FILL_0_INVX1_41 ( );
FILL FILL_1_INVX1_41 ( );
FILL FILL_2_INVX1_41 ( );
FILL FILL_3_INVX1_41 ( );
FILL FILL_0_DFFSR_45 ( );
FILL FILL_1_DFFSR_45 ( );
FILL FILL_2_DFFSR_45 ( );
FILL FILL_3_DFFSR_45 ( );
FILL FILL_4_DFFSR_45 ( );
FILL FILL_5_DFFSR_45 ( );
FILL FILL_6_DFFSR_45 ( );
FILL FILL_7_DFFSR_45 ( );
FILL FILL_8_DFFSR_45 ( );
FILL FILL_9_DFFSR_45 ( );
FILL FILL_10_DFFSR_45 ( );
FILL FILL_11_DFFSR_45 ( );
FILL FILL_12_DFFSR_45 ( );
FILL FILL_13_DFFSR_45 ( );
FILL FILL_14_DFFSR_45 ( );
FILL FILL_15_DFFSR_45 ( );
FILL FILL_16_DFFSR_45 ( );
FILL FILL_17_DFFSR_45 ( );
FILL FILL_18_DFFSR_45 ( );
FILL FILL_19_DFFSR_45 ( );
FILL FILL_20_DFFSR_45 ( );
FILL FILL_21_DFFSR_45 ( );
FILL FILL_22_DFFSR_45 ( );
FILL FILL_23_DFFSR_45 ( );
FILL FILL_24_DFFSR_45 ( );
FILL FILL_25_DFFSR_45 ( );
FILL FILL_26_DFFSR_45 ( );
FILL FILL_27_DFFSR_45 ( );
FILL FILL_28_DFFSR_45 ( );
FILL FILL_29_DFFSR_45 ( );
FILL FILL_30_DFFSR_45 ( );
FILL FILL_31_DFFSR_45 ( );
FILL FILL_32_DFFSR_45 ( );
FILL FILL_33_DFFSR_45 ( );
FILL FILL_34_DFFSR_45 ( );
FILL FILL_35_DFFSR_45 ( );
FILL FILL_36_DFFSR_45 ( );
FILL FILL_37_DFFSR_45 ( );
FILL FILL_38_DFFSR_45 ( );
FILL FILL_39_DFFSR_45 ( );
FILL FILL_40_DFFSR_45 ( );
FILL FILL_41_DFFSR_45 ( );
FILL FILL_42_DFFSR_45 ( );
FILL FILL_43_DFFSR_45 ( );
FILL FILL_44_DFFSR_45 ( );
FILL FILL_45_DFFSR_45 ( );
FILL FILL_46_DFFSR_45 ( );
FILL FILL_47_DFFSR_45 ( );
FILL FILL_48_DFFSR_45 ( );
FILL FILL_49_DFFSR_45 ( );
FILL FILL_50_DFFSR_45 ( );
FILL FILL_51_DFFSR_45 ( );
FILL FILL_0_XOR2X1_1 ( );
FILL FILL_1_XOR2X1_1 ( );
FILL FILL_2_XOR2X1_1 ( );
FILL FILL_3_XOR2X1_1 ( );
FILL FILL_4_XOR2X1_1 ( );
FILL FILL_5_XOR2X1_1 ( );
FILL FILL_6_XOR2X1_1 ( );
FILL FILL_7_XOR2X1_1 ( );
FILL FILL_8_XOR2X1_1 ( );
FILL FILL_9_XOR2X1_1 ( );
FILL FILL_10_XOR2X1_1 ( );
FILL FILL_11_XOR2X1_1 ( );
FILL FILL_12_XOR2X1_1 ( );
FILL FILL_13_XOR2X1_1 ( );
FILL FILL_14_XOR2X1_1 ( );
FILL FILL_15_XOR2X1_1 ( );
FILL FILL_0_INVX1_230 ( );
FILL FILL_1_INVX1_230 ( );
FILL FILL_2_INVX1_230 ( );
FILL FILL_3_INVX1_230 ( );
FILL FILL_0_NAND3X1_17 ( );
FILL FILL_1_NAND3X1_17 ( );
FILL FILL_2_NAND3X1_17 ( );
FILL FILL_3_NAND3X1_17 ( );
FILL FILL_4_NAND3X1_17 ( );
FILL FILL_5_NAND3X1_17 ( );
FILL FILL_6_NAND3X1_17 ( );
FILL FILL_7_NAND3X1_17 ( );
FILL FILL_8_NAND3X1_17 ( );
FILL FILL_9_NAND3X1_17 ( );
FILL FILL_0_AOI21X1_3 ( );
FILL FILL_1_AOI21X1_3 ( );
FILL FILL_2_AOI21X1_3 ( );
FILL FILL_3_AOI21X1_3 ( );
FILL FILL_4_AOI21X1_3 ( );
FILL FILL_5_AOI21X1_3 ( );
FILL FILL_6_AOI21X1_3 ( );
FILL FILL_7_AOI21X1_3 ( );
FILL FILL_8_AOI21X1_3 ( );
FILL FILL_9_AOI21X1_3 ( );
FILL FILL_0_OAI22X1_3 ( );
FILL FILL_1_OAI22X1_3 ( );
FILL FILL_2_OAI22X1_3 ( );
FILL FILL_3_OAI22X1_3 ( );
FILL FILL_4_OAI22X1_3 ( );
FILL FILL_5_OAI22X1_3 ( );
FILL FILL_6_OAI22X1_3 ( );
FILL FILL_7_OAI22X1_3 ( );
FILL FILL_8_OAI22X1_3 ( );
FILL FILL_9_OAI22X1_3 ( );
FILL FILL_10_OAI22X1_3 ( );
FILL FILL_0_NAND3X1_61 ( );
FILL FILL_1_NAND3X1_61 ( );
FILL FILL_2_NAND3X1_61 ( );
FILL FILL_3_NAND3X1_61 ( );
FILL FILL_4_NAND3X1_61 ( );
FILL FILL_5_NAND3X1_61 ( );
FILL FILL_6_NAND3X1_61 ( );
FILL FILL_7_NAND3X1_61 ( );
FILL FILL_8_NAND3X1_61 ( );
FILL FILL_0_DFFSR_79 ( );
FILL FILL_1_DFFSR_79 ( );
FILL FILL_2_DFFSR_79 ( );
FILL FILL_3_DFFSR_79 ( );
FILL FILL_4_DFFSR_79 ( );
FILL FILL_5_DFFSR_79 ( );
FILL FILL_6_DFFSR_79 ( );
FILL FILL_7_DFFSR_79 ( );
FILL FILL_8_DFFSR_79 ( );
FILL FILL_9_DFFSR_79 ( );
FILL FILL_10_DFFSR_79 ( );
FILL FILL_11_DFFSR_79 ( );
FILL FILL_12_DFFSR_79 ( );
FILL FILL_13_DFFSR_79 ( );
FILL FILL_14_DFFSR_79 ( );
FILL FILL_15_DFFSR_79 ( );
FILL FILL_16_DFFSR_79 ( );
FILL FILL_17_DFFSR_79 ( );
FILL FILL_18_DFFSR_79 ( );
FILL FILL_19_DFFSR_79 ( );
FILL FILL_20_DFFSR_79 ( );
FILL FILL_21_DFFSR_79 ( );
FILL FILL_22_DFFSR_79 ( );
FILL FILL_23_DFFSR_79 ( );
FILL FILL_24_DFFSR_79 ( );
FILL FILL_25_DFFSR_79 ( );
FILL FILL_26_DFFSR_79 ( );
FILL FILL_27_DFFSR_79 ( );
FILL FILL_28_DFFSR_79 ( );
FILL FILL_29_DFFSR_79 ( );
FILL FILL_30_DFFSR_79 ( );
FILL FILL_31_DFFSR_79 ( );
FILL FILL_32_DFFSR_79 ( );
FILL FILL_33_DFFSR_79 ( );
FILL FILL_34_DFFSR_79 ( );
FILL FILL_35_DFFSR_79 ( );
FILL FILL_36_DFFSR_79 ( );
FILL FILL_37_DFFSR_79 ( );
FILL FILL_38_DFFSR_79 ( );
FILL FILL_39_DFFSR_79 ( );
FILL FILL_40_DFFSR_79 ( );
FILL FILL_41_DFFSR_79 ( );
FILL FILL_42_DFFSR_79 ( );
FILL FILL_43_DFFSR_79 ( );
FILL FILL_44_DFFSR_79 ( );
FILL FILL_45_DFFSR_79 ( );
FILL FILL_46_DFFSR_79 ( );
FILL FILL_47_DFFSR_79 ( );
FILL FILL_48_DFFSR_79 ( );
FILL FILL_49_DFFSR_79 ( );
FILL FILL_50_DFFSR_79 ( );
FILL FILL_0_OAI22X1_50 ( );
FILL FILL_1_OAI22X1_50 ( );
FILL FILL_2_OAI22X1_50 ( );
FILL FILL_3_OAI22X1_50 ( );
FILL FILL_4_OAI22X1_50 ( );
FILL FILL_5_OAI22X1_50 ( );
FILL FILL_6_OAI22X1_50 ( );
FILL FILL_7_OAI22X1_50 ( );
FILL FILL_8_OAI22X1_50 ( );
FILL FILL_9_OAI22X1_50 ( );
FILL FILL_10_OAI22X1_50 ( );
FILL FILL_11_OAI22X1_50 ( );
FILL FILL_0_INVX1_359 ( );
FILL FILL_1_INVX1_359 ( );
FILL FILL_2_INVX1_359 ( );
FILL FILL_3_INVX1_359 ( );
FILL FILL_0_INVX1_368 ( );
FILL FILL_1_INVX1_368 ( );
FILL FILL_2_INVX1_368 ( );
FILL FILL_3_INVX1_368 ( );
FILL FILL_4_INVX1_368 ( );
FILL FILL_0_OAI22X1_55 ( );
FILL FILL_1_OAI22X1_55 ( );
FILL FILL_2_OAI22X1_55 ( );
FILL FILL_3_OAI22X1_55 ( );
FILL FILL_4_OAI22X1_55 ( );
FILL FILL_5_OAI22X1_55 ( );
FILL FILL_6_OAI22X1_55 ( );
FILL FILL_7_OAI22X1_55 ( );
FILL FILL_8_OAI22X1_55 ( );
FILL FILL_9_OAI22X1_55 ( );
FILL FILL_10_OAI22X1_55 ( );
FILL FILL_11_OAI22X1_55 ( );
FILL FILL_0_NAND2X1_124 ( );
FILL FILL_1_NAND2X1_124 ( );
FILL FILL_2_NAND2X1_124 ( );
FILL FILL_3_NAND2X1_124 ( );
FILL FILL_4_NAND2X1_124 ( );
FILL FILL_5_NAND2X1_124 ( );
FILL FILL_6_NAND2X1_124 ( );
FILL FILL_0_OAI21X1_124 ( );
FILL FILL_1_OAI21X1_124 ( );
FILL FILL_2_OAI21X1_124 ( );
FILL FILL_3_OAI21X1_124 ( );
FILL FILL_4_OAI21X1_124 ( );
FILL FILL_5_OAI21X1_124 ( );
FILL FILL_6_OAI21X1_124 ( );
FILL FILL_7_OAI21X1_124 ( );
FILL FILL_8_OAI21X1_124 ( );
FILL FILL_0_INVX1_96 ( );
FILL FILL_1_INVX1_96 ( );
FILL FILL_2_INVX1_96 ( );
FILL FILL_3_INVX1_96 ( );
FILL FILL_0_NAND2X1_142 ( );
FILL FILL_1_NAND2X1_142 ( );
FILL FILL_2_NAND2X1_142 ( );
FILL FILL_3_NAND2X1_142 ( );
FILL FILL_4_NAND2X1_142 ( );
FILL FILL_5_NAND2X1_142 ( );
FILL FILL_6_NAND2X1_142 ( );
FILL FILL_0_NAND2X1_77 ( );
FILL FILL_1_NAND2X1_77 ( );
FILL FILL_2_NAND2X1_77 ( );
FILL FILL_3_NAND2X1_77 ( );
FILL FILL_4_NAND2X1_77 ( );
FILL FILL_5_NAND2X1_77 ( );
FILL FILL_6_NAND2X1_77 ( );
FILL FILL_0_CLKBUF1_3 ( );
FILL FILL_1_CLKBUF1_3 ( );
FILL FILL_2_CLKBUF1_3 ( );
FILL FILL_3_CLKBUF1_3 ( );
FILL FILL_4_CLKBUF1_3 ( );
FILL FILL_5_CLKBUF1_3 ( );
FILL FILL_6_CLKBUF1_3 ( );
FILL FILL_7_CLKBUF1_3 ( );
FILL FILL_8_CLKBUF1_3 ( );
FILL FILL_9_CLKBUF1_3 ( );
FILL FILL_10_CLKBUF1_3 ( );
FILL FILL_11_CLKBUF1_3 ( );
FILL FILL_12_CLKBUF1_3 ( );
FILL FILL_13_CLKBUF1_3 ( );
FILL FILL_14_CLKBUF1_3 ( );
FILL FILL_15_CLKBUF1_3 ( );
FILL FILL_16_CLKBUF1_3 ( );
FILL FILL_17_CLKBUF1_3 ( );
FILL FILL_18_CLKBUF1_3 ( );
FILL FILL_19_CLKBUF1_3 ( );
FILL FILL_20_CLKBUF1_3 ( );
FILL FILL_21_CLKBUF1_3 ( );
FILL FILL_0_INVX1_158 ( );
FILL FILL_1_INVX1_158 ( );
FILL FILL_2_INVX1_158 ( );
FILL FILL_3_INVX1_158 ( );
FILL FILL_4_INVX1_158 ( );
FILL FILL_0_INVX1_151 ( );
FILL FILL_1_INVX1_151 ( );
FILL FILL_2_INVX1_151 ( );
FILL FILL_3_INVX1_151 ( );
FILL FILL_0_OAI21X1_134 ( );
FILL FILL_1_OAI21X1_134 ( );
FILL FILL_2_OAI21X1_134 ( );
FILL FILL_3_OAI21X1_134 ( );
FILL FILL_4_OAI21X1_134 ( );
FILL FILL_5_OAI21X1_134 ( );
FILL FILL_6_OAI21X1_134 ( );
FILL FILL_7_OAI21X1_134 ( );
FILL FILL_8_OAI21X1_134 ( );
FILL FILL_9_OAI21X1_134 ( );
FILL FILL_0_NAND2X1_134 ( );
FILL FILL_1_NAND2X1_134 ( );
FILL FILL_2_NAND2X1_134 ( );
FILL FILL_3_NAND2X1_134 ( );
FILL FILL_4_NAND2X1_134 ( );
FILL FILL_5_NAND2X1_134 ( );
FILL FILL_6_NAND2X1_134 ( );
FILL FILL_0_NAND2X1_16 ( );
FILL FILL_1_NAND2X1_16 ( );
FILL FILL_2_NAND2X1_16 ( );
FILL FILL_3_NAND2X1_16 ( );
FILL FILL_4_NAND2X1_16 ( );
FILL FILL_5_NAND2X1_16 ( );
FILL FILL_6_NAND2X1_16 ( );
FILL FILL_0_OAI21X1_261 ( );
FILL FILL_1_OAI21X1_261 ( );
FILL FILL_2_OAI21X1_261 ( );
FILL FILL_3_OAI21X1_261 ( );
FILL FILL_4_OAI21X1_261 ( );
FILL FILL_5_OAI21X1_261 ( );
FILL FILL_6_OAI21X1_261 ( );
FILL FILL_7_OAI21X1_261 ( );
FILL FILL_8_OAI21X1_261 ( );
FILL FILL_0_XOR2X1_15 ( );
FILL FILL_1_XOR2X1_15 ( );
FILL FILL_2_XOR2X1_15 ( );
FILL FILL_3_XOR2X1_15 ( );
FILL FILL_4_XOR2X1_15 ( );
FILL FILL_5_XOR2X1_15 ( );
FILL FILL_6_XOR2X1_15 ( );
FILL FILL_7_XOR2X1_15 ( );
FILL FILL_8_XOR2X1_15 ( );
FILL FILL_9_XOR2X1_15 ( );
FILL FILL_10_XOR2X1_15 ( );
FILL FILL_11_XOR2X1_15 ( );
FILL FILL_12_XOR2X1_15 ( );
FILL FILL_13_XOR2X1_15 ( );
FILL FILL_14_XOR2X1_15 ( );
FILL FILL_15_XOR2X1_15 ( );
FILL FILL_0_AOI22X1_14 ( );
FILL FILL_1_AOI22X1_14 ( );
FILL FILL_2_AOI22X1_14 ( );
FILL FILL_3_AOI22X1_14 ( );
FILL FILL_4_AOI22X1_14 ( );
FILL FILL_5_AOI22X1_14 ( );
FILL FILL_6_AOI22X1_14 ( );
FILL FILL_7_AOI22X1_14 ( );
FILL FILL_8_AOI22X1_14 ( );
FILL FILL_9_AOI22X1_14 ( );
FILL FILL_10_AOI22X1_14 ( );
FILL FILL_11_AOI22X1_14 ( );
FILL FILL_0_NAND2X1_30 ( );
FILL FILL_1_NAND2X1_30 ( );
FILL FILL_2_NAND2X1_30 ( );
FILL FILL_3_NAND2X1_30 ( );
FILL FILL_4_NAND2X1_30 ( );
FILL FILL_5_NAND2X1_30 ( );
FILL FILL_6_NAND2X1_30 ( );
FILL FILL_0_NOR2X1_52 ( );
FILL FILL_1_NOR2X1_52 ( );
FILL FILL_2_NOR2X1_52 ( );
FILL FILL_3_NOR2X1_52 ( );
FILL FILL_4_NOR2X1_52 ( );
FILL FILL_5_NOR2X1_52 ( );
FILL FILL_6_NOR2X1_52 ( );
FILL FILL_0_OAI22X1_27 ( );
FILL FILL_1_OAI22X1_27 ( );
FILL FILL_2_OAI22X1_27 ( );
FILL FILL_3_OAI22X1_27 ( );
FILL FILL_4_OAI22X1_27 ( );
FILL FILL_5_OAI22X1_27 ( );
FILL FILL_6_OAI22X1_27 ( );
FILL FILL_7_OAI22X1_27 ( );
FILL FILL_8_OAI22X1_27 ( );
FILL FILL_9_OAI22X1_27 ( );
FILL FILL_10_OAI22X1_27 ( );
FILL FILL_0_INVX1_309 ( );
FILL FILL_1_INVX1_309 ( );
FILL FILL_2_INVX1_309 ( );
FILL FILL_3_INVX1_309 ( );
FILL FILL_4_INVX1_309 ( );
FILL FILL_0_INVX1_310 ( );
FILL FILL_1_INVX1_310 ( );
FILL FILL_2_INVX1_310 ( );
FILL FILL_3_INVX1_310 ( );
FILL FILL_4_INVX1_310 ( );
FILL FILL_0_NAND2X1_238 ( );
FILL FILL_1_NAND2X1_238 ( );
FILL FILL_2_NAND2X1_238 ( );
FILL FILL_3_NAND2X1_238 ( );
FILL FILL_4_NAND2X1_238 ( );
FILL FILL_5_NAND2X1_238 ( );
FILL FILL_6_NAND2X1_238 ( );
FILL FILL_0_INVX1_44 ( );
FILL FILL_1_INVX1_44 ( );
FILL FILL_2_INVX1_44 ( );
FILL FILL_3_INVX1_44 ( );
FILL FILL_0_NOR2X1_21 ( );
FILL FILL_1_NOR2X1_21 ( );
FILL FILL_2_NOR2X1_21 ( );
FILL FILL_3_NOR2X1_21 ( );
FILL FILL_4_NOR2X1_21 ( );
FILL FILL_5_NOR2X1_21 ( );
FILL FILL_6_NOR2X1_21 ( );
FILL FILL_0_OAI22X1_24 ( );
FILL FILL_1_OAI22X1_24 ( );
FILL FILL_2_OAI22X1_24 ( );
FILL FILL_3_OAI22X1_24 ( );
FILL FILL_4_OAI22X1_24 ( );
FILL FILL_5_OAI22X1_24 ( );
FILL FILL_6_OAI22X1_24 ( );
FILL FILL_7_OAI22X1_24 ( );
FILL FILL_8_OAI22X1_24 ( );
FILL FILL_9_OAI22X1_24 ( );
FILL FILL_10_OAI22X1_24 ( );
FILL FILL_0_INVX1_270 ( );
FILL FILL_1_INVX1_270 ( );
FILL FILL_2_INVX1_270 ( );
FILL FILL_3_INVX1_270 ( );
FILL FILL_4_INVX1_270 ( );
FILL FILL_0_INVX1_304 ( );
FILL FILL_1_INVX1_304 ( );
FILL FILL_2_INVX1_304 ( );
FILL FILL_3_INVX1_304 ( );
FILL FILL_4_INVX1_304 ( );
FILL FILL_0_DFFSR_36 ( );
FILL FILL_1_DFFSR_36 ( );
FILL FILL_2_DFFSR_36 ( );
FILL FILL_3_DFFSR_36 ( );
FILL FILL_4_DFFSR_36 ( );
FILL FILL_5_DFFSR_36 ( );
FILL FILL_6_DFFSR_36 ( );
FILL FILL_7_DFFSR_36 ( );
FILL FILL_8_DFFSR_36 ( );
FILL FILL_9_DFFSR_36 ( );
FILL FILL_10_DFFSR_36 ( );
FILL FILL_11_DFFSR_36 ( );
FILL FILL_12_DFFSR_36 ( );
FILL FILL_13_DFFSR_36 ( );
FILL FILL_14_DFFSR_36 ( );
FILL FILL_15_DFFSR_36 ( );
FILL FILL_16_DFFSR_36 ( );
FILL FILL_17_DFFSR_36 ( );
FILL FILL_18_DFFSR_36 ( );
FILL FILL_19_DFFSR_36 ( );
FILL FILL_20_DFFSR_36 ( );
FILL FILL_21_DFFSR_36 ( );
FILL FILL_22_DFFSR_36 ( );
FILL FILL_23_DFFSR_36 ( );
FILL FILL_24_DFFSR_36 ( );
FILL FILL_25_DFFSR_36 ( );
FILL FILL_26_DFFSR_36 ( );
FILL FILL_27_DFFSR_36 ( );
FILL FILL_28_DFFSR_36 ( );
FILL FILL_29_DFFSR_36 ( );
FILL FILL_30_DFFSR_36 ( );
FILL FILL_31_DFFSR_36 ( );
FILL FILL_32_DFFSR_36 ( );
FILL FILL_33_DFFSR_36 ( );
FILL FILL_34_DFFSR_36 ( );
FILL FILL_35_DFFSR_36 ( );
FILL FILL_36_DFFSR_36 ( );
FILL FILL_37_DFFSR_36 ( );
FILL FILL_38_DFFSR_36 ( );
FILL FILL_39_DFFSR_36 ( );
FILL FILL_40_DFFSR_36 ( );
FILL FILL_41_DFFSR_36 ( );
FILL FILL_42_DFFSR_36 ( );
FILL FILL_43_DFFSR_36 ( );
FILL FILL_44_DFFSR_36 ( );
FILL FILL_45_DFFSR_36 ( );
FILL FILL_46_DFFSR_36 ( );
FILL FILL_47_DFFSR_36 ( );
FILL FILL_48_DFFSR_36 ( );
FILL FILL_49_DFFSR_36 ( );
FILL FILL_50_DFFSR_36 ( );
FILL FILL_51_DFFSR_36 ( );
FILL FILL_0_OAI21X1_45 ( );
FILL FILL_1_OAI21X1_45 ( );
FILL FILL_2_OAI21X1_45 ( );
FILL FILL_3_OAI21X1_45 ( );
FILL FILL_4_OAI21X1_45 ( );
FILL FILL_5_OAI21X1_45 ( );
FILL FILL_6_OAI21X1_45 ( );
FILL FILL_7_OAI21X1_45 ( );
FILL FILL_8_OAI21X1_45 ( );
FILL FILL_0_INVX1_51 ( );
FILL FILL_1_INVX1_51 ( );
FILL FILL_2_INVX1_51 ( );
FILL FILL_3_INVX1_51 ( );
FILL FILL_4_INVX1_51 ( );
FILL FILL_0_DFFSR_167 ( );
FILL FILL_1_DFFSR_167 ( );
FILL FILL_2_DFFSR_167 ( );
FILL FILL_3_DFFSR_167 ( );
FILL FILL_4_DFFSR_167 ( );
FILL FILL_5_DFFSR_167 ( );
FILL FILL_6_DFFSR_167 ( );
FILL FILL_7_DFFSR_167 ( );
FILL FILL_8_DFFSR_167 ( );
FILL FILL_9_DFFSR_167 ( );
FILL FILL_10_DFFSR_167 ( );
FILL FILL_11_DFFSR_167 ( );
FILL FILL_12_DFFSR_167 ( );
FILL FILL_13_DFFSR_167 ( );
FILL FILL_14_DFFSR_167 ( );
FILL FILL_15_DFFSR_167 ( );
FILL FILL_16_DFFSR_167 ( );
FILL FILL_17_DFFSR_167 ( );
FILL FILL_18_DFFSR_167 ( );
FILL FILL_19_DFFSR_167 ( );
FILL FILL_20_DFFSR_167 ( );
FILL FILL_21_DFFSR_167 ( );
FILL FILL_22_DFFSR_167 ( );
FILL FILL_23_DFFSR_167 ( );
FILL FILL_24_DFFSR_167 ( );
FILL FILL_25_DFFSR_167 ( );
FILL FILL_26_DFFSR_167 ( );
FILL FILL_27_DFFSR_167 ( );
FILL FILL_28_DFFSR_167 ( );
FILL FILL_29_DFFSR_167 ( );
FILL FILL_30_DFFSR_167 ( );
FILL FILL_31_DFFSR_167 ( );
FILL FILL_32_DFFSR_167 ( );
FILL FILL_33_DFFSR_167 ( );
FILL FILL_34_DFFSR_167 ( );
FILL FILL_35_DFFSR_167 ( );
FILL FILL_36_DFFSR_167 ( );
FILL FILL_37_DFFSR_167 ( );
FILL FILL_38_DFFSR_167 ( );
FILL FILL_39_DFFSR_167 ( );
FILL FILL_40_DFFSR_167 ( );
FILL FILL_41_DFFSR_167 ( );
FILL FILL_42_DFFSR_167 ( );
FILL FILL_43_DFFSR_167 ( );
FILL FILL_44_DFFSR_167 ( );
FILL FILL_45_DFFSR_167 ( );
FILL FILL_46_DFFSR_167 ( );
FILL FILL_47_DFFSR_167 ( );
FILL FILL_48_DFFSR_167 ( );
FILL FILL_49_DFFSR_167 ( );
FILL FILL_50_DFFSR_167 ( );
FILL FILL_51_DFFSR_167 ( );
FILL FILL_0_INVX1_412 ( );
FILL FILL_1_INVX1_412 ( );
FILL FILL_2_INVX1_412 ( );
FILL FILL_3_INVX1_412 ( );
FILL FILL_0_OAI21X1_250 ( );
FILL FILL_1_OAI21X1_250 ( );
FILL FILL_2_OAI21X1_250 ( );
FILL FILL_3_OAI21X1_250 ( );
FILL FILL_4_OAI21X1_250 ( );
FILL FILL_5_OAI21X1_250 ( );
FILL FILL_6_OAI21X1_250 ( );
FILL FILL_7_OAI21X1_250 ( );
FILL FILL_8_OAI21X1_250 ( );
FILL FILL_9_OAI21X1_250 ( );
FILL FILL_0_DFFPOSX1_8 ( );
FILL FILL_1_DFFPOSX1_8 ( );
FILL FILL_2_DFFPOSX1_8 ( );
FILL FILL_3_DFFPOSX1_8 ( );
FILL FILL_4_DFFPOSX1_8 ( );
FILL FILL_5_DFFPOSX1_8 ( );
FILL FILL_6_DFFPOSX1_8 ( );
FILL FILL_7_DFFPOSX1_8 ( );
FILL FILL_8_DFFPOSX1_8 ( );
FILL FILL_9_DFFPOSX1_8 ( );
FILL FILL_10_DFFPOSX1_8 ( );
FILL FILL_11_DFFPOSX1_8 ( );
FILL FILL_12_DFFPOSX1_8 ( );
FILL FILL_13_DFFPOSX1_8 ( );
FILL FILL_14_DFFPOSX1_8 ( );
FILL FILL_15_DFFPOSX1_8 ( );
FILL FILL_16_DFFPOSX1_8 ( );
FILL FILL_17_DFFPOSX1_8 ( );
FILL FILL_18_DFFPOSX1_8 ( );
FILL FILL_19_DFFPOSX1_8 ( );
FILL FILL_20_DFFPOSX1_8 ( );
FILL FILL_21_DFFPOSX1_8 ( );
FILL FILL_22_DFFPOSX1_8 ( );
FILL FILL_23_DFFPOSX1_8 ( );
FILL FILL_24_DFFPOSX1_8 ( );
FILL FILL_25_DFFPOSX1_8 ( );
FILL FILL_26_DFFPOSX1_8 ( );
FILL FILL_27_DFFPOSX1_8 ( );
FILL FILL_0_NAND2X1_95 ( );
FILL FILL_1_NAND2X1_95 ( );
FILL FILL_2_NAND2X1_95 ( );
FILL FILL_3_NAND2X1_95 ( );
FILL FILL_4_NAND2X1_95 ( );
FILL FILL_5_NAND2X1_95 ( );
FILL FILL_6_NAND2X1_95 ( );
FILL FILL_0_OAI21X1_95 ( );
FILL FILL_1_OAI21X1_95 ( );
FILL FILL_2_OAI21X1_95 ( );
FILL FILL_3_OAI21X1_95 ( );
FILL FILL_4_OAI21X1_95 ( );
FILL FILL_5_OAI21X1_95 ( );
FILL FILL_6_OAI21X1_95 ( );
FILL FILL_7_OAI21X1_95 ( );
FILL FILL_8_OAI21X1_95 ( );
FILL FILL_0_INVX1_107 ( );
FILL FILL_1_INVX1_107 ( );
FILL FILL_2_INVX1_107 ( );
FILL FILL_3_INVX1_107 ( );
FILL FILL_4_INVX1_107 ( );
FILL FILL_0_NAND2X1_79 ( );
FILL FILL_1_NAND2X1_79 ( );
FILL FILL_2_NAND2X1_79 ( );
FILL FILL_3_NAND2X1_79 ( );
FILL FILL_4_NAND2X1_79 ( );
FILL FILL_5_NAND2X1_79 ( );
FILL FILL_6_NAND2X1_79 ( );
FILL FILL_0_OAI21X1_79 ( );
FILL FILL_1_OAI21X1_79 ( );
FILL FILL_2_OAI21X1_79 ( );
FILL FILL_3_OAI21X1_79 ( );
FILL FILL_4_OAI21X1_79 ( );
FILL FILL_5_OAI21X1_79 ( );
FILL FILL_6_OAI21X1_79 ( );
FILL FILL_7_OAI21X1_79 ( );
FILL FILL_8_OAI21X1_79 ( );
FILL FILL_0_OAI21X1_114 ( );
FILL FILL_1_OAI21X1_114 ( );
FILL FILL_2_OAI21X1_114 ( );
FILL FILL_3_OAI21X1_114 ( );
FILL FILL_4_OAI21X1_114 ( );
FILL FILL_5_OAI21X1_114 ( );
FILL FILL_6_OAI21X1_114 ( );
FILL FILL_7_OAI21X1_114 ( );
FILL FILL_8_OAI21X1_114 ( );
FILL FILL_0_INVX1_129 ( );
FILL FILL_1_INVX1_129 ( );
FILL FILL_2_INVX1_129 ( );
FILL FILL_3_INVX1_129 ( );
FILL FILL_4_INVX1_129 ( );
FILL FILL_0_INVX1_131 ( );
FILL FILL_1_INVX1_131 ( );
FILL FILL_2_INVX1_131 ( );
FILL FILL_3_INVX1_131 ( );
FILL FILL_4_INVX1_131 ( );
FILL FILL_0_INVX1_358 ( );
FILL FILL_1_INVX1_358 ( );
FILL FILL_2_INVX1_358 ( );
FILL FILL_3_INVX1_358 ( );
FILL FILL_4_INVX1_358 ( );
FILL FILL_0_NAND2X1_116 ( );
FILL FILL_1_NAND2X1_116 ( );
FILL FILL_2_NAND2X1_116 ( );
FILL FILL_3_NAND2X1_116 ( );
FILL FILL_4_NAND2X1_116 ( );
FILL FILL_5_NAND2X1_116 ( );
FILL FILL_6_NAND2X1_116 ( );
FILL FILL_0_DFFSR_124 ( );
FILL FILL_1_DFFSR_124 ( );
FILL FILL_2_DFFSR_124 ( );
FILL FILL_3_DFFSR_124 ( );
FILL FILL_4_DFFSR_124 ( );
FILL FILL_5_DFFSR_124 ( );
FILL FILL_6_DFFSR_124 ( );
FILL FILL_7_DFFSR_124 ( );
FILL FILL_8_DFFSR_124 ( );
FILL FILL_9_DFFSR_124 ( );
FILL FILL_10_DFFSR_124 ( );
FILL FILL_11_DFFSR_124 ( );
FILL FILL_12_DFFSR_124 ( );
FILL FILL_13_DFFSR_124 ( );
FILL FILL_14_DFFSR_124 ( );
FILL FILL_15_DFFSR_124 ( );
FILL FILL_16_DFFSR_124 ( );
FILL FILL_17_DFFSR_124 ( );
FILL FILL_18_DFFSR_124 ( );
FILL FILL_19_DFFSR_124 ( );
FILL FILL_20_DFFSR_124 ( );
FILL FILL_21_DFFSR_124 ( );
FILL FILL_22_DFFSR_124 ( );
FILL FILL_23_DFFSR_124 ( );
FILL FILL_24_DFFSR_124 ( );
FILL FILL_25_DFFSR_124 ( );
FILL FILL_26_DFFSR_124 ( );
FILL FILL_27_DFFSR_124 ( );
FILL FILL_28_DFFSR_124 ( );
FILL FILL_29_DFFSR_124 ( );
FILL FILL_30_DFFSR_124 ( );
FILL FILL_31_DFFSR_124 ( );
FILL FILL_32_DFFSR_124 ( );
FILL FILL_33_DFFSR_124 ( );
FILL FILL_34_DFFSR_124 ( );
FILL FILL_35_DFFSR_124 ( );
FILL FILL_36_DFFSR_124 ( );
FILL FILL_37_DFFSR_124 ( );
FILL FILL_38_DFFSR_124 ( );
FILL FILL_39_DFFSR_124 ( );
FILL FILL_40_DFFSR_124 ( );
FILL FILL_41_DFFSR_124 ( );
FILL FILL_42_DFFSR_124 ( );
FILL FILL_43_DFFSR_124 ( );
FILL FILL_44_DFFSR_124 ( );
FILL FILL_45_DFFSR_124 ( );
FILL FILL_46_DFFSR_124 ( );
FILL FILL_47_DFFSR_124 ( );
FILL FILL_48_DFFSR_124 ( );
FILL FILL_49_DFFSR_124 ( );
FILL FILL_50_DFFSR_124 ( );
FILL FILL_0_INVX1_397 ( );
FILL FILL_1_INVX1_397 ( );
FILL FILL_2_INVX1_397 ( );
FILL FILL_3_INVX1_397 ( );
FILL FILL_0_INVX1_87 ( );
FILL FILL_1_INVX1_87 ( );
FILL FILL_2_INVX1_87 ( );
FILL FILL_3_INVX1_87 ( );
FILL FILL_4_INVX1_87 ( );
FILL FILL_0_OAI21X1_77 ( );
FILL FILL_1_OAI21X1_77 ( );
FILL FILL_2_OAI21X1_77 ( );
FILL FILL_3_OAI21X1_77 ( );
FILL FILL_4_OAI21X1_77 ( );
FILL FILL_5_OAI21X1_77 ( );
FILL FILL_6_OAI21X1_77 ( );
FILL FILL_7_OAI21X1_77 ( );
FILL FILL_8_OAI21X1_77 ( );
FILL FILL_0_INVX1_430 ( );
FILL FILL_1_INVX1_430 ( );
FILL FILL_2_INVX1_430 ( );
FILL FILL_3_INVX1_430 ( );
FILL FILL_4_INVX1_430 ( );
FILL FILL_0_NOR2X1_49 ( );
FILL FILL_1_NOR2X1_49 ( );
FILL FILL_2_NOR2X1_49 ( );
FILL FILL_3_NOR2X1_49 ( );
FILL FILL_4_NOR2X1_49 ( );
FILL FILL_5_NOR2X1_49 ( );
FILL FILL_6_NOR2X1_49 ( );
FILL FILL_0_OAI21X1_16 ( );
FILL FILL_1_OAI21X1_16 ( );
FILL FILL_2_OAI21X1_16 ( );
FILL FILL_3_OAI21X1_16 ( );
FILL FILL_4_OAI21X1_16 ( );
FILL FILL_5_OAI21X1_16 ( );
FILL FILL_6_OAI21X1_16 ( );
FILL FILL_7_OAI21X1_16 ( );
FILL FILL_8_OAI21X1_16 ( );
FILL FILL_9_OAI21X1_16 ( );
FILL FILL_0_NOR2X1_48 ( );
FILL FILL_1_NOR2X1_48 ( );
FILL FILL_2_NOR2X1_48 ( );
FILL FILL_3_NOR2X1_48 ( );
FILL FILL_4_NOR2X1_48 ( );
FILL FILL_5_NOR2X1_48 ( );
FILL FILL_6_NOR2X1_48 ( );
FILL FILL_0_NOR2X1_50 ( );
FILL FILL_1_NOR2X1_50 ( );
FILL FILL_2_NOR2X1_50 ( );
FILL FILL_3_NOR2X1_50 ( );
FILL FILL_4_NOR2X1_50 ( );
FILL FILL_5_NOR2X1_50 ( );
FILL FILL_6_NOR2X1_50 ( );
FILL FILL_0_INVX1_431 ( );
FILL FILL_1_INVX1_431 ( );
FILL FILL_2_INVX1_431 ( );
FILL FILL_3_INVX1_431 ( );
FILL FILL_0_AOI21X1_45 ( );
FILL FILL_1_AOI21X1_45 ( );
FILL FILL_2_AOI21X1_45 ( );
FILL FILL_3_AOI21X1_45 ( );
FILL FILL_4_AOI21X1_45 ( );
FILL FILL_5_AOI21X1_45 ( );
FILL FILL_6_AOI21X1_45 ( );
FILL FILL_7_AOI21X1_45 ( );
FILL FILL_8_AOI21X1_45 ( );
FILL FILL_9_AOI21X1_45 ( );
FILL FILL_0_OAI21X1_262 ( );
FILL FILL_1_OAI21X1_262 ( );
FILL FILL_2_OAI21X1_262 ( );
FILL FILL_3_OAI21X1_262 ( );
FILL FILL_4_OAI21X1_262 ( );
FILL FILL_5_OAI21X1_262 ( );
FILL FILL_6_OAI21X1_262 ( );
FILL FILL_7_OAI21X1_262 ( );
FILL FILL_8_OAI21X1_262 ( );
FILL FILL_0_INVX1_436 ( );
FILL FILL_1_INVX1_436 ( );
FILL FILL_2_INVX1_436 ( );
FILL FILL_3_INVX1_436 ( );
FILL FILL_4_INVX1_436 ( );
FILL FILL_0_NAND2X1_283 ( );
FILL FILL_1_NAND2X1_283 ( );
FILL FILL_2_NAND2X1_283 ( );
FILL FILL_3_NAND2X1_283 ( );
FILL FILL_4_NAND2X1_283 ( );
FILL FILL_5_NAND2X1_283 ( );
FILL FILL_6_NAND2X1_283 ( );
FILL FILL_0_NOR2X1_51 ( );
FILL FILL_1_NOR2X1_51 ( );
FILL FILL_2_NOR2X1_51 ( );
FILL FILL_3_NOR2X1_51 ( );
FILL FILL_4_NOR2X1_51 ( );
FILL FILL_5_NOR2X1_51 ( );
FILL FILL_6_NOR2X1_51 ( );
FILL FILL_0_DFFSR_55 ( );
FILL FILL_1_DFFSR_55 ( );
FILL FILL_2_DFFSR_55 ( );
FILL FILL_3_DFFSR_55 ( );
FILL FILL_4_DFFSR_55 ( );
FILL FILL_5_DFFSR_55 ( );
FILL FILL_6_DFFSR_55 ( );
FILL FILL_7_DFFSR_55 ( );
FILL FILL_8_DFFSR_55 ( );
FILL FILL_9_DFFSR_55 ( );
FILL FILL_10_DFFSR_55 ( );
FILL FILL_11_DFFSR_55 ( );
FILL FILL_12_DFFSR_55 ( );
FILL FILL_13_DFFSR_55 ( );
FILL FILL_14_DFFSR_55 ( );
FILL FILL_15_DFFSR_55 ( );
FILL FILL_16_DFFSR_55 ( );
FILL FILL_17_DFFSR_55 ( );
FILL FILL_18_DFFSR_55 ( );
FILL FILL_19_DFFSR_55 ( );
FILL FILL_20_DFFSR_55 ( );
FILL FILL_21_DFFSR_55 ( );
FILL FILL_22_DFFSR_55 ( );
FILL FILL_23_DFFSR_55 ( );
FILL FILL_24_DFFSR_55 ( );
FILL FILL_25_DFFSR_55 ( );
FILL FILL_26_DFFSR_55 ( );
FILL FILL_27_DFFSR_55 ( );
FILL FILL_28_DFFSR_55 ( );
FILL FILL_29_DFFSR_55 ( );
FILL FILL_30_DFFSR_55 ( );
FILL FILL_31_DFFSR_55 ( );
FILL FILL_32_DFFSR_55 ( );
FILL FILL_33_DFFSR_55 ( );
FILL FILL_34_DFFSR_55 ( );
FILL FILL_35_DFFSR_55 ( );
FILL FILL_36_DFFSR_55 ( );
FILL FILL_37_DFFSR_55 ( );
FILL FILL_38_DFFSR_55 ( );
FILL FILL_39_DFFSR_55 ( );
FILL FILL_40_DFFSR_55 ( );
FILL FILL_41_DFFSR_55 ( );
FILL FILL_42_DFFSR_55 ( );
FILL FILL_43_DFFSR_55 ( );
FILL FILL_44_DFFSR_55 ( );
FILL FILL_45_DFFSR_55 ( );
FILL FILL_46_DFFSR_55 ( );
FILL FILL_47_DFFSR_55 ( );
FILL FILL_48_DFFSR_55 ( );
FILL FILL_49_DFFSR_55 ( );
FILL FILL_50_DFFSR_55 ( );
FILL FILL_0_INVX1_299 ( );
FILL FILL_1_INVX1_299 ( );
FILL FILL_2_INVX1_299 ( );
FILL FILL_3_INVX1_299 ( );
FILL FILL_4_INVX1_299 ( );
FILL FILL_0_OAI21X1_30 ( );
FILL FILL_1_OAI21X1_30 ( );
FILL FILL_2_OAI21X1_30 ( );
FILL FILL_3_OAI21X1_30 ( );
FILL FILL_4_OAI21X1_30 ( );
FILL FILL_5_OAI21X1_30 ( );
FILL FILL_6_OAI21X1_30 ( );
FILL FILL_7_OAI21X1_30 ( );
FILL FILL_8_OAI21X1_30 ( );
FILL FILL_0_INVX1_34 ( );
FILL FILL_1_INVX1_34 ( );
FILL FILL_2_INVX1_34 ( );
FILL FILL_3_INVX1_34 ( );
FILL FILL_4_INVX1_34 ( );
FILL FILL_0_DFFSR_30 ( );
FILL FILL_1_DFFSR_30 ( );
FILL FILL_2_DFFSR_30 ( );
FILL FILL_3_DFFSR_30 ( );
FILL FILL_4_DFFSR_30 ( );
FILL FILL_5_DFFSR_30 ( );
FILL FILL_6_DFFSR_30 ( );
FILL FILL_7_DFFSR_30 ( );
FILL FILL_8_DFFSR_30 ( );
FILL FILL_9_DFFSR_30 ( );
FILL FILL_10_DFFSR_30 ( );
FILL FILL_11_DFFSR_30 ( );
FILL FILL_12_DFFSR_30 ( );
FILL FILL_13_DFFSR_30 ( );
FILL FILL_14_DFFSR_30 ( );
FILL FILL_15_DFFSR_30 ( );
FILL FILL_16_DFFSR_30 ( );
FILL FILL_17_DFFSR_30 ( );
FILL FILL_18_DFFSR_30 ( );
FILL FILL_19_DFFSR_30 ( );
FILL FILL_20_DFFSR_30 ( );
FILL FILL_21_DFFSR_30 ( );
FILL FILL_22_DFFSR_30 ( );
FILL FILL_23_DFFSR_30 ( );
FILL FILL_24_DFFSR_30 ( );
FILL FILL_25_DFFSR_30 ( );
FILL FILL_26_DFFSR_30 ( );
FILL FILL_27_DFFSR_30 ( );
FILL FILL_28_DFFSR_30 ( );
FILL FILL_29_DFFSR_30 ( );
FILL FILL_30_DFFSR_30 ( );
FILL FILL_31_DFFSR_30 ( );
FILL FILL_32_DFFSR_30 ( );
FILL FILL_33_DFFSR_30 ( );
FILL FILL_34_DFFSR_30 ( );
FILL FILL_35_DFFSR_30 ( );
FILL FILL_36_DFFSR_30 ( );
FILL FILL_37_DFFSR_30 ( );
FILL FILL_38_DFFSR_30 ( );
FILL FILL_39_DFFSR_30 ( );
FILL FILL_40_DFFSR_30 ( );
FILL FILL_41_DFFSR_30 ( );
FILL FILL_42_DFFSR_30 ( );
FILL FILL_43_DFFSR_30 ( );
FILL FILL_44_DFFSR_30 ( );
FILL FILL_45_DFFSR_30 ( );
FILL FILL_46_DFFSR_30 ( );
FILL FILL_47_DFFSR_30 ( );
FILL FILL_48_DFFSR_30 ( );
FILL FILL_49_DFFSR_30 ( );
FILL FILL_50_DFFSR_30 ( );
FILL FILL_0_NAND2X1_45 ( );
FILL FILL_1_NAND2X1_45 ( );
FILL FILL_2_NAND2X1_45 ( );
FILL FILL_3_NAND2X1_45 ( );
FILL FILL_4_NAND2X1_45 ( );
FILL FILL_5_NAND2X1_45 ( );
FILL FILL_6_NAND2X1_45 ( );
FILL FILL_0_NAND2X1_7 ( );
FILL FILL_1_NAND2X1_7 ( );
FILL FILL_2_NAND2X1_7 ( );
FILL FILL_3_NAND2X1_7 ( );
FILL FILL_4_NAND2X1_7 ( );
FILL FILL_5_NAND2X1_7 ( );
FILL FILL_6_NAND2X1_7 ( );
FILL FILL_0_INVX1_42 ( );
FILL FILL_1_INVX1_42 ( );
FILL FILL_2_INVX1_42 ( );
FILL FILL_3_INVX1_42 ( );
FILL FILL_0_DFFPOSX1_2 ( );
FILL FILL_1_DFFPOSX1_2 ( );
FILL FILL_2_DFFPOSX1_2 ( );
FILL FILL_3_DFFPOSX1_2 ( );
FILL FILL_4_DFFPOSX1_2 ( );
FILL FILL_5_DFFPOSX1_2 ( );
FILL FILL_6_DFFPOSX1_2 ( );
FILL FILL_7_DFFPOSX1_2 ( );
FILL FILL_8_DFFPOSX1_2 ( );
FILL FILL_9_DFFPOSX1_2 ( );
FILL FILL_10_DFFPOSX1_2 ( );
FILL FILL_11_DFFPOSX1_2 ( );
FILL FILL_12_DFFPOSX1_2 ( );
FILL FILL_13_DFFPOSX1_2 ( );
FILL FILL_14_DFFPOSX1_2 ( );
FILL FILL_15_DFFPOSX1_2 ( );
FILL FILL_16_DFFPOSX1_2 ( );
FILL FILL_17_DFFPOSX1_2 ( );
FILL FILL_18_DFFPOSX1_2 ( );
FILL FILL_19_DFFPOSX1_2 ( );
FILL FILL_20_DFFPOSX1_2 ( );
FILL FILL_21_DFFPOSX1_2 ( );
FILL FILL_22_DFFPOSX1_2 ( );
FILL FILL_23_DFFPOSX1_2 ( );
FILL FILL_24_DFFPOSX1_2 ( );
FILL FILL_25_DFFPOSX1_2 ( );
FILL FILL_26_DFFPOSX1_2 ( );
FILL FILL_27_DFFPOSX1_2 ( );
FILL FILL_0_NAND2X1_177 ( );
FILL FILL_1_NAND2X1_177 ( );
FILL FILL_2_NAND2X1_177 ( );
FILL FILL_3_NAND2X1_177 ( );
FILL FILL_4_NAND2X1_177 ( );
FILL FILL_5_NAND2X1_177 ( );
FILL FILL_6_NAND2X1_177 ( );
FILL FILL_0_DFFSR_182 ( );
FILL FILL_1_DFFSR_182 ( );
FILL FILL_2_DFFSR_182 ( );
FILL FILL_3_DFFSR_182 ( );
FILL FILL_4_DFFSR_182 ( );
FILL FILL_5_DFFSR_182 ( );
FILL FILL_6_DFFSR_182 ( );
FILL FILL_7_DFFSR_182 ( );
FILL FILL_8_DFFSR_182 ( );
FILL FILL_9_DFFSR_182 ( );
FILL FILL_10_DFFSR_182 ( );
FILL FILL_11_DFFSR_182 ( );
FILL FILL_12_DFFSR_182 ( );
FILL FILL_13_DFFSR_182 ( );
FILL FILL_14_DFFSR_182 ( );
FILL FILL_15_DFFSR_182 ( );
FILL FILL_16_DFFSR_182 ( );
FILL FILL_17_DFFSR_182 ( );
FILL FILL_18_DFFSR_182 ( );
FILL FILL_19_DFFSR_182 ( );
FILL FILL_20_DFFSR_182 ( );
FILL FILL_21_DFFSR_182 ( );
FILL FILL_22_DFFSR_182 ( );
FILL FILL_23_DFFSR_182 ( );
FILL FILL_24_DFFSR_182 ( );
FILL FILL_25_DFFSR_182 ( );
FILL FILL_26_DFFSR_182 ( );
FILL FILL_27_DFFSR_182 ( );
FILL FILL_28_DFFSR_182 ( );
FILL FILL_29_DFFSR_182 ( );
FILL FILL_30_DFFSR_182 ( );
FILL FILL_31_DFFSR_182 ( );
FILL FILL_32_DFFSR_182 ( );
FILL FILL_33_DFFSR_182 ( );
FILL FILL_34_DFFSR_182 ( );
FILL FILL_35_DFFSR_182 ( );
FILL FILL_36_DFFSR_182 ( );
FILL FILL_37_DFFSR_182 ( );
FILL FILL_38_DFFSR_182 ( );
FILL FILL_39_DFFSR_182 ( );
FILL FILL_40_DFFSR_182 ( );
FILL FILL_41_DFFSR_182 ( );
FILL FILL_42_DFFSR_182 ( );
FILL FILL_43_DFFSR_182 ( );
FILL FILL_44_DFFSR_182 ( );
FILL FILL_45_DFFSR_182 ( );
FILL FILL_46_DFFSR_182 ( );
FILL FILL_47_DFFSR_182 ( );
FILL FILL_48_DFFSR_182 ( );
FILL FILL_49_DFFSR_182 ( );
FILL FILL_50_DFFSR_182 ( );
FILL FILL_51_DFFSR_182 ( );
FILL FILL_0_CLKBUF1_5 ( );
FILL FILL_1_CLKBUF1_5 ( );
FILL FILL_2_CLKBUF1_5 ( );
FILL FILL_3_CLKBUF1_5 ( );
FILL FILL_4_CLKBUF1_5 ( );
FILL FILL_5_CLKBUF1_5 ( );
FILL FILL_6_CLKBUF1_5 ( );
FILL FILL_7_CLKBUF1_5 ( );
FILL FILL_8_CLKBUF1_5 ( );
FILL FILL_9_CLKBUF1_5 ( );
FILL FILL_10_CLKBUF1_5 ( );
FILL FILL_11_CLKBUF1_5 ( );
FILL FILL_12_CLKBUF1_5 ( );
FILL FILL_13_CLKBUF1_5 ( );
FILL FILL_14_CLKBUF1_5 ( );
FILL FILL_15_CLKBUF1_5 ( );
FILL FILL_16_CLKBUF1_5 ( );
FILL FILL_17_CLKBUF1_5 ( );
FILL FILL_18_CLKBUF1_5 ( );
FILL FILL_19_CLKBUF1_5 ( );
FILL FILL_20_CLKBUF1_5 ( );
FILL FILL_0_NAND2X1_128 ( );
FILL FILL_1_NAND2X1_128 ( );
FILL FILL_2_NAND2X1_128 ( );
FILL FILL_3_NAND2X1_128 ( );
FILL FILL_4_NAND2X1_128 ( );
FILL FILL_5_NAND2X1_128 ( );
FILL FILL_6_NAND2X1_128 ( );
FILL FILL_0_INVX1_89 ( );
FILL FILL_1_INVX1_89 ( );
FILL FILL_2_INVX1_89 ( );
FILL FILL_3_INVX1_89 ( );
FILL FILL_4_INVX1_89 ( );
FILL FILL_0_INVX1_394 ( );
FILL FILL_1_INVX1_394 ( );
FILL FILL_2_INVX1_394 ( );
FILL FILL_3_INVX1_394 ( );
FILL FILL_4_INVX1_394 ( );
FILL FILL_0_INVX1_383 ( );
FILL FILL_1_INVX1_383 ( );
FILL FILL_2_INVX1_383 ( );
FILL FILL_3_INVX1_383 ( );
FILL FILL_0_OAI21X1_116 ( );
FILL FILL_1_OAI21X1_116 ( );
FILL FILL_2_OAI21X1_116 ( );
FILL FILL_3_OAI21X1_116 ( );
FILL FILL_4_OAI21X1_116 ( );
FILL FILL_5_OAI21X1_116 ( );
FILL FILL_6_OAI21X1_116 ( );
FILL FILL_7_OAI21X1_116 ( );
FILL FILL_8_OAI21X1_116 ( );
FILL FILL_0_DFFSR_108 ( );
FILL FILL_1_DFFSR_108 ( );
FILL FILL_2_DFFSR_108 ( );
FILL FILL_3_DFFSR_108 ( );
FILL FILL_4_DFFSR_108 ( );
FILL FILL_5_DFFSR_108 ( );
FILL FILL_6_DFFSR_108 ( );
FILL FILL_7_DFFSR_108 ( );
FILL FILL_8_DFFSR_108 ( );
FILL FILL_9_DFFSR_108 ( );
FILL FILL_10_DFFSR_108 ( );
FILL FILL_11_DFFSR_108 ( );
FILL FILL_12_DFFSR_108 ( );
FILL FILL_13_DFFSR_108 ( );
FILL FILL_14_DFFSR_108 ( );
FILL FILL_15_DFFSR_108 ( );
FILL FILL_16_DFFSR_108 ( );
FILL FILL_17_DFFSR_108 ( );
FILL FILL_18_DFFSR_108 ( );
FILL FILL_19_DFFSR_108 ( );
FILL FILL_20_DFFSR_108 ( );
FILL FILL_21_DFFSR_108 ( );
FILL FILL_22_DFFSR_108 ( );
FILL FILL_23_DFFSR_108 ( );
FILL FILL_24_DFFSR_108 ( );
FILL FILL_25_DFFSR_108 ( );
FILL FILL_26_DFFSR_108 ( );
FILL FILL_27_DFFSR_108 ( );
FILL FILL_28_DFFSR_108 ( );
FILL FILL_29_DFFSR_108 ( );
FILL FILL_30_DFFSR_108 ( );
FILL FILL_31_DFFSR_108 ( );
FILL FILL_32_DFFSR_108 ( );
FILL FILL_33_DFFSR_108 ( );
FILL FILL_34_DFFSR_108 ( );
FILL FILL_35_DFFSR_108 ( );
FILL FILL_36_DFFSR_108 ( );
FILL FILL_37_DFFSR_108 ( );
FILL FILL_38_DFFSR_108 ( );
FILL FILL_39_DFFSR_108 ( );
FILL FILL_40_DFFSR_108 ( );
FILL FILL_41_DFFSR_108 ( );
FILL FILL_42_DFFSR_108 ( );
FILL FILL_43_DFFSR_108 ( );
FILL FILL_44_DFFSR_108 ( );
FILL FILL_45_DFFSR_108 ( );
FILL FILL_46_DFFSR_108 ( );
FILL FILL_47_DFFSR_108 ( );
FILL FILL_48_DFFSR_108 ( );
FILL FILL_49_DFFSR_108 ( );
FILL FILL_50_DFFSR_108 ( );
FILL FILL_0_INVX1_349 ( );
FILL FILL_1_INVX1_349 ( );
FILL FILL_2_INVX1_349 ( );
FILL FILL_3_INVX1_349 ( );
FILL FILL_0_OAI22X1_45 ( );
FILL FILL_1_OAI22X1_45 ( );
FILL FILL_2_OAI22X1_45 ( );
FILL FILL_3_OAI22X1_45 ( );
FILL FILL_4_OAI22X1_45 ( );
FILL FILL_5_OAI22X1_45 ( );
FILL FILL_6_OAI22X1_45 ( );
FILL FILL_7_OAI22X1_45 ( );
FILL FILL_8_OAI22X1_45 ( );
FILL FILL_9_OAI22X1_45 ( );
FILL FILL_10_OAI22X1_45 ( );
FILL FILL_11_OAI22X1_45 ( );
FILL FILL_0_DFFSR_77 ( );
FILL FILL_1_DFFSR_77 ( );
FILL FILL_2_DFFSR_77 ( );
FILL FILL_3_DFFSR_77 ( );
FILL FILL_4_DFFSR_77 ( );
FILL FILL_5_DFFSR_77 ( );
FILL FILL_6_DFFSR_77 ( );
FILL FILL_7_DFFSR_77 ( );
FILL FILL_8_DFFSR_77 ( );
FILL FILL_9_DFFSR_77 ( );
FILL FILL_10_DFFSR_77 ( );
FILL FILL_11_DFFSR_77 ( );
FILL FILL_12_DFFSR_77 ( );
FILL FILL_13_DFFSR_77 ( );
FILL FILL_14_DFFSR_77 ( );
FILL FILL_15_DFFSR_77 ( );
FILL FILL_16_DFFSR_77 ( );
FILL FILL_17_DFFSR_77 ( );
FILL FILL_18_DFFSR_77 ( );
FILL FILL_19_DFFSR_77 ( );
FILL FILL_20_DFFSR_77 ( );
FILL FILL_21_DFFSR_77 ( );
FILL FILL_22_DFFSR_77 ( );
FILL FILL_23_DFFSR_77 ( );
FILL FILL_24_DFFSR_77 ( );
FILL FILL_25_DFFSR_77 ( );
FILL FILL_26_DFFSR_77 ( );
FILL FILL_27_DFFSR_77 ( );
FILL FILL_28_DFFSR_77 ( );
FILL FILL_29_DFFSR_77 ( );
FILL FILL_30_DFFSR_77 ( );
FILL FILL_31_DFFSR_77 ( );
FILL FILL_32_DFFSR_77 ( );
FILL FILL_33_DFFSR_77 ( );
FILL FILL_34_DFFSR_77 ( );
FILL FILL_35_DFFSR_77 ( );
FILL FILL_36_DFFSR_77 ( );
FILL FILL_37_DFFSR_77 ( );
FILL FILL_38_DFFSR_77 ( );
FILL FILL_39_DFFSR_77 ( );
FILL FILL_40_DFFSR_77 ( );
FILL FILL_41_DFFSR_77 ( );
FILL FILL_42_DFFSR_77 ( );
FILL FILL_43_DFFSR_77 ( );
FILL FILL_44_DFFSR_77 ( );
FILL FILL_45_DFFSR_77 ( );
FILL FILL_46_DFFSR_77 ( );
FILL FILL_47_DFFSR_77 ( );
FILL FILL_48_DFFSR_77 ( );
FILL FILL_49_DFFSR_77 ( );
FILL FILL_50_DFFSR_77 ( );
FILL FILL_51_DFFSR_77 ( );
FILL FILL_0_INVX1_429 ( );
FILL FILL_1_INVX1_429 ( );
FILL FILL_2_INVX1_429 ( );
FILL FILL_3_INVX1_429 ( );
FILL FILL_4_INVX1_429 ( );
FILL FILL_0_NAND2X1_271 ( );
FILL FILL_1_NAND2X1_271 ( );
FILL FILL_2_NAND2X1_271 ( );
FILL FILL_3_NAND2X1_271 ( );
FILL FILL_4_NAND2X1_271 ( );
FILL FILL_5_NAND2X1_271 ( );
FILL FILL_6_NAND2X1_271 ( );
FILL FILL_0_INVX1_18 ( );
FILL FILL_1_INVX1_18 ( );
FILL FILL_2_INVX1_18 ( );
FILL FILL_3_INVX1_18 ( );
FILL FILL_0_NAND2X1_282 ( );
FILL FILL_1_NAND2X1_282 ( );
FILL FILL_2_NAND2X1_282 ( );
FILL FILL_3_NAND2X1_282 ( );
FILL FILL_4_NAND2X1_282 ( );
FILL FILL_5_NAND2X1_282 ( );
FILL FILL_6_NAND2X1_282 ( );
FILL FILL_0_NOR3X1_2 ( );
FILL FILL_1_NOR3X1_2 ( );
FILL FILL_2_NOR3X1_2 ( );
FILL FILL_3_NOR3X1_2 ( );
FILL FILL_4_NOR3X1_2 ( );
FILL FILL_5_NOR3X1_2 ( );
FILL FILL_6_NOR3X1_2 ( );
FILL FILL_7_NOR3X1_2 ( );
FILL FILL_8_NOR3X1_2 ( );
FILL FILL_9_NOR3X1_2 ( );
FILL FILL_10_NOR3X1_2 ( );
FILL FILL_11_NOR3X1_2 ( );
FILL FILL_12_NOR3X1_2 ( );
FILL FILL_13_NOR3X1_2 ( );
FILL FILL_14_NOR3X1_2 ( );
FILL FILL_15_NOR3X1_2 ( );
FILL FILL_16_NOR3X1_2 ( );
FILL FILL_17_NOR3X1_2 ( );
FILL FILL_18_NOR3X1_2 ( );
FILL FILL_0_NAND2X1_279 ( );
FILL FILL_1_NAND2X1_279 ( );
FILL FILL_2_NAND2X1_279 ( );
FILL FILL_3_NAND2X1_279 ( );
FILL FILL_4_NAND2X1_279 ( );
FILL FILL_5_NAND2X1_279 ( );
FILL FILL_6_NAND2X1_279 ( );
FILL FILL_0_XOR2X1_14 ( );
FILL FILL_1_XOR2X1_14 ( );
FILL FILL_2_XOR2X1_14 ( );
FILL FILL_3_XOR2X1_14 ( );
FILL FILL_4_XOR2X1_14 ( );
FILL FILL_5_XOR2X1_14 ( );
FILL FILL_6_XOR2X1_14 ( );
FILL FILL_7_XOR2X1_14 ( );
FILL FILL_8_XOR2X1_14 ( );
FILL FILL_9_XOR2X1_14 ( );
FILL FILL_10_XOR2X1_14 ( );
FILL FILL_11_XOR2X1_14 ( );
FILL FILL_12_XOR2X1_14 ( );
FILL FILL_13_XOR2X1_14 ( );
FILL FILL_14_XOR2X1_14 ( );
FILL FILL_15_XOR2X1_14 ( );
FILL FILL_16_XOR2X1_14 ( );
FILL FILL_0_INVX1_320 ( );
FILL FILL_1_INVX1_320 ( );
FILL FILL_2_INVX1_320 ( );
FILL FILL_3_INVX1_320 ( );
FILL FILL_4_INVX1_320 ( );
FILL FILL_0_INVX1_62 ( );
FILL FILL_1_INVX1_62 ( );
FILL FILL_2_INVX1_62 ( );
FILL FILL_3_INVX1_62 ( );
FILL FILL_4_INVX1_62 ( );
FILL FILL_0_OAI21X1_55 ( );
FILL FILL_1_OAI21X1_55 ( );
FILL FILL_2_OAI21X1_55 ( );
FILL FILL_3_OAI21X1_55 ( );
FILL FILL_4_OAI21X1_55 ( );
FILL FILL_5_OAI21X1_55 ( );
FILL FILL_6_OAI21X1_55 ( );
FILL FILL_7_OAI21X1_55 ( );
FILL FILL_8_OAI21X1_55 ( );
FILL FILL_0_NAND2X1_55 ( );
FILL FILL_1_NAND2X1_55 ( );
FILL FILL_2_NAND2X1_55 ( );
FILL FILL_3_NAND2X1_55 ( );
FILL FILL_4_NAND2X1_55 ( );
FILL FILL_5_NAND2X1_55 ( );
FILL FILL_6_NAND2X1_55 ( );
FILL FILL_0_OAI21X1_47 ( );
FILL FILL_1_OAI21X1_47 ( );
FILL FILL_2_OAI21X1_47 ( );
FILL FILL_3_OAI21X1_47 ( );
FILL FILL_4_OAI21X1_47 ( );
FILL FILL_5_OAI21X1_47 ( );
FILL FILL_6_OAI21X1_47 ( );
FILL FILL_7_OAI21X1_47 ( );
FILL FILL_8_OAI21X1_47 ( );
FILL FILL_0_INVX1_53 ( );
FILL FILL_1_INVX1_53 ( );
FILL FILL_2_INVX1_53 ( );
FILL FILL_3_INVX1_53 ( );
FILL FILL_4_INVX1_53 ( );
FILL FILL_0_NAND2X1_43 ( );
FILL FILL_1_NAND2X1_43 ( );
FILL FILL_2_NAND2X1_43 ( );
FILL FILL_3_NAND2X1_43 ( );
FILL FILL_4_NAND2X1_43 ( );
FILL FILL_5_NAND2X1_43 ( );
FILL FILL_6_NAND2X1_43 ( );
FILL FILL_0_OAI22X1_23 ( );
FILL FILL_1_OAI22X1_23 ( );
FILL FILL_2_OAI22X1_23 ( );
FILL FILL_3_OAI22X1_23 ( );
FILL FILL_4_OAI22X1_23 ( );
FILL FILL_5_OAI22X1_23 ( );
FILL FILL_6_OAI22X1_23 ( );
FILL FILL_7_OAI22X1_23 ( );
FILL FILL_8_OAI22X1_23 ( );
FILL FILL_9_OAI22X1_23 ( );
FILL FILL_10_OAI22X1_23 ( );
FILL FILL_0_INVX1_301 ( );
FILL FILL_1_INVX1_301 ( );
FILL FILL_2_INVX1_301 ( );
FILL FILL_3_INVX1_301 ( );
FILL FILL_4_INVX1_301 ( );
FILL FILL_0_DFFSR_37 ( );
FILL FILL_1_DFFSR_37 ( );
FILL FILL_2_DFFSR_37 ( );
FILL FILL_3_DFFSR_37 ( );
FILL FILL_4_DFFSR_37 ( );
FILL FILL_5_DFFSR_37 ( );
FILL FILL_6_DFFSR_37 ( );
FILL FILL_7_DFFSR_37 ( );
FILL FILL_8_DFFSR_37 ( );
FILL FILL_9_DFFSR_37 ( );
FILL FILL_10_DFFSR_37 ( );
FILL FILL_11_DFFSR_37 ( );
FILL FILL_12_DFFSR_37 ( );
FILL FILL_13_DFFSR_37 ( );
FILL FILL_14_DFFSR_37 ( );
FILL FILL_15_DFFSR_37 ( );
FILL FILL_16_DFFSR_37 ( );
FILL FILL_17_DFFSR_37 ( );
FILL FILL_18_DFFSR_37 ( );
FILL FILL_19_DFFSR_37 ( );
FILL FILL_20_DFFSR_37 ( );
FILL FILL_21_DFFSR_37 ( );
FILL FILL_22_DFFSR_37 ( );
FILL FILL_23_DFFSR_37 ( );
FILL FILL_24_DFFSR_37 ( );
FILL FILL_25_DFFSR_37 ( );
FILL FILL_26_DFFSR_37 ( );
FILL FILL_27_DFFSR_37 ( );
FILL FILL_28_DFFSR_37 ( );
FILL FILL_29_DFFSR_37 ( );
FILL FILL_30_DFFSR_37 ( );
FILL FILL_31_DFFSR_37 ( );
FILL FILL_32_DFFSR_37 ( );
FILL FILL_33_DFFSR_37 ( );
FILL FILL_34_DFFSR_37 ( );
FILL FILL_35_DFFSR_37 ( );
FILL FILL_36_DFFSR_37 ( );
FILL FILL_37_DFFSR_37 ( );
FILL FILL_38_DFFSR_37 ( );
FILL FILL_39_DFFSR_37 ( );
FILL FILL_40_DFFSR_37 ( );
FILL FILL_41_DFFSR_37 ( );
FILL FILL_42_DFFSR_37 ( );
FILL FILL_43_DFFSR_37 ( );
FILL FILL_44_DFFSR_37 ( );
FILL FILL_45_DFFSR_37 ( );
FILL FILL_46_DFFSR_37 ( );
FILL FILL_47_DFFSR_37 ( );
FILL FILL_48_DFFSR_37 ( );
FILL FILL_49_DFFSR_37 ( );
FILL FILL_50_DFFSR_37 ( );
FILL FILL_0_OAI21X1_37 ( );
FILL FILL_1_OAI21X1_37 ( );
FILL FILL_2_OAI21X1_37 ( );
FILL FILL_3_OAI21X1_37 ( );
FILL FILL_4_OAI21X1_37 ( );
FILL FILL_5_OAI21X1_37 ( );
FILL FILL_6_OAI21X1_37 ( );
FILL FILL_7_OAI21X1_37 ( );
FILL FILL_8_OAI21X1_37 ( );
FILL FILL_9_OAI21X1_37 ( );
FILL FILL_0_CLKBUF1_23 ( );
FILL FILL_1_CLKBUF1_23 ( );
FILL FILL_2_CLKBUF1_23 ( );
FILL FILL_3_CLKBUF1_23 ( );
FILL FILL_4_CLKBUF1_23 ( );
FILL FILL_5_CLKBUF1_23 ( );
FILL FILL_6_CLKBUF1_23 ( );
FILL FILL_7_CLKBUF1_23 ( );
FILL FILL_8_CLKBUF1_23 ( );
FILL FILL_9_CLKBUF1_23 ( );
FILL FILL_10_CLKBUF1_23 ( );
FILL FILL_11_CLKBUF1_23 ( );
FILL FILL_12_CLKBUF1_23 ( );
FILL FILL_13_CLKBUF1_23 ( );
FILL FILL_14_CLKBUF1_23 ( );
FILL FILL_15_CLKBUF1_23 ( );
FILL FILL_16_CLKBUF1_23 ( );
FILL FILL_17_CLKBUF1_23 ( );
FILL FILL_18_CLKBUF1_23 ( );
FILL FILL_19_CLKBUF1_23 ( );
FILL FILL_20_CLKBUF1_23 ( );
FILL FILL_0_OAI21X1_188 ( );
FILL FILL_1_OAI21X1_188 ( );
FILL FILL_2_OAI21X1_188 ( );
FILL FILL_3_OAI21X1_188 ( );
FILL FILL_4_OAI21X1_188 ( );
FILL FILL_5_OAI21X1_188 ( );
FILL FILL_6_OAI21X1_188 ( );
FILL FILL_7_OAI21X1_188 ( );
FILL FILL_8_OAI21X1_188 ( );
FILL FILL_9_OAI21X1_188 ( );
FILL FILL_0_DFFSR_164 ( );
FILL FILL_1_DFFSR_164 ( );
FILL FILL_2_DFFSR_164 ( );
FILL FILL_3_DFFSR_164 ( );
FILL FILL_4_DFFSR_164 ( );
FILL FILL_5_DFFSR_164 ( );
FILL FILL_6_DFFSR_164 ( );
FILL FILL_7_DFFSR_164 ( );
FILL FILL_8_DFFSR_164 ( );
FILL FILL_9_DFFSR_164 ( );
FILL FILL_10_DFFSR_164 ( );
FILL FILL_11_DFFSR_164 ( );
FILL FILL_12_DFFSR_164 ( );
FILL FILL_13_DFFSR_164 ( );
FILL FILL_14_DFFSR_164 ( );
FILL FILL_15_DFFSR_164 ( );
FILL FILL_16_DFFSR_164 ( );
FILL FILL_17_DFFSR_164 ( );
FILL FILL_18_DFFSR_164 ( );
FILL FILL_19_DFFSR_164 ( );
FILL FILL_20_DFFSR_164 ( );
FILL FILL_21_DFFSR_164 ( );
FILL FILL_22_DFFSR_164 ( );
FILL FILL_23_DFFSR_164 ( );
FILL FILL_24_DFFSR_164 ( );
FILL FILL_25_DFFSR_164 ( );
FILL FILL_26_DFFSR_164 ( );
FILL FILL_27_DFFSR_164 ( );
FILL FILL_28_DFFSR_164 ( );
FILL FILL_29_DFFSR_164 ( );
FILL FILL_30_DFFSR_164 ( );
FILL FILL_31_DFFSR_164 ( );
FILL FILL_32_DFFSR_164 ( );
FILL FILL_33_DFFSR_164 ( );
FILL FILL_34_DFFSR_164 ( );
FILL FILL_35_DFFSR_164 ( );
FILL FILL_36_DFFSR_164 ( );
FILL FILL_37_DFFSR_164 ( );
FILL FILL_38_DFFSR_164 ( );
FILL FILL_39_DFFSR_164 ( );
FILL FILL_40_DFFSR_164 ( );
FILL FILL_41_DFFSR_164 ( );
FILL FILL_42_DFFSR_164 ( );
FILL FILL_43_DFFSR_164 ( );
FILL FILL_44_DFFSR_164 ( );
FILL FILL_45_DFFSR_164 ( );
FILL FILL_46_DFFSR_164 ( );
FILL FILL_47_DFFSR_164 ( );
FILL FILL_48_DFFSR_164 ( );
FILL FILL_49_DFFSR_164 ( );
FILL FILL_50_DFFSR_164 ( );
FILL FILL_51_DFFSR_164 ( );
FILL FILL_0_BUFX2_22 ( );
FILL FILL_1_BUFX2_22 ( );
FILL FILL_2_BUFX2_22 ( );
FILL FILL_3_BUFX2_22 ( );
FILL FILL_4_BUFX2_22 ( );
FILL FILL_5_BUFX2_22 ( );
FILL FILL_6_BUFX2_22 ( );
FILL FILL_0_NAND2X1_103 ( );
FILL FILL_1_NAND2X1_103 ( );
FILL FILL_2_NAND2X1_103 ( );
FILL FILL_3_NAND2X1_103 ( );
FILL FILL_4_NAND2X1_103 ( );
FILL FILL_5_NAND2X1_103 ( );
FILL FILL_6_NAND2X1_103 ( );
FILL FILL_0_NAND2X1_87 ( );
FILL FILL_1_NAND2X1_87 ( );
FILL FILL_2_NAND2X1_87 ( );
FILL FILL_3_NAND2X1_87 ( );
FILL FILL_4_NAND2X1_87 ( );
FILL FILL_5_NAND2X1_87 ( );
FILL FILL_6_NAND2X1_87 ( );
FILL FILL_0_DFFSR_116 ( );
FILL FILL_1_DFFSR_116 ( );
FILL FILL_2_DFFSR_116 ( );
FILL FILL_3_DFFSR_116 ( );
FILL FILL_4_DFFSR_116 ( );
FILL FILL_5_DFFSR_116 ( );
FILL FILL_6_DFFSR_116 ( );
FILL FILL_7_DFFSR_116 ( );
FILL FILL_8_DFFSR_116 ( );
FILL FILL_9_DFFSR_116 ( );
FILL FILL_10_DFFSR_116 ( );
FILL FILL_11_DFFSR_116 ( );
FILL FILL_12_DFFSR_116 ( );
FILL FILL_13_DFFSR_116 ( );
FILL FILL_14_DFFSR_116 ( );
FILL FILL_15_DFFSR_116 ( );
FILL FILL_16_DFFSR_116 ( );
FILL FILL_17_DFFSR_116 ( );
FILL FILL_18_DFFSR_116 ( );
FILL FILL_19_DFFSR_116 ( );
FILL FILL_20_DFFSR_116 ( );
FILL FILL_21_DFFSR_116 ( );
FILL FILL_22_DFFSR_116 ( );
FILL FILL_23_DFFSR_116 ( );
FILL FILL_24_DFFSR_116 ( );
FILL FILL_25_DFFSR_116 ( );
FILL FILL_26_DFFSR_116 ( );
FILL FILL_27_DFFSR_116 ( );
FILL FILL_28_DFFSR_116 ( );
FILL FILL_29_DFFSR_116 ( );
FILL FILL_30_DFFSR_116 ( );
FILL FILL_31_DFFSR_116 ( );
FILL FILL_32_DFFSR_116 ( );
FILL FILL_33_DFFSR_116 ( );
FILL FILL_34_DFFSR_116 ( );
FILL FILL_35_DFFSR_116 ( );
FILL FILL_36_DFFSR_116 ( );
FILL FILL_37_DFFSR_116 ( );
FILL FILL_38_DFFSR_116 ( );
FILL FILL_39_DFFSR_116 ( );
FILL FILL_40_DFFSR_116 ( );
FILL FILL_41_DFFSR_116 ( );
FILL FILL_42_DFFSR_116 ( );
FILL FILL_43_DFFSR_116 ( );
FILL FILL_44_DFFSR_116 ( );
FILL FILL_45_DFFSR_116 ( );
FILL FILL_46_DFFSR_116 ( );
FILL FILL_47_DFFSR_116 ( );
FILL FILL_48_DFFSR_116 ( );
FILL FILL_49_DFFSR_116 ( );
FILL FILL_50_DFFSR_116 ( );
FILL FILL_0_INVX1_369 ( );
FILL FILL_1_INVX1_369 ( );
FILL FILL_2_INVX1_369 ( );
FILL FILL_3_INVX1_369 ( );
FILL FILL_0_NAND3X1_123 ( );
FILL FILL_1_NAND3X1_123 ( );
FILL FILL_2_NAND3X1_123 ( );
FILL FILL_3_NAND3X1_123 ( );
FILL FILL_4_NAND3X1_123 ( );
FILL FILL_5_NAND3X1_123 ( );
FILL FILL_6_NAND3X1_123 ( );
FILL FILL_7_NAND3X1_123 ( );
FILL FILL_8_NAND3X1_123 ( );
FILL FILL_0_INVX1_332 ( );
FILL FILL_1_INVX1_332 ( );
FILL FILL_2_INVX1_332 ( );
FILL FILL_3_INVX1_332 ( );
FILL FILL_4_INVX1_332 ( );
FILL FILL_0_INVX1_333 ( );
FILL FILL_1_INVX1_333 ( );
FILL FILL_2_INVX1_333 ( );
FILL FILL_3_INVX1_333 ( );
FILL FILL_4_INVX1_333 ( );
FILL FILL_0_NAND3X1_119 ( );
FILL FILL_1_NAND3X1_119 ( );
FILL FILL_2_NAND3X1_119 ( );
FILL FILL_3_NAND3X1_119 ( );
FILL FILL_4_NAND3X1_119 ( );
FILL FILL_5_NAND3X1_119 ( );
FILL FILL_6_NAND3X1_119 ( );
FILL FILL_7_NAND3X1_119 ( );
FILL FILL_8_NAND3X1_119 ( );
FILL FILL_0_INVX1_331 ( );
FILL FILL_1_INVX1_331 ( );
FILL FILL_2_INVX1_331 ( );
FILL FILL_3_INVX1_331 ( );
FILL FILL_0_INVX1_399 ( );
FILL FILL_1_INVX1_399 ( );
FILL FILL_2_INVX1_399 ( );
FILL FILL_3_INVX1_399 ( );
FILL FILL_4_INVX1_399 ( );
FILL FILL_0_NAND3X1_127 ( );
FILL FILL_1_NAND3X1_127 ( );
FILL FILL_2_NAND3X1_127 ( );
FILL FILL_3_NAND3X1_127 ( );
FILL FILL_4_NAND3X1_127 ( );
FILL FILL_5_NAND3X1_127 ( );
FILL FILL_6_NAND3X1_127 ( );
FILL FILL_7_NAND3X1_127 ( );
FILL FILL_8_NAND3X1_127 ( );
FILL FILL_0_INVX1_398 ( );
FILL FILL_1_INVX1_398 ( );
FILL FILL_2_INVX1_398 ( );
FILL FILL_3_INVX1_398 ( );
FILL FILL_4_INVX1_398 ( );
FILL FILL_0_INVX1_81 ( );
FILL FILL_1_INVX1_81 ( );
FILL FILL_2_INVX1_81 ( );
FILL FILL_3_INVX1_81 ( );
FILL FILL_4_INVX1_81 ( );
FILL FILL_0_OAI21X1_72 ( );
FILL FILL_1_OAI21X1_72 ( );
FILL FILL_2_OAI21X1_72 ( );
FILL FILL_3_OAI21X1_72 ( );
FILL FILL_4_OAI21X1_72 ( );
FILL FILL_5_OAI21X1_72 ( );
FILL FILL_6_OAI21X1_72 ( );
FILL FILL_7_OAI21X1_72 ( );
FILL FILL_8_OAI21X1_72 ( );
FILL FILL_0_NAND2X1_70 ( );
FILL FILL_1_NAND2X1_70 ( );
FILL FILL_2_NAND2X1_70 ( );
FILL FILL_3_NAND2X1_70 ( );
FILL FILL_4_NAND2X1_70 ( );
FILL FILL_5_NAND2X1_70 ( );
FILL FILL_6_NAND2X1_70 ( );
FILL FILL_0_NAND2X1_72 ( );
FILL FILL_1_NAND2X1_72 ( );
FILL FILL_2_NAND2X1_72 ( );
FILL FILL_3_NAND2X1_72 ( );
FILL FILL_4_NAND2X1_72 ( );
FILL FILL_5_NAND2X1_72 ( );
FILL FILL_6_NAND2X1_72 ( );
FILL FILL_0_NAND2X1_136 ( );
FILL FILL_1_NAND2X1_136 ( );
FILL FILL_2_NAND2X1_136 ( );
FILL FILL_3_NAND2X1_136 ( );
FILL FILL_4_NAND2X1_136 ( );
FILL FILL_5_NAND2X1_136 ( );
FILL FILL_6_NAND2X1_136 ( );
FILL FILL_0_OAI21X1_136 ( );
FILL FILL_1_OAI21X1_136 ( );
FILL FILL_2_OAI21X1_136 ( );
FILL FILL_3_OAI21X1_136 ( );
FILL FILL_4_OAI21X1_136 ( );
FILL FILL_5_OAI21X1_136 ( );
FILL FILL_6_OAI21X1_136 ( );
FILL FILL_7_OAI21X1_136 ( );
FILL FILL_8_OAI21X1_136 ( );
FILL FILL_9_OAI21X1_136 ( );
FILL FILL_0_INVX1_153 ( );
FILL FILL_1_INVX1_153 ( );
FILL FILL_2_INVX1_153 ( );
FILL FILL_3_INVX1_153 ( );
FILL FILL_0_DFFSR_40 ( );
FILL FILL_1_DFFSR_40 ( );
FILL FILL_2_DFFSR_40 ( );
FILL FILL_3_DFFSR_40 ( );
FILL FILL_4_DFFSR_40 ( );
FILL FILL_5_DFFSR_40 ( );
FILL FILL_6_DFFSR_40 ( );
FILL FILL_7_DFFSR_40 ( );
FILL FILL_8_DFFSR_40 ( );
FILL FILL_9_DFFSR_40 ( );
FILL FILL_10_DFFSR_40 ( );
FILL FILL_11_DFFSR_40 ( );
FILL FILL_12_DFFSR_40 ( );
FILL FILL_13_DFFSR_40 ( );
FILL FILL_14_DFFSR_40 ( );
FILL FILL_15_DFFSR_40 ( );
FILL FILL_16_DFFSR_40 ( );
FILL FILL_17_DFFSR_40 ( );
FILL FILL_18_DFFSR_40 ( );
FILL FILL_19_DFFSR_40 ( );
FILL FILL_20_DFFSR_40 ( );
FILL FILL_21_DFFSR_40 ( );
FILL FILL_22_DFFSR_40 ( );
FILL FILL_23_DFFSR_40 ( );
FILL FILL_24_DFFSR_40 ( );
FILL FILL_25_DFFSR_40 ( );
FILL FILL_26_DFFSR_40 ( );
FILL FILL_27_DFFSR_40 ( );
FILL FILL_28_DFFSR_40 ( );
FILL FILL_29_DFFSR_40 ( );
FILL FILL_30_DFFSR_40 ( );
FILL FILL_31_DFFSR_40 ( );
FILL FILL_32_DFFSR_40 ( );
FILL FILL_33_DFFSR_40 ( );
FILL FILL_34_DFFSR_40 ( );
FILL FILL_35_DFFSR_40 ( );
FILL FILL_36_DFFSR_40 ( );
FILL FILL_37_DFFSR_40 ( );
FILL FILL_38_DFFSR_40 ( );
FILL FILL_39_DFFSR_40 ( );
FILL FILL_40_DFFSR_40 ( );
FILL FILL_41_DFFSR_40 ( );
FILL FILL_42_DFFSR_40 ( );
FILL FILL_43_DFFSR_40 ( );
FILL FILL_44_DFFSR_40 ( );
FILL FILL_45_DFFSR_40 ( );
FILL FILL_46_DFFSR_40 ( );
FILL FILL_47_DFFSR_40 ( );
FILL FILL_48_DFFSR_40 ( );
FILL FILL_49_DFFSR_40 ( );
FILL FILL_50_DFFSR_40 ( );
FILL FILL_0_DFFSR_47 ( );
FILL FILL_1_DFFSR_47 ( );
FILL FILL_2_DFFSR_47 ( );
FILL FILL_3_DFFSR_47 ( );
FILL FILL_4_DFFSR_47 ( );
FILL FILL_5_DFFSR_47 ( );
FILL FILL_6_DFFSR_47 ( );
FILL FILL_7_DFFSR_47 ( );
FILL FILL_8_DFFSR_47 ( );
FILL FILL_9_DFFSR_47 ( );
FILL FILL_10_DFFSR_47 ( );
FILL FILL_11_DFFSR_47 ( );
FILL FILL_12_DFFSR_47 ( );
FILL FILL_13_DFFSR_47 ( );
FILL FILL_14_DFFSR_47 ( );
FILL FILL_15_DFFSR_47 ( );
FILL FILL_16_DFFSR_47 ( );
FILL FILL_17_DFFSR_47 ( );
FILL FILL_18_DFFSR_47 ( );
FILL FILL_19_DFFSR_47 ( );
FILL FILL_20_DFFSR_47 ( );
FILL FILL_21_DFFSR_47 ( );
FILL FILL_22_DFFSR_47 ( );
FILL FILL_23_DFFSR_47 ( );
FILL FILL_24_DFFSR_47 ( );
FILL FILL_25_DFFSR_47 ( );
FILL FILL_26_DFFSR_47 ( );
FILL FILL_27_DFFSR_47 ( );
FILL FILL_28_DFFSR_47 ( );
FILL FILL_29_DFFSR_47 ( );
FILL FILL_30_DFFSR_47 ( );
FILL FILL_31_DFFSR_47 ( );
FILL FILL_32_DFFSR_47 ( );
FILL FILL_33_DFFSR_47 ( );
FILL FILL_34_DFFSR_47 ( );
FILL FILL_35_DFFSR_47 ( );
FILL FILL_36_DFFSR_47 ( );
FILL FILL_37_DFFSR_47 ( );
FILL FILL_38_DFFSR_47 ( );
FILL FILL_39_DFFSR_47 ( );
FILL FILL_40_DFFSR_47 ( );
FILL FILL_41_DFFSR_47 ( );
FILL FILL_42_DFFSR_47 ( );
FILL FILL_43_DFFSR_47 ( );
FILL FILL_44_DFFSR_47 ( );
FILL FILL_45_DFFSR_47 ( );
FILL FILL_46_DFFSR_47 ( );
FILL FILL_47_DFFSR_47 ( );
FILL FILL_48_DFFSR_47 ( );
FILL FILL_49_DFFSR_47 ( );
FILL FILL_50_DFFSR_47 ( );
FILL FILL_0_DFFSR_35 ( );
FILL FILL_1_DFFSR_35 ( );
FILL FILL_2_DFFSR_35 ( );
FILL FILL_3_DFFSR_35 ( );
FILL FILL_4_DFFSR_35 ( );
FILL FILL_5_DFFSR_35 ( );
FILL FILL_6_DFFSR_35 ( );
FILL FILL_7_DFFSR_35 ( );
FILL FILL_8_DFFSR_35 ( );
FILL FILL_9_DFFSR_35 ( );
FILL FILL_10_DFFSR_35 ( );
FILL FILL_11_DFFSR_35 ( );
FILL FILL_12_DFFSR_35 ( );
FILL FILL_13_DFFSR_35 ( );
FILL FILL_14_DFFSR_35 ( );
FILL FILL_15_DFFSR_35 ( );
FILL FILL_16_DFFSR_35 ( );
FILL FILL_17_DFFSR_35 ( );
FILL FILL_18_DFFSR_35 ( );
FILL FILL_19_DFFSR_35 ( );
FILL FILL_20_DFFSR_35 ( );
FILL FILL_21_DFFSR_35 ( );
FILL FILL_22_DFFSR_35 ( );
FILL FILL_23_DFFSR_35 ( );
FILL FILL_24_DFFSR_35 ( );
FILL FILL_25_DFFSR_35 ( );
FILL FILL_26_DFFSR_35 ( );
FILL FILL_27_DFFSR_35 ( );
FILL FILL_28_DFFSR_35 ( );
FILL FILL_29_DFFSR_35 ( );
FILL FILL_30_DFFSR_35 ( );
FILL FILL_31_DFFSR_35 ( );
FILL FILL_32_DFFSR_35 ( );
FILL FILL_33_DFFSR_35 ( );
FILL FILL_34_DFFSR_35 ( );
FILL FILL_35_DFFSR_35 ( );
FILL FILL_36_DFFSR_35 ( );
FILL FILL_37_DFFSR_35 ( );
FILL FILL_38_DFFSR_35 ( );
FILL FILL_39_DFFSR_35 ( );
FILL FILL_40_DFFSR_35 ( );
FILL FILL_41_DFFSR_35 ( );
FILL FILL_42_DFFSR_35 ( );
FILL FILL_43_DFFSR_35 ( );
FILL FILL_44_DFFSR_35 ( );
FILL FILL_45_DFFSR_35 ( );
FILL FILL_46_DFFSR_35 ( );
FILL FILL_47_DFFSR_35 ( );
FILL FILL_48_DFFSR_35 ( );
FILL FILL_49_DFFSR_35 ( );
FILL FILL_50_DFFSR_35 ( );
FILL FILL_0_DFFSR_2 ( );
FILL FILL_1_DFFSR_2 ( );
FILL FILL_2_DFFSR_2 ( );
FILL FILL_3_DFFSR_2 ( );
FILL FILL_4_DFFSR_2 ( );
FILL FILL_5_DFFSR_2 ( );
FILL FILL_6_DFFSR_2 ( );
FILL FILL_7_DFFSR_2 ( );
FILL FILL_8_DFFSR_2 ( );
FILL FILL_9_DFFSR_2 ( );
FILL FILL_10_DFFSR_2 ( );
FILL FILL_11_DFFSR_2 ( );
FILL FILL_12_DFFSR_2 ( );
FILL FILL_13_DFFSR_2 ( );
FILL FILL_14_DFFSR_2 ( );
FILL FILL_15_DFFSR_2 ( );
FILL FILL_16_DFFSR_2 ( );
FILL FILL_17_DFFSR_2 ( );
FILL FILL_18_DFFSR_2 ( );
FILL FILL_19_DFFSR_2 ( );
FILL FILL_20_DFFSR_2 ( );
FILL FILL_21_DFFSR_2 ( );
FILL FILL_22_DFFSR_2 ( );
FILL FILL_23_DFFSR_2 ( );
FILL FILL_24_DFFSR_2 ( );
FILL FILL_25_DFFSR_2 ( );
FILL FILL_26_DFFSR_2 ( );
FILL FILL_27_DFFSR_2 ( );
FILL FILL_28_DFFSR_2 ( );
FILL FILL_29_DFFSR_2 ( );
FILL FILL_30_DFFSR_2 ( );
FILL FILL_31_DFFSR_2 ( );
FILL FILL_32_DFFSR_2 ( );
FILL FILL_33_DFFSR_2 ( );
FILL FILL_34_DFFSR_2 ( );
FILL FILL_35_DFFSR_2 ( );
FILL FILL_36_DFFSR_2 ( );
FILL FILL_37_DFFSR_2 ( );
FILL FILL_38_DFFSR_2 ( );
FILL FILL_39_DFFSR_2 ( );
FILL FILL_40_DFFSR_2 ( );
FILL FILL_41_DFFSR_2 ( );
FILL FILL_42_DFFSR_2 ( );
FILL FILL_43_DFFSR_2 ( );
FILL FILL_44_DFFSR_2 ( );
FILL FILL_45_DFFSR_2 ( );
FILL FILL_46_DFFSR_2 ( );
FILL FILL_47_DFFSR_2 ( );
FILL FILL_48_DFFSR_2 ( );
FILL FILL_49_DFFSR_2 ( );
FILL FILL_50_DFFSR_2 ( );
FILL FILL_0_BUFX2_1 ( );
FILL FILL_1_BUFX2_1 ( );
FILL FILL_2_BUFX2_1 ( );
FILL FILL_3_BUFX2_1 ( );
FILL FILL_4_BUFX2_1 ( );
FILL FILL_5_BUFX2_1 ( );
FILL FILL_6_BUFX2_1 ( );
FILL FILL_0_INVX1_229 ( );
FILL FILL_1_INVX1_229 ( );
FILL FILL_2_INVX1_229 ( );
FILL FILL_3_INVX1_229 ( );
FILL FILL_4_INVX1_229 ( );
FILL FILL_0_BUFX2_3 ( );
FILL FILL_1_BUFX2_3 ( );
FILL FILL_2_BUFX2_3 ( );
FILL FILL_3_BUFX2_3 ( );
FILL FILL_4_BUFX2_3 ( );
FILL FILL_5_BUFX2_3 ( );
FILL FILL_6_BUFX2_3 ( );
FILL FILL_0_INVX1_212 ( );
FILL FILL_1_INVX1_212 ( );
FILL FILL_2_INVX1_212 ( );
FILL FILL_3_INVX1_212 ( );
FILL FILL_4_INVX1_212 ( );
FILL FILL_0_INVX1_228 ( );
FILL FILL_1_INVX1_228 ( );
FILL FILL_2_INVX1_228 ( );
FILL FILL_3_INVX1_228 ( );
FILL FILL_0_INVX1_407 ( );
FILL FILL_1_INVX1_407 ( );
FILL FILL_2_INVX1_407 ( );
FILL FILL_3_INVX1_407 ( );
FILL FILL_0_OAI21X1_164 ( );
FILL FILL_1_OAI21X1_164 ( );
FILL FILL_2_OAI21X1_164 ( );
FILL FILL_3_OAI21X1_164 ( );
FILL FILL_4_OAI21X1_164 ( );
FILL FILL_5_OAI21X1_164 ( );
FILL FILL_6_OAI21X1_164 ( );
FILL FILL_7_OAI21X1_164 ( );
FILL FILL_8_OAI21X1_164 ( );
FILL FILL_0_INVX1_198 ( );
FILL FILL_1_INVX1_198 ( );
FILL FILL_2_INVX1_198 ( );
FILL FILL_3_INVX1_198 ( );
FILL FILL_4_INVX1_198 ( );
FILL FILL_0_OAI21X1_245 ( );
FILL FILL_1_OAI21X1_245 ( );
FILL FILL_2_OAI21X1_245 ( );
FILL FILL_3_OAI21X1_245 ( );
FILL FILL_4_OAI21X1_245 ( );
FILL FILL_5_OAI21X1_245 ( );
FILL FILL_6_OAI21X1_245 ( );
FILL FILL_7_OAI21X1_245 ( );
FILL FILL_8_OAI21X1_245 ( );
FILL FILL_9_OAI21X1_245 ( );
FILL FILL_0_NAND2X1_256 ( );
FILL FILL_1_NAND2X1_256 ( );
FILL FILL_2_NAND2X1_256 ( );
FILL FILL_3_NAND2X1_256 ( );
FILL FILL_4_NAND2X1_256 ( );
FILL FILL_5_NAND2X1_256 ( );
FILL FILL_6_NAND2X1_256 ( );
FILL FILL_0_OAI21X1_103 ( );
FILL FILL_1_OAI21X1_103 ( );
FILL FILL_2_OAI21X1_103 ( );
FILL FILL_3_OAI21X1_103 ( );
FILL FILL_4_OAI21X1_103 ( );
FILL FILL_5_OAI21X1_103 ( );
FILL FILL_6_OAI21X1_103 ( );
FILL FILL_7_OAI21X1_103 ( );
FILL FILL_8_OAI21X1_103 ( );
FILL FILL_9_OAI21X1_103 ( );
FILL FILL_0_INVX1_116 ( );
FILL FILL_1_INVX1_116 ( );
FILL FILL_2_INVX1_116 ( );
FILL FILL_3_INVX1_116 ( );
FILL FILL_0_NAND2X1_111 ( );
FILL FILL_1_NAND2X1_111 ( );
FILL FILL_2_NAND2X1_111 ( );
FILL FILL_3_NAND2X1_111 ( );
FILL FILL_4_NAND2X1_111 ( );
FILL FILL_5_NAND2X1_111 ( );
FILL FILL_6_NAND2X1_111 ( );
FILL FILL_0_OAI21X1_111 ( );
FILL FILL_1_OAI21X1_111 ( );
FILL FILL_2_OAI21X1_111 ( );
FILL FILL_3_OAI21X1_111 ( );
FILL FILL_4_OAI21X1_111 ( );
FILL FILL_5_OAI21X1_111 ( );
FILL FILL_6_OAI21X1_111 ( );
FILL FILL_7_OAI21X1_111 ( );
FILL FILL_8_OAI21X1_111 ( );
FILL FILL_0_INVX1_125 ( );
FILL FILL_1_INVX1_125 ( );
FILL FILL_2_INVX1_125 ( );
FILL FILL_3_INVX1_125 ( );
FILL FILL_4_INVX1_125 ( );
FILL FILL_0_INVX1_384 ( );
FILL FILL_1_INVX1_384 ( );
FILL FILL_2_INVX1_384 ( );
FILL FILL_3_INVX1_384 ( );
FILL FILL_4_INVX1_384 ( );
FILL FILL_0_NAND2X1_114 ( );
FILL FILL_1_NAND2X1_114 ( );
FILL FILL_2_NAND2X1_114 ( );
FILL FILL_3_NAND2X1_114 ( );
FILL FILL_4_NAND2X1_114 ( );
FILL FILL_5_NAND2X1_114 ( );
FILL FILL_6_NAND2X1_114 ( );
FILL FILL_0_OAI22X1_68 ( );
FILL FILL_1_OAI22X1_68 ( );
FILL FILL_2_OAI22X1_68 ( );
FILL FILL_3_OAI22X1_68 ( );
FILL FILL_4_OAI22X1_68 ( );
FILL FILL_5_OAI22X1_68 ( );
FILL FILL_6_OAI22X1_68 ( );
FILL FILL_7_OAI22X1_68 ( );
FILL FILL_8_OAI22X1_68 ( );
FILL FILL_9_OAI22X1_68 ( );
FILL FILL_10_OAI22X1_68 ( );
FILL FILL_11_OAI22X1_68 ( );
FILL FILL_0_INVX1_395 ( );
FILL FILL_1_INVX1_395 ( );
FILL FILL_2_INVX1_395 ( );
FILL FILL_3_INVX1_395 ( );
FILL FILL_0_NAND3X1_121 ( );
FILL FILL_1_NAND3X1_121 ( );
FILL FILL_2_NAND3X1_121 ( );
FILL FILL_3_NAND3X1_121 ( );
FILL FILL_4_NAND3X1_121 ( );
FILL FILL_5_NAND3X1_121 ( );
FILL FILL_6_NAND3X1_121 ( );
FILL FILL_7_NAND3X1_121 ( );
FILL FILL_8_NAND3X1_121 ( );
FILL FILL_9_NAND3X1_121 ( );
FILL FILL_0_NAND3X1_122 ( );
FILL FILL_1_NAND3X1_122 ( );
FILL FILL_2_NAND3X1_122 ( );
FILL FILL_3_NAND3X1_122 ( );
FILL FILL_4_NAND3X1_122 ( );
FILL FILL_5_NAND3X1_122 ( );
FILL FILL_6_NAND3X1_122 ( );
FILL FILL_7_NAND3X1_122 ( );
FILL FILL_8_NAND3X1_122 ( );
FILL FILL_0_NAND3X1_124 ( );
FILL FILL_1_NAND3X1_124 ( );
FILL FILL_2_NAND3X1_124 ( );
FILL FILL_3_NAND3X1_124 ( );
FILL FILL_4_NAND3X1_124 ( );
FILL FILL_5_NAND3X1_124 ( );
FILL FILL_6_NAND3X1_124 ( );
FILL FILL_7_NAND3X1_124 ( );
FILL FILL_8_NAND3X1_124 ( );
FILL FILL_9_NAND3X1_124 ( );
FILL FILL_0_NAND3X1_120 ( );
FILL FILL_1_NAND3X1_120 ( );
FILL FILL_2_NAND3X1_120 ( );
FILL FILL_3_NAND3X1_120 ( );
FILL FILL_4_NAND3X1_120 ( );
FILL FILL_5_NAND3X1_120 ( );
FILL FILL_6_NAND3X1_120 ( );
FILL FILL_7_NAND3X1_120 ( );
FILL FILL_8_NAND3X1_120 ( );
FILL FILL_0_NAND3X1_126 ( );
FILL FILL_1_NAND3X1_126 ( );
FILL FILL_2_NAND3X1_126 ( );
FILL FILL_3_NAND3X1_126 ( );
FILL FILL_4_NAND3X1_126 ( );
FILL FILL_5_NAND3X1_126 ( );
FILL FILL_6_NAND3X1_126 ( );
FILL FILL_7_NAND3X1_126 ( );
FILL FILL_8_NAND3X1_126 ( );
FILL FILL_0_NAND3X1_128 ( );
FILL FILL_1_NAND3X1_128 ( );
FILL FILL_2_NAND3X1_128 ( );
FILL FILL_3_NAND3X1_128 ( );
FILL FILL_4_NAND3X1_128 ( );
FILL FILL_5_NAND3X1_128 ( );
FILL FILL_6_NAND3X1_128 ( );
FILL FILL_7_NAND3X1_128 ( );
FILL FILL_8_NAND3X1_128 ( );
FILL FILL_0_OAI21X1_240 ( );
FILL FILL_1_OAI21X1_240 ( );
FILL FILL_2_OAI21X1_240 ( );
FILL FILL_3_OAI21X1_240 ( );
FILL FILL_4_OAI21X1_240 ( );
FILL FILL_5_OAI21X1_240 ( );
FILL FILL_6_OAI21X1_240 ( );
FILL FILL_7_OAI21X1_240 ( );
FILL FILL_8_OAI21X1_240 ( );
FILL FILL_9_OAI21X1_240 ( );
FILL FILL_0_INVX1_396 ( );
FILL FILL_1_INVX1_396 ( );
FILL FILL_2_INVX1_396 ( );
FILL FILL_3_INVX1_396 ( );
FILL FILL_4_INVX1_396 ( );
FILL FILL_0_DFFSR_136 ( );
FILL FILL_1_DFFSR_136 ( );
FILL FILL_2_DFFSR_136 ( );
FILL FILL_3_DFFSR_136 ( );
FILL FILL_4_DFFSR_136 ( );
FILL FILL_5_DFFSR_136 ( );
FILL FILL_6_DFFSR_136 ( );
FILL FILL_7_DFFSR_136 ( );
FILL FILL_8_DFFSR_136 ( );
FILL FILL_9_DFFSR_136 ( );
FILL FILL_10_DFFSR_136 ( );
FILL FILL_11_DFFSR_136 ( );
FILL FILL_12_DFFSR_136 ( );
FILL FILL_13_DFFSR_136 ( );
FILL FILL_14_DFFSR_136 ( );
FILL FILL_15_DFFSR_136 ( );
FILL FILL_16_DFFSR_136 ( );
FILL FILL_17_DFFSR_136 ( );
FILL FILL_18_DFFSR_136 ( );
FILL FILL_19_DFFSR_136 ( );
FILL FILL_20_DFFSR_136 ( );
FILL FILL_21_DFFSR_136 ( );
FILL FILL_22_DFFSR_136 ( );
FILL FILL_23_DFFSR_136 ( );
FILL FILL_24_DFFSR_136 ( );
FILL FILL_25_DFFSR_136 ( );
FILL FILL_26_DFFSR_136 ( );
FILL FILL_27_DFFSR_136 ( );
FILL FILL_28_DFFSR_136 ( );
FILL FILL_29_DFFSR_136 ( );
FILL FILL_30_DFFSR_136 ( );
FILL FILL_31_DFFSR_136 ( );
FILL FILL_32_DFFSR_136 ( );
FILL FILL_33_DFFSR_136 ( );
FILL FILL_34_DFFSR_136 ( );
FILL FILL_35_DFFSR_136 ( );
FILL FILL_36_DFFSR_136 ( );
FILL FILL_37_DFFSR_136 ( );
FILL FILL_38_DFFSR_136 ( );
FILL FILL_39_DFFSR_136 ( );
FILL FILL_40_DFFSR_136 ( );
FILL FILL_41_DFFSR_136 ( );
FILL FILL_42_DFFSR_136 ( );
FILL FILL_43_DFFSR_136 ( );
FILL FILL_44_DFFSR_136 ( );
FILL FILL_45_DFFSR_136 ( );
FILL FILL_46_DFFSR_136 ( );
FILL FILL_47_DFFSR_136 ( );
FILL FILL_48_DFFSR_136 ( );
FILL FILL_49_DFFSR_136 ( );
FILL FILL_50_DFFSR_136 ( );
FILL FILL_0_AND2X2_17 ( );
FILL FILL_1_AND2X2_17 ( );
FILL FILL_2_AND2X2_17 ( );
FILL FILL_3_AND2X2_17 ( );
FILL FILL_4_AND2X2_17 ( );
FILL FILL_5_AND2X2_17 ( );
FILL FILL_6_AND2X2_17 ( );
FILL FILL_7_AND2X2_17 ( );
FILL FILL_8_AND2X2_17 ( );
FILL FILL_0_AOI21X1_46 ( );
FILL FILL_1_AOI21X1_46 ( );
FILL FILL_2_AOI21X1_46 ( );
FILL FILL_3_AOI21X1_46 ( );
FILL FILL_4_AOI21X1_46 ( );
FILL FILL_5_AOI21X1_46 ( );
FILL FILL_6_AOI21X1_46 ( );
FILL FILL_7_AOI21X1_46 ( );
FILL FILL_8_AOI21X1_46 ( );
FILL FILL_0_OAI21X1_264 ( );
FILL FILL_1_OAI21X1_264 ( );
FILL FILL_2_OAI21X1_264 ( );
FILL FILL_3_OAI21X1_264 ( );
FILL FILL_4_OAI21X1_264 ( );
FILL FILL_5_OAI21X1_264 ( );
FILL FILL_6_OAI21X1_264 ( );
FILL FILL_7_OAI21X1_264 ( );
FILL FILL_8_OAI21X1_264 ( );
FILL FILL_0_NAND2X1_275 ( );
FILL FILL_1_NAND2X1_275 ( );
FILL FILL_2_NAND2X1_275 ( );
FILL FILL_3_NAND2X1_275 ( );
FILL FILL_4_NAND2X1_275 ( );
FILL FILL_5_NAND2X1_275 ( );
FILL FILL_6_NAND2X1_275 ( );
FILL FILL_0_OAI21X1_263 ( );
FILL FILL_1_OAI21X1_263 ( );
FILL FILL_2_OAI21X1_263 ( );
FILL FILL_3_OAI21X1_263 ( );
FILL FILL_4_OAI21X1_263 ( );
FILL FILL_5_OAI21X1_263 ( );
FILL FILL_6_OAI21X1_263 ( );
FILL FILL_7_OAI21X1_263 ( );
FILL FILL_8_OAI21X1_263 ( );
FILL FILL_0_OAI21X1_38 ( );
FILL FILL_1_OAI21X1_38 ( );
FILL FILL_2_OAI21X1_38 ( );
FILL FILL_3_OAI21X1_38 ( );
FILL FILL_4_OAI21X1_38 ( );
FILL FILL_5_OAI21X1_38 ( );
FILL FILL_6_OAI21X1_38 ( );
FILL FILL_7_OAI21X1_38 ( );
FILL FILL_8_OAI21X1_38 ( );
FILL FILL_9_OAI21X1_38 ( );
FILL FILL_0_NAND2X1_38 ( );
FILL FILL_1_NAND2X1_38 ( );
FILL FILL_2_NAND2X1_38 ( );
FILL FILL_3_NAND2X1_38 ( );
FILL FILL_4_NAND2X1_38 ( );
FILL FILL_5_NAND2X1_38 ( );
FILL FILL_6_NAND2X1_38 ( );
FILL FILL_0_INVX1_43 ( );
FILL FILL_1_INVX1_43 ( );
FILL FILL_2_INVX1_43 ( );
FILL FILL_3_INVX1_43 ( );
FILL FILL_0_INVX1_269 ( );
FILL FILL_1_INVX1_269 ( );
FILL FILL_2_INVX1_269 ( );
FILL FILL_3_INVX1_269 ( );
FILL FILL_4_INVX1_269 ( );
FILL FILL_0_OAI22X1_7 ( );
FILL FILL_1_OAI22X1_7 ( );
FILL FILL_2_OAI22X1_7 ( );
FILL FILL_3_OAI22X1_7 ( );
FILL FILL_4_OAI22X1_7 ( );
FILL FILL_5_OAI22X1_7 ( );
FILL FILL_6_OAI22X1_7 ( );
FILL FILL_7_OAI22X1_7 ( );
FILL FILL_8_OAI22X1_7 ( );
FILL FILL_9_OAI22X1_7 ( );
FILL FILL_10_OAI22X1_7 ( );
FILL FILL_11_OAI22X1_7 ( );
FILL FILL_0_NAND2X1_41 ( );
FILL FILL_1_NAND2X1_41 ( );
FILL FILL_2_NAND2X1_41 ( );
FILL FILL_3_NAND2X1_41 ( );
FILL FILL_4_NAND2X1_41 ( );
FILL FILL_5_NAND2X1_41 ( );
FILL FILL_6_NAND2X1_41 ( );
FILL FILL_0_DFFSR_17 ( );
FILL FILL_1_DFFSR_17 ( );
FILL FILL_2_DFFSR_17 ( );
FILL FILL_3_DFFSR_17 ( );
FILL FILL_4_DFFSR_17 ( );
FILL FILL_5_DFFSR_17 ( );
FILL FILL_6_DFFSR_17 ( );
FILL FILL_7_DFFSR_17 ( );
FILL FILL_8_DFFSR_17 ( );
FILL FILL_9_DFFSR_17 ( );
FILL FILL_10_DFFSR_17 ( );
FILL FILL_11_DFFSR_17 ( );
FILL FILL_12_DFFSR_17 ( );
FILL FILL_13_DFFSR_17 ( );
FILL FILL_14_DFFSR_17 ( );
FILL FILL_15_DFFSR_17 ( );
FILL FILL_16_DFFSR_17 ( );
FILL FILL_17_DFFSR_17 ( );
FILL FILL_18_DFFSR_17 ( );
FILL FILL_19_DFFSR_17 ( );
FILL FILL_20_DFFSR_17 ( );
FILL FILL_21_DFFSR_17 ( );
FILL FILL_22_DFFSR_17 ( );
FILL FILL_23_DFFSR_17 ( );
FILL FILL_24_DFFSR_17 ( );
FILL FILL_25_DFFSR_17 ( );
FILL FILL_26_DFFSR_17 ( );
FILL FILL_27_DFFSR_17 ( );
FILL FILL_28_DFFSR_17 ( );
FILL FILL_29_DFFSR_17 ( );
FILL FILL_30_DFFSR_17 ( );
FILL FILL_31_DFFSR_17 ( );
FILL FILL_32_DFFSR_17 ( );
FILL FILL_33_DFFSR_17 ( );
FILL FILL_34_DFFSR_17 ( );
FILL FILL_35_DFFSR_17 ( );
FILL FILL_36_DFFSR_17 ( );
FILL FILL_37_DFFSR_17 ( );
FILL FILL_38_DFFSR_17 ( );
FILL FILL_39_DFFSR_17 ( );
FILL FILL_40_DFFSR_17 ( );
FILL FILL_41_DFFSR_17 ( );
FILL FILL_42_DFFSR_17 ( );
FILL FILL_43_DFFSR_17 ( );
FILL FILL_44_DFFSR_17 ( );
FILL FILL_45_DFFSR_17 ( );
FILL FILL_46_DFFSR_17 ( );
FILL FILL_47_DFFSR_17 ( );
FILL FILL_48_DFFSR_17 ( );
FILL FILL_49_DFFSR_17 ( );
FILL FILL_50_DFFSR_17 ( );
FILL FILL_0_NAND2X1_10 ( );
FILL FILL_1_NAND2X1_10 ( );
FILL FILL_2_NAND2X1_10 ( );
FILL FILL_3_NAND2X1_10 ( );
FILL FILL_4_NAND2X1_10 ( );
FILL FILL_5_NAND2X1_10 ( );
FILL FILL_6_NAND2X1_10 ( );
FILL FILL_0_DFFSR_5 ( );
FILL FILL_1_DFFSR_5 ( );
FILL FILL_2_DFFSR_5 ( );
FILL FILL_3_DFFSR_5 ( );
FILL FILL_4_DFFSR_5 ( );
FILL FILL_5_DFFSR_5 ( );
FILL FILL_6_DFFSR_5 ( );
FILL FILL_7_DFFSR_5 ( );
FILL FILL_8_DFFSR_5 ( );
FILL FILL_9_DFFSR_5 ( );
FILL FILL_10_DFFSR_5 ( );
FILL FILL_11_DFFSR_5 ( );
FILL FILL_12_DFFSR_5 ( );
FILL FILL_13_DFFSR_5 ( );
FILL FILL_14_DFFSR_5 ( );
FILL FILL_15_DFFSR_5 ( );
FILL FILL_16_DFFSR_5 ( );
FILL FILL_17_DFFSR_5 ( );
FILL FILL_18_DFFSR_5 ( );
FILL FILL_19_DFFSR_5 ( );
FILL FILL_20_DFFSR_5 ( );
FILL FILL_21_DFFSR_5 ( );
FILL FILL_22_DFFSR_5 ( );
FILL FILL_23_DFFSR_5 ( );
FILL FILL_24_DFFSR_5 ( );
FILL FILL_25_DFFSR_5 ( );
FILL FILL_26_DFFSR_5 ( );
FILL FILL_27_DFFSR_5 ( );
FILL FILL_28_DFFSR_5 ( );
FILL FILL_29_DFFSR_5 ( );
FILL FILL_30_DFFSR_5 ( );
FILL FILL_31_DFFSR_5 ( );
FILL FILL_32_DFFSR_5 ( );
FILL FILL_33_DFFSR_5 ( );
FILL FILL_34_DFFSR_5 ( );
FILL FILL_35_DFFSR_5 ( );
FILL FILL_36_DFFSR_5 ( );
FILL FILL_37_DFFSR_5 ( );
FILL FILL_38_DFFSR_5 ( );
FILL FILL_39_DFFSR_5 ( );
FILL FILL_40_DFFSR_5 ( );
FILL FILL_41_DFFSR_5 ( );
FILL FILL_42_DFFSR_5 ( );
FILL FILL_43_DFFSR_5 ( );
FILL FILL_44_DFFSR_5 ( );
FILL FILL_45_DFFSR_5 ( );
FILL FILL_46_DFFSR_5 ( );
FILL FILL_47_DFFSR_5 ( );
FILL FILL_48_DFFSR_5 ( );
FILL FILL_49_DFFSR_5 ( );
FILL FILL_50_DFFSR_5 ( );
FILL FILL_51_DFFSR_5 ( );
FILL FILL_0_NAND3X1_18 ( );
FILL FILL_1_NAND3X1_18 ( );
FILL FILL_2_NAND3X1_18 ( );
FILL FILL_3_NAND3X1_18 ( );
FILL FILL_4_NAND3X1_18 ( );
FILL FILL_5_NAND3X1_18 ( );
FILL FILL_6_NAND3X1_18 ( );
FILL FILL_7_NAND3X1_18 ( );
FILL FILL_8_NAND3X1_18 ( );
FILL FILL_0_DFFSR_177 ( );
FILL FILL_1_DFFSR_177 ( );
FILL FILL_2_DFFSR_177 ( );
FILL FILL_3_DFFSR_177 ( );
FILL FILL_4_DFFSR_177 ( );
FILL FILL_5_DFFSR_177 ( );
FILL FILL_6_DFFSR_177 ( );
FILL FILL_7_DFFSR_177 ( );
FILL FILL_8_DFFSR_177 ( );
FILL FILL_9_DFFSR_177 ( );
FILL FILL_10_DFFSR_177 ( );
FILL FILL_11_DFFSR_177 ( );
FILL FILL_12_DFFSR_177 ( );
FILL FILL_13_DFFSR_177 ( );
FILL FILL_14_DFFSR_177 ( );
FILL FILL_15_DFFSR_177 ( );
FILL FILL_16_DFFSR_177 ( );
FILL FILL_17_DFFSR_177 ( );
FILL FILL_18_DFFSR_177 ( );
FILL FILL_19_DFFSR_177 ( );
FILL FILL_20_DFFSR_177 ( );
FILL FILL_21_DFFSR_177 ( );
FILL FILL_22_DFFSR_177 ( );
FILL FILL_23_DFFSR_177 ( );
FILL FILL_24_DFFSR_177 ( );
FILL FILL_25_DFFSR_177 ( );
FILL FILL_26_DFFSR_177 ( );
FILL FILL_27_DFFSR_177 ( );
FILL FILL_28_DFFSR_177 ( );
FILL FILL_29_DFFSR_177 ( );
FILL FILL_30_DFFSR_177 ( );
FILL FILL_31_DFFSR_177 ( );
FILL FILL_32_DFFSR_177 ( );
FILL FILL_33_DFFSR_177 ( );
FILL FILL_34_DFFSR_177 ( );
FILL FILL_35_DFFSR_177 ( );
FILL FILL_36_DFFSR_177 ( );
FILL FILL_37_DFFSR_177 ( );
FILL FILL_38_DFFSR_177 ( );
FILL FILL_39_DFFSR_177 ( );
FILL FILL_40_DFFSR_177 ( );
FILL FILL_41_DFFSR_177 ( );
FILL FILL_42_DFFSR_177 ( );
FILL FILL_43_DFFSR_177 ( );
FILL FILL_44_DFFSR_177 ( );
FILL FILL_45_DFFSR_177 ( );
FILL FILL_46_DFFSR_177 ( );
FILL FILL_47_DFFSR_177 ( );
FILL FILL_48_DFFSR_177 ( );
FILL FILL_49_DFFSR_177 ( );
FILL FILL_50_DFFSR_177 ( );
FILL FILL_0_DFFSR_111 ( );
FILL FILL_1_DFFSR_111 ( );
FILL FILL_2_DFFSR_111 ( );
FILL FILL_3_DFFSR_111 ( );
FILL FILL_4_DFFSR_111 ( );
FILL FILL_5_DFFSR_111 ( );
FILL FILL_6_DFFSR_111 ( );
FILL FILL_7_DFFSR_111 ( );
FILL FILL_8_DFFSR_111 ( );
FILL FILL_9_DFFSR_111 ( );
FILL FILL_10_DFFSR_111 ( );
FILL FILL_11_DFFSR_111 ( );
FILL FILL_12_DFFSR_111 ( );
FILL FILL_13_DFFSR_111 ( );
FILL FILL_14_DFFSR_111 ( );
FILL FILL_15_DFFSR_111 ( );
FILL FILL_16_DFFSR_111 ( );
FILL FILL_17_DFFSR_111 ( );
FILL FILL_18_DFFSR_111 ( );
FILL FILL_19_DFFSR_111 ( );
FILL FILL_20_DFFSR_111 ( );
FILL FILL_21_DFFSR_111 ( );
FILL FILL_22_DFFSR_111 ( );
FILL FILL_23_DFFSR_111 ( );
FILL FILL_24_DFFSR_111 ( );
FILL FILL_25_DFFSR_111 ( );
FILL FILL_26_DFFSR_111 ( );
FILL FILL_27_DFFSR_111 ( );
FILL FILL_28_DFFSR_111 ( );
FILL FILL_29_DFFSR_111 ( );
FILL FILL_30_DFFSR_111 ( );
FILL FILL_31_DFFSR_111 ( );
FILL FILL_32_DFFSR_111 ( );
FILL FILL_33_DFFSR_111 ( );
FILL FILL_34_DFFSR_111 ( );
FILL FILL_35_DFFSR_111 ( );
FILL FILL_36_DFFSR_111 ( );
FILL FILL_37_DFFSR_111 ( );
FILL FILL_38_DFFSR_111 ( );
FILL FILL_39_DFFSR_111 ( );
FILL FILL_40_DFFSR_111 ( );
FILL FILL_41_DFFSR_111 ( );
FILL FILL_42_DFFSR_111 ( );
FILL FILL_43_DFFSR_111 ( );
FILL FILL_44_DFFSR_111 ( );
FILL FILL_45_DFFSR_111 ( );
FILL FILL_46_DFFSR_111 ( );
FILL FILL_47_DFFSR_111 ( );
FILL FILL_48_DFFSR_111 ( );
FILL FILL_49_DFFSR_111 ( );
FILL FILL_50_DFFSR_111 ( );
FILL FILL_51_DFFSR_111 ( );
FILL FILL_0_OAI22X1_60 ( );
FILL FILL_1_OAI22X1_60 ( );
FILL FILL_2_OAI22X1_60 ( );
FILL FILL_3_OAI22X1_60 ( );
FILL FILL_4_OAI22X1_60 ( );
FILL FILL_5_OAI22X1_60 ( );
FILL FILL_6_OAI22X1_60 ( );
FILL FILL_7_OAI22X1_60 ( );
FILL FILL_8_OAI22X1_60 ( );
FILL FILL_9_OAI22X1_60 ( );
FILL FILL_10_OAI22X1_60 ( );
FILL FILL_11_OAI22X1_60 ( );
FILL FILL_0_NOR2X1_39 ( );
FILL FILL_1_NOR2X1_39 ( );
FILL FILL_2_NOR2X1_39 ( );
FILL FILL_3_NOR2X1_39 ( );
FILL FILL_4_NOR2X1_39 ( );
FILL FILL_5_NOR2X1_39 ( );
FILL FILL_6_NOR2X1_39 ( );
FILL FILL_0_NAND2X1_247 ( );
FILL FILL_1_NAND2X1_247 ( );
FILL FILL_2_NAND2X1_247 ( );
FILL FILL_3_NAND2X1_247 ( );
FILL FILL_4_NAND2X1_247 ( );
FILL FILL_5_NAND2X1_247 ( );
FILL FILL_6_NAND2X1_247 ( );
FILL FILL_0_NAND3X1_125 ( );
FILL FILL_1_NAND3X1_125 ( );
FILL FILL_2_NAND3X1_125 ( );
FILL FILL_3_NAND3X1_125 ( );
FILL FILL_4_NAND3X1_125 ( );
FILL FILL_5_NAND3X1_125 ( );
FILL FILL_6_NAND3X1_125 ( );
FILL FILL_7_NAND3X1_125 ( );
FILL FILL_8_NAND3X1_125 ( );
FILL FILL_0_DFFPOSX1_12 ( );
FILL FILL_1_DFFPOSX1_12 ( );
FILL FILL_2_DFFPOSX1_12 ( );
FILL FILL_3_DFFPOSX1_12 ( );
FILL FILL_4_DFFPOSX1_12 ( );
FILL FILL_5_DFFPOSX1_12 ( );
FILL FILL_6_DFFPOSX1_12 ( );
FILL FILL_7_DFFPOSX1_12 ( );
FILL FILL_8_DFFPOSX1_12 ( );
FILL FILL_9_DFFPOSX1_12 ( );
FILL FILL_10_DFFPOSX1_12 ( );
FILL FILL_11_DFFPOSX1_12 ( );
FILL FILL_12_DFFPOSX1_12 ( );
FILL FILL_13_DFFPOSX1_12 ( );
FILL FILL_14_DFFPOSX1_12 ( );
FILL FILL_15_DFFPOSX1_12 ( );
FILL FILL_16_DFFPOSX1_12 ( );
FILL FILL_17_DFFPOSX1_12 ( );
FILL FILL_18_DFFPOSX1_12 ( );
FILL FILL_19_DFFPOSX1_12 ( );
FILL FILL_20_DFFPOSX1_12 ( );
FILL FILL_21_DFFPOSX1_12 ( );
FILL FILL_22_DFFPOSX1_12 ( );
FILL FILL_23_DFFPOSX1_12 ( );
FILL FILL_24_DFFPOSX1_12 ( );
FILL FILL_25_DFFPOSX1_12 ( );
FILL FILL_26_DFFPOSX1_12 ( );
FILL FILL_27_DFFPOSX1_12 ( );
FILL FILL_0_NAND2X1_250 ( );
FILL FILL_1_NAND2X1_250 ( );
FILL FILL_2_NAND2X1_250 ( );
FILL FILL_3_NAND2X1_250 ( );
FILL FILL_4_NAND2X1_250 ( );
FILL FILL_5_NAND2X1_250 ( );
FILL FILL_6_NAND2X1_250 ( );
FILL FILL_0_DFFPOSX1_10 ( );
FILL FILL_1_DFFPOSX1_10 ( );
FILL FILL_2_DFFPOSX1_10 ( );
FILL FILL_3_DFFPOSX1_10 ( );
FILL FILL_4_DFFPOSX1_10 ( );
FILL FILL_5_DFFPOSX1_10 ( );
FILL FILL_6_DFFPOSX1_10 ( );
FILL FILL_7_DFFPOSX1_10 ( );
FILL FILL_8_DFFPOSX1_10 ( );
FILL FILL_9_DFFPOSX1_10 ( );
FILL FILL_10_DFFPOSX1_10 ( );
FILL FILL_11_DFFPOSX1_10 ( );
FILL FILL_12_DFFPOSX1_10 ( );
FILL FILL_13_DFFPOSX1_10 ( );
FILL FILL_14_DFFPOSX1_10 ( );
FILL FILL_15_DFFPOSX1_10 ( );
FILL FILL_16_DFFPOSX1_10 ( );
FILL FILL_17_DFFPOSX1_10 ( );
FILL FILL_18_DFFPOSX1_10 ( );
FILL FILL_19_DFFPOSX1_10 ( );
FILL FILL_20_DFFPOSX1_10 ( );
FILL FILL_21_DFFPOSX1_10 ( );
FILL FILL_22_DFFPOSX1_10 ( );
FILL FILL_23_DFFPOSX1_10 ( );
FILL FILL_24_DFFPOSX1_10 ( );
FILL FILL_25_DFFPOSX1_10 ( );
FILL FILL_26_DFFPOSX1_10 ( );
FILL FILL_27_DFFPOSX1_10 ( );
FILL FILL_0_DFFSR_144 ( );
FILL FILL_1_DFFSR_144 ( );
FILL FILL_2_DFFSR_144 ( );
FILL FILL_3_DFFSR_144 ( );
FILL FILL_4_DFFSR_144 ( );
FILL FILL_5_DFFSR_144 ( );
FILL FILL_6_DFFSR_144 ( );
FILL FILL_7_DFFSR_144 ( );
FILL FILL_8_DFFSR_144 ( );
FILL FILL_9_DFFSR_144 ( );
FILL FILL_10_DFFSR_144 ( );
FILL FILL_11_DFFSR_144 ( );
FILL FILL_12_DFFSR_144 ( );
FILL FILL_13_DFFSR_144 ( );
FILL FILL_14_DFFSR_144 ( );
FILL FILL_15_DFFSR_144 ( );
FILL FILL_16_DFFSR_144 ( );
FILL FILL_17_DFFSR_144 ( );
FILL FILL_18_DFFSR_144 ( );
FILL FILL_19_DFFSR_144 ( );
FILL FILL_20_DFFSR_144 ( );
FILL FILL_21_DFFSR_144 ( );
FILL FILL_22_DFFSR_144 ( );
FILL FILL_23_DFFSR_144 ( );
FILL FILL_24_DFFSR_144 ( );
FILL FILL_25_DFFSR_144 ( );
FILL FILL_26_DFFSR_144 ( );
FILL FILL_27_DFFSR_144 ( );
FILL FILL_28_DFFSR_144 ( );
FILL FILL_29_DFFSR_144 ( );
FILL FILL_30_DFFSR_144 ( );
FILL FILL_31_DFFSR_144 ( );
FILL FILL_32_DFFSR_144 ( );
FILL FILL_33_DFFSR_144 ( );
FILL FILL_34_DFFSR_144 ( );
FILL FILL_35_DFFSR_144 ( );
FILL FILL_36_DFFSR_144 ( );
FILL FILL_37_DFFSR_144 ( );
FILL FILL_38_DFFSR_144 ( );
FILL FILL_39_DFFSR_144 ( );
FILL FILL_40_DFFSR_144 ( );
FILL FILL_41_DFFSR_144 ( );
FILL FILL_42_DFFSR_144 ( );
FILL FILL_43_DFFSR_144 ( );
FILL FILL_44_DFFSR_144 ( );
FILL FILL_45_DFFSR_144 ( );
FILL FILL_46_DFFSR_144 ( );
FILL FILL_47_DFFSR_144 ( );
FILL FILL_48_DFFSR_144 ( );
FILL FILL_49_DFFSR_144 ( );
FILL FILL_50_DFFSR_144 ( );
FILL FILL_0_NAND2X1_132 ( );
FILL FILL_1_NAND2X1_132 ( );
FILL FILL_2_NAND2X1_132 ( );
FILL FILL_3_NAND2X1_132 ( );
FILL FILL_4_NAND2X1_132 ( );
FILL FILL_5_NAND2X1_132 ( );
FILL FILL_6_NAND2X1_132 ( );
FILL FILL_0_INVX1_45 ( );
FILL FILL_1_INVX1_45 ( );
FILL FILL_2_INVX1_45 ( );
FILL FILL_3_INVX1_45 ( );
FILL FILL_0_XOR2X1_16 ( );
FILL FILL_1_XOR2X1_16 ( );
FILL FILL_2_XOR2X1_16 ( );
FILL FILL_3_XOR2X1_16 ( );
FILL FILL_4_XOR2X1_16 ( );
FILL FILL_5_XOR2X1_16 ( );
FILL FILL_6_XOR2X1_16 ( );
FILL FILL_7_XOR2X1_16 ( );
FILL FILL_8_XOR2X1_16 ( );
FILL FILL_9_XOR2X1_16 ( );
FILL FILL_10_XOR2X1_16 ( );
FILL FILL_11_XOR2X1_16 ( );
FILL FILL_12_XOR2X1_16 ( );
FILL FILL_13_XOR2X1_16 ( );
FILL FILL_14_XOR2X1_16 ( );
FILL FILL_15_XOR2X1_16 ( );
FILL FILL_0_INVX1_435 ( );
FILL FILL_1_INVX1_435 ( );
FILL FILL_2_INVX1_435 ( );
FILL FILL_3_INVX1_435 ( );
FILL FILL_4_INVX1_435 ( );
FILL FILL_0_INVX1_434 ( );
FILL FILL_1_INVX1_434 ( );
FILL FILL_2_INVX1_434 ( );
FILL FILL_3_INVX1_434 ( );
FILL FILL_4_INVX1_434 ( );
FILL FILL_0_NAND3X1_133 ( );
FILL FILL_1_NAND3X1_133 ( );
FILL FILL_2_NAND3X1_133 ( );
FILL FILL_3_NAND3X1_133 ( );
FILL FILL_4_NAND3X1_133 ( );
FILL FILL_5_NAND3X1_133 ( );
FILL FILL_6_NAND3X1_133 ( );
FILL FILL_7_NAND3X1_133 ( );
FILL FILL_8_NAND3X1_133 ( );
FILL FILL_9_NAND3X1_133 ( );
FILL FILL_0_NAND2X1_284 ( );
FILL FILL_1_NAND2X1_284 ( );
FILL FILL_2_NAND2X1_284 ( );
FILL FILL_3_NAND2X1_284 ( );
FILL FILL_4_NAND2X1_284 ( );
FILL FILL_5_NAND2X1_284 ( );
FILL FILL_6_NAND2X1_284 ( );
FILL FILL_0_INVX1_314 ( );
FILL FILL_1_INVX1_314 ( );
FILL FILL_2_INVX1_314 ( );
FILL FILL_3_INVX1_314 ( );
FILL FILL_4_INVX1_314 ( );
FILL FILL_0_OAI22X1_29 ( );
FILL FILL_1_OAI22X1_29 ( );
FILL FILL_2_OAI22X1_29 ( );
FILL FILL_3_OAI22X1_29 ( );
FILL FILL_4_OAI22X1_29 ( );
FILL FILL_5_OAI22X1_29 ( );
FILL FILL_6_OAI22X1_29 ( );
FILL FILL_7_OAI22X1_29 ( );
FILL FILL_8_OAI22X1_29 ( );
FILL FILL_9_OAI22X1_29 ( );
FILL FILL_10_OAI22X1_29 ( );
FILL FILL_0_INVX1_313 ( );
FILL FILL_1_INVX1_313 ( );
FILL FILL_2_INVX1_313 ( );
FILL FILL_3_INVX1_313 ( );
FILL FILL_4_INVX1_313 ( );
FILL FILL_0_INVX1_274 ( );
FILL FILL_1_INVX1_274 ( );
FILL FILL_2_INVX1_274 ( );
FILL FILL_3_INVX1_274 ( );
FILL FILL_4_INVX1_274 ( );
FILL FILL_0_OAI22X1_9 ( );
FILL FILL_1_OAI22X1_9 ( );
FILL FILL_2_OAI22X1_9 ( );
FILL FILL_3_OAI22X1_9 ( );
FILL FILL_4_OAI22X1_9 ( );
FILL FILL_5_OAI22X1_9 ( );
FILL FILL_6_OAI22X1_9 ( );
FILL FILL_7_OAI22X1_9 ( );
FILL FILL_8_OAI22X1_9 ( );
FILL FILL_9_OAI22X1_9 ( );
FILL FILL_10_OAI22X1_9 ( );
FILL FILL_11_OAI22X1_9 ( );
FILL FILL_0_INVX1_40 ( );
FILL FILL_1_INVX1_40 ( );
FILL FILL_2_INVX1_40 ( );
FILL FILL_3_INVX1_40 ( );
FILL FILL_0_OAI21X1_35 ( );
FILL FILL_1_OAI21X1_35 ( );
FILL FILL_2_OAI21X1_35 ( );
FILL FILL_3_OAI21X1_35 ( );
FILL FILL_4_OAI21X1_35 ( );
FILL FILL_5_OAI21X1_35 ( );
FILL FILL_6_OAI21X1_35 ( );
FILL FILL_7_OAI21X1_35 ( );
FILL FILL_8_OAI21X1_35 ( );
FILL FILL_9_OAI21X1_35 ( );
FILL FILL_0_OAI21X1_17 ( );
FILL FILL_1_OAI21X1_17 ( );
FILL FILL_2_OAI21X1_17 ( );
FILL FILL_3_OAI21X1_17 ( );
FILL FILL_4_OAI21X1_17 ( );
FILL FILL_5_OAI21X1_17 ( );
FILL FILL_6_OAI21X1_17 ( );
FILL FILL_7_OAI21X1_17 ( );
FILL FILL_8_OAI21X1_17 ( );
FILL FILL_0_INVX1_20 ( );
FILL FILL_1_INVX1_20 ( );
FILL FILL_2_INVX1_20 ( );
FILL FILL_3_INVX1_20 ( );
FILL FILL_4_INVX1_20 ( );
FILL FILL_0_INVX1_273 ( );
FILL FILL_1_INVX1_273 ( );
FILL FILL_2_INVX1_273 ( );
FILL FILL_3_INVX1_273 ( );
FILL FILL_0_INVX1_8 ( );
FILL FILL_1_INVX1_8 ( );
FILL FILL_2_INVX1_8 ( );
FILL FILL_3_INVX1_8 ( );
FILL FILL_4_INVX1_8 ( );
FILL FILL_0_OAI21X1_7 ( );
FILL FILL_1_OAI21X1_7 ( );
FILL FILL_2_OAI21X1_7 ( );
FILL FILL_3_OAI21X1_7 ( );
FILL FILL_4_OAI21X1_7 ( );
FILL FILL_5_OAI21X1_7 ( );
FILL FILL_6_OAI21X1_7 ( );
FILL FILL_7_OAI21X1_7 ( );
FILL FILL_8_OAI21X1_7 ( );
FILL FILL_9_OAI21X1_7 ( );
FILL FILL_0_NAND2X1_37 ( );
FILL FILL_1_NAND2X1_37 ( );
FILL FILL_2_NAND2X1_37 ( );
FILL FILL_3_NAND2X1_37 ( );
FILL FILL_4_NAND2X1_37 ( );
FILL FILL_5_NAND2X1_37 ( );
FILL FILL_6_NAND2X1_37 ( );
FILL FILL_0_INVX1_3 ( );
FILL FILL_1_INVX1_3 ( );
FILL FILL_2_INVX1_3 ( );
FILL FILL_3_INVX1_3 ( );
FILL FILL_4_INVX1_3 ( );
FILL FILL_0_OAI21X1_2 ( );
FILL FILL_1_OAI21X1_2 ( );
FILL FILL_2_OAI21X1_2 ( );
FILL FILL_3_OAI21X1_2 ( );
FILL FILL_4_OAI21X1_2 ( );
FILL FILL_5_OAI21X1_2 ( );
FILL FILL_6_OAI21X1_2 ( );
FILL FILL_7_OAI21X1_2 ( );
FILL FILL_8_OAI21X1_2 ( );
FILL FILL_0_AOI21X1_1 ( );
FILL FILL_1_AOI21X1_1 ( );
FILL FILL_2_AOI21X1_1 ( );
FILL FILL_3_AOI21X1_1 ( );
FILL FILL_4_AOI21X1_1 ( );
FILL FILL_5_AOI21X1_1 ( );
FILL FILL_6_AOI21X1_1 ( );
FILL FILL_7_AOI21X1_1 ( );
FILL FILL_8_AOI21X1_1 ( );
FILL FILL_0_OAI21X1_5 ( );
FILL FILL_1_OAI21X1_5 ( );
FILL FILL_2_OAI21X1_5 ( );
FILL FILL_3_OAI21X1_5 ( );
FILL FILL_4_OAI21X1_5 ( );
FILL FILL_5_OAI21X1_5 ( );
FILL FILL_6_OAI21X1_5 ( );
FILL FILL_7_OAI21X1_5 ( );
FILL FILL_8_OAI21X1_5 ( );
FILL FILL_0_INVX1_6 ( );
FILL FILL_1_INVX1_6 ( );
FILL FILL_2_INVX1_6 ( );
FILL FILL_3_INVX1_6 ( );
FILL FILL_4_INVX1_6 ( );
FILL FILL_0_NAND2X1_2 ( );
FILL FILL_1_NAND2X1_2 ( );
FILL FILL_2_NAND2X1_2 ( );
FILL FILL_3_NAND2X1_2 ( );
FILL FILL_4_NAND2X1_2 ( );
FILL FILL_5_NAND2X1_2 ( );
FILL FILL_6_NAND2X1_2 ( );
FILL FILL_0_NAND3X1_19 ( );
FILL FILL_1_NAND3X1_19 ( );
FILL FILL_2_NAND3X1_19 ( );
FILL FILL_3_NAND3X1_19 ( );
FILL FILL_4_NAND3X1_19 ( );
FILL FILL_5_NAND3X1_19 ( );
FILL FILL_6_NAND3X1_19 ( );
FILL FILL_7_NAND3X1_19 ( );
FILL FILL_8_NAND3X1_19 ( );
FILL FILL_0_NAND2X1_160 ( );
FILL FILL_1_NAND2X1_160 ( );
FILL FILL_2_NAND2X1_160 ( );
FILL FILL_3_NAND2X1_160 ( );
FILL FILL_4_NAND2X1_160 ( );
FILL FILL_5_NAND2X1_160 ( );
FILL FILL_6_NAND2X1_160 ( );
FILL FILL_0_AOI21X1_11 ( );
FILL FILL_1_AOI21X1_11 ( );
FILL FILL_2_AOI21X1_11 ( );
FILL FILL_3_AOI21X1_11 ( );
FILL FILL_4_AOI21X1_11 ( );
FILL FILL_5_AOI21X1_11 ( );
FILL FILL_6_AOI21X1_11 ( );
FILL FILL_7_AOI21X1_11 ( );
FILL FILL_8_AOI21X1_11 ( );
FILL FILL_0_NAND2X1_164 ( );
FILL FILL_1_NAND2X1_164 ( );
FILL FILL_2_NAND2X1_164 ( );
FILL FILL_3_NAND2X1_164 ( );
FILL FILL_4_NAND2X1_164 ( );
FILL FILL_5_NAND2X1_164 ( );
FILL FILL_6_NAND2X1_164 ( );
FILL FILL_0_AOI21X1_17 ( );
FILL FILL_1_AOI21X1_17 ( );
FILL FILL_2_AOI21X1_17 ( );
FILL FILL_3_AOI21X1_17 ( );
FILL FILL_4_AOI21X1_17 ( );
FILL FILL_5_AOI21X1_17 ( );
FILL FILL_6_AOI21X1_17 ( );
FILL FILL_7_AOI21X1_17 ( );
FILL FILL_8_AOI21X1_17 ( );
FILL FILL_0_NAND2X1_197 ( );
FILL FILL_1_NAND2X1_197 ( );
FILL FILL_2_NAND2X1_197 ( );
FILL FILL_3_NAND2X1_197 ( );
FILL FILL_4_NAND2X1_197 ( );
FILL FILL_5_NAND2X1_197 ( );
FILL FILL_6_NAND2X1_197 ( );
FILL FILL_0_DFFSR_103 ( );
FILL FILL_1_DFFSR_103 ( );
FILL FILL_2_DFFSR_103 ( );
FILL FILL_3_DFFSR_103 ( );
FILL FILL_4_DFFSR_103 ( );
FILL FILL_5_DFFSR_103 ( );
FILL FILL_6_DFFSR_103 ( );
FILL FILL_7_DFFSR_103 ( );
FILL FILL_8_DFFSR_103 ( );
FILL FILL_9_DFFSR_103 ( );
FILL FILL_10_DFFSR_103 ( );
FILL FILL_11_DFFSR_103 ( );
FILL FILL_12_DFFSR_103 ( );
FILL FILL_13_DFFSR_103 ( );
FILL FILL_14_DFFSR_103 ( );
FILL FILL_15_DFFSR_103 ( );
FILL FILL_16_DFFSR_103 ( );
FILL FILL_17_DFFSR_103 ( );
FILL FILL_18_DFFSR_103 ( );
FILL FILL_19_DFFSR_103 ( );
FILL FILL_20_DFFSR_103 ( );
FILL FILL_21_DFFSR_103 ( );
FILL FILL_22_DFFSR_103 ( );
FILL FILL_23_DFFSR_103 ( );
FILL FILL_24_DFFSR_103 ( );
FILL FILL_25_DFFSR_103 ( );
FILL FILL_26_DFFSR_103 ( );
FILL FILL_27_DFFSR_103 ( );
FILL FILL_28_DFFSR_103 ( );
FILL FILL_29_DFFSR_103 ( );
FILL FILL_30_DFFSR_103 ( );
FILL FILL_31_DFFSR_103 ( );
FILL FILL_32_DFFSR_103 ( );
FILL FILL_33_DFFSR_103 ( );
FILL FILL_34_DFFSR_103 ( );
FILL FILL_35_DFFSR_103 ( );
FILL FILL_36_DFFSR_103 ( );
FILL FILL_37_DFFSR_103 ( );
FILL FILL_38_DFFSR_103 ( );
FILL FILL_39_DFFSR_103 ( );
FILL FILL_40_DFFSR_103 ( );
FILL FILL_41_DFFSR_103 ( );
FILL FILL_42_DFFSR_103 ( );
FILL FILL_43_DFFSR_103 ( );
FILL FILL_44_DFFSR_103 ( );
FILL FILL_45_DFFSR_103 ( );
FILL FILL_46_DFFSR_103 ( );
FILL FILL_47_DFFSR_103 ( );
FILL FILL_48_DFFSR_103 ( );
FILL FILL_49_DFFSR_103 ( );
FILL FILL_50_DFFSR_103 ( );
FILL FILL_51_DFFSR_103 ( );
FILL FILL_0_INVX1_378 ( );
FILL FILL_1_INVX1_378 ( );
FILL FILL_2_INVX1_378 ( );
FILL FILL_3_INVX1_378 ( );
FILL FILL_4_INVX1_378 ( );
FILL FILL_0_OAI22X1_59 ( );
FILL FILL_1_OAI22X1_59 ( );
FILL FILL_2_OAI22X1_59 ( );
FILL FILL_3_OAI22X1_59 ( );
FILL FILL_4_OAI22X1_59 ( );
FILL FILL_5_OAI22X1_59 ( );
FILL FILL_6_OAI22X1_59 ( );
FILL FILL_7_OAI22X1_59 ( );
FILL FILL_8_OAI22X1_59 ( );
FILL FILL_9_OAI22X1_59 ( );
FILL FILL_10_OAI22X1_59 ( );
FILL FILL_11_OAI22X1_59 ( );
FILL FILL_0_INVX1_376 ( );
FILL FILL_1_INVX1_376 ( );
FILL FILL_2_INVX1_376 ( );
FILL FILL_3_INVX1_376 ( );
FILL FILL_4_INVX1_376 ( );
FILL FILL_0_OAI22X1_42 ( );
FILL FILL_1_OAI22X1_42 ( );
FILL FILL_2_OAI22X1_42 ( );
FILL FILL_3_OAI22X1_42 ( );
FILL FILL_4_OAI22X1_42 ( );
FILL FILL_5_OAI22X1_42 ( );
FILL FILL_6_OAI22X1_42 ( );
FILL FILL_7_OAI22X1_42 ( );
FILL FILL_8_OAI22X1_42 ( );
FILL FILL_9_OAI22X1_42 ( );
FILL FILL_10_OAI22X1_42 ( );
FILL FILL_11_OAI22X1_42 ( );
FILL FILL_0_INVX1_342 ( );
FILL FILL_1_INVX1_342 ( );
FILL FILL_2_INVX1_342 ( );
FILL FILL_3_INVX1_342 ( );
FILL FILL_4_INVX1_342 ( );
FILL FILL_0_DFFSR_102 ( );
FILL FILL_1_DFFSR_102 ( );
FILL FILL_2_DFFSR_102 ( );
FILL FILL_3_DFFSR_102 ( );
FILL FILL_4_DFFSR_102 ( );
FILL FILL_5_DFFSR_102 ( );
FILL FILL_6_DFFSR_102 ( );
FILL FILL_7_DFFSR_102 ( );
FILL FILL_8_DFFSR_102 ( );
FILL FILL_9_DFFSR_102 ( );
FILL FILL_10_DFFSR_102 ( );
FILL FILL_11_DFFSR_102 ( );
FILL FILL_12_DFFSR_102 ( );
FILL FILL_13_DFFSR_102 ( );
FILL FILL_14_DFFSR_102 ( );
FILL FILL_15_DFFSR_102 ( );
FILL FILL_16_DFFSR_102 ( );
FILL FILL_17_DFFSR_102 ( );
FILL FILL_18_DFFSR_102 ( );
FILL FILL_19_DFFSR_102 ( );
FILL FILL_20_DFFSR_102 ( );
FILL FILL_21_DFFSR_102 ( );
FILL FILL_22_DFFSR_102 ( );
FILL FILL_23_DFFSR_102 ( );
FILL FILL_24_DFFSR_102 ( );
FILL FILL_25_DFFSR_102 ( );
FILL FILL_26_DFFSR_102 ( );
FILL FILL_27_DFFSR_102 ( );
FILL FILL_28_DFFSR_102 ( );
FILL FILL_29_DFFSR_102 ( );
FILL FILL_30_DFFSR_102 ( );
FILL FILL_31_DFFSR_102 ( );
FILL FILL_32_DFFSR_102 ( );
FILL FILL_33_DFFSR_102 ( );
FILL FILL_34_DFFSR_102 ( );
FILL FILL_35_DFFSR_102 ( );
FILL FILL_36_DFFSR_102 ( );
FILL FILL_37_DFFSR_102 ( );
FILL FILL_38_DFFSR_102 ( );
FILL FILL_39_DFFSR_102 ( );
FILL FILL_40_DFFSR_102 ( );
FILL FILL_41_DFFSR_102 ( );
FILL FILL_42_DFFSR_102 ( );
FILL FILL_43_DFFSR_102 ( );
FILL FILL_44_DFFSR_102 ( );
FILL FILL_45_DFFSR_102 ( );
FILL FILL_46_DFFSR_102 ( );
FILL FILL_47_DFFSR_102 ( );
FILL FILL_48_DFFSR_102 ( );
FILL FILL_49_DFFSR_102 ( );
FILL FILL_50_DFFSR_102 ( );
FILL FILL_0_INVX1_154 ( );
FILL FILL_1_INVX1_154 ( );
FILL FILL_2_INVX1_154 ( );
FILL FILL_3_INVX1_154 ( );
FILL FILL_0_NAND2X1_144 ( );
FILL FILL_1_NAND2X1_144 ( );
FILL FILL_2_NAND2X1_144 ( );
FILL FILL_3_NAND2X1_144 ( );
FILL FILL_4_NAND2X1_144 ( );
FILL FILL_5_NAND2X1_144 ( );
FILL FILL_6_NAND2X1_144 ( );
FILL FILL_0_OAI21X1_144 ( );
FILL FILL_1_OAI21X1_144 ( );
FILL FILL_2_OAI21X1_144 ( );
FILL FILL_3_OAI21X1_144 ( );
FILL FILL_4_OAI21X1_144 ( );
FILL FILL_5_OAI21X1_144 ( );
FILL FILL_6_OAI21X1_144 ( );
FILL FILL_7_OAI21X1_144 ( );
FILL FILL_8_OAI21X1_144 ( );
FILL FILL_0_INVX1_162 ( );
FILL FILL_1_INVX1_162 ( );
FILL FILL_2_INVX1_162 ( );
FILL FILL_3_INVX1_162 ( );
FILL FILL_4_INVX1_162 ( );
FILL FILL_0_XOR2X1_13 ( );
FILL FILL_1_XOR2X1_13 ( );
FILL FILL_2_XOR2X1_13 ( );
FILL FILL_3_XOR2X1_13 ( );
FILL FILL_4_XOR2X1_13 ( );
FILL FILL_5_XOR2X1_13 ( );
FILL FILL_6_XOR2X1_13 ( );
FILL FILL_7_XOR2X1_13 ( );
FILL FILL_8_XOR2X1_13 ( );
FILL FILL_9_XOR2X1_13 ( );
FILL FILL_10_XOR2X1_13 ( );
FILL FILL_11_XOR2X1_13 ( );
FILL FILL_12_XOR2X1_13 ( );
FILL FILL_13_XOR2X1_13 ( );
FILL FILL_14_XOR2X1_13 ( );
FILL FILL_15_XOR2X1_13 ( );
FILL FILL_0_NAND3X1_132 ( );
FILL FILL_1_NAND3X1_132 ( );
FILL FILL_2_NAND3X1_132 ( );
FILL FILL_3_NAND3X1_132 ( );
FILL FILL_4_NAND3X1_132 ( );
FILL FILL_5_NAND3X1_132 ( );
FILL FILL_6_NAND3X1_132 ( );
FILL FILL_7_NAND3X1_132 ( );
FILL FILL_8_NAND3X1_132 ( );
FILL FILL_0_XNOR2X1_4 ( );
FILL FILL_1_XNOR2X1_4 ( );
FILL FILL_2_XNOR2X1_4 ( );
FILL FILL_3_XNOR2X1_4 ( );
FILL FILL_4_XNOR2X1_4 ( );
FILL FILL_5_XNOR2X1_4 ( );
FILL FILL_6_XNOR2X1_4 ( );
FILL FILL_7_XNOR2X1_4 ( );
FILL FILL_8_XNOR2X1_4 ( );
FILL FILL_9_XNOR2X1_4 ( );
FILL FILL_10_XNOR2X1_4 ( );
FILL FILL_11_XNOR2X1_4 ( );
FILL FILL_12_XNOR2X1_4 ( );
FILL FILL_13_XNOR2X1_4 ( );
FILL FILL_14_XNOR2X1_4 ( );
FILL FILL_15_XNOR2X1_4 ( );
FILL FILL_16_XNOR2X1_4 ( );
FILL FILL_0_OAI21X1_40 ( );
FILL FILL_1_OAI21X1_40 ( );
FILL FILL_2_OAI21X1_40 ( );
FILL FILL_3_OAI21X1_40 ( );
FILL FILL_4_OAI21X1_40 ( );
FILL FILL_5_OAI21X1_40 ( );
FILL FILL_6_OAI21X1_40 ( );
FILL FILL_7_OAI21X1_40 ( );
FILL FILL_8_OAI21X1_40 ( );
FILL FILL_9_OAI21X1_40 ( );
FILL FILL_0_INVX1_328 ( );
FILL FILL_1_INVX1_328 ( );
FILL FILL_2_INVX1_328 ( );
FILL FILL_3_INVX1_328 ( );
FILL FILL_4_INVX1_328 ( );
FILL FILL_0_DFFSR_15 ( );
FILL FILL_1_DFFSR_15 ( );
FILL FILL_2_DFFSR_15 ( );
FILL FILL_3_DFFSR_15 ( );
FILL FILL_4_DFFSR_15 ( );
FILL FILL_5_DFFSR_15 ( );
FILL FILL_6_DFFSR_15 ( );
FILL FILL_7_DFFSR_15 ( );
FILL FILL_8_DFFSR_15 ( );
FILL FILL_9_DFFSR_15 ( );
FILL FILL_10_DFFSR_15 ( );
FILL FILL_11_DFFSR_15 ( );
FILL FILL_12_DFFSR_15 ( );
FILL FILL_13_DFFSR_15 ( );
FILL FILL_14_DFFSR_15 ( );
FILL FILL_15_DFFSR_15 ( );
FILL FILL_16_DFFSR_15 ( );
FILL FILL_17_DFFSR_15 ( );
FILL FILL_18_DFFSR_15 ( );
FILL FILL_19_DFFSR_15 ( );
FILL FILL_20_DFFSR_15 ( );
FILL FILL_21_DFFSR_15 ( );
FILL FILL_22_DFFSR_15 ( );
FILL FILL_23_DFFSR_15 ( );
FILL FILL_24_DFFSR_15 ( );
FILL FILL_25_DFFSR_15 ( );
FILL FILL_26_DFFSR_15 ( );
FILL FILL_27_DFFSR_15 ( );
FILL FILL_28_DFFSR_15 ( );
FILL FILL_29_DFFSR_15 ( );
FILL FILL_30_DFFSR_15 ( );
FILL FILL_31_DFFSR_15 ( );
FILL FILL_32_DFFSR_15 ( );
FILL FILL_33_DFFSR_15 ( );
FILL FILL_34_DFFSR_15 ( );
FILL FILL_35_DFFSR_15 ( );
FILL FILL_36_DFFSR_15 ( );
FILL FILL_37_DFFSR_15 ( );
FILL FILL_38_DFFSR_15 ( );
FILL FILL_39_DFFSR_15 ( );
FILL FILL_40_DFFSR_15 ( );
FILL FILL_41_DFFSR_15 ( );
FILL FILL_42_DFFSR_15 ( );
FILL FILL_43_DFFSR_15 ( );
FILL FILL_44_DFFSR_15 ( );
FILL FILL_45_DFFSR_15 ( );
FILL FILL_46_DFFSR_15 ( );
FILL FILL_47_DFFSR_15 ( );
FILL FILL_48_DFFSR_15 ( );
FILL FILL_49_DFFSR_15 ( );
FILL FILL_50_DFFSR_15 ( );
FILL FILL_51_DFFSR_15 ( );
FILL FILL_0_INVX1_268 ( );
FILL FILL_1_INVX1_268 ( );
FILL FILL_2_INVX1_268 ( );
FILL FILL_3_INVX1_268 ( );
FILL FILL_4_INVX1_268 ( );
FILL FILL_0_OAI21X1_41 ( );
FILL FILL_1_OAI21X1_41 ( );
FILL FILL_2_OAI21X1_41 ( );
FILL FILL_3_OAI21X1_41 ( );
FILL FILL_4_OAI21X1_41 ( );
FILL FILL_5_OAI21X1_41 ( );
FILL FILL_6_OAI21X1_41 ( );
FILL FILL_7_OAI21X1_41 ( );
FILL FILL_8_OAI21X1_41 ( );
FILL FILL_0_INVX1_302 ( );
FILL FILL_1_INVX1_302 ( );
FILL FILL_2_INVX1_302 ( );
FILL FILL_3_INVX1_302 ( );
FILL FILL_4_INVX1_302 ( );
FILL FILL_0_NAND2X1_17 ( );
FILL FILL_1_NAND2X1_17 ( );
FILL FILL_2_NAND2X1_17 ( );
FILL FILL_3_NAND2X1_17 ( );
FILL FILL_4_NAND2X1_17 ( );
FILL FILL_5_NAND2X1_17 ( );
FILL FILL_6_NAND2X1_17 ( );
FILL FILL_0_DFFSR_7 ( );
FILL FILL_1_DFFSR_7 ( );
FILL FILL_2_DFFSR_7 ( );
FILL FILL_3_DFFSR_7 ( );
FILL FILL_4_DFFSR_7 ( );
FILL FILL_5_DFFSR_7 ( );
FILL FILL_6_DFFSR_7 ( );
FILL FILL_7_DFFSR_7 ( );
FILL FILL_8_DFFSR_7 ( );
FILL FILL_9_DFFSR_7 ( );
FILL FILL_10_DFFSR_7 ( );
FILL FILL_11_DFFSR_7 ( );
FILL FILL_12_DFFSR_7 ( );
FILL FILL_13_DFFSR_7 ( );
FILL FILL_14_DFFSR_7 ( );
FILL FILL_15_DFFSR_7 ( );
FILL FILL_16_DFFSR_7 ( );
FILL FILL_17_DFFSR_7 ( );
FILL FILL_18_DFFSR_7 ( );
FILL FILL_19_DFFSR_7 ( );
FILL FILL_20_DFFSR_7 ( );
FILL FILL_21_DFFSR_7 ( );
FILL FILL_22_DFFSR_7 ( );
FILL FILL_23_DFFSR_7 ( );
FILL FILL_24_DFFSR_7 ( );
FILL FILL_25_DFFSR_7 ( );
FILL FILL_26_DFFSR_7 ( );
FILL FILL_27_DFFSR_7 ( );
FILL FILL_28_DFFSR_7 ( );
FILL FILL_29_DFFSR_7 ( );
FILL FILL_30_DFFSR_7 ( );
FILL FILL_31_DFFSR_7 ( );
FILL FILL_32_DFFSR_7 ( );
FILL FILL_33_DFFSR_7 ( );
FILL FILL_34_DFFSR_7 ( );
FILL FILL_35_DFFSR_7 ( );
FILL FILL_36_DFFSR_7 ( );
FILL FILL_37_DFFSR_7 ( );
FILL FILL_38_DFFSR_7 ( );
FILL FILL_39_DFFSR_7 ( );
FILL FILL_40_DFFSR_7 ( );
FILL FILL_41_DFFSR_7 ( );
FILL FILL_42_DFFSR_7 ( );
FILL FILL_43_DFFSR_7 ( );
FILL FILL_44_DFFSR_7 ( );
FILL FILL_45_DFFSR_7 ( );
FILL FILL_46_DFFSR_7 ( );
FILL FILL_47_DFFSR_7 ( );
FILL FILL_48_DFFSR_7 ( );
FILL FILL_49_DFFSR_7 ( );
FILL FILL_50_DFFSR_7 ( );
FILL FILL_0_NAND2X1_183 ( );
FILL FILL_1_NAND2X1_183 ( );
FILL FILL_2_NAND2X1_183 ( );
FILL FILL_3_NAND2X1_183 ( );
FILL FILL_4_NAND2X1_183 ( );
FILL FILL_5_NAND2X1_183 ( );
FILL FILL_6_NAND2X1_183 ( );
FILL FILL_0_NAND3X1_6 ( );
FILL FILL_1_NAND3X1_6 ( );
FILL FILL_2_NAND3X1_6 ( );
FILL FILL_3_NAND3X1_6 ( );
FILL FILL_4_NAND3X1_6 ( );
FILL FILL_5_NAND3X1_6 ( );
FILL FILL_6_NAND3X1_6 ( );
FILL FILL_7_NAND3X1_6 ( );
FILL FILL_8_NAND3X1_6 ( );
FILL FILL_0_NAND2X1_5 ( );
FILL FILL_1_NAND2X1_5 ( );
FILL FILL_2_NAND2X1_5 ( );
FILL FILL_3_NAND2X1_5 ( );
FILL FILL_4_NAND2X1_5 ( );
FILL FILL_5_NAND2X1_5 ( );
FILL FILL_6_NAND2X1_5 ( );
FILL FILL_0_NAND2X1_188 ( );
FILL FILL_1_NAND2X1_188 ( );
FILL FILL_2_NAND2X1_188 ( );
FILL FILL_3_NAND2X1_188 ( );
FILL FILL_4_NAND2X1_188 ( );
FILL FILL_5_NAND2X1_188 ( );
FILL FILL_6_NAND2X1_188 ( );
FILL FILL_0_OAI21X1_197 ( );
FILL FILL_1_OAI21X1_197 ( );
FILL FILL_2_OAI21X1_197 ( );
FILL FILL_3_OAI21X1_197 ( );
FILL FILL_4_OAI21X1_197 ( );
FILL FILL_5_OAI21X1_197 ( );
FILL FILL_6_OAI21X1_197 ( );
FILL FILL_7_OAI21X1_197 ( );
FILL FILL_8_OAI21X1_197 ( );
FILL FILL_0_INVX1_236 ( );
FILL FILL_1_INVX1_236 ( );
FILL FILL_2_INVX1_236 ( );
FILL FILL_3_INVX1_236 ( );
FILL FILL_0_AOI21X1_12 ( );
FILL FILL_1_AOI21X1_12 ( );
FILL FILL_2_AOI21X1_12 ( );
FILL FILL_3_AOI21X1_12 ( );
FILL FILL_4_AOI21X1_12 ( );
FILL FILL_5_AOI21X1_12 ( );
FILL FILL_6_AOI21X1_12 ( );
FILL FILL_7_AOI21X1_12 ( );
FILL FILL_8_AOI21X1_12 ( );
FILL FILL_9_AOI21X1_12 ( );
FILL FILL_0_AOI21X1_13 ( );
FILL FILL_1_AOI21X1_13 ( );
FILL FILL_2_AOI21X1_13 ( );
FILL FILL_3_AOI21X1_13 ( );
FILL FILL_4_AOI21X1_13 ( );
FILL FILL_5_AOI21X1_13 ( );
FILL FILL_6_AOI21X1_13 ( );
FILL FILL_7_AOI21X1_13 ( );
FILL FILL_8_AOI21X1_13 ( );
FILL FILL_9_AOI21X1_13 ( );
FILL FILL_0_OAI21X1_198 ( );
FILL FILL_1_OAI21X1_198 ( );
FILL FILL_2_OAI21X1_198 ( );
FILL FILL_3_OAI21X1_198 ( );
FILL FILL_4_OAI21X1_198 ( );
FILL FILL_5_OAI21X1_198 ( );
FILL FILL_6_OAI21X1_198 ( );
FILL FILL_7_OAI21X1_198 ( );
FILL FILL_8_OAI21X1_198 ( );
FILL FILL_0_INVX1_237 ( );
FILL FILL_1_INVX1_237 ( );
FILL FILL_2_INVX1_237 ( );
FILL FILL_3_INVX1_237 ( );
FILL FILL_0_NAND3X1_33 ( );
FILL FILL_1_NAND3X1_33 ( );
FILL FILL_2_NAND3X1_33 ( );
FILL FILL_3_NAND3X1_33 ( );
FILL FILL_4_NAND3X1_33 ( );
FILL FILL_5_NAND3X1_33 ( );
FILL FILL_6_NAND3X1_33 ( );
FILL FILL_7_NAND3X1_33 ( );
FILL FILL_8_NAND3X1_33 ( );
FILL FILL_9_NAND3X1_33 ( );
FILL FILL_0_NAND2X1_101 ( );
FILL FILL_1_NAND2X1_101 ( );
FILL FILL_2_NAND2X1_101 ( );
FILL FILL_3_NAND2X1_101 ( );
FILL FILL_4_NAND2X1_101 ( );
FILL FILL_5_NAND2X1_101 ( );
FILL FILL_6_NAND2X1_101 ( );
FILL FILL_0_OAI21X1_101 ( );
FILL FILL_1_OAI21X1_101 ( );
FILL FILL_2_OAI21X1_101 ( );
FILL FILL_3_OAI21X1_101 ( );
FILL FILL_4_OAI21X1_101 ( );
FILL FILL_5_OAI21X1_101 ( );
FILL FILL_6_OAI21X1_101 ( );
FILL FILL_7_OAI21X1_101 ( );
FILL FILL_8_OAI21X1_101 ( );
FILL FILL_9_OAI21X1_101 ( );
FILL FILL_0_INVX1_114 ( );
FILL FILL_1_INVX1_114 ( );
FILL FILL_2_INVX1_114 ( );
FILL FILL_3_INVX1_114 ( );
FILL FILL_0_INVX1_390 ( );
FILL FILL_1_INVX1_390 ( );
FILL FILL_2_INVX1_390 ( );
FILL FILL_3_INVX1_390 ( );
FILL FILL_4_INVX1_390 ( );
FILL FILL_0_INVX1_391 ( );
FILL FILL_1_INVX1_391 ( );
FILL FILL_2_INVX1_391 ( );
FILL FILL_3_INVX1_391 ( );
FILL FILL_0_OAI22X1_66 ( );
FILL FILL_1_OAI22X1_66 ( );
FILL FILL_2_OAI22X1_66 ( );
FILL FILL_3_OAI22X1_66 ( );
FILL FILL_4_OAI22X1_66 ( );
FILL FILL_5_OAI22X1_66 ( );
FILL FILL_6_OAI22X1_66 ( );
FILL FILL_7_OAI22X1_66 ( );
FILL FILL_8_OAI22X1_66 ( );
FILL FILL_9_OAI22X1_66 ( );
FILL FILL_10_OAI22X1_66 ( );
FILL FILL_11_OAI22X1_66 ( );
FILL FILL_0_INVX1_142 ( );
FILL FILL_1_INVX1_142 ( );
FILL FILL_2_INVX1_142 ( );
FILL FILL_3_INVX1_142 ( );
FILL FILL_4_INVX1_142 ( );
FILL FILL_0_OAI21X1_126 ( );
FILL FILL_1_OAI21X1_126 ( );
FILL FILL_2_OAI21X1_126 ( );
FILL FILL_3_OAI21X1_126 ( );
FILL FILL_4_OAI21X1_126 ( );
FILL FILL_5_OAI21X1_126 ( );
FILL FILL_6_OAI21X1_126 ( );
FILL FILL_7_OAI21X1_126 ( );
FILL FILL_8_OAI21X1_126 ( );
FILL FILL_0_NAND2X1_126 ( );
FILL FILL_1_NAND2X1_126 ( );
FILL FILL_2_NAND2X1_126 ( );
FILL FILL_3_NAND2X1_126 ( );
FILL FILL_4_NAND2X1_126 ( );
FILL FILL_5_NAND2X1_126 ( );
FILL FILL_6_NAND2X1_126 ( );
FILL FILL_0_NOR2X1_43 ( );
FILL FILL_1_NOR2X1_43 ( );
FILL FILL_2_NOR2X1_43 ( );
FILL FILL_3_NOR2X1_43 ( );
FILL FILL_4_NOR2X1_43 ( );
FILL FILL_5_NOR2X1_43 ( );
FILL FILL_6_NOR2X1_43 ( );
FILL FILL_0_NOR2X1_38 ( );
FILL FILL_1_NOR2X1_38 ( );
FILL FILL_2_NOR2X1_38 ( );
FILL FILL_3_NOR2X1_38 ( );
FILL FILL_4_NOR2X1_38 ( );
FILL FILL_5_NOR2X1_38 ( );
FILL FILL_6_NOR2X1_38 ( );
FILL FILL_0_NAND2X1_249 ( );
FILL FILL_1_NAND2X1_249 ( );
FILL FILL_2_NAND2X1_249 ( );
FILL FILL_3_NAND2X1_249 ( );
FILL FILL_4_NAND2X1_249 ( );
FILL FILL_5_NAND2X1_249 ( );
FILL FILL_6_NAND2X1_249 ( );
FILL FILL_0_INVX1_374 ( );
FILL FILL_1_INVX1_374 ( );
FILL FILL_2_INVX1_374 ( );
FILL FILL_3_INVX1_374 ( );
FILL FILL_4_INVX1_374 ( );
FILL FILL_0_OAI22X1_58 ( );
FILL FILL_1_OAI22X1_58 ( );
FILL FILL_2_OAI22X1_58 ( );
FILL FILL_3_OAI22X1_58 ( );
FILL FILL_4_OAI22X1_58 ( );
FILL FILL_5_OAI22X1_58 ( );
FILL FILL_6_OAI22X1_58 ( );
FILL FILL_7_OAI22X1_58 ( );
FILL FILL_8_OAI22X1_58 ( );
FILL FILL_9_OAI22X1_58 ( );
FILL FILL_10_OAI22X1_58 ( );
FILL FILL_11_OAI22X1_58 ( );
FILL FILL_0_DFFSR_72 ( );
FILL FILL_1_DFFSR_72 ( );
FILL FILL_2_DFFSR_72 ( );
FILL FILL_3_DFFSR_72 ( );
FILL FILL_4_DFFSR_72 ( );
FILL FILL_5_DFFSR_72 ( );
FILL FILL_6_DFFSR_72 ( );
FILL FILL_7_DFFSR_72 ( );
FILL FILL_8_DFFSR_72 ( );
FILL FILL_9_DFFSR_72 ( );
FILL FILL_10_DFFSR_72 ( );
FILL FILL_11_DFFSR_72 ( );
FILL FILL_12_DFFSR_72 ( );
FILL FILL_13_DFFSR_72 ( );
FILL FILL_14_DFFSR_72 ( );
FILL FILL_15_DFFSR_72 ( );
FILL FILL_16_DFFSR_72 ( );
FILL FILL_17_DFFSR_72 ( );
FILL FILL_18_DFFSR_72 ( );
FILL FILL_19_DFFSR_72 ( );
FILL FILL_20_DFFSR_72 ( );
FILL FILL_21_DFFSR_72 ( );
FILL FILL_22_DFFSR_72 ( );
FILL FILL_23_DFFSR_72 ( );
FILL FILL_24_DFFSR_72 ( );
FILL FILL_25_DFFSR_72 ( );
FILL FILL_26_DFFSR_72 ( );
FILL FILL_27_DFFSR_72 ( );
FILL FILL_28_DFFSR_72 ( );
FILL FILL_29_DFFSR_72 ( );
FILL FILL_30_DFFSR_72 ( );
FILL FILL_31_DFFSR_72 ( );
FILL FILL_32_DFFSR_72 ( );
FILL FILL_33_DFFSR_72 ( );
FILL FILL_34_DFFSR_72 ( );
FILL FILL_35_DFFSR_72 ( );
FILL FILL_36_DFFSR_72 ( );
FILL FILL_37_DFFSR_72 ( );
FILL FILL_38_DFFSR_72 ( );
FILL FILL_39_DFFSR_72 ( );
FILL FILL_40_DFFSR_72 ( );
FILL FILL_41_DFFSR_72 ( );
FILL FILL_42_DFFSR_72 ( );
FILL FILL_43_DFFSR_72 ( );
FILL FILL_44_DFFSR_72 ( );
FILL FILL_45_DFFSR_72 ( );
FILL FILL_46_DFFSR_72 ( );
FILL FILL_47_DFFSR_72 ( );
FILL FILL_48_DFFSR_72 ( );
FILL FILL_49_DFFSR_72 ( );
FILL FILL_50_DFFSR_72 ( );
FILL FILL_0_CLKBUF1_9 ( );
FILL FILL_1_CLKBUF1_9 ( );
FILL FILL_2_CLKBUF1_9 ( );
FILL FILL_3_CLKBUF1_9 ( );
FILL FILL_4_CLKBUF1_9 ( );
FILL FILL_5_CLKBUF1_9 ( );
FILL FILL_6_CLKBUF1_9 ( );
FILL FILL_7_CLKBUF1_9 ( );
FILL FILL_8_CLKBUF1_9 ( );
FILL FILL_9_CLKBUF1_9 ( );
FILL FILL_10_CLKBUF1_9 ( );
FILL FILL_11_CLKBUF1_9 ( );
FILL FILL_12_CLKBUF1_9 ( );
FILL FILL_13_CLKBUF1_9 ( );
FILL FILL_14_CLKBUF1_9 ( );
FILL FILL_15_CLKBUF1_9 ( );
FILL FILL_16_CLKBUF1_9 ( );
FILL FILL_17_CLKBUF1_9 ( );
FILL FILL_18_CLKBUF1_9 ( );
FILL FILL_19_CLKBUF1_9 ( );
FILL FILL_20_CLKBUF1_9 ( );
FILL FILL_0_AOI21X1_44 ( );
FILL FILL_1_AOI21X1_44 ( );
FILL FILL_2_AOI21X1_44 ( );
FILL FILL_3_AOI21X1_44 ( );
FILL FILL_4_AOI21X1_44 ( );
FILL FILL_5_AOI21X1_44 ( );
FILL FILL_6_AOI21X1_44 ( );
FILL FILL_7_AOI21X1_44 ( );
FILL FILL_8_AOI21X1_44 ( );
FILL FILL_9_AOI21X1_44 ( );
FILL FILL_0_AOI21X1_43 ( );
FILL FILL_1_AOI21X1_43 ( );
FILL FILL_2_AOI21X1_43 ( );
FILL FILL_3_AOI21X1_43 ( );
FILL FILL_4_AOI21X1_43 ( );
FILL FILL_5_AOI21X1_43 ( );
FILL FILL_6_AOI21X1_43 ( );
FILL FILL_7_AOI21X1_43 ( );
FILL FILL_8_AOI21X1_43 ( );
FILL FILL_0_XOR2X1_12 ( );
FILL FILL_1_XOR2X1_12 ( );
FILL FILL_2_XOR2X1_12 ( );
FILL FILL_3_XOR2X1_12 ( );
FILL FILL_4_XOR2X1_12 ( );
FILL FILL_5_XOR2X1_12 ( );
FILL FILL_6_XOR2X1_12 ( );
FILL FILL_7_XOR2X1_12 ( );
FILL FILL_8_XOR2X1_12 ( );
FILL FILL_9_XOR2X1_12 ( );
FILL FILL_10_XOR2X1_12 ( );
FILL FILL_11_XOR2X1_12 ( );
FILL FILL_12_XOR2X1_12 ( );
FILL FILL_13_XOR2X1_12 ( );
FILL FILL_14_XOR2X1_12 ( );
FILL FILL_15_XOR2X1_12 ( );
FILL FILL_0_INVX1_325 ( );
FILL FILL_1_INVX1_325 ( );
FILL FILL_2_INVX1_325 ( );
FILL FILL_3_INVX1_325 ( );
FILL FILL_4_INVX1_325 ( );
FILL FILL_0_INVX1_322 ( );
FILL FILL_1_INVX1_322 ( );
FILL FILL_2_INVX1_322 ( );
FILL FILL_3_INVX1_322 ( );
FILL FILL_4_INVX1_322 ( );
FILL FILL_0_INVX1_326 ( );
FILL FILL_1_INVX1_326 ( );
FILL FILL_2_INVX1_326 ( );
FILL FILL_3_INVX1_326 ( );
FILL FILL_4_INVX1_326 ( );
FILL FILL_0_OAI22X1_35 ( );
FILL FILL_1_OAI22X1_35 ( );
FILL FILL_2_OAI22X1_35 ( );
FILL FILL_3_OAI22X1_35 ( );
FILL FILL_4_OAI22X1_35 ( );
FILL FILL_5_OAI22X1_35 ( );
FILL FILL_6_OAI22X1_35 ( );
FILL FILL_7_OAI22X1_35 ( );
FILL FILL_8_OAI22X1_35 ( );
FILL FILL_9_OAI22X1_35 ( );
FILL FILL_10_OAI22X1_35 ( );
FILL FILL_0_NAND2X1_50 ( );
FILL FILL_1_NAND2X1_50 ( );
FILL FILL_2_NAND2X1_50 ( );
FILL FILL_3_NAND2X1_50 ( );
FILL FILL_4_NAND2X1_50 ( );
FILL FILL_5_NAND2X1_50 ( );
FILL FILL_6_NAND2X1_50 ( );
FILL FILL_0_OAI21X1_50 ( );
FILL FILL_1_OAI21X1_50 ( );
FILL FILL_2_OAI21X1_50 ( );
FILL FILL_3_OAI21X1_50 ( );
FILL FILL_4_OAI21X1_50 ( );
FILL FILL_5_OAI21X1_50 ( );
FILL FILL_6_OAI21X1_50 ( );
FILL FILL_7_OAI21X1_50 ( );
FILL FILL_8_OAI21X1_50 ( );
FILL FILL_9_OAI21X1_50 ( );
FILL FILL_0_INVX1_17 ( );
FILL FILL_1_INVX1_17 ( );
FILL FILL_2_INVX1_17 ( );
FILL FILL_3_INVX1_17 ( );
FILL FILL_0_NAND2X1_15 ( );
FILL FILL_1_NAND2X1_15 ( );
FILL FILL_2_NAND2X1_15 ( );
FILL FILL_3_NAND2X1_15 ( );
FILL FILL_4_NAND2X1_15 ( );
FILL FILL_5_NAND2X1_15 ( );
FILL FILL_6_NAND2X1_15 ( );
FILL FILL_0_CLKBUF1_21 ( );
FILL FILL_1_CLKBUF1_21 ( );
FILL FILL_2_CLKBUF1_21 ( );
FILL FILL_3_CLKBUF1_21 ( );
FILL FILL_4_CLKBUF1_21 ( );
FILL FILL_5_CLKBUF1_21 ( );
FILL FILL_6_CLKBUF1_21 ( );
FILL FILL_7_CLKBUF1_21 ( );
FILL FILL_8_CLKBUF1_21 ( );
FILL FILL_9_CLKBUF1_21 ( );
FILL FILL_10_CLKBUF1_21 ( );
FILL FILL_11_CLKBUF1_21 ( );
FILL FILL_12_CLKBUF1_21 ( );
FILL FILL_13_CLKBUF1_21 ( );
FILL FILL_14_CLKBUF1_21 ( );
FILL FILL_15_CLKBUF1_21 ( );
FILL FILL_16_CLKBUF1_21 ( );
FILL FILL_17_CLKBUF1_21 ( );
FILL FILL_18_CLKBUF1_21 ( );
FILL FILL_19_CLKBUF1_21 ( );
FILL FILL_20_CLKBUF1_21 ( );
FILL FILL_0_NAND2X1_35 ( );
FILL FILL_1_NAND2X1_35 ( );
FILL FILL_2_NAND2X1_35 ( );
FILL FILL_3_NAND2X1_35 ( );
FILL FILL_4_NAND2X1_35 ( );
FILL FILL_5_NAND2X1_35 ( );
FILL FILL_6_NAND2X1_35 ( );
FILL FILL_0_INVX1_47 ( );
FILL FILL_1_INVX1_47 ( );
FILL FILL_2_INVX1_47 ( );
FILL FILL_3_INVX1_47 ( );
FILL FILL_4_INVX1_47 ( );
FILL FILL_0_CLKBUF1_15 ( );
FILL FILL_1_CLKBUF1_15 ( );
FILL FILL_2_CLKBUF1_15 ( );
FILL FILL_3_CLKBUF1_15 ( );
FILL FILL_4_CLKBUF1_15 ( );
FILL FILL_5_CLKBUF1_15 ( );
FILL FILL_6_CLKBUF1_15 ( );
FILL FILL_7_CLKBUF1_15 ( );
FILL FILL_8_CLKBUF1_15 ( );
FILL FILL_9_CLKBUF1_15 ( );
FILL FILL_10_CLKBUF1_15 ( );
FILL FILL_11_CLKBUF1_15 ( );
FILL FILL_12_CLKBUF1_15 ( );
FILL FILL_13_CLKBUF1_15 ( );
FILL FILL_14_CLKBUF1_15 ( );
FILL FILL_15_CLKBUF1_15 ( );
FILL FILL_16_CLKBUF1_15 ( );
FILL FILL_17_CLKBUF1_15 ( );
FILL FILL_18_CLKBUF1_15 ( );
FILL FILL_19_CLKBUF1_15 ( );
FILL FILL_20_CLKBUF1_15 ( );
FILL FILL_0_DFFPOSX1_4 ( );
FILL FILL_1_DFFPOSX1_4 ( );
FILL FILL_2_DFFPOSX1_4 ( );
FILL FILL_3_DFFPOSX1_4 ( );
FILL FILL_4_DFFPOSX1_4 ( );
FILL FILL_5_DFFPOSX1_4 ( );
FILL FILL_6_DFFPOSX1_4 ( );
FILL FILL_7_DFFPOSX1_4 ( );
FILL FILL_8_DFFPOSX1_4 ( );
FILL FILL_9_DFFPOSX1_4 ( );
FILL FILL_10_DFFPOSX1_4 ( );
FILL FILL_11_DFFPOSX1_4 ( );
FILL FILL_12_DFFPOSX1_4 ( );
FILL FILL_13_DFFPOSX1_4 ( );
FILL FILL_14_DFFPOSX1_4 ( );
FILL FILL_15_DFFPOSX1_4 ( );
FILL FILL_16_DFFPOSX1_4 ( );
FILL FILL_17_DFFPOSX1_4 ( );
FILL FILL_18_DFFPOSX1_4 ( );
FILL FILL_19_DFFPOSX1_4 ( );
FILL FILL_20_DFFPOSX1_4 ( );
FILL FILL_21_DFFPOSX1_4 ( );
FILL FILL_22_DFFPOSX1_4 ( );
FILL FILL_23_DFFPOSX1_4 ( );
FILL FILL_24_DFFPOSX1_4 ( );
FILL FILL_25_DFFPOSX1_4 ( );
FILL FILL_26_DFFPOSX1_4 ( );
FILL FILL_27_DFFPOSX1_4 ( );
FILL FILL_0_OAI21X1_182 ( );
FILL FILL_1_OAI21X1_182 ( );
FILL FILL_2_OAI21X1_182 ( );
FILL FILL_3_OAI21X1_182 ( );
FILL FILL_4_OAI21X1_182 ( );
FILL FILL_5_OAI21X1_182 ( );
FILL FILL_6_OAI21X1_182 ( );
FILL FILL_7_OAI21X1_182 ( );
FILL FILL_8_OAI21X1_182 ( );
FILL FILL_0_INVX1_222 ( );
FILL FILL_1_INVX1_222 ( );
FILL FILL_2_INVX1_222 ( );
FILL FILL_3_INVX1_222 ( );
FILL FILL_4_INVX1_222 ( );
FILL FILL_0_OAI21X1_183 ( );
FILL FILL_1_OAI21X1_183 ( );
FILL FILL_2_OAI21X1_183 ( );
FILL FILL_3_OAI21X1_183 ( );
FILL FILL_4_OAI21X1_183 ( );
FILL FILL_5_OAI21X1_183 ( );
FILL FILL_6_OAI21X1_183 ( );
FILL FILL_7_OAI21X1_183 ( );
FILL FILL_8_OAI21X1_183 ( );
FILL FILL_0_INVX1_221 ( );
FILL FILL_1_INVX1_221 ( );
FILL FILL_2_INVX1_221 ( );
FILL FILL_3_INVX1_221 ( );
FILL FILL_4_INVX1_221 ( );
FILL FILL_0_XOR2X1_3 ( );
FILL FILL_1_XOR2X1_3 ( );
FILL FILL_2_XOR2X1_3 ( );
FILL FILL_3_XOR2X1_3 ( );
FILL FILL_4_XOR2X1_3 ( );
FILL FILL_5_XOR2X1_3 ( );
FILL FILL_6_XOR2X1_3 ( );
FILL FILL_7_XOR2X1_3 ( );
FILL FILL_8_XOR2X1_3 ( );
FILL FILL_9_XOR2X1_3 ( );
FILL FILL_10_XOR2X1_3 ( );
FILL FILL_11_XOR2X1_3 ( );
FILL FILL_12_XOR2X1_3 ( );
FILL FILL_13_XOR2X1_3 ( );
FILL FILL_14_XOR2X1_3 ( );
FILL FILL_15_XOR2X1_3 ( );
FILL FILL_0_DFFSR_180 ( );
FILL FILL_1_DFFSR_180 ( );
FILL FILL_2_DFFSR_180 ( );
FILL FILL_3_DFFSR_180 ( );
FILL FILL_4_DFFSR_180 ( );
FILL FILL_5_DFFSR_180 ( );
FILL FILL_6_DFFSR_180 ( );
FILL FILL_7_DFFSR_180 ( );
FILL FILL_8_DFFSR_180 ( );
FILL FILL_9_DFFSR_180 ( );
FILL FILL_10_DFFSR_180 ( );
FILL FILL_11_DFFSR_180 ( );
FILL FILL_12_DFFSR_180 ( );
FILL FILL_13_DFFSR_180 ( );
FILL FILL_14_DFFSR_180 ( );
FILL FILL_15_DFFSR_180 ( );
FILL FILL_16_DFFSR_180 ( );
FILL FILL_17_DFFSR_180 ( );
FILL FILL_18_DFFSR_180 ( );
FILL FILL_19_DFFSR_180 ( );
FILL FILL_20_DFFSR_180 ( );
FILL FILL_21_DFFSR_180 ( );
FILL FILL_22_DFFSR_180 ( );
FILL FILL_23_DFFSR_180 ( );
FILL FILL_24_DFFSR_180 ( );
FILL FILL_25_DFFSR_180 ( );
FILL FILL_26_DFFSR_180 ( );
FILL FILL_27_DFFSR_180 ( );
FILL FILL_28_DFFSR_180 ( );
FILL FILL_29_DFFSR_180 ( );
FILL FILL_30_DFFSR_180 ( );
FILL FILL_31_DFFSR_180 ( );
FILL FILL_32_DFFSR_180 ( );
FILL FILL_33_DFFSR_180 ( );
FILL FILL_34_DFFSR_180 ( );
FILL FILL_35_DFFSR_180 ( );
FILL FILL_36_DFFSR_180 ( );
FILL FILL_37_DFFSR_180 ( );
FILL FILL_38_DFFSR_180 ( );
FILL FILL_39_DFFSR_180 ( );
FILL FILL_40_DFFSR_180 ( );
FILL FILL_41_DFFSR_180 ( );
FILL FILL_42_DFFSR_180 ( );
FILL FILL_43_DFFSR_180 ( );
FILL FILL_44_DFFSR_180 ( );
FILL FILL_45_DFFSR_180 ( );
FILL FILL_46_DFFSR_180 ( );
FILL FILL_47_DFFSR_180 ( );
FILL FILL_48_DFFSR_180 ( );
FILL FILL_49_DFFSR_180 ( );
FILL FILL_50_DFFSR_180 ( );
FILL FILL_0_DFFSR_126 ( );
FILL FILL_1_DFFSR_126 ( );
FILL FILL_2_DFFSR_126 ( );
FILL FILL_3_DFFSR_126 ( );
FILL FILL_4_DFFSR_126 ( );
FILL FILL_5_DFFSR_126 ( );
FILL FILL_6_DFFSR_126 ( );
FILL FILL_7_DFFSR_126 ( );
FILL FILL_8_DFFSR_126 ( );
FILL FILL_9_DFFSR_126 ( );
FILL FILL_10_DFFSR_126 ( );
FILL FILL_11_DFFSR_126 ( );
FILL FILL_12_DFFSR_126 ( );
FILL FILL_13_DFFSR_126 ( );
FILL FILL_14_DFFSR_126 ( );
FILL FILL_15_DFFSR_126 ( );
FILL FILL_16_DFFSR_126 ( );
FILL FILL_17_DFFSR_126 ( );
FILL FILL_18_DFFSR_126 ( );
FILL FILL_19_DFFSR_126 ( );
FILL FILL_20_DFFSR_126 ( );
FILL FILL_21_DFFSR_126 ( );
FILL FILL_22_DFFSR_126 ( );
FILL FILL_23_DFFSR_126 ( );
FILL FILL_24_DFFSR_126 ( );
FILL FILL_25_DFFSR_126 ( );
FILL FILL_26_DFFSR_126 ( );
FILL FILL_27_DFFSR_126 ( );
FILL FILL_28_DFFSR_126 ( );
FILL FILL_29_DFFSR_126 ( );
FILL FILL_30_DFFSR_126 ( );
FILL FILL_31_DFFSR_126 ( );
FILL FILL_32_DFFSR_126 ( );
FILL FILL_33_DFFSR_126 ( );
FILL FILL_34_DFFSR_126 ( );
FILL FILL_35_DFFSR_126 ( );
FILL FILL_36_DFFSR_126 ( );
FILL FILL_37_DFFSR_126 ( );
FILL FILL_38_DFFSR_126 ( );
FILL FILL_39_DFFSR_126 ( );
FILL FILL_40_DFFSR_126 ( );
FILL FILL_41_DFFSR_126 ( );
FILL FILL_42_DFFSR_126 ( );
FILL FILL_43_DFFSR_126 ( );
FILL FILL_44_DFFSR_126 ( );
FILL FILL_45_DFFSR_126 ( );
FILL FILL_46_DFFSR_126 ( );
FILL FILL_47_DFFSR_126 ( );
FILL FILL_48_DFFSR_126 ( );
FILL FILL_49_DFFSR_126 ( );
FILL FILL_50_DFFSR_126 ( );
FILL FILL_0_OAI22X1_57 ( );
FILL FILL_1_OAI22X1_57 ( );
FILL FILL_2_OAI22X1_57 ( );
FILL FILL_3_OAI22X1_57 ( );
FILL FILL_4_OAI22X1_57 ( );
FILL FILL_5_OAI22X1_57 ( );
FILL FILL_6_OAI22X1_57 ( );
FILL FILL_7_OAI22X1_57 ( );
FILL FILL_8_OAI22X1_57 ( );
FILL FILL_9_OAI22X1_57 ( );
FILL FILL_10_OAI22X1_57 ( );
FILL FILL_11_OAI22X1_57 ( );
FILL FILL_0_INVX1_379 ( );
FILL FILL_1_INVX1_379 ( );
FILL FILL_2_INVX1_379 ( );
FILL FILL_3_INVX1_379 ( );
FILL FILL_0_BUFX2_17 ( );
FILL FILL_1_BUFX2_17 ( );
FILL FILL_2_BUFX2_17 ( );
FILL FILL_3_BUFX2_17 ( );
FILL FILL_4_BUFX2_17 ( );
FILL FILL_5_BUFX2_17 ( );
FILL FILL_6_BUFX2_17 ( );
FILL FILL_0_NOR2X1_42 ( );
FILL FILL_1_NOR2X1_42 ( );
FILL FILL_2_NOR2X1_42 ( );
FILL FILL_3_NOR2X1_42 ( );
FILL FILL_4_NOR2X1_42 ( );
FILL FILL_5_NOR2X1_42 ( );
FILL FILL_6_NOR2X1_42 ( );
FILL FILL_0_NAND2X1_102 ( );
FILL FILL_1_NAND2X1_102 ( );
FILL FILL_2_NAND2X1_102 ( );
FILL FILL_3_NAND2X1_102 ( );
FILL FILL_4_NAND2X1_102 ( );
FILL FILL_5_NAND2X1_102 ( );
FILL FILL_6_NAND2X1_102 ( );
FILL FILL_0_NAND2X1_80 ( );
FILL FILL_1_NAND2X1_80 ( );
FILL FILL_2_NAND2X1_80 ( );
FILL FILL_3_NAND2X1_80 ( );
FILL FILL_4_NAND2X1_80 ( );
FILL FILL_5_NAND2X1_80 ( );
FILL FILL_6_NAND2X1_80 ( );
FILL FILL_0_INVX1_115 ( );
FILL FILL_1_INVX1_115 ( );
FILL FILL_2_INVX1_115 ( );
FILL FILL_3_INVX1_115 ( );
FILL FILL_0_OAI21X1_102 ( );
FILL FILL_1_OAI21X1_102 ( );
FILL FILL_2_OAI21X1_102 ( );
FILL FILL_3_OAI21X1_102 ( );
FILL FILL_4_OAI21X1_102 ( );
FILL FILL_5_OAI21X1_102 ( );
FILL FILL_6_OAI21X1_102 ( );
FILL FILL_7_OAI21X1_102 ( );
FILL FILL_8_OAI21X1_102 ( );
FILL FILL_9_OAI21X1_102 ( );
FILL FILL_0_DFFSR_70 ( );
FILL FILL_1_DFFSR_70 ( );
FILL FILL_2_DFFSR_70 ( );
FILL FILL_3_DFFSR_70 ( );
FILL FILL_4_DFFSR_70 ( );
FILL FILL_5_DFFSR_70 ( );
FILL FILL_6_DFFSR_70 ( );
FILL FILL_7_DFFSR_70 ( );
FILL FILL_8_DFFSR_70 ( );
FILL FILL_9_DFFSR_70 ( );
FILL FILL_10_DFFSR_70 ( );
FILL FILL_11_DFFSR_70 ( );
FILL FILL_12_DFFSR_70 ( );
FILL FILL_13_DFFSR_70 ( );
FILL FILL_14_DFFSR_70 ( );
FILL FILL_15_DFFSR_70 ( );
FILL FILL_16_DFFSR_70 ( );
FILL FILL_17_DFFSR_70 ( );
FILL FILL_18_DFFSR_70 ( );
FILL FILL_19_DFFSR_70 ( );
FILL FILL_20_DFFSR_70 ( );
FILL FILL_21_DFFSR_70 ( );
FILL FILL_22_DFFSR_70 ( );
FILL FILL_23_DFFSR_70 ( );
FILL FILL_24_DFFSR_70 ( );
FILL FILL_25_DFFSR_70 ( );
FILL FILL_26_DFFSR_70 ( );
FILL FILL_27_DFFSR_70 ( );
FILL FILL_28_DFFSR_70 ( );
FILL FILL_29_DFFSR_70 ( );
FILL FILL_30_DFFSR_70 ( );
FILL FILL_31_DFFSR_70 ( );
FILL FILL_32_DFFSR_70 ( );
FILL FILL_33_DFFSR_70 ( );
FILL FILL_34_DFFSR_70 ( );
FILL FILL_35_DFFSR_70 ( );
FILL FILL_36_DFFSR_70 ( );
FILL FILL_37_DFFSR_70 ( );
FILL FILL_38_DFFSR_70 ( );
FILL FILL_39_DFFSR_70 ( );
FILL FILL_40_DFFSR_70 ( );
FILL FILL_41_DFFSR_70 ( );
FILL FILL_42_DFFSR_70 ( );
FILL FILL_43_DFFSR_70 ( );
FILL FILL_44_DFFSR_70 ( );
FILL FILL_45_DFFSR_70 ( );
FILL FILL_46_DFFSR_70 ( );
FILL FILL_47_DFFSR_70 ( );
FILL FILL_48_DFFSR_70 ( );
FILL FILL_49_DFFSR_70 ( );
FILL FILL_50_DFFSR_70 ( );
FILL FILL_51_DFFSR_70 ( );
FILL FILL_0_NAND2X1_139 ( );
FILL FILL_1_NAND2X1_139 ( );
FILL FILL_2_NAND2X1_139 ( );
FILL FILL_3_NAND2X1_139 ( );
FILL FILL_4_NAND2X1_139 ( );
FILL FILL_5_NAND2X1_139 ( );
FILL FILL_6_NAND2X1_139 ( );
FILL FILL_0_INVX1_426 ( );
FILL FILL_1_INVX1_426 ( );
FILL FILL_2_INVX1_426 ( );
FILL FILL_3_INVX1_426 ( );
FILL FILL_0_NOR2X1_47 ( );
FILL FILL_1_NOR2X1_47 ( );
FILL FILL_2_NOR2X1_47 ( );
FILL FILL_3_NOR2X1_47 ( );
FILL FILL_4_NOR2X1_47 ( );
FILL FILL_5_NOR2X1_47 ( );
FILL FILL_6_NOR2X1_47 ( );
FILL FILL_0_NAND2X1_274 ( );
FILL FILL_1_NAND2X1_274 ( );
FILL FILL_2_NAND2X1_274 ( );
FILL FILL_3_NAND2X1_274 ( );
FILL FILL_4_NAND2X1_274 ( );
FILL FILL_5_NAND2X1_274 ( );
FILL FILL_6_NAND2X1_274 ( );
FILL FILL_0_INVX1_425 ( );
FILL FILL_1_INVX1_425 ( );
FILL FILL_2_INVX1_425 ( );
FILL FILL_3_INVX1_425 ( );
FILL FILL_4_INVX1_425 ( );
FILL FILL_0_DFFPOSX1_31 ( );
FILL FILL_1_DFFPOSX1_31 ( );
FILL FILL_2_DFFPOSX1_31 ( );
FILL FILL_3_DFFPOSX1_31 ( );
FILL FILL_4_DFFPOSX1_31 ( );
FILL FILL_5_DFFPOSX1_31 ( );
FILL FILL_6_DFFPOSX1_31 ( );
FILL FILL_7_DFFPOSX1_31 ( );
FILL FILL_8_DFFPOSX1_31 ( );
FILL FILL_9_DFFPOSX1_31 ( );
FILL FILL_10_DFFPOSX1_31 ( );
FILL FILL_11_DFFPOSX1_31 ( );
FILL FILL_12_DFFPOSX1_31 ( );
FILL FILL_13_DFFPOSX1_31 ( );
FILL FILL_14_DFFPOSX1_31 ( );
FILL FILL_15_DFFPOSX1_31 ( );
FILL FILL_16_DFFPOSX1_31 ( );
FILL FILL_17_DFFPOSX1_31 ( );
FILL FILL_18_DFFPOSX1_31 ( );
FILL FILL_19_DFFPOSX1_31 ( );
FILL FILL_20_DFFPOSX1_31 ( );
FILL FILL_21_DFFPOSX1_31 ( );
FILL FILL_22_DFFPOSX1_31 ( );
FILL FILL_23_DFFPOSX1_31 ( );
FILL FILL_24_DFFPOSX1_31 ( );
FILL FILL_25_DFFPOSX1_31 ( );
FILL FILL_26_DFFPOSX1_31 ( );
FILL FILL_27_DFFPOSX1_31 ( );
FILL FILL_0_NAND2X1_241 ( );
FILL FILL_1_NAND2X1_241 ( );
FILL FILL_2_NAND2X1_241 ( );
FILL FILL_3_NAND2X1_241 ( );
FILL FILL_4_NAND2X1_241 ( );
FILL FILL_5_NAND2X1_241 ( );
FILL FILL_6_NAND2X1_241 ( );
FILL FILL_0_NOR2X1_27 ( );
FILL FILL_1_NOR2X1_27 ( );
FILL FILL_2_NOR2X1_27 ( );
FILL FILL_3_NOR2X1_27 ( );
FILL FILL_4_NOR2X1_27 ( );
FILL FILL_5_NOR2X1_27 ( );
FILL FILL_6_NOR2X1_27 ( );
FILL FILL_0_OAI22X1_36 ( );
FILL FILL_1_OAI22X1_36 ( );
FILL FILL_2_OAI22X1_36 ( );
FILL FILL_3_OAI22X1_36 ( );
FILL FILL_4_OAI22X1_36 ( );
FILL FILL_5_OAI22X1_36 ( );
FILL FILL_6_OAI22X1_36 ( );
FILL FILL_7_OAI22X1_36 ( );
FILL FILL_8_OAI22X1_36 ( );
FILL FILL_9_OAI22X1_36 ( );
FILL FILL_10_OAI22X1_36 ( );
FILL FILL_0_INVX1_57 ( );
FILL FILL_1_INVX1_57 ( );
FILL FILL_2_INVX1_57 ( );
FILL FILL_3_INVX1_57 ( );
FILL FILL_0_OAI21X1_15 ( );
FILL FILL_1_OAI21X1_15 ( );
FILL FILL_2_OAI21X1_15 ( );
FILL FILL_3_OAI21X1_15 ( );
FILL FILL_4_OAI21X1_15 ( );
FILL FILL_5_OAI21X1_15 ( );
FILL FILL_6_OAI21X1_15 ( );
FILL FILL_7_OAI21X1_15 ( );
FILL FILL_8_OAI21X1_15 ( );
FILL FILL_9_OAI21X1_15 ( );
FILL FILL_0_NOR2X1_13 ( );
FILL FILL_1_NOR2X1_13 ( );
FILL FILL_2_NOR2X1_13 ( );
FILL FILL_3_NOR2X1_13 ( );
FILL FILL_4_NOR2X1_13 ( );
FILL FILL_5_NOR2X1_13 ( );
FILL FILL_6_NOR2X1_13 ( );
FILL FILL_0_DFFSR_41 ( );
FILL FILL_1_DFFSR_41 ( );
FILL FILL_2_DFFSR_41 ( );
FILL FILL_3_DFFSR_41 ( );
FILL FILL_4_DFFSR_41 ( );
FILL FILL_5_DFFSR_41 ( );
FILL FILL_6_DFFSR_41 ( );
FILL FILL_7_DFFSR_41 ( );
FILL FILL_8_DFFSR_41 ( );
FILL FILL_9_DFFSR_41 ( );
FILL FILL_10_DFFSR_41 ( );
FILL FILL_11_DFFSR_41 ( );
FILL FILL_12_DFFSR_41 ( );
FILL FILL_13_DFFSR_41 ( );
FILL FILL_14_DFFSR_41 ( );
FILL FILL_15_DFFSR_41 ( );
FILL FILL_16_DFFSR_41 ( );
FILL FILL_17_DFFSR_41 ( );
FILL FILL_18_DFFSR_41 ( );
FILL FILL_19_DFFSR_41 ( );
FILL FILL_20_DFFSR_41 ( );
FILL FILL_21_DFFSR_41 ( );
FILL FILL_22_DFFSR_41 ( );
FILL FILL_23_DFFSR_41 ( );
FILL FILL_24_DFFSR_41 ( );
FILL FILL_25_DFFSR_41 ( );
FILL FILL_26_DFFSR_41 ( );
FILL FILL_27_DFFSR_41 ( );
FILL FILL_28_DFFSR_41 ( );
FILL FILL_29_DFFSR_41 ( );
FILL FILL_30_DFFSR_41 ( );
FILL FILL_31_DFFSR_41 ( );
FILL FILL_32_DFFSR_41 ( );
FILL FILL_33_DFFSR_41 ( );
FILL FILL_34_DFFSR_41 ( );
FILL FILL_35_DFFSR_41 ( );
FILL FILL_36_DFFSR_41 ( );
FILL FILL_37_DFFSR_41 ( );
FILL FILL_38_DFFSR_41 ( );
FILL FILL_39_DFFSR_41 ( );
FILL FILL_40_DFFSR_41 ( );
FILL FILL_41_DFFSR_41 ( );
FILL FILL_42_DFFSR_41 ( );
FILL FILL_43_DFFSR_41 ( );
FILL FILL_44_DFFSR_41 ( );
FILL FILL_45_DFFSR_41 ( );
FILL FILL_46_DFFSR_41 ( );
FILL FILL_47_DFFSR_41 ( );
FILL FILL_48_DFFSR_41 ( );
FILL FILL_49_DFFSR_41 ( );
FILL FILL_50_DFFSR_41 ( );
FILL FILL_0_INVX1_267 ( );
FILL FILL_1_INVX1_267 ( );
FILL FILL_2_INVX1_267 ( );
FILL FILL_3_INVX1_267 ( );
FILL FILL_0_NAND2X1_57 ( );
FILL FILL_1_NAND2X1_57 ( );
FILL FILL_2_NAND2X1_57 ( );
FILL FILL_3_NAND2X1_57 ( );
FILL FILL_4_NAND2X1_57 ( );
FILL FILL_5_NAND2X1_57 ( );
FILL FILL_6_NAND2X1_57 ( );
FILL FILL_0_AND2X2_3 ( );
FILL FILL_1_AND2X2_3 ( );
FILL FILL_2_AND2X2_3 ( );
FILL FILL_3_AND2X2_3 ( );
FILL FILL_4_AND2X2_3 ( );
FILL FILL_5_AND2X2_3 ( );
FILL FILL_6_AND2X2_3 ( );
FILL FILL_7_AND2X2_3 ( );
FILL FILL_8_AND2X2_3 ( );
FILL FILL_0_NOR2X1_6 ( );
FILL FILL_1_NOR2X1_6 ( );
FILL FILL_2_NOR2X1_6 ( );
FILL FILL_3_NOR2X1_6 ( );
FILL FILL_4_NOR2X1_6 ( );
FILL FILL_5_NOR2X1_6 ( );
FILL FILL_6_NOR2X1_6 ( );
FILL FILL_0_OAI21X1_181 ( );
FILL FILL_1_OAI21X1_181 ( );
FILL FILL_2_OAI21X1_181 ( );
FILL FILL_3_OAI21X1_181 ( );
FILL FILL_4_OAI21X1_181 ( );
FILL FILL_5_OAI21X1_181 ( );
FILL FILL_6_OAI21X1_181 ( );
FILL FILL_7_OAI21X1_181 ( );
FILL FILL_8_OAI21X1_181 ( );
FILL FILL_9_OAI21X1_181 ( );
FILL FILL_0_NOR2X1_5 ( );
FILL FILL_1_NOR2X1_5 ( );
FILL FILL_2_NOR2X1_5 ( );
FILL FILL_3_NOR2X1_5 ( );
FILL FILL_4_NOR2X1_5 ( );
FILL FILL_5_NOR2X1_5 ( );
FILL FILL_6_NOR2X1_5 ( );
FILL FILL_0_INVX1_234 ( );
FILL FILL_1_INVX1_234 ( );
FILL FILL_2_INVX1_234 ( );
FILL FILL_3_INVX1_234 ( );
FILL FILL_0_AOI21X1_10 ( );
FILL FILL_1_AOI21X1_10 ( );
FILL FILL_2_AOI21X1_10 ( );
FILL FILL_3_AOI21X1_10 ( );
FILL FILL_4_AOI21X1_10 ( );
FILL FILL_5_AOI21X1_10 ( );
FILL FILL_6_AOI21X1_10 ( );
FILL FILL_7_AOI21X1_10 ( );
FILL FILL_8_AOI21X1_10 ( );
FILL FILL_9_AOI21X1_10 ( );
FILL FILL_0_DFFSR_160 ( );
FILL FILL_1_DFFSR_160 ( );
FILL FILL_2_DFFSR_160 ( );
FILL FILL_3_DFFSR_160 ( );
FILL FILL_4_DFFSR_160 ( );
FILL FILL_5_DFFSR_160 ( );
FILL FILL_6_DFFSR_160 ( );
FILL FILL_7_DFFSR_160 ( );
FILL FILL_8_DFFSR_160 ( );
FILL FILL_9_DFFSR_160 ( );
FILL FILL_10_DFFSR_160 ( );
FILL FILL_11_DFFSR_160 ( );
FILL FILL_12_DFFSR_160 ( );
FILL FILL_13_DFFSR_160 ( );
FILL FILL_14_DFFSR_160 ( );
FILL FILL_15_DFFSR_160 ( );
FILL FILL_16_DFFSR_160 ( );
FILL FILL_17_DFFSR_160 ( );
FILL FILL_18_DFFSR_160 ( );
FILL FILL_19_DFFSR_160 ( );
FILL FILL_20_DFFSR_160 ( );
FILL FILL_21_DFFSR_160 ( );
FILL FILL_22_DFFSR_160 ( );
FILL FILL_23_DFFSR_160 ( );
FILL FILL_24_DFFSR_160 ( );
FILL FILL_25_DFFSR_160 ( );
FILL FILL_26_DFFSR_160 ( );
FILL FILL_27_DFFSR_160 ( );
FILL FILL_28_DFFSR_160 ( );
FILL FILL_29_DFFSR_160 ( );
FILL FILL_30_DFFSR_160 ( );
FILL FILL_31_DFFSR_160 ( );
FILL FILL_32_DFFSR_160 ( );
FILL FILL_33_DFFSR_160 ( );
FILL FILL_34_DFFSR_160 ( );
FILL FILL_35_DFFSR_160 ( );
FILL FILL_36_DFFSR_160 ( );
FILL FILL_37_DFFSR_160 ( );
FILL FILL_38_DFFSR_160 ( );
FILL FILL_39_DFFSR_160 ( );
FILL FILL_40_DFFSR_160 ( );
FILL FILL_41_DFFSR_160 ( );
FILL FILL_42_DFFSR_160 ( );
FILL FILL_43_DFFSR_160 ( );
FILL FILL_44_DFFSR_160 ( );
FILL FILL_45_DFFSR_160 ( );
FILL FILL_46_DFFSR_160 ( );
FILL FILL_47_DFFSR_160 ( );
FILL FILL_48_DFFSR_160 ( );
FILL FILL_49_DFFSR_160 ( );
FILL FILL_50_DFFSR_160 ( );
FILL FILL_0_NAND2X1_198 ( );
FILL FILL_1_NAND2X1_198 ( );
FILL FILL_2_NAND2X1_198 ( );
FILL FILL_3_NAND2X1_198 ( );
FILL FILL_4_NAND2X1_198 ( );
FILL FILL_5_NAND2X1_198 ( );
FILL FILL_6_NAND2X1_198 ( );
FILL FILL_0_OAI21X1_209 ( );
FILL FILL_1_OAI21X1_209 ( );
FILL FILL_2_OAI21X1_209 ( );
FILL FILL_3_OAI21X1_209 ( );
FILL FILL_4_OAI21X1_209 ( );
FILL FILL_5_OAI21X1_209 ( );
FILL FILL_6_OAI21X1_209 ( );
FILL FILL_7_OAI21X1_209 ( );
FILL FILL_8_OAI21X1_209 ( );
FILL FILL_9_OAI21X1_209 ( );
FILL FILL_0_DFFSR_101 ( );
FILL FILL_1_DFFSR_101 ( );
FILL FILL_2_DFFSR_101 ( );
FILL FILL_3_DFFSR_101 ( );
FILL FILL_4_DFFSR_101 ( );
FILL FILL_5_DFFSR_101 ( );
FILL FILL_6_DFFSR_101 ( );
FILL FILL_7_DFFSR_101 ( );
FILL FILL_8_DFFSR_101 ( );
FILL FILL_9_DFFSR_101 ( );
FILL FILL_10_DFFSR_101 ( );
FILL FILL_11_DFFSR_101 ( );
FILL FILL_12_DFFSR_101 ( );
FILL FILL_13_DFFSR_101 ( );
FILL FILL_14_DFFSR_101 ( );
FILL FILL_15_DFFSR_101 ( );
FILL FILL_16_DFFSR_101 ( );
FILL FILL_17_DFFSR_101 ( );
FILL FILL_18_DFFSR_101 ( );
FILL FILL_19_DFFSR_101 ( );
FILL FILL_20_DFFSR_101 ( );
FILL FILL_21_DFFSR_101 ( );
FILL FILL_22_DFFSR_101 ( );
FILL FILL_23_DFFSR_101 ( );
FILL FILL_24_DFFSR_101 ( );
FILL FILL_25_DFFSR_101 ( );
FILL FILL_26_DFFSR_101 ( );
FILL FILL_27_DFFSR_101 ( );
FILL FILL_28_DFFSR_101 ( );
FILL FILL_29_DFFSR_101 ( );
FILL FILL_30_DFFSR_101 ( );
FILL FILL_31_DFFSR_101 ( );
FILL FILL_32_DFFSR_101 ( );
FILL FILL_33_DFFSR_101 ( );
FILL FILL_34_DFFSR_101 ( );
FILL FILL_35_DFFSR_101 ( );
FILL FILL_36_DFFSR_101 ( );
FILL FILL_37_DFFSR_101 ( );
FILL FILL_38_DFFSR_101 ( );
FILL FILL_39_DFFSR_101 ( );
FILL FILL_40_DFFSR_101 ( );
FILL FILL_41_DFFSR_101 ( );
FILL FILL_42_DFFSR_101 ( );
FILL FILL_43_DFFSR_101 ( );
FILL FILL_44_DFFSR_101 ( );
FILL FILL_45_DFFSR_101 ( );
FILL FILL_46_DFFSR_101 ( );
FILL FILL_47_DFFSR_101 ( );
FILL FILL_48_DFFSR_101 ( );
FILL FILL_49_DFFSR_101 ( );
FILL FILL_50_DFFSR_101 ( );
FILL FILL_0_INVX1_372 ( );
FILL FILL_1_INVX1_372 ( );
FILL FILL_2_INVX1_372 ( );
FILL FILL_3_INVX1_372 ( );
FILL FILL_4_INVX1_372 ( );
FILL FILL_0_INVX1_377 ( );
FILL FILL_1_INVX1_377 ( );
FILL FILL_2_INVX1_377 ( );
FILL FILL_3_INVX1_377 ( );
FILL FILL_0_OAI22X1_41 ( );
FILL FILL_1_OAI22X1_41 ( );
FILL FILL_2_OAI22X1_41 ( );
FILL FILL_3_OAI22X1_41 ( );
FILL FILL_4_OAI22X1_41 ( );
FILL FILL_5_OAI22X1_41 ( );
FILL FILL_6_OAI22X1_41 ( );
FILL FILL_7_OAI22X1_41 ( );
FILL FILL_8_OAI22X1_41 ( );
FILL FILL_9_OAI22X1_41 ( );
FILL FILL_10_OAI22X1_41 ( );
FILL FILL_11_OAI22X1_41 ( );
FILL FILL_0_NOR2X1_30 ( );
FILL FILL_1_NOR2X1_30 ( );
FILL FILL_2_NOR2X1_30 ( );
FILL FILL_3_NOR2X1_30 ( );
FILL FILL_4_NOR2X1_30 ( );
FILL FILL_5_NOR2X1_30 ( );
FILL FILL_6_NOR2X1_30 ( );
FILL FILL_0_NAND2X1_243 ( );
FILL FILL_1_NAND2X1_243 ( );
FILL FILL_2_NAND2X1_243 ( );
FILL FILL_3_NAND2X1_243 ( );
FILL FILL_4_NAND2X1_243 ( );
FILL FILL_5_NAND2X1_243 ( );
FILL FILL_6_NAND2X1_243 ( );
FILL FILL_0_OAI22X1_65 ( );
FILL FILL_1_OAI22X1_65 ( );
FILL FILL_2_OAI22X1_65 ( );
FILL FILL_3_OAI22X1_65 ( );
FILL FILL_4_OAI22X1_65 ( );
FILL FILL_5_OAI22X1_65 ( );
FILL FILL_6_OAI22X1_65 ( );
FILL FILL_7_OAI22X1_65 ( );
FILL FILL_8_OAI22X1_65 ( );
FILL FILL_9_OAI22X1_65 ( );
FILL FILL_10_OAI22X1_65 ( );
FILL FILL_11_OAI22X1_65 ( );
FILL FILL_0_INVX1_389 ( );
FILL FILL_1_INVX1_389 ( );
FILL FILL_2_INVX1_389 ( );
FILL FILL_3_INVX1_389 ( );
FILL FILL_0_INVX1_375 ( );
FILL FILL_1_INVX1_375 ( );
FILL FILL_2_INVX1_375 ( );
FILL FILL_3_INVX1_375 ( );
FILL FILL_0_INVX1_79 ( );
FILL FILL_1_INVX1_79 ( );
FILL FILL_2_INVX1_79 ( );
FILL FILL_3_INVX1_79 ( );
FILL FILL_4_INVX1_79 ( );
FILL FILL_0_OAI21X1_70 ( );
FILL FILL_1_OAI21X1_70 ( );
FILL FILL_2_OAI21X1_70 ( );
FILL FILL_3_OAI21X1_70 ( );
FILL FILL_4_OAI21X1_70 ( );
FILL FILL_5_OAI21X1_70 ( );
FILL FILL_6_OAI21X1_70 ( );
FILL FILL_7_OAI21X1_70 ( );
FILL FILL_8_OAI21X1_70 ( );
FILL FILL_0_INVX1_124 ( );
FILL FILL_1_INVX1_124 ( );
FILL FILL_2_INVX1_124 ( );
FILL FILL_3_INVX1_124 ( );
FILL FILL_4_INVX1_124 ( );
FILL FILL_0_DFFSR_110 ( );
FILL FILL_1_DFFSR_110 ( );
FILL FILL_2_DFFSR_110 ( );
FILL FILL_3_DFFSR_110 ( );
FILL FILL_4_DFFSR_110 ( );
FILL FILL_5_DFFSR_110 ( );
FILL FILL_6_DFFSR_110 ( );
FILL FILL_7_DFFSR_110 ( );
FILL FILL_8_DFFSR_110 ( );
FILL FILL_9_DFFSR_110 ( );
FILL FILL_10_DFFSR_110 ( );
FILL FILL_11_DFFSR_110 ( );
FILL FILL_12_DFFSR_110 ( );
FILL FILL_13_DFFSR_110 ( );
FILL FILL_14_DFFSR_110 ( );
FILL FILL_15_DFFSR_110 ( );
FILL FILL_16_DFFSR_110 ( );
FILL FILL_17_DFFSR_110 ( );
FILL FILL_18_DFFSR_110 ( );
FILL FILL_19_DFFSR_110 ( );
FILL FILL_20_DFFSR_110 ( );
FILL FILL_21_DFFSR_110 ( );
FILL FILL_22_DFFSR_110 ( );
FILL FILL_23_DFFSR_110 ( );
FILL FILL_24_DFFSR_110 ( );
FILL FILL_25_DFFSR_110 ( );
FILL FILL_26_DFFSR_110 ( );
FILL FILL_27_DFFSR_110 ( );
FILL FILL_28_DFFSR_110 ( );
FILL FILL_29_DFFSR_110 ( );
FILL FILL_30_DFFSR_110 ( );
FILL FILL_31_DFFSR_110 ( );
FILL FILL_32_DFFSR_110 ( );
FILL FILL_33_DFFSR_110 ( );
FILL FILL_34_DFFSR_110 ( );
FILL FILL_35_DFFSR_110 ( );
FILL FILL_36_DFFSR_110 ( );
FILL FILL_37_DFFSR_110 ( );
FILL FILL_38_DFFSR_110 ( );
FILL FILL_39_DFFSR_110 ( );
FILL FILL_40_DFFSR_110 ( );
FILL FILL_41_DFFSR_110 ( );
FILL FILL_42_DFFSR_110 ( );
FILL FILL_43_DFFSR_110 ( );
FILL FILL_44_DFFSR_110 ( );
FILL FILL_45_DFFSR_110 ( );
FILL FILL_46_DFFSR_110 ( );
FILL FILL_47_DFFSR_110 ( );
FILL FILL_48_DFFSR_110 ( );
FILL FILL_49_DFFSR_110 ( );
FILL FILL_50_DFFSR_110 ( );
FILL FILL_0_NAND2X1_138 ( );
FILL FILL_1_NAND2X1_138 ( );
FILL FILL_2_NAND2X1_138 ( );
FILL FILL_3_NAND2X1_138 ( );
FILL FILL_4_NAND2X1_138 ( );
FILL FILL_5_NAND2X1_138 ( );
FILL FILL_6_NAND2X1_138 ( );
FILL FILL_0_OAI21X1_138 ( );
FILL FILL_1_OAI21X1_138 ( );
FILL FILL_2_OAI21X1_138 ( );
FILL FILL_3_OAI21X1_138 ( );
FILL FILL_4_OAI21X1_138 ( );
FILL FILL_5_OAI21X1_138 ( );
FILL FILL_6_OAI21X1_138 ( );
FILL FILL_7_OAI21X1_138 ( );
FILL FILL_8_OAI21X1_138 ( );
FILL FILL_0_INVX1_156 ( );
FILL FILL_1_INVX1_156 ( );
FILL FILL_2_INVX1_156 ( );
FILL FILL_3_INVX1_156 ( );
FILL FILL_4_INVX1_156 ( );
FILL FILL_0_XOR2X1_11 ( );
FILL FILL_1_XOR2X1_11 ( );
FILL FILL_2_XOR2X1_11 ( );
FILL FILL_3_XOR2X1_11 ( );
FILL FILL_4_XOR2X1_11 ( );
FILL FILL_5_XOR2X1_11 ( );
FILL FILL_6_XOR2X1_11 ( );
FILL FILL_7_XOR2X1_11 ( );
FILL FILL_8_XOR2X1_11 ( );
FILL FILL_9_XOR2X1_11 ( );
FILL FILL_10_XOR2X1_11 ( );
FILL FILL_11_XOR2X1_11 ( );
FILL FILL_12_XOR2X1_11 ( );
FILL FILL_13_XOR2X1_11 ( );
FILL FILL_14_XOR2X1_11 ( );
FILL FILL_15_XOR2X1_11 ( );
FILL FILL_0_NAND2X1_24 ( );
FILL FILL_1_NAND2X1_24 ( );
FILL FILL_2_NAND2X1_24 ( );
FILL FILL_3_NAND2X1_24 ( );
FILL FILL_4_NAND2X1_24 ( );
FILL FILL_5_NAND2X1_24 ( );
FILL FILL_6_NAND2X1_24 ( );
FILL FILL_0_INVX1_321 ( );
FILL FILL_1_INVX1_321 ( );
FILL FILL_2_INVX1_321 ( );
FILL FILL_3_INVX1_321 ( );
FILL FILL_4_INVX1_321 ( );
FILL FILL_0_OAI22X1_33 ( );
FILL FILL_1_OAI22X1_33 ( );
FILL FILL_2_OAI22X1_33 ( );
FILL FILL_3_OAI22X1_33 ( );
FILL FILL_4_OAI22X1_33 ( );
FILL FILL_5_OAI22X1_33 ( );
FILL FILL_6_OAI22X1_33 ( );
FILL FILL_7_OAI22X1_33 ( );
FILL FILL_8_OAI22X1_33 ( );
FILL FILL_9_OAI22X1_33 ( );
FILL FILL_10_OAI22X1_33 ( );
FILL FILL_0_DFFSR_38 ( );
FILL FILL_1_DFFSR_38 ( );
FILL FILL_2_DFFSR_38 ( );
FILL FILL_3_DFFSR_38 ( );
FILL FILL_4_DFFSR_38 ( );
FILL FILL_5_DFFSR_38 ( );
FILL FILL_6_DFFSR_38 ( );
FILL FILL_7_DFFSR_38 ( );
FILL FILL_8_DFFSR_38 ( );
FILL FILL_9_DFFSR_38 ( );
FILL FILL_10_DFFSR_38 ( );
FILL FILL_11_DFFSR_38 ( );
FILL FILL_12_DFFSR_38 ( );
FILL FILL_13_DFFSR_38 ( );
FILL FILL_14_DFFSR_38 ( );
FILL FILL_15_DFFSR_38 ( );
FILL FILL_16_DFFSR_38 ( );
FILL FILL_17_DFFSR_38 ( );
FILL FILL_18_DFFSR_38 ( );
FILL FILL_19_DFFSR_38 ( );
FILL FILL_20_DFFSR_38 ( );
FILL FILL_21_DFFSR_38 ( );
FILL FILL_22_DFFSR_38 ( );
FILL FILL_23_DFFSR_38 ( );
FILL FILL_24_DFFSR_38 ( );
FILL FILL_25_DFFSR_38 ( );
FILL FILL_26_DFFSR_38 ( );
FILL FILL_27_DFFSR_38 ( );
FILL FILL_28_DFFSR_38 ( );
FILL FILL_29_DFFSR_38 ( );
FILL FILL_30_DFFSR_38 ( );
FILL FILL_31_DFFSR_38 ( );
FILL FILL_32_DFFSR_38 ( );
FILL FILL_33_DFFSR_38 ( );
FILL FILL_34_DFFSR_38 ( );
FILL FILL_35_DFFSR_38 ( );
FILL FILL_36_DFFSR_38 ( );
FILL FILL_37_DFFSR_38 ( );
FILL FILL_38_DFFSR_38 ( );
FILL FILL_39_DFFSR_38 ( );
FILL FILL_40_DFFSR_38 ( );
FILL FILL_41_DFFSR_38 ( );
FILL FILL_42_DFFSR_38 ( );
FILL FILL_43_DFFSR_38 ( );
FILL FILL_44_DFFSR_38 ( );
FILL FILL_45_DFFSR_38 ( );
FILL FILL_46_DFFSR_38 ( );
FILL FILL_47_DFFSR_38 ( );
FILL FILL_48_DFFSR_38 ( );
FILL FILL_49_DFFSR_38 ( );
FILL FILL_50_DFFSR_38 ( );
FILL FILL_0_OAI22X1_8 ( );
FILL FILL_1_OAI22X1_8 ( );
FILL FILL_2_OAI22X1_8 ( );
FILL FILL_3_OAI22X1_8 ( );
FILL FILL_4_OAI22X1_8 ( );
FILL FILL_5_OAI22X1_8 ( );
FILL FILL_6_OAI22X1_8 ( );
FILL FILL_7_OAI22X1_8 ( );
FILL FILL_8_OAI22X1_8 ( );
FILL FILL_9_OAI22X1_8 ( );
FILL FILL_10_OAI22X1_8 ( );
FILL FILL_11_OAI22X1_8 ( );
FILL FILL_0_CLKBUF1_10 ( );
FILL FILL_1_CLKBUF1_10 ( );
FILL FILL_2_CLKBUF1_10 ( );
FILL FILL_3_CLKBUF1_10 ( );
FILL FILL_4_CLKBUF1_10 ( );
FILL FILL_5_CLKBUF1_10 ( );
FILL FILL_6_CLKBUF1_10 ( );
FILL FILL_7_CLKBUF1_10 ( );
FILL FILL_8_CLKBUF1_10 ( );
FILL FILL_9_CLKBUF1_10 ( );
FILL FILL_10_CLKBUF1_10 ( );
FILL FILL_11_CLKBUF1_10 ( );
FILL FILL_12_CLKBUF1_10 ( );
FILL FILL_13_CLKBUF1_10 ( );
FILL FILL_14_CLKBUF1_10 ( );
FILL FILL_15_CLKBUF1_10 ( );
FILL FILL_16_CLKBUF1_10 ( );
FILL FILL_17_CLKBUF1_10 ( );
FILL FILL_18_CLKBUF1_10 ( );
FILL FILL_19_CLKBUF1_10 ( );
FILL FILL_20_CLKBUF1_10 ( );
FILL FILL_0_INVX1_271 ( );
FILL FILL_1_INVX1_271 ( );
FILL FILL_2_INVX1_271 ( );
FILL FILL_3_INVX1_271 ( );
FILL FILL_4_INVX1_271 ( );
FILL FILL_0_DFFSR_57 ( );
FILL FILL_1_DFFSR_57 ( );
FILL FILL_2_DFFSR_57 ( );
FILL FILL_3_DFFSR_57 ( );
FILL FILL_4_DFFSR_57 ( );
FILL FILL_5_DFFSR_57 ( );
FILL FILL_6_DFFSR_57 ( );
FILL FILL_7_DFFSR_57 ( );
FILL FILL_8_DFFSR_57 ( );
FILL FILL_9_DFFSR_57 ( );
FILL FILL_10_DFFSR_57 ( );
FILL FILL_11_DFFSR_57 ( );
FILL FILL_12_DFFSR_57 ( );
FILL FILL_13_DFFSR_57 ( );
FILL FILL_14_DFFSR_57 ( );
FILL FILL_15_DFFSR_57 ( );
FILL FILL_16_DFFSR_57 ( );
FILL FILL_17_DFFSR_57 ( );
FILL FILL_18_DFFSR_57 ( );
FILL FILL_19_DFFSR_57 ( );
FILL FILL_20_DFFSR_57 ( );
FILL FILL_21_DFFSR_57 ( );
FILL FILL_22_DFFSR_57 ( );
FILL FILL_23_DFFSR_57 ( );
FILL FILL_24_DFFSR_57 ( );
FILL FILL_25_DFFSR_57 ( );
FILL FILL_26_DFFSR_57 ( );
FILL FILL_27_DFFSR_57 ( );
FILL FILL_28_DFFSR_57 ( );
FILL FILL_29_DFFSR_57 ( );
FILL FILL_30_DFFSR_57 ( );
FILL FILL_31_DFFSR_57 ( );
FILL FILL_32_DFFSR_57 ( );
FILL FILL_33_DFFSR_57 ( );
FILL FILL_34_DFFSR_57 ( );
FILL FILL_35_DFFSR_57 ( );
FILL FILL_36_DFFSR_57 ( );
FILL FILL_37_DFFSR_57 ( );
FILL FILL_38_DFFSR_57 ( );
FILL FILL_39_DFFSR_57 ( );
FILL FILL_40_DFFSR_57 ( );
FILL FILL_41_DFFSR_57 ( );
FILL FILL_42_DFFSR_57 ( );
FILL FILL_43_DFFSR_57 ( );
FILL FILL_44_DFFSR_57 ( );
FILL FILL_45_DFFSR_57 ( );
FILL FILL_46_DFFSR_57 ( );
FILL FILL_47_DFFSR_57 ( );
FILL FILL_48_DFFSR_57 ( );
FILL FILL_49_DFFSR_57 ( );
FILL FILL_50_DFFSR_57 ( );
FILL FILL_51_DFFSR_57 ( );
FILL FILL_0_NAND2X1_163 ( );
FILL FILL_1_NAND2X1_163 ( );
FILL FILL_2_NAND2X1_163 ( );
FILL FILL_3_NAND2X1_163 ( );
FILL FILL_4_NAND2X1_163 ( );
FILL FILL_5_NAND2X1_163 ( );
FILL FILL_6_NAND2X1_163 ( );
FILL FILL_0_OAI21X1_189 ( );
FILL FILL_1_OAI21X1_189 ( );
FILL FILL_2_OAI21X1_189 ( );
FILL FILL_3_OAI21X1_189 ( );
FILL FILL_4_OAI21X1_189 ( );
FILL FILL_5_OAI21X1_189 ( );
FILL FILL_6_OAI21X1_189 ( );
FILL FILL_7_OAI21X1_189 ( );
FILL FILL_8_OAI21X1_189 ( );
FILL FILL_9_OAI21X1_189 ( );
FILL FILL_0_INVX1_194 ( );
FILL FILL_1_INVX1_194 ( );
FILL FILL_2_INVX1_194 ( );
FILL FILL_3_INVX1_194 ( );
FILL FILL_4_INVX1_194 ( );
FILL FILL_0_OAI21X1_160 ( );
FILL FILL_1_OAI21X1_160 ( );
FILL FILL_2_OAI21X1_160 ( );
FILL FILL_3_OAI21X1_160 ( );
FILL FILL_4_OAI21X1_160 ( );
FILL FILL_5_OAI21X1_160 ( );
FILL FILL_6_OAI21X1_160 ( );
FILL FILL_7_OAI21X1_160 ( );
FILL FILL_8_OAI21X1_160 ( );
FILL FILL_0_OAI21X1_248 ( );
FILL FILL_1_OAI21X1_248 ( );
FILL FILL_2_OAI21X1_248 ( );
FILL FILL_3_OAI21X1_248 ( );
FILL FILL_4_OAI21X1_248 ( );
FILL FILL_5_OAI21X1_248 ( );
FILL FILL_6_OAI21X1_248 ( );
FILL FILL_7_OAI21X1_248 ( );
FILL FILL_8_OAI21X1_248 ( );
FILL FILL_9_OAI21X1_248 ( );
FILL FILL_0_OAI21X1_199 ( );
FILL FILL_1_OAI21X1_199 ( );
FILL FILL_2_OAI21X1_199 ( );
FILL FILL_3_OAI21X1_199 ( );
FILL FILL_4_OAI21X1_199 ( );
FILL FILL_5_OAI21X1_199 ( );
FILL FILL_6_OAI21X1_199 ( );
FILL FILL_7_OAI21X1_199 ( );
FILL FILL_8_OAI21X1_199 ( );
FILL FILL_9_OAI21X1_199 ( );
FILL FILL_0_NAND2X1_218 ( );
FILL FILL_1_NAND2X1_218 ( );
FILL FILL_2_NAND2X1_218 ( );
FILL FILL_3_NAND2X1_218 ( );
FILL FILL_4_NAND2X1_218 ( );
FILL FILL_5_NAND2X1_218 ( );
FILL FILL_6_NAND2X1_218 ( );
FILL FILL_0_NAND3X1_32 ( );
FILL FILL_1_NAND3X1_32 ( );
FILL FILL_2_NAND3X1_32 ( );
FILL FILL_3_NAND3X1_32 ( );
FILL FILL_4_NAND3X1_32 ( );
FILL FILL_5_NAND3X1_32 ( );
FILL FILL_6_NAND3X1_32 ( );
FILL FILL_7_NAND3X1_32 ( );
FILL FILL_8_NAND3X1_32 ( );
FILL FILL_9_NAND3X1_32 ( );
FILL FILL_0_DFFSR_73 ( );
FILL FILL_1_DFFSR_73 ( );
FILL FILL_2_DFFSR_73 ( );
FILL FILL_3_DFFSR_73 ( );
FILL FILL_4_DFFSR_73 ( );
FILL FILL_5_DFFSR_73 ( );
FILL FILL_6_DFFSR_73 ( );
FILL FILL_7_DFFSR_73 ( );
FILL FILL_8_DFFSR_73 ( );
FILL FILL_9_DFFSR_73 ( );
FILL FILL_10_DFFSR_73 ( );
FILL FILL_11_DFFSR_73 ( );
FILL FILL_12_DFFSR_73 ( );
FILL FILL_13_DFFSR_73 ( );
FILL FILL_14_DFFSR_73 ( );
FILL FILL_15_DFFSR_73 ( );
FILL FILL_16_DFFSR_73 ( );
FILL FILL_17_DFFSR_73 ( );
FILL FILL_18_DFFSR_73 ( );
FILL FILL_19_DFFSR_73 ( );
FILL FILL_20_DFFSR_73 ( );
FILL FILL_21_DFFSR_73 ( );
FILL FILL_22_DFFSR_73 ( );
FILL FILL_23_DFFSR_73 ( );
FILL FILL_24_DFFSR_73 ( );
FILL FILL_25_DFFSR_73 ( );
FILL FILL_26_DFFSR_73 ( );
FILL FILL_27_DFFSR_73 ( );
FILL FILL_28_DFFSR_73 ( );
FILL FILL_29_DFFSR_73 ( );
FILL FILL_30_DFFSR_73 ( );
FILL FILL_31_DFFSR_73 ( );
FILL FILL_32_DFFSR_73 ( );
FILL FILL_33_DFFSR_73 ( );
FILL FILL_34_DFFSR_73 ( );
FILL FILL_35_DFFSR_73 ( );
FILL FILL_36_DFFSR_73 ( );
FILL FILL_37_DFFSR_73 ( );
FILL FILL_38_DFFSR_73 ( );
FILL FILL_39_DFFSR_73 ( );
FILL FILL_40_DFFSR_73 ( );
FILL FILL_41_DFFSR_73 ( );
FILL FILL_42_DFFSR_73 ( );
FILL FILL_43_DFFSR_73 ( );
FILL FILL_44_DFFSR_73 ( );
FILL FILL_45_DFFSR_73 ( );
FILL FILL_46_DFFSR_73 ( );
FILL FILL_47_DFFSR_73 ( );
FILL FILL_48_DFFSR_73 ( );
FILL FILL_49_DFFSR_73 ( );
FILL FILL_50_DFFSR_73 ( );
FILL FILL_0_INVX1_83 ( );
FILL FILL_1_INVX1_83 ( );
FILL FILL_2_INVX1_83 ( );
FILL FILL_3_INVX1_83 ( );
FILL FILL_4_INVX1_83 ( );
FILL FILL_0_OAI21X1_73 ( );
FILL FILL_1_OAI21X1_73 ( );
FILL FILL_2_OAI21X1_73 ( );
FILL FILL_3_OAI21X1_73 ( );
FILL FILL_4_OAI21X1_73 ( );
FILL FILL_5_OAI21X1_73 ( );
FILL FILL_6_OAI21X1_73 ( );
FILL FILL_7_OAI21X1_73 ( );
FILL FILL_8_OAI21X1_73 ( );
FILL FILL_0_NAND2X1_78 ( );
FILL FILL_1_NAND2X1_78 ( );
FILL FILL_2_NAND2X1_78 ( );
FILL FILL_3_NAND2X1_78 ( );
FILL FILL_4_NAND2X1_78 ( );
FILL FILL_5_NAND2X1_78 ( );
FILL FILL_6_NAND2X1_78 ( );
FILL FILL_0_NAND2X1_73 ( );
FILL FILL_1_NAND2X1_73 ( );
FILL FILL_2_NAND2X1_73 ( );
FILL FILL_3_NAND2X1_73 ( );
FILL FILL_4_NAND2X1_73 ( );
FILL FILL_5_NAND2X1_73 ( );
FILL FILL_6_NAND2X1_73 ( );
FILL FILL_0_NOR2X1_31 ( );
FILL FILL_1_NOR2X1_31 ( );
FILL FILL_2_NOR2X1_31 ( );
FILL FILL_3_NOR2X1_31 ( );
FILL FILL_4_NOR2X1_31 ( );
FILL FILL_5_NOR2X1_31 ( );
FILL FILL_6_NOR2X1_31 ( );
FILL FILL_0_OAI21X1_80 ( );
FILL FILL_1_OAI21X1_80 ( );
FILL FILL_2_OAI21X1_80 ( );
FILL FILL_3_OAI21X1_80 ( );
FILL FILL_4_OAI21X1_80 ( );
FILL FILL_5_OAI21X1_80 ( );
FILL FILL_6_OAI21X1_80 ( );
FILL FILL_7_OAI21X1_80 ( );
FILL FILL_8_OAI21X1_80 ( );
FILL FILL_0_INVX1_90 ( );
FILL FILL_1_INVX1_90 ( );
FILL FILL_2_INVX1_90 ( );
FILL FILL_3_INVX1_90 ( );
FILL FILL_4_INVX1_90 ( );
FILL FILL_0_INVX1_133 ( );
FILL FILL_1_INVX1_133 ( );
FILL FILL_2_INVX1_133 ( );
FILL FILL_3_INVX1_133 ( );
FILL FILL_4_INVX1_133 ( );
FILL FILL_0_OAI21X1_118 ( );
FILL FILL_1_OAI21X1_118 ( );
FILL FILL_2_OAI21X1_118 ( );
FILL FILL_3_OAI21X1_118 ( );
FILL FILL_4_OAI21X1_118 ( );
FILL FILL_5_OAI21X1_118 ( );
FILL FILL_6_OAI21X1_118 ( );
FILL FILL_7_OAI21X1_118 ( );
FILL FILL_8_OAI21X1_118 ( );
FILL FILL_0_NAND2X1_118 ( );
FILL FILL_1_NAND2X1_118 ( );
FILL FILL_2_NAND2X1_118 ( );
FILL FILL_3_NAND2X1_118 ( );
FILL FILL_4_NAND2X1_118 ( );
FILL FILL_5_NAND2X1_118 ( );
FILL FILL_6_NAND2X1_118 ( );
FILL FILL_0_BUFX2_24 ( );
FILL FILL_1_BUFX2_24 ( );
FILL FILL_2_BUFX2_24 ( );
FILL FILL_3_BUFX2_24 ( );
FILL FILL_4_BUFX2_24 ( );
FILL FILL_5_BUFX2_24 ( );
FILL FILL_6_BUFX2_24 ( );
FILL FILL_0_NAND2X1_110 ( );
FILL FILL_1_NAND2X1_110 ( );
FILL FILL_2_NAND2X1_110 ( );
FILL FILL_3_NAND2X1_110 ( );
FILL FILL_4_NAND2X1_110 ( );
FILL FILL_5_NAND2X1_110 ( );
FILL FILL_6_NAND2X1_110 ( );
FILL FILL_0_OAI21X1_110 ( );
FILL FILL_1_OAI21X1_110 ( );
FILL FILL_2_OAI21X1_110 ( );
FILL FILL_3_OAI21X1_110 ( );
FILL FILL_4_OAI21X1_110 ( );
FILL FILL_5_OAI21X1_110 ( );
FILL FILL_6_OAI21X1_110 ( );
FILL FILL_7_OAI21X1_110 ( );
FILL FILL_8_OAI21X1_110 ( );
FILL FILL_0_DFFSR_138 ( );
FILL FILL_1_DFFSR_138 ( );
FILL FILL_2_DFFSR_138 ( );
FILL FILL_3_DFFSR_138 ( );
FILL FILL_4_DFFSR_138 ( );
FILL FILL_5_DFFSR_138 ( );
FILL FILL_6_DFFSR_138 ( );
FILL FILL_7_DFFSR_138 ( );
FILL FILL_8_DFFSR_138 ( );
FILL FILL_9_DFFSR_138 ( );
FILL FILL_10_DFFSR_138 ( );
FILL FILL_11_DFFSR_138 ( );
FILL FILL_12_DFFSR_138 ( );
FILL FILL_13_DFFSR_138 ( );
FILL FILL_14_DFFSR_138 ( );
FILL FILL_15_DFFSR_138 ( );
FILL FILL_16_DFFSR_138 ( );
FILL FILL_17_DFFSR_138 ( );
FILL FILL_18_DFFSR_138 ( );
FILL FILL_19_DFFSR_138 ( );
FILL FILL_20_DFFSR_138 ( );
FILL FILL_21_DFFSR_138 ( );
FILL FILL_22_DFFSR_138 ( );
FILL FILL_23_DFFSR_138 ( );
FILL FILL_24_DFFSR_138 ( );
FILL FILL_25_DFFSR_138 ( );
FILL FILL_26_DFFSR_138 ( );
FILL FILL_27_DFFSR_138 ( );
FILL FILL_28_DFFSR_138 ( );
FILL FILL_29_DFFSR_138 ( );
FILL FILL_30_DFFSR_138 ( );
FILL FILL_31_DFFSR_138 ( );
FILL FILL_32_DFFSR_138 ( );
FILL FILL_33_DFFSR_138 ( );
FILL FILL_34_DFFSR_138 ( );
FILL FILL_35_DFFSR_138 ( );
FILL FILL_36_DFFSR_138 ( );
FILL FILL_37_DFFSR_138 ( );
FILL FILL_38_DFFSR_138 ( );
FILL FILL_39_DFFSR_138 ( );
FILL FILL_40_DFFSR_138 ( );
FILL FILL_41_DFFSR_138 ( );
FILL FILL_42_DFFSR_138 ( );
FILL FILL_43_DFFSR_138 ( );
FILL FILL_44_DFFSR_138 ( );
FILL FILL_45_DFFSR_138 ( );
FILL FILL_46_DFFSR_138 ( );
FILL FILL_47_DFFSR_138 ( );
FILL FILL_48_DFFSR_138 ( );
FILL FILL_49_DFFSR_138 ( );
FILL FILL_50_DFFSR_138 ( );
FILL FILL_0_OAI21X1_24 ( );
FILL FILL_1_OAI21X1_24 ( );
FILL FILL_2_OAI21X1_24 ( );
FILL FILL_3_OAI21X1_24 ( );
FILL FILL_4_OAI21X1_24 ( );
FILL FILL_5_OAI21X1_24 ( );
FILL FILL_6_OAI21X1_24 ( );
FILL FILL_7_OAI21X1_24 ( );
FILL FILL_8_OAI21X1_24 ( );
FILL FILL_0_INVX1_27 ( );
FILL FILL_1_INVX1_27 ( );
FILL FILL_2_INVX1_27 ( );
FILL FILL_3_INVX1_27 ( );
FILL FILL_4_INVX1_27 ( );
FILL FILL_0_NAND2X1_40 ( );
FILL FILL_1_NAND2X1_40 ( );
FILL FILL_2_NAND2X1_40 ( );
FILL FILL_3_NAND2X1_40 ( );
FILL FILL_4_NAND2X1_40 ( );
FILL FILL_5_NAND2X1_40 ( );
FILL FILL_6_NAND2X1_40 ( );
FILL FILL_0_NOR2X1_26 ( );
FILL FILL_1_NOR2X1_26 ( );
FILL FILL_2_NOR2X1_26 ( );
FILL FILL_3_NOR2X1_26 ( );
FILL FILL_4_NOR2X1_26 ( );
FILL FILL_5_NOR2X1_26 ( );
FILL FILL_6_NOR2X1_26 ( );
FILL FILL_0_DFFSR_50 ( );
FILL FILL_1_DFFSR_50 ( );
FILL FILL_2_DFFSR_50 ( );
FILL FILL_3_DFFSR_50 ( );
FILL FILL_4_DFFSR_50 ( );
FILL FILL_5_DFFSR_50 ( );
FILL FILL_6_DFFSR_50 ( );
FILL FILL_7_DFFSR_50 ( );
FILL FILL_8_DFFSR_50 ( );
FILL FILL_9_DFFSR_50 ( );
FILL FILL_10_DFFSR_50 ( );
FILL FILL_11_DFFSR_50 ( );
FILL FILL_12_DFFSR_50 ( );
FILL FILL_13_DFFSR_50 ( );
FILL FILL_14_DFFSR_50 ( );
FILL FILL_15_DFFSR_50 ( );
FILL FILL_16_DFFSR_50 ( );
FILL FILL_17_DFFSR_50 ( );
FILL FILL_18_DFFSR_50 ( );
FILL FILL_19_DFFSR_50 ( );
FILL FILL_20_DFFSR_50 ( );
FILL FILL_21_DFFSR_50 ( );
FILL FILL_22_DFFSR_50 ( );
FILL FILL_23_DFFSR_50 ( );
FILL FILL_24_DFFSR_50 ( );
FILL FILL_25_DFFSR_50 ( );
FILL FILL_26_DFFSR_50 ( );
FILL FILL_27_DFFSR_50 ( );
FILL FILL_28_DFFSR_50 ( );
FILL FILL_29_DFFSR_50 ( );
FILL FILL_30_DFFSR_50 ( );
FILL FILL_31_DFFSR_50 ( );
FILL FILL_32_DFFSR_50 ( );
FILL FILL_33_DFFSR_50 ( );
FILL FILL_34_DFFSR_50 ( );
FILL FILL_35_DFFSR_50 ( );
FILL FILL_36_DFFSR_50 ( );
FILL FILL_37_DFFSR_50 ( );
FILL FILL_38_DFFSR_50 ( );
FILL FILL_39_DFFSR_50 ( );
FILL FILL_40_DFFSR_50 ( );
FILL FILL_41_DFFSR_50 ( );
FILL FILL_42_DFFSR_50 ( );
FILL FILL_43_DFFSR_50 ( );
FILL FILL_44_DFFSR_50 ( );
FILL FILL_45_DFFSR_50 ( );
FILL FILL_46_DFFSR_50 ( );
FILL FILL_47_DFFSR_50 ( );
FILL FILL_48_DFFSR_50 ( );
FILL FILL_49_DFFSR_50 ( );
FILL FILL_50_DFFSR_50 ( );
FILL FILL_51_DFFSR_50 ( );
FILL FILL_0_OAI22X1_6 ( );
FILL FILL_1_OAI22X1_6 ( );
FILL FILL_2_OAI22X1_6 ( );
FILL FILL_3_OAI22X1_6 ( );
FILL FILL_4_OAI22X1_6 ( );
FILL FILL_5_OAI22X1_6 ( );
FILL FILL_6_OAI22X1_6 ( );
FILL FILL_7_OAI22X1_6 ( );
FILL FILL_8_OAI22X1_6 ( );
FILL FILL_9_OAI22X1_6 ( );
FILL FILL_10_OAI22X1_6 ( );
FILL FILL_0_OAI22X1_21 ( );
FILL FILL_1_OAI22X1_21 ( );
FILL FILL_2_OAI22X1_21 ( );
FILL FILL_3_OAI22X1_21 ( );
FILL FILL_4_OAI22X1_21 ( );
FILL FILL_5_OAI22X1_21 ( );
FILL FILL_6_OAI22X1_21 ( );
FILL FILL_7_OAI22X1_21 ( );
FILL FILL_8_OAI22X1_21 ( );
FILL FILL_9_OAI22X1_21 ( );
FILL FILL_10_OAI22X1_21 ( );
FILL FILL_0_INVX1_272 ( );
FILL FILL_1_INVX1_272 ( );
FILL FILL_2_INVX1_272 ( );
FILL FILL_3_INVX1_272 ( );
FILL FILL_0_NAND2X1_49 ( );
FILL FILL_1_NAND2X1_49 ( );
FILL FILL_2_NAND2X1_49 ( );
FILL FILL_3_NAND2X1_49 ( );
FILL FILL_4_NAND2X1_49 ( );
FILL FILL_5_NAND2X1_49 ( );
FILL FILL_6_NAND2X1_49 ( );
FILL FILL_0_DFFSR_49 ( );
FILL FILL_1_DFFSR_49 ( );
FILL FILL_2_DFFSR_49 ( );
FILL FILL_3_DFFSR_49 ( );
FILL FILL_4_DFFSR_49 ( );
FILL FILL_5_DFFSR_49 ( );
FILL FILL_6_DFFSR_49 ( );
FILL FILL_7_DFFSR_49 ( );
FILL FILL_8_DFFSR_49 ( );
FILL FILL_9_DFFSR_49 ( );
FILL FILL_10_DFFSR_49 ( );
FILL FILL_11_DFFSR_49 ( );
FILL FILL_12_DFFSR_49 ( );
FILL FILL_13_DFFSR_49 ( );
FILL FILL_14_DFFSR_49 ( );
FILL FILL_15_DFFSR_49 ( );
FILL FILL_16_DFFSR_49 ( );
FILL FILL_17_DFFSR_49 ( );
FILL FILL_18_DFFSR_49 ( );
FILL FILL_19_DFFSR_49 ( );
FILL FILL_20_DFFSR_49 ( );
FILL FILL_21_DFFSR_49 ( );
FILL FILL_22_DFFSR_49 ( );
FILL FILL_23_DFFSR_49 ( );
FILL FILL_24_DFFSR_49 ( );
FILL FILL_25_DFFSR_49 ( );
FILL FILL_26_DFFSR_49 ( );
FILL FILL_27_DFFSR_49 ( );
FILL FILL_28_DFFSR_49 ( );
FILL FILL_29_DFFSR_49 ( );
FILL FILL_30_DFFSR_49 ( );
FILL FILL_31_DFFSR_49 ( );
FILL FILL_32_DFFSR_49 ( );
FILL FILL_33_DFFSR_49 ( );
FILL FILL_34_DFFSR_49 ( );
FILL FILL_35_DFFSR_49 ( );
FILL FILL_36_DFFSR_49 ( );
FILL FILL_37_DFFSR_49 ( );
FILL FILL_38_DFFSR_49 ( );
FILL FILL_39_DFFSR_49 ( );
FILL FILL_40_DFFSR_49 ( );
FILL FILL_41_DFFSR_49 ( );
FILL FILL_42_DFFSR_49 ( );
FILL FILL_43_DFFSR_49 ( );
FILL FILL_44_DFFSR_49 ( );
FILL FILL_45_DFFSR_49 ( );
FILL FILL_46_DFFSR_49 ( );
FILL FILL_47_DFFSR_49 ( );
FILL FILL_48_DFFSR_49 ( );
FILL FILL_49_DFFSR_49 ( );
FILL FILL_50_DFFSR_49 ( );
FILL FILL_0_INVX1_56 ( );
FILL FILL_1_INVX1_56 ( );
FILL FILL_2_INVX1_56 ( );
FILL FILL_3_INVX1_56 ( );
FILL FILL_0_OAI21X1_49 ( );
FILL FILL_1_OAI21X1_49 ( );
FILL FILL_2_OAI21X1_49 ( );
FILL FILL_3_OAI21X1_49 ( );
FILL FILL_4_OAI21X1_49 ( );
FILL FILL_5_OAI21X1_49 ( );
FILL FILL_6_OAI21X1_49 ( );
FILL FILL_7_OAI21X1_49 ( );
FILL FILL_8_OAI21X1_49 ( );
FILL FILL_9_OAI21X1_49 ( );
FILL FILL_0_OAI21X1_57 ( );
FILL FILL_1_OAI21X1_57 ( );
FILL FILL_2_OAI21X1_57 ( );
FILL FILL_3_OAI21X1_57 ( );
FILL FILL_4_OAI21X1_57 ( );
FILL FILL_5_OAI21X1_57 ( );
FILL FILL_6_OAI21X1_57 ( );
FILL FILL_7_OAI21X1_57 ( );
FILL FILL_8_OAI21X1_57 ( );
FILL FILL_9_OAI21X1_57 ( );
FILL FILL_0_INVX1_65 ( );
FILL FILL_1_INVX1_65 ( );
FILL FILL_2_INVX1_65 ( );
FILL FILL_3_INVX1_65 ( );
FILL FILL_0_INVX1_297 ( );
FILL FILL_1_INVX1_297 ( );
FILL FILL_2_INVX1_297 ( );
FILL FILL_3_INVX1_297 ( );
FILL FILL_4_INVX1_297 ( );
FILL FILL_0_NAND2X1_13 ( );
FILL FILL_1_NAND2X1_13 ( );
FILL FILL_2_NAND2X1_13 ( );
FILL FILL_3_NAND2X1_13 ( );
FILL FILL_4_NAND2X1_13 ( );
FILL FILL_5_NAND2X1_13 ( );
FILL FILL_6_NAND2X1_13 ( );
FILL FILL_0_INVX1_410 ( );
FILL FILL_1_INVX1_410 ( );
FILL FILL_2_INVX1_410 ( );
FILL FILL_3_INVX1_410 ( );
FILL FILL_0_DFFPOSX1_5 ( );
FILL FILL_1_DFFPOSX1_5 ( );
FILL FILL_2_DFFPOSX1_5 ( );
FILL FILL_3_DFFPOSX1_5 ( );
FILL FILL_4_DFFPOSX1_5 ( );
FILL FILL_5_DFFPOSX1_5 ( );
FILL FILL_6_DFFPOSX1_5 ( );
FILL FILL_7_DFFPOSX1_5 ( );
FILL FILL_8_DFFPOSX1_5 ( );
FILL FILL_9_DFFPOSX1_5 ( );
FILL FILL_10_DFFPOSX1_5 ( );
FILL FILL_11_DFFPOSX1_5 ( );
FILL FILL_12_DFFPOSX1_5 ( );
FILL FILL_13_DFFPOSX1_5 ( );
FILL FILL_14_DFFPOSX1_5 ( );
FILL FILL_15_DFFPOSX1_5 ( );
FILL FILL_16_DFFPOSX1_5 ( );
FILL FILL_17_DFFPOSX1_5 ( );
FILL FILL_18_DFFPOSX1_5 ( );
FILL FILL_19_DFFPOSX1_5 ( );
FILL FILL_20_DFFPOSX1_5 ( );
FILL FILL_21_DFFPOSX1_5 ( );
FILL FILL_22_DFFPOSX1_5 ( );
FILL FILL_23_DFFPOSX1_5 ( );
FILL FILL_24_DFFPOSX1_5 ( );
FILL FILL_25_DFFPOSX1_5 ( );
FILL FILL_26_DFFPOSX1_5 ( );
FILL FILL_27_DFFPOSX1_5 ( );
FILL FILL_0_NAND2X1_259 ( );
FILL FILL_1_NAND2X1_259 ( );
FILL FILL_2_NAND2X1_259 ( );
FILL FILL_3_NAND2X1_259 ( );
FILL FILL_4_NAND2X1_259 ( );
FILL FILL_5_NAND2X1_259 ( );
FILL FILL_6_NAND2X1_259 ( );
FILL FILL_0_INVX1_135 ( );
FILL FILL_1_INVX1_135 ( );
FILL FILL_2_INVX1_135 ( );
FILL FILL_3_INVX1_135 ( );
FILL FILL_4_INVX1_135 ( );
FILL FILL_0_DFFSR_120 ( );
FILL FILL_1_DFFSR_120 ( );
FILL FILL_2_DFFSR_120 ( );
FILL FILL_3_DFFSR_120 ( );
FILL FILL_4_DFFSR_120 ( );
FILL FILL_5_DFFSR_120 ( );
FILL FILL_6_DFFSR_120 ( );
FILL FILL_7_DFFSR_120 ( );
FILL FILL_8_DFFSR_120 ( );
FILL FILL_9_DFFSR_120 ( );
FILL FILL_10_DFFSR_120 ( );
FILL FILL_11_DFFSR_120 ( );
FILL FILL_12_DFFSR_120 ( );
FILL FILL_13_DFFSR_120 ( );
FILL FILL_14_DFFSR_120 ( );
FILL FILL_15_DFFSR_120 ( );
FILL FILL_16_DFFSR_120 ( );
FILL FILL_17_DFFSR_120 ( );
FILL FILL_18_DFFSR_120 ( );
FILL FILL_19_DFFSR_120 ( );
FILL FILL_20_DFFSR_120 ( );
FILL FILL_21_DFFSR_120 ( );
FILL FILL_22_DFFSR_120 ( );
FILL FILL_23_DFFSR_120 ( );
FILL FILL_24_DFFSR_120 ( );
FILL FILL_25_DFFSR_120 ( );
FILL FILL_26_DFFSR_120 ( );
FILL FILL_27_DFFSR_120 ( );
FILL FILL_28_DFFSR_120 ( );
FILL FILL_29_DFFSR_120 ( );
FILL FILL_30_DFFSR_120 ( );
FILL FILL_31_DFFSR_120 ( );
FILL FILL_32_DFFSR_120 ( );
FILL FILL_33_DFFSR_120 ( );
FILL FILL_34_DFFSR_120 ( );
FILL FILL_35_DFFSR_120 ( );
FILL FILL_36_DFFSR_120 ( );
FILL FILL_37_DFFSR_120 ( );
FILL FILL_38_DFFSR_120 ( );
FILL FILL_39_DFFSR_120 ( );
FILL FILL_40_DFFSR_120 ( );
FILL FILL_41_DFFSR_120 ( );
FILL FILL_42_DFFSR_120 ( );
FILL FILL_43_DFFSR_120 ( );
FILL FILL_44_DFFSR_120 ( );
FILL FILL_45_DFFSR_120 ( );
FILL FILL_46_DFFSR_120 ( );
FILL FILL_47_DFFSR_120 ( );
FILL FILL_48_DFFSR_120 ( );
FILL FILL_49_DFFSR_120 ( );
FILL FILL_50_DFFSR_120 ( );
FILL FILL_0_NAND2X1_94 ( );
FILL FILL_1_NAND2X1_94 ( );
FILL FILL_2_NAND2X1_94 ( );
FILL FILL_3_NAND2X1_94 ( );
FILL FILL_4_NAND2X1_94 ( );
FILL FILL_5_NAND2X1_94 ( );
FILL FILL_6_NAND2X1_94 ( );
FILL FILL_0_OAI21X1_94 ( );
FILL FILL_1_OAI21X1_94 ( );
FILL FILL_2_OAI21X1_94 ( );
FILL FILL_3_OAI21X1_94 ( );
FILL FILL_4_OAI21X1_94 ( );
FILL FILL_5_OAI21X1_94 ( );
FILL FILL_6_OAI21X1_94 ( );
FILL FILL_7_OAI21X1_94 ( );
FILL FILL_8_OAI21X1_94 ( );
FILL FILL_0_INVX1_106 ( );
FILL FILL_1_INVX1_106 ( );
FILL FILL_2_INVX1_106 ( );
FILL FILL_3_INVX1_106 ( );
FILL FILL_4_INVX1_106 ( );
FILL FILL_0_OAI22X1_44 ( );
FILL FILL_1_OAI22X1_44 ( );
FILL FILL_2_OAI22X1_44 ( );
FILL FILL_3_OAI22X1_44 ( );
FILL FILL_4_OAI22X1_44 ( );
FILL FILL_5_OAI22X1_44 ( );
FILL FILL_6_OAI22X1_44 ( );
FILL FILL_7_OAI22X1_44 ( );
FILL FILL_8_OAI22X1_44 ( );
FILL FILL_9_OAI22X1_44 ( );
FILL FILL_10_OAI22X1_44 ( );
FILL FILL_11_OAI22X1_44 ( );
FILL FILL_0_INVX1_100 ( );
FILL FILL_1_INVX1_100 ( );
FILL FILL_2_INVX1_100 ( );
FILL FILL_3_INVX1_100 ( );
FILL FILL_0_DFFSR_118 ( );
FILL FILL_1_DFFSR_118 ( );
FILL FILL_2_DFFSR_118 ( );
FILL FILL_3_DFFSR_118 ( );
FILL FILL_4_DFFSR_118 ( );
FILL FILL_5_DFFSR_118 ( );
FILL FILL_6_DFFSR_118 ( );
FILL FILL_7_DFFSR_118 ( );
FILL FILL_8_DFFSR_118 ( );
FILL FILL_9_DFFSR_118 ( );
FILL FILL_10_DFFSR_118 ( );
FILL FILL_11_DFFSR_118 ( );
FILL FILL_12_DFFSR_118 ( );
FILL FILL_13_DFFSR_118 ( );
FILL FILL_14_DFFSR_118 ( );
FILL FILL_15_DFFSR_118 ( );
FILL FILL_16_DFFSR_118 ( );
FILL FILL_17_DFFSR_118 ( );
FILL FILL_18_DFFSR_118 ( );
FILL FILL_19_DFFSR_118 ( );
FILL FILL_20_DFFSR_118 ( );
FILL FILL_21_DFFSR_118 ( );
FILL FILL_22_DFFSR_118 ( );
FILL FILL_23_DFFSR_118 ( );
FILL FILL_24_DFFSR_118 ( );
FILL FILL_25_DFFSR_118 ( );
FILL FILL_26_DFFSR_118 ( );
FILL FILL_27_DFFSR_118 ( );
FILL FILL_28_DFFSR_118 ( );
FILL FILL_29_DFFSR_118 ( );
FILL FILL_30_DFFSR_118 ( );
FILL FILL_31_DFFSR_118 ( );
FILL FILL_32_DFFSR_118 ( );
FILL FILL_33_DFFSR_118 ( );
FILL FILL_34_DFFSR_118 ( );
FILL FILL_35_DFFSR_118 ( );
FILL FILL_36_DFFSR_118 ( );
FILL FILL_37_DFFSR_118 ( );
FILL FILL_38_DFFSR_118 ( );
FILL FILL_39_DFFSR_118 ( );
FILL FILL_40_DFFSR_118 ( );
FILL FILL_41_DFFSR_118 ( );
FILL FILL_42_DFFSR_118 ( );
FILL FILL_43_DFFSR_118 ( );
FILL FILL_44_DFFSR_118 ( );
FILL FILL_45_DFFSR_118 ( );
FILL FILL_46_DFFSR_118 ( );
FILL FILL_47_DFFSR_118 ( );
FILL FILL_48_DFFSR_118 ( );
FILL FILL_49_DFFSR_118 ( );
FILL FILL_50_DFFSR_118 ( );
FILL FILL_51_DFFSR_118 ( );
FILL FILL_0_XOR2X1_10 ( );
FILL FILL_1_XOR2X1_10 ( );
FILL FILL_2_XOR2X1_10 ( );
FILL FILL_3_XOR2X1_10 ( );
FILL FILL_4_XOR2X1_10 ( );
FILL FILL_5_XOR2X1_10 ( );
FILL FILL_6_XOR2X1_10 ( );
FILL FILL_7_XOR2X1_10 ( );
FILL FILL_8_XOR2X1_10 ( );
FILL FILL_9_XOR2X1_10 ( );
FILL FILL_10_XOR2X1_10 ( );
FILL FILL_11_XOR2X1_10 ( );
FILL FILL_12_XOR2X1_10 ( );
FILL FILL_13_XOR2X1_10 ( );
FILL FILL_14_XOR2X1_10 ( );
FILL FILL_15_XOR2X1_10 ( );
FILL FILL_0_NAND2X1_272 ( );
FILL FILL_1_NAND2X1_272 ( );
FILL FILL_2_NAND2X1_272 ( );
FILL FILL_3_NAND2X1_272 ( );
FILL FILL_4_NAND2X1_272 ( );
FILL FILL_5_NAND2X1_272 ( );
FILL FILL_6_NAND2X1_272 ( );
FILL FILL_0_OAI21X1_260 ( );
FILL FILL_1_OAI21X1_260 ( );
FILL FILL_2_OAI21X1_260 ( );
FILL FILL_3_OAI21X1_260 ( );
FILL FILL_4_OAI21X1_260 ( );
FILL FILL_5_OAI21X1_260 ( );
FILL FILL_6_OAI21X1_260 ( );
FILL FILL_7_OAI21X1_260 ( );
FILL FILL_8_OAI21X1_260 ( );
FILL FILL_9_OAI21X1_260 ( );
FILL FILL_0_DFFPOSX1_22 ( );
FILL FILL_1_DFFPOSX1_22 ( );
FILL FILL_2_DFFPOSX1_22 ( );
FILL FILL_3_DFFPOSX1_22 ( );
FILL FILL_4_DFFPOSX1_22 ( );
FILL FILL_5_DFFPOSX1_22 ( );
FILL FILL_6_DFFPOSX1_22 ( );
FILL FILL_7_DFFPOSX1_22 ( );
FILL FILL_8_DFFPOSX1_22 ( );
FILL FILL_9_DFFPOSX1_22 ( );
FILL FILL_10_DFFPOSX1_22 ( );
FILL FILL_11_DFFPOSX1_22 ( );
FILL FILL_12_DFFPOSX1_22 ( );
FILL FILL_13_DFFPOSX1_22 ( );
FILL FILL_14_DFFPOSX1_22 ( );
FILL FILL_15_DFFPOSX1_22 ( );
FILL FILL_16_DFFPOSX1_22 ( );
FILL FILL_17_DFFPOSX1_22 ( );
FILL FILL_18_DFFPOSX1_22 ( );
FILL FILL_19_DFFPOSX1_22 ( );
FILL FILL_20_DFFPOSX1_22 ( );
FILL FILL_21_DFFPOSX1_22 ( );
FILL FILL_22_DFFPOSX1_22 ( );
FILL FILL_23_DFFPOSX1_22 ( );
FILL FILL_24_DFFPOSX1_22 ( );
FILL FILL_25_DFFPOSX1_22 ( );
FILL FILL_26_DFFPOSX1_22 ( );
FILL FILL_27_DFFPOSX1_22 ( );
FILL FILL_0_NAND2X1_48 ( );
FILL FILL_1_NAND2X1_48 ( );
FILL FILL_2_NAND2X1_48 ( );
FILL FILL_3_NAND2X1_48 ( );
FILL FILL_4_NAND2X1_48 ( );
FILL FILL_5_NAND2X1_48 ( );
FILL FILL_6_NAND2X1_48 ( );
FILL FILL_0_INVX1_324 ( );
FILL FILL_1_INVX1_324 ( );
FILL FILL_2_INVX1_324 ( );
FILL FILL_3_INVX1_324 ( );
FILL FILL_4_INVX1_324 ( );
FILL FILL_0_OAI22X1_34 ( );
FILL FILL_1_OAI22X1_34 ( );
FILL FILL_2_OAI22X1_34 ( );
FILL FILL_3_OAI22X1_34 ( );
FILL FILL_4_OAI22X1_34 ( );
FILL FILL_5_OAI22X1_34 ( );
FILL FILL_6_OAI22X1_34 ( );
FILL FILL_7_OAI22X1_34 ( );
FILL FILL_8_OAI22X1_34 ( );
FILL FILL_9_OAI22X1_34 ( );
FILL FILL_10_OAI22X1_34 ( );
FILL FILL_0_INVX1_275 ( );
FILL FILL_1_INVX1_275 ( );
FILL FILL_2_INVX1_275 ( );
FILL FILL_3_INVX1_275 ( );
FILL FILL_0_INVX1_72 ( );
FILL FILL_1_INVX1_72 ( );
FILL FILL_2_INVX1_72 ( );
FILL FILL_3_INVX1_72 ( );
FILL FILL_0_INVX1_327 ( );
FILL FILL_1_INVX1_327 ( );
FILL FILL_2_INVX1_327 ( );
FILL FILL_3_INVX1_327 ( );
FILL FILL_4_INVX1_327 ( );
FILL FILL_0_NOR2X1_20 ( );
FILL FILL_1_NOR2X1_20 ( );
FILL FILL_2_NOR2X1_20 ( );
FILL FILL_3_NOR2X1_20 ( );
FILL FILL_4_NOR2X1_20 ( );
FILL FILL_5_NOR2X1_20 ( );
FILL FILL_6_NOR2X1_20 ( );
FILL FILL_0_OAI22X1_22 ( );
FILL FILL_1_OAI22X1_22 ( );
FILL FILL_2_OAI22X1_22 ( );
FILL FILL_3_OAI22X1_22 ( );
FILL FILL_4_OAI22X1_22 ( );
FILL FILL_5_OAI22X1_22 ( );
FILL FILL_6_OAI22X1_22 ( );
FILL FILL_7_OAI22X1_22 ( );
FILL FILL_8_OAI22X1_22 ( );
FILL FILL_9_OAI22X1_22 ( );
FILL FILL_10_OAI22X1_22 ( );
FILL FILL_0_DFFSR_64 ( );
FILL FILL_1_DFFSR_64 ( );
FILL FILL_2_DFFSR_64 ( );
FILL FILL_3_DFFSR_64 ( );
FILL FILL_4_DFFSR_64 ( );
FILL FILL_5_DFFSR_64 ( );
FILL FILL_6_DFFSR_64 ( );
FILL FILL_7_DFFSR_64 ( );
FILL FILL_8_DFFSR_64 ( );
FILL FILL_9_DFFSR_64 ( );
FILL FILL_10_DFFSR_64 ( );
FILL FILL_11_DFFSR_64 ( );
FILL FILL_12_DFFSR_64 ( );
FILL FILL_13_DFFSR_64 ( );
FILL FILL_14_DFFSR_64 ( );
FILL FILL_15_DFFSR_64 ( );
FILL FILL_16_DFFSR_64 ( );
FILL FILL_17_DFFSR_64 ( );
FILL FILL_18_DFFSR_64 ( );
FILL FILL_19_DFFSR_64 ( );
FILL FILL_20_DFFSR_64 ( );
FILL FILL_21_DFFSR_64 ( );
FILL FILL_22_DFFSR_64 ( );
FILL FILL_23_DFFSR_64 ( );
FILL FILL_24_DFFSR_64 ( );
FILL FILL_25_DFFSR_64 ( );
FILL FILL_26_DFFSR_64 ( );
FILL FILL_27_DFFSR_64 ( );
FILL FILL_28_DFFSR_64 ( );
FILL FILL_29_DFFSR_64 ( );
FILL FILL_30_DFFSR_64 ( );
FILL FILL_31_DFFSR_64 ( );
FILL FILL_32_DFFSR_64 ( );
FILL FILL_33_DFFSR_64 ( );
FILL FILL_34_DFFSR_64 ( );
FILL FILL_35_DFFSR_64 ( );
FILL FILL_36_DFFSR_64 ( );
FILL FILL_37_DFFSR_64 ( );
FILL FILL_38_DFFSR_64 ( );
FILL FILL_39_DFFSR_64 ( );
FILL FILL_40_DFFSR_64 ( );
FILL FILL_41_DFFSR_64 ( );
FILL FILL_42_DFFSR_64 ( );
FILL FILL_43_DFFSR_64 ( );
FILL FILL_44_DFFSR_64 ( );
FILL FILL_45_DFFSR_64 ( );
FILL FILL_46_DFFSR_64 ( );
FILL FILL_47_DFFSR_64 ( );
FILL FILL_48_DFFSR_64 ( );
FILL FILL_49_DFFSR_64 ( );
FILL FILL_50_DFFSR_64 ( );
FILL FILL_0_NAND2X1_170 ( );
FILL FILL_1_NAND2X1_170 ( );
FILL FILL_2_NAND2X1_170 ( );
FILL FILL_3_NAND2X1_170 ( );
FILL FILL_4_NAND2X1_170 ( );
FILL FILL_5_NAND2X1_170 ( );
FILL FILL_6_NAND2X1_170 ( );
FILL FILL_0_INVX1_300 ( );
FILL FILL_1_INVX1_300 ( );
FILL FILL_2_INVX1_300 ( );
FILL FILL_3_INVX1_300 ( );
FILL FILL_4_INVX1_300 ( );
FILL FILL_0_INVX1_13 ( );
FILL FILL_1_INVX1_13 ( );
FILL FILL_2_INVX1_13 ( );
FILL FILL_3_INVX1_13 ( );
FILL FILL_0_OAI21X1_11 ( );
FILL FILL_1_OAI21X1_11 ( );
FILL FILL_2_OAI21X1_11 ( );
FILL FILL_3_OAI21X1_11 ( );
FILL FILL_4_OAI21X1_11 ( );
FILL FILL_5_OAI21X1_11 ( );
FILL FILL_6_OAI21X1_11 ( );
FILL FILL_7_OAI21X1_11 ( );
FILL FILL_8_OAI21X1_11 ( );
FILL FILL_9_OAI21X1_11 ( );
FILL FILL_0_DFFSR_11 ( );
FILL FILL_1_DFFSR_11 ( );
FILL FILL_2_DFFSR_11 ( );
FILL FILL_3_DFFSR_11 ( );
FILL FILL_4_DFFSR_11 ( );
FILL FILL_5_DFFSR_11 ( );
FILL FILL_6_DFFSR_11 ( );
FILL FILL_7_DFFSR_11 ( );
FILL FILL_8_DFFSR_11 ( );
FILL FILL_9_DFFSR_11 ( );
FILL FILL_10_DFFSR_11 ( );
FILL FILL_11_DFFSR_11 ( );
FILL FILL_12_DFFSR_11 ( );
FILL FILL_13_DFFSR_11 ( );
FILL FILL_14_DFFSR_11 ( );
FILL FILL_15_DFFSR_11 ( );
FILL FILL_16_DFFSR_11 ( );
FILL FILL_17_DFFSR_11 ( );
FILL FILL_18_DFFSR_11 ( );
FILL FILL_19_DFFSR_11 ( );
FILL FILL_20_DFFSR_11 ( );
FILL FILL_21_DFFSR_11 ( );
FILL FILL_22_DFFSR_11 ( );
FILL FILL_23_DFFSR_11 ( );
FILL FILL_24_DFFSR_11 ( );
FILL FILL_25_DFFSR_11 ( );
FILL FILL_26_DFFSR_11 ( );
FILL FILL_27_DFFSR_11 ( );
FILL FILL_28_DFFSR_11 ( );
FILL FILL_29_DFFSR_11 ( );
FILL FILL_30_DFFSR_11 ( );
FILL FILL_31_DFFSR_11 ( );
FILL FILL_32_DFFSR_11 ( );
FILL FILL_33_DFFSR_11 ( );
FILL FILL_34_DFFSR_11 ( );
FILL FILL_35_DFFSR_11 ( );
FILL FILL_36_DFFSR_11 ( );
FILL FILL_37_DFFSR_11 ( );
FILL FILL_38_DFFSR_11 ( );
FILL FILL_39_DFFSR_11 ( );
FILL FILL_40_DFFSR_11 ( );
FILL FILL_41_DFFSR_11 ( );
FILL FILL_42_DFFSR_11 ( );
FILL FILL_43_DFFSR_11 ( );
FILL FILL_44_DFFSR_11 ( );
FILL FILL_45_DFFSR_11 ( );
FILL FILL_46_DFFSR_11 ( );
FILL FILL_47_DFFSR_11 ( );
FILL FILL_48_DFFSR_11 ( );
FILL FILL_49_DFFSR_11 ( );
FILL FILL_50_DFFSR_11 ( );
FILL FILL_0_DFFSR_187 ( );
FILL FILL_1_DFFSR_187 ( );
FILL FILL_2_DFFSR_187 ( );
FILL FILL_3_DFFSR_187 ( );
FILL FILL_4_DFFSR_187 ( );
FILL FILL_5_DFFSR_187 ( );
FILL FILL_6_DFFSR_187 ( );
FILL FILL_7_DFFSR_187 ( );
FILL FILL_8_DFFSR_187 ( );
FILL FILL_9_DFFSR_187 ( );
FILL FILL_10_DFFSR_187 ( );
FILL FILL_11_DFFSR_187 ( );
FILL FILL_12_DFFSR_187 ( );
FILL FILL_13_DFFSR_187 ( );
FILL FILL_14_DFFSR_187 ( );
FILL FILL_15_DFFSR_187 ( );
FILL FILL_16_DFFSR_187 ( );
FILL FILL_17_DFFSR_187 ( );
FILL FILL_18_DFFSR_187 ( );
FILL FILL_19_DFFSR_187 ( );
FILL FILL_20_DFFSR_187 ( );
FILL FILL_21_DFFSR_187 ( );
FILL FILL_22_DFFSR_187 ( );
FILL FILL_23_DFFSR_187 ( );
FILL FILL_24_DFFSR_187 ( );
FILL FILL_25_DFFSR_187 ( );
FILL FILL_26_DFFSR_187 ( );
FILL FILL_27_DFFSR_187 ( );
FILL FILL_28_DFFSR_187 ( );
FILL FILL_29_DFFSR_187 ( );
FILL FILL_30_DFFSR_187 ( );
FILL FILL_31_DFFSR_187 ( );
FILL FILL_32_DFFSR_187 ( );
FILL FILL_33_DFFSR_187 ( );
FILL FILL_34_DFFSR_187 ( );
FILL FILL_35_DFFSR_187 ( );
FILL FILL_36_DFFSR_187 ( );
FILL FILL_37_DFFSR_187 ( );
FILL FILL_38_DFFSR_187 ( );
FILL FILL_39_DFFSR_187 ( );
FILL FILL_40_DFFSR_187 ( );
FILL FILL_41_DFFSR_187 ( );
FILL FILL_42_DFFSR_187 ( );
FILL FILL_43_DFFSR_187 ( );
FILL FILL_44_DFFSR_187 ( );
FILL FILL_45_DFFSR_187 ( );
FILL FILL_46_DFFSR_187 ( );
FILL FILL_47_DFFSR_187 ( );
FILL FILL_48_DFFSR_187 ( );
FILL FILL_49_DFFSR_187 ( );
FILL FILL_50_DFFSR_187 ( );
FILL FILL_0_BUFX2_16 ( );
FILL FILL_1_BUFX2_16 ( );
FILL FILL_2_BUFX2_16 ( );
FILL FILL_3_BUFX2_16 ( );
FILL FILL_4_BUFX2_16 ( );
FILL FILL_5_BUFX2_16 ( );
FILL FILL_6_BUFX2_16 ( );
FILL FILL_0_OAI21X1_120 ( );
FILL FILL_1_OAI21X1_120 ( );
FILL FILL_2_OAI21X1_120 ( );
FILL FILL_3_OAI21X1_120 ( );
FILL FILL_4_OAI21X1_120 ( );
FILL FILL_5_OAI21X1_120 ( );
FILL FILL_6_OAI21X1_120 ( );
FILL FILL_7_OAI21X1_120 ( );
FILL FILL_8_OAI21X1_120 ( );
FILL FILL_0_BUFX2_15 ( );
FILL FILL_1_BUFX2_15 ( );
FILL FILL_2_BUFX2_15 ( );
FILL FILL_3_BUFX2_15 ( );
FILL FILL_4_BUFX2_15 ( );
FILL FILL_5_BUFX2_15 ( );
FILL FILL_6_BUFX2_15 ( );
FILL FILL_0_INVX1_126 ( );
FILL FILL_1_INVX1_126 ( );
FILL FILL_2_INVX1_126 ( );
FILL FILL_3_INVX1_126 ( );
FILL FILL_4_INVX1_126 ( );
FILL FILL_0_NAND2X1_120 ( );
FILL FILL_1_NAND2X1_120 ( );
FILL FILL_2_NAND2X1_120 ( );
FILL FILL_3_NAND2X1_120 ( );
FILL FILL_4_NAND2X1_120 ( );
FILL FILL_5_NAND2X1_120 ( );
FILL FILL_6_NAND2X1_120 ( );
FILL FILL_0_DFFSR_94 ( );
FILL FILL_1_DFFSR_94 ( );
FILL FILL_2_DFFSR_94 ( );
FILL FILL_3_DFFSR_94 ( );
FILL FILL_4_DFFSR_94 ( );
FILL FILL_5_DFFSR_94 ( );
FILL FILL_6_DFFSR_94 ( );
FILL FILL_7_DFFSR_94 ( );
FILL FILL_8_DFFSR_94 ( );
FILL FILL_9_DFFSR_94 ( );
FILL FILL_10_DFFSR_94 ( );
FILL FILL_11_DFFSR_94 ( );
FILL FILL_12_DFFSR_94 ( );
FILL FILL_13_DFFSR_94 ( );
FILL FILL_14_DFFSR_94 ( );
FILL FILL_15_DFFSR_94 ( );
FILL FILL_16_DFFSR_94 ( );
FILL FILL_17_DFFSR_94 ( );
FILL FILL_18_DFFSR_94 ( );
FILL FILL_19_DFFSR_94 ( );
FILL FILL_20_DFFSR_94 ( );
FILL FILL_21_DFFSR_94 ( );
FILL FILL_22_DFFSR_94 ( );
FILL FILL_23_DFFSR_94 ( );
FILL FILL_24_DFFSR_94 ( );
FILL FILL_25_DFFSR_94 ( );
FILL FILL_26_DFFSR_94 ( );
FILL FILL_27_DFFSR_94 ( );
FILL FILL_28_DFFSR_94 ( );
FILL FILL_29_DFFSR_94 ( );
FILL FILL_30_DFFSR_94 ( );
FILL FILL_31_DFFSR_94 ( );
FILL FILL_32_DFFSR_94 ( );
FILL FILL_33_DFFSR_94 ( );
FILL FILL_34_DFFSR_94 ( );
FILL FILL_35_DFFSR_94 ( );
FILL FILL_36_DFFSR_94 ( );
FILL FILL_37_DFFSR_94 ( );
FILL FILL_38_DFFSR_94 ( );
FILL FILL_39_DFFSR_94 ( );
FILL FILL_40_DFFSR_94 ( );
FILL FILL_41_DFFSR_94 ( );
FILL FILL_42_DFFSR_94 ( );
FILL FILL_43_DFFSR_94 ( );
FILL FILL_44_DFFSR_94 ( );
FILL FILL_45_DFFSR_94 ( );
FILL FILL_46_DFFSR_94 ( );
FILL FILL_47_DFFSR_94 ( );
FILL FILL_48_DFFSR_94 ( );
FILL FILL_49_DFFSR_94 ( );
FILL FILL_50_DFFSR_94 ( );
FILL FILL_0_DFFSR_80 ( );
FILL FILL_1_DFFSR_80 ( );
FILL FILL_2_DFFSR_80 ( );
FILL FILL_3_DFFSR_80 ( );
FILL FILL_4_DFFSR_80 ( );
FILL FILL_5_DFFSR_80 ( );
FILL FILL_6_DFFSR_80 ( );
FILL FILL_7_DFFSR_80 ( );
FILL FILL_8_DFFSR_80 ( );
FILL FILL_9_DFFSR_80 ( );
FILL FILL_10_DFFSR_80 ( );
FILL FILL_11_DFFSR_80 ( );
FILL FILL_12_DFFSR_80 ( );
FILL FILL_13_DFFSR_80 ( );
FILL FILL_14_DFFSR_80 ( );
FILL FILL_15_DFFSR_80 ( );
FILL FILL_16_DFFSR_80 ( );
FILL FILL_17_DFFSR_80 ( );
FILL FILL_18_DFFSR_80 ( );
FILL FILL_19_DFFSR_80 ( );
FILL FILL_20_DFFSR_80 ( );
FILL FILL_21_DFFSR_80 ( );
FILL FILL_22_DFFSR_80 ( );
FILL FILL_23_DFFSR_80 ( );
FILL FILL_24_DFFSR_80 ( );
FILL FILL_25_DFFSR_80 ( );
FILL FILL_26_DFFSR_80 ( );
FILL FILL_27_DFFSR_80 ( );
FILL FILL_28_DFFSR_80 ( );
FILL FILL_29_DFFSR_80 ( );
FILL FILL_30_DFFSR_80 ( );
FILL FILL_31_DFFSR_80 ( );
FILL FILL_32_DFFSR_80 ( );
FILL FILL_33_DFFSR_80 ( );
FILL FILL_34_DFFSR_80 ( );
FILL FILL_35_DFFSR_80 ( );
FILL FILL_36_DFFSR_80 ( );
FILL FILL_37_DFFSR_80 ( );
FILL FILL_38_DFFSR_80 ( );
FILL FILL_39_DFFSR_80 ( );
FILL FILL_40_DFFSR_80 ( );
FILL FILL_41_DFFSR_80 ( );
FILL FILL_42_DFFSR_80 ( );
FILL FILL_43_DFFSR_80 ( );
FILL FILL_44_DFFSR_80 ( );
FILL FILL_45_DFFSR_80 ( );
FILL FILL_46_DFFSR_80 ( );
FILL FILL_47_DFFSR_80 ( );
FILL FILL_48_DFFSR_80 ( );
FILL FILL_49_DFFSR_80 ( );
FILL FILL_50_DFFSR_80 ( );
FILL FILL_51_DFFSR_80 ( );
FILL FILL_0_INVX1_424 ( );
FILL FILL_1_INVX1_424 ( );
FILL FILL_2_INVX1_424 ( );
FILL FILL_3_INVX1_424 ( );
FILL FILL_4_INVX1_424 ( );
FILL FILL_0_NAND2X1_273 ( );
FILL FILL_1_NAND2X1_273 ( );
FILL FILL_2_NAND2X1_273 ( );
FILL FILL_3_NAND2X1_273 ( );
FILL FILL_4_NAND2X1_273 ( );
FILL FILL_5_NAND2X1_273 ( );
FILL FILL_6_NAND2X1_273 ( );
FILL FILL_0_NOR2X1_46 ( );
FILL FILL_1_NOR2X1_46 ( );
FILL FILL_2_NOR2X1_46 ( );
FILL FILL_3_NOR2X1_46 ( );
FILL FILL_4_NOR2X1_46 ( );
FILL FILL_5_NOR2X1_46 ( );
FILL FILL_6_NOR2X1_46 ( );
FILL FILL_0_INVX1_157 ( );
FILL FILL_1_INVX1_157 ( );
FILL FILL_2_INVX1_157 ( );
FILL FILL_3_INVX1_157 ( );
FILL FILL_4_INVX1_157 ( );
FILL FILL_0_DFFSR_24 ( );
FILL FILL_1_DFFSR_24 ( );
FILL FILL_2_DFFSR_24 ( );
FILL FILL_3_DFFSR_24 ( );
FILL FILL_4_DFFSR_24 ( );
FILL FILL_5_DFFSR_24 ( );
FILL FILL_6_DFFSR_24 ( );
FILL FILL_7_DFFSR_24 ( );
FILL FILL_8_DFFSR_24 ( );
FILL FILL_9_DFFSR_24 ( );
FILL FILL_10_DFFSR_24 ( );
FILL FILL_11_DFFSR_24 ( );
FILL FILL_12_DFFSR_24 ( );
FILL FILL_13_DFFSR_24 ( );
FILL FILL_14_DFFSR_24 ( );
FILL FILL_15_DFFSR_24 ( );
FILL FILL_16_DFFSR_24 ( );
FILL FILL_17_DFFSR_24 ( );
FILL FILL_18_DFFSR_24 ( );
FILL FILL_19_DFFSR_24 ( );
FILL FILL_20_DFFSR_24 ( );
FILL FILL_21_DFFSR_24 ( );
FILL FILL_22_DFFSR_24 ( );
FILL FILL_23_DFFSR_24 ( );
FILL FILL_24_DFFSR_24 ( );
FILL FILL_25_DFFSR_24 ( );
FILL FILL_26_DFFSR_24 ( );
FILL FILL_27_DFFSR_24 ( );
FILL FILL_28_DFFSR_24 ( );
FILL FILL_29_DFFSR_24 ( );
FILL FILL_30_DFFSR_24 ( );
FILL FILL_31_DFFSR_24 ( );
FILL FILL_32_DFFSR_24 ( );
FILL FILL_33_DFFSR_24 ( );
FILL FILL_34_DFFSR_24 ( );
FILL FILL_35_DFFSR_24 ( );
FILL FILL_36_DFFSR_24 ( );
FILL FILL_37_DFFSR_24 ( );
FILL FILL_38_DFFSR_24 ( );
FILL FILL_39_DFFSR_24 ( );
FILL FILL_40_DFFSR_24 ( );
FILL FILL_41_DFFSR_24 ( );
FILL FILL_42_DFFSR_24 ( );
FILL FILL_43_DFFSR_24 ( );
FILL FILL_44_DFFSR_24 ( );
FILL FILL_45_DFFSR_24 ( );
FILL FILL_46_DFFSR_24 ( );
FILL FILL_47_DFFSR_24 ( );
FILL FILL_48_DFFSR_24 ( );
FILL FILL_49_DFFSR_24 ( );
FILL FILL_50_DFFSR_24 ( );
FILL FILL_0_OAI21X1_42 ( );
FILL FILL_1_OAI21X1_42 ( );
FILL FILL_2_OAI21X1_42 ( );
FILL FILL_3_OAI21X1_42 ( );
FILL FILL_4_OAI21X1_42 ( );
FILL FILL_5_OAI21X1_42 ( );
FILL FILL_6_OAI21X1_42 ( );
FILL FILL_7_OAI21X1_42 ( );
FILL FILL_8_OAI21X1_42 ( );
FILL FILL_0_INVX1_48 ( );
FILL FILL_1_INVX1_48 ( );
FILL FILL_2_INVX1_48 ( );
FILL FILL_3_INVX1_48 ( );
FILL FILL_4_INVX1_48 ( );
FILL FILL_0_INVX1_323 ( );
FILL FILL_1_INVX1_323 ( );
FILL FILL_2_INVX1_323 ( );
FILL FILL_3_INVX1_323 ( );
FILL FILL_4_INVX1_323 ( );
FILL FILL_0_NAND2X1_64 ( );
FILL FILL_1_NAND2X1_64 ( );
FILL FILL_2_NAND2X1_64 ( );
FILL FILL_3_NAND2X1_64 ( );
FILL FILL_4_NAND2X1_64 ( );
FILL FILL_5_NAND2X1_64 ( );
FILL FILL_6_NAND2X1_64 ( );
FILL FILL_0_OAI21X1_64 ( );
FILL FILL_1_OAI21X1_64 ( );
FILL FILL_2_OAI21X1_64 ( );
FILL FILL_3_OAI21X1_64 ( );
FILL FILL_4_OAI21X1_64 ( );
FILL FILL_5_OAI21X1_64 ( );
FILL FILL_6_OAI21X1_64 ( );
FILL FILL_7_OAI21X1_64 ( );
FILL FILL_8_OAI21X1_64 ( );
FILL FILL_9_OAI21X1_64 ( );
FILL FILL_0_NAND2X1_234 ( );
FILL FILL_1_NAND2X1_234 ( );
FILL FILL_2_NAND2X1_234 ( );
FILL FILL_3_NAND2X1_234 ( );
FILL FILL_4_NAND2X1_234 ( );
FILL FILL_5_NAND2X1_234 ( );
FILL FILL_6_NAND2X1_234 ( );
FILL FILL_0_NOR2X1_12 ( );
FILL FILL_1_NOR2X1_12 ( );
FILL FILL_2_NOR2X1_12 ( );
FILL FILL_3_NOR2X1_12 ( );
FILL FILL_4_NOR2X1_12 ( );
FILL FILL_5_NOR2X1_12 ( );
FILL FILL_6_NOR2X1_12 ( );
FILL FILL_0_OAI22X1_5 ( );
FILL FILL_1_OAI22X1_5 ( );
FILL FILL_2_OAI22X1_5 ( );
FILL FILL_3_OAI22X1_5 ( );
FILL FILL_4_OAI22X1_5 ( );
FILL FILL_5_OAI22X1_5 ( );
FILL FILL_6_OAI22X1_5 ( );
FILL FILL_7_OAI22X1_5 ( );
FILL FILL_8_OAI22X1_5 ( );
FILL FILL_9_OAI22X1_5 ( );
FILL FILL_10_OAI22X1_5 ( );
FILL FILL_11_OAI22X1_5 ( );
FILL FILL_0_INVX1_285 ( );
FILL FILL_1_INVX1_285 ( );
FILL FILL_2_INVX1_285 ( );
FILL FILL_3_INVX1_285 ( );
FILL FILL_0_INVX1_263 ( );
FILL FILL_1_INVX1_263 ( );
FILL FILL_2_INVX1_263 ( );
FILL FILL_3_INVX1_263 ( );
FILL FILL_0_INVX1_58 ( );
FILL FILL_1_INVX1_58 ( );
FILL FILL_2_INVX1_58 ( );
FILL FILL_3_INVX1_58 ( );
FILL FILL_0_DFFPOSX1_19 ( );
FILL FILL_1_DFFPOSX1_19 ( );
FILL FILL_2_DFFPOSX1_19 ( );
FILL FILL_3_DFFPOSX1_19 ( );
FILL FILL_4_DFFPOSX1_19 ( );
FILL FILL_5_DFFPOSX1_19 ( );
FILL FILL_6_DFFPOSX1_19 ( );
FILL FILL_7_DFFPOSX1_19 ( );
FILL FILL_8_DFFPOSX1_19 ( );
FILL FILL_9_DFFPOSX1_19 ( );
FILL FILL_10_DFFPOSX1_19 ( );
FILL FILL_11_DFFPOSX1_19 ( );
FILL FILL_12_DFFPOSX1_19 ( );
FILL FILL_13_DFFPOSX1_19 ( );
FILL FILL_14_DFFPOSX1_19 ( );
FILL FILL_15_DFFPOSX1_19 ( );
FILL FILL_16_DFFPOSX1_19 ( );
FILL FILL_17_DFFPOSX1_19 ( );
FILL FILL_18_DFFPOSX1_19 ( );
FILL FILL_19_DFFPOSX1_19 ( );
FILL FILL_20_DFFPOSX1_19 ( );
FILL FILL_21_DFFPOSX1_19 ( );
FILL FILL_22_DFFPOSX1_19 ( );
FILL FILL_23_DFFPOSX1_19 ( );
FILL FILL_24_DFFPOSX1_19 ( );
FILL FILL_25_DFFPOSX1_19 ( );
FILL FILL_26_DFFPOSX1_19 ( );
FILL FILL_27_DFFPOSX1_19 ( );
FILL FILL_0_NAND2X1_11 ( );
FILL FILL_1_NAND2X1_11 ( );
FILL FILL_2_NAND2X1_11 ( );
FILL FILL_3_NAND2X1_11 ( );
FILL FILL_4_NAND2X1_11 ( );
FILL FILL_5_NAND2X1_11 ( );
FILL FILL_6_NAND2X1_11 ( );
FILL FILL_0_DFFSR_13 ( );
FILL FILL_1_DFFSR_13 ( );
FILL FILL_2_DFFSR_13 ( );
FILL FILL_3_DFFSR_13 ( );
FILL FILL_4_DFFSR_13 ( );
FILL FILL_5_DFFSR_13 ( );
FILL FILL_6_DFFSR_13 ( );
FILL FILL_7_DFFSR_13 ( );
FILL FILL_8_DFFSR_13 ( );
FILL FILL_9_DFFSR_13 ( );
FILL FILL_10_DFFSR_13 ( );
FILL FILL_11_DFFSR_13 ( );
FILL FILL_12_DFFSR_13 ( );
FILL FILL_13_DFFSR_13 ( );
FILL FILL_14_DFFSR_13 ( );
FILL FILL_15_DFFSR_13 ( );
FILL FILL_16_DFFSR_13 ( );
FILL FILL_17_DFFSR_13 ( );
FILL FILL_18_DFFSR_13 ( );
FILL FILL_19_DFFSR_13 ( );
FILL FILL_20_DFFSR_13 ( );
FILL FILL_21_DFFSR_13 ( );
FILL FILL_22_DFFSR_13 ( );
FILL FILL_23_DFFSR_13 ( );
FILL FILL_24_DFFSR_13 ( );
FILL FILL_25_DFFSR_13 ( );
FILL FILL_26_DFFSR_13 ( );
FILL FILL_27_DFFSR_13 ( );
FILL FILL_28_DFFSR_13 ( );
FILL FILL_29_DFFSR_13 ( );
FILL FILL_30_DFFSR_13 ( );
FILL FILL_31_DFFSR_13 ( );
FILL FILL_32_DFFSR_13 ( );
FILL FILL_33_DFFSR_13 ( );
FILL FILL_34_DFFSR_13 ( );
FILL FILL_35_DFFSR_13 ( );
FILL FILL_36_DFFSR_13 ( );
FILL FILL_37_DFFSR_13 ( );
FILL FILL_38_DFFSR_13 ( );
FILL FILL_39_DFFSR_13 ( );
FILL FILL_40_DFFSR_13 ( );
FILL FILL_41_DFFSR_13 ( );
FILL FILL_42_DFFSR_13 ( );
FILL FILL_43_DFFSR_13 ( );
FILL FILL_44_DFFSR_13 ( );
FILL FILL_45_DFFSR_13 ( );
FILL FILL_46_DFFSR_13 ( );
FILL FILL_47_DFFSR_13 ( );
FILL FILL_48_DFFSR_13 ( );
FILL FILL_49_DFFSR_13 ( );
FILL FILL_50_DFFSR_13 ( );
FILL FILL_0_OAI21X1_13 ( );
FILL FILL_1_OAI21X1_13 ( );
FILL FILL_2_OAI21X1_13 ( );
FILL FILL_3_OAI21X1_13 ( );
FILL FILL_4_OAI21X1_13 ( );
FILL FILL_5_OAI21X1_13 ( );
FILL FILL_6_OAI21X1_13 ( );
FILL FILL_7_OAI21X1_13 ( );
FILL FILL_8_OAI21X1_13 ( );
FILL FILL_9_OAI21X1_13 ( );
FILL FILL_0_DFFSR_176 ( );
FILL FILL_1_DFFSR_176 ( );
FILL FILL_2_DFFSR_176 ( );
FILL FILL_3_DFFSR_176 ( );
FILL FILL_4_DFFSR_176 ( );
FILL FILL_5_DFFSR_176 ( );
FILL FILL_6_DFFSR_176 ( );
FILL FILL_7_DFFSR_176 ( );
FILL FILL_8_DFFSR_176 ( );
FILL FILL_9_DFFSR_176 ( );
FILL FILL_10_DFFSR_176 ( );
FILL FILL_11_DFFSR_176 ( );
FILL FILL_12_DFFSR_176 ( );
FILL FILL_13_DFFSR_176 ( );
FILL FILL_14_DFFSR_176 ( );
FILL FILL_15_DFFSR_176 ( );
FILL FILL_16_DFFSR_176 ( );
FILL FILL_17_DFFSR_176 ( );
FILL FILL_18_DFFSR_176 ( );
FILL FILL_19_DFFSR_176 ( );
FILL FILL_20_DFFSR_176 ( );
FILL FILL_21_DFFSR_176 ( );
FILL FILL_22_DFFSR_176 ( );
FILL FILL_23_DFFSR_176 ( );
FILL FILL_24_DFFSR_176 ( );
FILL FILL_25_DFFSR_176 ( );
FILL FILL_26_DFFSR_176 ( );
FILL FILL_27_DFFSR_176 ( );
FILL FILL_28_DFFSR_176 ( );
FILL FILL_29_DFFSR_176 ( );
FILL FILL_30_DFFSR_176 ( );
FILL FILL_31_DFFSR_176 ( );
FILL FILL_32_DFFSR_176 ( );
FILL FILL_33_DFFSR_176 ( );
FILL FILL_34_DFFSR_176 ( );
FILL FILL_35_DFFSR_176 ( );
FILL FILL_36_DFFSR_176 ( );
FILL FILL_37_DFFSR_176 ( );
FILL FILL_38_DFFSR_176 ( );
FILL FILL_39_DFFSR_176 ( );
FILL FILL_40_DFFSR_176 ( );
FILL FILL_41_DFFSR_176 ( );
FILL FILL_42_DFFSR_176 ( );
FILL FILL_43_DFFSR_176 ( );
FILL FILL_44_DFFSR_176 ( );
FILL FILL_45_DFFSR_176 ( );
FILL FILL_46_DFFSR_176 ( );
FILL FILL_47_DFFSR_176 ( );
FILL FILL_48_DFFSR_176 ( );
FILL FILL_49_DFFSR_176 ( );
FILL FILL_50_DFFSR_176 ( );
FILL FILL_51_DFFSR_176 ( );
FILL FILL_0_BUFX2_29 ( );
FILL FILL_1_BUFX2_29 ( );
FILL FILL_2_BUFX2_29 ( );
FILL FILL_3_BUFX2_29 ( );
FILL FILL_4_BUFX2_29 ( );
FILL FILL_5_BUFX2_29 ( );
FILL FILL_6_BUFX2_29 ( );
FILL FILL_0_DFFSR_112 ( );
FILL FILL_1_DFFSR_112 ( );
FILL FILL_2_DFFSR_112 ( );
FILL FILL_3_DFFSR_112 ( );
FILL FILL_4_DFFSR_112 ( );
FILL FILL_5_DFFSR_112 ( );
FILL FILL_6_DFFSR_112 ( );
FILL FILL_7_DFFSR_112 ( );
FILL FILL_8_DFFSR_112 ( );
FILL FILL_9_DFFSR_112 ( );
FILL FILL_10_DFFSR_112 ( );
FILL FILL_11_DFFSR_112 ( );
FILL FILL_12_DFFSR_112 ( );
FILL FILL_13_DFFSR_112 ( );
FILL FILL_14_DFFSR_112 ( );
FILL FILL_15_DFFSR_112 ( );
FILL FILL_16_DFFSR_112 ( );
FILL FILL_17_DFFSR_112 ( );
FILL FILL_18_DFFSR_112 ( );
FILL FILL_19_DFFSR_112 ( );
FILL FILL_20_DFFSR_112 ( );
FILL FILL_21_DFFSR_112 ( );
FILL FILL_22_DFFSR_112 ( );
FILL FILL_23_DFFSR_112 ( );
FILL FILL_24_DFFSR_112 ( );
FILL FILL_25_DFFSR_112 ( );
FILL FILL_26_DFFSR_112 ( );
FILL FILL_27_DFFSR_112 ( );
FILL FILL_28_DFFSR_112 ( );
FILL FILL_29_DFFSR_112 ( );
FILL FILL_30_DFFSR_112 ( );
FILL FILL_31_DFFSR_112 ( );
FILL FILL_32_DFFSR_112 ( );
FILL FILL_33_DFFSR_112 ( );
FILL FILL_34_DFFSR_112 ( );
FILL FILL_35_DFFSR_112 ( );
FILL FILL_36_DFFSR_112 ( );
FILL FILL_37_DFFSR_112 ( );
FILL FILL_38_DFFSR_112 ( );
FILL FILL_39_DFFSR_112 ( );
FILL FILL_40_DFFSR_112 ( );
FILL FILL_41_DFFSR_112 ( );
FILL FILL_42_DFFSR_112 ( );
FILL FILL_43_DFFSR_112 ( );
FILL FILL_44_DFFSR_112 ( );
FILL FILL_45_DFFSR_112 ( );
FILL FILL_46_DFFSR_112 ( );
FILL FILL_47_DFFSR_112 ( );
FILL FILL_48_DFFSR_112 ( );
FILL FILL_49_DFFSR_112 ( );
FILL FILL_50_DFFSR_112 ( );
FILL FILL_0_INVX1_373 ( );
FILL FILL_1_INVX1_373 ( );
FILL FILL_2_INVX1_373 ( );
FILL FILL_3_INVX1_373 ( );
FILL FILL_0_INVX1_392 ( );
FILL FILL_1_INVX1_392 ( );
FILL FILL_2_INVX1_392 ( );
FILL FILL_3_INVX1_392 ( );
FILL FILL_4_INVX1_392 ( );
FILL FILL_0_OAI22X1_67 ( );
FILL FILL_1_OAI22X1_67 ( );
FILL FILL_2_OAI22X1_67 ( );
FILL FILL_3_OAI22X1_67 ( );
FILL FILL_4_OAI22X1_67 ( );
FILL FILL_5_OAI22X1_67 ( );
FILL FILL_6_OAI22X1_67 ( );
FILL FILL_7_OAI22X1_67 ( );
FILL FILL_8_OAI22X1_67 ( );
FILL FILL_9_OAI22X1_67 ( );
FILL FILL_10_OAI22X1_67 ( );
FILL FILL_11_OAI22X1_67 ( );
FILL FILL_0_INVX1_340 ( );
FILL FILL_1_INVX1_340 ( );
FILL FILL_2_INVX1_340 ( );
FILL FILL_3_INVX1_340 ( );
FILL FILL_4_INVX1_340 ( );
FILL FILL_0_INVX1_341 ( );
FILL FILL_1_INVX1_341 ( );
FILL FILL_2_INVX1_341 ( );
FILL FILL_3_INVX1_341 ( );
FILL FILL_0_NAND2X1_93 ( );
FILL FILL_1_NAND2X1_93 ( );
FILL FILL_2_NAND2X1_93 ( );
FILL FILL_3_NAND2X1_93 ( );
FILL FILL_4_NAND2X1_93 ( );
FILL FILL_5_NAND2X1_93 ( );
FILL FILL_6_NAND2X1_93 ( );
FILL FILL_0_INVX1_388 ( );
FILL FILL_1_INVX1_388 ( );
FILL FILL_2_INVX1_388 ( );
FILL FILL_3_INVX1_388 ( );
FILL FILL_4_INVX1_388 ( );
FILL FILL_0_NAND2X1_88 ( );
FILL FILL_1_NAND2X1_88 ( );
FILL FILL_2_NAND2X1_88 ( );
FILL FILL_3_NAND2X1_88 ( );
FILL FILL_4_NAND2X1_88 ( );
FILL FILL_5_NAND2X1_88 ( );
FILL FILL_6_NAND2X1_88 ( );
FILL FILL_0_INVX1_85 ( );
FILL FILL_1_INVX1_85 ( );
FILL FILL_2_INVX1_85 ( );
FILL FILL_3_INVX1_85 ( );
FILL FILL_4_INVX1_85 ( );
FILL FILL_0_BUFX2_18 ( );
FILL FILL_1_BUFX2_18 ( );
FILL FILL_2_BUFX2_18 ( );
FILL FILL_3_BUFX2_18 ( );
FILL FILL_4_BUFX2_18 ( );
FILL FILL_5_BUFX2_18 ( );
FILL FILL_6_BUFX2_18 ( );
FILL FILL_0_DFFSR_65 ( );
FILL FILL_1_DFFSR_65 ( );
FILL FILL_2_DFFSR_65 ( );
FILL FILL_3_DFFSR_65 ( );
FILL FILL_4_DFFSR_65 ( );
FILL FILL_5_DFFSR_65 ( );
FILL FILL_6_DFFSR_65 ( );
FILL FILL_7_DFFSR_65 ( );
FILL FILL_8_DFFSR_65 ( );
FILL FILL_9_DFFSR_65 ( );
FILL FILL_10_DFFSR_65 ( );
FILL FILL_11_DFFSR_65 ( );
FILL FILL_12_DFFSR_65 ( );
FILL FILL_13_DFFSR_65 ( );
FILL FILL_14_DFFSR_65 ( );
FILL FILL_15_DFFSR_65 ( );
FILL FILL_16_DFFSR_65 ( );
FILL FILL_17_DFFSR_65 ( );
FILL FILL_18_DFFSR_65 ( );
FILL FILL_19_DFFSR_65 ( );
FILL FILL_20_DFFSR_65 ( );
FILL FILL_21_DFFSR_65 ( );
FILL FILL_22_DFFSR_65 ( );
FILL FILL_23_DFFSR_65 ( );
FILL FILL_24_DFFSR_65 ( );
FILL FILL_25_DFFSR_65 ( );
FILL FILL_26_DFFSR_65 ( );
FILL FILL_27_DFFSR_65 ( );
FILL FILL_28_DFFSR_65 ( );
FILL FILL_29_DFFSR_65 ( );
FILL FILL_30_DFFSR_65 ( );
FILL FILL_31_DFFSR_65 ( );
FILL FILL_32_DFFSR_65 ( );
FILL FILL_33_DFFSR_65 ( );
FILL FILL_34_DFFSR_65 ( );
FILL FILL_35_DFFSR_65 ( );
FILL FILL_36_DFFSR_65 ( );
FILL FILL_37_DFFSR_65 ( );
FILL FILL_38_DFFSR_65 ( );
FILL FILL_39_DFFSR_65 ( );
FILL FILL_40_DFFSR_65 ( );
FILL FILL_41_DFFSR_65 ( );
FILL FILL_42_DFFSR_65 ( );
FILL FILL_43_DFFSR_65 ( );
FILL FILL_44_DFFSR_65 ( );
FILL FILL_45_DFFSR_65 ( );
FILL FILL_46_DFFSR_65 ( );
FILL FILL_47_DFFSR_65 ( );
FILL FILL_48_DFFSR_65 ( );
FILL FILL_49_DFFSR_65 ( );
FILL FILL_50_DFFSR_65 ( );
FILL FILL_0_OAI21X1_139 ( );
FILL FILL_1_OAI21X1_139 ( );
FILL FILL_2_OAI21X1_139 ( );
FILL FILL_3_OAI21X1_139 ( );
FILL FILL_4_OAI21X1_139 ( );
FILL FILL_5_OAI21X1_139 ( );
FILL FILL_6_OAI21X1_139 ( );
FILL FILL_7_OAI21X1_139 ( );
FILL FILL_8_OAI21X1_139 ( );
FILL FILL_0_AND2X2_15 ( );
FILL FILL_1_AND2X2_15 ( );
FILL FILL_2_AND2X2_15 ( );
FILL FILL_3_AND2X2_15 ( );
FILL FILL_4_AND2X2_15 ( );
FILL FILL_5_AND2X2_15 ( );
FILL FILL_6_AND2X2_15 ( );
FILL FILL_7_AND2X2_15 ( );
FILL FILL_8_AND2X2_15 ( );
FILL FILL_9_AND2X2_15 ( );
FILL FILL_0_INVX1_19 ( );
FILL FILL_1_INVX1_19 ( );
FILL FILL_2_INVX1_19 ( );
FILL FILL_3_INVX1_19 ( );
FILL FILL_0_NAND2X1_32 ( );
FILL FILL_1_NAND2X1_32 ( );
FILL FILL_2_NAND2X1_32 ( );
FILL FILL_3_NAND2X1_32 ( );
FILL FILL_4_NAND2X1_32 ( );
FILL FILL_5_NAND2X1_32 ( );
FILL FILL_6_NAND2X1_32 ( );
FILL FILL_0_INVX1_36 ( );
FILL FILL_1_INVX1_36 ( );
FILL FILL_2_INVX1_36 ( );
FILL FILL_3_INVX1_36 ( );
FILL FILL_4_INVX1_36 ( );
FILL FILL_0_DFFSR_42 ( );
FILL FILL_1_DFFSR_42 ( );
FILL FILL_2_DFFSR_42 ( );
FILL FILL_3_DFFSR_42 ( );
FILL FILL_4_DFFSR_42 ( );
FILL FILL_5_DFFSR_42 ( );
FILL FILL_6_DFFSR_42 ( );
FILL FILL_7_DFFSR_42 ( );
FILL FILL_8_DFFSR_42 ( );
FILL FILL_9_DFFSR_42 ( );
FILL FILL_10_DFFSR_42 ( );
FILL FILL_11_DFFSR_42 ( );
FILL FILL_12_DFFSR_42 ( );
FILL FILL_13_DFFSR_42 ( );
FILL FILL_14_DFFSR_42 ( );
FILL FILL_15_DFFSR_42 ( );
FILL FILL_16_DFFSR_42 ( );
FILL FILL_17_DFFSR_42 ( );
FILL FILL_18_DFFSR_42 ( );
FILL FILL_19_DFFSR_42 ( );
FILL FILL_20_DFFSR_42 ( );
FILL FILL_21_DFFSR_42 ( );
FILL FILL_22_DFFSR_42 ( );
FILL FILL_23_DFFSR_42 ( );
FILL FILL_24_DFFSR_42 ( );
FILL FILL_25_DFFSR_42 ( );
FILL FILL_26_DFFSR_42 ( );
FILL FILL_27_DFFSR_42 ( );
FILL FILL_28_DFFSR_42 ( );
FILL FILL_29_DFFSR_42 ( );
FILL FILL_30_DFFSR_42 ( );
FILL FILL_31_DFFSR_42 ( );
FILL FILL_32_DFFSR_42 ( );
FILL FILL_33_DFFSR_42 ( );
FILL FILL_34_DFFSR_42 ( );
FILL FILL_35_DFFSR_42 ( );
FILL FILL_36_DFFSR_42 ( );
FILL FILL_37_DFFSR_42 ( );
FILL FILL_38_DFFSR_42 ( );
FILL FILL_39_DFFSR_42 ( );
FILL FILL_40_DFFSR_42 ( );
FILL FILL_41_DFFSR_42 ( );
FILL FILL_42_DFFSR_42 ( );
FILL FILL_43_DFFSR_42 ( );
FILL FILL_44_DFFSR_42 ( );
FILL FILL_45_DFFSR_42 ( );
FILL FILL_46_DFFSR_42 ( );
FILL FILL_47_DFFSR_42 ( );
FILL FILL_48_DFFSR_42 ( );
FILL FILL_49_DFFSR_42 ( );
FILL FILL_50_DFFSR_42 ( );
FILL FILL_51_DFFSR_42 ( );
FILL FILL_0_NAND2X1_58 ( );
FILL FILL_1_NAND2X1_58 ( );
FILL FILL_2_NAND2X1_58 ( );
FILL FILL_3_NAND2X1_58 ( );
FILL FILL_4_NAND2X1_58 ( );
FILL FILL_5_NAND2X1_58 ( );
FILL FILL_6_NAND2X1_58 ( );
FILL FILL_0_NOR2X1_16 ( );
FILL FILL_1_NOR2X1_16 ( );
FILL FILL_2_NOR2X1_16 ( );
FILL FILL_3_NOR2X1_16 ( );
FILL FILL_4_NOR2X1_16 ( );
FILL FILL_5_NOR2X1_16 ( );
FILL FILL_6_NOR2X1_16 ( );
FILL FILL_0_INVX1_66 ( );
FILL FILL_1_INVX1_66 ( );
FILL FILL_2_INVX1_66 ( );
FILL FILL_3_INVX1_66 ( );
FILL FILL_0_OAI21X1_58 ( );
FILL FILL_1_OAI21X1_58 ( );
FILL FILL_2_OAI21X1_58 ( );
FILL FILL_3_OAI21X1_58 ( );
FILL FILL_4_OAI21X1_58 ( );
FILL FILL_5_OAI21X1_58 ( );
FILL FILL_6_OAI21X1_58 ( );
FILL FILL_7_OAI21X1_58 ( );
FILL FILL_8_OAI21X1_58 ( );
FILL FILL_9_OAI21X1_58 ( );
FILL FILL_0_OAI22X1_13 ( );
FILL FILL_1_OAI22X1_13 ( );
FILL FILL_2_OAI22X1_13 ( );
FILL FILL_3_OAI22X1_13 ( );
FILL FILL_4_OAI22X1_13 ( );
FILL FILL_5_OAI22X1_13 ( );
FILL FILL_6_OAI22X1_13 ( );
FILL FILL_7_OAI22X1_13 ( );
FILL FILL_8_OAI22X1_13 ( );
FILL FILL_9_OAI22X1_13 ( );
FILL FILL_10_OAI22X1_13 ( );
FILL FILL_11_OAI22X1_13 ( );
FILL FILL_0_INVX1_282 ( );
FILL FILL_1_INVX1_282 ( );
FILL FILL_2_INVX1_282 ( );
FILL FILL_3_INVX1_282 ( );
FILL FILL_4_INVX1_282 ( );
FILL FILL_0_INVX1_298 ( );
FILL FILL_1_INVX1_298 ( );
FILL FILL_2_INVX1_298 ( );
FILL FILL_3_INVX1_298 ( );
FILL FILL_4_INVX1_298 ( );
FILL FILL_0_INVX1_281 ( );
FILL FILL_1_INVX1_281 ( );
FILL FILL_2_INVX1_281 ( );
FILL FILL_3_INVX1_281 ( );
FILL FILL_0_INVX1_33 ( );
FILL FILL_1_INVX1_33 ( );
FILL FILL_2_INVX1_33 ( );
FILL FILL_3_INVX1_33 ( );
FILL FILL_4_INVX1_33 ( );
FILL FILL_0_OAI21X1_29 ( );
FILL FILL_1_OAI21X1_29 ( );
FILL FILL_2_OAI21X1_29 ( );
FILL FILL_3_OAI21X1_29 ( );
FILL FILL_4_OAI21X1_29 ( );
FILL FILL_5_OAI21X1_29 ( );
FILL FILL_6_OAI21X1_29 ( );
FILL FILL_7_OAI21X1_29 ( );
FILL FILL_8_OAI21X1_29 ( );
FILL FILL_0_DFFPOSX1_28 ( );
FILL FILL_1_DFFPOSX1_28 ( );
FILL FILL_2_DFFPOSX1_28 ( );
FILL FILL_3_DFFPOSX1_28 ( );
FILL FILL_4_DFFPOSX1_28 ( );
FILL FILL_5_DFFPOSX1_28 ( );
FILL FILL_6_DFFPOSX1_28 ( );
FILL FILL_7_DFFPOSX1_28 ( );
FILL FILL_8_DFFPOSX1_28 ( );
FILL FILL_9_DFFPOSX1_28 ( );
FILL FILL_10_DFFPOSX1_28 ( );
FILL FILL_11_DFFPOSX1_28 ( );
FILL FILL_12_DFFPOSX1_28 ( );
FILL FILL_13_DFFPOSX1_28 ( );
FILL FILL_14_DFFPOSX1_28 ( );
FILL FILL_15_DFFPOSX1_28 ( );
FILL FILL_16_DFFPOSX1_28 ( );
FILL FILL_17_DFFPOSX1_28 ( );
FILL FILL_18_DFFPOSX1_28 ( );
FILL FILL_19_DFFPOSX1_28 ( );
FILL FILL_20_DFFPOSX1_28 ( );
FILL FILL_21_DFFPOSX1_28 ( );
FILL FILL_22_DFFPOSX1_28 ( );
FILL FILL_23_DFFPOSX1_28 ( );
FILL FILL_24_DFFPOSX1_28 ( );
FILL FILL_25_DFFPOSX1_28 ( );
FILL FILL_26_DFFPOSX1_28 ( );
FILL FILL_27_DFFPOSX1_28 ( );
FILL FILL_0_INVX1_15 ( );
FILL FILL_1_INVX1_15 ( );
FILL FILL_2_INVX1_15 ( );
FILL FILL_3_INVX1_15 ( );
FILL FILL_0_DFFSR_163 ( );
FILL FILL_1_DFFSR_163 ( );
FILL FILL_2_DFFSR_163 ( );
FILL FILL_3_DFFSR_163 ( );
FILL FILL_4_DFFSR_163 ( );
FILL FILL_5_DFFSR_163 ( );
FILL FILL_6_DFFSR_163 ( );
FILL FILL_7_DFFSR_163 ( );
FILL FILL_8_DFFSR_163 ( );
FILL FILL_9_DFFSR_163 ( );
FILL FILL_10_DFFSR_163 ( );
FILL FILL_11_DFFSR_163 ( );
FILL FILL_12_DFFSR_163 ( );
FILL FILL_13_DFFSR_163 ( );
FILL FILL_14_DFFSR_163 ( );
FILL FILL_15_DFFSR_163 ( );
FILL FILL_16_DFFSR_163 ( );
FILL FILL_17_DFFSR_163 ( );
FILL FILL_18_DFFSR_163 ( );
FILL FILL_19_DFFSR_163 ( );
FILL FILL_20_DFFSR_163 ( );
FILL FILL_21_DFFSR_163 ( );
FILL FILL_22_DFFSR_163 ( );
FILL FILL_23_DFFSR_163 ( );
FILL FILL_24_DFFSR_163 ( );
FILL FILL_25_DFFSR_163 ( );
FILL FILL_26_DFFSR_163 ( );
FILL FILL_27_DFFSR_163 ( );
FILL FILL_28_DFFSR_163 ( );
FILL FILL_29_DFFSR_163 ( );
FILL FILL_30_DFFSR_163 ( );
FILL FILL_31_DFFSR_163 ( );
FILL FILL_32_DFFSR_163 ( );
FILL FILL_33_DFFSR_163 ( );
FILL FILL_34_DFFSR_163 ( );
FILL FILL_35_DFFSR_163 ( );
FILL FILL_36_DFFSR_163 ( );
FILL FILL_37_DFFSR_163 ( );
FILL FILL_38_DFFSR_163 ( );
FILL FILL_39_DFFSR_163 ( );
FILL FILL_40_DFFSR_163 ( );
FILL FILL_41_DFFSR_163 ( );
FILL FILL_42_DFFSR_163 ( );
FILL FILL_43_DFFSR_163 ( );
FILL FILL_44_DFFSR_163 ( );
FILL FILL_45_DFFSR_163 ( );
FILL FILL_46_DFFSR_163 ( );
FILL FILL_47_DFFSR_163 ( );
FILL FILL_48_DFFSR_163 ( );
FILL FILL_49_DFFSR_163 ( );
FILL FILL_50_DFFSR_163 ( );
FILL FILL_0_INVX1_406 ( );
FILL FILL_1_INVX1_406 ( );
FILL FILL_2_INVX1_406 ( );
FILL FILL_3_INVX1_406 ( );
FILL FILL_0_NAND2X1_166 ( );
FILL FILL_1_NAND2X1_166 ( );
FILL FILL_2_NAND2X1_166 ( );
FILL FILL_3_NAND2X1_166 ( );
FILL FILL_4_NAND2X1_166 ( );
FILL FILL_5_NAND2X1_166 ( );
FILL FILL_6_NAND2X1_166 ( );
FILL FILL_0_DFFPOSX1_6 ( );
FILL FILL_1_DFFPOSX1_6 ( );
FILL FILL_2_DFFPOSX1_6 ( );
FILL FILL_3_DFFPOSX1_6 ( );
FILL FILL_4_DFFPOSX1_6 ( );
FILL FILL_5_DFFPOSX1_6 ( );
FILL FILL_6_DFFPOSX1_6 ( );
FILL FILL_7_DFFPOSX1_6 ( );
FILL FILL_8_DFFPOSX1_6 ( );
FILL FILL_9_DFFPOSX1_6 ( );
FILL FILL_10_DFFPOSX1_6 ( );
FILL FILL_11_DFFPOSX1_6 ( );
FILL FILL_12_DFFPOSX1_6 ( );
FILL FILL_13_DFFPOSX1_6 ( );
FILL FILL_14_DFFPOSX1_6 ( );
FILL FILL_15_DFFPOSX1_6 ( );
FILL FILL_16_DFFPOSX1_6 ( );
FILL FILL_17_DFFPOSX1_6 ( );
FILL FILL_18_DFFPOSX1_6 ( );
FILL FILL_19_DFFPOSX1_6 ( );
FILL FILL_20_DFFPOSX1_6 ( );
FILL FILL_21_DFFPOSX1_6 ( );
FILL FILL_22_DFFPOSX1_6 ( );
FILL FILL_23_DFFPOSX1_6 ( );
FILL FILL_24_DFFPOSX1_6 ( );
FILL FILL_25_DFFPOSX1_6 ( );
FILL FILL_26_DFFPOSX1_6 ( );
FILL FILL_27_DFFPOSX1_6 ( );
FILL FILL_0_DFFSR_87 ( );
FILL FILL_1_DFFSR_87 ( );
FILL FILL_2_DFFSR_87 ( );
FILL FILL_3_DFFSR_87 ( );
FILL FILL_4_DFFSR_87 ( );
FILL FILL_5_DFFSR_87 ( );
FILL FILL_6_DFFSR_87 ( );
FILL FILL_7_DFFSR_87 ( );
FILL FILL_8_DFFSR_87 ( );
FILL FILL_9_DFFSR_87 ( );
FILL FILL_10_DFFSR_87 ( );
FILL FILL_11_DFFSR_87 ( );
FILL FILL_12_DFFSR_87 ( );
FILL FILL_13_DFFSR_87 ( );
FILL FILL_14_DFFSR_87 ( );
FILL FILL_15_DFFSR_87 ( );
FILL FILL_16_DFFSR_87 ( );
FILL FILL_17_DFFSR_87 ( );
FILL FILL_18_DFFSR_87 ( );
FILL FILL_19_DFFSR_87 ( );
FILL FILL_20_DFFSR_87 ( );
FILL FILL_21_DFFSR_87 ( );
FILL FILL_22_DFFSR_87 ( );
FILL FILL_23_DFFSR_87 ( );
FILL FILL_24_DFFSR_87 ( );
FILL FILL_25_DFFSR_87 ( );
FILL FILL_26_DFFSR_87 ( );
FILL FILL_27_DFFSR_87 ( );
FILL FILL_28_DFFSR_87 ( );
FILL FILL_29_DFFSR_87 ( );
FILL FILL_30_DFFSR_87 ( );
FILL FILL_31_DFFSR_87 ( );
FILL FILL_32_DFFSR_87 ( );
FILL FILL_33_DFFSR_87 ( );
FILL FILL_34_DFFSR_87 ( );
FILL FILL_35_DFFSR_87 ( );
FILL FILL_36_DFFSR_87 ( );
FILL FILL_37_DFFSR_87 ( );
FILL FILL_38_DFFSR_87 ( );
FILL FILL_39_DFFSR_87 ( );
FILL FILL_40_DFFSR_87 ( );
FILL FILL_41_DFFSR_87 ( );
FILL FILL_42_DFFSR_87 ( );
FILL FILL_43_DFFSR_87 ( );
FILL FILL_44_DFFSR_87 ( );
FILL FILL_45_DFFSR_87 ( );
FILL FILL_46_DFFSR_87 ( );
FILL FILL_47_DFFSR_87 ( );
FILL FILL_48_DFFSR_87 ( );
FILL FILL_49_DFFSR_87 ( );
FILL FILL_50_DFFSR_87 ( );
FILL FILL_51_DFFSR_87 ( );
FILL FILL_0_INVX1_393 ( );
FILL FILL_1_INVX1_393 ( );
FILL FILL_2_INVX1_393 ( );
FILL FILL_3_INVX1_393 ( );
FILL FILL_0_DFFSR_88 ( );
FILL FILL_1_DFFSR_88 ( );
FILL FILL_2_DFFSR_88 ( );
FILL FILL_3_DFFSR_88 ( );
FILL FILL_4_DFFSR_88 ( );
FILL FILL_5_DFFSR_88 ( );
FILL FILL_6_DFFSR_88 ( );
FILL FILL_7_DFFSR_88 ( );
FILL FILL_8_DFFSR_88 ( );
FILL FILL_9_DFFSR_88 ( );
FILL FILL_10_DFFSR_88 ( );
FILL FILL_11_DFFSR_88 ( );
FILL FILL_12_DFFSR_88 ( );
FILL FILL_13_DFFSR_88 ( );
FILL FILL_14_DFFSR_88 ( );
FILL FILL_15_DFFSR_88 ( );
FILL FILL_16_DFFSR_88 ( );
FILL FILL_17_DFFSR_88 ( );
FILL FILL_18_DFFSR_88 ( );
FILL FILL_19_DFFSR_88 ( );
FILL FILL_20_DFFSR_88 ( );
FILL FILL_21_DFFSR_88 ( );
FILL FILL_22_DFFSR_88 ( );
FILL FILL_23_DFFSR_88 ( );
FILL FILL_24_DFFSR_88 ( );
FILL FILL_25_DFFSR_88 ( );
FILL FILL_26_DFFSR_88 ( );
FILL FILL_27_DFFSR_88 ( );
FILL FILL_28_DFFSR_88 ( );
FILL FILL_29_DFFSR_88 ( );
FILL FILL_30_DFFSR_88 ( );
FILL FILL_31_DFFSR_88 ( );
FILL FILL_32_DFFSR_88 ( );
FILL FILL_33_DFFSR_88 ( );
FILL FILL_34_DFFSR_88 ( );
FILL FILL_35_DFFSR_88 ( );
FILL FILL_36_DFFSR_88 ( );
FILL FILL_37_DFFSR_88 ( );
FILL FILL_38_DFFSR_88 ( );
FILL FILL_39_DFFSR_88 ( );
FILL FILL_40_DFFSR_88 ( );
FILL FILL_41_DFFSR_88 ( );
FILL FILL_42_DFFSR_88 ( );
FILL FILL_43_DFFSR_88 ( );
FILL FILL_44_DFFSR_88 ( );
FILL FILL_45_DFFSR_88 ( );
FILL FILL_46_DFFSR_88 ( );
FILL FILL_47_DFFSR_88 ( );
FILL FILL_48_DFFSR_88 ( );
FILL FILL_49_DFFSR_88 ( );
FILL FILL_50_DFFSR_88 ( );
FILL FILL_0_AOI21X1_40 ( );
FILL FILL_1_AOI21X1_40 ( );
FILL FILL_2_AOI21X1_40 ( );
FILL FILL_3_AOI21X1_40 ( );
FILL FILL_4_AOI21X1_40 ( );
FILL FILL_5_AOI21X1_40 ( );
FILL FILL_6_AOI21X1_40 ( );
FILL FILL_7_AOI21X1_40 ( );
FILL FILL_8_AOI21X1_40 ( );
FILL FILL_0_INVX1_74 ( );
FILL FILL_1_INVX1_74 ( );
FILL FILL_2_INVX1_74 ( );
FILL FILL_3_INVX1_74 ( );
FILL FILL_4_INVX1_74 ( );
FILL FILL_0_OAI21X1_65 ( );
FILL FILL_1_OAI21X1_65 ( );
FILL FILL_2_OAI21X1_65 ( );
FILL FILL_3_OAI21X1_65 ( );
FILL FILL_4_OAI21X1_65 ( );
FILL FILL_5_OAI21X1_65 ( );
FILL FILL_6_OAI21X1_65 ( );
FILL FILL_7_OAI21X1_65 ( );
FILL FILL_8_OAI21X1_65 ( );
FILL FILL_0_NAND2X1_65 ( );
FILL FILL_1_NAND2X1_65 ( );
FILL FILL_2_NAND2X1_65 ( );
FILL FILL_3_NAND2X1_65 ( );
FILL FILL_4_NAND2X1_65 ( );
FILL FILL_5_NAND2X1_65 ( );
FILL FILL_6_NAND2X1_65 ( );
FILL FILL_0_DFFSR_139 ( );
FILL FILL_1_DFFSR_139 ( );
FILL FILL_2_DFFSR_139 ( );
FILL FILL_3_DFFSR_139 ( );
FILL FILL_4_DFFSR_139 ( );
FILL FILL_5_DFFSR_139 ( );
FILL FILL_6_DFFSR_139 ( );
FILL FILL_7_DFFSR_139 ( );
FILL FILL_8_DFFSR_139 ( );
FILL FILL_9_DFFSR_139 ( );
FILL FILL_10_DFFSR_139 ( );
FILL FILL_11_DFFSR_139 ( );
FILL FILL_12_DFFSR_139 ( );
FILL FILL_13_DFFSR_139 ( );
FILL FILL_14_DFFSR_139 ( );
FILL FILL_15_DFFSR_139 ( );
FILL FILL_16_DFFSR_139 ( );
FILL FILL_17_DFFSR_139 ( );
FILL FILL_18_DFFSR_139 ( );
FILL FILL_19_DFFSR_139 ( );
FILL FILL_20_DFFSR_139 ( );
FILL FILL_21_DFFSR_139 ( );
FILL FILL_22_DFFSR_139 ( );
FILL FILL_23_DFFSR_139 ( );
FILL FILL_24_DFFSR_139 ( );
FILL FILL_25_DFFSR_139 ( );
FILL FILL_26_DFFSR_139 ( );
FILL FILL_27_DFFSR_139 ( );
FILL FILL_28_DFFSR_139 ( );
FILL FILL_29_DFFSR_139 ( );
FILL FILL_30_DFFSR_139 ( );
FILL FILL_31_DFFSR_139 ( );
FILL FILL_32_DFFSR_139 ( );
FILL FILL_33_DFFSR_139 ( );
FILL FILL_34_DFFSR_139 ( );
FILL FILL_35_DFFSR_139 ( );
FILL FILL_36_DFFSR_139 ( );
FILL FILL_37_DFFSR_139 ( );
FILL FILL_38_DFFSR_139 ( );
FILL FILL_39_DFFSR_139 ( );
FILL FILL_40_DFFSR_139 ( );
FILL FILL_41_DFFSR_139 ( );
FILL FILL_42_DFFSR_139 ( );
FILL FILL_43_DFFSR_139 ( );
FILL FILL_44_DFFSR_139 ( );
FILL FILL_45_DFFSR_139 ( );
FILL FILL_46_DFFSR_139 ( );
FILL FILL_47_DFFSR_139 ( );
FILL FILL_48_DFFSR_139 ( );
FILL FILL_49_DFFSR_139 ( );
FILL FILL_50_DFFSR_139 ( );
FILL FILL_51_DFFSR_139 ( );
FILL FILL_0_OAI21X1_32 ( );
FILL FILL_1_OAI21X1_32 ( );
FILL FILL_2_OAI21X1_32 ( );
FILL FILL_3_OAI21X1_32 ( );
FILL FILL_4_OAI21X1_32 ( );
FILL FILL_5_OAI21X1_32 ( );
FILL FILL_6_OAI21X1_32 ( );
FILL FILL_7_OAI21X1_32 ( );
FILL FILL_8_OAI21X1_32 ( );
FILL FILL_0_NAND2X1_42 ( );
FILL FILL_1_NAND2X1_42 ( );
FILL FILL_2_NAND2X1_42 ( );
FILL FILL_3_NAND2X1_42 ( );
FILL FILL_4_NAND2X1_42 ( );
FILL FILL_5_NAND2X1_42 ( );
FILL FILL_6_NAND2X1_42 ( );
FILL FILL_0_OAI21X1_48 ( );
FILL FILL_1_OAI21X1_48 ( );
FILL FILL_2_OAI21X1_48 ( );
FILL FILL_3_OAI21X1_48 ( );
FILL FILL_4_OAI21X1_48 ( );
FILL FILL_5_OAI21X1_48 ( );
FILL FILL_6_OAI21X1_48 ( );
FILL FILL_7_OAI21X1_48 ( );
FILL FILL_8_OAI21X1_48 ( );
FILL FILL_0_INVX1_54 ( );
FILL FILL_1_INVX1_54 ( );
FILL FILL_2_INVX1_54 ( );
FILL FILL_3_INVX1_54 ( );
FILL FILL_4_INVX1_54 ( );
FILL FILL_0_OAI22X1_10 ( );
FILL FILL_1_OAI22X1_10 ( );
FILL FILL_2_OAI22X1_10 ( );
FILL FILL_3_OAI22X1_10 ( );
FILL FILL_4_OAI22X1_10 ( );
FILL FILL_5_OAI22X1_10 ( );
FILL FILL_6_OAI22X1_10 ( );
FILL FILL_7_OAI22X1_10 ( );
FILL FILL_8_OAI22X1_10 ( );
FILL FILL_9_OAI22X1_10 ( );
FILL FILL_10_OAI22X1_10 ( );
FILL FILL_11_OAI22X1_10 ( );
FILL FILL_0_NOR2X1_14 ( );
FILL FILL_1_NOR2X1_14 ( );
FILL FILL_2_NOR2X1_14 ( );
FILL FILL_3_NOR2X1_14 ( );
FILL FILL_4_NOR2X1_14 ( );
FILL FILL_5_NOR2X1_14 ( );
FILL FILL_6_NOR2X1_14 ( );
FILL FILL_0_OAI22X1_11 ( );
FILL FILL_1_OAI22X1_11 ( );
FILL FILL_2_OAI22X1_11 ( );
FILL FILL_3_OAI22X1_11 ( );
FILL FILL_4_OAI22X1_11 ( );
FILL FILL_5_OAI22X1_11 ( );
FILL FILL_6_OAI22X1_11 ( );
FILL FILL_7_OAI22X1_11 ( );
FILL FILL_8_OAI22X1_11 ( );
FILL FILL_9_OAI22X1_11 ( );
FILL FILL_10_OAI22X1_11 ( );
FILL FILL_11_OAI22X1_11 ( );
FILL FILL_0_INVX1_277 ( );
FILL FILL_1_INVX1_277 ( );
FILL FILL_2_INVX1_277 ( );
FILL FILL_3_INVX1_277 ( );
FILL FILL_0_INVX1_278 ( );
FILL FILL_1_INVX1_278 ( );
FILL FILL_2_INVX1_278 ( );
FILL FILL_3_INVX1_278 ( );
FILL FILL_4_INVX1_278 ( );
FILL FILL_0_OAI22X1_14 ( );
FILL FILL_1_OAI22X1_14 ( );
FILL FILL_2_OAI22X1_14 ( );
FILL FILL_3_OAI22X1_14 ( );
FILL FILL_4_OAI22X1_14 ( );
FILL FILL_5_OAI22X1_14 ( );
FILL FILL_6_OAI22X1_14 ( );
FILL FILL_7_OAI22X1_14 ( );
FILL FILL_8_OAI22X1_14 ( );
FILL FILL_9_OAI22X1_14 ( );
FILL FILL_10_OAI22X1_14 ( );
FILL FILL_11_OAI22X1_14 ( );
FILL FILL_0_DFFSR_58 ( );
FILL FILL_1_DFFSR_58 ( );
FILL FILL_2_DFFSR_58 ( );
FILL FILL_3_DFFSR_58 ( );
FILL FILL_4_DFFSR_58 ( );
FILL FILL_5_DFFSR_58 ( );
FILL FILL_6_DFFSR_58 ( );
FILL FILL_7_DFFSR_58 ( );
FILL FILL_8_DFFSR_58 ( );
FILL FILL_9_DFFSR_58 ( );
FILL FILL_10_DFFSR_58 ( );
FILL FILL_11_DFFSR_58 ( );
FILL FILL_12_DFFSR_58 ( );
FILL FILL_13_DFFSR_58 ( );
FILL FILL_14_DFFSR_58 ( );
FILL FILL_15_DFFSR_58 ( );
FILL FILL_16_DFFSR_58 ( );
FILL FILL_17_DFFSR_58 ( );
FILL FILL_18_DFFSR_58 ( );
FILL FILL_19_DFFSR_58 ( );
FILL FILL_20_DFFSR_58 ( );
FILL FILL_21_DFFSR_58 ( );
FILL FILL_22_DFFSR_58 ( );
FILL FILL_23_DFFSR_58 ( );
FILL FILL_24_DFFSR_58 ( );
FILL FILL_25_DFFSR_58 ( );
FILL FILL_26_DFFSR_58 ( );
FILL FILL_27_DFFSR_58 ( );
FILL FILL_28_DFFSR_58 ( );
FILL FILL_29_DFFSR_58 ( );
FILL FILL_30_DFFSR_58 ( );
FILL FILL_31_DFFSR_58 ( );
FILL FILL_32_DFFSR_58 ( );
FILL FILL_33_DFFSR_58 ( );
FILL FILL_34_DFFSR_58 ( );
FILL FILL_35_DFFSR_58 ( );
FILL FILL_36_DFFSR_58 ( );
FILL FILL_37_DFFSR_58 ( );
FILL FILL_38_DFFSR_58 ( );
FILL FILL_39_DFFSR_58 ( );
FILL FILL_40_DFFSR_58 ( );
FILL FILL_41_DFFSR_58 ( );
FILL FILL_42_DFFSR_58 ( );
FILL FILL_43_DFFSR_58 ( );
FILL FILL_44_DFFSR_58 ( );
FILL FILL_45_DFFSR_58 ( );
FILL FILL_46_DFFSR_58 ( );
FILL FILL_47_DFFSR_58 ( );
FILL FILL_48_DFFSR_58 ( );
FILL FILL_49_DFFSR_58 ( );
FILL FILL_50_DFFSR_58 ( );
FILL FILL_0_NAND2X1_29 ( );
FILL FILL_1_NAND2X1_29 ( );
FILL FILL_2_NAND2X1_29 ( );
FILL FILL_3_NAND2X1_29 ( );
FILL FILL_4_NAND2X1_29 ( );
FILL FILL_5_NAND2X1_29 ( );
FILL FILL_6_NAND2X1_29 ( );
FILL FILL_0_DFFSR_3 ( );
FILL FILL_1_DFFSR_3 ( );
FILL FILL_2_DFFSR_3 ( );
FILL FILL_3_DFFSR_3 ( );
FILL FILL_4_DFFSR_3 ( );
FILL FILL_5_DFFSR_3 ( );
FILL FILL_6_DFFSR_3 ( );
FILL FILL_7_DFFSR_3 ( );
FILL FILL_8_DFFSR_3 ( );
FILL FILL_9_DFFSR_3 ( );
FILL FILL_10_DFFSR_3 ( );
FILL FILL_11_DFFSR_3 ( );
FILL FILL_12_DFFSR_3 ( );
FILL FILL_13_DFFSR_3 ( );
FILL FILL_14_DFFSR_3 ( );
FILL FILL_15_DFFSR_3 ( );
FILL FILL_16_DFFSR_3 ( );
FILL FILL_17_DFFSR_3 ( );
FILL FILL_18_DFFSR_3 ( );
FILL FILL_19_DFFSR_3 ( );
FILL FILL_20_DFFSR_3 ( );
FILL FILL_21_DFFSR_3 ( );
FILL FILL_22_DFFSR_3 ( );
FILL FILL_23_DFFSR_3 ( );
FILL FILL_24_DFFSR_3 ( );
FILL FILL_25_DFFSR_3 ( );
FILL FILL_26_DFFSR_3 ( );
FILL FILL_27_DFFSR_3 ( );
FILL FILL_28_DFFSR_3 ( );
FILL FILL_29_DFFSR_3 ( );
FILL FILL_30_DFFSR_3 ( );
FILL FILL_31_DFFSR_3 ( );
FILL FILL_32_DFFSR_3 ( );
FILL FILL_33_DFFSR_3 ( );
FILL FILL_34_DFFSR_3 ( );
FILL FILL_35_DFFSR_3 ( );
FILL FILL_36_DFFSR_3 ( );
FILL FILL_37_DFFSR_3 ( );
FILL FILL_38_DFFSR_3 ( );
FILL FILL_39_DFFSR_3 ( );
FILL FILL_40_DFFSR_3 ( );
FILL FILL_41_DFFSR_3 ( );
FILL FILL_42_DFFSR_3 ( );
FILL FILL_43_DFFSR_3 ( );
FILL FILL_44_DFFSR_3 ( );
FILL FILL_45_DFFSR_3 ( );
FILL FILL_46_DFFSR_3 ( );
FILL FILL_47_DFFSR_3 ( );
FILL FILL_48_DFFSR_3 ( );
FILL FILL_49_DFFSR_3 ( );
FILL FILL_50_DFFSR_3 ( );
FILL FILL_0_OAI21X1_163 ( );
FILL FILL_1_OAI21X1_163 ( );
FILL FILL_2_OAI21X1_163 ( );
FILL FILL_3_OAI21X1_163 ( );
FILL FILL_4_OAI21X1_163 ( );
FILL FILL_5_OAI21X1_163 ( );
FILL FILL_6_OAI21X1_163 ( );
FILL FILL_7_OAI21X1_163 ( );
FILL FILL_8_OAI21X1_163 ( );
FILL FILL_0_INVX1_197 ( );
FILL FILL_1_INVX1_197 ( );
FILL FILL_2_INVX1_197 ( );
FILL FILL_3_INVX1_197 ( );
FILL FILL_4_INVX1_197 ( );
FILL FILL_0_OAI21X1_244 ( );
FILL FILL_1_OAI21X1_244 ( );
FILL FILL_2_OAI21X1_244 ( );
FILL FILL_3_OAI21X1_244 ( );
FILL FILL_4_OAI21X1_244 ( );
FILL FILL_5_OAI21X1_244 ( );
FILL FILL_6_OAI21X1_244 ( );
FILL FILL_7_OAI21X1_244 ( );
FILL FILL_8_OAI21X1_244 ( );
FILL FILL_9_OAI21X1_244 ( );
FILL FILL_0_OAI21X1_166 ( );
FILL FILL_1_OAI21X1_166 ( );
FILL FILL_2_OAI21X1_166 ( );
FILL FILL_3_OAI21X1_166 ( );
FILL FILL_4_OAI21X1_166 ( );
FILL FILL_5_OAI21X1_166 ( );
FILL FILL_6_OAI21X1_166 ( );
FILL FILL_7_OAI21X1_166 ( );
FILL FILL_8_OAI21X1_166 ( );
FILL FILL_0_NAND2X1_266 ( );
FILL FILL_1_NAND2X1_266 ( );
FILL FILL_2_NAND2X1_266 ( );
FILL FILL_3_NAND2X1_266 ( );
FILL FILL_4_NAND2X1_266 ( );
FILL FILL_5_NAND2X1_266 ( );
FILL FILL_6_NAND2X1_266 ( );
FILL FILL_0_OAI21X1_255 ( );
FILL FILL_1_OAI21X1_255 ( );
FILL FILL_2_OAI21X1_255 ( );
FILL FILL_3_OAI21X1_255 ( );
FILL FILL_4_OAI21X1_255 ( );
FILL FILL_5_OAI21X1_255 ( );
FILL FILL_6_OAI21X1_255 ( );
FILL FILL_7_OAI21X1_255 ( );
FILL FILL_8_OAI21X1_255 ( );
FILL FILL_0_INVX1_418 ( );
FILL FILL_1_INVX1_418 ( );
FILL FILL_2_INVX1_418 ( );
FILL FILL_3_INVX1_418 ( );
FILL FILL_4_INVX1_418 ( );
FILL FILL_0_NAND2X1_255 ( );
FILL FILL_1_NAND2X1_255 ( );
FILL FILL_2_NAND2X1_255 ( );
FILL FILL_3_NAND2X1_255 ( );
FILL FILL_4_NAND2X1_255 ( );
FILL FILL_5_NAND2X1_255 ( );
FILL FILL_6_NAND2X1_255 ( );
FILL FILL_0_OAI21X1_87 ( );
FILL FILL_1_OAI21X1_87 ( );
FILL FILL_2_OAI21X1_87 ( );
FILL FILL_3_OAI21X1_87 ( );
FILL FILL_4_OAI21X1_87 ( );
FILL FILL_5_OAI21X1_87 ( );
FILL FILL_6_OAI21X1_87 ( );
FILL FILL_7_OAI21X1_87 ( );
FILL FILL_8_OAI21X1_87 ( );
FILL FILL_9_OAI21X1_87 ( );
FILL FILL_0_INVX1_98 ( );
FILL FILL_1_INVX1_98 ( );
FILL FILL_2_INVX1_98 ( );
FILL FILL_3_INVX1_98 ( );
FILL FILL_0_INVX1_97 ( );
FILL FILL_1_INVX1_97 ( );
FILL FILL_2_INVX1_97 ( );
FILL FILL_3_INVX1_97 ( );
FILL FILL_0_OAI21X1_112 ( );
FILL FILL_1_OAI21X1_112 ( );
FILL FILL_2_OAI21X1_112 ( );
FILL FILL_3_OAI21X1_112 ( );
FILL FILL_4_OAI21X1_112 ( );
FILL FILL_5_OAI21X1_112 ( );
FILL FILL_6_OAI21X1_112 ( );
FILL FILL_7_OAI21X1_112 ( );
FILL FILL_8_OAI21X1_112 ( );
FILL FILL_0_NAND2X1_112 ( );
FILL FILL_1_NAND2X1_112 ( );
FILL FILL_2_NAND2X1_112 ( );
FILL FILL_3_NAND2X1_112 ( );
FILL FILL_4_NAND2X1_112 ( );
FILL FILL_5_NAND2X1_112 ( );
FILL FILL_6_NAND2X1_112 ( );
FILL FILL_0_DFFSR_104 ( );
FILL FILL_1_DFFSR_104 ( );
FILL FILL_2_DFFSR_104 ( );
FILL FILL_3_DFFSR_104 ( );
FILL FILL_4_DFFSR_104 ( );
FILL FILL_5_DFFSR_104 ( );
FILL FILL_6_DFFSR_104 ( );
FILL FILL_7_DFFSR_104 ( );
FILL FILL_8_DFFSR_104 ( );
FILL FILL_9_DFFSR_104 ( );
FILL FILL_10_DFFSR_104 ( );
FILL FILL_11_DFFSR_104 ( );
FILL FILL_12_DFFSR_104 ( );
FILL FILL_13_DFFSR_104 ( );
FILL FILL_14_DFFSR_104 ( );
FILL FILL_15_DFFSR_104 ( );
FILL FILL_16_DFFSR_104 ( );
FILL FILL_17_DFFSR_104 ( );
FILL FILL_18_DFFSR_104 ( );
FILL FILL_19_DFFSR_104 ( );
FILL FILL_20_DFFSR_104 ( );
FILL FILL_21_DFFSR_104 ( );
FILL FILL_22_DFFSR_104 ( );
FILL FILL_23_DFFSR_104 ( );
FILL FILL_24_DFFSR_104 ( );
FILL FILL_25_DFFSR_104 ( );
FILL FILL_26_DFFSR_104 ( );
FILL FILL_27_DFFSR_104 ( );
FILL FILL_28_DFFSR_104 ( );
FILL FILL_29_DFFSR_104 ( );
FILL FILL_30_DFFSR_104 ( );
FILL FILL_31_DFFSR_104 ( );
FILL FILL_32_DFFSR_104 ( );
FILL FILL_33_DFFSR_104 ( );
FILL FILL_34_DFFSR_104 ( );
FILL FILL_35_DFFSR_104 ( );
FILL FILL_36_DFFSR_104 ( );
FILL FILL_37_DFFSR_104 ( );
FILL FILL_38_DFFSR_104 ( );
FILL FILL_39_DFFSR_104 ( );
FILL FILL_40_DFFSR_104 ( );
FILL FILL_41_DFFSR_104 ( );
FILL FILL_42_DFFSR_104 ( );
FILL FILL_43_DFFSR_104 ( );
FILL FILL_44_DFFSR_104 ( );
FILL FILL_45_DFFSR_104 ( );
FILL FILL_46_DFFSR_104 ( );
FILL FILL_47_DFFSR_104 ( );
FILL FILL_48_DFFSR_104 ( );
FILL FILL_49_DFFSR_104 ( );
FILL FILL_50_DFFSR_104 ( );
FILL FILL_0_INVX1_99 ( );
FILL FILL_1_INVX1_99 ( );
FILL FILL_2_INVX1_99 ( );
FILL FILL_3_INVX1_99 ( );
FILL FILL_0_INVX1_347 ( );
FILL FILL_1_INVX1_347 ( );
FILL FILL_2_INVX1_347 ( );
FILL FILL_3_INVX1_347 ( );
FILL FILL_0_OAI21X1_88 ( );
FILL FILL_1_OAI21X1_88 ( );
FILL FILL_2_OAI21X1_88 ( );
FILL FILL_3_OAI21X1_88 ( );
FILL FILL_4_OAI21X1_88 ( );
FILL FILL_5_OAI21X1_88 ( );
FILL FILL_6_OAI21X1_88 ( );
FILL FILL_7_OAI21X1_88 ( );
FILL FILL_8_OAI21X1_88 ( );
FILL FILL_9_OAI21X1_88 ( );
FILL FILL_0_OAI21X1_75 ( );
FILL FILL_1_OAI21X1_75 ( );
FILL FILL_2_OAI21X1_75 ( );
FILL FILL_3_OAI21X1_75 ( );
FILL FILL_4_OAI21X1_75 ( );
FILL FILL_5_OAI21X1_75 ( );
FILL FILL_6_OAI21X1_75 ( );
FILL FILL_7_OAI21X1_75 ( );
FILL FILL_8_OAI21X1_75 ( );
FILL FILL_0_INVX1_348 ( );
FILL FILL_1_INVX1_348 ( );
FILL FILL_2_INVX1_348 ( );
FILL FILL_3_INVX1_348 ( );
FILL FILL_4_INVX1_348 ( );
FILL FILL_0_NAND2X1_75 ( );
FILL FILL_1_NAND2X1_75 ( );
FILL FILL_2_NAND2X1_75 ( );
FILL FILL_3_NAND2X1_75 ( );
FILL FILL_4_NAND2X1_75 ( );
FILL FILL_5_NAND2X1_75 ( );
FILL FILL_6_NAND2X1_75 ( );
FILL FILL_0_OAI21X1_239 ( );
FILL FILL_1_OAI21X1_239 ( );
FILL FILL_2_OAI21X1_239 ( );
FILL FILL_3_OAI21X1_239 ( );
FILL FILL_4_OAI21X1_239 ( );
FILL FILL_5_OAI21X1_239 ( );
FILL FILL_6_OAI21X1_239 ( );
FILL FILL_7_OAI21X1_239 ( );
FILL FILL_8_OAI21X1_239 ( );
FILL FILL_0_DFFPOSX1_11 ( );
FILL FILL_1_DFFPOSX1_11 ( );
FILL FILL_2_DFFPOSX1_11 ( );
FILL FILL_3_DFFPOSX1_11 ( );
FILL FILL_4_DFFPOSX1_11 ( );
FILL FILL_5_DFFPOSX1_11 ( );
FILL FILL_6_DFFPOSX1_11 ( );
FILL FILL_7_DFFPOSX1_11 ( );
FILL FILL_8_DFFPOSX1_11 ( );
FILL FILL_9_DFFPOSX1_11 ( );
FILL FILL_10_DFFPOSX1_11 ( );
FILL FILL_11_DFFPOSX1_11 ( );
FILL FILL_12_DFFPOSX1_11 ( );
FILL FILL_13_DFFPOSX1_11 ( );
FILL FILL_14_DFFPOSX1_11 ( );
FILL FILL_15_DFFPOSX1_11 ( );
FILL FILL_16_DFFPOSX1_11 ( );
FILL FILL_17_DFFPOSX1_11 ( );
FILL FILL_18_DFFPOSX1_11 ( );
FILL FILL_19_DFFPOSX1_11 ( );
FILL FILL_20_DFFPOSX1_11 ( );
FILL FILL_21_DFFPOSX1_11 ( );
FILL FILL_22_DFFPOSX1_11 ( );
FILL FILL_23_DFFPOSX1_11 ( );
FILL FILL_24_DFFPOSX1_11 ( );
FILL FILL_25_DFFPOSX1_11 ( );
FILL FILL_26_DFFPOSX1_11 ( );
FILL FILL_27_DFFPOSX1_11 ( );
FILL FILL_0_INVX1_147 ( );
FILL FILL_1_INVX1_147 ( );
FILL FILL_2_INVX1_147 ( );
FILL FILL_3_INVX1_147 ( );
FILL FILL_0_OAI21X1_130 ( );
FILL FILL_1_OAI21X1_130 ( );
FILL FILL_2_OAI21X1_130 ( );
FILL FILL_3_OAI21X1_130 ( );
FILL FILL_4_OAI21X1_130 ( );
FILL FILL_5_OAI21X1_130 ( );
FILL FILL_6_OAI21X1_130 ( );
FILL FILL_7_OAI21X1_130 ( );
FILL FILL_8_OAI21X1_130 ( );
FILL FILL_9_OAI21X1_130 ( );
FILL FILL_0_NAND2X1_130 ( );
FILL FILL_1_NAND2X1_130 ( );
FILL FILL_2_NAND2X1_130 ( );
FILL FILL_3_NAND2X1_130 ( );
FILL FILL_4_NAND2X1_130 ( );
FILL FILL_5_NAND2X1_130 ( );
FILL FILL_6_NAND2X1_130 ( );
FILL FILL_0_INVX1_146 ( );
FILL FILL_1_INVX1_146 ( );
FILL FILL_2_INVX1_146 ( );
FILL FILL_3_INVX1_146 ( );
FILL FILL_0_OAI21X1_129 ( );
FILL FILL_1_OAI21X1_129 ( );
FILL FILL_2_OAI21X1_129 ( );
FILL FILL_3_OAI21X1_129 ( );
FILL FILL_4_OAI21X1_129 ( );
FILL FILL_5_OAI21X1_129 ( );
FILL FILL_6_OAI21X1_129 ( );
FILL FILL_7_OAI21X1_129 ( );
FILL FILL_8_OAI21X1_129 ( );
FILL FILL_9_OAI21X1_129 ( );
FILL FILL_0_OAI21X1_132 ( );
FILL FILL_1_OAI21X1_132 ( );
FILL FILL_2_OAI21X1_132 ( );
FILL FILL_3_OAI21X1_132 ( );
FILL FILL_4_OAI21X1_132 ( );
FILL FILL_5_OAI21X1_132 ( );
FILL FILL_6_OAI21X1_132 ( );
FILL FILL_7_OAI21X1_132 ( );
FILL FILL_8_OAI21X1_132 ( );
FILL FILL_9_OAI21X1_132 ( );
FILL FILL_0_NAND2X1_129 ( );
FILL FILL_1_NAND2X1_129 ( );
FILL FILL_2_NAND2X1_129 ( );
FILL FILL_3_NAND2X1_129 ( );
FILL FILL_4_NAND2X1_129 ( );
FILL FILL_5_NAND2X1_129 ( );
FILL FILL_6_NAND2X1_129 ( );
FILL FILL_0_DFFSR_48 ( );
FILL FILL_1_DFFSR_48 ( );
FILL FILL_2_DFFSR_48 ( );
FILL FILL_3_DFFSR_48 ( );
FILL FILL_4_DFFSR_48 ( );
FILL FILL_5_DFFSR_48 ( );
FILL FILL_6_DFFSR_48 ( );
FILL FILL_7_DFFSR_48 ( );
FILL FILL_8_DFFSR_48 ( );
FILL FILL_9_DFFSR_48 ( );
FILL FILL_10_DFFSR_48 ( );
FILL FILL_11_DFFSR_48 ( );
FILL FILL_12_DFFSR_48 ( );
FILL FILL_13_DFFSR_48 ( );
FILL FILL_14_DFFSR_48 ( );
FILL FILL_15_DFFSR_48 ( );
FILL FILL_16_DFFSR_48 ( );
FILL FILL_17_DFFSR_48 ( );
FILL FILL_18_DFFSR_48 ( );
FILL FILL_19_DFFSR_48 ( );
FILL FILL_20_DFFSR_48 ( );
FILL FILL_21_DFFSR_48 ( );
FILL FILL_22_DFFSR_48 ( );
FILL FILL_23_DFFSR_48 ( );
FILL FILL_24_DFFSR_48 ( );
FILL FILL_25_DFFSR_48 ( );
FILL FILL_26_DFFSR_48 ( );
FILL FILL_27_DFFSR_48 ( );
FILL FILL_28_DFFSR_48 ( );
FILL FILL_29_DFFSR_48 ( );
FILL FILL_30_DFFSR_48 ( );
FILL FILL_31_DFFSR_48 ( );
FILL FILL_32_DFFSR_48 ( );
FILL FILL_33_DFFSR_48 ( );
FILL FILL_34_DFFSR_48 ( );
FILL FILL_35_DFFSR_48 ( );
FILL FILL_36_DFFSR_48 ( );
FILL FILL_37_DFFSR_48 ( );
FILL FILL_38_DFFSR_48 ( );
FILL FILL_39_DFFSR_48 ( );
FILL FILL_40_DFFSR_48 ( );
FILL FILL_41_DFFSR_48 ( );
FILL FILL_42_DFFSR_48 ( );
FILL FILL_43_DFFSR_48 ( );
FILL FILL_44_DFFSR_48 ( );
FILL FILL_45_DFFSR_48 ( );
FILL FILL_46_DFFSR_48 ( );
FILL FILL_47_DFFSR_48 ( );
FILL FILL_48_DFFSR_48 ( );
FILL FILL_49_DFFSR_48 ( );
FILL FILL_50_DFFSR_48 ( );
FILL FILL_51_DFFSR_48 ( );
FILL FILL_0_INVX1_283 ( );
FILL FILL_1_INVX1_283 ( );
FILL FILL_2_INVX1_283 ( );
FILL FILL_3_INVX1_283 ( );
FILL FILL_0_OAI22X1_15 ( );
FILL FILL_1_OAI22X1_15 ( );
FILL FILL_2_OAI22X1_15 ( );
FILL FILL_3_OAI22X1_15 ( );
FILL FILL_4_OAI22X1_15 ( );
FILL FILL_5_OAI22X1_15 ( );
FILL FILL_6_OAI22X1_15 ( );
FILL FILL_7_OAI22X1_15 ( );
FILL FILL_8_OAI22X1_15 ( );
FILL FILL_9_OAI22X1_15 ( );
FILL FILL_10_OAI22X1_15 ( );
FILL FILL_11_OAI22X1_15 ( );
FILL FILL_0_NOR2X1_17 ( );
FILL FILL_1_NOR2X1_17 ( );
FILL FILL_2_NOR2X1_17 ( );
FILL FILL_3_NOR2X1_17 ( );
FILL FILL_4_NOR2X1_17 ( );
FILL FILL_5_NOR2X1_17 ( );
FILL FILL_6_NOR2X1_17 ( );
FILL FILL_0_OAI22X1_16 ( );
FILL FILL_1_OAI22X1_16 ( );
FILL FILL_2_OAI22X1_16 ( );
FILL FILL_3_OAI22X1_16 ( );
FILL FILL_4_OAI22X1_16 ( );
FILL FILL_5_OAI22X1_16 ( );
FILL FILL_6_OAI22X1_16 ( );
FILL FILL_7_OAI22X1_16 ( );
FILL FILL_8_OAI22X1_16 ( );
FILL FILL_9_OAI22X1_16 ( );
FILL FILL_10_OAI22X1_16 ( );
FILL FILL_11_OAI22X1_16 ( );
FILL FILL_0_INVX1_288 ( );
FILL FILL_1_INVX1_288 ( );
FILL FILL_2_INVX1_288 ( );
FILL FILL_3_INVX1_288 ( );
FILL FILL_4_INVX1_288 ( );
FILL FILL_0_DFFSR_29 ( );
FILL FILL_1_DFFSR_29 ( );
FILL FILL_2_DFFSR_29 ( );
FILL FILL_3_DFFSR_29 ( );
FILL FILL_4_DFFSR_29 ( );
FILL FILL_5_DFFSR_29 ( );
FILL FILL_6_DFFSR_29 ( );
FILL FILL_7_DFFSR_29 ( );
FILL FILL_8_DFFSR_29 ( );
FILL FILL_9_DFFSR_29 ( );
FILL FILL_10_DFFSR_29 ( );
FILL FILL_11_DFFSR_29 ( );
FILL FILL_12_DFFSR_29 ( );
FILL FILL_13_DFFSR_29 ( );
FILL FILL_14_DFFSR_29 ( );
FILL FILL_15_DFFSR_29 ( );
FILL FILL_16_DFFSR_29 ( );
FILL FILL_17_DFFSR_29 ( );
FILL FILL_18_DFFSR_29 ( );
FILL FILL_19_DFFSR_29 ( );
FILL FILL_20_DFFSR_29 ( );
FILL FILL_21_DFFSR_29 ( );
FILL FILL_22_DFFSR_29 ( );
FILL FILL_23_DFFSR_29 ( );
FILL FILL_24_DFFSR_29 ( );
FILL FILL_25_DFFSR_29 ( );
FILL FILL_26_DFFSR_29 ( );
FILL FILL_27_DFFSR_29 ( );
FILL FILL_28_DFFSR_29 ( );
FILL FILL_29_DFFSR_29 ( );
FILL FILL_30_DFFSR_29 ( );
FILL FILL_31_DFFSR_29 ( );
FILL FILL_32_DFFSR_29 ( );
FILL FILL_33_DFFSR_29 ( );
FILL FILL_34_DFFSR_29 ( );
FILL FILL_35_DFFSR_29 ( );
FILL FILL_36_DFFSR_29 ( );
FILL FILL_37_DFFSR_29 ( );
FILL FILL_38_DFFSR_29 ( );
FILL FILL_39_DFFSR_29 ( );
FILL FILL_40_DFFSR_29 ( );
FILL FILL_41_DFFSR_29 ( );
FILL FILL_42_DFFSR_29 ( );
FILL FILL_43_DFFSR_29 ( );
FILL FILL_44_DFFSR_29 ( );
FILL FILL_45_DFFSR_29 ( );
FILL FILL_46_DFFSR_29 ( );
FILL FILL_47_DFFSR_29 ( );
FILL FILL_48_DFFSR_29 ( );
FILL FILL_49_DFFSR_29 ( );
FILL FILL_50_DFFSR_29 ( );
FILL FILL_51_DFFSR_29 ( );
FILL FILL_0_INVX1_4 ( );
FILL FILL_1_INVX1_4 ( );
FILL FILL_2_INVX1_4 ( );
FILL FILL_3_INVX1_4 ( );
FILL FILL_4_INVX1_4 ( );
FILL FILL_0_NAND2X1_21 ( );
FILL FILL_1_NAND2X1_21 ( );
FILL FILL_2_NAND2X1_21 ( );
FILL FILL_3_NAND2X1_21 ( );
FILL FILL_4_NAND2X1_21 ( );
FILL FILL_5_NAND2X1_21 ( );
FILL FILL_6_NAND2X1_21 ( );
FILL FILL_0_DFFSR_4 ( );
FILL FILL_1_DFFSR_4 ( );
FILL FILL_2_DFFSR_4 ( );
FILL FILL_3_DFFSR_4 ( );
FILL FILL_4_DFFSR_4 ( );
FILL FILL_5_DFFSR_4 ( );
FILL FILL_6_DFFSR_4 ( );
FILL FILL_7_DFFSR_4 ( );
FILL FILL_8_DFFSR_4 ( );
FILL FILL_9_DFFSR_4 ( );
FILL FILL_10_DFFSR_4 ( );
FILL FILL_11_DFFSR_4 ( );
FILL FILL_12_DFFSR_4 ( );
FILL FILL_13_DFFSR_4 ( );
FILL FILL_14_DFFSR_4 ( );
FILL FILL_15_DFFSR_4 ( );
FILL FILL_16_DFFSR_4 ( );
FILL FILL_17_DFFSR_4 ( );
FILL FILL_18_DFFSR_4 ( );
FILL FILL_19_DFFSR_4 ( );
FILL FILL_20_DFFSR_4 ( );
FILL FILL_21_DFFSR_4 ( );
FILL FILL_22_DFFSR_4 ( );
FILL FILL_23_DFFSR_4 ( );
FILL FILL_24_DFFSR_4 ( );
FILL FILL_25_DFFSR_4 ( );
FILL FILL_26_DFFSR_4 ( );
FILL FILL_27_DFFSR_4 ( );
FILL FILL_28_DFFSR_4 ( );
FILL FILL_29_DFFSR_4 ( );
FILL FILL_30_DFFSR_4 ( );
FILL FILL_31_DFFSR_4 ( );
FILL FILL_32_DFFSR_4 ( );
FILL FILL_33_DFFSR_4 ( );
FILL FILL_34_DFFSR_4 ( );
FILL FILL_35_DFFSR_4 ( );
FILL FILL_36_DFFSR_4 ( );
FILL FILL_37_DFFSR_4 ( );
FILL FILL_38_DFFSR_4 ( );
FILL FILL_39_DFFSR_4 ( );
FILL FILL_40_DFFSR_4 ( );
FILL FILL_41_DFFSR_4 ( );
FILL FILL_42_DFFSR_4 ( );
FILL FILL_43_DFFSR_4 ( );
FILL FILL_44_DFFSR_4 ( );
FILL FILL_45_DFFSR_4 ( );
FILL FILL_46_DFFSR_4 ( );
FILL FILL_47_DFFSR_4 ( );
FILL FILL_48_DFFSR_4 ( );
FILL FILL_49_DFFSR_4 ( );
FILL FILL_50_DFFSR_4 ( );
FILL FILL_0_INVX1_200 ( );
FILL FILL_1_INVX1_200 ( );
FILL FILL_2_INVX1_200 ( );
FILL FILL_3_INVX1_200 ( );
FILL FILL_4_INVX1_200 ( );
FILL FILL_0_NAND2X1_269 ( );
FILL FILL_1_NAND2X1_269 ( );
FILL FILL_2_NAND2X1_269 ( );
FILL FILL_3_NAND2X1_269 ( );
FILL FILL_4_NAND2X1_269 ( );
FILL FILL_5_NAND2X1_269 ( );
FILL FILL_6_NAND2X1_269 ( );
FILL FILL_0_NAND2X1_267 ( );
FILL FILL_1_NAND2X1_267 ( );
FILL FILL_2_NAND2X1_267 ( );
FILL FILL_3_NAND2X1_267 ( );
FILL FILL_4_NAND2X1_267 ( );
FILL FILL_5_NAND2X1_267 ( );
FILL FILL_6_NAND2X1_267 ( );
FILL FILL_0_NAND2X1_86 ( );
FILL FILL_1_NAND2X1_86 ( );
FILL FILL_2_NAND2X1_86 ( );
FILL FILL_3_NAND2X1_86 ( );
FILL FILL_4_NAND2X1_86 ( );
FILL FILL_5_NAND2X1_86 ( );
FILL FILL_6_NAND2X1_86 ( );
FILL FILL_0_OAI21X1_86 ( );
FILL FILL_1_OAI21X1_86 ( );
FILL FILL_2_OAI21X1_86 ( );
FILL FILL_3_OAI21X1_86 ( );
FILL FILL_4_OAI21X1_86 ( );
FILL FILL_5_OAI21X1_86 ( );
FILL FILL_6_OAI21X1_86 ( );
FILL FILL_7_OAI21X1_86 ( );
FILL FILL_8_OAI21X1_86 ( );
FILL FILL_9_OAI21X1_86 ( );
FILL FILL_0_OAI21X1_96 ( );
FILL FILL_1_OAI21X1_96 ( );
FILL FILL_2_OAI21X1_96 ( );
FILL FILL_3_OAI21X1_96 ( );
FILL FILL_4_OAI21X1_96 ( );
FILL FILL_5_OAI21X1_96 ( );
FILL FILL_6_OAI21X1_96 ( );
FILL FILL_7_OAI21X1_96 ( );
FILL FILL_8_OAI21X1_96 ( );
FILL FILL_0_NAND2X1_96 ( );
FILL FILL_1_NAND2X1_96 ( );
FILL FILL_2_NAND2X1_96 ( );
FILL FILL_3_NAND2X1_96 ( );
FILL FILL_4_NAND2X1_96 ( );
FILL FILL_5_NAND2X1_96 ( );
FILL FILL_6_NAND2X1_96 ( );
FILL FILL_0_INVX1_105 ( );
FILL FILL_1_INVX1_105 ( );
FILL FILL_2_INVX1_105 ( );
FILL FILL_3_INVX1_105 ( );
FILL FILL_4_INVX1_105 ( );
FILL FILL_0_OAI21X1_93 ( );
FILL FILL_1_OAI21X1_93 ( );
FILL FILL_2_OAI21X1_93 ( );
FILL FILL_3_OAI21X1_93 ( );
FILL FILL_4_OAI21X1_93 ( );
FILL FILL_5_OAI21X1_93 ( );
FILL FILL_6_OAI21X1_93 ( );
FILL FILL_7_OAI21X1_93 ( );
FILL FILL_8_OAI21X1_93 ( );
FILL FILL_0_NAND2X1_104 ( );
FILL FILL_1_NAND2X1_104 ( );
FILL FILL_2_NAND2X1_104 ( );
FILL FILL_3_NAND2X1_104 ( );
FILL FILL_4_NAND2X1_104 ( );
FILL FILL_5_NAND2X1_104 ( );
FILL FILL_6_NAND2X1_104 ( );
FILL FILL_0_INVX1_117 ( );
FILL FILL_1_INVX1_117 ( );
FILL FILL_2_INVX1_117 ( );
FILL FILL_3_INVX1_117 ( );
FILL FILL_0_OAI21X1_104 ( );
FILL FILL_1_OAI21X1_104 ( );
FILL FILL_2_OAI21X1_104 ( );
FILL FILL_3_OAI21X1_104 ( );
FILL FILL_4_OAI21X1_104 ( );
FILL FILL_5_OAI21X1_104 ( );
FILL FILL_6_OAI21X1_104 ( );
FILL FILL_7_OAI21X1_104 ( );
FILL FILL_8_OAI21X1_104 ( );
FILL FILL_9_OAI21X1_104 ( );
FILL FILL_0_INVX1_75 ( );
FILL FILL_1_INVX1_75 ( );
FILL FILL_2_INVX1_75 ( );
FILL FILL_3_INVX1_75 ( );
FILL FILL_4_INVX1_75 ( );
FILL FILL_0_OAI21X1_66 ( );
FILL FILL_1_OAI21X1_66 ( );
FILL FILL_2_OAI21X1_66 ( );
FILL FILL_3_OAI21X1_66 ( );
FILL FILL_4_OAI21X1_66 ( );
FILL FILL_5_OAI21X1_66 ( );
FILL FILL_6_OAI21X1_66 ( );
FILL FILL_7_OAI21X1_66 ( );
FILL FILL_8_OAI21X1_66 ( );
FILL FILL_0_DFFSR_75 ( );
FILL FILL_1_DFFSR_75 ( );
FILL FILL_2_DFFSR_75 ( );
FILL FILL_3_DFFSR_75 ( );
FILL FILL_4_DFFSR_75 ( );
FILL FILL_5_DFFSR_75 ( );
FILL FILL_6_DFFSR_75 ( );
FILL FILL_7_DFFSR_75 ( );
FILL FILL_8_DFFSR_75 ( );
FILL FILL_9_DFFSR_75 ( );
FILL FILL_10_DFFSR_75 ( );
FILL FILL_11_DFFSR_75 ( );
FILL FILL_12_DFFSR_75 ( );
FILL FILL_13_DFFSR_75 ( );
FILL FILL_14_DFFSR_75 ( );
FILL FILL_15_DFFSR_75 ( );
FILL FILL_16_DFFSR_75 ( );
FILL FILL_17_DFFSR_75 ( );
FILL FILL_18_DFFSR_75 ( );
FILL FILL_19_DFFSR_75 ( );
FILL FILL_20_DFFSR_75 ( );
FILL FILL_21_DFFSR_75 ( );
FILL FILL_22_DFFSR_75 ( );
FILL FILL_23_DFFSR_75 ( );
FILL FILL_24_DFFSR_75 ( );
FILL FILL_25_DFFSR_75 ( );
FILL FILL_26_DFFSR_75 ( );
FILL FILL_27_DFFSR_75 ( );
FILL FILL_28_DFFSR_75 ( );
FILL FILL_29_DFFSR_75 ( );
FILL FILL_30_DFFSR_75 ( );
FILL FILL_31_DFFSR_75 ( );
FILL FILL_32_DFFSR_75 ( );
FILL FILL_33_DFFSR_75 ( );
FILL FILL_34_DFFSR_75 ( );
FILL FILL_35_DFFSR_75 ( );
FILL FILL_36_DFFSR_75 ( );
FILL FILL_37_DFFSR_75 ( );
FILL FILL_38_DFFSR_75 ( );
FILL FILL_39_DFFSR_75 ( );
FILL FILL_40_DFFSR_75 ( );
FILL FILL_41_DFFSR_75 ( );
FILL FILL_42_DFFSR_75 ( );
FILL FILL_43_DFFSR_75 ( );
FILL FILL_44_DFFSR_75 ( );
FILL FILL_45_DFFSR_75 ( );
FILL FILL_46_DFFSR_75 ( );
FILL FILL_47_DFFSR_75 ( );
FILL FILL_48_DFFSR_75 ( );
FILL FILL_49_DFFSR_75 ( );
FILL FILL_50_DFFSR_75 ( );
FILL FILL_0_NAND2X1_66 ( );
FILL FILL_1_NAND2X1_66 ( );
FILL FILL_2_NAND2X1_66 ( );
FILL FILL_3_NAND2X1_66 ( );
FILL FILL_4_NAND2X1_66 ( );
FILL FILL_5_NAND2X1_66 ( );
FILL FILL_6_NAND2X1_66 ( );
FILL FILL_0_DFFSR_130 ( );
FILL FILL_1_DFFSR_130 ( );
FILL FILL_2_DFFSR_130 ( );
FILL FILL_3_DFFSR_130 ( );
FILL FILL_4_DFFSR_130 ( );
FILL FILL_5_DFFSR_130 ( );
FILL FILL_6_DFFSR_130 ( );
FILL FILL_7_DFFSR_130 ( );
FILL FILL_8_DFFSR_130 ( );
FILL FILL_9_DFFSR_130 ( );
FILL FILL_10_DFFSR_130 ( );
FILL FILL_11_DFFSR_130 ( );
FILL FILL_12_DFFSR_130 ( );
FILL FILL_13_DFFSR_130 ( );
FILL FILL_14_DFFSR_130 ( );
FILL FILL_15_DFFSR_130 ( );
FILL FILL_16_DFFSR_130 ( );
FILL FILL_17_DFFSR_130 ( );
FILL FILL_18_DFFSR_130 ( );
FILL FILL_19_DFFSR_130 ( );
FILL FILL_20_DFFSR_130 ( );
FILL FILL_21_DFFSR_130 ( );
FILL FILL_22_DFFSR_130 ( );
FILL FILL_23_DFFSR_130 ( );
FILL FILL_24_DFFSR_130 ( );
FILL FILL_25_DFFSR_130 ( );
FILL FILL_26_DFFSR_130 ( );
FILL FILL_27_DFFSR_130 ( );
FILL FILL_28_DFFSR_130 ( );
FILL FILL_29_DFFSR_130 ( );
FILL FILL_30_DFFSR_130 ( );
FILL FILL_31_DFFSR_130 ( );
FILL FILL_32_DFFSR_130 ( );
FILL FILL_33_DFFSR_130 ( );
FILL FILL_34_DFFSR_130 ( );
FILL FILL_35_DFFSR_130 ( );
FILL FILL_36_DFFSR_130 ( );
FILL FILL_37_DFFSR_130 ( );
FILL FILL_38_DFFSR_130 ( );
FILL FILL_39_DFFSR_130 ( );
FILL FILL_40_DFFSR_130 ( );
FILL FILL_41_DFFSR_130 ( );
FILL FILL_42_DFFSR_130 ( );
FILL FILL_43_DFFSR_130 ( );
FILL FILL_44_DFFSR_130 ( );
FILL FILL_45_DFFSR_130 ( );
FILL FILL_46_DFFSR_130 ( );
FILL FILL_47_DFFSR_130 ( );
FILL FILL_48_DFFSR_130 ( );
FILL FILL_49_DFFSR_130 ( );
FILL FILL_50_DFFSR_130 ( );
FILL FILL_0_INVX1_149 ( );
FILL FILL_1_INVX1_149 ( );
FILL FILL_2_INVX1_149 ( );
FILL FILL_3_INVX1_149 ( );
FILL FILL_0_CLKBUF1_13 ( );
FILL FILL_1_CLKBUF1_13 ( );
FILL FILL_2_CLKBUF1_13 ( );
FILL FILL_3_CLKBUF1_13 ( );
FILL FILL_4_CLKBUF1_13 ( );
FILL FILL_5_CLKBUF1_13 ( );
FILL FILL_6_CLKBUF1_13 ( );
FILL FILL_7_CLKBUF1_13 ( );
FILL FILL_8_CLKBUF1_13 ( );
FILL FILL_9_CLKBUF1_13 ( );
FILL FILL_10_CLKBUF1_13 ( );
FILL FILL_11_CLKBUF1_13 ( );
FILL FILL_12_CLKBUF1_13 ( );
FILL FILL_13_CLKBUF1_13 ( );
FILL FILL_14_CLKBUF1_13 ( );
FILL FILL_15_CLKBUF1_13 ( );
FILL FILL_16_CLKBUF1_13 ( );
FILL FILL_17_CLKBUF1_13 ( );
FILL FILL_18_CLKBUF1_13 ( );
FILL FILL_19_CLKBUF1_13 ( );
FILL FILL_20_CLKBUF1_13 ( );
FILL FILL_0_INVX1_279 ( );
FILL FILL_1_INVX1_279 ( );
FILL FILL_2_INVX1_279 ( );
FILL FILL_3_INVX1_279 ( );
FILL FILL_0_OAI22X1_12 ( );
FILL FILL_1_OAI22X1_12 ( );
FILL FILL_2_OAI22X1_12 ( );
FILL FILL_3_OAI22X1_12 ( );
FILL FILL_4_OAI22X1_12 ( );
FILL FILL_5_OAI22X1_12 ( );
FILL FILL_6_OAI22X1_12 ( );
FILL FILL_7_OAI22X1_12 ( );
FILL FILL_8_OAI22X1_12 ( );
FILL FILL_9_OAI22X1_12 ( );
FILL FILL_10_OAI22X1_12 ( );
FILL FILL_11_OAI22X1_12 ( );
FILL FILL_0_NAND2X1_235 ( );
FILL FILL_1_NAND2X1_235 ( );
FILL FILL_2_NAND2X1_235 ( );
FILL FILL_3_NAND2X1_235 ( );
FILL FILL_4_NAND2X1_235 ( );
FILL FILL_5_NAND2X1_235 ( );
FILL FILL_6_NAND2X1_235 ( );
FILL FILL_0_NOR2X1_15 ( );
FILL FILL_1_NOR2X1_15 ( );
FILL FILL_2_NOR2X1_15 ( );
FILL FILL_3_NOR2X1_15 ( );
FILL FILL_4_NOR2X1_15 ( );
FILL FILL_5_NOR2X1_15 ( );
FILL FILL_6_NOR2X1_15 ( );
FILL FILL_0_CLKBUF1_20 ( );
FILL FILL_1_CLKBUF1_20 ( );
FILL FILL_2_CLKBUF1_20 ( );
FILL FILL_3_CLKBUF1_20 ( );
FILL FILL_4_CLKBUF1_20 ( );
FILL FILL_5_CLKBUF1_20 ( );
FILL FILL_6_CLKBUF1_20 ( );
FILL FILL_7_CLKBUF1_20 ( );
FILL FILL_8_CLKBUF1_20 ( );
FILL FILL_9_CLKBUF1_20 ( );
FILL FILL_10_CLKBUF1_20 ( );
FILL FILL_11_CLKBUF1_20 ( );
FILL FILL_12_CLKBUF1_20 ( );
FILL FILL_13_CLKBUF1_20 ( );
FILL FILL_14_CLKBUF1_20 ( );
FILL FILL_15_CLKBUF1_20 ( );
FILL FILL_16_CLKBUF1_20 ( );
FILL FILL_17_CLKBUF1_20 ( );
FILL FILL_18_CLKBUF1_20 ( );
FILL FILL_19_CLKBUF1_20 ( );
FILL FILL_20_CLKBUF1_20 ( );
FILL FILL_0_NAND2X1_56 ( );
FILL FILL_1_NAND2X1_56 ( );
FILL FILL_2_NAND2X1_56 ( );
FILL FILL_3_NAND2X1_56 ( );
FILL FILL_4_NAND2X1_56 ( );
FILL FILL_5_NAND2X1_56 ( );
FILL FILL_6_NAND2X1_56 ( );
FILL FILL_0_INVX1_286 ( );
FILL FILL_1_INVX1_286 ( );
FILL FILL_2_INVX1_286 ( );
FILL FILL_3_INVX1_286 ( );
FILL FILL_4_INVX1_286 ( );
FILL FILL_0_OAI21X1_59 ( );
FILL FILL_1_OAI21X1_59 ( );
FILL FILL_2_OAI21X1_59 ( );
FILL FILL_3_OAI21X1_59 ( );
FILL FILL_4_OAI21X1_59 ( );
FILL FILL_5_OAI21X1_59 ( );
FILL FILL_6_OAI21X1_59 ( );
FILL FILL_7_OAI21X1_59 ( );
FILL FILL_8_OAI21X1_59 ( );
FILL FILL_9_OAI21X1_59 ( );
FILL FILL_0_INVX1_67 ( );
FILL FILL_1_INVX1_67 ( );
FILL FILL_2_INVX1_67 ( );
FILL FILL_3_INVX1_67 ( );
FILL FILL_0_INVX1_287 ( );
FILL FILL_1_INVX1_287 ( );
FILL FILL_2_INVX1_287 ( );
FILL FILL_3_INVX1_287 ( );
FILL FILL_0_DFFSR_59 ( );
FILL FILL_1_DFFSR_59 ( );
FILL FILL_2_DFFSR_59 ( );
FILL FILL_3_DFFSR_59 ( );
FILL FILL_4_DFFSR_59 ( );
FILL FILL_5_DFFSR_59 ( );
FILL FILL_6_DFFSR_59 ( );
FILL FILL_7_DFFSR_59 ( );
FILL FILL_8_DFFSR_59 ( );
FILL FILL_9_DFFSR_59 ( );
FILL FILL_10_DFFSR_59 ( );
FILL FILL_11_DFFSR_59 ( );
FILL FILL_12_DFFSR_59 ( );
FILL FILL_13_DFFSR_59 ( );
FILL FILL_14_DFFSR_59 ( );
FILL FILL_15_DFFSR_59 ( );
FILL FILL_16_DFFSR_59 ( );
FILL FILL_17_DFFSR_59 ( );
FILL FILL_18_DFFSR_59 ( );
FILL FILL_19_DFFSR_59 ( );
FILL FILL_20_DFFSR_59 ( );
FILL FILL_21_DFFSR_59 ( );
FILL FILL_22_DFFSR_59 ( );
FILL FILL_23_DFFSR_59 ( );
FILL FILL_24_DFFSR_59 ( );
FILL FILL_25_DFFSR_59 ( );
FILL FILL_26_DFFSR_59 ( );
FILL FILL_27_DFFSR_59 ( );
FILL FILL_28_DFFSR_59 ( );
FILL FILL_29_DFFSR_59 ( );
FILL FILL_30_DFFSR_59 ( );
FILL FILL_31_DFFSR_59 ( );
FILL FILL_32_DFFSR_59 ( );
FILL FILL_33_DFFSR_59 ( );
FILL FILL_34_DFFSR_59 ( );
FILL FILL_35_DFFSR_59 ( );
FILL FILL_36_DFFSR_59 ( );
FILL FILL_37_DFFSR_59 ( );
FILL FILL_38_DFFSR_59 ( );
FILL FILL_39_DFFSR_59 ( );
FILL FILL_40_DFFSR_59 ( );
FILL FILL_41_DFFSR_59 ( );
FILL FILL_42_DFFSR_59 ( );
FILL FILL_43_DFFSR_59 ( );
FILL FILL_44_DFFSR_59 ( );
FILL FILL_45_DFFSR_59 ( );
FILL FILL_46_DFFSR_59 ( );
FILL FILL_47_DFFSR_59 ( );
FILL FILL_48_DFFSR_59 ( );
FILL FILL_49_DFFSR_59 ( );
FILL FILL_50_DFFSR_59 ( );
FILL FILL_0_NAND2X1_3 ( );
FILL FILL_1_NAND2X1_3 ( );
FILL FILL_2_NAND2X1_3 ( );
FILL FILL_3_NAND2X1_3 ( );
FILL FILL_4_NAND2X1_3 ( );
FILL FILL_5_NAND2X1_3 ( );
FILL FILL_6_NAND2X1_3 ( );
FILL FILL_0_OAI21X1_3 ( );
FILL FILL_1_OAI21X1_3 ( );
FILL FILL_2_OAI21X1_3 ( );
FILL FILL_3_OAI21X1_3 ( );
FILL FILL_4_OAI21X1_3 ( );
FILL FILL_5_OAI21X1_3 ( );
FILL FILL_6_OAI21X1_3 ( );
FILL FILL_7_OAI21X1_3 ( );
FILL FILL_8_OAI21X1_3 ( );
FILL FILL_0_INVX1_5 ( );
FILL FILL_1_INVX1_5 ( );
FILL FILL_2_INVX1_5 ( );
FILL FILL_3_INVX1_5 ( );
FILL FILL_4_INVX1_5 ( );
FILL FILL_0_OAI21X1_4 ( );
FILL FILL_1_OAI21X1_4 ( );
FILL FILL_2_OAI21X1_4 ( );
FILL FILL_3_OAI21X1_4 ( );
FILL FILL_4_OAI21X1_4 ( );
FILL FILL_5_OAI21X1_4 ( );
FILL FILL_6_OAI21X1_4 ( );
FILL FILL_7_OAI21X1_4 ( );
FILL FILL_8_OAI21X1_4 ( );
FILL FILL_0_DFFSR_166 ( );
FILL FILL_1_DFFSR_166 ( );
FILL FILL_2_DFFSR_166 ( );
FILL FILL_3_DFFSR_166 ( );
FILL FILL_4_DFFSR_166 ( );
FILL FILL_5_DFFSR_166 ( );
FILL FILL_6_DFFSR_166 ( );
FILL FILL_7_DFFSR_166 ( );
FILL FILL_8_DFFSR_166 ( );
FILL FILL_9_DFFSR_166 ( );
FILL FILL_10_DFFSR_166 ( );
FILL FILL_11_DFFSR_166 ( );
FILL FILL_12_DFFSR_166 ( );
FILL FILL_13_DFFSR_166 ( );
FILL FILL_14_DFFSR_166 ( );
FILL FILL_15_DFFSR_166 ( );
FILL FILL_16_DFFSR_166 ( );
FILL FILL_17_DFFSR_166 ( );
FILL FILL_18_DFFSR_166 ( );
FILL FILL_19_DFFSR_166 ( );
FILL FILL_20_DFFSR_166 ( );
FILL FILL_21_DFFSR_166 ( );
FILL FILL_22_DFFSR_166 ( );
FILL FILL_23_DFFSR_166 ( );
FILL FILL_24_DFFSR_166 ( );
FILL FILL_25_DFFSR_166 ( );
FILL FILL_26_DFFSR_166 ( );
FILL FILL_27_DFFSR_166 ( );
FILL FILL_28_DFFSR_166 ( );
FILL FILL_29_DFFSR_166 ( );
FILL FILL_30_DFFSR_166 ( );
FILL FILL_31_DFFSR_166 ( );
FILL FILL_32_DFFSR_166 ( );
FILL FILL_33_DFFSR_166 ( );
FILL FILL_34_DFFSR_166 ( );
FILL FILL_35_DFFSR_166 ( );
FILL FILL_36_DFFSR_166 ( );
FILL FILL_37_DFFSR_166 ( );
FILL FILL_38_DFFSR_166 ( );
FILL FILL_39_DFFSR_166 ( );
FILL FILL_40_DFFSR_166 ( );
FILL FILL_41_DFFSR_166 ( );
FILL FILL_42_DFFSR_166 ( );
FILL FILL_43_DFFSR_166 ( );
FILL FILL_44_DFFSR_166 ( );
FILL FILL_45_DFFSR_166 ( );
FILL FILL_46_DFFSR_166 ( );
FILL FILL_47_DFFSR_166 ( );
FILL FILL_48_DFFSR_166 ( );
FILL FILL_49_DFFSR_166 ( );
FILL FILL_50_DFFSR_166 ( );
FILL FILL_0_BUFX2_30 ( );
FILL FILL_1_BUFX2_30 ( );
FILL FILL_2_BUFX2_30 ( );
FILL FILL_3_BUFX2_30 ( );
FILL FILL_4_BUFX2_30 ( );
FILL FILL_5_BUFX2_30 ( );
FILL FILL_6_BUFX2_30 ( );
FILL FILL_0_INVX1_235 ( );
FILL FILL_1_INVX1_235 ( );
FILL FILL_2_INVX1_235 ( );
FILL FILL_3_INVX1_235 ( );
FILL FILL_0_DFFSR_93 ( );
FILL FILL_1_DFFSR_93 ( );
FILL FILL_2_DFFSR_93 ( );
FILL FILL_3_DFFSR_93 ( );
FILL FILL_4_DFFSR_93 ( );
FILL FILL_5_DFFSR_93 ( );
FILL FILL_6_DFFSR_93 ( );
FILL FILL_7_DFFSR_93 ( );
FILL FILL_8_DFFSR_93 ( );
FILL FILL_9_DFFSR_93 ( );
FILL FILL_10_DFFSR_93 ( );
FILL FILL_11_DFFSR_93 ( );
FILL FILL_12_DFFSR_93 ( );
FILL FILL_13_DFFSR_93 ( );
FILL FILL_14_DFFSR_93 ( );
FILL FILL_15_DFFSR_93 ( );
FILL FILL_16_DFFSR_93 ( );
FILL FILL_17_DFFSR_93 ( );
FILL FILL_18_DFFSR_93 ( );
FILL FILL_19_DFFSR_93 ( );
FILL FILL_20_DFFSR_93 ( );
FILL FILL_21_DFFSR_93 ( );
FILL FILL_22_DFFSR_93 ( );
FILL FILL_23_DFFSR_93 ( );
FILL FILL_24_DFFSR_93 ( );
FILL FILL_25_DFFSR_93 ( );
FILL FILL_26_DFFSR_93 ( );
FILL FILL_27_DFFSR_93 ( );
FILL FILL_28_DFFSR_93 ( );
FILL FILL_29_DFFSR_93 ( );
FILL FILL_30_DFFSR_93 ( );
FILL FILL_31_DFFSR_93 ( );
FILL FILL_32_DFFSR_93 ( );
FILL FILL_33_DFFSR_93 ( );
FILL FILL_34_DFFSR_93 ( );
FILL FILL_35_DFFSR_93 ( );
FILL FILL_36_DFFSR_93 ( );
FILL FILL_37_DFFSR_93 ( );
FILL FILL_38_DFFSR_93 ( );
FILL FILL_39_DFFSR_93 ( );
FILL FILL_40_DFFSR_93 ( );
FILL FILL_41_DFFSR_93 ( );
FILL FILL_42_DFFSR_93 ( );
FILL FILL_43_DFFSR_93 ( );
FILL FILL_44_DFFSR_93 ( );
FILL FILL_45_DFFSR_93 ( );
FILL FILL_46_DFFSR_93 ( );
FILL FILL_47_DFFSR_93 ( );
FILL FILL_48_DFFSR_93 ( );
FILL FILL_49_DFFSR_93 ( );
FILL FILL_50_DFFSR_93 ( );
FILL FILL_51_DFFSR_93 ( );
FILL FILL_0_INVX1_108 ( );
FILL FILL_1_INVX1_108 ( );
FILL FILL_2_INVX1_108 ( );
FILL FILL_3_INVX1_108 ( );
FILL FILL_4_INVX1_108 ( );
FILL FILL_0_DFFSR_66 ( );
FILL FILL_1_DFFSR_66 ( );
FILL FILL_2_DFFSR_66 ( );
FILL FILL_3_DFFSR_66 ( );
FILL FILL_4_DFFSR_66 ( );
FILL FILL_5_DFFSR_66 ( );
FILL FILL_6_DFFSR_66 ( );
FILL FILL_7_DFFSR_66 ( );
FILL FILL_8_DFFSR_66 ( );
FILL FILL_9_DFFSR_66 ( );
FILL FILL_10_DFFSR_66 ( );
FILL FILL_11_DFFSR_66 ( );
FILL FILL_12_DFFSR_66 ( );
FILL FILL_13_DFFSR_66 ( );
FILL FILL_14_DFFSR_66 ( );
FILL FILL_15_DFFSR_66 ( );
FILL FILL_16_DFFSR_66 ( );
FILL FILL_17_DFFSR_66 ( );
FILL FILL_18_DFFSR_66 ( );
FILL FILL_19_DFFSR_66 ( );
FILL FILL_20_DFFSR_66 ( );
FILL FILL_21_DFFSR_66 ( );
FILL FILL_22_DFFSR_66 ( );
FILL FILL_23_DFFSR_66 ( );
FILL FILL_24_DFFSR_66 ( );
FILL FILL_25_DFFSR_66 ( );
FILL FILL_26_DFFSR_66 ( );
FILL FILL_27_DFFSR_66 ( );
FILL FILL_28_DFFSR_66 ( );
FILL FILL_29_DFFSR_66 ( );
FILL FILL_30_DFFSR_66 ( );
FILL FILL_31_DFFSR_66 ( );
FILL FILL_32_DFFSR_66 ( );
FILL FILL_33_DFFSR_66 ( );
FILL FILL_34_DFFSR_66 ( );
FILL FILL_35_DFFSR_66 ( );
FILL FILL_36_DFFSR_66 ( );
FILL FILL_37_DFFSR_66 ( );
FILL FILL_38_DFFSR_66 ( );
FILL FILL_39_DFFSR_66 ( );
FILL FILL_40_DFFSR_66 ( );
FILL FILL_41_DFFSR_66 ( );
FILL FILL_42_DFFSR_66 ( );
FILL FILL_43_DFFSR_66 ( );
FILL FILL_44_DFFSR_66 ( );
FILL FILL_45_DFFSR_66 ( );
FILL FILL_46_DFFSR_66 ( );
FILL FILL_47_DFFSR_66 ( );
FILL FILL_48_DFFSR_66 ( );
FILL FILL_49_DFFSR_66 ( );
FILL FILL_50_DFFSR_66 ( );
FILL FILL_0_DFFSR_67 ( );
FILL FILL_1_DFFSR_67 ( );
FILL FILL_2_DFFSR_67 ( );
FILL FILL_3_DFFSR_67 ( );
FILL FILL_4_DFFSR_67 ( );
FILL FILL_5_DFFSR_67 ( );
FILL FILL_6_DFFSR_67 ( );
FILL FILL_7_DFFSR_67 ( );
FILL FILL_8_DFFSR_67 ( );
FILL FILL_9_DFFSR_67 ( );
FILL FILL_10_DFFSR_67 ( );
FILL FILL_11_DFFSR_67 ( );
FILL FILL_12_DFFSR_67 ( );
FILL FILL_13_DFFSR_67 ( );
FILL FILL_14_DFFSR_67 ( );
FILL FILL_15_DFFSR_67 ( );
FILL FILL_16_DFFSR_67 ( );
FILL FILL_17_DFFSR_67 ( );
FILL FILL_18_DFFSR_67 ( );
FILL FILL_19_DFFSR_67 ( );
FILL FILL_20_DFFSR_67 ( );
FILL FILL_21_DFFSR_67 ( );
FILL FILL_22_DFFSR_67 ( );
FILL FILL_23_DFFSR_67 ( );
FILL FILL_24_DFFSR_67 ( );
FILL FILL_25_DFFSR_67 ( );
FILL FILL_26_DFFSR_67 ( );
FILL FILL_27_DFFSR_67 ( );
FILL FILL_28_DFFSR_67 ( );
FILL FILL_29_DFFSR_67 ( );
FILL FILL_30_DFFSR_67 ( );
FILL FILL_31_DFFSR_67 ( );
FILL FILL_32_DFFSR_67 ( );
FILL FILL_33_DFFSR_67 ( );
FILL FILL_34_DFFSR_67 ( );
FILL FILL_35_DFFSR_67 ( );
FILL FILL_36_DFFSR_67 ( );
FILL FILL_37_DFFSR_67 ( );
FILL FILL_38_DFFSR_67 ( );
FILL FILL_39_DFFSR_67 ( );
FILL FILL_40_DFFSR_67 ( );
FILL FILL_41_DFFSR_67 ( );
FILL FILL_42_DFFSR_67 ( );
FILL FILL_43_DFFSR_67 ( );
FILL FILL_44_DFFSR_67 ( );
FILL FILL_45_DFFSR_67 ( );
FILL FILL_46_DFFSR_67 ( );
FILL FILL_47_DFFSR_67 ( );
FILL FILL_48_DFFSR_67 ( );
FILL FILL_49_DFFSR_67 ( );
FILL FILL_50_DFFSR_67 ( );
FILL FILL_51_DFFSR_67 ( );
FILL FILL_0_DFFSR_132 ( );
FILL FILL_1_DFFSR_132 ( );
FILL FILL_2_DFFSR_132 ( );
FILL FILL_3_DFFSR_132 ( );
FILL FILL_4_DFFSR_132 ( );
FILL FILL_5_DFFSR_132 ( );
FILL FILL_6_DFFSR_132 ( );
FILL FILL_7_DFFSR_132 ( );
FILL FILL_8_DFFSR_132 ( );
FILL FILL_9_DFFSR_132 ( );
FILL FILL_10_DFFSR_132 ( );
FILL FILL_11_DFFSR_132 ( );
FILL FILL_12_DFFSR_132 ( );
FILL FILL_13_DFFSR_132 ( );
FILL FILL_14_DFFSR_132 ( );
FILL FILL_15_DFFSR_132 ( );
FILL FILL_16_DFFSR_132 ( );
FILL FILL_17_DFFSR_132 ( );
FILL FILL_18_DFFSR_132 ( );
FILL FILL_19_DFFSR_132 ( );
FILL FILL_20_DFFSR_132 ( );
FILL FILL_21_DFFSR_132 ( );
FILL FILL_22_DFFSR_132 ( );
FILL FILL_23_DFFSR_132 ( );
FILL FILL_24_DFFSR_132 ( );
FILL FILL_25_DFFSR_132 ( );
FILL FILL_26_DFFSR_132 ( );
FILL FILL_27_DFFSR_132 ( );
FILL FILL_28_DFFSR_132 ( );
FILL FILL_29_DFFSR_132 ( );
FILL FILL_30_DFFSR_132 ( );
FILL FILL_31_DFFSR_132 ( );
FILL FILL_32_DFFSR_132 ( );
FILL FILL_33_DFFSR_132 ( );
FILL FILL_34_DFFSR_132 ( );
FILL FILL_35_DFFSR_132 ( );
FILL FILL_36_DFFSR_132 ( );
FILL FILL_37_DFFSR_132 ( );
FILL FILL_38_DFFSR_132 ( );
FILL FILL_39_DFFSR_132 ( );
FILL FILL_40_DFFSR_132 ( );
FILL FILL_41_DFFSR_132 ( );
FILL FILL_42_DFFSR_132 ( );
FILL FILL_43_DFFSR_132 ( );
FILL FILL_44_DFFSR_132 ( );
FILL FILL_45_DFFSR_132 ( );
FILL FILL_46_DFFSR_132 ( );
FILL FILL_47_DFFSR_132 ( );
FILL FILL_48_DFFSR_132 ( );
FILL FILL_49_DFFSR_132 ( );
FILL FILL_50_DFFSR_132 ( );
FILL FILL_51_DFFSR_132 ( );
FILL FILL_0_INVX1_280 ( );
FILL FILL_1_INVX1_280 ( );
FILL FILL_2_INVX1_280 ( );
FILL FILL_3_INVX1_280 ( );
FILL FILL_4_INVX1_280 ( );
FILL FILL_0_DFFSR_56 ( );
FILL FILL_1_DFFSR_56 ( );
FILL FILL_2_DFFSR_56 ( );
FILL FILL_3_DFFSR_56 ( );
FILL FILL_4_DFFSR_56 ( );
FILL FILL_5_DFFSR_56 ( );
FILL FILL_6_DFFSR_56 ( );
FILL FILL_7_DFFSR_56 ( );
FILL FILL_8_DFFSR_56 ( );
FILL FILL_9_DFFSR_56 ( );
FILL FILL_10_DFFSR_56 ( );
FILL FILL_11_DFFSR_56 ( );
FILL FILL_12_DFFSR_56 ( );
FILL FILL_13_DFFSR_56 ( );
FILL FILL_14_DFFSR_56 ( );
FILL FILL_15_DFFSR_56 ( );
FILL FILL_16_DFFSR_56 ( );
FILL FILL_17_DFFSR_56 ( );
FILL FILL_18_DFFSR_56 ( );
FILL FILL_19_DFFSR_56 ( );
FILL FILL_20_DFFSR_56 ( );
FILL FILL_21_DFFSR_56 ( );
FILL FILL_22_DFFSR_56 ( );
FILL FILL_23_DFFSR_56 ( );
FILL FILL_24_DFFSR_56 ( );
FILL FILL_25_DFFSR_56 ( );
FILL FILL_26_DFFSR_56 ( );
FILL FILL_27_DFFSR_56 ( );
FILL FILL_28_DFFSR_56 ( );
FILL FILL_29_DFFSR_56 ( );
FILL FILL_30_DFFSR_56 ( );
FILL FILL_31_DFFSR_56 ( );
FILL FILL_32_DFFSR_56 ( );
FILL FILL_33_DFFSR_56 ( );
FILL FILL_34_DFFSR_56 ( );
FILL FILL_35_DFFSR_56 ( );
FILL FILL_36_DFFSR_56 ( );
FILL FILL_37_DFFSR_56 ( );
FILL FILL_38_DFFSR_56 ( );
FILL FILL_39_DFFSR_56 ( );
FILL FILL_40_DFFSR_56 ( );
FILL FILL_41_DFFSR_56 ( );
FILL FILL_42_DFFSR_56 ( );
FILL FILL_43_DFFSR_56 ( );
FILL FILL_44_DFFSR_56 ( );
FILL FILL_45_DFFSR_56 ( );
FILL FILL_46_DFFSR_56 ( );
FILL FILL_47_DFFSR_56 ( );
FILL FILL_48_DFFSR_56 ( );
FILL FILL_49_DFFSR_56 ( );
FILL FILL_50_DFFSR_56 ( );
FILL FILL_51_DFFSR_56 ( );
FILL FILL_0_OAI21X1_56 ( );
FILL FILL_1_OAI21X1_56 ( );
FILL FILL_2_OAI21X1_56 ( );
FILL FILL_3_OAI21X1_56 ( );
FILL FILL_4_OAI21X1_56 ( );
FILL FILL_5_OAI21X1_56 ( );
FILL FILL_6_OAI21X1_56 ( );
FILL FILL_7_OAI21X1_56 ( );
FILL FILL_8_OAI21X1_56 ( );
FILL FILL_0_INVX1_63 ( );
FILL FILL_1_INVX1_63 ( );
FILL FILL_2_INVX1_63 ( );
FILL FILL_3_INVX1_63 ( );
FILL FILL_4_INVX1_63 ( );
FILL FILL_0_OAI21X1_51 ( );
FILL FILL_1_OAI21X1_51 ( );
FILL FILL_2_OAI21X1_51 ( );
FILL FILL_3_OAI21X1_51 ( );
FILL FILL_4_OAI21X1_51 ( );
FILL FILL_5_OAI21X1_51 ( );
FILL FILL_6_OAI21X1_51 ( );
FILL FILL_7_OAI21X1_51 ( );
FILL FILL_8_OAI21X1_51 ( );
FILL FILL_0_NAND2X1_51 ( );
FILL FILL_1_NAND2X1_51 ( );
FILL FILL_2_NAND2X1_51 ( );
FILL FILL_3_NAND2X1_51 ( );
FILL FILL_4_NAND2X1_51 ( );
FILL FILL_5_NAND2X1_51 ( );
FILL FILL_6_NAND2X1_51 ( );
FILL FILL_0_DFFSR_51 ( );
FILL FILL_1_DFFSR_51 ( );
FILL FILL_2_DFFSR_51 ( );
FILL FILL_3_DFFSR_51 ( );
FILL FILL_4_DFFSR_51 ( );
FILL FILL_5_DFFSR_51 ( );
FILL FILL_6_DFFSR_51 ( );
FILL FILL_7_DFFSR_51 ( );
FILL FILL_8_DFFSR_51 ( );
FILL FILL_9_DFFSR_51 ( );
FILL FILL_10_DFFSR_51 ( );
FILL FILL_11_DFFSR_51 ( );
FILL FILL_12_DFFSR_51 ( );
FILL FILL_13_DFFSR_51 ( );
FILL FILL_14_DFFSR_51 ( );
FILL FILL_15_DFFSR_51 ( );
FILL FILL_16_DFFSR_51 ( );
FILL FILL_17_DFFSR_51 ( );
FILL FILL_18_DFFSR_51 ( );
FILL FILL_19_DFFSR_51 ( );
FILL FILL_20_DFFSR_51 ( );
FILL FILL_21_DFFSR_51 ( );
FILL FILL_22_DFFSR_51 ( );
FILL FILL_23_DFFSR_51 ( );
FILL FILL_24_DFFSR_51 ( );
FILL FILL_25_DFFSR_51 ( );
FILL FILL_26_DFFSR_51 ( );
FILL FILL_27_DFFSR_51 ( );
FILL FILL_28_DFFSR_51 ( );
FILL FILL_29_DFFSR_51 ( );
FILL FILL_30_DFFSR_51 ( );
FILL FILL_31_DFFSR_51 ( );
FILL FILL_32_DFFSR_51 ( );
FILL FILL_33_DFFSR_51 ( );
FILL FILL_34_DFFSR_51 ( );
FILL FILL_35_DFFSR_51 ( );
FILL FILL_36_DFFSR_51 ( );
FILL FILL_37_DFFSR_51 ( );
FILL FILL_38_DFFSR_51 ( );
FILL FILL_39_DFFSR_51 ( );
FILL FILL_40_DFFSR_51 ( );
FILL FILL_41_DFFSR_51 ( );
FILL FILL_42_DFFSR_51 ( );
FILL FILL_43_DFFSR_51 ( );
FILL FILL_44_DFFSR_51 ( );
FILL FILL_45_DFFSR_51 ( );
FILL FILL_46_DFFSR_51 ( );
FILL FILL_47_DFFSR_51 ( );
FILL FILL_48_DFFSR_51 ( );
FILL FILL_49_DFFSR_51 ( );
FILL FILL_50_DFFSR_51 ( );
FILL FILL_0_INVX1_24 ( );
FILL FILL_1_INVX1_24 ( );
FILL FILL_2_INVX1_24 ( );
FILL FILL_3_INVX1_24 ( );
FILL FILL_4_INVX1_24 ( );
FILL FILL_0_OAI21X1_21 ( );
FILL FILL_1_OAI21X1_21 ( );
FILL FILL_2_OAI21X1_21 ( );
FILL FILL_3_OAI21X1_21 ( );
FILL FILL_4_OAI21X1_21 ( );
FILL FILL_5_OAI21X1_21 ( );
FILL FILL_6_OAI21X1_21 ( );
FILL FILL_7_OAI21X1_21 ( );
FILL FILL_8_OAI21X1_21 ( );
FILL FILL_0_INVX1_409 ( );
FILL FILL_1_INVX1_409 ( );
FILL FILL_2_INVX1_409 ( );
FILL FILL_3_INVX1_409 ( );
FILL FILL_0_INVX1_2 ( );
FILL FILL_1_INVX1_2 ( );
FILL FILL_2_INVX1_2 ( );
FILL FILL_3_INVX1_2 ( );
FILL FILL_4_INVX1_2 ( );
FILL FILL_0_OAI21X1_1 ( );
FILL FILL_1_OAI21X1_1 ( );
FILL FILL_2_OAI21X1_1 ( );
FILL FILL_3_OAI21X1_1 ( );
FILL FILL_4_OAI21X1_1 ( );
FILL FILL_5_OAI21X1_1 ( );
FILL FILL_6_OAI21X1_1 ( );
FILL FILL_7_OAI21X1_1 ( );
FILL FILL_8_OAI21X1_1 ( );
FILL FILL_0_NAND2X1_4 ( );
FILL FILL_1_NAND2X1_4 ( );
FILL FILL_2_NAND2X1_4 ( );
FILL FILL_3_NAND2X1_4 ( );
FILL FILL_4_NAND2X1_4 ( );
FILL FILL_5_NAND2X1_4 ( );
FILL FILL_6_NAND2X1_4 ( );
FILL FILL_0_NAND2X1_263 ( );
FILL FILL_1_NAND2X1_263 ( );
FILL FILL_2_NAND2X1_263 ( );
FILL FILL_3_NAND2X1_263 ( );
FILL FILL_4_NAND2X1_263 ( );
FILL FILL_5_NAND2X1_263 ( );
FILL FILL_6_NAND2X1_263 ( );
FILL FILL_0_NAND2X1_1 ( );
FILL FILL_1_NAND2X1_1 ( );
FILL FILL_2_NAND2X1_1 ( );
FILL FILL_3_NAND2X1_1 ( );
FILL FILL_4_NAND2X1_1 ( );
FILL FILL_5_NAND2X1_1 ( );
FILL FILL_6_NAND2X1_1 ( );
FILL FILL_0_OAI21X1_258 ( );
FILL FILL_1_OAI21X1_258 ( );
FILL FILL_2_OAI21X1_258 ( );
FILL FILL_3_OAI21X1_258 ( );
FILL FILL_4_OAI21X1_258 ( );
FILL FILL_5_OAI21X1_258 ( );
FILL FILL_6_OAI21X1_258 ( );
FILL FILL_7_OAI21X1_258 ( );
FILL FILL_8_OAI21X1_258 ( );
FILL FILL_0_OAI21X1_257 ( );
FILL FILL_1_OAI21X1_257 ( );
FILL FILL_2_OAI21X1_257 ( );
FILL FILL_3_OAI21X1_257 ( );
FILL FILL_4_OAI21X1_257 ( );
FILL FILL_5_OAI21X1_257 ( );
FILL FILL_6_OAI21X1_257 ( );
FILL FILL_7_OAI21X1_257 ( );
FILL FILL_8_OAI21X1_257 ( );
FILL FILL_0_INVX1_420 ( );
FILL FILL_1_INVX1_420 ( );
FILL FILL_2_INVX1_420 ( );
FILL FILL_3_INVX1_420 ( );
FILL FILL_4_INVX1_420 ( );
FILL FILL_0_INVX1_419 ( );
FILL FILL_1_INVX1_419 ( );
FILL FILL_2_INVX1_419 ( );
FILL FILL_3_INVX1_419 ( );
FILL FILL_4_INVX1_419 ( );
FILL FILL_0_OAI21X1_256 ( );
FILL FILL_1_OAI21X1_256 ( );
FILL FILL_2_OAI21X1_256 ( );
FILL FILL_3_OAI21X1_256 ( );
FILL FILL_4_OAI21X1_256 ( );
FILL FILL_5_OAI21X1_256 ( );
FILL FILL_6_OAI21X1_256 ( );
FILL FILL_7_OAI21X1_256 ( );
FILL FILL_8_OAI21X1_256 ( );
FILL FILL_0_DFFSR_96 ( );
FILL FILL_1_DFFSR_96 ( );
FILL FILL_2_DFFSR_96 ( );
FILL FILL_3_DFFSR_96 ( );
FILL FILL_4_DFFSR_96 ( );
FILL FILL_5_DFFSR_96 ( );
FILL FILL_6_DFFSR_96 ( );
FILL FILL_7_DFFSR_96 ( );
FILL FILL_8_DFFSR_96 ( );
FILL FILL_9_DFFSR_96 ( );
FILL FILL_10_DFFSR_96 ( );
FILL FILL_11_DFFSR_96 ( );
FILL FILL_12_DFFSR_96 ( );
FILL FILL_13_DFFSR_96 ( );
FILL FILL_14_DFFSR_96 ( );
FILL FILL_15_DFFSR_96 ( );
FILL FILL_16_DFFSR_96 ( );
FILL FILL_17_DFFSR_96 ( );
FILL FILL_18_DFFSR_96 ( );
FILL FILL_19_DFFSR_96 ( );
FILL FILL_20_DFFSR_96 ( );
FILL FILL_21_DFFSR_96 ( );
FILL FILL_22_DFFSR_96 ( );
FILL FILL_23_DFFSR_96 ( );
FILL FILL_24_DFFSR_96 ( );
FILL FILL_25_DFFSR_96 ( );
FILL FILL_26_DFFSR_96 ( );
FILL FILL_27_DFFSR_96 ( );
FILL FILL_28_DFFSR_96 ( );
FILL FILL_29_DFFSR_96 ( );
FILL FILL_30_DFFSR_96 ( );
FILL FILL_31_DFFSR_96 ( );
FILL FILL_32_DFFSR_96 ( );
FILL FILL_33_DFFSR_96 ( );
FILL FILL_34_DFFSR_96 ( );
FILL FILL_35_DFFSR_96 ( );
FILL FILL_36_DFFSR_96 ( );
FILL FILL_37_DFFSR_96 ( );
FILL FILL_38_DFFSR_96 ( );
FILL FILL_39_DFFSR_96 ( );
FILL FILL_40_DFFSR_96 ( );
FILL FILL_41_DFFSR_96 ( );
FILL FILL_42_DFFSR_96 ( );
FILL FILL_43_DFFSR_96 ( );
FILL FILL_44_DFFSR_96 ( );
FILL FILL_45_DFFSR_96 ( );
FILL FILL_46_DFFSR_96 ( );
FILL FILL_47_DFFSR_96 ( );
FILL FILL_48_DFFSR_96 ( );
FILL FILL_49_DFFSR_96 ( );
FILL FILL_50_DFFSR_96 ( );
FILL FILL_51_DFFSR_96 ( );
FILL FILL_0_INVX1_88 ( );
FILL FILL_1_INVX1_88 ( );
FILL FILL_2_INVX1_88 ( );
FILL FILL_3_INVX1_88 ( );
FILL FILL_4_INVX1_88 ( );
FILL FILL_0_NAND2X1_74 ( );
FILL FILL_1_NAND2X1_74 ( );
FILL FILL_2_NAND2X1_74 ( );
FILL FILL_3_NAND2X1_74 ( );
FILL FILL_4_NAND2X1_74 ( );
FILL FILL_5_NAND2X1_74 ( );
FILL FILL_6_NAND2X1_74 ( );
FILL FILL_0_DFFSR_90 ( );
FILL FILL_1_DFFSR_90 ( );
FILL FILL_2_DFFSR_90 ( );
FILL FILL_3_DFFSR_90 ( );
FILL FILL_4_DFFSR_90 ( );
FILL FILL_5_DFFSR_90 ( );
FILL FILL_6_DFFSR_90 ( );
FILL FILL_7_DFFSR_90 ( );
FILL FILL_8_DFFSR_90 ( );
FILL FILL_9_DFFSR_90 ( );
FILL FILL_10_DFFSR_90 ( );
FILL FILL_11_DFFSR_90 ( );
FILL FILL_12_DFFSR_90 ( );
FILL FILL_13_DFFSR_90 ( );
FILL FILL_14_DFFSR_90 ( );
FILL FILL_15_DFFSR_90 ( );
FILL FILL_16_DFFSR_90 ( );
FILL FILL_17_DFFSR_90 ( );
FILL FILL_18_DFFSR_90 ( );
FILL FILL_19_DFFSR_90 ( );
FILL FILL_20_DFFSR_90 ( );
FILL FILL_21_DFFSR_90 ( );
FILL FILL_22_DFFSR_90 ( );
FILL FILL_23_DFFSR_90 ( );
FILL FILL_24_DFFSR_90 ( );
FILL FILL_25_DFFSR_90 ( );
FILL FILL_26_DFFSR_90 ( );
FILL FILL_27_DFFSR_90 ( );
FILL FILL_28_DFFSR_90 ( );
FILL FILL_29_DFFSR_90 ( );
FILL FILL_30_DFFSR_90 ( );
FILL FILL_31_DFFSR_90 ( );
FILL FILL_32_DFFSR_90 ( );
FILL FILL_33_DFFSR_90 ( );
FILL FILL_34_DFFSR_90 ( );
FILL FILL_35_DFFSR_90 ( );
FILL FILL_36_DFFSR_90 ( );
FILL FILL_37_DFFSR_90 ( );
FILL FILL_38_DFFSR_90 ( );
FILL FILL_39_DFFSR_90 ( );
FILL FILL_40_DFFSR_90 ( );
FILL FILL_41_DFFSR_90 ( );
FILL FILL_42_DFFSR_90 ( );
FILL FILL_43_DFFSR_90 ( );
FILL FILL_44_DFFSR_90 ( );
FILL FILL_45_DFFSR_90 ( );
FILL FILL_46_DFFSR_90 ( );
FILL FILL_47_DFFSR_90 ( );
FILL FILL_48_DFFSR_90 ( );
FILL FILL_49_DFFSR_90 ( );
FILL FILL_50_DFFSR_90 ( );
FILL FILL_0_INVX1_127 ( );
FILL FILL_1_INVX1_127 ( );
FILL FILL_2_INVX1_127 ( );
FILL FILL_3_INVX1_127 ( );
FILL FILL_4_INVX1_127 ( );
FILL FILL_0_INVX1_76 ( );
FILL FILL_1_INVX1_76 ( );
FILL FILL_2_INVX1_76 ( );
FILL FILL_3_INVX1_76 ( );
FILL FILL_4_INVX1_76 ( );
FILL FILL_0_NAND2X1_67 ( );
FILL FILL_1_NAND2X1_67 ( );
FILL FILL_2_NAND2X1_67 ( );
FILL FILL_3_NAND2X1_67 ( );
FILL FILL_4_NAND2X1_67 ( );
FILL FILL_5_NAND2X1_67 ( );
FILL FILL_6_NAND2X1_67 ( );
FILL FILL_0_OAI21X1_67 ( );
FILL FILL_1_OAI21X1_67 ( );
FILL FILL_2_OAI21X1_67 ( );
FILL FILL_3_OAI21X1_67 ( );
FILL FILL_4_OAI21X1_67 ( );
FILL FILL_5_OAI21X1_67 ( );
FILL FILL_6_OAI21X1_67 ( );
FILL FILL_7_OAI21X1_67 ( );
FILL FILL_8_OAI21X1_67 ( );
FILL FILL_0_INVX1_414 ( );
FILL FILL_1_INVX1_414 ( );
FILL FILL_2_INVX1_414 ( );
FILL FILL_3_INVX1_414 ( );
FILL FILL_0_DFFSR_129 ( );
FILL FILL_1_DFFSR_129 ( );
FILL FILL_2_DFFSR_129 ( );
FILL FILL_3_DFFSR_129 ( );
FILL FILL_4_DFFSR_129 ( );
FILL FILL_5_DFFSR_129 ( );
FILL FILL_6_DFFSR_129 ( );
FILL FILL_7_DFFSR_129 ( );
FILL FILL_8_DFFSR_129 ( );
FILL FILL_9_DFFSR_129 ( );
FILL FILL_10_DFFSR_129 ( );
FILL FILL_11_DFFSR_129 ( );
FILL FILL_12_DFFSR_129 ( );
FILL FILL_13_DFFSR_129 ( );
FILL FILL_14_DFFSR_129 ( );
FILL FILL_15_DFFSR_129 ( );
FILL FILL_16_DFFSR_129 ( );
FILL FILL_17_DFFSR_129 ( );
FILL FILL_18_DFFSR_129 ( );
FILL FILL_19_DFFSR_129 ( );
FILL FILL_20_DFFSR_129 ( );
FILL FILL_21_DFFSR_129 ( );
FILL FILL_22_DFFSR_129 ( );
FILL FILL_23_DFFSR_129 ( );
FILL FILL_24_DFFSR_129 ( );
FILL FILL_25_DFFSR_129 ( );
FILL FILL_26_DFFSR_129 ( );
FILL FILL_27_DFFSR_129 ( );
FILL FILL_28_DFFSR_129 ( );
FILL FILL_29_DFFSR_129 ( );
FILL FILL_30_DFFSR_129 ( );
FILL FILL_31_DFFSR_129 ( );
FILL FILL_32_DFFSR_129 ( );
FILL FILL_33_DFFSR_129 ( );
FILL FILL_34_DFFSR_129 ( );
FILL FILL_35_DFFSR_129 ( );
FILL FILL_36_DFFSR_129 ( );
FILL FILL_37_DFFSR_129 ( );
FILL FILL_38_DFFSR_129 ( );
FILL FILL_39_DFFSR_129 ( );
FILL FILL_40_DFFSR_129 ( );
FILL FILL_41_DFFSR_129 ( );
FILL FILL_42_DFFSR_129 ( );
FILL FILL_43_DFFSR_129 ( );
FILL FILL_44_DFFSR_129 ( );
FILL FILL_45_DFFSR_129 ( );
FILL FILL_46_DFFSR_129 ( );
FILL FILL_47_DFFSR_129 ( );
FILL FILL_48_DFFSR_129 ( );
FILL FILL_49_DFFSR_129 ( );
FILL FILL_50_DFFSR_129 ( );
FILL FILL_51_DFFSR_129 ( );
FILL FILL_0_NAND2X1_34 ( );
FILL FILL_1_NAND2X1_34 ( );
FILL FILL_2_NAND2X1_34 ( );
FILL FILL_3_NAND2X1_34 ( );
FILL FILL_4_NAND2X1_34 ( );
FILL FILL_5_NAND2X1_34 ( );
FILL FILL_6_NAND2X1_34 ( );
FILL FILL_0_DFFSR_32 ( );
FILL FILL_1_DFFSR_32 ( );
FILL FILL_2_DFFSR_32 ( );
FILL FILL_3_DFFSR_32 ( );
FILL FILL_4_DFFSR_32 ( );
FILL FILL_5_DFFSR_32 ( );
FILL FILL_6_DFFSR_32 ( );
FILL FILL_7_DFFSR_32 ( );
FILL FILL_8_DFFSR_32 ( );
FILL FILL_9_DFFSR_32 ( );
FILL FILL_10_DFFSR_32 ( );
FILL FILL_11_DFFSR_32 ( );
FILL FILL_12_DFFSR_32 ( );
FILL FILL_13_DFFSR_32 ( );
FILL FILL_14_DFFSR_32 ( );
FILL FILL_15_DFFSR_32 ( );
FILL FILL_16_DFFSR_32 ( );
FILL FILL_17_DFFSR_32 ( );
FILL FILL_18_DFFSR_32 ( );
FILL FILL_19_DFFSR_32 ( );
FILL FILL_20_DFFSR_32 ( );
FILL FILL_21_DFFSR_32 ( );
FILL FILL_22_DFFSR_32 ( );
FILL FILL_23_DFFSR_32 ( );
FILL FILL_24_DFFSR_32 ( );
FILL FILL_25_DFFSR_32 ( );
FILL FILL_26_DFFSR_32 ( );
FILL FILL_27_DFFSR_32 ( );
FILL FILL_28_DFFSR_32 ( );
FILL FILL_29_DFFSR_32 ( );
FILL FILL_30_DFFSR_32 ( );
FILL FILL_31_DFFSR_32 ( );
FILL FILL_32_DFFSR_32 ( );
FILL FILL_33_DFFSR_32 ( );
FILL FILL_34_DFFSR_32 ( );
FILL FILL_35_DFFSR_32 ( );
FILL FILL_36_DFFSR_32 ( );
FILL FILL_37_DFFSR_32 ( );
FILL FILL_38_DFFSR_32 ( );
FILL FILL_39_DFFSR_32 ( );
FILL FILL_40_DFFSR_32 ( );
FILL FILL_41_DFFSR_32 ( );
FILL FILL_42_DFFSR_32 ( );
FILL FILL_43_DFFSR_32 ( );
FILL FILL_44_DFFSR_32 ( );
FILL FILL_45_DFFSR_32 ( );
FILL FILL_46_DFFSR_32 ( );
FILL FILL_47_DFFSR_32 ( );
FILL FILL_48_DFFSR_32 ( );
FILL FILL_49_DFFSR_32 ( );
FILL FILL_50_DFFSR_32 ( );
FILL FILL_51_DFFSR_32 ( );
FILL FILL_0_NAND2X1_236 ( );
FILL FILL_1_NAND2X1_236 ( );
FILL FILL_2_NAND2X1_236 ( );
FILL FILL_3_NAND2X1_236 ( );
FILL FILL_4_NAND2X1_236 ( );
FILL FILL_5_NAND2X1_236 ( );
FILL FILL_0_INVX1_31 ( );
FILL FILL_1_INVX1_31 ( );
FILL FILL_2_INVX1_31 ( );
FILL FILL_3_INVX1_31 ( );
FILL FILL_4_INVX1_31 ( );
FILL FILL_0_INVX1_262 ( );
FILL FILL_1_INVX1_262 ( );
FILL FILL_2_INVX1_262 ( );
FILL FILL_3_INVX1_262 ( );
FILL FILL_4_INVX1_262 ( );
FILL FILL_0_NAND2X1_59 ( );
FILL FILL_1_NAND2X1_59 ( );
FILL FILL_2_NAND2X1_59 ( );
FILL FILL_3_NAND2X1_59 ( );
FILL FILL_4_NAND2X1_59 ( );
FILL FILL_5_NAND2X1_59 ( );
FILL FILL_6_NAND2X1_59 ( );
FILL FILL_0_DFFSR_21 ( );
FILL FILL_1_DFFSR_21 ( );
FILL FILL_2_DFFSR_21 ( );
FILL FILL_3_DFFSR_21 ( );
FILL FILL_4_DFFSR_21 ( );
FILL FILL_5_DFFSR_21 ( );
FILL FILL_6_DFFSR_21 ( );
FILL FILL_7_DFFSR_21 ( );
FILL FILL_8_DFFSR_21 ( );
FILL FILL_9_DFFSR_21 ( );
FILL FILL_10_DFFSR_21 ( );
FILL FILL_11_DFFSR_21 ( );
FILL FILL_12_DFFSR_21 ( );
FILL FILL_13_DFFSR_21 ( );
FILL FILL_14_DFFSR_21 ( );
FILL FILL_15_DFFSR_21 ( );
FILL FILL_16_DFFSR_21 ( );
FILL FILL_17_DFFSR_21 ( );
FILL FILL_18_DFFSR_21 ( );
FILL FILL_19_DFFSR_21 ( );
FILL FILL_20_DFFSR_21 ( );
FILL FILL_21_DFFSR_21 ( );
FILL FILL_22_DFFSR_21 ( );
FILL FILL_23_DFFSR_21 ( );
FILL FILL_24_DFFSR_21 ( );
FILL FILL_25_DFFSR_21 ( );
FILL FILL_26_DFFSR_21 ( );
FILL FILL_27_DFFSR_21 ( );
FILL FILL_28_DFFSR_21 ( );
FILL FILL_29_DFFSR_21 ( );
FILL FILL_30_DFFSR_21 ( );
FILL FILL_31_DFFSR_21 ( );
FILL FILL_32_DFFSR_21 ( );
FILL FILL_33_DFFSR_21 ( );
FILL FILL_34_DFFSR_21 ( );
FILL FILL_35_DFFSR_21 ( );
FILL FILL_36_DFFSR_21 ( );
FILL FILL_37_DFFSR_21 ( );
FILL FILL_38_DFFSR_21 ( );
FILL FILL_39_DFFSR_21 ( );
FILL FILL_40_DFFSR_21 ( );
FILL FILL_41_DFFSR_21 ( );
FILL FILL_42_DFFSR_21 ( );
FILL FILL_43_DFFSR_21 ( );
FILL FILL_44_DFFSR_21 ( );
FILL FILL_45_DFFSR_21 ( );
FILL FILL_46_DFFSR_21 ( );
FILL FILL_47_DFFSR_21 ( );
FILL FILL_48_DFFSR_21 ( );
FILL FILL_49_DFFSR_21 ( );
FILL FILL_50_DFFSR_21 ( );
FILL FILL_0_DFFSR_179 ( );
FILL FILL_1_DFFSR_179 ( );
FILL FILL_2_DFFSR_179 ( );
FILL FILL_3_DFFSR_179 ( );
FILL FILL_4_DFFSR_179 ( );
FILL FILL_5_DFFSR_179 ( );
FILL FILL_6_DFFSR_179 ( );
FILL FILL_7_DFFSR_179 ( );
FILL FILL_8_DFFSR_179 ( );
FILL FILL_9_DFFSR_179 ( );
FILL FILL_10_DFFSR_179 ( );
FILL FILL_11_DFFSR_179 ( );
FILL FILL_12_DFFSR_179 ( );
FILL FILL_13_DFFSR_179 ( );
FILL FILL_14_DFFSR_179 ( );
FILL FILL_15_DFFSR_179 ( );
FILL FILL_16_DFFSR_179 ( );
FILL FILL_17_DFFSR_179 ( );
FILL FILL_18_DFFSR_179 ( );
FILL FILL_19_DFFSR_179 ( );
FILL FILL_20_DFFSR_179 ( );
FILL FILL_21_DFFSR_179 ( );
FILL FILL_22_DFFSR_179 ( );
FILL FILL_23_DFFSR_179 ( );
FILL FILL_24_DFFSR_179 ( );
FILL FILL_25_DFFSR_179 ( );
FILL FILL_26_DFFSR_179 ( );
FILL FILL_27_DFFSR_179 ( );
FILL FILL_28_DFFSR_179 ( );
FILL FILL_29_DFFSR_179 ( );
FILL FILL_30_DFFSR_179 ( );
FILL FILL_31_DFFSR_179 ( );
FILL FILL_32_DFFSR_179 ( );
FILL FILL_33_DFFSR_179 ( );
FILL FILL_34_DFFSR_179 ( );
FILL FILL_35_DFFSR_179 ( );
FILL FILL_36_DFFSR_179 ( );
FILL FILL_37_DFFSR_179 ( );
FILL FILL_38_DFFSR_179 ( );
FILL FILL_39_DFFSR_179 ( );
FILL FILL_40_DFFSR_179 ( );
FILL FILL_41_DFFSR_179 ( );
FILL FILL_42_DFFSR_179 ( );
FILL FILL_43_DFFSR_179 ( );
FILL FILL_44_DFFSR_179 ( );
FILL FILL_45_DFFSR_179 ( );
FILL FILL_46_DFFSR_179 ( );
FILL FILL_47_DFFSR_179 ( );
FILL FILL_48_DFFSR_179 ( );
FILL FILL_49_DFFSR_179 ( );
FILL FILL_50_DFFSR_179 ( );
FILL FILL_51_DFFSR_179 ( );
FILL FILL_0_DFFSR_188 ( );
FILL FILL_1_DFFSR_188 ( );
FILL FILL_2_DFFSR_188 ( );
FILL FILL_3_DFFSR_188 ( );
FILL FILL_4_DFFSR_188 ( );
FILL FILL_5_DFFSR_188 ( );
FILL FILL_6_DFFSR_188 ( );
FILL FILL_7_DFFSR_188 ( );
FILL FILL_8_DFFSR_188 ( );
FILL FILL_9_DFFSR_188 ( );
FILL FILL_10_DFFSR_188 ( );
FILL FILL_11_DFFSR_188 ( );
FILL FILL_12_DFFSR_188 ( );
FILL FILL_13_DFFSR_188 ( );
FILL FILL_14_DFFSR_188 ( );
FILL FILL_15_DFFSR_188 ( );
FILL FILL_16_DFFSR_188 ( );
FILL FILL_17_DFFSR_188 ( );
FILL FILL_18_DFFSR_188 ( );
FILL FILL_19_DFFSR_188 ( );
FILL FILL_20_DFFSR_188 ( );
FILL FILL_21_DFFSR_188 ( );
FILL FILL_22_DFFSR_188 ( );
FILL FILL_23_DFFSR_188 ( );
FILL FILL_24_DFFSR_188 ( );
FILL FILL_25_DFFSR_188 ( );
FILL FILL_26_DFFSR_188 ( );
FILL FILL_27_DFFSR_188 ( );
FILL FILL_28_DFFSR_188 ( );
FILL FILL_29_DFFSR_188 ( );
FILL FILL_30_DFFSR_188 ( );
FILL FILL_31_DFFSR_188 ( );
FILL FILL_32_DFFSR_188 ( );
FILL FILL_33_DFFSR_188 ( );
FILL FILL_34_DFFSR_188 ( );
FILL FILL_35_DFFSR_188 ( );
FILL FILL_36_DFFSR_188 ( );
FILL FILL_37_DFFSR_188 ( );
FILL FILL_38_DFFSR_188 ( );
FILL FILL_39_DFFSR_188 ( );
FILL FILL_40_DFFSR_188 ( );
FILL FILL_41_DFFSR_188 ( );
FILL FILL_42_DFFSR_188 ( );
FILL FILL_43_DFFSR_188 ( );
FILL FILL_44_DFFSR_188 ( );
FILL FILL_45_DFFSR_188 ( );
FILL FILL_46_DFFSR_188 ( );
FILL FILL_47_DFFSR_188 ( );
FILL FILL_48_DFFSR_188 ( );
FILL FILL_49_DFFSR_188 ( );
FILL FILL_50_DFFSR_188 ( );
FILL FILL_0_NAND3X1_34 ( );
FILL FILL_1_NAND3X1_34 ( );
FILL FILL_2_NAND3X1_34 ( );
FILL FILL_3_NAND3X1_34 ( );
FILL FILL_4_NAND3X1_34 ( );
FILL FILL_5_NAND3X1_34 ( );
FILL FILL_6_NAND3X1_34 ( );
FILL FILL_7_NAND3X1_34 ( );
FILL FILL_8_NAND3X1_34 ( );
FILL FILL_0_DFFSR_78 ( );
FILL FILL_1_DFFSR_78 ( );
FILL FILL_2_DFFSR_78 ( );
FILL FILL_3_DFFSR_78 ( );
FILL FILL_4_DFFSR_78 ( );
FILL FILL_5_DFFSR_78 ( );
FILL FILL_6_DFFSR_78 ( );
FILL FILL_7_DFFSR_78 ( );
FILL FILL_8_DFFSR_78 ( );
FILL FILL_9_DFFSR_78 ( );
FILL FILL_10_DFFSR_78 ( );
FILL FILL_11_DFFSR_78 ( );
FILL FILL_12_DFFSR_78 ( );
FILL FILL_13_DFFSR_78 ( );
FILL FILL_14_DFFSR_78 ( );
FILL FILL_15_DFFSR_78 ( );
FILL FILL_16_DFFSR_78 ( );
FILL FILL_17_DFFSR_78 ( );
FILL FILL_18_DFFSR_78 ( );
FILL FILL_19_DFFSR_78 ( );
FILL FILL_20_DFFSR_78 ( );
FILL FILL_21_DFFSR_78 ( );
FILL FILL_22_DFFSR_78 ( );
FILL FILL_23_DFFSR_78 ( );
FILL FILL_24_DFFSR_78 ( );
FILL FILL_25_DFFSR_78 ( );
FILL FILL_26_DFFSR_78 ( );
FILL FILL_27_DFFSR_78 ( );
FILL FILL_28_DFFSR_78 ( );
FILL FILL_29_DFFSR_78 ( );
FILL FILL_30_DFFSR_78 ( );
FILL FILL_31_DFFSR_78 ( );
FILL FILL_32_DFFSR_78 ( );
FILL FILL_33_DFFSR_78 ( );
FILL FILL_34_DFFSR_78 ( );
FILL FILL_35_DFFSR_78 ( );
FILL FILL_36_DFFSR_78 ( );
FILL FILL_37_DFFSR_78 ( );
FILL FILL_38_DFFSR_78 ( );
FILL FILL_39_DFFSR_78 ( );
FILL FILL_40_DFFSR_78 ( );
FILL FILL_41_DFFSR_78 ( );
FILL FILL_42_DFFSR_78 ( );
FILL FILL_43_DFFSR_78 ( );
FILL FILL_44_DFFSR_78 ( );
FILL FILL_45_DFFSR_78 ( );
FILL FILL_46_DFFSR_78 ( );
FILL FILL_47_DFFSR_78 ( );
FILL FILL_48_DFFSR_78 ( );
FILL FILL_49_DFFSR_78 ( );
FILL FILL_50_DFFSR_78 ( );
FILL FILL_0_OAI21X1_78 ( );
FILL FILL_1_OAI21X1_78 ( );
FILL FILL_2_OAI21X1_78 ( );
FILL FILL_3_OAI21X1_78 ( );
FILL FILL_4_OAI21X1_78 ( );
FILL FILL_5_OAI21X1_78 ( );
FILL FILL_6_OAI21X1_78 ( );
FILL FILL_7_OAI21X1_78 ( );
FILL FILL_8_OAI21X1_78 ( );
FILL FILL_0_NAND2X1_90 ( );
FILL FILL_1_NAND2X1_90 ( );
FILL FILL_2_NAND2X1_90 ( );
FILL FILL_3_NAND2X1_90 ( );
FILL FILL_4_NAND2X1_90 ( );
FILL FILL_5_NAND2X1_90 ( );
FILL FILL_6_NAND2X1_90 ( );
FILL FILL_0_OAI21X1_90 ( );
FILL FILL_1_OAI21X1_90 ( );
FILL FILL_2_OAI21X1_90 ( );
FILL FILL_3_OAI21X1_90 ( );
FILL FILL_4_OAI21X1_90 ( );
FILL FILL_5_OAI21X1_90 ( );
FILL FILL_6_OAI21X1_90 ( );
FILL FILL_7_OAI21X1_90 ( );
FILL FILL_8_OAI21X1_90 ( );
FILL FILL_0_INVX1_343 ( );
FILL FILL_1_INVX1_343 ( );
FILL FILL_2_INVX1_343 ( );
FILL FILL_3_INVX1_343 ( );
FILL FILL_0_INVX1_102 ( );
FILL FILL_1_INVX1_102 ( );
FILL FILL_2_INVX1_102 ( );
FILL FILL_3_INVX1_102 ( );
FILL FILL_4_INVX1_102 ( );
FILL FILL_0_INVX1_346 ( );
FILL FILL_1_INVX1_346 ( );
FILL FILL_2_INVX1_346 ( );
FILL FILL_3_INVX1_346 ( );
FILL FILL_4_INVX1_346 ( );
FILL FILL_0_INVX1_120 ( );
FILL FILL_1_INVX1_120 ( );
FILL FILL_2_INVX1_120 ( );
FILL FILL_3_INVX1_120 ( );
FILL FILL_4_INVX1_120 ( );
FILL FILL_0_DFFSR_106 ( );
FILL FILL_1_DFFSR_106 ( );
FILL FILL_2_DFFSR_106 ( );
FILL FILL_3_DFFSR_106 ( );
FILL FILL_4_DFFSR_106 ( );
FILL FILL_5_DFFSR_106 ( );
FILL FILL_6_DFFSR_106 ( );
FILL FILL_7_DFFSR_106 ( );
FILL FILL_8_DFFSR_106 ( );
FILL FILL_9_DFFSR_106 ( );
FILL FILL_10_DFFSR_106 ( );
FILL FILL_11_DFFSR_106 ( );
FILL FILL_12_DFFSR_106 ( );
FILL FILL_13_DFFSR_106 ( );
FILL FILL_14_DFFSR_106 ( );
FILL FILL_15_DFFSR_106 ( );
FILL FILL_16_DFFSR_106 ( );
FILL FILL_17_DFFSR_106 ( );
FILL FILL_18_DFFSR_106 ( );
FILL FILL_19_DFFSR_106 ( );
FILL FILL_20_DFFSR_106 ( );
FILL FILL_21_DFFSR_106 ( );
FILL FILL_22_DFFSR_106 ( );
FILL FILL_23_DFFSR_106 ( );
FILL FILL_24_DFFSR_106 ( );
FILL FILL_25_DFFSR_106 ( );
FILL FILL_26_DFFSR_106 ( );
FILL FILL_27_DFFSR_106 ( );
FILL FILL_28_DFFSR_106 ( );
FILL FILL_29_DFFSR_106 ( );
FILL FILL_30_DFFSR_106 ( );
FILL FILL_31_DFFSR_106 ( );
FILL FILL_32_DFFSR_106 ( );
FILL FILL_33_DFFSR_106 ( );
FILL FILL_34_DFFSR_106 ( );
FILL FILL_35_DFFSR_106 ( );
FILL FILL_36_DFFSR_106 ( );
FILL FILL_37_DFFSR_106 ( );
FILL FILL_38_DFFSR_106 ( );
FILL FILL_39_DFFSR_106 ( );
FILL FILL_40_DFFSR_106 ( );
FILL FILL_41_DFFSR_106 ( );
FILL FILL_42_DFFSR_106 ( );
FILL FILL_43_DFFSR_106 ( );
FILL FILL_44_DFFSR_106 ( );
FILL FILL_45_DFFSR_106 ( );
FILL FILL_46_DFFSR_106 ( );
FILL FILL_47_DFFSR_106 ( );
FILL FILL_48_DFFSR_106 ( );
FILL FILL_49_DFFSR_106 ( );
FILL FILL_50_DFFSR_106 ( );
FILL FILL_0_DFFSR_131 ( );
FILL FILL_1_DFFSR_131 ( );
FILL FILL_2_DFFSR_131 ( );
FILL FILL_3_DFFSR_131 ( );
FILL FILL_4_DFFSR_131 ( );
FILL FILL_5_DFFSR_131 ( );
FILL FILL_6_DFFSR_131 ( );
FILL FILL_7_DFFSR_131 ( );
FILL FILL_8_DFFSR_131 ( );
FILL FILL_9_DFFSR_131 ( );
FILL FILL_10_DFFSR_131 ( );
FILL FILL_11_DFFSR_131 ( );
FILL FILL_12_DFFSR_131 ( );
FILL FILL_13_DFFSR_131 ( );
FILL FILL_14_DFFSR_131 ( );
FILL FILL_15_DFFSR_131 ( );
FILL FILL_16_DFFSR_131 ( );
FILL FILL_17_DFFSR_131 ( );
FILL FILL_18_DFFSR_131 ( );
FILL FILL_19_DFFSR_131 ( );
FILL FILL_20_DFFSR_131 ( );
FILL FILL_21_DFFSR_131 ( );
FILL FILL_22_DFFSR_131 ( );
FILL FILL_23_DFFSR_131 ( );
FILL FILL_24_DFFSR_131 ( );
FILL FILL_25_DFFSR_131 ( );
FILL FILL_26_DFFSR_131 ( );
FILL FILL_27_DFFSR_131 ( );
FILL FILL_28_DFFSR_131 ( );
FILL FILL_29_DFFSR_131 ( );
FILL FILL_30_DFFSR_131 ( );
FILL FILL_31_DFFSR_131 ( );
FILL FILL_32_DFFSR_131 ( );
FILL FILL_33_DFFSR_131 ( );
FILL FILL_34_DFFSR_131 ( );
FILL FILL_35_DFFSR_131 ( );
FILL FILL_36_DFFSR_131 ( );
FILL FILL_37_DFFSR_131 ( );
FILL FILL_38_DFFSR_131 ( );
FILL FILL_39_DFFSR_131 ( );
FILL FILL_40_DFFSR_131 ( );
FILL FILL_41_DFFSR_131 ( );
FILL FILL_42_DFFSR_131 ( );
FILL FILL_43_DFFSR_131 ( );
FILL FILL_44_DFFSR_131 ( );
FILL FILL_45_DFFSR_131 ( );
FILL FILL_46_DFFSR_131 ( );
FILL FILL_47_DFFSR_131 ( );
FILL FILL_48_DFFSR_131 ( );
FILL FILL_49_DFFSR_131 ( );
FILL FILL_50_DFFSR_131 ( );
FILL FILL_0_OAI21X1_34 ( );
FILL FILL_1_OAI21X1_34 ( );
FILL FILL_2_OAI21X1_34 ( );
FILL FILL_3_OAI21X1_34 ( );
FILL FILL_4_OAI21X1_34 ( );
FILL FILL_5_OAI21X1_34 ( );
FILL FILL_6_OAI21X1_34 ( );
FILL FILL_7_OAI21X1_34 ( );
FILL FILL_8_OAI21X1_34 ( );
FILL FILL_9_OAI21X1_34 ( );
FILL FILL_0_INVX1_39 ( );
FILL FILL_1_INVX1_39 ( );
FILL FILL_2_INVX1_39 ( );
FILL FILL_3_INVX1_39 ( );
FILL FILL_0_INVX1_276 ( );
FILL FILL_1_INVX1_276 ( );
FILL FILL_2_INVX1_276 ( );
FILL FILL_3_INVX1_276 ( );
FILL FILL_4_INVX1_276 ( );
FILL FILL_0_DFFSR_27 ( );
FILL FILL_1_DFFSR_27 ( );
FILL FILL_2_DFFSR_27 ( );
FILL FILL_3_DFFSR_27 ( );
FILL FILL_4_DFFSR_27 ( );
FILL FILL_5_DFFSR_27 ( );
FILL FILL_6_DFFSR_27 ( );
FILL FILL_7_DFFSR_27 ( );
FILL FILL_8_DFFSR_27 ( );
FILL FILL_9_DFFSR_27 ( );
FILL FILL_10_DFFSR_27 ( );
FILL FILL_11_DFFSR_27 ( );
FILL FILL_12_DFFSR_27 ( );
FILL FILL_13_DFFSR_27 ( );
FILL FILL_14_DFFSR_27 ( );
FILL FILL_15_DFFSR_27 ( );
FILL FILL_16_DFFSR_27 ( );
FILL FILL_17_DFFSR_27 ( );
FILL FILL_18_DFFSR_27 ( );
FILL FILL_19_DFFSR_27 ( );
FILL FILL_20_DFFSR_27 ( );
FILL FILL_21_DFFSR_27 ( );
FILL FILL_22_DFFSR_27 ( );
FILL FILL_23_DFFSR_27 ( );
FILL FILL_24_DFFSR_27 ( );
FILL FILL_25_DFFSR_27 ( );
FILL FILL_26_DFFSR_27 ( );
FILL FILL_27_DFFSR_27 ( );
FILL FILL_28_DFFSR_27 ( );
FILL FILL_29_DFFSR_27 ( );
FILL FILL_30_DFFSR_27 ( );
FILL FILL_31_DFFSR_27 ( );
FILL FILL_32_DFFSR_27 ( );
FILL FILL_33_DFFSR_27 ( );
FILL FILL_34_DFFSR_27 ( );
FILL FILL_35_DFFSR_27 ( );
FILL FILL_36_DFFSR_27 ( );
FILL FILL_37_DFFSR_27 ( );
FILL FILL_38_DFFSR_27 ( );
FILL FILL_39_DFFSR_27 ( );
FILL FILL_40_DFFSR_27 ( );
FILL FILL_41_DFFSR_27 ( );
FILL FILL_42_DFFSR_27 ( );
FILL FILL_43_DFFSR_27 ( );
FILL FILL_44_DFFSR_27 ( );
FILL FILL_45_DFFSR_27 ( );
FILL FILL_46_DFFSR_27 ( );
FILL FILL_47_DFFSR_27 ( );
FILL FILL_48_DFFSR_27 ( );
FILL FILL_49_DFFSR_27 ( );
FILL FILL_50_DFFSR_27 ( );
FILL FILL_0_OAI21X1_27 ( );
FILL FILL_1_OAI21X1_27 ( );
FILL FILL_2_OAI21X1_27 ( );
FILL FILL_3_OAI21X1_27 ( );
FILL FILL_4_OAI21X1_27 ( );
FILL FILL_5_OAI21X1_27 ( );
FILL FILL_6_OAI21X1_27 ( );
FILL FILL_7_OAI21X1_27 ( );
FILL FILL_8_OAI21X1_27 ( );
FILL FILL_0_INVX1_284 ( );
FILL FILL_1_INVX1_284 ( );
FILL FILL_2_INVX1_284 ( );
FILL FILL_3_INVX1_284 ( );
FILL FILL_4_INVX1_284 ( );
FILL FILL_0_NAND2X1_27 ( );
FILL FILL_1_NAND2X1_27 ( );
FILL FILL_2_NAND2X1_27 ( );
FILL FILL_3_NAND2X1_27 ( );
FILL FILL_4_NAND2X1_27 ( );
FILL FILL_5_NAND2X1_27 ( );
FILL FILL_6_NAND2X1_27 ( );
FILL FILL_0_INVX1_22 ( );
FILL FILL_1_INVX1_22 ( );
FILL FILL_2_INVX1_22 ( );
FILL FILL_3_INVX1_22 ( );
FILL FILL_4_INVX1_22 ( );
FILL FILL_0_OAI21X1_19 ( );
FILL FILL_1_OAI21X1_19 ( );
FILL FILL_2_OAI21X1_19 ( );
FILL FILL_3_OAI21X1_19 ( );
FILL FILL_4_OAI21X1_19 ( );
FILL FILL_5_OAI21X1_19 ( );
FILL FILL_6_OAI21X1_19 ( );
FILL FILL_7_OAI21X1_19 ( );
FILL FILL_8_OAI21X1_19 ( );
FILL FILL_0_NAND2X1_19 ( );
FILL FILL_1_NAND2X1_19 ( );
FILL FILL_2_NAND2X1_19 ( );
FILL FILL_3_NAND2X1_19 ( );
FILL FILL_4_NAND2X1_19 ( );
FILL FILL_5_NAND2X1_19 ( );
FILL FILL_6_NAND2X1_19 ( );
FILL FILL_0_INVX1_11 ( );
FILL FILL_1_INVX1_11 ( );
FILL FILL_2_INVX1_11 ( );
FILL FILL_3_INVX1_11 ( );
FILL FILL_0_NAND2X1_9 ( );
FILL FILL_1_NAND2X1_9 ( );
FILL FILL_2_NAND2X1_9 ( );
FILL FILL_3_NAND2X1_9 ( );
FILL FILL_4_NAND2X1_9 ( );
FILL FILL_5_NAND2X1_9 ( );
FILL FILL_6_NAND2X1_9 ( );
FILL FILL_0_DFFSR_1 ( );
FILL FILL_1_DFFSR_1 ( );
FILL FILL_2_DFFSR_1 ( );
FILL FILL_3_DFFSR_1 ( );
FILL FILL_4_DFFSR_1 ( );
FILL FILL_5_DFFSR_1 ( );
FILL FILL_6_DFFSR_1 ( );
FILL FILL_7_DFFSR_1 ( );
FILL FILL_8_DFFSR_1 ( );
FILL FILL_9_DFFSR_1 ( );
FILL FILL_10_DFFSR_1 ( );
FILL FILL_11_DFFSR_1 ( );
FILL FILL_12_DFFSR_1 ( );
FILL FILL_13_DFFSR_1 ( );
FILL FILL_14_DFFSR_1 ( );
FILL FILL_15_DFFSR_1 ( );
FILL FILL_16_DFFSR_1 ( );
FILL FILL_17_DFFSR_1 ( );
FILL FILL_18_DFFSR_1 ( );
FILL FILL_19_DFFSR_1 ( );
FILL FILL_20_DFFSR_1 ( );
FILL FILL_21_DFFSR_1 ( );
FILL FILL_22_DFFSR_1 ( );
FILL FILL_23_DFFSR_1 ( );
FILL FILL_24_DFFSR_1 ( );
FILL FILL_25_DFFSR_1 ( );
FILL FILL_26_DFFSR_1 ( );
FILL FILL_27_DFFSR_1 ( );
FILL FILL_28_DFFSR_1 ( );
FILL FILL_29_DFFSR_1 ( );
FILL FILL_30_DFFSR_1 ( );
FILL FILL_31_DFFSR_1 ( );
FILL FILL_32_DFFSR_1 ( );
FILL FILL_33_DFFSR_1 ( );
FILL FILL_34_DFFSR_1 ( );
FILL FILL_35_DFFSR_1 ( );
FILL FILL_36_DFFSR_1 ( );
FILL FILL_37_DFFSR_1 ( );
FILL FILL_38_DFFSR_1 ( );
FILL FILL_39_DFFSR_1 ( );
FILL FILL_40_DFFSR_1 ( );
FILL FILL_41_DFFSR_1 ( );
FILL FILL_42_DFFSR_1 ( );
FILL FILL_43_DFFSR_1 ( );
FILL FILL_44_DFFSR_1 ( );
FILL FILL_45_DFFSR_1 ( );
FILL FILL_46_DFFSR_1 ( );
FILL FILL_47_DFFSR_1 ( );
FILL FILL_48_DFFSR_1 ( );
FILL FILL_49_DFFSR_1 ( );
FILL FILL_50_DFFSR_1 ( );
FILL FILL_51_DFFSR_1 ( );
FILL FILL_0_OAI21X1_247 ( );
FILL FILL_1_OAI21X1_247 ( );
FILL FILL_2_OAI21X1_247 ( );
FILL FILL_3_OAI21X1_247 ( );
FILL FILL_4_OAI21X1_247 ( );
FILL FILL_5_OAI21X1_247 ( );
FILL FILL_6_OAI21X1_247 ( );
FILL FILL_7_OAI21X1_247 ( );
FILL FILL_8_OAI21X1_247 ( );
FILL FILL_9_OAI21X1_247 ( );
FILL FILL_0_OAI21X1_252 ( );
FILL FILL_1_OAI21X1_252 ( );
FILL FILL_2_OAI21X1_252 ( );
FILL FILL_3_OAI21X1_252 ( );
FILL FILL_4_OAI21X1_252 ( );
FILL FILL_5_OAI21X1_252 ( );
FILL FILL_6_OAI21X1_252 ( );
FILL FILL_7_OAI21X1_252 ( );
FILL FILL_8_OAI21X1_252 ( );
FILL FILL_0_DFFSR_189 ( );
FILL FILL_1_DFFSR_189 ( );
FILL FILL_2_DFFSR_189 ( );
FILL FILL_3_DFFSR_189 ( );
FILL FILL_4_DFFSR_189 ( );
FILL FILL_5_DFFSR_189 ( );
FILL FILL_6_DFFSR_189 ( );
FILL FILL_7_DFFSR_189 ( );
FILL FILL_8_DFFSR_189 ( );
FILL FILL_9_DFFSR_189 ( );
FILL FILL_10_DFFSR_189 ( );
FILL FILL_11_DFFSR_189 ( );
FILL FILL_12_DFFSR_189 ( );
FILL FILL_13_DFFSR_189 ( );
FILL FILL_14_DFFSR_189 ( );
FILL FILL_15_DFFSR_189 ( );
FILL FILL_16_DFFSR_189 ( );
FILL FILL_17_DFFSR_189 ( );
FILL FILL_18_DFFSR_189 ( );
FILL FILL_19_DFFSR_189 ( );
FILL FILL_20_DFFSR_189 ( );
FILL FILL_21_DFFSR_189 ( );
FILL FILL_22_DFFSR_189 ( );
FILL FILL_23_DFFSR_189 ( );
FILL FILL_24_DFFSR_189 ( );
FILL FILL_25_DFFSR_189 ( );
FILL FILL_26_DFFSR_189 ( );
FILL FILL_27_DFFSR_189 ( );
FILL FILL_28_DFFSR_189 ( );
FILL FILL_29_DFFSR_189 ( );
FILL FILL_30_DFFSR_189 ( );
FILL FILL_31_DFFSR_189 ( );
FILL FILL_32_DFFSR_189 ( );
FILL FILL_33_DFFSR_189 ( );
FILL FILL_34_DFFSR_189 ( );
FILL FILL_35_DFFSR_189 ( );
FILL FILL_36_DFFSR_189 ( );
FILL FILL_37_DFFSR_189 ( );
FILL FILL_38_DFFSR_189 ( );
FILL FILL_39_DFFSR_189 ( );
FILL FILL_40_DFFSR_189 ( );
FILL FILL_41_DFFSR_189 ( );
FILL FILL_42_DFFSR_189 ( );
FILL FILL_43_DFFSR_189 ( );
FILL FILL_44_DFFSR_189 ( );
FILL FILL_45_DFFSR_189 ( );
FILL FILL_46_DFFSR_189 ( );
FILL FILL_47_DFFSR_189 ( );
FILL FILL_48_DFFSR_189 ( );
FILL FILL_49_DFFSR_189 ( );
FILL FILL_50_DFFSR_189 ( );
FILL FILL_51_DFFSR_189 ( );
FILL FILL_0_DFFSR_86 ( );
FILL FILL_1_DFFSR_86 ( );
FILL FILL_2_DFFSR_86 ( );
FILL FILL_3_DFFSR_86 ( );
FILL FILL_4_DFFSR_86 ( );
FILL FILL_5_DFFSR_86 ( );
FILL FILL_6_DFFSR_86 ( );
FILL FILL_7_DFFSR_86 ( );
FILL FILL_8_DFFSR_86 ( );
FILL FILL_9_DFFSR_86 ( );
FILL FILL_10_DFFSR_86 ( );
FILL FILL_11_DFFSR_86 ( );
FILL FILL_12_DFFSR_86 ( );
FILL FILL_13_DFFSR_86 ( );
FILL FILL_14_DFFSR_86 ( );
FILL FILL_15_DFFSR_86 ( );
FILL FILL_16_DFFSR_86 ( );
FILL FILL_17_DFFSR_86 ( );
FILL FILL_18_DFFSR_86 ( );
FILL FILL_19_DFFSR_86 ( );
FILL FILL_20_DFFSR_86 ( );
FILL FILL_21_DFFSR_86 ( );
FILL FILL_22_DFFSR_86 ( );
FILL FILL_23_DFFSR_86 ( );
FILL FILL_24_DFFSR_86 ( );
FILL FILL_25_DFFSR_86 ( );
FILL FILL_26_DFFSR_86 ( );
FILL FILL_27_DFFSR_86 ( );
FILL FILL_28_DFFSR_86 ( );
FILL FILL_29_DFFSR_86 ( );
FILL FILL_30_DFFSR_86 ( );
FILL FILL_31_DFFSR_86 ( );
FILL FILL_32_DFFSR_86 ( );
FILL FILL_33_DFFSR_86 ( );
FILL FILL_34_DFFSR_86 ( );
FILL FILL_35_DFFSR_86 ( );
FILL FILL_36_DFFSR_86 ( );
FILL FILL_37_DFFSR_86 ( );
FILL FILL_38_DFFSR_86 ( );
FILL FILL_39_DFFSR_86 ( );
FILL FILL_40_DFFSR_86 ( );
FILL FILL_41_DFFSR_86 ( );
FILL FILL_42_DFFSR_86 ( );
FILL FILL_43_DFFSR_86 ( );
FILL FILL_44_DFFSR_86 ( );
FILL FILL_45_DFFSR_86 ( );
FILL FILL_46_DFFSR_86 ( );
FILL FILL_47_DFFSR_86 ( );
FILL FILL_48_DFFSR_86 ( );
FILL FILL_49_DFFSR_86 ( );
FILL FILL_50_DFFSR_86 ( );
FILL FILL_0_DFFSR_82 ( );
FILL FILL_1_DFFSR_82 ( );
FILL FILL_2_DFFSR_82 ( );
FILL FILL_3_DFFSR_82 ( );
FILL FILL_4_DFFSR_82 ( );
FILL FILL_5_DFFSR_82 ( );
FILL FILL_6_DFFSR_82 ( );
FILL FILL_7_DFFSR_82 ( );
FILL FILL_8_DFFSR_82 ( );
FILL FILL_9_DFFSR_82 ( );
FILL FILL_10_DFFSR_82 ( );
FILL FILL_11_DFFSR_82 ( );
FILL FILL_12_DFFSR_82 ( );
FILL FILL_13_DFFSR_82 ( );
FILL FILL_14_DFFSR_82 ( );
FILL FILL_15_DFFSR_82 ( );
FILL FILL_16_DFFSR_82 ( );
FILL FILL_17_DFFSR_82 ( );
FILL FILL_18_DFFSR_82 ( );
FILL FILL_19_DFFSR_82 ( );
FILL FILL_20_DFFSR_82 ( );
FILL FILL_21_DFFSR_82 ( );
FILL FILL_22_DFFSR_82 ( );
FILL FILL_23_DFFSR_82 ( );
FILL FILL_24_DFFSR_82 ( );
FILL FILL_25_DFFSR_82 ( );
FILL FILL_26_DFFSR_82 ( );
FILL FILL_27_DFFSR_82 ( );
FILL FILL_28_DFFSR_82 ( );
FILL FILL_29_DFFSR_82 ( );
FILL FILL_30_DFFSR_82 ( );
FILL FILL_31_DFFSR_82 ( );
FILL FILL_32_DFFSR_82 ( );
FILL FILL_33_DFFSR_82 ( );
FILL FILL_34_DFFSR_82 ( );
FILL FILL_35_DFFSR_82 ( );
FILL FILL_36_DFFSR_82 ( );
FILL FILL_37_DFFSR_82 ( );
FILL FILL_38_DFFSR_82 ( );
FILL FILL_39_DFFSR_82 ( );
FILL FILL_40_DFFSR_82 ( );
FILL FILL_41_DFFSR_82 ( );
FILL FILL_42_DFFSR_82 ( );
FILL FILL_43_DFFSR_82 ( );
FILL FILL_44_DFFSR_82 ( );
FILL FILL_45_DFFSR_82 ( );
FILL FILL_46_DFFSR_82 ( );
FILL FILL_47_DFFSR_82 ( );
FILL FILL_48_DFFSR_82 ( );
FILL FILL_49_DFFSR_82 ( );
FILL FILL_50_DFFSR_82 ( );
FILL FILL_0_NAND2X1_98 ( );
FILL FILL_1_NAND2X1_98 ( );
FILL FILL_2_NAND2X1_98 ( );
FILL FILL_3_NAND2X1_98 ( );
FILL FILL_4_NAND2X1_98 ( );
FILL FILL_5_NAND2X1_98 ( );
FILL FILL_6_NAND2X1_98 ( );
FILL FILL_0_OAI21X1_98 ( );
FILL FILL_1_OAI21X1_98 ( );
FILL FILL_2_OAI21X1_98 ( );
FILL FILL_3_OAI21X1_98 ( );
FILL FILL_4_OAI21X1_98 ( );
FILL FILL_5_OAI21X1_98 ( );
FILL FILL_6_OAI21X1_98 ( );
FILL FILL_7_OAI21X1_98 ( );
FILL FILL_8_OAI21X1_98 ( );
FILL FILL_9_OAI21X1_98 ( );
FILL FILL_0_INVX1_111 ( );
FILL FILL_1_INVX1_111 ( );
FILL FILL_2_INVX1_111 ( );
FILL FILL_3_INVX1_111 ( );
FILL FILL_0_OAI21X1_106 ( );
FILL FILL_1_OAI21X1_106 ( );
FILL FILL_2_OAI21X1_106 ( );
FILL FILL_3_OAI21X1_106 ( );
FILL FILL_4_OAI21X1_106 ( );
FILL FILL_5_OAI21X1_106 ( );
FILL FILL_6_OAI21X1_106 ( );
FILL FILL_7_OAI21X1_106 ( );
FILL FILL_8_OAI21X1_106 ( );
FILL FILL_0_NAND2X1_106 ( );
FILL FILL_1_NAND2X1_106 ( );
FILL FILL_2_NAND2X1_106 ( );
FILL FILL_3_NAND2X1_106 ( );
FILL FILL_4_NAND2X1_106 ( );
FILL FILL_5_NAND2X1_106 ( );
FILL FILL_6_NAND2X1_106 ( );
FILL FILL_0_DFFPOSX1_29 ( );
FILL FILL_1_DFFPOSX1_29 ( );
FILL FILL_2_DFFPOSX1_29 ( );
FILL FILL_3_DFFPOSX1_29 ( );
FILL FILL_4_DFFPOSX1_29 ( );
FILL FILL_5_DFFPOSX1_29 ( );
FILL FILL_6_DFFPOSX1_29 ( );
FILL FILL_7_DFFPOSX1_29 ( );
FILL FILL_8_DFFPOSX1_29 ( );
FILL FILL_9_DFFPOSX1_29 ( );
FILL FILL_10_DFFPOSX1_29 ( );
FILL FILL_11_DFFPOSX1_29 ( );
FILL FILL_12_DFFPOSX1_29 ( );
FILL FILL_13_DFFPOSX1_29 ( );
FILL FILL_14_DFFPOSX1_29 ( );
FILL FILL_15_DFFPOSX1_29 ( );
FILL FILL_16_DFFPOSX1_29 ( );
FILL FILL_17_DFFPOSX1_29 ( );
FILL FILL_18_DFFPOSX1_29 ( );
FILL FILL_19_DFFPOSX1_29 ( );
FILL FILL_20_DFFPOSX1_29 ( );
FILL FILL_21_DFFPOSX1_29 ( );
FILL FILL_22_DFFPOSX1_29 ( );
FILL FILL_23_DFFPOSX1_29 ( );
FILL FILL_24_DFFPOSX1_29 ( );
FILL FILL_25_DFFPOSX1_29 ( );
FILL FILL_26_DFFPOSX1_29 ( );
FILL FILL_27_DFFPOSX1_29 ( );
FILL FILL_0_NOR2X1_54 ( );
FILL FILL_1_NOR2X1_54 ( );
FILL FILL_2_NOR2X1_54 ( );
FILL FILL_3_NOR2X1_54 ( );
FILL FILL_4_NOR2X1_54 ( );
FILL FILL_5_NOR2X1_54 ( );
FILL FILL_6_NOR2X1_54 ( );
FILL FILL_0_INVX1_148 ( );
FILL FILL_1_INVX1_148 ( );
FILL FILL_2_INVX1_148 ( );
FILL FILL_3_INVX1_148 ( );
FILL FILL_0_OAI21X1_26 ( );
FILL FILL_1_OAI21X1_26 ( );
FILL FILL_2_OAI21X1_26 ( );
FILL FILL_3_OAI21X1_26 ( );
FILL FILL_4_OAI21X1_26 ( );
FILL FILL_5_OAI21X1_26 ( );
FILL FILL_6_OAI21X1_26 ( );
FILL FILL_7_OAI21X1_26 ( );
FILL FILL_8_OAI21X1_26 ( );
FILL FILL_0_INVX1_30 ( );
FILL FILL_1_INVX1_30 ( );
FILL FILL_2_INVX1_30 ( );
FILL FILL_3_INVX1_30 ( );
FILL FILL_4_INVX1_30 ( );
FILL FILL_0_NAND2X1_26 ( );
FILL FILL_1_NAND2X1_26 ( );
FILL FILL_2_NAND2X1_26 ( );
FILL FILL_3_NAND2X1_26 ( );
FILL FILL_4_NAND2X1_26 ( );
FILL FILL_5_NAND2X1_26 ( );
FILL FILL_6_NAND2X1_26 ( );
FILL FILL_0_DFFSR_34 ( );
FILL FILL_1_DFFSR_34 ( );
FILL FILL_2_DFFSR_34 ( );
FILL FILL_3_DFFSR_34 ( );
FILL FILL_4_DFFSR_34 ( );
FILL FILL_5_DFFSR_34 ( );
FILL FILL_6_DFFSR_34 ( );
FILL FILL_7_DFFSR_34 ( );
FILL FILL_8_DFFSR_34 ( );
FILL FILL_9_DFFSR_34 ( );
FILL FILL_10_DFFSR_34 ( );
FILL FILL_11_DFFSR_34 ( );
FILL FILL_12_DFFSR_34 ( );
FILL FILL_13_DFFSR_34 ( );
FILL FILL_14_DFFSR_34 ( );
FILL FILL_15_DFFSR_34 ( );
FILL FILL_16_DFFSR_34 ( );
FILL FILL_17_DFFSR_34 ( );
FILL FILL_18_DFFSR_34 ( );
FILL FILL_19_DFFSR_34 ( );
FILL FILL_20_DFFSR_34 ( );
FILL FILL_21_DFFSR_34 ( );
FILL FILL_22_DFFSR_34 ( );
FILL FILL_23_DFFSR_34 ( );
FILL FILL_24_DFFSR_34 ( );
FILL FILL_25_DFFSR_34 ( );
FILL FILL_26_DFFSR_34 ( );
FILL FILL_27_DFFSR_34 ( );
FILL FILL_28_DFFSR_34 ( );
FILL FILL_29_DFFSR_34 ( );
FILL FILL_30_DFFSR_34 ( );
FILL FILL_31_DFFSR_34 ( );
FILL FILL_32_DFFSR_34 ( );
FILL FILL_33_DFFSR_34 ( );
FILL FILL_34_DFFSR_34 ( );
FILL FILL_35_DFFSR_34 ( );
FILL FILL_36_DFFSR_34 ( );
FILL FILL_37_DFFSR_34 ( );
FILL FILL_38_DFFSR_34 ( );
FILL FILL_39_DFFSR_34 ( );
FILL FILL_40_DFFSR_34 ( );
FILL FILL_41_DFFSR_34 ( );
FILL FILL_42_DFFSR_34 ( );
FILL FILL_43_DFFSR_34 ( );
FILL FILL_44_DFFSR_34 ( );
FILL FILL_45_DFFSR_34 ( );
FILL FILL_46_DFFSR_34 ( );
FILL FILL_47_DFFSR_34 ( );
FILL FILL_48_DFFSR_34 ( );
FILL FILL_49_DFFSR_34 ( );
FILL FILL_50_DFFSR_34 ( );
FILL FILL_0_INVX1_21 ( );
FILL FILL_1_INVX1_21 ( );
FILL FILL_2_INVX1_21 ( );
FILL FILL_3_INVX1_21 ( );
FILL FILL_4_INVX1_21 ( );
FILL FILL_0_NAND2X1_18 ( );
FILL FILL_1_NAND2X1_18 ( );
FILL FILL_2_NAND2X1_18 ( );
FILL FILL_3_NAND2X1_18 ( );
FILL FILL_4_NAND2X1_18 ( );
FILL FILL_5_NAND2X1_18 ( );
FILL FILL_6_NAND2X1_18 ( );
FILL FILL_0_DFFSR_19 ( );
FILL FILL_1_DFFSR_19 ( );
FILL FILL_2_DFFSR_19 ( );
FILL FILL_3_DFFSR_19 ( );
FILL FILL_4_DFFSR_19 ( );
FILL FILL_5_DFFSR_19 ( );
FILL FILL_6_DFFSR_19 ( );
FILL FILL_7_DFFSR_19 ( );
FILL FILL_8_DFFSR_19 ( );
FILL FILL_9_DFFSR_19 ( );
FILL FILL_10_DFFSR_19 ( );
FILL FILL_11_DFFSR_19 ( );
FILL FILL_12_DFFSR_19 ( );
FILL FILL_13_DFFSR_19 ( );
FILL FILL_14_DFFSR_19 ( );
FILL FILL_15_DFFSR_19 ( );
FILL FILL_16_DFFSR_19 ( );
FILL FILL_17_DFFSR_19 ( );
FILL FILL_18_DFFSR_19 ( );
FILL FILL_19_DFFSR_19 ( );
FILL FILL_20_DFFSR_19 ( );
FILL FILL_21_DFFSR_19 ( );
FILL FILL_22_DFFSR_19 ( );
FILL FILL_23_DFFSR_19 ( );
FILL FILL_24_DFFSR_19 ( );
FILL FILL_25_DFFSR_19 ( );
FILL FILL_26_DFFSR_19 ( );
FILL FILL_27_DFFSR_19 ( );
FILL FILL_28_DFFSR_19 ( );
FILL FILL_29_DFFSR_19 ( );
FILL FILL_30_DFFSR_19 ( );
FILL FILL_31_DFFSR_19 ( );
FILL FILL_32_DFFSR_19 ( );
FILL FILL_33_DFFSR_19 ( );
FILL FILL_34_DFFSR_19 ( );
FILL FILL_35_DFFSR_19 ( );
FILL FILL_36_DFFSR_19 ( );
FILL FILL_37_DFFSR_19 ( );
FILL FILL_38_DFFSR_19 ( );
FILL FILL_39_DFFSR_19 ( );
FILL FILL_40_DFFSR_19 ( );
FILL FILL_41_DFFSR_19 ( );
FILL FILL_42_DFFSR_19 ( );
FILL FILL_43_DFFSR_19 ( );
FILL FILL_44_DFFSR_19 ( );
FILL FILL_45_DFFSR_19 ( );
FILL FILL_46_DFFSR_19 ( );
FILL FILL_47_DFFSR_19 ( );
FILL FILL_48_DFFSR_19 ( );
FILL FILL_49_DFFSR_19 ( );
FILL FILL_50_DFFSR_19 ( );
FILL FILL_51_DFFSR_19 ( );
FILL FILL_0_OAI21X1_9 ( );
FILL FILL_1_OAI21X1_9 ( );
FILL FILL_2_OAI21X1_9 ( );
FILL FILL_3_OAI21X1_9 ( );
FILL FILL_4_OAI21X1_9 ( );
FILL FILL_5_OAI21X1_9 ( );
FILL FILL_6_OAI21X1_9 ( );
FILL FILL_7_OAI21X1_9 ( );
FILL FILL_8_OAI21X1_9 ( );
FILL FILL_9_OAI21X1_9 ( );
FILL FILL_0_DFFSR_178 ( );
FILL FILL_1_DFFSR_178 ( );
FILL FILL_2_DFFSR_178 ( );
FILL FILL_3_DFFSR_178 ( );
FILL FILL_4_DFFSR_178 ( );
FILL FILL_5_DFFSR_178 ( );
FILL FILL_6_DFFSR_178 ( );
FILL FILL_7_DFFSR_178 ( );
FILL FILL_8_DFFSR_178 ( );
FILL FILL_9_DFFSR_178 ( );
FILL FILL_10_DFFSR_178 ( );
FILL FILL_11_DFFSR_178 ( );
FILL FILL_12_DFFSR_178 ( );
FILL FILL_13_DFFSR_178 ( );
FILL FILL_14_DFFSR_178 ( );
FILL FILL_15_DFFSR_178 ( );
FILL FILL_16_DFFSR_178 ( );
FILL FILL_17_DFFSR_178 ( );
FILL FILL_18_DFFSR_178 ( );
FILL FILL_19_DFFSR_178 ( );
FILL FILL_20_DFFSR_178 ( );
FILL FILL_21_DFFSR_178 ( );
FILL FILL_22_DFFSR_178 ( );
FILL FILL_23_DFFSR_178 ( );
FILL FILL_24_DFFSR_178 ( );
FILL FILL_25_DFFSR_178 ( );
FILL FILL_26_DFFSR_178 ( );
FILL FILL_27_DFFSR_178 ( );
FILL FILL_28_DFFSR_178 ( );
FILL FILL_29_DFFSR_178 ( );
FILL FILL_30_DFFSR_178 ( );
FILL FILL_31_DFFSR_178 ( );
FILL FILL_32_DFFSR_178 ( );
FILL FILL_33_DFFSR_178 ( );
FILL FILL_34_DFFSR_178 ( );
FILL FILL_35_DFFSR_178 ( );
FILL FILL_36_DFFSR_178 ( );
FILL FILL_37_DFFSR_178 ( );
FILL FILL_38_DFFSR_178 ( );
FILL FILL_39_DFFSR_178 ( );
FILL FILL_40_DFFSR_178 ( );
FILL FILL_41_DFFSR_178 ( );
FILL FILL_42_DFFSR_178 ( );
FILL FILL_43_DFFSR_178 ( );
FILL FILL_44_DFFSR_178 ( );
FILL FILL_45_DFFSR_178 ( );
FILL FILL_46_DFFSR_178 ( );
FILL FILL_47_DFFSR_178 ( );
FILL FILL_48_DFFSR_178 ( );
FILL FILL_49_DFFSR_178 ( );
FILL FILL_50_DFFSR_178 ( );
FILL FILL_0_DFFSR_184 ( );
FILL FILL_1_DFFSR_184 ( );
FILL FILL_2_DFFSR_184 ( );
FILL FILL_3_DFFSR_184 ( );
FILL FILL_4_DFFSR_184 ( );
FILL FILL_5_DFFSR_184 ( );
FILL FILL_6_DFFSR_184 ( );
FILL FILL_7_DFFSR_184 ( );
FILL FILL_8_DFFSR_184 ( );
FILL FILL_9_DFFSR_184 ( );
FILL FILL_10_DFFSR_184 ( );
FILL FILL_11_DFFSR_184 ( );
FILL FILL_12_DFFSR_184 ( );
FILL FILL_13_DFFSR_184 ( );
FILL FILL_14_DFFSR_184 ( );
FILL FILL_15_DFFSR_184 ( );
FILL FILL_16_DFFSR_184 ( );
FILL FILL_17_DFFSR_184 ( );
FILL FILL_18_DFFSR_184 ( );
FILL FILL_19_DFFSR_184 ( );
FILL FILL_20_DFFSR_184 ( );
FILL FILL_21_DFFSR_184 ( );
FILL FILL_22_DFFSR_184 ( );
FILL FILL_23_DFFSR_184 ( );
FILL FILL_24_DFFSR_184 ( );
FILL FILL_25_DFFSR_184 ( );
FILL FILL_26_DFFSR_184 ( );
FILL FILL_27_DFFSR_184 ( );
FILL FILL_28_DFFSR_184 ( );
FILL FILL_29_DFFSR_184 ( );
FILL FILL_30_DFFSR_184 ( );
FILL FILL_31_DFFSR_184 ( );
FILL FILL_32_DFFSR_184 ( );
FILL FILL_33_DFFSR_184 ( );
FILL FILL_34_DFFSR_184 ( );
FILL FILL_35_DFFSR_184 ( );
FILL FILL_36_DFFSR_184 ( );
FILL FILL_37_DFFSR_184 ( );
FILL FILL_38_DFFSR_184 ( );
FILL FILL_39_DFFSR_184 ( );
FILL FILL_40_DFFSR_184 ( );
FILL FILL_41_DFFSR_184 ( );
FILL FILL_42_DFFSR_184 ( );
FILL FILL_43_DFFSR_184 ( );
FILL FILL_44_DFFSR_184 ( );
FILL FILL_45_DFFSR_184 ( );
FILL FILL_46_DFFSR_184 ( );
FILL FILL_47_DFFSR_184 ( );
FILL FILL_48_DFFSR_184 ( );
FILL FILL_49_DFFSR_184 ( );
FILL FILL_50_DFFSR_184 ( );
FILL FILL_0_INVX1_421 ( );
FILL FILL_1_INVX1_421 ( );
FILL FILL_2_INVX1_421 ( );
FILL FILL_3_INVX1_421 ( );
FILL FILL_4_INVX1_421 ( );
FILL FILL_0_BUFX2_31 ( );
FILL FILL_1_BUFX2_31 ( );
FILL FILL_2_BUFX2_31 ( );
FILL FILL_3_BUFX2_31 ( );
FILL FILL_4_BUFX2_31 ( );
FILL FILL_5_BUFX2_31 ( );
FILL FILL_6_BUFX2_31 ( );
FILL FILL_0_DFFSR_74 ( );
FILL FILL_1_DFFSR_74 ( );
FILL FILL_2_DFFSR_74 ( );
FILL FILL_3_DFFSR_74 ( );
FILL FILL_4_DFFSR_74 ( );
FILL FILL_5_DFFSR_74 ( );
FILL FILL_6_DFFSR_74 ( );
FILL FILL_7_DFFSR_74 ( );
FILL FILL_8_DFFSR_74 ( );
FILL FILL_9_DFFSR_74 ( );
FILL FILL_10_DFFSR_74 ( );
FILL FILL_11_DFFSR_74 ( );
FILL FILL_12_DFFSR_74 ( );
FILL FILL_13_DFFSR_74 ( );
FILL FILL_14_DFFSR_74 ( );
FILL FILL_15_DFFSR_74 ( );
FILL FILL_16_DFFSR_74 ( );
FILL FILL_17_DFFSR_74 ( );
FILL FILL_18_DFFSR_74 ( );
FILL FILL_19_DFFSR_74 ( );
FILL FILL_20_DFFSR_74 ( );
FILL FILL_21_DFFSR_74 ( );
FILL FILL_22_DFFSR_74 ( );
FILL FILL_23_DFFSR_74 ( );
FILL FILL_24_DFFSR_74 ( );
FILL FILL_25_DFFSR_74 ( );
FILL FILL_26_DFFSR_74 ( );
FILL FILL_27_DFFSR_74 ( );
FILL FILL_28_DFFSR_74 ( );
FILL FILL_29_DFFSR_74 ( );
FILL FILL_30_DFFSR_74 ( );
FILL FILL_31_DFFSR_74 ( );
FILL FILL_32_DFFSR_74 ( );
FILL FILL_33_DFFSR_74 ( );
FILL FILL_34_DFFSR_74 ( );
FILL FILL_35_DFFSR_74 ( );
FILL FILL_36_DFFSR_74 ( );
FILL FILL_37_DFFSR_74 ( );
FILL FILL_38_DFFSR_74 ( );
FILL FILL_39_DFFSR_74 ( );
FILL FILL_40_DFFSR_74 ( );
FILL FILL_41_DFFSR_74 ( );
FILL FILL_42_DFFSR_74 ( );
FILL FILL_43_DFFSR_74 ( );
FILL FILL_44_DFFSR_74 ( );
FILL FILL_45_DFFSR_74 ( );
FILL FILL_46_DFFSR_74 ( );
FILL FILL_47_DFFSR_74 ( );
FILL FILL_48_DFFSR_74 ( );
FILL FILL_49_DFFSR_74 ( );
FILL FILL_50_DFFSR_74 ( );
FILL FILL_51_DFFSR_74 ( );
FILL FILL_0_INVX1_84 ( );
FILL FILL_1_INVX1_84 ( );
FILL FILL_2_INVX1_84 ( );
FILL FILL_3_INVX1_84 ( );
FILL FILL_4_INVX1_84 ( );
FILL FILL_0_OAI21X1_74 ( );
FILL FILL_1_OAI21X1_74 ( );
FILL FILL_2_OAI21X1_74 ( );
FILL FILL_3_OAI21X1_74 ( );
FILL FILL_4_OAI21X1_74 ( );
FILL FILL_5_OAI21X1_74 ( );
FILL FILL_6_OAI21X1_74 ( );
FILL FILL_7_OAI21X1_74 ( );
FILL FILL_8_OAI21X1_74 ( );
FILL FILL_0_NAND2X1_82 ( );
FILL FILL_1_NAND2X1_82 ( );
FILL FILL_2_NAND2X1_82 ( );
FILL FILL_3_NAND2X1_82 ( );
FILL FILL_4_NAND2X1_82 ( );
FILL FILL_5_NAND2X1_82 ( );
FILL FILL_6_NAND2X1_82 ( );
FILL FILL_0_INVX1_93 ( );
FILL FILL_1_INVX1_93 ( );
FILL FILL_2_INVX1_93 ( );
FILL FILL_3_INVX1_93 ( );
FILL FILL_0_OAI21X1_82 ( );
FILL FILL_1_OAI21X1_82 ( );
FILL FILL_2_OAI21X1_82 ( );
FILL FILL_3_OAI21X1_82 ( );
FILL FILL_4_OAI21X1_82 ( );
FILL FILL_5_OAI21X1_82 ( );
FILL FILL_6_OAI21X1_82 ( );
FILL FILL_7_OAI21X1_82 ( );
FILL FILL_8_OAI21X1_82 ( );
FILL FILL_9_OAI21X1_82 ( );
FILL FILL_0_DFFSR_98 ( );
FILL FILL_1_DFFSR_98 ( );
FILL FILL_2_DFFSR_98 ( );
FILL FILL_3_DFFSR_98 ( );
FILL FILL_4_DFFSR_98 ( );
FILL FILL_5_DFFSR_98 ( );
FILL FILL_6_DFFSR_98 ( );
FILL FILL_7_DFFSR_98 ( );
FILL FILL_8_DFFSR_98 ( );
FILL FILL_9_DFFSR_98 ( );
FILL FILL_10_DFFSR_98 ( );
FILL FILL_11_DFFSR_98 ( );
FILL FILL_12_DFFSR_98 ( );
FILL FILL_13_DFFSR_98 ( );
FILL FILL_14_DFFSR_98 ( );
FILL FILL_15_DFFSR_98 ( );
FILL FILL_16_DFFSR_98 ( );
FILL FILL_17_DFFSR_98 ( );
FILL FILL_18_DFFSR_98 ( );
FILL FILL_19_DFFSR_98 ( );
FILL FILL_20_DFFSR_98 ( );
FILL FILL_21_DFFSR_98 ( );
FILL FILL_22_DFFSR_98 ( );
FILL FILL_23_DFFSR_98 ( );
FILL FILL_24_DFFSR_98 ( );
FILL FILL_25_DFFSR_98 ( );
FILL FILL_26_DFFSR_98 ( );
FILL FILL_27_DFFSR_98 ( );
FILL FILL_28_DFFSR_98 ( );
FILL FILL_29_DFFSR_98 ( );
FILL FILL_30_DFFSR_98 ( );
FILL FILL_31_DFFSR_98 ( );
FILL FILL_32_DFFSR_98 ( );
FILL FILL_33_DFFSR_98 ( );
FILL FILL_34_DFFSR_98 ( );
FILL FILL_35_DFFSR_98 ( );
FILL FILL_36_DFFSR_98 ( );
FILL FILL_37_DFFSR_98 ( );
FILL FILL_38_DFFSR_98 ( );
FILL FILL_39_DFFSR_98 ( );
FILL FILL_40_DFFSR_98 ( );
FILL FILL_41_DFFSR_98 ( );
FILL FILL_42_DFFSR_98 ( );
FILL FILL_43_DFFSR_98 ( );
FILL FILL_44_DFFSR_98 ( );
FILL FILL_45_DFFSR_98 ( );
FILL FILL_46_DFFSR_98 ( );
FILL FILL_47_DFFSR_98 ( );
FILL FILL_48_DFFSR_98 ( );
FILL FILL_49_DFFSR_98 ( );
FILL FILL_50_DFFSR_98 ( );
FILL FILL_0_NAND2X1_131 ( );
FILL FILL_1_NAND2X1_131 ( );
FILL FILL_2_NAND2X1_131 ( );
FILL FILL_3_NAND2X1_131 ( );
FILL FILL_4_NAND2X1_131 ( );
FILL FILL_5_NAND2X1_131 ( );
FILL FILL_6_NAND2X1_131 ( );
FILL FILL_0_OAI21X1_131 ( );
FILL FILL_1_OAI21X1_131 ( );
FILL FILL_2_OAI21X1_131 ( );
FILL FILL_3_OAI21X1_131 ( );
FILL FILL_4_OAI21X1_131 ( );
FILL FILL_5_OAI21X1_131 ( );
FILL FILL_6_OAI21X1_131 ( );
FILL FILL_7_OAI21X1_131 ( );
FILL FILL_8_OAI21X1_131 ( );
FILL FILL_9_OAI21X1_131 ( );
FILL FILL_0_DFFSR_26 ( );
FILL FILL_1_DFFSR_26 ( );
FILL FILL_2_DFFSR_26 ( );
FILL FILL_3_DFFSR_26 ( );
FILL FILL_4_DFFSR_26 ( );
FILL FILL_5_DFFSR_26 ( );
FILL FILL_6_DFFSR_26 ( );
FILL FILL_7_DFFSR_26 ( );
FILL FILL_8_DFFSR_26 ( );
FILL FILL_9_DFFSR_26 ( );
FILL FILL_10_DFFSR_26 ( );
FILL FILL_11_DFFSR_26 ( );
FILL FILL_12_DFFSR_26 ( );
FILL FILL_13_DFFSR_26 ( );
FILL FILL_14_DFFSR_26 ( );
FILL FILL_15_DFFSR_26 ( );
FILL FILL_16_DFFSR_26 ( );
FILL FILL_17_DFFSR_26 ( );
FILL FILL_18_DFFSR_26 ( );
FILL FILL_19_DFFSR_26 ( );
FILL FILL_20_DFFSR_26 ( );
FILL FILL_21_DFFSR_26 ( );
FILL FILL_22_DFFSR_26 ( );
FILL FILL_23_DFFSR_26 ( );
FILL FILL_24_DFFSR_26 ( );
FILL FILL_25_DFFSR_26 ( );
FILL FILL_26_DFFSR_26 ( );
FILL FILL_27_DFFSR_26 ( );
FILL FILL_28_DFFSR_26 ( );
FILL FILL_29_DFFSR_26 ( );
FILL FILL_30_DFFSR_26 ( );
FILL FILL_31_DFFSR_26 ( );
FILL FILL_32_DFFSR_26 ( );
FILL FILL_33_DFFSR_26 ( );
FILL FILL_34_DFFSR_26 ( );
FILL FILL_35_DFFSR_26 ( );
FILL FILL_36_DFFSR_26 ( );
FILL FILL_37_DFFSR_26 ( );
FILL FILL_38_DFFSR_26 ( );
FILL FILL_39_DFFSR_26 ( );
FILL FILL_40_DFFSR_26 ( );
FILL FILL_41_DFFSR_26 ( );
FILL FILL_42_DFFSR_26 ( );
FILL FILL_43_DFFSR_26 ( );
FILL FILL_44_DFFSR_26 ( );
FILL FILL_45_DFFSR_26 ( );
FILL FILL_46_DFFSR_26 ( );
FILL FILL_47_DFFSR_26 ( );
FILL FILL_48_DFFSR_26 ( );
FILL FILL_49_DFFSR_26 ( );
FILL FILL_50_DFFSR_26 ( );
FILL FILL_51_DFFSR_26 ( );
FILL FILL_0_DFFSR_18 ( );
FILL FILL_1_DFFSR_18 ( );
FILL FILL_2_DFFSR_18 ( );
FILL FILL_3_DFFSR_18 ( );
FILL FILL_4_DFFSR_18 ( );
FILL FILL_5_DFFSR_18 ( );
FILL FILL_6_DFFSR_18 ( );
FILL FILL_7_DFFSR_18 ( );
FILL FILL_8_DFFSR_18 ( );
FILL FILL_9_DFFSR_18 ( );
FILL FILL_10_DFFSR_18 ( );
FILL FILL_11_DFFSR_18 ( );
FILL FILL_12_DFFSR_18 ( );
FILL FILL_13_DFFSR_18 ( );
FILL FILL_14_DFFSR_18 ( );
FILL FILL_15_DFFSR_18 ( );
FILL FILL_16_DFFSR_18 ( );
FILL FILL_17_DFFSR_18 ( );
FILL FILL_18_DFFSR_18 ( );
FILL FILL_19_DFFSR_18 ( );
FILL FILL_20_DFFSR_18 ( );
FILL FILL_21_DFFSR_18 ( );
FILL FILL_22_DFFSR_18 ( );
FILL FILL_23_DFFSR_18 ( );
FILL FILL_24_DFFSR_18 ( );
FILL FILL_25_DFFSR_18 ( );
FILL FILL_26_DFFSR_18 ( );
FILL FILL_27_DFFSR_18 ( );
FILL FILL_28_DFFSR_18 ( );
FILL FILL_29_DFFSR_18 ( );
FILL FILL_30_DFFSR_18 ( );
FILL FILL_31_DFFSR_18 ( );
FILL FILL_32_DFFSR_18 ( );
FILL FILL_33_DFFSR_18 ( );
FILL FILL_34_DFFSR_18 ( );
FILL FILL_35_DFFSR_18 ( );
FILL FILL_36_DFFSR_18 ( );
FILL FILL_37_DFFSR_18 ( );
FILL FILL_38_DFFSR_18 ( );
FILL FILL_39_DFFSR_18 ( );
FILL FILL_40_DFFSR_18 ( );
FILL FILL_41_DFFSR_18 ( );
FILL FILL_42_DFFSR_18 ( );
FILL FILL_43_DFFSR_18 ( );
FILL FILL_44_DFFSR_18 ( );
FILL FILL_45_DFFSR_18 ( );
FILL FILL_46_DFFSR_18 ( );
FILL FILL_47_DFFSR_18 ( );
FILL FILL_48_DFFSR_18 ( );
FILL FILL_49_DFFSR_18 ( );
FILL FILL_50_DFFSR_18 ( );
FILL FILL_0_OAI21X1_18 ( );
FILL FILL_1_OAI21X1_18 ( );
FILL FILL_2_OAI21X1_18 ( );
FILL FILL_3_OAI21X1_18 ( );
FILL FILL_4_OAI21X1_18 ( );
FILL FILL_5_OAI21X1_18 ( );
FILL FILL_6_OAI21X1_18 ( );
FILL FILL_7_OAI21X1_18 ( );
FILL FILL_8_OAI21X1_18 ( );
FILL FILL_0_DFFSR_9 ( );
FILL FILL_1_DFFSR_9 ( );
FILL FILL_2_DFFSR_9 ( );
FILL FILL_3_DFFSR_9 ( );
FILL FILL_4_DFFSR_9 ( );
FILL FILL_5_DFFSR_9 ( );
FILL FILL_6_DFFSR_9 ( );
FILL FILL_7_DFFSR_9 ( );
FILL FILL_8_DFFSR_9 ( );
FILL FILL_9_DFFSR_9 ( );
FILL FILL_10_DFFSR_9 ( );
FILL FILL_11_DFFSR_9 ( );
FILL FILL_12_DFFSR_9 ( );
FILL FILL_13_DFFSR_9 ( );
FILL FILL_14_DFFSR_9 ( );
FILL FILL_15_DFFSR_9 ( );
FILL FILL_16_DFFSR_9 ( );
FILL FILL_17_DFFSR_9 ( );
FILL FILL_18_DFFSR_9 ( );
FILL FILL_19_DFFSR_9 ( );
FILL FILL_20_DFFSR_9 ( );
FILL FILL_21_DFFSR_9 ( );
FILL FILL_22_DFFSR_9 ( );
FILL FILL_23_DFFSR_9 ( );
FILL FILL_24_DFFSR_9 ( );
FILL FILL_25_DFFSR_9 ( );
FILL FILL_26_DFFSR_9 ( );
FILL FILL_27_DFFSR_9 ( );
FILL FILL_28_DFFSR_9 ( );
FILL FILL_29_DFFSR_9 ( );
FILL FILL_30_DFFSR_9 ( );
FILL FILL_31_DFFSR_9 ( );
FILL FILL_32_DFFSR_9 ( );
FILL FILL_33_DFFSR_9 ( );
FILL FILL_34_DFFSR_9 ( );
FILL FILL_35_DFFSR_9 ( );
FILL FILL_36_DFFSR_9 ( );
FILL FILL_37_DFFSR_9 ( );
FILL FILL_38_DFFSR_9 ( );
FILL FILL_39_DFFSR_9 ( );
FILL FILL_40_DFFSR_9 ( );
FILL FILL_41_DFFSR_9 ( );
FILL FILL_42_DFFSR_9 ( );
FILL FILL_43_DFFSR_9 ( );
FILL FILL_44_DFFSR_9 ( );
FILL FILL_45_DFFSR_9 ( );
FILL FILL_46_DFFSR_9 ( );
FILL FILL_47_DFFSR_9 ( );
FILL FILL_48_DFFSR_9 ( );
FILL FILL_49_DFFSR_9 ( );
FILL FILL_50_DFFSR_9 ( );
FILL FILL_51_DFFSR_9 ( );
FILL FILL_0_NAND2X1_257 ( );
FILL FILL_1_NAND2X1_257 ( );
FILL FILL_2_NAND2X1_257 ( );
FILL FILL_3_NAND2X1_257 ( );
FILL FILL_4_NAND2X1_257 ( );
FILL FILL_5_NAND2X1_257 ( );
FILL FILL_6_NAND2X1_257 ( );
FILL FILL_0_OAI21X1_246 ( );
FILL FILL_1_OAI21X1_246 ( );
FILL FILL_2_OAI21X1_246 ( );
FILL FILL_3_OAI21X1_246 ( );
FILL FILL_4_OAI21X1_246 ( );
FILL FILL_5_OAI21X1_246 ( );
FILL FILL_6_OAI21X1_246 ( );
FILL FILL_7_OAI21X1_246 ( );
FILL FILL_8_OAI21X1_246 ( );
FILL FILL_9_OAI21X1_246 ( );
FILL FILL_0_INVX1_408 ( );
FILL FILL_1_INVX1_408 ( );
FILL FILL_2_INVX1_408 ( );
FILL FILL_3_INVX1_408 ( );
FILL FILL_0_CLKBUF1_19 ( );
FILL FILL_1_CLKBUF1_19 ( );
FILL FILL_2_CLKBUF1_19 ( );
FILL FILL_3_CLKBUF1_19 ( );
FILL FILL_4_CLKBUF1_19 ( );
FILL FILL_5_CLKBUF1_19 ( );
FILL FILL_6_CLKBUF1_19 ( );
FILL FILL_7_CLKBUF1_19 ( );
FILL FILL_8_CLKBUF1_19 ( );
FILL FILL_9_CLKBUF1_19 ( );
FILL FILL_10_CLKBUF1_19 ( );
FILL FILL_11_CLKBUF1_19 ( );
FILL FILL_12_CLKBUF1_19 ( );
FILL FILL_13_CLKBUF1_19 ( );
FILL FILL_14_CLKBUF1_19 ( );
FILL FILL_15_CLKBUF1_19 ( );
FILL FILL_16_CLKBUF1_19 ( );
FILL FILL_17_CLKBUF1_19 ( );
FILL FILL_18_CLKBUF1_19 ( );
FILL FILL_19_CLKBUF1_19 ( );
FILL FILL_20_CLKBUF1_19 ( );
FILL FILL_0_BUFX2_26 ( );
FILL FILL_1_BUFX2_26 ( );
FILL FILL_2_BUFX2_26 ( );
FILL FILL_3_BUFX2_26 ( );
FILL FILL_4_BUFX2_26 ( );
FILL FILL_5_BUFX2_26 ( );
FILL FILL_6_BUFX2_26 ( );
FILL FILL_0_NAND2X1_258 ( );
FILL FILL_1_NAND2X1_258 ( );
FILL FILL_2_NAND2X1_258 ( );
FILL FILL_3_NAND2X1_258 ( );
FILL FILL_4_NAND2X1_258 ( );
FILL FILL_5_NAND2X1_258 ( );
FILL FILL_6_NAND2X1_258 ( );
FILL FILL_0_INVX1_415 ( );
FILL FILL_1_INVX1_415 ( );
FILL FILL_2_INVX1_415 ( );
FILL FILL_3_INVX1_415 ( );
FILL FILL_4_INVX1_415 ( );
FILL FILL_0_DFFSR_190 ( );
FILL FILL_1_DFFSR_190 ( );
FILL FILL_2_DFFSR_190 ( );
FILL FILL_3_DFFSR_190 ( );
FILL FILL_4_DFFSR_190 ( );
FILL FILL_5_DFFSR_190 ( );
FILL FILL_6_DFFSR_190 ( );
FILL FILL_7_DFFSR_190 ( );
FILL FILL_8_DFFSR_190 ( );
FILL FILL_9_DFFSR_190 ( );
FILL FILL_10_DFFSR_190 ( );
FILL FILL_11_DFFSR_190 ( );
FILL FILL_12_DFFSR_190 ( );
FILL FILL_13_DFFSR_190 ( );
FILL FILL_14_DFFSR_190 ( );
FILL FILL_15_DFFSR_190 ( );
FILL FILL_16_DFFSR_190 ( );
FILL FILL_17_DFFSR_190 ( );
FILL FILL_18_DFFSR_190 ( );
FILL FILL_19_DFFSR_190 ( );
FILL FILL_20_DFFSR_190 ( );
FILL FILL_21_DFFSR_190 ( );
FILL FILL_22_DFFSR_190 ( );
FILL FILL_23_DFFSR_190 ( );
FILL FILL_24_DFFSR_190 ( );
FILL FILL_25_DFFSR_190 ( );
FILL FILL_26_DFFSR_190 ( );
FILL FILL_27_DFFSR_190 ( );
FILL FILL_28_DFFSR_190 ( );
FILL FILL_29_DFFSR_190 ( );
FILL FILL_30_DFFSR_190 ( );
FILL FILL_31_DFFSR_190 ( );
FILL FILL_32_DFFSR_190 ( );
FILL FILL_33_DFFSR_190 ( );
FILL FILL_34_DFFSR_190 ( );
FILL FILL_35_DFFSR_190 ( );
FILL FILL_36_DFFSR_190 ( );
FILL FILL_37_DFFSR_190 ( );
FILL FILL_38_DFFSR_190 ( );
FILL FILL_39_DFFSR_190 ( );
FILL FILL_40_DFFSR_190 ( );
FILL FILL_41_DFFSR_190 ( );
FILL FILL_42_DFFSR_190 ( );
FILL FILL_43_DFFSR_190 ( );
FILL FILL_44_DFFSR_190 ( );
FILL FILL_45_DFFSR_190 ( );
FILL FILL_46_DFFSR_190 ( );
FILL FILL_47_DFFSR_190 ( );
FILL FILL_48_DFFSR_190 ( );
FILL FILL_49_DFFSR_190 ( );
FILL FILL_50_DFFSR_190 ( );
FILL FILL_0_BUFX2_32 ( );
FILL FILL_1_BUFX2_32 ( );
FILL FILL_2_BUFX2_32 ( );
FILL FILL_3_BUFX2_32 ( );
FILL FILL_4_BUFX2_32 ( );
FILL FILL_5_BUFX2_32 ( );
FILL FILL_6_BUFX2_32 ( );
FILL FILL_0_NAND2X1_167 ( );
FILL FILL_1_NAND2X1_167 ( );
FILL FILL_2_NAND2X1_167 ( );
FILL FILL_3_NAND2X1_167 ( );
FILL FILL_4_NAND2X1_167 ( );
FILL FILL_5_NAND2X1_167 ( );
FILL FILL_6_NAND2X1_167 ( );
FILL FILL_0_0_0 ( );
FILL FILL_0_0_1 ( );
FILL FILL_0_0_2 ( );
FILL FILL_0_1_0 ( );
FILL FILL_0_1_1 ( );
FILL FILL_0_1_2 ( );
FILL FILL_0_2_0 ( );
FILL FILL_0_2_1 ( );
FILL FILL_0_2_2 ( );
FILL FILL_0_3_0 ( );
FILL FILL_0_3_1 ( );
FILL FILL_0_3_2 ( );
FILL FILL_0_4_0 ( );
FILL FILL_0_4_1 ( );
FILL FILL_0_4_2 ( );
FILL FILL_0_5_0 ( );
FILL FILL_0_5_1 ( );
FILL FILL_0_5_2 ( );
FILL FILL_1_1 ( );
FILL FILL_1_2 ( );
FILL FILL_1_3 ( );
FILL FILL_1_0_0 ( );
FILL FILL_1_0_1 ( );
FILL FILL_1_0_2 ( );
FILL FILL_1_1_0 ( );
FILL FILL_1_1_1 ( );
FILL FILL_1_1_2 ( );
FILL FILL_1_2_0 ( );
FILL FILL_1_2_1 ( );
FILL FILL_1_2_2 ( );
FILL FILL_1_3_0 ( );
FILL FILL_1_3_1 ( );
FILL FILL_1_3_2 ( );
FILL FILL_1_4_0 ( );
FILL FILL_1_4_1 ( );
FILL FILL_1_4_2 ( );
FILL FILL_1_5_0 ( );
FILL FILL_1_5_1 ( );
FILL FILL_1_5_2 ( );
FILL FILL_2_1 ( );
FILL FILL_2_2 ( );
FILL FILL_2_3 ( );
FILL FILL_2_4 ( );
FILL FILL_2_0_0 ( );
FILL FILL_2_0_1 ( );
FILL FILL_2_0_2 ( );
FILL FILL_2_1_0 ( );
FILL FILL_2_1_1 ( );
FILL FILL_2_1_2 ( );
FILL FILL_2_2_0 ( );
FILL FILL_2_2_1 ( );
FILL FILL_2_2_2 ( );
FILL FILL_2_3_0 ( );
FILL FILL_2_3_1 ( );
FILL FILL_2_3_2 ( );
FILL FILL_2_4_0 ( );
FILL FILL_2_4_1 ( );
FILL FILL_2_4_2 ( );
FILL FILL_2_5_0 ( );
FILL FILL_2_5_1 ( );
FILL FILL_2_5_2 ( );
FILL FILL_3_1 ( );
FILL FILL_3_2 ( );
FILL FILL_3_3 ( );
FILL FILL_3_0_0 ( );
FILL FILL_3_0_1 ( );
FILL FILL_3_0_2 ( );
FILL FILL_3_1_0 ( );
FILL FILL_3_1_1 ( );
FILL FILL_3_1_2 ( );
FILL FILL_3_2_0 ( );
FILL FILL_3_2_1 ( );
FILL FILL_3_2_2 ( );
FILL FILL_3_3_0 ( );
FILL FILL_3_3_1 ( );
FILL FILL_3_3_2 ( );
FILL FILL_3_4_0 ( );
FILL FILL_3_4_1 ( );
FILL FILL_3_4_2 ( );
FILL FILL_3_5_0 ( );
FILL FILL_3_5_1 ( );
FILL FILL_3_5_2 ( );
FILL FILL_4_1 ( );
FILL FILL_4_2 ( );
FILL FILL_4_3 ( );
FILL FILL_4_4 ( );
FILL FILL_4_5 ( );
FILL FILL_4_6 ( );
FILL FILL_4_7 ( );
FILL FILL_4_0_0 ( );
FILL FILL_4_0_1 ( );
FILL FILL_4_0_2 ( );
FILL FILL_4_1_0 ( );
FILL FILL_4_1_1 ( );
FILL FILL_4_1_2 ( );
FILL FILL_4_2_0 ( );
FILL FILL_4_2_1 ( );
FILL FILL_4_2_2 ( );
FILL FILL_4_3_0 ( );
FILL FILL_4_3_1 ( );
FILL FILL_4_3_2 ( );
FILL FILL_4_4_0 ( );
FILL FILL_4_4_1 ( );
FILL FILL_4_4_2 ( );
FILL FILL_4_5_0 ( );
FILL FILL_4_5_1 ( );
FILL FILL_4_5_2 ( );
FILL FILL_5_1 ( );
FILL FILL_5_2 ( );
FILL FILL_5_3 ( );
FILL FILL_5_4 ( );
FILL FILL_5_5 ( );
FILL FILL_5_6 ( );
FILL FILL_5_7 ( );
FILL FILL_5_8 ( );
FILL FILL_5_0_0 ( );
FILL FILL_5_0_1 ( );
FILL FILL_5_0_2 ( );
FILL FILL_5_1_0 ( );
FILL FILL_5_1_1 ( );
FILL FILL_5_1_2 ( );
FILL FILL_5_2_0 ( );
FILL FILL_5_2_1 ( );
FILL FILL_5_2_2 ( );
FILL FILL_5_3_0 ( );
FILL FILL_5_3_1 ( );
FILL FILL_5_3_2 ( );
FILL FILL_5_4_0 ( );
FILL FILL_5_4_1 ( );
FILL FILL_5_4_2 ( );
FILL FILL_5_5_0 ( );
FILL FILL_5_5_1 ( );
FILL FILL_5_5_2 ( );
FILL FILL_6_1 ( );
FILL FILL_6_2 ( );
FILL FILL_6_0_0 ( );
FILL FILL_6_0_1 ( );
FILL FILL_6_0_2 ( );
FILL FILL_6_1_0 ( );
FILL FILL_6_1_1 ( );
FILL FILL_6_1_2 ( );
FILL FILL_6_2_0 ( );
FILL FILL_6_2_1 ( );
FILL FILL_6_2_2 ( );
FILL FILL_6_3_0 ( );
FILL FILL_6_3_1 ( );
FILL FILL_6_3_2 ( );
FILL FILL_6_4_0 ( );
FILL FILL_6_4_1 ( );
FILL FILL_6_4_2 ( );
FILL FILL_6_5_0 ( );
FILL FILL_6_5_1 ( );
FILL FILL_6_5_2 ( );
FILL FILL_7_1 ( );
FILL FILL_7_2 ( );
FILL FILL_7_3 ( );
FILL FILL_7_4 ( );
FILL FILL_7_5 ( );
FILL FILL_7_6 ( );
FILL FILL_7_7 ( );
FILL FILL_7_0_0 ( );
FILL FILL_7_0_1 ( );
FILL FILL_7_0_2 ( );
FILL FILL_7_1_0 ( );
FILL FILL_7_1_1 ( );
FILL FILL_7_1_2 ( );
FILL FILL_7_2_0 ( );
FILL FILL_7_2_1 ( );
FILL FILL_7_2_2 ( );
FILL FILL_7_3_0 ( );
FILL FILL_7_3_1 ( );
FILL FILL_7_3_2 ( );
FILL FILL_7_4_0 ( );
FILL FILL_7_4_1 ( );
FILL FILL_7_4_2 ( );
FILL FILL_7_5_0 ( );
FILL FILL_7_5_1 ( );
FILL FILL_7_5_2 ( );
FILL FILL_8_1 ( );
FILL FILL_8_2 ( );
FILL FILL_8_0_0 ( );
FILL FILL_8_0_1 ( );
FILL FILL_8_0_2 ( );
FILL FILL_8_1_0 ( );
FILL FILL_8_1_1 ( );
FILL FILL_8_1_2 ( );
FILL FILL_8_2_0 ( );
FILL FILL_8_2_1 ( );
FILL FILL_8_2_2 ( );
FILL FILL_8_3_0 ( );
FILL FILL_8_3_1 ( );
FILL FILL_8_3_2 ( );
FILL FILL_8_4_0 ( );
FILL FILL_8_4_1 ( );
FILL FILL_8_4_2 ( );
FILL FILL_8_5_0 ( );
FILL FILL_8_5_1 ( );
FILL FILL_8_5_2 ( );
FILL FILL_9_1 ( );
FILL FILL_9_2 ( );
FILL FILL_9_3 ( );
FILL FILL_9_4 ( );
FILL FILL_9_0_0 ( );
FILL FILL_9_0_1 ( );
FILL FILL_9_0_2 ( );
FILL FILL_9_1_0 ( );
FILL FILL_9_1_1 ( );
FILL FILL_9_1_2 ( );
FILL FILL_9_2_0 ( );
FILL FILL_9_2_1 ( );
FILL FILL_9_2_2 ( );
FILL FILL_9_3_0 ( );
FILL FILL_9_3_1 ( );
FILL FILL_9_3_2 ( );
FILL FILL_9_4_0 ( );
FILL FILL_9_4_1 ( );
FILL FILL_9_4_2 ( );
FILL FILL_9_5_0 ( );
FILL FILL_9_5_1 ( );
FILL FILL_9_5_2 ( );
FILL FILL_10_1 ( );
FILL FILL_10_2 ( );
FILL FILL_10_3 ( );
FILL FILL_10_4 ( );
FILL FILL_10_5 ( );
FILL FILL_10_6 ( );
FILL FILL_10_7 ( );
FILL FILL_10_0_0 ( );
FILL FILL_10_0_1 ( );
FILL FILL_10_0_2 ( );
FILL FILL_10_1_0 ( );
FILL FILL_10_1_1 ( );
FILL FILL_10_1_2 ( );
FILL FILL_10_2_0 ( );
FILL FILL_10_2_1 ( );
FILL FILL_10_2_2 ( );
FILL FILL_10_3_0 ( );
FILL FILL_10_3_1 ( );
FILL FILL_10_3_2 ( );
FILL FILL_10_4_0 ( );
FILL FILL_10_4_1 ( );
FILL FILL_10_4_2 ( );
FILL FILL_10_5_0 ( );
FILL FILL_10_5_1 ( );
FILL FILL_10_5_2 ( );
FILL FILL_11_1 ( );
FILL FILL_11_2 ( );
FILL FILL_11_3 ( );
FILL FILL_11_4 ( );
FILL FILL_11_5 ( );
FILL FILL_11_6 ( );
FILL FILL_11_7 ( );
FILL FILL_11_0_0 ( );
FILL FILL_11_0_1 ( );
FILL FILL_11_0_2 ( );
FILL FILL_11_1_0 ( );
FILL FILL_11_1_1 ( );
FILL FILL_11_1_2 ( );
FILL FILL_11_2_0 ( );
FILL FILL_11_2_1 ( );
FILL FILL_11_2_2 ( );
FILL FILL_11_3_0 ( );
FILL FILL_11_3_1 ( );
FILL FILL_11_3_2 ( );
FILL FILL_11_4_0 ( );
FILL FILL_11_4_1 ( );
FILL FILL_11_4_2 ( );
FILL FILL_11_5_0 ( );
FILL FILL_11_5_1 ( );
FILL FILL_11_5_2 ( );
FILL FILL_12_0_0 ( );
FILL FILL_12_0_1 ( );
FILL FILL_12_0_2 ( );
FILL FILL_12_1_0 ( );
FILL FILL_12_1_1 ( );
FILL FILL_12_1_2 ( );
FILL FILL_12_2_0 ( );
FILL FILL_12_2_1 ( );
FILL FILL_12_2_2 ( );
FILL FILL_12_3_0 ( );
FILL FILL_12_3_1 ( );
FILL FILL_12_3_2 ( );
FILL FILL_12_4_0 ( );
FILL FILL_12_4_1 ( );
FILL FILL_12_4_2 ( );
FILL FILL_12_5_0 ( );
FILL FILL_12_5_1 ( );
FILL FILL_12_5_2 ( );
FILL FILL_13_1 ( );
FILL FILL_13_2 ( );
FILL FILL_13_0_0 ( );
FILL FILL_13_0_1 ( );
FILL FILL_13_0_2 ( );
FILL FILL_13_1_0 ( );
FILL FILL_13_1_1 ( );
FILL FILL_13_1_2 ( );
FILL FILL_13_2_0 ( );
FILL FILL_13_2_1 ( );
FILL FILL_13_2_2 ( );
FILL FILL_13_3_0 ( );
FILL FILL_13_3_1 ( );
FILL FILL_13_3_2 ( );
FILL FILL_13_4_0 ( );
FILL FILL_13_4_1 ( );
FILL FILL_13_4_2 ( );
FILL FILL_13_5_0 ( );
FILL FILL_13_5_1 ( );
FILL FILL_13_5_2 ( );
FILL FILL_14_1 ( );
FILL FILL_14_2 ( );
FILL FILL_14_3 ( );
FILL FILL_14_4 ( );
FILL FILL_14_5 ( );
FILL FILL_14_6 ( );
FILL FILL_14_7 ( );
FILL FILL_14_0_0 ( );
FILL FILL_14_0_1 ( );
FILL FILL_14_0_2 ( );
FILL FILL_14_1_0 ( );
FILL FILL_14_1_1 ( );
FILL FILL_14_1_2 ( );
FILL FILL_14_2_0 ( );
FILL FILL_14_2_1 ( );
FILL FILL_14_2_2 ( );
FILL FILL_14_3_0 ( );
FILL FILL_14_3_1 ( );
FILL FILL_14_3_2 ( );
FILL FILL_14_4_0 ( );
FILL FILL_14_4_1 ( );
FILL FILL_14_4_2 ( );
FILL FILL_14_5_0 ( );
FILL FILL_14_5_1 ( );
FILL FILL_14_5_2 ( );
FILL FILL_15_1 ( );
FILL FILL_15_2 ( );
FILL FILL_15_0_0 ( );
FILL FILL_15_0_1 ( );
FILL FILL_15_0_2 ( );
FILL FILL_15_1_0 ( );
FILL FILL_15_1_1 ( );
FILL FILL_15_1_2 ( );
FILL FILL_15_2_0 ( );
FILL FILL_15_2_1 ( );
FILL FILL_15_2_2 ( );
FILL FILL_15_3_0 ( );
FILL FILL_15_3_1 ( );
FILL FILL_15_3_2 ( );
FILL FILL_15_4_0 ( );
FILL FILL_15_4_1 ( );
FILL FILL_15_4_2 ( );
FILL FILL_15_5_0 ( );
FILL FILL_15_5_1 ( );
FILL FILL_15_5_2 ( );
FILL FILL_16_1 ( );
FILL FILL_16_2 ( );
FILL FILL_16_3 ( );
FILL FILL_16_4 ( );
FILL FILL_16_0_0 ( );
FILL FILL_16_0_1 ( );
FILL FILL_16_0_2 ( );
FILL FILL_16_1_0 ( );
FILL FILL_16_1_1 ( );
FILL FILL_16_1_2 ( );
FILL FILL_16_2_0 ( );
FILL FILL_16_2_1 ( );
FILL FILL_16_2_2 ( );
FILL FILL_16_3_0 ( );
FILL FILL_16_3_1 ( );
FILL FILL_16_3_2 ( );
FILL FILL_16_4_0 ( );
FILL FILL_16_4_1 ( );
FILL FILL_16_4_2 ( );
FILL FILL_16_5_0 ( );
FILL FILL_16_5_1 ( );
FILL FILL_16_5_2 ( );
FILL FILL_17_1 ( );
FILL FILL_17_2 ( );
FILL FILL_17_3 ( );
FILL FILL_17_4 ( );
FILL FILL_17_5 ( );
FILL FILL_17_6 ( );
FILL FILL_17_7 ( );
FILL FILL_17_0_0 ( );
FILL FILL_17_0_1 ( );
FILL FILL_17_0_2 ( );
FILL FILL_17_1_0 ( );
FILL FILL_17_1_1 ( );
FILL FILL_17_1_2 ( );
FILL FILL_17_2_0 ( );
FILL FILL_17_2_1 ( );
FILL FILL_17_2_2 ( );
FILL FILL_17_3_0 ( );
FILL FILL_17_3_1 ( );
FILL FILL_17_3_2 ( );
FILL FILL_17_4_0 ( );
FILL FILL_17_4_1 ( );
FILL FILL_17_4_2 ( );
FILL FILL_17_5_0 ( );
FILL FILL_17_5_1 ( );
FILL FILL_17_5_2 ( );
FILL FILL_18_0_0 ( );
FILL FILL_18_0_1 ( );
FILL FILL_18_0_2 ( );
FILL FILL_18_1_0 ( );
FILL FILL_18_1_1 ( );
FILL FILL_18_1_2 ( );
FILL FILL_18_2_0 ( );
FILL FILL_18_2_1 ( );
FILL FILL_18_2_2 ( );
FILL FILL_18_3_0 ( );
FILL FILL_18_3_1 ( );
FILL FILL_18_3_2 ( );
FILL FILL_18_4_0 ( );
FILL FILL_18_4_1 ( );
FILL FILL_18_4_2 ( );
FILL FILL_18_5_0 ( );
FILL FILL_18_5_1 ( );
FILL FILL_18_5_2 ( );
FILL FILL_19_1 ( );
FILL FILL_19_2 ( );
FILL FILL_19_3 ( );
FILL FILL_19_4 ( );
FILL FILL_19_5 ( );
FILL FILL_19_6 ( );
FILL FILL_19_7 ( );
FILL FILL_19_8 ( );
FILL FILL_19_0_0 ( );
FILL FILL_19_0_1 ( );
FILL FILL_19_0_2 ( );
FILL FILL_19_1_0 ( );
FILL FILL_19_1_1 ( );
FILL FILL_19_1_2 ( );
FILL FILL_19_2_0 ( );
FILL FILL_19_2_1 ( );
FILL FILL_19_2_2 ( );
FILL FILL_19_3_0 ( );
FILL FILL_19_3_1 ( );
FILL FILL_19_3_2 ( );
FILL FILL_19_4_0 ( );
FILL FILL_19_4_1 ( );
FILL FILL_19_4_2 ( );
FILL FILL_19_5_0 ( );
FILL FILL_19_5_1 ( );
FILL FILL_19_5_2 ( );
FILL FILL_20_1 ( );
FILL FILL_20_2 ( );
FILL FILL_20_3 ( );
FILL FILL_20_4 ( );
FILL FILL_20_5 ( );
FILL FILL_20_6 ( );
FILL FILL_20_7 ( );
FILL FILL_20_8 ( );
FILL FILL_20_9 ( );
FILL FILL_20_0_0 ( );
FILL FILL_20_0_1 ( );
FILL FILL_20_0_2 ( );
FILL FILL_20_1_0 ( );
FILL FILL_20_1_1 ( );
FILL FILL_20_1_2 ( );
FILL FILL_20_2_0 ( );
FILL FILL_20_2_1 ( );
FILL FILL_20_2_2 ( );
FILL FILL_20_3_0 ( );
FILL FILL_20_3_1 ( );
FILL FILL_20_3_2 ( );
FILL FILL_20_4_0 ( );
FILL FILL_20_4_1 ( );
FILL FILL_20_4_2 ( );
FILL FILL_20_5_0 ( );
FILL FILL_20_5_1 ( );
FILL FILL_20_5_2 ( );
FILL FILL_21_1 ( );
FILL FILL_21_2 ( );
FILL FILL_21_3 ( );
FILL FILL_21_4 ( );
FILL FILL_21_5 ( );
FILL FILL_21_6 ( );
FILL FILL_21_7 ( );
FILL FILL_21_8 ( );
FILL FILL_21_0_0 ( );
FILL FILL_21_0_1 ( );
FILL FILL_21_0_2 ( );
FILL FILL_21_1_0 ( );
FILL FILL_21_1_1 ( );
FILL FILL_21_1_2 ( );
FILL FILL_21_2_0 ( );
FILL FILL_21_2_1 ( );
FILL FILL_21_2_2 ( );
FILL FILL_21_3_0 ( );
FILL FILL_21_3_1 ( );
FILL FILL_21_3_2 ( );
FILL FILL_21_4_0 ( );
FILL FILL_21_4_1 ( );
FILL FILL_21_4_2 ( );
FILL FILL_21_5_0 ( );
FILL FILL_21_5_1 ( );
FILL FILL_21_5_2 ( );
FILL FILL_22_1 ( );
FILL FILL_22_2 ( );
FILL FILL_22_3 ( );
FILL FILL_22_4 ( );
FILL FILL_22_5 ( );
FILL FILL_22_6 ( );
FILL FILL_22_7 ( );
FILL FILL_22_8 ( );
FILL FILL_22_0_0 ( );
FILL FILL_22_0_1 ( );
FILL FILL_22_0_2 ( );
FILL FILL_22_1_0 ( );
FILL FILL_22_1_1 ( );
FILL FILL_22_1_2 ( );
FILL FILL_22_2_0 ( );
FILL FILL_22_2_1 ( );
FILL FILL_22_2_2 ( );
FILL FILL_22_3_0 ( );
FILL FILL_22_3_1 ( );
FILL FILL_22_3_2 ( );
FILL FILL_22_4_0 ( );
FILL FILL_22_4_1 ( );
FILL FILL_22_4_2 ( );
FILL FILL_22_5_0 ( );
FILL FILL_22_5_1 ( );
FILL FILL_22_5_2 ( );
FILL FILL_23_1 ( );
FILL FILL_23_2 ( );
FILL FILL_23_3 ( );
FILL FILL_23_4 ( );
FILL FILL_23_5 ( );
FILL FILL_23_0_0 ( );
FILL FILL_23_0_1 ( );
FILL FILL_23_0_2 ( );
FILL FILL_23_1_0 ( );
FILL FILL_23_1_1 ( );
FILL FILL_23_1_2 ( );
FILL FILL_23_2_0 ( );
FILL FILL_23_2_1 ( );
FILL FILL_23_2_2 ( );
FILL FILL_23_3_0 ( );
FILL FILL_23_3_1 ( );
FILL FILL_23_3_2 ( );
FILL FILL_23_4_0 ( );
FILL FILL_23_4_1 ( );
FILL FILL_23_4_2 ( );
FILL FILL_23_5_0 ( );
FILL FILL_23_5_1 ( );
FILL FILL_23_5_2 ( );
FILL FILL_24_0_0 ( );
FILL FILL_24_0_1 ( );
FILL FILL_24_0_2 ( );
FILL FILL_24_1_0 ( );
FILL FILL_24_1_1 ( );
FILL FILL_24_1_2 ( );
FILL FILL_24_2_0 ( );
FILL FILL_24_2_1 ( );
FILL FILL_24_2_2 ( );
FILL FILL_24_3_0 ( );
FILL FILL_24_3_1 ( );
FILL FILL_24_3_2 ( );
FILL FILL_24_4_0 ( );
FILL FILL_24_4_1 ( );
FILL FILL_24_4_2 ( );
FILL FILL_24_5_0 ( );
FILL FILL_24_5_1 ( );
FILL FILL_24_5_2 ( );
FILL FILL_25_1 ( );
FILL FILL_25_2 ( );
FILL FILL_25_3 ( );
FILL FILL_25_4 ( );
FILL FILL_25_5 ( );
FILL FILL_25_0_0 ( );
FILL FILL_25_0_1 ( );
FILL FILL_25_0_2 ( );
FILL FILL_25_1_0 ( );
FILL FILL_25_1_1 ( );
FILL FILL_25_1_2 ( );
FILL FILL_25_2_0 ( );
FILL FILL_25_2_1 ( );
FILL FILL_25_2_2 ( );
FILL FILL_25_3_0 ( );
FILL FILL_25_3_1 ( );
FILL FILL_25_3_2 ( );
FILL FILL_25_4_0 ( );
FILL FILL_25_4_1 ( );
FILL FILL_25_4_2 ( );
FILL FILL_25_5_0 ( );
FILL FILL_25_5_1 ( );
FILL FILL_25_5_2 ( );
FILL FILL_26_1 ( );
FILL FILL_26_2 ( );
FILL FILL_26_3 ( );
FILL FILL_26_4 ( );
FILL FILL_26_5 ( );
FILL FILL_26_6 ( );
FILL FILL_26_0_0 ( );
FILL FILL_26_0_1 ( );
FILL FILL_26_0_2 ( );
FILL FILL_26_1_0 ( );
FILL FILL_26_1_1 ( );
FILL FILL_26_1_2 ( );
FILL FILL_26_2_0 ( );
FILL FILL_26_2_1 ( );
FILL FILL_26_2_2 ( );
FILL FILL_26_3_0 ( );
FILL FILL_26_3_1 ( );
FILL FILL_26_3_2 ( );
FILL FILL_26_4_0 ( );
FILL FILL_26_4_1 ( );
FILL FILL_26_4_2 ( );
FILL FILL_26_5_0 ( );
FILL FILL_26_5_1 ( );
FILL FILL_26_5_2 ( );
FILL FILL_27_1 ( );
FILL FILL_27_0_0 ( );
FILL FILL_27_0_1 ( );
FILL FILL_27_0_2 ( );
FILL FILL_27_1_0 ( );
FILL FILL_27_1_1 ( );
FILL FILL_27_1_2 ( );
FILL FILL_27_2_0 ( );
FILL FILL_27_2_1 ( );
FILL FILL_27_2_2 ( );
FILL FILL_27_3_0 ( );
FILL FILL_27_3_1 ( );
FILL FILL_27_3_2 ( );
FILL FILL_27_4_0 ( );
FILL FILL_27_4_1 ( );
FILL FILL_27_4_2 ( );
FILL FILL_27_5_0 ( );
FILL FILL_27_5_1 ( );
FILL FILL_27_5_2 ( );
FILL FILL_28_1 ( );
FILL FILL_28_0_0 ( );
FILL FILL_28_0_1 ( );
FILL FILL_28_0_2 ( );
FILL FILL_28_1_0 ( );
FILL FILL_28_1_1 ( );
FILL FILL_28_1_2 ( );
FILL FILL_28_2_0 ( );
FILL FILL_28_2_1 ( );
FILL FILL_28_2_2 ( );
FILL FILL_28_3_0 ( );
FILL FILL_28_3_1 ( );
FILL FILL_28_3_2 ( );
FILL FILL_28_4_0 ( );
FILL FILL_28_4_1 ( );
FILL FILL_28_4_2 ( );
FILL FILL_28_5_0 ( );
FILL FILL_28_5_1 ( );
FILL FILL_28_5_2 ( );
FILL FILL_29_1 ( );
FILL FILL_29_2 ( );
FILL FILL_29_3 ( );
FILL FILL_29_4 ( );
FILL FILL_29_5 ( );
FILL FILL_29_0_0 ( );
FILL FILL_29_0_1 ( );
FILL FILL_29_0_2 ( );
FILL FILL_29_1_0 ( );
FILL FILL_29_1_1 ( );
FILL FILL_29_1_2 ( );
FILL FILL_29_2_0 ( );
FILL FILL_29_2_1 ( );
FILL FILL_29_2_2 ( );
FILL FILL_29_3_0 ( );
FILL FILL_29_3_1 ( );
FILL FILL_29_3_2 ( );
FILL FILL_29_4_0 ( );
FILL FILL_29_4_1 ( );
FILL FILL_29_4_2 ( );
FILL FILL_29_5_0 ( );
FILL FILL_29_5_1 ( );
FILL FILL_29_5_2 ( );
FILL FILL_30_1 ( );
FILL FILL_30_2 ( );
FILL FILL_30_3 ( );
FILL FILL_30_0_0 ( );
FILL FILL_30_0_1 ( );
FILL FILL_30_0_2 ( );
FILL FILL_30_1_0 ( );
FILL FILL_30_1_1 ( );
FILL FILL_30_1_2 ( );
FILL FILL_30_2_0 ( );
FILL FILL_30_2_1 ( );
FILL FILL_30_2_2 ( );
FILL FILL_30_3_0 ( );
FILL FILL_30_3_1 ( );
FILL FILL_30_3_2 ( );
FILL FILL_30_4_0 ( );
FILL FILL_30_4_1 ( );
FILL FILL_30_4_2 ( );
FILL FILL_30_5_0 ( );
FILL FILL_30_5_1 ( );
FILL FILL_30_5_2 ( );
FILL FILL_31_1 ( );
FILL FILL_31_0_0 ( );
FILL FILL_31_0_1 ( );
FILL FILL_31_0_2 ( );
FILL FILL_31_1_0 ( );
FILL FILL_31_1_1 ( );
FILL FILL_31_1_2 ( );
FILL FILL_31_2_0 ( );
FILL FILL_31_2_1 ( );
FILL FILL_31_2_2 ( );
FILL FILL_31_3_0 ( );
FILL FILL_31_3_1 ( );
FILL FILL_31_3_2 ( );
FILL FILL_31_4_0 ( );
FILL FILL_31_4_1 ( );
FILL FILL_31_4_2 ( );
FILL FILL_31_5_0 ( );
FILL FILL_31_5_1 ( );
FILL FILL_31_5_2 ( );
FILL FILL_32_1 ( );
FILL FILL_32_2 ( );
FILL FILL_32_0_0 ( );
FILL FILL_32_0_1 ( );
FILL FILL_32_0_2 ( );
FILL FILL_32_1_0 ( );
FILL FILL_32_1_1 ( );
FILL FILL_32_1_2 ( );
FILL FILL_32_2_0 ( );
FILL FILL_32_2_1 ( );
FILL FILL_32_2_2 ( );
FILL FILL_32_3_0 ( );
FILL FILL_32_3_1 ( );
FILL FILL_32_3_2 ( );
FILL FILL_32_4_0 ( );
FILL FILL_32_4_1 ( );
FILL FILL_32_4_2 ( );
FILL FILL_32_5_0 ( );
FILL FILL_32_5_1 ( );
FILL FILL_32_5_2 ( );
FILL FILL_33_1 ( );
FILL FILL_33_2 ( );
FILL FILL_33_3 ( );
FILL FILL_33_4 ( );
FILL FILL_33_5 ( );
FILL FILL_33_6 ( );
FILL FILL_33_7 ( );
FILL FILL_33_8 ( );
FILL FILL_33_0_0 ( );
FILL FILL_33_0_1 ( );
FILL FILL_33_0_2 ( );
FILL FILL_33_1_0 ( );
FILL FILL_33_1_1 ( );
FILL FILL_33_1_2 ( );
FILL FILL_33_2_0 ( );
FILL FILL_33_2_1 ( );
FILL FILL_33_2_2 ( );
FILL FILL_33_3_0 ( );
FILL FILL_33_3_1 ( );
FILL FILL_33_3_2 ( );
FILL FILL_33_4_0 ( );
FILL FILL_33_4_1 ( );
FILL FILL_33_4_2 ( );
FILL FILL_33_5_0 ( );
FILL FILL_33_5_1 ( );
FILL FILL_33_5_2 ( );
FILL FILL_34_1 ( );
FILL FILL_34_2 ( );
FILL FILL_34_3 ( );
FILL FILL_34_4 ( );
FILL FILL_34_5 ( );
FILL FILL_34_6 ( );
FILL FILL_34_7 ( );
FILL FILL_34_8 ( );
FILL FILL_34_9 ( );
FILL FILL_34_0_0 ( );
FILL FILL_34_0_1 ( );
FILL FILL_34_0_2 ( );
FILL FILL_34_1_0 ( );
FILL FILL_34_1_1 ( );
FILL FILL_34_1_2 ( );
FILL FILL_34_2_0 ( );
FILL FILL_34_2_1 ( );
FILL FILL_34_2_2 ( );
FILL FILL_34_3_0 ( );
FILL FILL_34_3_1 ( );
FILL FILL_34_3_2 ( );
FILL FILL_34_4_0 ( );
FILL FILL_34_4_1 ( );
FILL FILL_34_4_2 ( );
FILL FILL_34_5_0 ( );
FILL FILL_34_5_1 ( );
FILL FILL_34_5_2 ( );
FILL FILL_35_1 ( );
FILL FILL_35_2 ( );
FILL FILL_35_3 ( );
FILL FILL_35_4 ( );
FILL FILL_35_5 ( );
FILL FILL_35_6 ( );
FILL FILL_35_7 ( );
FILL FILL_35_8 ( );
FILL FILL_35_0_0 ( );
FILL FILL_35_0_1 ( );
FILL FILL_35_0_2 ( );
FILL FILL_35_1_0 ( );
FILL FILL_35_1_1 ( );
FILL FILL_35_1_2 ( );
FILL FILL_35_2_0 ( );
FILL FILL_35_2_1 ( );
FILL FILL_35_2_2 ( );
FILL FILL_35_3_0 ( );
FILL FILL_35_3_1 ( );
FILL FILL_35_3_2 ( );
FILL FILL_35_4_0 ( );
FILL FILL_35_4_1 ( );
FILL FILL_35_4_2 ( );
FILL FILL_35_5_0 ( );
FILL FILL_35_5_1 ( );
FILL FILL_35_5_2 ( );
FILL FILL_36_1 ( );
FILL FILL_36_2 ( );
FILL FILL_36_3 ( );
FILL FILL_36_0_0 ( );
FILL FILL_36_0_1 ( );
FILL FILL_36_0_2 ( );
FILL FILL_36_1_0 ( );
FILL FILL_36_1_1 ( );
FILL FILL_36_1_2 ( );
FILL FILL_36_2_0 ( );
FILL FILL_36_2_1 ( );
FILL FILL_36_2_2 ( );
FILL FILL_36_3_0 ( );
FILL FILL_36_3_1 ( );
FILL FILL_36_3_2 ( );
FILL FILL_36_4_0 ( );
FILL FILL_36_4_1 ( );
FILL FILL_36_4_2 ( );
FILL FILL_36_5_0 ( );
FILL FILL_36_5_1 ( );
FILL FILL_36_5_2 ( );
FILL FILL_37_0_0 ( );
FILL FILL_37_0_1 ( );
FILL FILL_37_0_2 ( );
FILL FILL_37_1_0 ( );
FILL FILL_37_1_1 ( );
FILL FILL_37_1_2 ( );
FILL FILL_37_2_0 ( );
FILL FILL_37_2_1 ( );
FILL FILL_37_2_2 ( );
FILL FILL_37_3_0 ( );
FILL FILL_37_3_1 ( );
FILL FILL_37_3_2 ( );
FILL FILL_37_4_0 ( );
FILL FILL_37_4_1 ( );
FILL FILL_37_4_2 ( );
FILL FILL_37_5_0 ( );
FILL FILL_37_5_1 ( );
FILL FILL_37_5_2 ( );
FILL FILL_38_1 ( );
FILL FILL_38_2 ( );
FILL FILL_38_3 ( );
FILL FILL_38_4 ( );
FILL FILL_38_5 ( );
FILL FILL_38_6 ( );
FILL FILL_38_7 ( );
FILL FILL_38_8 ( );
FILL FILL_38_0_0 ( );
FILL FILL_38_0_1 ( );
FILL FILL_38_0_2 ( );
FILL FILL_38_1_0 ( );
FILL FILL_38_1_1 ( );
FILL FILL_38_1_2 ( );
FILL FILL_38_2_0 ( );
FILL FILL_38_2_1 ( );
FILL FILL_38_2_2 ( );
FILL FILL_38_3_0 ( );
FILL FILL_38_3_1 ( );
FILL FILL_38_3_2 ( );
FILL FILL_38_4_0 ( );
FILL FILL_38_4_1 ( );
FILL FILL_38_4_2 ( );
FILL FILL_38_5_0 ( );
FILL FILL_38_5_1 ( );
FILL FILL_38_5_2 ( );
FILL FILL_39_1 ( );
FILL FILL_39_2 ( );
FILL FILL_39_3 ( );
FILL FILL_39_4 ( );
FILL FILL_39_5 ( );
FILL FILL_39_6 ( );
FILL FILL_39_7 ( );
FILL FILL_39_0_0 ( );
FILL FILL_39_0_1 ( );
FILL FILL_39_0_2 ( );
FILL FILL_39_1_0 ( );
FILL FILL_39_1_1 ( );
FILL FILL_39_1_2 ( );
FILL FILL_39_2_0 ( );
FILL FILL_39_2_1 ( );
FILL FILL_39_2_2 ( );
FILL FILL_39_3_0 ( );
FILL FILL_39_3_1 ( );
FILL FILL_39_3_2 ( );
FILL FILL_39_4_0 ( );
FILL FILL_39_4_1 ( );
FILL FILL_39_4_2 ( );
FILL FILL_39_5_0 ( );
FILL FILL_39_5_1 ( );
FILL FILL_39_5_2 ( );
FILL FILL_40_1 ( );
FILL FILL_40_2 ( );
FILL FILL_40_3 ( );
FILL FILL_40_4 ( );
FILL FILL_40_0_0 ( );
FILL FILL_40_0_1 ( );
FILL FILL_40_0_2 ( );
FILL FILL_40_1_0 ( );
FILL FILL_40_1_1 ( );
FILL FILL_40_1_2 ( );
FILL FILL_40_2_0 ( );
FILL FILL_40_2_1 ( );
FILL FILL_40_2_2 ( );
FILL FILL_40_3_0 ( );
FILL FILL_40_3_1 ( );
FILL FILL_40_3_2 ( );
FILL FILL_40_4_0 ( );
FILL FILL_40_4_1 ( );
FILL FILL_40_4_2 ( );
FILL FILL_40_5_0 ( );
FILL FILL_40_5_1 ( );
FILL FILL_40_5_2 ( );
FILL FILL_41_1 ( );
FILL FILL_41_2 ( );
FILL FILL_41_3 ( );
FILL FILL_41_4 ( );
FILL FILL_41_5 ( );
FILL FILL_41_6 ( );
FILL FILL_41_0_0 ( );
FILL FILL_41_0_1 ( );
FILL FILL_41_0_2 ( );
FILL FILL_41_1_0 ( );
FILL FILL_41_1_1 ( );
FILL FILL_41_1_2 ( );
FILL FILL_41_2_0 ( );
FILL FILL_41_2_1 ( );
FILL FILL_41_2_2 ( );
FILL FILL_41_3_0 ( );
FILL FILL_41_3_1 ( );
FILL FILL_41_3_2 ( );
FILL FILL_41_4_0 ( );
FILL FILL_41_4_1 ( );
FILL FILL_41_4_2 ( );
FILL FILL_41_5_0 ( );
FILL FILL_41_5_1 ( );
FILL FILL_41_5_2 ( );
FILL FILL_42_1 ( );
FILL FILL_42_2 ( );
FILL FILL_42_3 ( );
FILL FILL_42_4 ( );
FILL FILL_42_5 ( );
FILL FILL_42_0_0 ( );
FILL FILL_42_0_1 ( );
FILL FILL_42_0_2 ( );
FILL FILL_42_1_0 ( );
FILL FILL_42_1_1 ( );
FILL FILL_42_1_2 ( );
FILL FILL_42_2_0 ( );
FILL FILL_42_2_1 ( );
FILL FILL_42_2_2 ( );
FILL FILL_42_3_0 ( );
FILL FILL_42_3_1 ( );
FILL FILL_42_3_2 ( );
FILL FILL_42_4_0 ( );
FILL FILL_42_4_1 ( );
FILL FILL_42_4_2 ( );
FILL FILL_42_5_0 ( );
FILL FILL_42_5_1 ( );
FILL FILL_42_5_2 ( );
FILL FILL_43_1 ( );
FILL FILL_43_2 ( );
FILL FILL_43_3 ( );
FILL FILL_43_4 ( );
FILL FILL_43_5 ( );
FILL FILL_43_6 ( );
FILL FILL_43_7 ( );
FILL FILL_43_8 ( );
FILL FILL_43_0_0 ( );
FILL FILL_43_0_1 ( );
FILL FILL_43_0_2 ( );
FILL FILL_43_1_0 ( );
FILL FILL_43_1_1 ( );
FILL FILL_43_1_2 ( );
FILL FILL_43_2_0 ( );
FILL FILL_43_2_1 ( );
FILL FILL_43_2_2 ( );
FILL FILL_43_3_0 ( );
FILL FILL_43_3_1 ( );
FILL FILL_43_3_2 ( );
FILL FILL_43_4_0 ( );
FILL FILL_43_4_1 ( );
FILL FILL_43_4_2 ( );
FILL FILL_43_5_0 ( );
FILL FILL_43_5_1 ( );
FILL FILL_43_5_2 ( );
FILL FILL_44_1 ( );
FILL FILL_44_2 ( );
FILL FILL_44_3 ( );
FILL FILL_44_4 ( );
FILL FILL_44_5 ( );
FILL FILL_44_0_0 ( );
FILL FILL_44_0_1 ( );
FILL FILL_44_0_2 ( );
FILL FILL_44_1_0 ( );
FILL FILL_44_1_1 ( );
FILL FILL_44_1_2 ( );
FILL FILL_44_2_0 ( );
FILL FILL_44_2_1 ( );
FILL FILL_44_2_2 ( );
FILL FILL_44_3_0 ( );
FILL FILL_44_3_1 ( );
FILL FILL_44_3_2 ( );
FILL FILL_44_4_0 ( );
FILL FILL_44_4_1 ( );
FILL FILL_44_4_2 ( );
FILL FILL_44_5_0 ( );
FILL FILL_44_5_1 ( );
FILL FILL_44_5_2 ( );
FILL FILL_45_1 ( );
FILL FILL_45_2 ( );
FILL FILL_45_3 ( );
FILL FILL_45_4 ( );
FILL FILL_45_5 ( );
FILL FILL_45_6 ( );
FILL FILL_45_7 ( );
FILL FILL_45_0_0 ( );
FILL FILL_45_0_1 ( );
FILL FILL_45_0_2 ( );
FILL FILL_45_1_0 ( );
FILL FILL_45_1_1 ( );
FILL FILL_45_1_2 ( );
FILL FILL_45_2_0 ( );
FILL FILL_45_2_1 ( );
FILL FILL_45_2_2 ( );
FILL FILL_45_3_0 ( );
FILL FILL_45_3_1 ( );
FILL FILL_45_3_2 ( );
FILL FILL_45_4_0 ( );
FILL FILL_45_4_1 ( );
FILL FILL_45_4_2 ( );
FILL FILL_45_5_0 ( );
FILL FILL_45_5_1 ( );
FILL FILL_45_5_2 ( );
FILL FILL_46_1 ( );
FILL FILL_46_2 ( );
FILL FILL_46_3 ( );
FILL FILL_46_4 ( );
FILL FILL_46_0_0 ( );
FILL FILL_46_0_1 ( );
FILL FILL_46_0_2 ( );
FILL FILL_46_1_0 ( );
FILL FILL_46_1_1 ( );
FILL FILL_46_1_2 ( );
FILL FILL_46_2_0 ( );
FILL FILL_46_2_1 ( );
FILL FILL_46_2_2 ( );
FILL FILL_46_3_0 ( );
FILL FILL_46_3_1 ( );
FILL FILL_46_3_2 ( );
FILL FILL_46_4_0 ( );
FILL FILL_46_4_1 ( );
FILL FILL_46_4_2 ( );
FILL FILL_46_5_0 ( );
FILL FILL_46_5_1 ( );
FILL FILL_46_5_2 ( );
FILL FILL_47_1 ( );
FILL FILL_47_2 ( );
FILL FILL_47_0_0 ( );
FILL FILL_47_0_1 ( );
FILL FILL_47_0_2 ( );
FILL FILL_47_1_0 ( );
FILL FILL_47_1_1 ( );
FILL FILL_47_1_2 ( );
FILL FILL_47_2_0 ( );
FILL FILL_47_2_1 ( );
FILL FILL_47_2_2 ( );
FILL FILL_47_3_0 ( );
FILL FILL_47_3_1 ( );
FILL FILL_47_3_2 ( );
FILL FILL_47_4_0 ( );
FILL FILL_47_4_1 ( );
FILL FILL_47_4_2 ( );
FILL FILL_47_5_0 ( );
FILL FILL_47_5_1 ( );
FILL FILL_47_5_2 ( );
FILL FILL_48_1 ( );
FILL FILL_48_2 ( );
FILL FILL_48_3 ( );
FILL FILL_48_4 ( );
FILL FILL_48_5 ( );
FILL FILL_48_6 ( );
FILL FILL_48_7 ( );
FILL FILL_48_8 ( );
FILL FILL_48_9 ( );
FILL FILL_48_0_0 ( );
FILL FILL_48_0_1 ( );
FILL FILL_48_0_2 ( );
FILL FILL_48_1_0 ( );
FILL FILL_48_1_1 ( );
FILL FILL_48_1_2 ( );
FILL FILL_48_2_0 ( );
FILL FILL_48_2_1 ( );
FILL FILL_48_2_2 ( );
FILL FILL_48_3_0 ( );
FILL FILL_48_3_1 ( );
FILL FILL_48_3_2 ( );
FILL FILL_48_4_0 ( );
FILL FILL_48_4_1 ( );
FILL FILL_48_4_2 ( );
FILL FILL_48_5_0 ( );
FILL FILL_48_5_1 ( );
FILL FILL_48_5_2 ( );
endmodule
